magic
tech sky130A
magscale 1 2
timestamp 1608446478
<< metal1 >>
rect 58618 700952 58624 701004
rect 58676 700992 58682 701004
rect 137830 700992 137836 701004
rect 58676 700964 137836 700992
rect 58676 700952 58682 700964
rect 137830 700952 137836 700964
rect 137888 700952 137894 701004
rect 137922 700952 137928 701004
rect 137980 700992 137986 701004
rect 235166 700992 235172 701004
rect 137980 700964 235172 700992
rect 137980 700952 137986 700964
rect 235166 700952 235172 700964
rect 235224 700952 235230 701004
rect 58710 700884 58716 700936
rect 58768 700924 58774 700936
rect 202782 700924 202788 700936
rect 58768 700896 202788 700924
rect 58768 700884 58774 700896
rect 202782 700884 202788 700896
rect 202840 700884 202846 700936
rect 57790 700816 57796 700868
rect 57848 700856 57854 700868
rect 218974 700856 218980 700868
rect 57848 700828 218980 700856
rect 57848 700816 57854 700828
rect 218974 700816 218980 700828
rect 219032 700816 219038 700868
rect 58894 700748 58900 700800
rect 58952 700788 58958 700800
rect 267642 700788 267648 700800
rect 58952 700760 267648 700788
rect 58952 700748 58958 700760
rect 267642 700748 267648 700760
rect 267700 700748 267706 700800
rect 58802 700680 58808 700732
rect 58860 700720 58866 700732
rect 283834 700720 283840 700732
rect 58860 700692 283840 700720
rect 58860 700680 58866 700692
rect 283834 700680 283840 700692
rect 283892 700680 283898 700732
rect 58986 700612 58992 700664
rect 59044 700652 59050 700664
rect 332502 700652 332508 700664
rect 59044 700624 332508 700652
rect 59044 700612 59050 700624
rect 332502 700612 332508 700624
rect 332560 700612 332566 700664
rect 57882 700544 57888 700596
rect 57940 700584 57946 700596
rect 348786 700584 348792 700596
rect 57940 700556 348792 700584
rect 57940 700544 57946 700556
rect 348786 700544 348792 700556
rect 348844 700544 348850 700596
rect 59170 700476 59176 700528
rect 59228 700516 59234 700528
rect 397454 700516 397460 700528
rect 59228 700488 397460 700516
rect 59228 700476 59234 700488
rect 397454 700476 397460 700488
rect 397512 700476 397518 700528
rect 59078 700408 59084 700460
rect 59136 700448 59142 700460
rect 413646 700448 413652 700460
rect 59136 700420 413652 700448
rect 59136 700408 59142 700420
rect 413646 700408 413652 700420
rect 413704 700408 413710 700460
rect 59262 700340 59268 700392
rect 59320 700380 59326 700392
rect 478506 700380 478512 700392
rect 59320 700352 478512 700380
rect 59320 700340 59326 700352
rect 478506 700340 478512 700352
rect 478564 700340 478570 700392
rect 59354 700272 59360 700324
rect 59412 700312 59418 700324
rect 527174 700312 527180 700324
rect 59412 700284 527180 700312
rect 59412 700272 59418 700284
rect 527174 700272 527180 700284
rect 527232 700272 527238 700324
rect 58526 700204 58532 700256
rect 58584 700244 58590 700256
rect 154114 700244 154120 700256
rect 58584 700216 154120 700244
rect 58584 700204 58590 700216
rect 154114 700204 154120 700216
rect 154172 700204 154178 700256
rect 58342 700136 58348 700188
rect 58400 700176 58406 700188
rect 89162 700176 89168 700188
rect 58400 700148 89168 700176
rect 58400 700136 58406 700148
rect 89162 700136 89168 700148
rect 89220 700136 89226 700188
rect 58434 700068 58440 700120
rect 58492 700108 58498 700120
rect 72970 700108 72976 700120
rect 58492 700080 72976 700108
rect 58492 700068 58498 700080
rect 72970 700068 72976 700080
rect 73028 700068 73034 700120
rect 40494 699932 40500 699984
rect 40552 699972 40558 699984
rect 42058 699972 42064 699984
rect 40552 699944 42064 699972
rect 40552 699932 40558 699944
rect 42058 699932 42064 699944
rect 42116 699932 42122 699984
rect 8110 699660 8116 699712
rect 8168 699700 8174 699712
rect 10318 699700 10324 699712
rect 8168 699672 10324 699700
rect 8168 699660 8174 699672
rect 10318 699660 10324 699672
rect 10376 699660 10382 699712
rect 24302 699660 24308 699712
rect 24360 699700 24366 699712
rect 24762 699700 24768 699712
rect 24360 699672 24768 699700
rect 24360 699660 24366 699672
rect 24762 699660 24768 699672
rect 24820 699660 24826 699712
rect 137278 699660 137284 699712
rect 137336 699700 137342 699712
rect 137922 699700 137928 699712
rect 137336 699672 137928 699700
rect 137336 699660 137342 699672
rect 137922 699660 137928 699672
rect 137980 699660 137986 699712
rect 104986 698232 104992 698284
rect 105044 698272 105050 698284
rect 105538 698272 105544 698284
rect 105044 698244 105544 698272
rect 105044 698232 105050 698244
rect 105538 698232 105544 698244
rect 105596 698232 105602 698284
rect 364426 698232 364432 698284
rect 364484 698272 364490 698284
rect 365070 698272 365076 698284
rect 364484 698244 365076 698272
rect 364484 698232 364490 698244
rect 365070 698232 365076 698244
rect 365128 698232 365134 698284
rect 560294 697280 560300 697332
rect 560352 697320 560358 697332
rect 565170 697320 565176 697332
rect 560352 697292 565176 697320
rect 560352 697280 560358 697292
rect 565170 697280 565176 697292
rect 565228 697280 565234 697332
rect 540974 697144 540980 697196
rect 541032 697184 541038 697196
rect 548610 697184 548616 697196
rect 541032 697156 548616 697184
rect 541032 697144 541038 697156
rect 548610 697144 548616 697156
rect 548668 697144 548674 697196
rect 70302 697076 70308 697128
rect 70360 697116 70366 697128
rect 77202 697116 77208 697128
rect 70360 697088 77208 697116
rect 70360 697076 70366 697088
rect 77202 697076 77208 697088
rect 77260 697076 77266 697128
rect 89622 697076 89628 697128
rect 89680 697116 89686 697128
rect 96522 697116 96528 697128
rect 89680 697088 96528 697116
rect 89680 697076 89686 697088
rect 96522 697076 96528 697088
rect 96580 697076 96586 697128
rect 108942 697076 108948 697128
rect 109000 697116 109006 697128
rect 115842 697116 115848 697128
rect 109000 697088 115848 697116
rect 109000 697076 109006 697088
rect 115842 697076 115848 697088
rect 115900 697076 115906 697128
rect 128262 697076 128268 697128
rect 128320 697116 128326 697128
rect 135162 697116 135168 697128
rect 128320 697088 135168 697116
rect 128320 697076 128326 697088
rect 135162 697076 135168 697088
rect 135220 697076 135226 697128
rect 147582 697076 147588 697128
rect 147640 697116 147646 697128
rect 154482 697116 154488 697128
rect 147640 697088 154488 697116
rect 147640 697076 147646 697088
rect 154482 697076 154488 697088
rect 154540 697076 154546 697128
rect 166902 697076 166908 697128
rect 166960 697116 166966 697128
rect 173802 697116 173808 697128
rect 166960 697088 173808 697116
rect 166960 697076 166966 697088
rect 173802 697076 173808 697088
rect 173860 697076 173866 697128
rect 186222 697076 186228 697128
rect 186280 697116 186286 697128
rect 193122 697116 193128 697128
rect 186280 697088 193128 697116
rect 186280 697076 186286 697088
rect 193122 697076 193128 697088
rect 193180 697076 193186 697128
rect 205542 697076 205548 697128
rect 205600 697116 205606 697128
rect 212442 697116 212448 697128
rect 205600 697088 212448 697116
rect 205600 697076 205606 697088
rect 212442 697076 212448 697088
rect 212500 697076 212506 697128
rect 224862 697076 224868 697128
rect 224920 697116 224926 697128
rect 231762 697116 231768 697128
rect 224920 697088 231768 697116
rect 224920 697076 224926 697088
rect 231762 697076 231768 697088
rect 231820 697076 231826 697128
rect 244182 697076 244188 697128
rect 244240 697116 244246 697128
rect 251082 697116 251088 697128
rect 244240 697088 251088 697116
rect 244240 697076 244246 697088
rect 251082 697076 251088 697088
rect 251140 697076 251146 697128
rect 263502 697076 263508 697128
rect 263560 697116 263566 697128
rect 270402 697116 270408 697128
rect 263560 697088 270408 697116
rect 263560 697076 263566 697088
rect 270402 697076 270408 697088
rect 270460 697076 270466 697128
rect 282822 697076 282828 697128
rect 282880 697116 282886 697128
rect 289722 697116 289728 697128
rect 282880 697088 289728 697116
rect 282880 697076 282886 697088
rect 289722 697076 289728 697088
rect 289780 697076 289786 697128
rect 302142 697076 302148 697128
rect 302200 697116 302206 697128
rect 309042 697116 309048 697128
rect 302200 697088 309048 697116
rect 302200 697076 302206 697088
rect 309042 697076 309048 697088
rect 309100 697076 309106 697128
rect 321462 697076 321468 697128
rect 321520 697116 321526 697128
rect 328362 697116 328368 697128
rect 321520 697088 328368 697116
rect 321520 697076 321526 697088
rect 328362 697076 328368 697088
rect 328420 697076 328426 697128
rect 170122 695444 170128 695496
rect 170180 695484 170186 695496
rect 170306 695484 170312 695496
rect 170180 695456 170312 695484
rect 170180 695444 170186 695456
rect 170306 695444 170312 695456
rect 170364 695444 170370 695496
rect 429194 692792 429200 692844
rect 429252 692832 429258 692844
rect 429930 692832 429936 692844
rect 429252 692804 429936 692832
rect 429252 692792 429258 692804
rect 429930 692792 429936 692804
rect 429988 692792 429994 692844
rect 494054 692792 494060 692844
rect 494112 692832 494118 692844
rect 494882 692832 494888 692844
rect 494112 692804 494888 692832
rect 494112 692792 494118 692804
rect 494882 692792 494888 692804
rect 494940 692792 494946 692844
rect 173894 686264 173900 686316
rect 173952 686304 173958 686316
rect 178770 686304 178776 686316
rect 173952 686276 178776 686304
rect 173952 686264 173958 686276
rect 178770 686264 178776 686276
rect 178828 686264 178834 686316
rect 367094 686264 367100 686316
rect 367152 686304 367158 686316
rect 371970 686304 371976 686316
rect 367152 686276 371976 686304
rect 367152 686264 367158 686276
rect 371970 686264 371976 686276
rect 372028 686264 372034 686316
rect 560294 686264 560300 686316
rect 560352 686304 560358 686316
rect 565170 686304 565176 686316
rect 560352 686276 565176 686304
rect 560352 686264 560358 686276
rect 565170 686264 565176 686276
rect 565228 686264 565234 686316
rect 154574 686128 154580 686180
rect 154632 686168 154638 686180
rect 162210 686168 162216 686180
rect 154632 686140 162216 686168
rect 154632 686128 154638 686140
rect 162210 686128 162216 686140
rect 162268 686128 162274 686180
rect 289814 686128 289820 686180
rect 289872 686168 289878 686180
rect 294506 686168 294512 686180
rect 289872 686140 294512 686168
rect 289872 686128 289878 686140
rect 294506 686128 294512 686140
rect 294564 686128 294570 686180
rect 347774 686128 347780 686180
rect 347832 686168 347838 686180
rect 355410 686168 355416 686180
rect 347832 686140 355416 686168
rect 347832 686128 347838 686140
rect 355410 686128 355416 686140
rect 355468 686128 355474 686180
rect 540974 686128 540980 686180
rect 541032 686168 541038 686180
rect 548610 686168 548616 686180
rect 541032 686140 548616 686168
rect 541032 686128 541038 686140
rect 548610 686128 548616 686140
rect 548668 686128 548674 686180
rect 169846 685924 169852 685976
rect 169904 685964 169910 685976
rect 170122 685964 170128 685976
rect 169904 685936 170128 685964
rect 169904 685924 169910 685936
rect 170122 685924 170128 685936
rect 170180 685924 170186 685976
rect 299566 685856 299572 685908
rect 299624 685896 299630 685908
rect 300118 685896 300124 685908
rect 299624 685868 300124 685896
rect 299624 685856 299630 685868
rect 300118 685856 300124 685868
rect 300176 685856 300182 685908
rect 559006 684496 559012 684548
rect 559064 684536 559070 684548
rect 559650 684536 559656 684548
rect 559064 684508 559656 684536
rect 559064 684496 559070 684508
rect 559650 684496 559656 684508
rect 559708 684496 559714 684548
rect 169846 684428 169852 684480
rect 169904 684468 169910 684480
rect 170214 684468 170220 684480
rect 169904 684440 170220 684468
rect 169904 684428 169910 684440
rect 170214 684428 170220 684440
rect 170272 684428 170278 684480
rect 299566 684428 299572 684480
rect 299624 684468 299630 684480
rect 299658 684468 299664 684480
rect 299624 684440 299664 684468
rect 299624 684428 299630 684440
rect 299658 684428 299664 684440
rect 299716 684428 299722 684480
rect 299658 678988 299664 679040
rect 299716 678988 299722 679040
rect 299676 678904 299704 678988
rect 299658 678852 299664 678904
rect 299716 678852 299722 678904
rect 559006 674840 559012 674892
rect 559064 674880 559070 674892
rect 559374 674880 559380 674892
rect 559064 674852 559380 674880
rect 559064 674840 559070 674852
rect 559374 674840 559380 674852
rect 559432 674840 559438 674892
rect 173894 673888 173900 673940
rect 173952 673928 173958 673940
rect 178770 673928 178776 673940
rect 173952 673900 178776 673928
rect 173952 673888 173958 673900
rect 178770 673888 178776 673900
rect 178828 673888 178834 673940
rect 367094 673888 367100 673940
rect 367152 673928 367158 673940
rect 371970 673928 371976 673940
rect 367152 673900 371976 673928
rect 367152 673888 367158 673900
rect 371970 673888 371976 673900
rect 372028 673888 372034 673940
rect 560294 673888 560300 673940
rect 560352 673928 560358 673940
rect 565170 673928 565176 673940
rect 560352 673900 565176 673928
rect 560352 673888 560358 673900
rect 565170 673888 565176 673900
rect 565228 673888 565234 673940
rect 154574 673752 154580 673804
rect 154632 673792 154638 673804
rect 162210 673792 162216 673804
rect 154632 673764 162216 673792
rect 154632 673752 154638 673764
rect 162210 673752 162216 673764
rect 162268 673752 162274 673804
rect 289814 673752 289820 673804
rect 289872 673792 289878 673804
rect 292666 673792 292672 673804
rect 289872 673764 292672 673792
rect 289872 673752 289878 673764
rect 292666 673752 292672 673764
rect 292724 673752 292730 673804
rect 347774 673752 347780 673804
rect 347832 673792 347838 673804
rect 355410 673792 355416 673804
rect 347832 673764 355416 673792
rect 347832 673752 347838 673764
rect 355410 673752 355416 673764
rect 355468 673752 355474 673804
rect 540974 673752 540980 673804
rect 541032 673792 541038 673804
rect 548610 673792 548616 673804
rect 541032 673764 548616 673792
rect 541032 673752 541038 673764
rect 548610 673752 548616 673764
rect 548668 673752 548674 673804
rect 104894 673480 104900 673532
rect 104952 673520 104958 673532
rect 105078 673520 105084 673532
rect 104952 673492 105084 673520
rect 104952 673480 104958 673492
rect 105078 673480 105084 673492
rect 105136 673480 105142 673532
rect 494054 673480 494060 673532
rect 494112 673520 494118 673532
rect 494238 673520 494244 673532
rect 494112 673492 494244 673520
rect 494112 673480 494118 673492
rect 494238 673480 494244 673492
rect 494296 673480 494302 673532
rect 429194 673412 429200 673464
rect 429252 673452 429258 673464
rect 429470 673452 429476 673464
rect 429252 673424 429476 673452
rect 429252 673412 429258 673424
rect 429470 673412 429476 673424
rect 429528 673412 429534 673464
rect 364426 669400 364432 669452
rect 364484 669400 364490 669452
rect 364444 669316 364472 669400
rect 364426 669264 364432 669316
rect 364484 669264 364490 669316
rect 494054 669264 494060 669316
rect 494112 669304 494118 669316
rect 494238 669304 494244 669316
rect 494112 669276 494244 669304
rect 494112 669264 494118 669276
rect 494238 669264 494244 669276
rect 494296 669264 494302 669316
rect 3510 667904 3516 667956
rect 3568 667944 3574 667956
rect 21358 667944 21364 667956
rect 3568 667916 21364 667944
rect 3568 667904 3574 667916
rect 21358 667904 21364 667916
rect 21416 667904 21422 667956
rect 299658 666544 299664 666596
rect 299716 666584 299722 666596
rect 299934 666584 299940 666596
rect 299716 666556 299940 666584
rect 299716 666544 299722 666556
rect 299934 666544 299940 666556
rect 299992 666544 299998 666596
rect 493962 666476 493968 666528
rect 494020 666516 494026 666528
rect 494238 666516 494244 666528
rect 494020 666488 494244 666516
rect 494020 666476 494026 666488
rect 494238 666476 494244 666488
rect 494296 666476 494302 666528
rect 169938 661716 169944 661768
rect 169996 661756 170002 661768
rect 170214 661756 170220 661768
rect 169996 661728 170220 661756
rect 169996 661716 170002 661728
rect 170214 661716 170220 661728
rect 170272 661716 170278 661768
rect 559098 661716 559104 661768
rect 559156 661756 559162 661768
rect 559374 661756 559380 661768
rect 559156 661728 559380 661756
rect 559156 661716 559162 661728
rect 559374 661716 559380 661728
rect 559432 661716 559438 661768
rect 169938 656888 169944 656940
rect 169996 656928 170002 656940
rect 170030 656928 170036 656940
rect 169996 656900 170036 656928
rect 169996 656888 170002 656900
rect 170030 656888 170036 656900
rect 170088 656888 170094 656940
rect 493962 656888 493968 656940
rect 494020 656928 494026 656940
rect 494146 656928 494152 656940
rect 494020 656900 494152 656928
rect 494020 656888 494026 656900
rect 494146 656888 494152 656900
rect 494204 656888 494210 656940
rect 559098 656888 559104 656940
rect 559156 656928 559162 656940
rect 559190 656928 559196 656940
rect 559156 656900 559196 656928
rect 559156 656888 559162 656900
rect 559190 656888 559196 656900
rect 559248 656888 559254 656940
rect 299474 656820 299480 656872
rect 299532 656860 299538 656872
rect 299750 656860 299756 656872
rect 299532 656832 299756 656860
rect 299532 656820 299538 656832
rect 299750 656820 299756 656832
rect 299808 656820 299814 656872
rect 263502 653352 263508 653404
rect 263560 653392 263566 653404
rect 378134 653392 378140 653404
rect 263560 653364 378140 653392
rect 263560 653352 263566 653364
rect 378134 653352 378140 653364
rect 378192 653352 378198 653404
rect 139394 652848 139400 652860
rect 135272 652820 139400 652848
rect 3050 652740 3056 652792
rect 3108 652780 3114 652792
rect 13078 652780 13084 652792
rect 3108 652752 13084 652780
rect 3108 652740 3114 652752
rect 13078 652740 13084 652752
rect 13136 652740 13142 652792
rect 129274 652740 129280 652792
rect 129332 652780 129338 652792
rect 133690 652780 133696 652792
rect 129332 652752 133696 652780
rect 129332 652740 129338 652752
rect 133690 652740 133696 652752
rect 133748 652780 133754 652792
rect 135272 652780 135300 652820
rect 139394 652808 139400 652820
rect 139452 652848 139458 652860
rect 139452 652820 139716 652848
rect 139452 652808 139458 652820
rect 133748 652752 135300 652780
rect 139688 652780 139716 652820
rect 378134 652808 378140 652860
rect 378192 652848 378198 652860
rect 383470 652848 383476 652860
rect 378192 652820 383476 652848
rect 378192 652808 378198 652820
rect 383470 652808 383476 652820
rect 383528 652848 383534 652860
rect 387794 652848 387800 652860
rect 383528 652820 387800 652848
rect 383528 652808 383534 652820
rect 387794 652808 387800 652820
rect 387852 652808 387858 652860
rect 258626 652780 258632 652792
rect 139688 652752 258632 652780
rect 133748 652740 133754 652752
rect 258626 652740 258632 652752
rect 258684 652780 258690 652792
rect 263502 652780 263508 652792
rect 258684 652752 263508 652780
rect 258684 652740 258690 652752
rect 263502 652740 263508 652752
rect 263560 652740 263566 652792
rect 197354 650904 197360 650956
rect 197412 650944 197418 650956
rect 206922 650944 206928 650956
rect 197412 650916 206928 650944
rect 197412 650904 197418 650916
rect 206922 650904 206928 650916
rect 206980 650904 206986 650956
rect 195238 650768 195244 650820
rect 195296 650808 195302 650820
rect 197354 650808 197360 650820
rect 195296 650780 197360 650808
rect 195296 650768 195302 650780
rect 197354 650768 197360 650780
rect 197412 650768 197418 650820
rect 367094 650768 367100 650820
rect 367152 650808 367158 650820
rect 370406 650808 370412 650820
rect 367152 650780 370412 650808
rect 367152 650768 367158 650780
rect 370406 650768 370412 650780
rect 370464 650768 370470 650820
rect 57698 650700 57704 650752
rect 57756 650740 57762 650752
rect 105078 650740 105084 650752
rect 57756 650712 105084 650740
rect 57756 650700 57762 650712
rect 105078 650700 105084 650712
rect 105136 650700 105142 650752
rect 278774 650700 278780 650752
rect 278832 650740 278838 650752
rect 288342 650740 288348 650752
rect 278832 650712 288348 650740
rect 278832 650700 278838 650712
rect 288342 650700 288348 650712
rect 288400 650700 288406 650752
rect 572622 650700 572628 650752
rect 572680 650740 572686 650752
rect 579522 650740 579528 650752
rect 572680 650712 579528 650740
rect 572680 650700 572686 650712
rect 579522 650700 579528 650712
rect 579580 650700 579586 650752
rect 59446 650632 59452 650684
rect 59504 650672 59510 650684
rect 364518 650672 364524 650684
rect 59504 650644 364524 650672
rect 59504 650632 59510 650644
rect 364518 650632 364524 650644
rect 364576 650632 364582 650684
rect 89622 650564 89628 650616
rect 89680 650604 89686 650616
rect 96522 650604 96528 650616
rect 89680 650576 96528 650604
rect 89680 650564 89686 650576
rect 96522 650564 96528 650576
rect 96580 650564 96586 650616
rect 106734 650564 106740 650616
rect 106792 650604 106798 650616
rect 115750 650604 115756 650616
rect 106792 650576 115756 650604
rect 106792 650564 106798 650576
rect 115750 650564 115756 650576
rect 115808 650564 115814 650616
rect 207014 650564 207020 650616
rect 207072 650604 207078 650616
rect 207072 650576 215432 650604
rect 207072 650564 207078 650576
rect 115934 650496 115940 650548
rect 115992 650536 115998 650548
rect 120718 650536 120724 650548
rect 115992 650508 120724 650536
rect 115992 650496 115998 650508
rect 120718 650496 120724 650508
rect 120776 650496 120782 650548
rect 215404 650536 215432 650576
rect 219360 650576 225000 650604
rect 219360 650536 219388 650576
rect 177316 650508 186912 650536
rect 215404 650508 219388 650536
rect 137646 650428 137652 650480
rect 137704 650468 137710 650480
rect 147582 650468 147588 650480
rect 137704 650440 147588 650468
rect 137704 650428 137710 650440
rect 147582 650428 147588 650440
rect 147640 650428 147646 650480
rect 147674 650360 147680 650412
rect 147732 650400 147738 650412
rect 157242 650400 157248 650412
rect 147732 650372 157248 650400
rect 147732 650360 147738 650372
rect 157242 650360 157248 650372
rect 157300 650360 157306 650412
rect 157334 650360 157340 650412
rect 157392 650400 157398 650412
rect 157392 650372 157472 650400
rect 157392 650360 157398 650372
rect 157444 650332 157472 650372
rect 164142 650332 164148 650344
rect 157444 650304 164148 650332
rect 164142 650292 164148 650304
rect 164200 650292 164206 650344
rect 164234 650292 164240 650344
rect 164292 650332 164298 650344
rect 164292 650304 173756 650332
rect 164292 650292 164298 650304
rect 173728 650264 173756 650304
rect 177316 650264 177344 650508
rect 186884 650400 186912 650508
rect 224972 650468 225000 650576
rect 254044 650576 258120 650604
rect 237374 650536 237380 650548
rect 234724 650508 237380 650536
rect 224972 650440 228956 650468
rect 195238 650400 195244 650412
rect 186884 650372 195244 650400
rect 195238 650360 195244 650372
rect 195296 650360 195302 650412
rect 228928 650400 228956 650440
rect 234724 650400 234752 650508
rect 237374 650496 237380 650508
rect 237432 650496 237438 650548
rect 228928 650372 234752 650400
rect 237558 650360 237564 650412
rect 237616 650400 237622 650412
rect 254044 650400 254072 650576
rect 258092 650468 258120 650576
rect 340782 650564 340788 650616
rect 340840 650604 340846 650616
rect 347682 650604 347688 650616
rect 340840 650576 347688 650604
rect 340840 650564 340846 650576
rect 347682 650564 347688 650576
rect 347740 650564 347746 650616
rect 560294 650564 560300 650616
rect 560352 650604 560358 650616
rect 563146 650604 563152 650616
rect 560352 650576 563152 650604
rect 560352 650564 560358 650576
rect 563146 650564 563152 650576
rect 563204 650564 563210 650616
rect 289814 650496 289820 650548
rect 289872 650536 289878 650548
rect 292666 650536 292672 650548
rect 289872 650508 292672 650536
rect 289872 650496 289878 650508
rect 292666 650496 292672 650508
rect 292724 650496 292730 650548
rect 405734 650496 405740 650548
rect 405792 650536 405798 650548
rect 413370 650536 413376 650548
rect 405792 650508 413376 650536
rect 405792 650496 405798 650508
rect 413370 650496 413376 650508
rect 413428 650496 413434 650548
rect 533982 650496 533988 650548
rect 534040 650536 534046 650548
rect 540882 650536 540888 650548
rect 534040 650508 540888 650536
rect 534040 650496 534046 650508
rect 540882 650496 540888 650508
rect 540940 650496 540946 650548
rect 266354 650468 266360 650480
rect 258092 650440 266360 650468
rect 266354 650428 266360 650440
rect 266412 650428 266418 650480
rect 456702 650428 456708 650480
rect 456760 650468 456766 650480
rect 463602 650468 463608 650480
rect 456760 650440 463608 650468
rect 456760 650428 456766 650440
rect 463602 650428 463608 650440
rect 463660 650428 463666 650480
rect 476022 650428 476028 650480
rect 476080 650468 476086 650480
rect 482922 650468 482928 650480
rect 476080 650440 482928 650468
rect 476080 650428 476086 650440
rect 482922 650428 482928 650440
rect 482980 650428 482986 650480
rect 495342 650428 495348 650480
rect 495400 650468 495406 650480
rect 502242 650468 502248 650480
rect 495400 650440 502248 650468
rect 495400 650428 495406 650440
rect 502242 650428 502248 650440
rect 502300 650428 502306 650480
rect 514662 650428 514668 650480
rect 514720 650468 514726 650480
rect 521562 650468 521568 650480
rect 514720 650440 521568 650468
rect 514720 650428 514726 650440
rect 521562 650428 521568 650440
rect 521620 650428 521626 650480
rect 237616 650372 254072 650400
rect 237616 650360 237622 650372
rect 285582 650292 285588 650344
rect 285640 650332 285646 650344
rect 386414 650332 386420 650344
rect 285640 650304 386420 650332
rect 285640 650292 285646 650304
rect 386414 650292 386420 650304
rect 386472 650292 386478 650344
rect 173728 650236 177344 650264
rect 285582 650196 285588 650208
rect 282840 650168 285588 650196
rect 280062 650088 280068 650140
rect 280120 650128 280126 650140
rect 282840 650128 282868 650168
rect 285582 650156 285588 650168
rect 285640 650156 285646 650208
rect 280120 650100 282868 650128
rect 280120 650088 280126 650100
rect 266354 650020 266360 650072
rect 266412 650060 266418 650072
rect 270494 650060 270500 650072
rect 266412 650032 270500 650060
rect 266412 650020 266418 650032
rect 270494 650020 270500 650032
rect 270552 650020 270558 650072
rect 169938 647232 169944 647284
rect 169996 647272 170002 647284
rect 170030 647272 170036 647284
rect 169996 647244 170036 647272
rect 169996 647232 170002 647244
rect 170030 647232 170036 647244
rect 170088 647232 170094 647284
rect 299474 647232 299480 647284
rect 299532 647272 299538 647284
rect 299658 647272 299664 647284
rect 299532 647244 299664 647272
rect 299532 647232 299538 647244
rect 299658 647232 299664 647244
rect 299716 647232 299722 647284
rect 429378 647232 429384 647284
rect 429436 647272 429442 647284
rect 429470 647272 429476 647284
rect 429436 647244 429476 647272
rect 429436 647232 429442 647244
rect 429470 647232 429476 647244
rect 429528 647232 429534 647284
rect 559098 647232 559104 647284
rect 559156 647272 559162 647284
rect 559190 647272 559196 647284
rect 559156 647244 559196 647272
rect 559156 647232 559162 647244
rect 559190 647232 559196 647244
rect 559248 647232 559254 647284
rect 297358 645872 297364 645924
rect 297416 645912 297422 645924
rect 307110 645912 307116 645924
rect 297416 645884 307116 645912
rect 297416 645872 297422 645884
rect 307110 645872 307116 645884
rect 307168 645872 307174 645924
rect 294598 644444 294604 644496
rect 294656 644484 294662 644496
rect 307110 644484 307116 644496
rect 294656 644456 307116 644484
rect 294656 644444 294662 644456
rect 307110 644444 307116 644456
rect 307168 644444 307174 644496
rect 291838 643084 291844 643136
rect 291896 643124 291902 643136
rect 307110 643124 307116 643136
rect 291896 643096 307116 643124
rect 291896 643084 291902 643096
rect 307110 643084 307116 643096
rect 307168 643084 307174 643136
rect 290458 641724 290464 641776
rect 290516 641764 290522 641776
rect 307662 641764 307668 641776
rect 290516 641736 307668 641764
rect 290516 641724 290522 641736
rect 307662 641724 307668 641736
rect 307720 641724 307726 641776
rect 169938 640364 169944 640416
rect 169996 640404 170002 640416
rect 170030 640404 170036 640416
rect 169996 640376 170036 640404
rect 169996 640364 170002 640376
rect 170030 640364 170036 640376
rect 170088 640364 170094 640416
rect 429378 640364 429384 640416
rect 429436 640404 429442 640416
rect 429470 640404 429476 640416
rect 429436 640376 429476 640404
rect 429436 640364 429442 640376
rect 429470 640364 429476 640376
rect 429528 640364 429534 640416
rect 559098 640364 559104 640416
rect 559156 640404 559162 640416
rect 559190 640404 559196 640416
rect 559156 640376 559196 640404
rect 559156 640364 559162 640376
rect 559190 640364 559196 640376
rect 559248 640364 559254 640416
rect 287698 640296 287704 640348
rect 287756 640336 287762 640348
rect 307662 640336 307668 640348
rect 287756 640308 307668 640336
rect 287756 640296 287762 640308
rect 307662 640296 307668 640308
rect 307720 640296 307726 640348
rect 286318 638936 286324 638988
rect 286376 638976 286382 638988
rect 306650 638976 306656 638988
rect 286376 638948 306656 638976
rect 286376 638936 286382 638948
rect 306650 638936 306656 638948
rect 306708 638936 306714 638988
rect 301498 637576 301504 637628
rect 301556 637616 301562 637628
rect 306834 637616 306840 637628
rect 301556 637588 306840 637616
rect 301556 637576 301562 637588
rect 306834 637576 306840 637588
rect 306892 637576 306898 637628
rect 494054 634788 494060 634840
rect 494112 634828 494118 634840
rect 494238 634828 494244 634840
rect 494112 634800 494244 634828
rect 494112 634788 494118 634800
rect 494238 634788 494244 634800
rect 494296 634788 494302 634840
rect 299658 630708 299664 630760
rect 299716 630748 299722 630760
rect 299750 630748 299756 630760
rect 299716 630720 299756 630748
rect 299716 630708 299722 630720
rect 299750 630708 299756 630720
rect 299808 630708 299814 630760
rect 169846 630640 169852 630692
rect 169904 630680 169910 630692
rect 170030 630680 170036 630692
rect 169904 630652 170036 630680
rect 169904 630640 169910 630652
rect 170030 630640 170036 630652
rect 170088 630640 170094 630692
rect 429286 630640 429292 630692
rect 429344 630680 429350 630692
rect 429470 630680 429476 630692
rect 429344 630652 429476 630680
rect 429344 630640 429350 630652
rect 429470 630640 429476 630652
rect 429528 630640 429534 630692
rect 559006 630640 559012 630692
rect 559064 630680 559070 630692
rect 559190 630680 559196 630692
rect 559064 630652 559196 630680
rect 559064 630640 559070 630652
rect 559190 630640 559196 630652
rect 559248 630640 559254 630692
rect 494054 615476 494060 615528
rect 494112 615516 494118 615528
rect 494238 615516 494244 615528
rect 494112 615488 494244 615516
rect 494112 615476 494118 615488
rect 494238 615476 494244 615488
rect 494296 615476 494302 615528
rect 169846 611328 169852 611380
rect 169904 611368 169910 611380
rect 170030 611368 170036 611380
rect 169904 611340 170036 611368
rect 169904 611328 169910 611340
rect 170030 611328 170036 611340
rect 170088 611328 170094 611380
rect 299566 611328 299572 611380
rect 299624 611368 299630 611380
rect 299750 611368 299756 611380
rect 299624 611340 299756 611368
rect 299624 611328 299630 611340
rect 299750 611328 299756 611340
rect 299808 611328 299814 611380
rect 429286 611328 429292 611380
rect 429344 611368 429350 611380
rect 429470 611368 429476 611380
rect 429344 611340 429476 611368
rect 429344 611328 429350 611340
rect 429470 611328 429476 611340
rect 429528 611328 429534 611380
rect 559006 611328 559012 611380
rect 559064 611368 559070 611380
rect 559190 611368 559196 611380
rect 559064 611340 559196 611368
rect 559064 611328 559070 611340
rect 559190 611328 559196 611340
rect 559248 611328 559254 611380
rect 3602 609968 3608 610020
rect 3660 610008 3666 610020
rect 31018 610008 31024 610020
rect 3660 609980 31024 610008
rect 3660 609968 3666 609980
rect 31018 609968 31024 609980
rect 31076 609968 31082 610020
rect 169846 608540 169852 608592
rect 169904 608580 169910 608592
rect 169938 608580 169944 608592
rect 169904 608552 169944 608580
rect 169904 608540 169910 608552
rect 169938 608540 169944 608552
rect 169996 608540 170002 608592
rect 299566 608540 299572 608592
rect 299624 608580 299630 608592
rect 299658 608580 299664 608592
rect 299624 608552 299664 608580
rect 299624 608540 299630 608552
rect 299658 608540 299664 608552
rect 299716 608540 299722 608592
rect 429286 608540 429292 608592
rect 429344 608580 429350 608592
rect 429378 608580 429384 608592
rect 429344 608552 429384 608580
rect 429344 608540 429350 608552
rect 429378 608540 429384 608552
rect 429436 608540 429442 608592
rect 559006 608540 559012 608592
rect 559064 608580 559070 608592
rect 559098 608580 559104 608592
rect 559064 608552 559104 608580
rect 559064 608540 559070 608552
rect 559098 608540 559104 608552
rect 559156 608540 559162 608592
rect 169846 601672 169852 601724
rect 169904 601712 169910 601724
rect 170122 601712 170128 601724
rect 169904 601684 170128 601712
rect 169904 601672 169910 601684
rect 170122 601672 170128 601684
rect 170180 601672 170186 601724
rect 299566 601672 299572 601724
rect 299624 601712 299630 601724
rect 299842 601712 299848 601724
rect 299624 601684 299848 601712
rect 299624 601672 299630 601684
rect 299842 601672 299848 601684
rect 299900 601672 299906 601724
rect 429286 601672 429292 601724
rect 429344 601712 429350 601724
rect 429562 601712 429568 601724
rect 429344 601684 429568 601712
rect 429344 601672 429350 601684
rect 429562 601672 429568 601684
rect 429620 601672 429626 601724
rect 559006 601672 559012 601724
rect 559064 601712 559070 601724
rect 559282 601712 559288 601724
rect 559064 601684 559288 601712
rect 559064 601672 559070 601684
rect 559282 601672 559288 601684
rect 559340 601672 559346 601724
rect 169938 598884 169944 598936
rect 169996 598924 170002 598936
rect 170122 598924 170128 598936
rect 169996 598896 170128 598924
rect 169996 598884 170002 598896
rect 170122 598884 170128 598896
rect 170180 598884 170186 598936
rect 299658 598884 299664 598936
rect 299716 598924 299722 598936
rect 299842 598924 299848 598936
rect 299716 598896 299848 598924
rect 299716 598884 299722 598896
rect 299842 598884 299848 598896
rect 299900 598884 299906 598936
rect 559098 598884 559104 598936
rect 559156 598924 559162 598936
rect 559282 598924 559288 598936
rect 559156 598896 559288 598924
rect 559156 598884 559162 598896
rect 559282 598884 559288 598896
rect 559340 598884 559346 598936
rect 494054 596164 494060 596216
rect 494112 596204 494118 596216
rect 494238 596204 494244 596216
rect 494112 596176 494244 596204
rect 494112 596164 494118 596176
rect 494238 596164 494244 596176
rect 494296 596164 494302 596216
rect 3326 594804 3332 594856
rect 3384 594844 3390 594856
rect 14458 594844 14464 594856
rect 3384 594816 14464 594844
rect 3384 594804 3390 594816
rect 14458 594804 14464 594816
rect 14516 594804 14522 594856
rect 429562 592016 429568 592068
rect 429620 592016 429626 592068
rect 429580 591920 429608 592016
rect 429654 591920 429660 591932
rect 429580 591892 429660 591920
rect 429654 591880 429660 591892
rect 429712 591880 429718 591932
rect 169938 589296 169944 589348
rect 169996 589336 170002 589348
rect 170214 589336 170220 589348
rect 169996 589308 170220 589336
rect 169996 589296 170002 589308
rect 170214 589296 170220 589308
rect 170272 589296 170278 589348
rect 270402 589296 270408 589348
rect 270460 589336 270466 589348
rect 309778 589336 309784 589348
rect 270460 589308 309784 589336
rect 270460 589296 270466 589308
rect 309778 589296 309784 589308
rect 309836 589296 309842 589348
rect 559098 589296 559104 589348
rect 559156 589336 559162 589348
rect 559374 589336 559380 589348
rect 559156 589308 559380 589336
rect 559156 589296 559162 589308
rect 559374 589296 559380 589308
rect 559432 589296 559438 589348
rect 493870 589228 493876 589280
rect 493928 589268 493934 589280
rect 494146 589268 494152 589280
rect 493928 589240 494152 589268
rect 493928 589228 493934 589240
rect 494146 589228 494152 589240
rect 494204 589228 494210 589280
rect 429286 583040 429292 583092
rect 429344 583080 429350 583092
rect 429562 583080 429568 583092
rect 429344 583052 429568 583080
rect 429344 583040 429350 583052
rect 429562 583040 429568 583052
rect 429620 583040 429626 583092
rect 170214 582468 170220 582480
rect 170140 582440 170220 582468
rect 170140 582344 170168 582440
rect 170214 582428 170220 582440
rect 170272 582428 170278 582480
rect 299934 582468 299940 582480
rect 299860 582440 299940 582468
rect 299860 582344 299888 582440
rect 299934 582428 299940 582440
rect 299992 582428 299998 582480
rect 559374 582468 559380 582480
rect 559300 582440 559380 582468
rect 559300 582344 559328 582440
rect 559374 582428 559380 582440
rect 559432 582428 559438 582480
rect 170122 582292 170128 582344
rect 170180 582292 170186 582344
rect 299842 582292 299848 582344
rect 299900 582292 299906 582344
rect 559282 582292 559288 582344
rect 559340 582292 559346 582344
rect 493870 579640 493876 579692
rect 493928 579680 493934 579692
rect 494054 579680 494060 579692
rect 493928 579652 494060 579680
rect 493928 579640 493934 579652
rect 494054 579640 494060 579652
rect 494112 579640 494118 579692
rect 429286 578212 429292 578264
rect 429344 578252 429350 578264
rect 429378 578252 429384 578264
rect 429344 578224 429384 578252
rect 429344 578212 429350 578224
rect 429378 578212 429384 578224
rect 429436 578212 429442 578264
rect 429378 572568 429384 572620
rect 429436 572608 429442 572620
rect 429654 572608 429660 572620
rect 429436 572580 429660 572608
rect 429436 572568 429442 572580
rect 429654 572568 429660 572580
rect 429712 572568 429718 572620
rect 494146 569848 494152 569900
rect 494204 569888 494210 569900
rect 494330 569888 494336 569900
rect 494204 569860 494336 569888
rect 494204 569848 494210 569860
rect 494330 569848 494336 569860
rect 494388 569848 494394 569900
rect 494330 563184 494336 563236
rect 494388 563184 494394 563236
rect 494348 563100 494376 563184
rect 494330 563048 494336 563100
rect 494388 563048 494394 563100
rect 56870 560872 56876 560924
rect 56928 560912 56934 560924
rect 188982 560912 188988 560924
rect 56928 560884 188988 560912
rect 56928 560872 56934 560884
rect 188982 560872 188988 560884
rect 189040 560912 189046 560924
rect 305638 560912 305644 560924
rect 189040 560884 305644 560912
rect 189040 560872 189046 560884
rect 305638 560872 305644 560884
rect 305696 560872 305702 560924
rect 429470 560260 429476 560312
rect 429528 560300 429534 560312
rect 429654 560300 429660 560312
rect 429528 560272 429660 560300
rect 429528 560260 429534 560272
rect 429654 560260 429660 560272
rect 429712 560260 429718 560312
rect 559006 560260 559012 560312
rect 559064 560300 559070 560312
rect 559098 560300 559104 560312
rect 559064 560272 559104 560300
rect 559064 560260 559070 560272
rect 559098 560260 559104 560272
rect 559156 560260 559162 560312
rect 309778 560192 309784 560244
rect 309836 560232 309842 560244
rect 310422 560232 310428 560244
rect 309836 560204 310428 560232
rect 309836 560192 309842 560204
rect 310422 560192 310428 560204
rect 310480 560232 310486 560244
rect 389174 560232 389180 560244
rect 310480 560204 389180 560232
rect 310480 560192 310486 560204
rect 389174 560192 389180 560204
rect 389232 560192 389238 560244
rect 62022 558832 62028 558884
rect 62080 558872 62086 558884
rect 197354 558872 197360 558884
rect 62080 558844 197360 558872
rect 62080 558832 62086 558844
rect 197354 558832 197360 558844
rect 197412 558832 197418 558884
rect 215294 558832 215300 558884
rect 215352 558872 215358 558884
rect 224494 558872 224500 558884
rect 215352 558844 224500 558872
rect 215352 558832 215358 558844
rect 224494 558832 224500 558844
rect 224552 558832 224558 558884
rect 335446 558832 335452 558884
rect 335504 558872 335510 558884
rect 344830 558872 344836 558884
rect 335504 558844 344836 558872
rect 335504 558832 335510 558844
rect 344830 558832 344836 558844
rect 344888 558832 344894 558884
rect 67450 558764 67456 558816
rect 67508 558804 67514 558816
rect 201494 558804 201500 558816
rect 67508 558776 201500 558804
rect 67508 558764 67514 558776
rect 201494 558764 201500 558776
rect 201552 558764 201558 558816
rect 328454 558764 328460 558816
rect 328512 558804 328518 558816
rect 338022 558804 338028 558816
rect 328512 558776 338028 558804
rect 328512 558764 328518 558776
rect 338022 558764 338028 558776
rect 338080 558764 338086 558816
rect 77386 558696 77392 558748
rect 77444 558736 77450 558748
rect 86402 558736 86408 558748
rect 77444 558708 86408 558736
rect 77444 558696 77450 558708
rect 86402 558696 86408 558708
rect 86460 558736 86466 558748
rect 95786 558736 95792 558748
rect 86460 558708 95792 558736
rect 86460 558696 86466 558708
rect 95786 558696 95792 558708
rect 95844 558736 95850 558748
rect 105538 558736 105544 558748
rect 95844 558708 105544 558736
rect 95844 558696 95850 558708
rect 105538 558696 105544 558708
rect 105596 558696 105602 558748
rect 125502 558696 125508 558748
rect 125560 558736 125566 558748
rect 208394 558736 208400 558748
rect 125560 558708 208400 558736
rect 125560 558696 125566 558708
rect 208394 558696 208400 558708
rect 208452 558736 208458 558748
rect 209682 558736 209688 558748
rect 208452 558708 209688 558736
rect 208452 558696 208458 558708
rect 209682 558696 209688 558708
rect 209740 558696 209746 558748
rect 223574 558696 223580 558748
rect 223632 558736 223638 558748
rect 231854 558736 231860 558748
rect 223632 558708 231860 558736
rect 223632 558696 223638 558708
rect 231854 558696 231860 558708
rect 231912 558696 231918 558748
rect 328546 558696 328552 558748
rect 328604 558736 328610 558748
rect 337930 558736 337936 558748
rect 328604 558708 337936 558736
rect 328604 558696 328610 558708
rect 337930 558696 337936 558708
rect 337988 558696 337994 558748
rect 76006 558628 76012 558680
rect 76064 558668 76070 558680
rect 76064 558640 84240 558668
rect 76064 558628 76070 558640
rect 84212 558600 84240 558640
rect 84286 558628 84292 558680
rect 84344 558668 84350 558680
rect 93302 558668 93308 558680
rect 84344 558640 93308 558668
rect 84344 558628 84350 558640
rect 93302 558628 93308 558640
rect 93360 558628 93366 558680
rect 97810 558628 97816 558680
rect 97868 558668 97874 558680
rect 133138 558668 133144 558680
rect 97868 558640 133144 558668
rect 97868 558628 97874 558640
rect 133138 558628 133144 558640
rect 133196 558628 133202 558680
rect 224494 558628 224500 558680
rect 224552 558668 224558 558680
rect 233234 558668 233240 558680
rect 224552 558640 233240 558668
rect 224552 558628 224558 558640
rect 233234 558628 233240 558640
rect 233292 558628 233298 558680
rect 344830 558628 344836 558680
rect 344888 558668 344894 558680
rect 353294 558668 353300 558680
rect 344888 558640 353300 558668
rect 344888 558628 344894 558640
rect 353294 558628 353300 558640
rect 353352 558628 353358 558680
rect 85206 558600 85212 558612
rect 84212 558572 85212 558600
rect 85206 558560 85212 558572
rect 85264 558600 85270 558612
rect 94866 558600 94872 558612
rect 85264 558572 94872 558600
rect 85264 558560 85270 558572
rect 94866 558560 94872 558572
rect 94924 558600 94930 558612
rect 103882 558600 103888 558612
rect 94924 558572 103888 558600
rect 94924 558560 94930 558572
rect 103882 558560 103888 558572
rect 103940 558600 103946 558612
rect 104158 558600 104164 558612
rect 103940 558572 104164 558600
rect 103940 558560 103946 558572
rect 104158 558560 104164 558572
rect 104216 558560 104222 558612
rect 104802 558560 104808 558612
rect 104860 558600 104866 558612
rect 137370 558600 137376 558612
rect 104860 558572 137376 558600
rect 104860 558560 104866 558572
rect 137370 558560 137376 558572
rect 137428 558560 137434 558612
rect 217778 558560 217784 558612
rect 217836 558600 217842 558612
rect 225874 558600 225880 558612
rect 217836 558572 225880 558600
rect 217836 558560 217842 558572
rect 225874 558560 225880 558572
rect 225932 558600 225938 558612
rect 234890 558600 234896 558612
rect 225932 558572 234896 558600
rect 225932 558560 225938 558572
rect 234890 558560 234896 558572
rect 234948 558560 234954 558612
rect 336458 558560 336464 558612
rect 336516 558600 336522 558612
rect 345750 558600 345756 558612
rect 336516 558572 345756 558600
rect 336516 558560 336522 558572
rect 345750 558560 345756 558572
rect 345808 558600 345814 558612
rect 354674 558600 354680 558612
rect 345808 558572 354680 558600
rect 345808 558560 345814 558572
rect 354674 558560 354680 558572
rect 354732 558560 354738 558612
rect 79594 558492 79600 558544
rect 79652 558532 79658 558544
rect 88886 558532 88892 558544
rect 79652 558504 88892 558532
rect 79652 558492 79658 558504
rect 88886 558492 88892 558504
rect 88944 558532 88950 558544
rect 98086 558532 98092 558544
rect 88944 558504 98092 558532
rect 88944 558492 88950 558504
rect 98086 558492 98092 558504
rect 98144 558492 98150 558544
rect 99558 558492 99564 558544
rect 99616 558532 99622 558544
rect 108298 558532 108304 558544
rect 99616 558504 108304 558532
rect 99616 558492 99622 558504
rect 108298 558492 108304 558504
rect 108356 558492 108362 558544
rect 209682 558492 209688 558544
rect 209740 558532 209746 558544
rect 217962 558532 217968 558544
rect 209740 558504 217968 558532
rect 209740 558492 209746 558504
rect 217962 558492 217968 558504
rect 218020 558492 218026 558544
rect 223574 558532 223580 558544
rect 221292 558504 223580 558532
rect 78490 558424 78496 558476
rect 78548 558464 78554 558476
rect 87874 558464 87880 558476
rect 78548 558436 87880 558464
rect 78548 558424 78554 558436
rect 87874 558424 87880 558436
rect 87932 558464 87938 558476
rect 96982 558464 96988 558476
rect 87932 558436 96988 558464
rect 87932 558424 87938 558436
rect 96982 558424 96988 558436
rect 97040 558464 97046 558476
rect 106918 558464 106924 558476
rect 97040 558436 106924 558464
rect 97040 558424 97046 558436
rect 106918 558424 106924 558436
rect 106976 558424 106982 558476
rect 108482 558424 108488 558476
rect 108540 558464 108546 558476
rect 144178 558464 144184 558476
rect 108540 558436 144184 558464
rect 108540 558424 108546 558436
rect 144178 558424 144184 558436
rect 144236 558424 144242 558476
rect 213914 558424 213920 558476
rect 213972 558464 213978 558476
rect 221292 558464 221320 558504
rect 223574 558492 223580 558504
rect 223632 558492 223638 558544
rect 330478 558492 330484 558544
rect 330536 558532 330542 558544
rect 339862 558532 339868 558544
rect 330536 558504 339868 558532
rect 330536 558492 330542 558504
rect 339862 558492 339868 558504
rect 339920 558532 339926 558544
rect 349522 558532 349528 558544
rect 339920 558504 349528 558532
rect 339920 558492 339926 558504
rect 349522 558492 349528 558504
rect 349580 558532 349586 558544
rect 357710 558532 357716 558544
rect 349580 558504 357716 558532
rect 349580 558492 349586 558504
rect 357710 558492 357716 558504
rect 357768 558492 357774 558544
rect 227162 558464 227168 558476
rect 213972 558436 221320 558464
rect 221384 558436 227168 558464
rect 213972 558424 213978 558436
rect 80790 558356 80796 558408
rect 80848 558396 80854 558408
rect 89806 558396 89812 558408
rect 80848 558368 89812 558396
rect 80848 558356 80854 558368
rect 89806 558356 89812 558368
rect 89864 558396 89870 558408
rect 99558 558396 99564 558408
rect 89864 558368 99564 558396
rect 89864 558356 89870 558368
rect 99558 558356 99564 558368
rect 99616 558356 99622 558408
rect 100570 558396 100576 558408
rect 100312 558368 100576 558396
rect 72602 558288 72608 558340
rect 72660 558328 72666 558340
rect 81894 558328 81900 558340
rect 72660 558300 81900 558328
rect 72660 558288 72666 558300
rect 81894 558288 81900 558300
rect 81952 558328 81958 558340
rect 91094 558328 91100 558340
rect 81952 558300 91100 558328
rect 81952 558288 81958 558300
rect 91094 558288 91100 558300
rect 91152 558288 91158 558340
rect 92474 558288 92480 558340
rect 92532 558328 92538 558340
rect 97994 558328 98000 558340
rect 92532 558300 98000 558328
rect 92532 558288 92538 558300
rect 97994 558288 98000 558300
rect 98052 558288 98058 558340
rect 98086 558288 98092 558340
rect 98144 558328 98150 558340
rect 100312 558328 100340 558368
rect 100570 558356 100576 558368
rect 100628 558356 100634 558408
rect 101950 558356 101956 558408
rect 102008 558396 102014 558408
rect 140038 558396 140044 558408
rect 102008 558368 140044 558396
rect 102008 558356 102014 558368
rect 140038 558356 140044 558368
rect 140096 558356 140102 558408
rect 208578 558356 208584 558408
rect 208636 558396 208642 558408
rect 210602 558396 210608 558408
rect 208636 558368 210608 558396
rect 208636 558356 208642 558368
rect 210602 558356 210608 558368
rect 210660 558396 210666 558408
rect 210660 558368 217916 558396
rect 210660 558356 210666 558368
rect 98144 558300 100340 558328
rect 98144 558288 98150 558300
rect 100386 558288 100392 558340
rect 100444 558328 100450 558340
rect 140130 558328 140136 558340
rect 100444 558300 140136 558328
rect 100444 558288 100450 558300
rect 140130 558288 140136 558300
rect 140188 558288 140194 558340
rect 211154 558288 211160 558340
rect 211212 558328 211218 558340
rect 211798 558328 211804 558340
rect 211212 558300 211804 558328
rect 211212 558288 211218 558300
rect 211798 558288 211804 558300
rect 211856 558328 211862 558340
rect 215110 558328 215116 558340
rect 211856 558300 215116 558328
rect 211856 558288 211862 558300
rect 215110 558288 215116 558300
rect 215168 558288 215174 558340
rect 217888 558328 217916 558368
rect 217962 558356 217968 558408
rect 218020 558396 218026 558408
rect 221384 558396 221412 558436
rect 227162 558424 227168 558436
rect 227220 558464 227226 558476
rect 231854 558464 231860 558476
rect 227220 558436 231860 558464
rect 227220 558424 227226 558436
rect 231854 558424 231860 558436
rect 231912 558424 231918 558476
rect 337746 558424 337752 558476
rect 337804 558464 337810 558476
rect 346854 558464 346860 558476
rect 337804 558436 346860 558464
rect 337804 558424 337810 558436
rect 346854 558424 346860 558436
rect 346912 558464 346918 558476
rect 356054 558464 356060 558476
rect 346912 558436 356060 558464
rect 346912 558424 346918 558436
rect 356054 558424 356060 558436
rect 356112 558424 356118 558476
rect 229554 558396 229560 558408
rect 218020 558368 221412 558396
rect 221476 558368 229560 558396
rect 218020 558356 218026 558368
rect 220078 558328 220084 558340
rect 217888 558300 220084 558328
rect 220078 558288 220084 558300
rect 220136 558328 220142 558340
rect 220814 558328 220820 558340
rect 220136 558300 220820 558328
rect 220136 558288 220142 558300
rect 220814 558288 220820 558300
rect 220872 558288 220878 558340
rect 221090 558288 221096 558340
rect 221148 558328 221154 558340
rect 221476 558328 221504 558368
rect 229554 558356 229560 558368
rect 229612 558396 229618 558408
rect 238754 558396 238760 558408
rect 229612 558368 238760 558396
rect 229612 558356 229618 558368
rect 238754 558356 238760 558368
rect 238812 558356 238818 558408
rect 329282 558356 329288 558408
rect 329340 558396 329346 558408
rect 339034 558396 339040 558408
rect 329340 558368 339040 558396
rect 329340 558356 329346 558368
rect 339034 558356 339040 558368
rect 339092 558396 339098 558408
rect 348234 558396 348240 558408
rect 339092 558368 348240 558396
rect 339092 558356 339098 558368
rect 348234 558356 348240 558368
rect 348292 558396 348298 558408
rect 357434 558396 357440 558408
rect 348292 558368 357440 558396
rect 348292 558356 348298 558368
rect 357434 558356 357440 558368
rect 357492 558356 357498 558408
rect 221148 558300 221504 558328
rect 221148 558288 221154 558300
rect 221550 558288 221556 558340
rect 221608 558328 221614 558340
rect 230474 558328 230480 558340
rect 221608 558300 230480 558328
rect 221608 558288 221614 558300
rect 230474 558288 230480 558300
rect 230532 558288 230538 558340
rect 332686 558288 332692 558340
rect 332744 558328 332750 558340
rect 342530 558328 342536 558340
rect 332744 558300 342536 558328
rect 332744 558288 332750 558300
rect 342530 558288 342536 558300
rect 342588 558328 342594 558340
rect 348142 558328 348148 558340
rect 342588 558300 348148 558328
rect 342588 558288 342594 558300
rect 348142 558288 348148 558300
rect 348200 558288 348206 558340
rect 81250 558220 81256 558272
rect 81308 558260 81314 558272
rect 145558 558260 145564 558272
rect 81308 558232 145564 558260
rect 81308 558220 81314 558232
rect 145558 558220 145564 558232
rect 145616 558220 145622 558272
rect 222378 558260 222384 558272
rect 221660 558232 222384 558260
rect 76834 558152 76840 558204
rect 76892 558192 76898 558204
rect 141418 558192 141424 558204
rect 76892 558164 141424 558192
rect 76892 558152 76898 558164
rect 141418 558152 141424 558164
rect 141476 558152 141482 558204
rect 206922 558152 206928 558204
rect 206980 558192 206986 558204
rect 215294 558192 215300 558204
rect 206980 558164 215300 558192
rect 206980 558152 206986 558164
rect 215294 558152 215300 558164
rect 215352 558152 215358 558204
rect 221660 558192 221688 558232
rect 222378 558220 222384 558232
rect 222436 558260 222442 558272
rect 231854 558260 231860 558272
rect 222436 558232 231860 558260
rect 222436 558220 222442 558232
rect 231854 558220 231860 558232
rect 231912 558220 231918 558272
rect 331306 558220 331312 558272
rect 331364 558260 331370 558272
rect 331766 558260 331772 558272
rect 331364 558232 331772 558260
rect 331364 558220 331370 558232
rect 331766 558220 331772 558232
rect 331824 558260 331830 558272
rect 341242 558260 341248 558272
rect 331824 558232 341248 558260
rect 331824 558220 331830 558232
rect 341242 558220 341248 558232
rect 341300 558260 341306 558272
rect 350534 558260 350540 558272
rect 341300 558232 350540 558260
rect 341300 558220 341306 558232
rect 350534 558220 350540 558232
rect 350592 558220 350598 558272
rect 228174 558192 228180 558204
rect 218900 558164 221688 558192
rect 224972 558164 228180 558192
rect 73798 558084 73804 558136
rect 73856 558124 73862 558136
rect 82814 558124 82820 558136
rect 73856 558096 82820 558124
rect 73856 558084 73862 558096
rect 82814 558084 82820 558096
rect 82872 558084 82878 558136
rect 83826 558084 83832 558136
rect 83884 558124 83890 558136
rect 152458 558124 152464 558136
rect 83884 558096 152464 558124
rect 83884 558084 83890 558096
rect 152458 558084 152464 558096
rect 152516 558084 152522 558136
rect 79410 558016 79416 558068
rect 79468 558056 79474 558068
rect 148318 558056 148324 558068
rect 79468 558028 148324 558056
rect 79468 558016 79474 558028
rect 148318 558016 148324 558028
rect 148376 558016 148382 558068
rect 200114 558016 200120 558068
rect 200172 558056 200178 558068
rect 213638 558056 213644 558068
rect 200172 558028 213644 558056
rect 200172 558016 200178 558028
rect 213638 558016 213644 558028
rect 213696 558016 213702 558068
rect 74258 557948 74264 558000
rect 74316 557988 74322 558000
rect 135898 557988 135904 558000
rect 74316 557960 135904 557988
rect 74316 557948 74322 557960
rect 135898 557948 135904 557960
rect 135956 557948 135962 558000
rect 194410 557948 194416 558000
rect 194468 557988 194474 558000
rect 200022 557988 200028 558000
rect 194468 557960 200028 557988
rect 194468 557948 194474 557960
rect 200022 557948 200028 557960
rect 200080 557948 200086 558000
rect 203518 557948 203524 558000
rect 203576 557988 203582 558000
rect 213086 557988 213092 558000
rect 203576 557960 213092 557988
rect 203576 557948 203582 557960
rect 213086 557948 213092 557960
rect 213144 557988 213150 558000
rect 218900 557988 218928 558164
rect 218974 558016 218980 558068
rect 219032 558056 219038 558068
rect 224972 558056 225000 558164
rect 228174 558152 228180 558164
rect 228232 558192 228238 558204
rect 237374 558192 237380 558204
rect 228232 558164 237380 558192
rect 228232 558152 228238 558164
rect 237374 558152 237380 558164
rect 237432 558152 237438 558204
rect 288526 558152 288532 558204
rect 288584 558192 288590 558204
rect 298002 558192 298008 558204
rect 288584 558164 298008 558192
rect 288584 558152 288590 558164
rect 298002 558152 298008 558164
rect 298060 558152 298066 558204
rect 302234 558152 302240 558204
rect 302292 558192 302298 558204
rect 313366 558192 313372 558204
rect 302292 558164 313372 558192
rect 302292 558152 302298 558164
rect 313366 558152 313372 558164
rect 313424 558152 313430 558204
rect 334066 558152 334072 558204
rect 334124 558192 334130 558204
rect 343634 558192 343640 558204
rect 334124 558164 343640 558192
rect 334124 558152 334130 558164
rect 343634 558152 343640 558164
rect 343692 558192 343698 558204
rect 351914 558192 351920 558204
rect 343692 558164 351920 558192
rect 343692 558152 343698 558164
rect 351914 558152 351920 558164
rect 351972 558152 351978 558204
rect 283742 558084 283748 558136
rect 283800 558124 283806 558136
rect 354674 558124 354680 558136
rect 283800 558096 354680 558124
rect 283800 558084 283806 558096
rect 354674 558084 354680 558096
rect 354732 558084 354738 558136
rect 219032 558028 225000 558056
rect 219032 558016 219038 558028
rect 213144 557960 218928 557988
rect 213144 557948 213150 557960
rect 298002 557948 298008 558000
rect 298060 557988 298066 558000
rect 302142 557988 302148 558000
rect 298060 557960 302148 557988
rect 298060 557948 298066 557960
rect 302142 557948 302148 557960
rect 302200 557948 302206 558000
rect 326338 557948 326344 558000
rect 326396 557988 326402 558000
rect 335446 557988 335452 558000
rect 326396 557960 335452 557988
rect 326396 557948 326402 557960
rect 335446 557948 335452 557960
rect 335504 557948 335510 558000
rect 82814 557880 82820 557932
rect 82872 557920 82878 557932
rect 92474 557920 92480 557932
rect 82872 557892 92480 557920
rect 82872 557880 82878 557892
rect 92474 557880 92480 557892
rect 92532 557880 92538 557932
rect 93762 557880 93768 557932
rect 93820 557920 93826 557932
rect 127250 557920 127256 557932
rect 93820 557892 127256 557920
rect 93820 557880 93826 557892
rect 127250 557880 127256 557892
rect 127308 557880 127314 557932
rect 129642 557880 129648 557932
rect 129700 557920 129706 557932
rect 208578 557920 208584 557932
rect 129700 557892 208584 557920
rect 129700 557880 129706 557892
rect 208578 557880 208584 557892
rect 208636 557880 208642 557932
rect 302878 557880 302884 557932
rect 302936 557920 302942 557932
rect 317414 557920 317420 557932
rect 302936 557892 317420 557920
rect 302936 557880 302942 557892
rect 317414 557880 317420 557892
rect 317472 557880 317478 557932
rect 323578 557880 323584 557932
rect 323636 557920 323642 557932
rect 332686 557920 332692 557932
rect 323636 557892 332692 557920
rect 323636 557880 323642 557892
rect 332686 557880 332692 557892
rect 332744 557880 332750 557932
rect 79962 557812 79968 557864
rect 80020 557852 80026 557864
rect 102870 557852 102876 557864
rect 80020 557824 102876 557852
rect 80020 557812 80026 557824
rect 102870 557812 102876 557824
rect 102928 557812 102934 557864
rect 121362 557812 121368 557864
rect 121420 557852 121426 557864
rect 206094 557852 206100 557864
rect 121420 557824 206100 557852
rect 121420 557812 121426 557824
rect 206094 557812 206100 557824
rect 206152 557852 206158 557864
rect 206922 557852 206928 557864
rect 206152 557824 206928 557852
rect 206152 557812 206158 557824
rect 206922 557812 206928 557824
rect 206980 557812 206986 557864
rect 209038 557812 209044 557864
rect 209096 557852 209102 557864
rect 218974 557852 218980 557864
rect 209096 557824 218980 557852
rect 209096 557812 209102 557824
rect 218974 557812 218980 557824
rect 219032 557812 219038 557864
rect 288434 557852 288440 557864
rect 288360 557824 288440 557852
rect 288360 557796 288388 557824
rect 288434 557812 288440 557824
rect 288492 557812 288498 557864
rect 297450 557812 297456 557864
rect 297508 557852 297514 557864
rect 320174 557852 320180 557864
rect 297508 557824 320180 557852
rect 297508 557812 297514 557824
rect 320174 557812 320180 557824
rect 320232 557812 320238 557864
rect 322198 557812 322204 557864
rect 322256 557852 322262 557864
rect 331306 557852 331312 557864
rect 322256 557824 331312 557852
rect 322256 557812 322262 557824
rect 331306 557812 331312 557824
rect 331364 557812 331370 557864
rect 66162 557744 66168 557796
rect 66220 557784 66226 557796
rect 200206 557784 200212 557796
rect 66220 557756 200212 557784
rect 66220 557744 66226 557756
rect 200206 557744 200212 557756
rect 200264 557744 200270 557796
rect 202138 557744 202144 557796
rect 202196 557784 202202 557796
rect 211154 557784 211160 557796
rect 202196 557756 211160 557784
rect 202196 557744 202202 557756
rect 211154 557744 211160 557756
rect 211212 557744 211218 557796
rect 213638 557744 213644 557796
rect 213696 557784 213702 557796
rect 222102 557784 222108 557796
rect 213696 557756 222108 557784
rect 213696 557744 213702 557756
rect 222102 557744 222108 557756
rect 222160 557744 222166 557796
rect 222194 557744 222200 557796
rect 222252 557784 222258 557796
rect 229094 557784 229100 557796
rect 222252 557756 229100 557784
rect 222252 557744 222258 557756
rect 229094 557744 229100 557756
rect 229152 557744 229158 557796
rect 288342 557744 288348 557796
rect 288400 557744 288406 557796
rect 302142 557744 302148 557796
rect 302200 557784 302206 557796
rect 302234 557784 302240 557796
rect 302200 557756 302240 557784
rect 302200 557744 302206 557756
rect 302234 557744 302240 557756
rect 302292 557744 302298 557796
rect 324958 557744 324964 557796
rect 325016 557784 325022 557796
rect 334066 557784 334072 557796
rect 325016 557756 334072 557784
rect 325016 557744 325022 557756
rect 334066 557744 334072 557756
rect 334124 557744 334130 557796
rect 74994 557676 75000 557728
rect 75052 557716 75058 557728
rect 84194 557716 84200 557728
rect 75052 557688 84200 557716
rect 75052 557676 75058 557688
rect 84194 557676 84200 557688
rect 84252 557676 84258 557728
rect 93302 557676 93308 557728
rect 93360 557716 93366 557728
rect 99834 557716 99840 557728
rect 93360 557688 99840 557716
rect 93360 557676 93366 557688
rect 99834 557676 99840 557688
rect 99892 557676 99898 557728
rect 107470 557676 107476 557728
rect 107528 557716 107534 557728
rect 141510 557716 141516 557728
rect 107528 557688 141516 557716
rect 107528 557676 107534 557688
rect 141510 557676 141516 557688
rect 141568 557676 141574 557728
rect 204898 557676 204904 557728
rect 204956 557716 204962 557728
rect 213914 557716 213920 557728
rect 204956 557688 213920 557716
rect 204956 557676 204962 557688
rect 213914 557676 213920 557688
rect 213972 557676 213978 557728
rect 241606 557716 241612 557728
rect 240060 557688 241612 557716
rect 63402 557608 63408 557660
rect 63460 557648 63466 557660
rect 198734 557648 198740 557660
rect 63460 557620 198740 557648
rect 63460 557608 63466 557620
rect 198734 557608 198740 557620
rect 198792 557608 198798 557660
rect 207658 557608 207664 557660
rect 207716 557648 207722 557660
rect 217778 557648 217784 557660
rect 207716 557620 217784 557648
rect 207716 557608 207722 557620
rect 217778 557608 217784 557620
rect 217836 557608 217842 557660
rect 238662 557608 238668 557660
rect 238720 557608 238726 557660
rect 91094 557540 91100 557592
rect 91152 557580 91158 557592
rect 100018 557580 100024 557592
rect 91152 557552 100024 557580
rect 91152 557540 91158 557552
rect 100018 557540 100024 557552
rect 100076 557540 100082 557592
rect 102778 557580 102784 557592
rect 100128 557552 102784 557580
rect 99834 557472 99840 557524
rect 99892 557512 99898 557524
rect 100128 557512 100156 557552
rect 102778 557540 102784 557552
rect 102836 557540 102842 557592
rect 107746 557580 107752 557592
rect 102888 557552 107752 557580
rect 99892 557484 100156 557512
rect 99892 557472 99898 557484
rect 100570 557472 100576 557524
rect 100628 557512 100634 557524
rect 102888 557512 102916 557552
rect 107746 557540 107752 557552
rect 107804 557580 107810 557592
rect 108482 557580 108488 557592
rect 107804 557552 108488 557580
rect 107804 557540 107810 557552
rect 108482 557540 108488 557552
rect 108540 557540 108546 557592
rect 127250 557540 127256 557592
rect 127308 557580 127314 557592
rect 131758 557580 131764 557592
rect 127308 557552 131764 557580
rect 127308 557540 127314 557552
rect 131758 557540 131764 557552
rect 131816 557540 131822 557592
rect 200022 557540 200028 557592
rect 200080 557580 200086 557592
rect 200114 557580 200120 557592
rect 200080 557552 200120 557580
rect 200080 557540 200086 557552
rect 200114 557540 200120 557552
rect 200172 557540 200178 557592
rect 238680 557580 238708 557608
rect 240060 557580 240088 557688
rect 241606 557676 241612 557688
rect 241664 557676 241670 557728
rect 283650 557676 283656 557728
rect 283708 557716 283714 557728
rect 351914 557716 351920 557728
rect 283708 557688 351920 557716
rect 283708 557676 283714 557688
rect 351914 557676 351920 557688
rect 351972 557676 351978 557728
rect 251082 557608 251088 557660
rect 251140 557648 251146 557660
rect 253842 557648 253848 557660
rect 251140 557620 253848 557648
rect 251140 557608 251146 557620
rect 253842 557608 253848 557620
rect 253900 557608 253906 557660
rect 253934 557608 253940 557660
rect 253992 557648 253998 557660
rect 253992 557620 255176 557648
rect 253992 557608 253998 557620
rect 238680 557552 240088 557580
rect 255148 557580 255176 557620
rect 270402 557608 270408 557660
rect 270460 557648 270466 557660
rect 273162 557648 273168 557660
rect 270460 557620 273168 557648
rect 270460 557608 270466 557620
rect 273162 557608 273168 557620
rect 273220 557608 273226 557660
rect 273254 557608 273260 557660
rect 273312 557648 273318 557660
rect 273312 557620 274496 557648
rect 273312 557608 273318 557620
rect 260834 557580 260840 557592
rect 255148 557552 260840 557580
rect 260834 557540 260840 557552
rect 260892 557540 260898 557592
rect 274468 557580 274496 557620
rect 283558 557608 283564 557660
rect 283616 557648 283622 557660
rect 353294 557648 353300 557660
rect 283616 557620 353300 557648
rect 283616 557608 283622 557620
rect 353294 557608 353300 557620
rect 353352 557608 353358 557660
rect 282362 557580 282368 557592
rect 274468 557552 282368 557580
rect 282362 557540 282368 557552
rect 282420 557580 282426 557592
rect 288342 557580 288348 557592
rect 282420 557552 288348 557580
rect 282420 557540 282426 557552
rect 288342 557540 288348 557552
rect 288400 557540 288406 557592
rect 327718 557540 327724 557592
rect 327776 557580 327782 557592
rect 336458 557580 336464 557592
rect 327776 557552 336464 557580
rect 327776 557540 327782 557552
rect 336458 557540 336464 557552
rect 336516 557540 336522 557592
rect 100628 557484 102916 557512
rect 100628 557472 100634 557484
rect 58250 556180 58256 556232
rect 58308 556220 58314 556232
rect 580166 556220 580172 556232
rect 58308 556192 580172 556220
rect 58308 556180 58314 556192
rect 580166 556180 580172 556192
rect 580224 556180 580230 556232
rect 282362 549244 282368 549296
rect 282420 549284 282426 549296
rect 282454 549284 282460 549296
rect 282420 549256 282460 549284
rect 282420 549244 282426 549256
rect 282454 549244 282460 549256
rect 282512 549244 282518 549296
rect 77570 545708 77576 545760
rect 77628 545748 77634 545760
rect 188798 545748 188804 545760
rect 77628 545720 188804 545748
rect 77628 545708 77634 545720
rect 188798 545708 188804 545720
rect 188856 545708 188862 545760
rect 560294 545504 560300 545556
rect 560352 545544 560358 545556
rect 563146 545544 563152 545556
rect 560352 545516 563152 545544
rect 560352 545504 560358 545516
rect 563146 545504 563152 545516
rect 563204 545504 563210 545556
rect 302142 545436 302148 545488
rect 302200 545476 302206 545488
rect 309042 545476 309048 545488
rect 302200 545448 309048 545476
rect 302200 545436 302206 545448
rect 309042 545436 309048 545448
rect 309100 545436 309106 545488
rect 572622 545436 572628 545488
rect 572680 545476 572686 545488
rect 579522 545476 579528 545488
rect 572680 545448 579528 545476
rect 572680 545436 572686 545448
rect 579522 545436 579528 545448
rect 579580 545436 579586 545488
rect 115934 545368 115940 545420
rect 115992 545408 115998 545420
rect 125410 545408 125416 545420
rect 115992 545380 125416 545408
rect 115992 545368 115998 545380
rect 125410 545368 125416 545380
rect 125468 545368 125474 545420
rect 135254 545368 135260 545420
rect 135312 545408 135318 545420
rect 144822 545408 144828 545420
rect 135312 545380 144828 545408
rect 135312 545368 135318 545380
rect 144822 545368 144828 545380
rect 144880 545368 144886 545420
rect 195882 545368 195888 545420
rect 195940 545408 195946 545420
rect 201402 545408 201408 545420
rect 195940 545380 201408 545408
rect 195940 545368 195946 545380
rect 201402 545368 201408 545380
rect 201460 545368 201466 545420
rect 212534 545368 212540 545420
rect 212592 545408 212598 545420
rect 222010 545408 222016 545420
rect 212592 545380 222016 545408
rect 212592 545368 212598 545380
rect 222010 545368 222016 545380
rect 222068 545368 222074 545420
rect 231854 545368 231860 545420
rect 231912 545408 231918 545420
rect 241422 545408 241428 545420
rect 231912 545380 241428 545408
rect 231912 545368 231918 545380
rect 241422 545368 241428 545380
rect 241480 545368 241486 545420
rect 251174 545368 251180 545420
rect 251232 545408 251238 545420
rect 260742 545408 260748 545420
rect 251232 545380 260748 545408
rect 251232 545368 251238 545380
rect 260742 545368 260748 545380
rect 260800 545368 260806 545420
rect 483014 545368 483020 545420
rect 483072 545408 483078 545420
rect 485866 545408 485872 545420
rect 483072 545380 485872 545408
rect 483072 545368 483078 545380
rect 485866 545368 485872 545380
rect 485924 545368 485930 545420
rect 540974 545368 540980 545420
rect 541032 545408 541038 545420
rect 548610 545408 548616 545420
rect 541032 545380 548616 545408
rect 541032 545368 541038 545380
rect 548610 545368 548616 545380
rect 548668 545368 548674 545420
rect 85574 545300 85580 545352
rect 85632 545340 85638 545352
rect 95050 545340 95056 545352
rect 85632 545312 95056 545340
rect 85632 545300 85638 545312
rect 95050 545300 95056 545312
rect 95108 545300 95114 545352
rect 166902 545300 166908 545352
rect 166960 545340 166966 545352
rect 177298 545340 177304 545352
rect 166960 545312 177304 545340
rect 166960 545300 166966 545312
rect 177298 545300 177304 545312
rect 177356 545300 177362 545352
rect 321462 545300 321468 545352
rect 321520 545340 321526 545352
rect 328362 545340 328368 545352
rect 321520 545312 328368 545340
rect 321520 545300 321526 545312
rect 328362 545300 328368 545312
rect 328420 545300 328426 545352
rect 96614 545232 96620 545284
rect 96672 545272 96678 545284
rect 104802 545272 104808 545284
rect 96672 545244 104808 545272
rect 96672 545232 96678 545244
rect 104802 545232 104808 545244
rect 104860 545232 104866 545284
rect 57606 545028 57612 545080
rect 57664 545068 57670 545080
rect 112806 545068 112812 545080
rect 57664 545040 112812 545068
rect 57664 545028 57670 545040
rect 112806 545028 112812 545040
rect 112864 545028 112870 545080
rect 114922 545028 114928 545080
rect 114980 545068 114986 545080
rect 202138 545068 202144 545080
rect 114980 545040 202144 545068
rect 114980 545028 114986 545040
rect 202138 545028 202144 545040
rect 202196 545028 202202 545080
rect 89622 544960 89628 545012
rect 89680 545000 89686 545012
rect 177206 545000 177212 545012
rect 89680 544972 177212 545000
rect 89680 544960 89686 544972
rect 177206 544960 177212 544972
rect 177264 544960 177270 545012
rect 92382 544892 92388 544944
rect 92440 544932 92446 544944
rect 181346 544932 181352 544944
rect 92440 544904 181352 544932
rect 92440 544892 92446 544904
rect 181346 544892 181352 544904
rect 181404 544892 181410 544944
rect 96246 544824 96252 544876
rect 96304 544864 96310 544876
rect 188338 544864 188344 544876
rect 96304 544836 188344 544864
rect 96304 544824 96310 544836
rect 188338 544824 188344 544836
rect 188396 544824 188402 544876
rect 91002 544756 91008 544808
rect 91060 544796 91066 544808
rect 179230 544796 179236 544808
rect 91060 544768 179236 544796
rect 91060 544756 91066 544768
rect 179230 544756 179236 544768
rect 179288 544756 179294 544808
rect 96522 544688 96528 544740
rect 96580 544728 96586 544740
rect 189626 544728 189632 544740
rect 96580 544700 189632 544728
rect 96580 544688 96586 544700
rect 189626 544688 189632 544700
rect 189684 544688 189690 544740
rect 94130 544620 94136 544672
rect 94188 544660 94194 544672
rect 188430 544660 188436 544672
rect 94188 544632 188436 544660
rect 94188 544620 94194 544632
rect 188430 544620 188436 544632
rect 188488 544620 188494 544672
rect 89990 544552 89996 544604
rect 90048 544592 90054 544604
rect 188614 544592 188620 544604
rect 90048 544564 188620 544592
rect 90048 544552 90054 544564
rect 188614 544552 188620 544564
rect 188672 544552 188678 544604
rect 57054 544484 57060 544536
rect 57112 544524 57118 544536
rect 102502 544524 102508 544536
rect 57112 544496 102508 544524
rect 57112 544484 57118 544496
rect 102502 544484 102508 544496
rect 102560 544484 102566 544536
rect 103422 544484 103428 544536
rect 103480 544524 103486 544536
rect 202046 544524 202052 544536
rect 103480 544496 202052 544524
rect 103480 544484 103486 544496
rect 202046 544484 202052 544496
rect 202104 544484 202110 544536
rect 57422 544416 57428 544468
rect 57480 544456 57486 544468
rect 108666 544456 108672 544468
rect 57480 544428 108672 544456
rect 57480 544416 57486 544428
rect 108666 544416 108672 544428
rect 108724 544416 108730 544468
rect 110322 544416 110328 544468
rect 110380 544456 110386 544468
rect 212166 544456 212172 544468
rect 110380 544428 212172 544456
rect 110380 544416 110386 544428
rect 212166 544416 212172 544428
rect 212224 544416 212230 544468
rect 81710 544348 81716 544400
rect 81768 544388 81774 544400
rect 195974 544388 195980 544400
rect 81768 544360 195980 544388
rect 81768 544348 81774 544360
rect 195974 544348 195980 544360
rect 196032 544348 196038 544400
rect 86862 544280 86868 544332
rect 86920 544320 86926 544332
rect 173066 544320 173072 544332
rect 86920 544292 173072 544320
rect 86920 544280 86926 544292
rect 173066 544280 173072 544292
rect 173124 544280 173130 544332
rect 88242 544212 88248 544264
rect 88300 544252 88306 544264
rect 175090 544252 175096 544264
rect 88300 544224 175096 544252
rect 88300 544212 88306 544224
rect 175090 544212 175096 544224
rect 175148 544212 175154 544264
rect 86770 544144 86776 544196
rect 86828 544184 86834 544196
rect 170950 544184 170956 544196
rect 86828 544156 170956 544184
rect 86828 544144 86834 544156
rect 170950 544144 170956 544156
rect 171008 544144 171014 544196
rect 85482 544076 85488 544128
rect 85540 544116 85546 544128
rect 168834 544116 168840 544128
rect 85540 544088 168840 544116
rect 85540 544076 85546 544088
rect 168834 544076 168840 544088
rect 168892 544076 168898 544128
rect 73062 544008 73068 544060
rect 73120 544048 73126 544060
rect 148134 544048 148140 544060
rect 73120 544020 148140 544048
rect 73120 544008 73126 544020
rect 148134 544008 148140 544020
rect 148192 544008 148198 544060
rect 102870 543940 102876 543992
rect 102928 543980 102934 543992
rect 160554 543980 160560 543992
rect 102928 543952 160560 543980
rect 102928 543940 102934 543952
rect 160554 543940 160560 543952
rect 160612 543940 160618 543992
rect 57514 543872 57520 543924
rect 57572 543912 57578 543924
rect 110782 543912 110788 543924
rect 57572 543884 110788 543912
rect 57572 543872 57578 543884
rect 110782 543872 110788 543884
rect 110840 543872 110846 543924
rect 57330 543804 57336 543856
rect 57388 543844 57394 543856
rect 106642 543844 106648 543856
rect 57388 543816 106648 543844
rect 57388 543804 57394 543816
rect 106642 543804 106648 543816
rect 106700 543804 106706 543856
rect 57238 543736 57244 543788
rect 57296 543776 57302 543788
rect 104526 543776 104532 543788
rect 57296 543748 104532 543776
rect 57296 543736 57302 543748
rect 104526 543736 104532 543748
rect 104584 543736 104590 543788
rect 429378 543736 429384 543788
rect 429436 543776 429442 543788
rect 429436 543748 429516 543776
rect 429436 543736 429442 543748
rect 429488 543720 429516 543748
rect 71682 543668 71688 543720
rect 71740 543708 71746 543720
rect 75454 543708 75460 543720
rect 71740 543680 75460 543708
rect 71740 543668 71746 543680
rect 75454 543668 75460 543680
rect 75512 543668 75518 543720
rect 75822 543668 75828 543720
rect 75880 543708 75886 543720
rect 152274 543708 152280 543720
rect 75880 543680 152280 543708
rect 75880 543668 75886 543680
rect 152274 543668 152280 543680
rect 152332 543668 152338 543720
rect 152458 543668 152464 543720
rect 152516 543708 152522 543720
rect 166810 543708 166816 543720
rect 152516 543680 166816 543708
rect 152516 543668 152522 543680
rect 166810 543668 166816 543680
rect 166868 543668 166874 543720
rect 206922 543668 206928 543720
rect 206980 543708 206986 543720
rect 220446 543708 220452 543720
rect 206980 543680 220452 543708
rect 206980 543668 206986 543680
rect 220446 543668 220452 543680
rect 220504 543668 220510 543720
rect 229002 543668 229008 543720
rect 229060 543708 229066 543720
rect 260190 543708 260196 543720
rect 229060 543680 260196 543708
rect 229060 543668 229066 543680
rect 260190 543668 260196 543680
rect 260248 543668 260254 543720
rect 429470 543668 429476 543720
rect 429528 543668 429534 543720
rect 78582 543600 78588 543652
rect 78640 543640 78646 543652
rect 156414 543640 156420 543652
rect 78640 543612 156420 543640
rect 78640 543600 78646 543612
rect 156414 543600 156420 543612
rect 156472 543600 156478 543652
rect 205542 543600 205548 543652
rect 205600 543640 205606 543652
rect 218698 543640 218704 543652
rect 205600 543612 218704 543640
rect 205600 543600 205606 543612
rect 218698 543600 218704 543612
rect 218756 543600 218762 543652
rect 227622 543600 227628 543652
rect 227680 543640 227686 543652
rect 258074 543640 258080 543652
rect 227680 543612 258080 543640
rect 227680 543600 227686 543612
rect 258074 543600 258080 543612
rect 258132 543600 258138 543652
rect 61010 543532 61016 543584
rect 61068 543572 61074 543584
rect 62022 543572 62028 543584
rect 61068 543544 62028 543572
rect 61068 543532 61074 543544
rect 62022 543532 62028 543544
rect 62080 543532 62086 543584
rect 70210 543532 70216 543584
rect 70268 543572 70274 543584
rect 71314 543572 71320 543584
rect 70268 543544 71320 543572
rect 70268 543532 70274 543544
rect 71314 543532 71320 543544
rect 71372 543532 71378 543584
rect 82722 543532 82728 543584
rect 82780 543572 82786 543584
rect 164694 543572 164700 543584
rect 82780 543544 164700 543572
rect 82780 543532 82786 543544
rect 164694 543532 164700 543544
rect 164752 543532 164758 543584
rect 208302 543532 208308 543584
rect 208360 543572 208366 543584
rect 222838 543572 222844 543584
rect 208360 543544 222844 543572
rect 208360 543532 208366 543544
rect 222838 543532 222844 543544
rect 222896 543532 222902 543584
rect 230382 543532 230388 543584
rect 230440 543572 230446 543584
rect 262214 543572 262220 543584
rect 230440 543544 262220 543572
rect 230440 543532 230446 543544
rect 262214 543532 262220 543544
rect 262272 543532 262278 543584
rect 127342 543464 127348 543516
rect 127400 543504 127406 543516
rect 209038 543504 209044 543516
rect 127400 543476 209044 543504
rect 127400 543464 127406 543476
rect 209038 543464 209044 543476
rect 209096 543464 209102 543516
rect 209682 543464 209688 543516
rect 209740 543504 209746 543516
rect 224494 543504 224500 543516
rect 209740 543476 224500 543504
rect 209740 543464 209746 543476
rect 224494 543464 224500 543476
rect 224552 543464 224558 543516
rect 231762 543464 231768 543516
rect 231820 543504 231826 543516
rect 264330 543504 264336 543516
rect 231820 543476 264336 543504
rect 231820 543464 231826 543476
rect 264330 543464 264336 543476
rect 264388 543464 264394 543516
rect 123202 543396 123208 543448
rect 123260 543436 123266 543448
rect 207658 543436 207664 543448
rect 123260 543408 207664 543436
rect 123260 543396 123266 543408
rect 207658 543396 207664 543408
rect 207716 543396 207722 543448
rect 211062 543396 211068 543448
rect 211120 543436 211126 543448
rect 226978 543436 226984 543448
rect 211120 543408 226984 543436
rect 211120 543396 211126 543408
rect 226978 543396 226984 543408
rect 227036 543396 227042 543448
rect 233142 543396 233148 543448
rect 233200 543436 233206 543448
rect 266446 543436 266452 543448
rect 233200 543408 266452 543436
rect 233200 543396 233206 543408
rect 266446 543396 266452 543408
rect 266504 543396 266510 543448
rect 119062 543328 119068 543380
rect 119120 543368 119126 543380
rect 204898 543368 204904 543380
rect 119120 543340 204904 543368
rect 119120 543328 119126 543340
rect 204898 543328 204904 543340
rect 204956 543328 204962 543380
rect 212442 543328 212448 543380
rect 212500 543368 212506 543380
rect 231118 543368 231124 543380
rect 212500 543340 231124 543368
rect 212500 543328 212506 543340
rect 231118 543328 231124 543340
rect 231176 543328 231182 543380
rect 233050 543328 233056 543380
rect 233108 543368 233114 543380
rect 268470 543368 268476 543380
rect 233108 543340 268476 543368
rect 233108 543328 233114 543340
rect 268470 543328 268476 543340
rect 268528 543328 268534 543380
rect 117038 543260 117044 543312
rect 117096 543300 117102 543312
rect 203518 543300 203524 543312
rect 117096 543272 203524 543300
rect 117096 543260 117102 543272
rect 203518 543260 203524 543272
rect 203576 543260 203582 543312
rect 215202 543260 215208 543312
rect 215260 543300 215266 543312
rect 235258 543300 235264 543312
rect 215260 543272 235264 543300
rect 215260 543260 215266 543272
rect 235258 543260 235264 543272
rect 235316 543260 235322 543312
rect 235902 543260 235908 543312
rect 235960 543300 235966 543312
rect 272610 543300 272616 543312
rect 235960 543272 272616 543300
rect 235960 543260 235966 543272
rect 272610 543260 272616 543272
rect 272668 543260 272674 543312
rect 93670 543192 93676 543244
rect 93728 543232 93734 543244
rect 183370 543232 183376 543244
rect 93728 543204 183376 543232
rect 93728 543192 93734 543204
rect 183370 543192 183376 543204
rect 183428 543192 183434 543244
rect 210970 543192 210976 543244
rect 211028 543232 211034 543244
rect 229094 543232 229100 543244
rect 211028 543204 229100 543232
rect 211028 543192 211034 543204
rect 229094 543192 229100 543204
rect 229152 543192 229158 543244
rect 234522 543192 234528 543244
rect 234580 543232 234586 543244
rect 270586 543232 270592 543244
rect 234580 543204 270592 543232
rect 234580 543192 234586 543204
rect 270586 543192 270592 543204
rect 270644 543192 270650 543244
rect 56962 543124 56968 543176
rect 57020 543164 57026 543176
rect 79686 543164 79692 543176
rect 57020 543136 79692 543164
rect 57020 543124 57026 543136
rect 79686 543124 79692 543136
rect 79744 543124 79750 543176
rect 95142 543124 95148 543176
rect 95200 543164 95206 543176
rect 187510 543164 187516 543176
rect 95200 543136 187516 543164
rect 95200 543124 95206 543136
rect 187510 543124 187516 543136
rect 187568 543124 187574 543176
rect 204162 543124 204168 543176
rect 204220 543164 204226 543176
rect 216214 543164 216220 543176
rect 204220 543136 216220 543164
rect 204220 543124 204226 543136
rect 216214 543124 216220 543136
rect 216272 543124 216278 543176
rect 216582 543124 216588 543176
rect 216640 543164 216646 543176
rect 237374 543164 237380 543176
rect 216640 543136 237380 543164
rect 216640 543124 216646 543136
rect 237374 543124 237380 543136
rect 237432 543124 237438 543176
rect 238662 543124 238668 543176
rect 238720 543164 238726 543176
rect 276750 543164 276756 543176
rect 238720 543136 276756 543164
rect 238720 543124 238726 543136
rect 276750 543124 276756 543136
rect 276808 543124 276814 543176
rect 67542 543056 67548 543108
rect 67600 543096 67606 543108
rect 98362 543096 98368 543108
rect 67600 543068 98368 543096
rect 67600 543056 67606 543068
rect 98362 543056 98368 543068
rect 98420 543056 98426 543108
rect 99282 543056 99288 543108
rect 99340 543096 99346 543108
rect 193766 543096 193772 543108
rect 99340 543068 193772 543096
rect 99340 543056 99346 543068
rect 193766 543056 193772 543068
rect 193824 543056 193830 543108
rect 213822 543056 213828 543108
rect 213880 543096 213886 543108
rect 233234 543096 233240 543108
rect 213880 543068 233240 543096
rect 213880 543056 213886 543068
rect 233234 543056 233240 543068
rect 233292 543056 233298 543108
rect 237282 543056 237288 543108
rect 237340 543096 237346 543108
rect 274726 543096 274732 543108
rect 237340 543068 274732 543096
rect 237340 543056 237346 543068
rect 274726 543056 274732 543068
rect 274784 543056 274790 543108
rect 57146 542988 57152 543040
rect 57204 543028 57210 543040
rect 100386 543028 100392 543040
rect 57204 543000 100392 543028
rect 57204 542988 57210 543000
rect 100386 542988 100392 543000
rect 100444 542988 100450 543040
rect 102042 542988 102048 543040
rect 102100 543028 102106 543040
rect 197906 543028 197912 543040
rect 102100 543000 197912 543028
rect 102100 542988 102106 543000
rect 197906 542988 197912 543000
rect 197964 542988 197970 543040
rect 202782 542988 202788 543040
rect 202840 543028 202846 543040
rect 214558 543028 214564 543040
rect 202840 543000 214564 543028
rect 202840 542988 202846 543000
rect 214558 542988 214564 543000
rect 214616 542988 214622 543040
rect 217870 542988 217876 543040
rect 217928 543028 217934 543040
rect 239398 543028 239404 543040
rect 217928 543000 239404 543028
rect 217928 542988 217934 543000
rect 239398 542988 239404 543000
rect 239456 542988 239462 543040
rect 240042 542988 240048 543040
rect 240100 543028 240106 543040
rect 278866 543028 278872 543040
rect 240100 543000 278872 543028
rect 240100 542988 240106 543000
rect 278866 542988 278872 543000
rect 278924 542988 278930 543040
rect 104158 542920 104164 542972
rect 104216 542960 104222 542972
rect 137738 542960 137744 542972
rect 104216 542932 137744 542960
rect 104216 542920 104222 542932
rect 137738 542920 137744 542932
rect 137796 542920 137802 542972
rect 204162 542960 204168 542972
rect 139964 542932 204168 542960
rect 70302 542852 70308 542904
rect 70360 542892 70366 542904
rect 73430 542892 73436 542904
rect 70360 542864 73436 542892
rect 70360 542852 70366 542864
rect 73430 542852 73436 542864
rect 73488 542852 73494 542904
rect 105538 542852 105544 542904
rect 105596 542892 105602 542904
rect 139854 542892 139860 542904
rect 105596 542864 139860 542892
rect 105596 542852 105602 542864
rect 139854 542852 139860 542864
rect 139912 542852 139918 542904
rect 100018 542784 100024 542836
rect 100076 542824 100082 542836
rect 131482 542824 131488 542836
rect 100076 542796 131488 542824
rect 100076 542784 100082 542796
rect 131482 542784 131488 542796
rect 131540 542784 131546 542836
rect 133138 542784 133144 542836
rect 133196 542824 133202 542836
rect 133196 542796 135852 542824
rect 133196 542784 133202 542796
rect 102778 542716 102784 542768
rect 102836 542756 102842 542768
rect 135714 542756 135720 542768
rect 102836 542728 135720 542756
rect 102836 542716 102842 542728
rect 135714 542716 135720 542728
rect 135772 542716 135778 542768
rect 135824 542756 135852 542796
rect 137370 542784 137376 542836
rect 137428 542824 137434 542836
rect 139964 542824 139992 542932
rect 204162 542920 204168 542932
rect 204220 542920 204226 542972
rect 226242 542920 226248 542972
rect 226300 542960 226306 542972
rect 256050 542960 256056 542972
rect 226300 542932 256056 542960
rect 226300 542920 226306 542932
rect 256050 542920 256056 542932
rect 256108 542920 256114 542972
rect 140038 542852 140044 542904
rect 140096 542892 140102 542904
rect 200022 542892 200028 542904
rect 140096 542864 200028 542892
rect 140096 542852 140102 542864
rect 200022 542852 200028 542864
rect 200080 542852 200086 542904
rect 226150 542852 226156 542904
rect 226208 542892 226214 542904
rect 253934 542892 253940 542904
rect 226208 542864 253940 542892
rect 226208 542852 226214 542864
rect 253934 542852 253940 542864
rect 253992 542852 253998 542904
rect 191742 542824 191748 542836
rect 137428 542796 139992 542824
rect 140056 542796 191748 542824
rect 137428 542784 137434 542796
rect 140056 542756 140084 542796
rect 191742 542784 191748 542796
rect 191800 542784 191806 542836
rect 223482 542784 223488 542836
rect 223540 542824 223546 542836
rect 249794 542824 249800 542836
rect 223540 542796 249800 542824
rect 223540 542784 223546 542796
rect 249794 542784 249800 542796
rect 249852 542784 249858 542836
rect 135824 542728 140084 542756
rect 140130 542716 140136 542768
rect 140188 542756 140194 542768
rect 195882 542756 195888 542768
rect 140188 542728 195888 542756
rect 140188 542716 140194 542728
rect 195882 542716 195888 542728
rect 195940 542716 195946 542768
rect 224862 542716 224868 542768
rect 224920 542756 224926 542768
rect 251910 542756 251916 542768
rect 224920 542728 251916 542756
rect 224920 542716 224926 542728
rect 251910 542716 251916 542728
rect 251968 542716 251974 542768
rect 131758 542648 131764 542700
rect 131816 542688 131822 542700
rect 185486 542688 185492 542700
rect 131816 542660 185492 542688
rect 131816 542648 131822 542660
rect 185486 542648 185492 542660
rect 185544 542648 185550 542700
rect 222102 542648 222108 542700
rect 222160 542688 222166 542700
rect 247770 542688 247776 542700
rect 222160 542660 247776 542688
rect 222160 542648 222166 542660
rect 247770 542648 247776 542660
rect 247828 542648 247834 542700
rect 108298 542580 108304 542632
rect 108356 542620 108362 542632
rect 146018 542620 146024 542632
rect 108356 542592 146024 542620
rect 108356 542580 108362 542592
rect 146018 542580 146024 542592
rect 146076 542580 146082 542632
rect 162670 542620 162676 542632
rect 146128 542592 162676 542620
rect 65150 542512 65156 542564
rect 65208 542552 65214 542564
rect 66162 542552 66168 542564
rect 65208 542524 66168 542552
rect 65208 542512 65214 542524
rect 66162 542512 66168 542524
rect 66220 542512 66226 542564
rect 108482 542512 108488 542564
rect 108540 542552 108546 542564
rect 143994 542552 144000 542564
rect 108540 542524 144000 542552
rect 108540 542512 108546 542524
rect 143994 542512 144000 542524
rect 144052 542512 144058 542564
rect 145558 542512 145564 542564
rect 145616 542552 145622 542564
rect 146128 542552 146156 542592
rect 162670 542580 162676 542592
rect 162728 542580 162734 542632
rect 220722 542580 220728 542632
rect 220780 542620 220786 542632
rect 245654 542620 245660 542632
rect 220780 542592 245660 542620
rect 220780 542580 220786 542592
rect 245654 542580 245660 542592
rect 245712 542580 245718 542632
rect 145616 542524 146156 542552
rect 145616 542512 145622 542524
rect 148318 542512 148324 542564
rect 148376 542552 148382 542564
rect 158530 542552 158536 542564
rect 148376 542524 158536 542552
rect 148376 542512 148382 542524
rect 158530 542512 158536 542524
rect 158588 542512 158594 542564
rect 217962 542512 217968 542564
rect 218020 542552 218026 542564
rect 241514 542552 241520 542564
rect 218020 542524 241520 542552
rect 218020 542512 218026 542524
rect 241514 542512 241520 542524
rect 241572 542512 241578 542564
rect 106918 542444 106924 542496
rect 106976 542484 106982 542496
rect 141878 542484 141884 542496
rect 106976 542456 141884 542484
rect 106976 542444 106982 542456
rect 141878 542444 141884 542456
rect 141936 542444 141942 542496
rect 154390 542484 154396 542496
rect 141988 542456 154396 542484
rect 101398 542376 101404 542428
rect 101456 542416 101462 542428
rect 133598 542416 133604 542428
rect 101456 542388 133604 542416
rect 101456 542376 101462 542388
rect 133598 542376 133604 542388
rect 133656 542376 133662 542428
rect 135898 542376 135904 542428
rect 135956 542416 135962 542428
rect 135956 542388 141372 542416
rect 135956 542376 135962 542388
rect 141344 542348 141372 542388
rect 141418 542376 141424 542428
rect 141476 542416 141482 542428
rect 141988 542416 142016 542456
rect 154390 542444 154396 542456
rect 154448 542444 154454 542496
rect 219342 542444 219348 542496
rect 219400 542484 219406 542496
rect 243538 542484 243544 542496
rect 219400 542456 243544 542484
rect 219400 542444 219406 542456
rect 243538 542444 243544 542456
rect 243596 542444 243602 542496
rect 150158 542416 150164 542428
rect 141476 542388 142016 542416
rect 142080 542388 150164 542416
rect 141476 542376 141482 542388
rect 142080 542348 142108 542388
rect 150158 542376 150164 542388
rect 150216 542376 150222 542428
rect 141344 542320 142108 542348
rect 429378 540948 429384 541000
rect 429436 540988 429442 541000
rect 429470 540988 429476 541000
rect 429436 540960 429476 540988
rect 429436 540948 429442 540960
rect 429470 540948 429476 540960
rect 429528 540948 429534 541000
rect 56870 540812 56876 540864
rect 56928 540852 56934 540864
rect 137278 540852 137284 540864
rect 56928 540824 137284 540852
rect 56928 540812 56934 540824
rect 137278 540812 137284 540824
rect 137336 540812 137342 540864
rect 56778 540744 56784 540796
rect 56836 540784 56842 540796
rect 170030 540784 170036 540796
rect 56836 540756 170036 540784
rect 56836 540744 56842 540756
rect 170030 540744 170036 540756
rect 170088 540744 170094 540796
rect 56962 540676 56968 540728
rect 57020 540716 57026 540728
rect 299750 540716 299756 540728
rect 57020 540688 299756 540716
rect 57020 540676 57026 540688
rect 299750 540676 299756 540688
rect 299808 540676 299814 540728
rect 59906 540608 59912 540660
rect 59964 540648 59970 540660
rect 429378 540648 429384 540660
rect 59964 540620 429384 540648
rect 59964 540608 59970 540620
rect 429378 540608 429384 540620
rect 429436 540608 429442 540660
rect 57974 540540 57980 540592
rect 58032 540580 58038 540592
rect 462314 540580 462320 540592
rect 58032 540552 462320 540580
rect 58032 540540 58038 540552
rect 462314 540540 462320 540552
rect 462372 540540 462378 540592
rect 59814 540472 59820 540524
rect 59872 540512 59878 540524
rect 491754 540512 491760 540524
rect 59872 540484 491760 540512
rect 59872 540472 59878 540484
rect 491754 540472 491760 540484
rect 491812 540472 491818 540524
rect 59722 540404 59728 540456
rect 59780 540444 59786 540456
rect 580350 540444 580356 540456
rect 59780 540416 580356 540444
rect 59780 540404 59786 540416
rect 580350 540404 580356 540416
rect 580408 540404 580414 540456
rect 59630 540336 59636 540388
rect 59688 540376 59694 540388
rect 580718 540376 580724 540388
rect 59688 540348 580724 540376
rect 59688 540336 59694 540348
rect 580718 540336 580724 540348
rect 580776 540336 580782 540388
rect 58066 540268 58072 540320
rect 58124 540308 58130 540320
rect 580258 540308 580264 540320
rect 58124 540280 580264 540308
rect 58124 540268 58130 540280
rect 580258 540268 580264 540280
rect 580316 540268 580322 540320
rect 58158 540200 58164 540252
rect 58216 540240 58222 540252
rect 580442 540240 580448 540252
rect 58216 540212 580448 540240
rect 58216 540200 58222 540212
rect 580442 540200 580448 540212
rect 580500 540200 580506 540252
rect 59538 539724 59544 539776
rect 59596 539764 59602 539776
rect 580902 539764 580908 539776
rect 59596 539736 580908 539764
rect 59596 539724 59602 539736
rect 580902 539724 580908 539736
rect 580960 539724 580966 539776
rect 57606 539656 57612 539708
rect 57664 539696 57670 539708
rect 580534 539696 580540 539708
rect 57664 539668 580540 539696
rect 57664 539656 57670 539668
rect 580534 539656 580540 539668
rect 580592 539656 580598 539708
rect 57514 539588 57520 539640
rect 57572 539628 57578 539640
rect 580810 539628 580816 539640
rect 57572 539600 580816 539628
rect 57572 539588 57578 539600
rect 580810 539588 580816 539600
rect 580868 539588 580874 539640
rect 57146 539180 57152 539232
rect 57204 539220 57210 539232
rect 580258 539220 580264 539232
rect 57204 539192 580264 539220
rect 57204 539180 57210 539192
rect 580258 539180 580264 539192
rect 580316 539180 580322 539232
rect 33778 538228 33784 538280
rect 33836 538268 33842 538280
rect 57422 538268 57428 538280
rect 33836 538240 57428 538268
rect 33836 538228 33842 538240
rect 57422 538228 57428 538240
rect 57480 538228 57486 538280
rect 19978 536800 19984 536852
rect 20036 536840 20042 536852
rect 57422 536840 57428 536852
rect 20036 536812 57428 536840
rect 20036 536800 20042 536812
rect 57422 536800 57428 536812
rect 57480 536800 57486 536852
rect 17218 534080 17224 534132
rect 17276 534120 17282 534132
rect 57422 534120 57428 534132
rect 17276 534092 57428 534120
rect 17276 534080 17282 534092
rect 57422 534080 57428 534092
rect 57480 534080 57486 534132
rect 28258 532720 28264 532772
rect 28316 532760 28322 532772
rect 57422 532760 57428 532772
rect 28316 532732 57428 532760
rect 28316 532720 28322 532732
rect 57422 532720 57428 532732
rect 57480 532720 57486 532772
rect 48958 531360 48964 531412
rect 49016 531400 49022 531412
rect 57422 531400 57428 531412
rect 49016 531372 57428 531400
rect 49016 531360 49022 531372
rect 57422 531360 57428 531372
rect 57480 531360 57486 531412
rect 4798 528572 4804 528624
rect 4856 528612 4862 528624
rect 57422 528612 57428 528624
rect 4856 528584 57428 528612
rect 4856 528572 4862 528584
rect 57422 528572 57428 528584
rect 57480 528572 57486 528624
rect 53098 527144 53104 527196
rect 53156 527184 53162 527196
rect 57422 527184 57428 527196
rect 53156 527156 57428 527184
rect 53156 527144 53162 527156
rect 57422 527144 57428 527156
rect 57480 527144 57486 527196
rect 46198 524424 46204 524476
rect 46256 524464 46262 524476
rect 57422 524464 57428 524476
rect 46256 524436 57428 524464
rect 46256 524424 46262 524436
rect 57422 524424 57428 524436
rect 57480 524424 57486 524476
rect 282546 524424 282552 524476
rect 282604 524424 282610 524476
rect 282564 524328 282592 524424
rect 282638 524328 282644 524340
rect 282564 524300 282644 524328
rect 282638 524288 282644 524300
rect 282696 524288 282702 524340
rect 4890 522996 4896 523048
rect 4948 523036 4954 523048
rect 57422 523036 57428 523048
rect 4948 523008 57428 523036
rect 4948 522996 4954 523008
rect 57422 522996 57428 523008
rect 57480 522996 57486 523048
rect 51718 521704 51724 521756
rect 51776 521744 51782 521756
rect 57422 521744 57428 521756
rect 51776 521716 57428 521744
rect 51776 521704 51782 521716
rect 57422 521704 57428 521716
rect 57480 521704 57486 521756
rect 43438 518916 43444 518968
rect 43496 518956 43502 518968
rect 57422 518956 57428 518968
rect 43496 518928 57428 518956
rect 43496 518916 43502 518928
rect 57422 518916 57428 518928
rect 57480 518916 57486 518968
rect 4982 517488 4988 517540
rect 5040 517528 5046 517540
rect 57422 517528 57428 517540
rect 5040 517500 57428 517528
rect 5040 517488 5046 517500
rect 57422 517488 57428 517500
rect 57480 517488 57486 517540
rect 50338 514768 50344 514820
rect 50396 514808 50402 514820
rect 57422 514808 57428 514820
rect 50396 514780 57428 514808
rect 50396 514768 50402 514780
rect 57422 514768 57428 514780
rect 57480 514768 57486 514820
rect 282546 514768 282552 514820
rect 282604 514768 282610 514820
rect 282564 514740 282592 514768
rect 282638 514740 282644 514752
rect 282564 514712 282644 514740
rect 282638 514700 282644 514712
rect 282696 514700 282702 514752
rect 35158 513340 35164 513392
rect 35216 513380 35222 513392
rect 57422 513380 57428 513392
rect 35216 513352 57428 513380
rect 35216 513340 35222 513352
rect 57422 513340 57428 513352
rect 57480 513340 57486 513392
rect 5074 511980 5080 512032
rect 5132 512020 5138 512032
rect 57422 512020 57428 512032
rect 5132 511992 57428 512020
rect 5132 511980 5138 511992
rect 57422 511980 57428 511992
rect 57480 511980 57486 512032
rect 282546 511980 282552 512032
rect 282604 512020 282610 512032
rect 282638 512020 282644 512032
rect 282604 511992 282644 512020
rect 282604 511980 282610 511992
rect 282638 511980 282644 511992
rect 282696 511980 282702 512032
rect 39390 509260 39396 509312
rect 39448 509300 39454 509312
rect 57422 509300 57428 509312
rect 39448 509272 57428 509300
rect 39448 509260 39454 509272
rect 57422 509260 57428 509272
rect 57480 509260 57486 509312
rect 33870 507832 33876 507884
rect 33928 507872 33934 507884
rect 57422 507872 57428 507884
rect 33928 507844 57428 507872
rect 33928 507832 33934 507844
rect 57422 507832 57428 507844
rect 57480 507832 57486 507884
rect 282546 505112 282552 505164
rect 282604 505112 282610 505164
rect 282564 505016 282592 505112
rect 282638 505016 282644 505028
rect 282564 504988 282644 505016
rect 282638 504976 282644 504988
rect 282696 504976 282702 505028
rect 37918 503684 37924 503736
rect 37976 503724 37982 503736
rect 57422 503724 57428 503736
rect 37976 503696 57428 503724
rect 37976 503684 37982 503696
rect 57422 503684 57428 503696
rect 57480 503684 57486 503736
rect 28350 502324 28356 502376
rect 28408 502364 28414 502376
rect 57422 502364 57428 502376
rect 28408 502336 57428 502364
rect 28408 502324 28414 502336
rect 57422 502324 57428 502336
rect 57480 502324 57486 502376
rect 32398 498176 32404 498228
rect 32456 498216 32462 498228
rect 57422 498216 57428 498228
rect 32456 498188 57428 498216
rect 32456 498176 32462 498188
rect 57422 498176 57428 498188
rect 57480 498176 57486 498228
rect 282362 497496 282368 497548
rect 282420 497536 282426 497548
rect 282546 497536 282552 497548
rect 282420 497508 282552 497536
rect 282420 497496 282426 497508
rect 282546 497496 282552 497508
rect 282604 497496 282610 497548
rect 3970 495456 3976 495508
rect 4028 495496 4034 495508
rect 5166 495496 5172 495508
rect 4028 495468 5172 495496
rect 4028 495456 4034 495468
rect 5166 495456 5172 495468
rect 5224 495456 5230 495508
rect 20070 495456 20076 495508
rect 20128 495496 20134 495508
rect 57422 495496 57428 495508
rect 20128 495468 57428 495496
rect 20128 495456 20134 495468
rect 57422 495456 57428 495468
rect 57480 495456 57486 495508
rect 15838 489880 15844 489932
rect 15896 489920 15902 489932
rect 56686 489920 56692 489932
rect 15896 489892 56692 489920
rect 15896 489880 15902 489892
rect 56686 489880 56692 489892
rect 56744 489880 56750 489932
rect 3970 485800 3976 485852
rect 4028 485840 4034 485852
rect 56686 485840 56692 485852
rect 4028 485812 56692 485840
rect 4028 485800 4034 485812
rect 56686 485800 56692 485812
rect 56744 485800 56750 485852
rect 282546 485800 282552 485852
rect 282604 485800 282610 485852
rect 282564 485704 282592 485800
rect 282638 485704 282644 485716
rect 282564 485676 282644 485704
rect 282638 485664 282644 485676
rect 282696 485664 282702 485716
rect 3878 484372 3884 484424
rect 3936 484412 3942 484424
rect 56686 484412 56692 484424
rect 3936 484384 56692 484412
rect 3936 484372 3942 484384
rect 56686 484372 56692 484384
rect 56744 484372 56750 484424
rect 282362 482944 282368 482996
rect 282420 482984 282426 482996
rect 282638 482984 282644 482996
rect 282420 482956 282644 482984
rect 282420 482944 282426 482956
rect 282638 482944 282644 482956
rect 282696 482944 282702 482996
rect 56686 481720 56692 481772
rect 56744 481760 56750 481772
rect 56744 481732 56824 481760
rect 56744 481720 56750 481732
rect 5166 481584 5172 481636
rect 5224 481624 5230 481636
rect 56686 481624 56692 481636
rect 5224 481596 56692 481624
rect 5224 481584 5230 481596
rect 56686 481584 56692 481596
rect 56744 481584 56750 481636
rect 56686 481108 56692 481160
rect 56744 481148 56750 481160
rect 56796 481148 56824 481732
rect 56744 481120 56824 481148
rect 56744 481108 56750 481120
rect 2866 480156 2872 480208
rect 2924 480196 2930 480208
rect 56502 480196 56508 480208
rect 2924 480168 56508 480196
rect 2924 480156 2930 480168
rect 56502 480156 56508 480168
rect 56560 480156 56566 480208
rect 4062 477436 4068 477488
rect 4120 477476 4126 477488
rect 56502 477476 56508 477488
rect 4120 477448 56508 477476
rect 4120 477436 4126 477448
rect 56502 477436 56508 477448
rect 56560 477436 56566 477488
rect 3694 476008 3700 476060
rect 3752 476048 3758 476060
rect 56502 476048 56508 476060
rect 3752 476020 56508 476048
rect 3752 476008 3758 476020
rect 56502 476008 56508 476020
rect 56560 476008 56566 476060
rect 3786 474648 3792 474700
rect 3844 474688 3850 474700
rect 56502 474688 56508 474700
rect 3844 474660 56508 474688
rect 3844 474648 3850 474660
rect 56502 474648 56508 474660
rect 56560 474648 56566 474700
rect 3602 471928 3608 471980
rect 3660 471968 3666 471980
rect 56502 471968 56508 471980
rect 3660 471940 56508 471968
rect 3660 471928 3666 471940
rect 56502 471928 56508 471940
rect 56560 471928 56566 471980
rect 31018 470500 31024 470552
rect 31076 470540 31082 470552
rect 56502 470540 56508 470552
rect 31076 470512 56508 470540
rect 31076 470500 31082 470512
rect 56502 470500 56508 470512
rect 56560 470500 56566 470552
rect 14458 467780 14464 467832
rect 14516 467820 14522 467832
rect 56502 467820 56508 467832
rect 14516 467792 56508 467820
rect 14516 467780 14522 467792
rect 56502 467780 56508 467792
rect 56560 467780 56566 467832
rect 282546 466420 282552 466472
rect 282604 466420 282610 466472
rect 3510 466352 3516 466404
rect 3568 466392 3574 466404
rect 56502 466392 56508 466404
rect 3568 466364 56508 466392
rect 3568 466352 3574 466364
rect 56502 466352 56508 466364
rect 56560 466352 56566 466404
rect 282564 466392 282592 466420
rect 282638 466392 282644 466404
rect 282564 466364 282644 466392
rect 282638 466352 282644 466364
rect 282696 466352 282702 466404
rect 21358 464992 21364 465044
rect 21416 465032 21422 465044
rect 56502 465032 56508 465044
rect 21416 465004 56508 465032
rect 21416 464992 21422 465004
rect 56502 464992 56508 465004
rect 56560 464992 56566 465044
rect 282362 463632 282368 463684
rect 282420 463672 282426 463684
rect 282638 463672 282644 463684
rect 282420 463644 282644 463672
rect 282420 463632 282426 463644
rect 282638 463632 282644 463644
rect 282696 463632 282702 463684
rect 13078 462272 13084 462324
rect 13136 462312 13142 462324
rect 56502 462312 56508 462324
rect 13136 462284 56508 462312
rect 13136 462272 13142 462284
rect 56502 462272 56508 462284
rect 56560 462272 56566 462324
rect 3418 460844 3424 460896
rect 3476 460884 3482 460896
rect 3476 460856 56732 460884
rect 3476 460844 3482 460856
rect 56594 460708 56600 460760
rect 56652 460748 56658 460760
rect 56704 460748 56732 460856
rect 56652 460720 56732 460748
rect 56652 460708 56658 460720
rect 24762 458124 24768 458176
rect 24820 458164 24826 458176
rect 56594 458164 56600 458176
rect 24820 458136 56600 458164
rect 24820 458124 24826 458136
rect 56594 458124 56600 458136
rect 56652 458124 56658 458176
rect 10318 456696 10324 456748
rect 10376 456736 10382 456748
rect 56594 456736 56600 456748
rect 10376 456708 56600 456736
rect 10376 456696 10382 456708
rect 56594 456696 56600 456708
rect 56652 456696 56658 456748
rect 42058 455336 42064 455388
rect 42116 455376 42122 455388
rect 56594 455376 56600 455388
rect 42116 455348 56600 455376
rect 42116 455336 42122 455348
rect 56594 455336 56600 455348
rect 56652 455336 56658 455388
rect 3418 452548 3424 452600
rect 3476 452588 3482 452600
rect 56594 452588 56600 452600
rect 3476 452560 56600 452588
rect 3476 452548 3482 452560
rect 56594 452548 56600 452560
rect 56652 452548 56658 452600
rect 282546 447108 282552 447160
rect 282604 447108 282610 447160
rect 282564 447080 282592 447108
rect 282638 447080 282644 447092
rect 282564 447052 282644 447080
rect 282638 447040 282644 447052
rect 282696 447040 282702 447092
rect 282822 434664 282828 434716
rect 282880 434704 282886 434716
rect 283006 434704 283012 434716
rect 282880 434676 283012 434704
rect 282880 434664 282886 434676
rect 283006 434664 283012 434676
rect 283064 434664 283070 434716
rect 281534 429156 281540 429208
rect 281592 429196 281598 429208
rect 367094 429196 367100 429208
rect 281592 429168 367100 429196
rect 281592 429156 281598 429168
rect 367094 429156 367100 429168
rect 367152 429156 367158 429208
rect 281534 427796 281540 427848
rect 281592 427836 281598 427848
rect 368474 427836 368480 427848
rect 281592 427808 368480 427836
rect 281592 427796 281598 427808
rect 368474 427796 368480 427808
rect 368532 427796 368538 427848
rect 281626 426504 281632 426556
rect 281684 426544 281690 426556
rect 369854 426544 369860 426556
rect 281684 426516 369860 426544
rect 281684 426504 281690 426516
rect 369854 426504 369860 426516
rect 369912 426504 369918 426556
rect 281534 426436 281540 426488
rect 281592 426476 281598 426488
rect 371234 426476 371240 426488
rect 281592 426448 371240 426476
rect 281592 426436 281598 426448
rect 371234 426436 371240 426448
rect 371292 426436 371298 426488
rect 281534 425076 281540 425128
rect 281592 425116 281598 425128
rect 372614 425116 372620 425128
rect 281592 425088 372620 425116
rect 281592 425076 281598 425088
rect 372614 425076 372620 425088
rect 372672 425076 372678 425128
rect 281534 423648 281540 423700
rect 281592 423688 281598 423700
rect 373994 423688 374000 423700
rect 281592 423660 374000 423688
rect 281592 423648 281598 423660
rect 373994 423648 374000 423660
rect 374052 423648 374058 423700
rect 281626 422356 281632 422408
rect 281684 422396 281690 422408
rect 374086 422396 374092 422408
rect 281684 422368 374092 422396
rect 281684 422356 281690 422368
rect 374086 422356 374092 422368
rect 374144 422356 374150 422408
rect 281534 422288 281540 422340
rect 281592 422328 281598 422340
rect 375374 422328 375380 422340
rect 281592 422300 375380 422328
rect 281592 422288 281598 422300
rect 375374 422288 375380 422300
rect 375432 422288 375438 422340
rect 281534 420928 281540 420980
rect 281592 420968 281598 420980
rect 376754 420968 376760 420980
rect 281592 420940 376760 420968
rect 281592 420928 281598 420940
rect 376754 420928 376760 420940
rect 376812 420928 376818 420980
rect 281534 419500 281540 419552
rect 281592 419540 281598 419552
rect 378134 419540 378140 419552
rect 281592 419512 378140 419540
rect 281592 419500 281598 419512
rect 378134 419500 378140 419512
rect 378192 419500 378198 419552
rect 59446 419432 59452 419484
rect 59504 419472 59510 419484
rect 59906 419472 59912 419484
rect 59504 419444 59912 419472
rect 59504 419432 59510 419444
rect 59906 419432 59912 419444
rect 59964 419432 59970 419484
rect 281626 418208 281632 418260
rect 281684 418248 281690 418260
rect 379514 418248 379520 418260
rect 281684 418220 379520 418248
rect 281684 418208 281690 418220
rect 379514 418208 379520 418220
rect 379572 418208 379578 418260
rect 281534 418140 281540 418192
rect 281592 418180 281598 418192
rect 380894 418180 380900 418192
rect 281592 418152 380900 418180
rect 281592 418140 281598 418152
rect 380894 418140 380900 418152
rect 380952 418140 380958 418192
rect 282822 416780 282828 416832
rect 282880 416820 282886 416832
rect 382274 416820 382280 416832
rect 282880 416792 382280 416820
rect 282880 416780 282886 416792
rect 382274 416780 382280 416792
rect 382332 416780 382338 416832
rect 282270 415420 282276 415472
rect 282328 415460 282334 415472
rect 382366 415460 382372 415472
rect 282328 415432 382372 415460
rect 282328 415420 282334 415432
rect 382366 415420 382372 415432
rect 382424 415420 382430 415472
rect 281718 414060 281724 414112
rect 281776 414100 281782 414112
rect 383838 414100 383844 414112
rect 281776 414072 383844 414100
rect 281776 414060 281782 414072
rect 383838 414060 383844 414072
rect 383896 414060 383902 414112
rect 282086 413992 282092 414044
rect 282144 414032 282150 414044
rect 385034 414032 385040 414044
rect 282144 414004 385040 414032
rect 282144 413992 282150 414004
rect 385034 413992 385040 414004
rect 385092 413992 385098 414044
rect 282638 413924 282644 413976
rect 282696 413964 282702 413976
rect 412634 413964 412640 413976
rect 282696 413936 412640 413964
rect 282696 413924 282702 413936
rect 412634 413924 412640 413936
rect 412692 413924 412698 413976
rect 383562 413856 383568 413908
rect 383620 413896 383626 413908
rect 393130 413896 393136 413908
rect 383620 413868 393136 413896
rect 383620 413856 383626 413868
rect 393130 413856 393136 413868
rect 393188 413856 393194 413908
rect 325878 413788 325884 413840
rect 325936 413828 325942 413840
rect 335170 413828 335176 413840
rect 325936 413800 335176 413828
rect 325936 413788 325942 413800
rect 335170 413788 335176 413800
rect 335228 413788 335234 413840
rect 345198 413788 345204 413840
rect 345256 413828 345262 413840
rect 354490 413828 354496 413840
rect 345256 413800 354496 413828
rect 345256 413788 345262 413800
rect 354490 413788 354496 413800
rect 354548 413788 354554 413840
rect 378042 413788 378048 413840
rect 378100 413828 378106 413840
rect 387334 413828 387340 413840
rect 378100 413800 387340 413828
rect 378100 413788 378106 413800
rect 387334 413788 387340 413800
rect 387392 413828 387398 413840
rect 396074 413828 396080 413840
rect 387392 413800 396080 413828
rect 387392 413788 387398 413800
rect 396074 413788 396080 413800
rect 396132 413788 396138 413840
rect 325786 413720 325792 413772
rect 325844 413760 325850 413772
rect 335262 413760 335268 413772
rect 325844 413732 335268 413760
rect 325844 413720 325850 413732
rect 335262 413720 335268 413732
rect 335320 413720 335326 413772
rect 345106 413720 345112 413772
rect 345164 413760 345170 413772
rect 354582 413760 354588 413772
rect 345164 413732 354588 413760
rect 345164 413720 345170 413732
rect 354582 413720 354588 413732
rect 354640 413720 354646 413772
rect 369762 413720 369768 413772
rect 369820 413760 369826 413772
rect 378778 413760 378784 413772
rect 369820 413732 378784 413760
rect 369820 413720 369826 413732
rect 378778 413720 378784 413732
rect 378836 413760 378842 413772
rect 388346 413760 388352 413772
rect 378836 413732 388352 413760
rect 378836 413720 378842 413732
rect 388346 413720 388352 413732
rect 388404 413760 388410 413772
rect 397454 413760 397460 413772
rect 388404 413732 397460 413760
rect 388404 413720 388410 413732
rect 397454 413720 397460 413732
rect 397512 413720 397518 413772
rect 282638 413652 282644 413704
rect 282696 413692 282702 413704
rect 368290 413692 368296 413704
rect 282696 413664 368296 413692
rect 282696 413652 282702 413664
rect 368290 413652 368296 413664
rect 368348 413692 368354 413704
rect 378042 413692 378048 413704
rect 368348 413664 378048 413692
rect 368348 413652 368354 413664
rect 378042 413652 378048 413664
rect 378100 413652 378106 413704
rect 386046 413652 386052 413704
rect 386104 413692 386110 413704
rect 394694 413692 394700 413704
rect 386104 413664 394700 413692
rect 386104 413652 386110 413664
rect 394694 413652 394700 413664
rect 394752 413652 394758 413704
rect 281534 413584 281540 413636
rect 281592 413624 281598 413636
rect 368750 413624 368756 413636
rect 281592 413596 368756 413624
rect 281592 413584 281598 413596
rect 368750 413584 368756 413596
rect 368808 413584 368814 413636
rect 368842 413584 368848 413636
rect 368900 413624 368906 413636
rect 369854 413624 369860 413636
rect 368900 413596 369860 413624
rect 368900 413584 368906 413596
rect 369854 413584 369860 413596
rect 369912 413624 369918 413636
rect 379606 413624 379612 413636
rect 369912 413596 379612 413624
rect 369912 413584 369918 413596
rect 379606 413584 379612 413596
rect 379664 413624 379670 413636
rect 389634 413624 389640 413636
rect 379664 413596 389640 413624
rect 379664 413584 379670 413596
rect 389634 413584 389640 413596
rect 389692 413584 389698 413636
rect 318242 413516 318248 413568
rect 318300 413556 318306 413568
rect 405734 413556 405740 413568
rect 318300 413528 405740 413556
rect 318300 413516 318306 413528
rect 405734 413516 405740 413528
rect 405792 413516 405798 413568
rect 281810 413448 281816 413500
rect 281868 413488 281874 413500
rect 368842 413488 368848 413500
rect 281868 413460 368848 413488
rect 281868 413448 281874 413460
rect 368842 413448 368848 413460
rect 368900 413448 368906 413500
rect 368934 413448 368940 413500
rect 368992 413488 368998 413500
rect 372982 413488 372988 413500
rect 368992 413460 372988 413488
rect 368992 413448 368998 413460
rect 372982 413448 372988 413460
rect 373040 413488 373046 413500
rect 382274 413488 382280 413500
rect 373040 413460 382280 413488
rect 373040 413448 373046 413460
rect 382274 413448 382280 413460
rect 382332 413448 382338 413500
rect 384942 413448 384948 413500
rect 385000 413488 385006 413500
rect 393958 413488 393964 413500
rect 385000 413460 393964 413488
rect 385000 413448 385006 413460
rect 393958 413448 393964 413460
rect 394016 413448 394022 413500
rect 394694 413448 394700 413500
rect 394752 413488 394758 413500
rect 395338 413488 395344 413500
rect 394752 413460 395344 413488
rect 394752 413448 394758 413460
rect 395338 413448 395344 413460
rect 395396 413488 395402 413500
rect 404354 413488 404360 413500
rect 395396 413460 404360 413488
rect 395396 413448 395402 413460
rect 404354 413448 404360 413460
rect 404412 413448 404418 413500
rect 287146 413380 287152 413432
rect 287204 413420 287210 413432
rect 296530 413420 296536 413432
rect 287204 413392 296536 413420
rect 287204 413380 287210 413392
rect 296530 413380 296536 413392
rect 296588 413380 296594 413432
rect 306466 413380 306472 413432
rect 306524 413420 306530 413432
rect 315850 413420 315856 413432
rect 306524 413392 315856 413420
rect 306524 413380 306530 413392
rect 315850 413380 315856 413392
rect 315908 413380 315914 413432
rect 318150 413380 318156 413432
rect 318208 413420 318214 413432
rect 407114 413420 407120 413432
rect 318208 413392 407120 413420
rect 318208 413380 318214 413392
rect 407114 413380 407120 413392
rect 407172 413380 407178 413432
rect 282178 413312 282184 413364
rect 282236 413352 282242 413364
rect 371970 413352 371976 413364
rect 282236 413324 371976 413352
rect 282236 413312 282242 413324
rect 371970 413312 371976 413324
rect 372028 413352 372034 413364
rect 381538 413352 381544 413364
rect 372028 413324 381544 413352
rect 372028 413312 372034 413324
rect 381538 413312 381544 413324
rect 381596 413352 381602 413364
rect 390922 413352 390928 413364
rect 381596 413324 390928 413352
rect 381596 413312 381602 413324
rect 390922 413312 390928 413324
rect 390980 413352 390986 413364
rect 391842 413352 391848 413364
rect 390980 413324 391848 413352
rect 390980 413312 390986 413324
rect 391842 413312 391848 413324
rect 391900 413312 391906 413364
rect 393130 413312 393136 413364
rect 393188 413352 393194 413364
rect 401594 413352 401600 413364
rect 393188 413324 401600 413352
rect 393188 413312 393194 413324
rect 401594 413312 401600 413324
rect 401652 413312 401658 413364
rect 282822 413244 282828 413296
rect 282880 413284 282886 413296
rect 386414 413284 386420 413296
rect 282880 413256 386420 413284
rect 282880 413244 282886 413256
rect 386414 413244 386420 413256
rect 386472 413244 386478 413296
rect 393958 413244 393964 413296
rect 394016 413284 394022 413296
rect 403158 413284 403164 413296
rect 394016 413256 403164 413284
rect 394016 413244 394022 413256
rect 403158 413244 403164 413256
rect 403216 413244 403222 413296
rect 287054 413176 287060 413228
rect 287112 413216 287118 413228
rect 296622 413216 296628 413228
rect 287112 413188 296628 413216
rect 287112 413176 287118 413188
rect 296622 413176 296628 413188
rect 296680 413176 296686 413228
rect 306374 413176 306380 413228
rect 306432 413216 306438 413228
rect 315942 413216 315948 413228
rect 306432 413188 315948 413216
rect 306432 413176 306438 413188
rect 315942 413176 315948 413188
rect 316000 413176 316006 413228
rect 318058 413176 318064 413228
rect 318116 413216 318122 413228
rect 408494 413216 408500 413228
rect 318116 413188 408500 413216
rect 318116 413176 318122 413188
rect 408494 413176 408500 413188
rect 408552 413176 408558 413228
rect 282362 413108 282368 413160
rect 282420 413148 282426 413160
rect 368934 413148 368940 413160
rect 282420 413120 368940 413148
rect 282420 413108 282426 413120
rect 368934 413108 368940 413120
rect 368992 413108 368998 413160
rect 369044 413120 369348 413148
rect 281994 413040 282000 413092
rect 282052 413080 282058 413092
rect 287146 413080 287152 413092
rect 282052 413052 287152 413080
rect 282052 413040 282058 413052
rect 287146 413040 287152 413052
rect 287204 413040 287210 413092
rect 296530 413040 296536 413092
rect 296588 413080 296594 413092
rect 306466 413080 306472 413092
rect 296588 413052 306472 413080
rect 296588 413040 296594 413052
rect 306466 413040 306472 413052
rect 306524 413040 306530 413092
rect 315850 413040 315856 413092
rect 315908 413080 315914 413092
rect 325878 413080 325884 413092
rect 315908 413052 325884 413080
rect 315908 413040 315914 413052
rect 325878 413040 325884 413052
rect 325936 413040 325942 413092
rect 335170 413040 335176 413092
rect 335228 413080 335234 413092
rect 345198 413080 345204 413092
rect 335228 413052 345204 413080
rect 335228 413040 335234 413052
rect 345198 413040 345204 413052
rect 345256 413040 345262 413092
rect 354490 413040 354496 413092
rect 354548 413080 354554 413092
rect 368842 413080 368848 413092
rect 354548 413052 368848 413080
rect 354548 413040 354554 413052
rect 368842 413040 368848 413052
rect 368900 413040 368906 413092
rect 282454 412972 282460 413024
rect 282512 413012 282518 413024
rect 287054 413012 287060 413024
rect 282512 412984 287060 413012
rect 282512 412972 282518 412984
rect 287054 412972 287060 412984
rect 287112 412972 287118 413024
rect 296622 412972 296628 413024
rect 296680 413012 296686 413024
rect 306374 413012 306380 413024
rect 296680 412984 306380 413012
rect 296680 412972 296686 412984
rect 306374 412972 306380 412984
rect 306432 412972 306438 413024
rect 315942 412972 315948 413024
rect 316000 413012 316006 413024
rect 325786 413012 325792 413024
rect 316000 412984 325792 413012
rect 316000 412972 316006 412984
rect 325786 412972 325792 412984
rect 325844 412972 325850 413024
rect 335262 412972 335268 413024
rect 335320 413012 335326 413024
rect 345106 413012 345112 413024
rect 335320 412984 345112 413012
rect 335320 412972 335326 412984
rect 345106 412972 345112 412984
rect 345164 412972 345170 413024
rect 354582 412972 354588 413024
rect 354640 413012 354646 413024
rect 369044 413012 369072 413120
rect 369320 413080 369348 413120
rect 382274 413108 382280 413160
rect 382332 413148 382338 413160
rect 391750 413148 391756 413160
rect 382332 413120 391756 413148
rect 382332 413108 382338 413120
rect 391750 413108 391756 413120
rect 391808 413108 391814 413160
rect 391842 413108 391848 413160
rect 391900 413148 391906 413160
rect 398834 413148 398840 413160
rect 391900 413120 398840 413148
rect 391900 413108 391906 413120
rect 398834 413108 398840 413120
rect 398892 413108 398898 413160
rect 375466 413080 375472 413092
rect 369320 413052 375472 413080
rect 375466 413040 375472 413052
rect 375524 413080 375530 413092
rect 391768 413080 391796 413108
rect 400214 413080 400220 413092
rect 375524 413052 383608 413080
rect 391768 413052 400220 413080
rect 375524 413040 375530 413052
rect 354640 412984 369072 413012
rect 354640 412972 354646 412984
rect 369302 412972 369308 413024
rect 369360 413012 369366 413024
rect 374362 413012 374368 413024
rect 369360 412984 374368 413012
rect 369360 412972 369366 412984
rect 374362 412972 374368 412984
rect 374420 413012 374426 413024
rect 383470 413012 383476 413024
rect 374420 412984 383476 413012
rect 374420 412972 374426 412984
rect 383470 412972 383476 412984
rect 383528 412972 383534 413024
rect 383580 413012 383608 413052
rect 400214 413040 400220 413052
rect 400272 413040 400278 413092
rect 384942 413012 384948 413024
rect 383580 412984 384948 413012
rect 384942 412972 384948 412984
rect 385000 412972 385006 413024
rect 282270 412904 282276 412956
rect 282328 412944 282334 412956
rect 376570 412944 376576 412956
rect 282328 412916 376576 412944
rect 282328 412904 282334 412916
rect 376570 412904 376576 412916
rect 376628 412944 376634 412956
rect 386046 412944 386052 412956
rect 376628 412916 386052 412944
rect 376628 412904 376634 412916
rect 386046 412904 386052 412916
rect 386104 412904 386110 412956
rect 389634 412904 389640 412956
rect 389692 412944 389698 412956
rect 397454 412944 397460 412956
rect 389692 412916 397460 412944
rect 389692 412904 389698 412916
rect 397454 412904 397460 412916
rect 397512 412904 397518 412956
rect 282730 412836 282736 412888
rect 282788 412876 282794 412888
rect 393314 412876 393320 412888
rect 282788 412848 393320 412876
rect 282788 412836 282794 412848
rect 393314 412836 393320 412848
rect 393372 412836 393378 412888
rect 282086 412768 282092 412820
rect 282144 412808 282150 412820
rect 394694 412808 394700 412820
rect 282144 412780 394700 412808
rect 282144 412768 282150 412780
rect 394694 412768 394700 412780
rect 394752 412768 394758 412820
rect 281534 412700 281540 412752
rect 281592 412700 281598 412752
rect 281626 412700 281632 412752
rect 281684 412740 281690 412752
rect 396074 412740 396080 412752
rect 281684 412712 396080 412740
rect 281684 412700 281690 412712
rect 396074 412700 396080 412712
rect 396132 412700 396138 412752
rect 281552 412672 281580 412700
rect 405734 412672 405740 412684
rect 281552 412644 405740 412672
rect 405734 412632 405740 412644
rect 405792 412632 405798 412684
rect 281534 412564 281540 412616
rect 281592 412564 281598 412616
rect 281552 412344 281580 412564
rect 281810 412496 281816 412548
rect 281868 412496 281874 412548
rect 281828 412468 281856 412496
rect 282730 412468 282736 412480
rect 281828 412440 282736 412468
rect 282730 412428 282736 412440
rect 282788 412428 282794 412480
rect 281810 412360 281816 412412
rect 281868 412400 281874 412412
rect 282086 412400 282092 412412
rect 281868 412372 282092 412400
rect 281868 412360 281874 412372
rect 282086 412360 282092 412372
rect 282144 412360 282150 412412
rect 284110 412360 284116 412412
rect 284168 412400 284174 412412
rect 343726 412400 343732 412412
rect 284168 412372 343732 412400
rect 284168 412360 284174 412372
rect 343726 412360 343732 412372
rect 343784 412360 343790 412412
rect 281534 412292 281540 412344
rect 281592 412292 281598 412344
rect 284018 412292 284024 412344
rect 284076 412332 284082 412344
rect 343634 412332 343640 412344
rect 284076 412304 343640 412332
rect 284076 412292 284082 412304
rect 343634 412292 343640 412304
rect 343692 412292 343698 412344
rect 284202 412224 284208 412276
rect 284260 412264 284266 412276
rect 345014 412264 345020 412276
rect 284260 412236 345020 412264
rect 284260 412224 284266 412236
rect 345014 412224 345020 412236
rect 345072 412224 345078 412276
rect 283466 412156 283472 412208
rect 283524 412196 283530 412208
rect 346394 412196 346400 412208
rect 283524 412168 346400 412196
rect 283524 412156 283530 412168
rect 346394 412156 346400 412168
rect 346452 412156 346458 412208
rect 283374 412088 283380 412140
rect 283432 412128 283438 412140
rect 347774 412128 347780 412140
rect 283432 412100 347780 412128
rect 283432 412088 283438 412100
rect 347774 412088 347780 412100
rect 347832 412088 347838 412140
rect 282914 412020 282920 412072
rect 282972 412060 282978 412072
rect 349154 412060 349160 412072
rect 282972 412032 349160 412060
rect 282972 412020 282978 412032
rect 349154 412020 349160 412032
rect 349212 412020 349218 412072
rect 281902 411952 281908 412004
rect 281960 411992 281966 412004
rect 350626 411992 350632 412004
rect 281960 411964 350632 411992
rect 281960 411952 281966 411964
rect 350626 411952 350632 411964
rect 350684 411952 350690 412004
rect 305638 411884 305644 411936
rect 305696 411924 305702 411936
rect 419534 411924 419540 411936
rect 305696 411896 419540 411924
rect 305696 411884 305702 411896
rect 419534 411884 419540 411896
rect 419592 411884 419598 411936
rect 311158 411816 311164 411868
rect 311216 411856 311222 411868
rect 397454 411856 397460 411868
rect 311216 411828 397460 411856
rect 311216 411816 311222 411828
rect 397454 411816 397460 411828
rect 397512 411816 397518 411868
rect 282086 411748 282092 411800
rect 282144 411788 282150 411800
rect 388070 411788 388076 411800
rect 282144 411760 388076 411788
rect 282144 411748 282150 411760
rect 388070 411748 388076 411760
rect 388128 411748 388134 411800
rect 283006 411680 283012 411732
rect 283064 411720 283070 411732
rect 391014 411720 391020 411732
rect 283064 411692 391020 411720
rect 283064 411680 283070 411692
rect 391014 411680 391020 411692
rect 391072 411680 391078 411732
rect 285030 411612 285036 411664
rect 285088 411652 285094 411664
rect 399110 411652 399116 411664
rect 285088 411624 399116 411652
rect 285088 411612 285094 411624
rect 399110 411612 399116 411624
rect 399168 411612 399174 411664
rect 282086 411544 282092 411596
rect 282144 411584 282150 411596
rect 398006 411584 398012 411596
rect 282144 411556 398012 411584
rect 282144 411544 282150 411556
rect 398006 411544 398012 411556
rect 398064 411544 398070 411596
rect 283098 411476 283104 411528
rect 283156 411516 283162 411528
rect 400950 411516 400956 411528
rect 283156 411488 400956 411516
rect 283156 411476 283162 411488
rect 400950 411476 400956 411488
rect 401008 411476 401014 411528
rect 283282 411408 283288 411460
rect 283340 411448 283346 411460
rect 401686 411448 401692 411460
rect 283340 411420 401692 411448
rect 283340 411408 283346 411420
rect 401686 411408 401692 411420
rect 401744 411408 401750 411460
rect 282454 411340 282460 411392
rect 282512 411380 282518 411392
rect 282822 411380 282828 411392
rect 282512 411352 282828 411380
rect 282512 411340 282518 411352
rect 282822 411340 282828 411352
rect 282880 411340 282886 411392
rect 284938 411340 284944 411392
rect 284996 411380 285002 411392
rect 404354 411380 404360 411392
rect 284996 411352 404360 411380
rect 284996 411340 285002 411352
rect 404354 411340 404360 411352
rect 404412 411340 404418 411392
rect 281902 411312 281908 411324
rect 281828 411284 281908 411312
rect 281828 410156 281856 411284
rect 281902 411272 281908 411284
rect 281960 411272 281966 411324
rect 283190 411272 283196 411324
rect 283248 411312 283254 411324
rect 403250 411312 403256 411324
rect 283248 411284 403256 411312
rect 283248 411272 283254 411284
rect 403250 411272 403256 411284
rect 403308 411272 403314 411324
rect 282822 411204 282828 411256
rect 282880 411244 282886 411256
rect 389266 411244 389272 411256
rect 282880 411216 389272 411244
rect 282880 411204 282886 411216
rect 389266 411204 389272 411216
rect 389324 411204 389330 411256
rect 281902 411136 281908 411188
rect 281960 411176 281966 411188
rect 389726 411176 389732 411188
rect 281960 411148 389732 411176
rect 281960 411136 281966 411148
rect 389726 411136 389732 411148
rect 389784 411136 389790 411188
rect 298738 410728 298744 410780
rect 298796 410768 298802 410780
rect 342254 410768 342260 410780
rect 298796 410740 342260 410768
rect 298796 410728 298802 410740
rect 342254 410728 342260 410740
rect 342312 410728 342318 410780
rect 283926 410660 283932 410712
rect 283984 410700 283990 410712
rect 340874 410700 340880 410712
rect 283984 410672 340880 410700
rect 283984 410660 283990 410672
rect 340874 410660 340880 410672
rect 340932 410660 340938 410712
rect 282914 410592 282920 410644
rect 282972 410632 282978 410644
rect 392302 410632 392308 410644
rect 282972 410604 392308 410632
rect 282972 410592 282978 410604
rect 392302 410592 392308 410604
rect 392360 410592 392366 410644
rect 283834 410524 283840 410576
rect 283892 410564 283898 410576
rect 409966 410564 409972 410576
rect 283892 410536 409972 410564
rect 283892 410524 283898 410536
rect 409966 410524 409972 410536
rect 410024 410524 410030 410576
rect 281902 410156 281908 410168
rect 281828 410128 281908 410156
rect 281902 410116 281908 410128
rect 281960 410116 281966 410168
rect 282086 407872 282092 407924
rect 282144 407872 282150 407924
rect 282178 407872 282184 407924
rect 282236 407912 282242 407924
rect 282638 407912 282644 407924
rect 282236 407884 282644 407912
rect 282236 407872 282242 407884
rect 282638 407872 282644 407884
rect 282696 407872 282702 407924
rect 281626 407804 281632 407856
rect 281684 407844 281690 407856
rect 281684 407816 282040 407844
rect 281684 407804 281690 407816
rect 282012 407720 282040 407816
rect 281626 407668 281632 407720
rect 281684 407708 281690 407720
rect 281902 407708 281908 407720
rect 281684 407680 281908 407708
rect 281684 407668 281690 407680
rect 281902 407668 281908 407680
rect 281960 407668 281966 407720
rect 281994 407668 282000 407720
rect 282052 407668 282058 407720
rect 282104 407640 282132 407872
rect 281920 407612 282132 407640
rect 281920 407584 281948 407612
rect 281902 407532 281908 407584
rect 281960 407532 281966 407584
rect 281994 407532 282000 407584
rect 282052 407572 282058 407584
rect 282730 407572 282736 407584
rect 282052 407544 282736 407572
rect 282052 407532 282058 407544
rect 282730 407532 282736 407544
rect 282788 407532 282794 407584
rect 282822 404268 282828 404320
rect 282880 404308 282886 404320
rect 311158 404308 311164 404320
rect 282880 404280 311164 404308
rect 282880 404268 282886 404280
rect 311158 404268 311164 404280
rect 311216 404268 311222 404320
rect 282270 402840 282276 402892
rect 282328 402840 282334 402892
rect 282288 402688 282316 402840
rect 282270 402636 282276 402688
rect 282328 402636 282334 402688
rect 282178 402568 282184 402620
rect 282236 402608 282242 402620
rect 285030 402608 285036 402620
rect 282236 402580 285036 402608
rect 282236 402568 282242 402580
rect 285030 402568 285036 402580
rect 285088 402568 285094 402620
rect 281626 401140 281632 401192
rect 281684 401180 281690 401192
rect 283098 401180 283104 401192
rect 281684 401152 283104 401180
rect 281684 401140 281690 401152
rect 283098 401140 283104 401152
rect 283156 401140 283162 401192
rect 281626 400120 281632 400172
rect 281684 400160 281690 400172
rect 283282 400160 283288 400172
rect 281684 400132 283288 400160
rect 281684 400120 281690 400132
rect 283282 400120 283288 400132
rect 283340 400120 283346 400172
rect 281626 399508 281632 399560
rect 281684 399548 281690 399560
rect 283190 399548 283196 399560
rect 281684 399520 283196 399548
rect 281684 399508 281690 399520
rect 283190 399508 283196 399520
rect 283248 399508 283254 399560
rect 282178 398148 282184 398200
rect 282236 398188 282242 398200
rect 284938 398188 284944 398200
rect 282236 398160 284944 398188
rect 282236 398148 282242 398160
rect 284938 398148 284944 398160
rect 284996 398148 285002 398200
rect 3142 395972 3148 396024
rect 3200 396012 3206 396024
rect 56686 396012 56692 396024
rect 3200 395984 56692 396012
rect 3200 395972 3206 395984
rect 56686 395972 56692 395984
rect 56744 395972 56750 396024
rect 281626 394544 281632 394596
rect 281684 394584 281690 394596
rect 283742 394584 283748 394596
rect 281684 394556 283748 394584
rect 281684 394544 281690 394556
rect 283742 394544 283748 394556
rect 283800 394544 283806 394596
rect 282178 393252 282184 393304
rect 282236 393292 282242 393304
rect 282546 393292 282552 393304
rect 282236 393264 282552 393292
rect 282236 393252 282242 393264
rect 282546 393252 282552 393264
rect 282604 393252 282610 393304
rect 281810 393184 281816 393236
rect 281868 393224 281874 393236
rect 282362 393224 282368 393236
rect 281868 393196 282368 393224
rect 281868 393184 281874 393196
rect 282362 393184 282368 393196
rect 282420 393184 282426 393236
rect 281626 393116 281632 393168
rect 281684 393156 281690 393168
rect 283558 393156 283564 393168
rect 281684 393128 283564 393156
rect 281684 393116 281690 393128
rect 283558 393116 283564 393128
rect 283616 393116 283622 393168
rect 281626 392368 281632 392420
rect 281684 392408 281690 392420
rect 283650 392408 283656 392420
rect 281684 392380 283656 392408
rect 281684 392368 281690 392380
rect 283650 392368 283656 392380
rect 283708 392368 283714 392420
rect 310422 389784 310428 389836
rect 310480 389824 310486 389836
rect 338022 389824 338028 389836
rect 310480 389796 338028 389824
rect 310480 389784 310486 389796
rect 338022 389784 338028 389796
rect 338080 389784 338086 389836
rect 281626 388152 281632 388204
rect 281684 388192 281690 388204
rect 283374 388192 283380 388204
rect 281684 388164 283380 388192
rect 281684 388152 281690 388164
rect 283374 388152 283380 388164
rect 283432 388152 283438 388204
rect 281626 386996 281632 387048
rect 281684 387036 281690 387048
rect 283466 387036 283472 387048
rect 281684 387008 283472 387036
rect 281684 386996 281690 387008
rect 283466 386996 283472 387008
rect 283524 386996 283530 387048
rect 281718 386044 281724 386096
rect 281776 386084 281782 386096
rect 284202 386084 284208 386096
rect 281776 386056 284208 386084
rect 281776 386044 281782 386056
rect 284202 386044 284208 386056
rect 284260 386044 284266 386096
rect 281626 385568 281632 385620
rect 281684 385608 281690 385620
rect 284110 385608 284116 385620
rect 281684 385580 284116 385608
rect 281684 385568 281690 385580
rect 284110 385568 284116 385580
rect 284168 385568 284174 385620
rect 281626 384888 281632 384940
rect 281684 384928 281690 384940
rect 284018 384928 284024 384940
rect 281684 384900 284024 384928
rect 281684 384888 281690 384900
rect 284018 384888 284024 384900
rect 284076 384888 284082 384940
rect 281718 383800 281724 383852
rect 281776 383840 281782 383852
rect 281776 383812 282500 383840
rect 281776 383800 281782 383812
rect 282472 383784 282500 383812
rect 281810 383732 281816 383784
rect 281868 383772 281874 383784
rect 282362 383772 282368 383784
rect 281868 383744 282368 383772
rect 281868 383732 281874 383744
rect 282362 383732 282368 383744
rect 282420 383732 282426 383784
rect 282454 383732 282460 383784
rect 282512 383732 282518 383784
rect 282178 383664 282184 383716
rect 282236 383704 282242 383716
rect 282546 383704 282552 383716
rect 282236 383676 282552 383704
rect 282236 383664 282242 383676
rect 282546 383664 282552 383676
rect 282604 383664 282610 383716
rect 282822 383596 282828 383648
rect 282880 383636 282886 383648
rect 298738 383636 298744 383648
rect 282880 383608 298744 383636
rect 282880 383596 282886 383608
rect 298738 383596 298744 383608
rect 298796 383596 298802 383648
rect 281718 382168 281724 382220
rect 281776 382208 281782 382220
rect 339494 382208 339500 382220
rect 281776 382180 339500 382208
rect 281776 382168 281782 382180
rect 339494 382168 339500 382180
rect 339552 382168 339558 382220
rect 281626 381964 281632 382016
rect 281684 382004 281690 382016
rect 283926 382004 283932 382016
rect 281684 381976 283932 382004
rect 281684 381964 281690 381976
rect 283926 381964 283932 381976
rect 283984 381964 283990 382016
rect 3234 380808 3240 380860
rect 3292 380848 3298 380860
rect 57054 380848 57060 380860
rect 3292 380820 57060 380848
rect 3292 380808 3298 380820
rect 57054 380808 57060 380820
rect 57112 380808 57118 380860
rect 282822 380808 282828 380860
rect 282880 380848 282886 380860
rect 338114 380848 338120 380860
rect 282880 380820 338120 380848
rect 282880 380808 282886 380820
rect 338114 380808 338120 380820
rect 338172 380808 338178 380860
rect 282822 379448 282828 379500
rect 282880 379488 282886 379500
rect 336826 379488 336832 379500
rect 282880 379460 336832 379488
rect 282880 379448 282886 379460
rect 336826 379448 336832 379460
rect 336884 379448 336890 379500
rect 282822 378088 282828 378140
rect 282880 378128 282886 378140
rect 336734 378128 336740 378140
rect 282880 378100 336740 378128
rect 282880 378088 282886 378100
rect 336734 378088 336740 378100
rect 336792 378088 336798 378140
rect 282178 378020 282184 378072
rect 282236 378060 282242 378072
rect 335354 378060 335360 378072
rect 282236 378032 335360 378060
rect 282236 378020 282242 378032
rect 335354 378020 335360 378032
rect 335412 378020 335418 378072
rect 282822 376660 282828 376712
rect 282880 376700 282886 376712
rect 333974 376700 333980 376712
rect 282880 376672 333980 376700
rect 282880 376660 282886 376672
rect 333974 376660 333980 376672
rect 334032 376660 334038 376712
rect 282822 375300 282828 375352
rect 282880 375340 282886 375352
rect 332594 375340 332600 375352
rect 282880 375312 332600 375340
rect 282880 375300 282886 375312
rect 332594 375300 332600 375312
rect 332652 375300 332658 375352
rect 281902 373940 281908 373992
rect 281960 373980 281966 373992
rect 282546 373980 282552 373992
rect 281960 373952 282552 373980
rect 281960 373940 281966 373952
rect 282546 373940 282552 373952
rect 282604 373940 282610 373992
rect 282822 373940 282828 373992
rect 282880 373980 282886 373992
rect 331214 373980 331220 373992
rect 282880 373952 331220 373980
rect 282880 373940 282886 373952
rect 331214 373940 331220 373952
rect 331272 373940 331278 373992
rect 282178 373872 282184 373924
rect 282236 373912 282242 373924
rect 329926 373912 329932 373924
rect 282236 373884 329932 373912
rect 282236 373872 282242 373884
rect 329926 373872 329932 373884
rect 329984 373872 329990 373924
rect 281810 373804 281816 373856
rect 281868 373844 281874 373856
rect 282362 373844 282368 373856
rect 281868 373816 282368 373844
rect 281868 373804 281874 373816
rect 282362 373804 282368 373816
rect 282420 373804 282426 373856
rect 282454 373804 282460 373856
rect 282512 373804 282518 373856
rect 281718 373736 281724 373788
rect 281776 373776 281782 373788
rect 282472 373776 282500 373804
rect 281776 373748 282500 373776
rect 281776 373736 281782 373748
rect 282822 372512 282828 372564
rect 282880 372552 282886 372564
rect 329834 372552 329840 372564
rect 282880 372524 329840 372552
rect 282880 372512 282886 372524
rect 329834 372512 329840 372524
rect 329892 372512 329898 372564
rect 282822 371152 282828 371204
rect 282880 371192 282886 371204
rect 328454 371192 328460 371204
rect 282880 371164 328460 371192
rect 282880 371152 282886 371164
rect 328454 371152 328460 371164
rect 328512 371152 328518 371204
rect 282178 371084 282184 371136
rect 282236 371124 282242 371136
rect 327074 371124 327080 371136
rect 282236 371096 327080 371124
rect 282236 371084 282242 371096
rect 327074 371084 327080 371096
rect 327132 371084 327138 371136
rect 282822 369792 282828 369844
rect 282880 369832 282886 369844
rect 325694 369832 325700 369844
rect 282880 369804 325700 369832
rect 282880 369792 282886 369804
rect 325694 369792 325700 369804
rect 325752 369792 325758 369844
rect 282822 368432 282828 368484
rect 282880 368472 282886 368484
rect 324314 368472 324320 368484
rect 282880 368444 324320 368472
rect 282880 368432 282886 368444
rect 324314 368432 324320 368444
rect 324372 368432 324378 368484
rect 3142 367004 3148 367056
rect 3200 367044 3206 367056
rect 15838 367044 15844 367056
rect 3200 367016 15844 367044
rect 3200 367004 3206 367016
rect 15838 367004 15844 367016
rect 15896 367004 15902 367056
rect 282822 367004 282828 367056
rect 282880 367044 282886 367056
rect 322934 367044 322940 367056
rect 282880 367016 322940 367044
rect 282880 367004 282886 367016
rect 322934 367004 322940 367016
rect 322992 367004 322998 367056
rect 282178 366936 282184 366988
rect 282236 366976 282242 366988
rect 321554 366976 321560 366988
rect 282236 366948 321560 366976
rect 282236 366936 282242 366948
rect 321554 366936 321560 366948
rect 321612 366936 321618 366988
rect 282822 365644 282828 365696
rect 282880 365684 282886 365696
rect 330478 365684 330484 365696
rect 282880 365656 330484 365684
rect 282880 365644 282886 365656
rect 330478 365644 330484 365656
rect 330536 365644 330542 365696
rect 281718 364488 281724 364540
rect 281776 364528 281782 364540
rect 281776 364500 282500 364528
rect 281776 364488 281782 364500
rect 282472 364472 282500 364500
rect 281810 364420 281816 364472
rect 281868 364460 281874 364472
rect 282362 364460 282368 364472
rect 281868 364432 282368 364460
rect 281868 364420 281874 364432
rect 282362 364420 282368 364432
rect 282420 364420 282426 364472
rect 282454 364420 282460 364472
rect 282512 364420 282518 364472
rect 281902 364352 281908 364404
rect 281960 364392 281966 364404
rect 282546 364392 282552 364404
rect 281960 364364 282552 364392
rect 281960 364352 281966 364364
rect 282546 364352 282552 364364
rect 282604 364352 282610 364404
rect 282822 364284 282828 364336
rect 282880 364324 282886 364336
rect 329282 364324 329288 364336
rect 282880 364296 329288 364324
rect 282880 364284 282886 364296
rect 329282 364284 329288 364296
rect 329340 364284 329346 364336
rect 282178 362924 282184 362976
rect 282236 362964 282242 362976
rect 282730 362964 282736 362976
rect 282236 362936 282736 362964
rect 282236 362924 282242 362936
rect 282730 362924 282736 362936
rect 282788 362924 282794 362976
rect 282822 362856 282828 362908
rect 282880 362896 282886 362908
rect 329098 362896 329104 362908
rect 282880 362868 329104 362896
rect 282880 362856 282886 362868
rect 329098 362856 329104 362868
rect 329156 362856 329162 362908
rect 282730 362788 282736 362840
rect 282788 362828 282794 362840
rect 327718 362828 327724 362840
rect 282788 362800 327724 362828
rect 282788 362788 282794 362800
rect 327718 362788 327724 362800
rect 327776 362788 327782 362840
rect 281718 361496 281724 361548
rect 281776 361536 281782 361548
rect 326338 361536 326344 361548
rect 281776 361508 326344 361536
rect 281776 361496 281782 361508
rect 326338 361496 326344 361508
rect 326396 361496 326402 361548
rect 282822 360136 282828 360188
rect 282880 360176 282886 360188
rect 324958 360176 324964 360188
rect 282880 360148 324964 360176
rect 282880 360136 282886 360148
rect 324958 360136 324964 360148
rect 325016 360136 325022 360188
rect 282730 360068 282736 360120
rect 282788 360108 282794 360120
rect 323578 360108 323584 360120
rect 282788 360080 323584 360108
rect 282788 360068 282794 360080
rect 323578 360068 323584 360080
rect 323636 360068 323642 360120
rect 281902 358708 281908 358760
rect 281960 358748 281966 358760
rect 322198 358748 322204 358760
rect 281960 358720 322204 358748
rect 281960 358708 281966 358720
rect 322198 358708 322204 358720
rect 322256 358708 322262 358760
rect 282086 354560 282092 354612
rect 282144 354600 282150 354612
rect 282454 354600 282460 354612
rect 282144 354572 282460 354600
rect 282144 354560 282150 354572
rect 282454 354560 282460 354572
rect 282512 354560 282518 354612
rect 282822 349052 282828 349104
rect 282880 349092 282886 349104
rect 297358 349092 297364 349104
rect 282880 349064 297364 349092
rect 282880 349052 282886 349064
rect 297358 349052 297364 349064
rect 297416 349052 297422 349104
rect 282822 347692 282828 347744
rect 282880 347732 282886 347744
rect 294598 347732 294604 347744
rect 282880 347704 294604 347732
rect 282880 347692 282886 347704
rect 294598 347692 294604 347704
rect 294656 347692 294662 347744
rect 282270 347624 282276 347676
rect 282328 347664 282334 347676
rect 291838 347664 291844 347676
rect 282328 347636 291844 347664
rect 282328 347624 282334 347636
rect 291838 347624 291844 347636
rect 291896 347624 291902 347676
rect 282086 346332 282092 346384
rect 282144 346372 282150 346384
rect 290458 346372 290464 346384
rect 282144 346344 290464 346372
rect 282144 346332 282150 346344
rect 290458 346332 290464 346344
rect 290516 346332 290522 346384
rect 282822 344496 282828 344548
rect 282880 344536 282886 344548
rect 287698 344536 287704 344548
rect 282880 344508 287704 344536
rect 282880 344496 282886 344508
rect 287698 344496 287704 344508
rect 287756 344496 287762 344548
rect 282546 343544 282552 343596
rect 282604 343584 282610 343596
rect 301498 343584 301504 343596
rect 282604 343556 301504 343584
rect 282604 343544 282610 343556
rect 301498 343544 301504 343556
rect 301556 343544 301562 343596
rect 282730 343476 282736 343528
rect 282788 343516 282794 343528
rect 286318 343516 286324 343528
rect 282788 343488 286324 343516
rect 282788 343476 282794 343488
rect 286318 343476 286324 343488
rect 286376 343476 286382 343528
rect 282822 342184 282828 342236
rect 282880 342224 282886 342236
rect 316034 342224 316040 342236
rect 282880 342196 316040 342224
rect 282880 342184 282886 342196
rect 316034 342184 316040 342196
rect 316092 342184 316098 342236
rect 3418 338036 3424 338088
rect 3476 338076 3482 338088
rect 57422 338076 57428 338088
rect 3476 338048 57428 338076
rect 3476 338036 3482 338048
rect 57422 338036 57428 338048
rect 57480 338036 57486 338088
rect 57790 336676 57796 336728
rect 57848 336716 57854 336728
rect 59722 336716 59728 336728
rect 57848 336688 59728 336716
rect 57848 336676 57854 336688
rect 59722 336676 59728 336688
rect 59780 336676 59786 336728
rect 282178 333888 282184 333940
rect 282236 333928 282242 333940
rect 307018 333928 307024 333940
rect 282236 333900 307024 333928
rect 282236 333888 282242 333900
rect 307018 333888 307024 333900
rect 307076 333888 307082 333940
rect 281626 333548 281632 333600
rect 281684 333588 281690 333600
rect 283834 333588 283840 333600
rect 281684 333560 283840 333588
rect 281684 333548 281690 333560
rect 283834 333548 283840 333560
rect 283892 333548 283898 333600
rect 281994 331780 282000 331832
rect 282052 331820 282058 331832
rect 282730 331820 282736 331832
rect 282052 331792 282736 331820
rect 282052 331780 282058 331792
rect 282730 331780 282736 331792
rect 282788 331780 282794 331832
rect 281626 331168 281632 331220
rect 281684 331208 281690 331220
rect 320266 331208 320272 331220
rect 281684 331180 320272 331208
rect 281684 331168 281690 331180
rect 320266 331168 320272 331180
rect 320324 331168 320330 331220
rect 56962 330828 56968 330880
rect 57020 330868 57026 330880
rect 59814 330868 59820 330880
rect 57020 330840 59820 330868
rect 57020 330828 57026 330840
rect 59814 330828 59820 330840
rect 59872 330828 59878 330880
rect 56594 330760 56600 330812
rect 56652 330800 56658 330812
rect 56652 330772 57100 330800
rect 56652 330760 56658 330772
rect 56594 330624 56600 330676
rect 56652 330664 56658 330676
rect 56870 330664 56876 330676
rect 56652 330636 56876 330664
rect 56652 330624 56658 330636
rect 56870 330624 56876 330636
rect 56928 330624 56934 330676
rect 57072 330472 57100 330772
rect 57054 330420 57060 330472
rect 57112 330420 57118 330472
rect 281626 329740 281632 329792
rect 281684 329780 281690 329792
rect 318794 329780 318800 329792
rect 281684 329752 318800 329780
rect 281684 329740 281690 329752
rect 318794 329740 318800 329752
rect 318852 329740 318858 329792
rect 281534 329672 281540 329724
rect 281592 329712 281598 329724
rect 297450 329712 297456 329724
rect 281592 329684 297456 329712
rect 281592 329672 281598 329684
rect 297450 329672 297456 329684
rect 297508 329672 297514 329724
rect 56962 329332 56968 329384
rect 57020 329372 57026 329384
rect 57790 329372 57796 329384
rect 57020 329344 57796 329372
rect 57020 329332 57026 329344
rect 57790 329332 57796 329344
rect 57848 329332 57854 329384
rect 57054 329196 57060 329248
rect 57112 329236 57118 329248
rect 57790 329236 57796 329248
rect 57112 329208 57796 329236
rect 57112 329196 57118 329208
rect 57790 329196 57796 329208
rect 57848 329196 57854 329248
rect 281534 328380 281540 328432
rect 281592 328420 281598 328432
rect 302878 328420 302884 328432
rect 281592 328392 302884 328420
rect 281592 328380 281598 328392
rect 302878 328380 302884 328392
rect 302936 328380 302942 328432
rect 281534 327020 281540 327072
rect 281592 327060 281598 327072
rect 318242 327060 318248 327072
rect 281592 327032 318248 327060
rect 281592 327020 281598 327032
rect 318242 327020 318248 327032
rect 318300 327020 318306 327072
rect 282086 326408 282092 326460
rect 282144 326448 282150 326460
rect 282730 326448 282736 326460
rect 282144 326420 282736 326448
rect 282144 326408 282150 326420
rect 282730 326408 282736 326420
rect 282788 326408 282794 326460
rect 281902 326340 281908 326392
rect 281960 326380 281966 326392
rect 282178 326380 282184 326392
rect 281960 326352 282184 326380
rect 281960 326340 281966 326352
rect 282178 326340 282184 326352
rect 282236 326340 282242 326392
rect 282270 326340 282276 326392
rect 282328 326380 282334 326392
rect 282638 326380 282644 326392
rect 282328 326352 282644 326380
rect 282328 326340 282334 326352
rect 282638 326340 282644 326352
rect 282696 326340 282702 326392
rect 281810 326272 281816 326324
rect 281868 326312 281874 326324
rect 282730 326312 282736 326324
rect 281868 326284 282736 326312
rect 281868 326272 281874 326284
rect 282730 326272 282736 326284
rect 282788 326272 282794 326324
rect 281534 325592 281540 325644
rect 281592 325632 281598 325644
rect 318150 325632 318156 325644
rect 281592 325604 318156 325632
rect 281592 325592 281598 325604
rect 318150 325592 318156 325604
rect 318208 325592 318214 325644
rect 56594 325456 56600 325508
rect 56652 325496 56658 325508
rect 57974 325496 57980 325508
rect 56652 325468 57980 325496
rect 56652 325456 56658 325468
rect 57974 325456 57980 325468
rect 58032 325456 58038 325508
rect 56594 325320 56600 325372
rect 56652 325360 56658 325372
rect 56870 325360 56876 325372
rect 56652 325332 56876 325360
rect 56652 325320 56658 325332
rect 56870 325320 56876 325332
rect 56928 325320 56934 325372
rect 56870 325184 56876 325236
rect 56928 325224 56934 325236
rect 57514 325224 57520 325236
rect 56928 325196 57520 325224
rect 56928 325184 56934 325196
rect 57514 325184 57520 325196
rect 57572 325184 57578 325236
rect 57882 325116 57888 325168
rect 57940 325156 57946 325168
rect 59538 325156 59544 325168
rect 57940 325128 59544 325156
rect 57940 325116 57946 325128
rect 59538 325116 59544 325128
rect 59596 325116 59602 325168
rect 57698 325048 57704 325100
rect 57756 325088 57762 325100
rect 59630 325088 59636 325100
rect 57756 325060 59636 325088
rect 57756 325048 57762 325060
rect 59630 325048 59636 325060
rect 59688 325048 59694 325100
rect 3234 324232 3240 324284
rect 3292 324272 3298 324284
rect 32398 324272 32404 324284
rect 3292 324244 32404 324272
rect 3292 324232 3298 324244
rect 32398 324232 32404 324244
rect 32456 324232 32462 324284
rect 281534 324232 281540 324284
rect 281592 324272 281598 324284
rect 318058 324272 318064 324284
rect 281592 324244 318064 324272
rect 281592 324232 281598 324244
rect 318058 324232 318064 324244
rect 318116 324232 318122 324284
rect 281534 322872 281540 322924
rect 281592 322912 281598 322924
rect 305638 322912 305644 322924
rect 281592 322884 305644 322912
rect 281592 322872 281598 322884
rect 305638 322872 305644 322884
rect 305696 322872 305702 322924
rect 284294 322192 284300 322244
rect 284352 322232 284358 322244
rect 285582 322232 285588 322244
rect 284352 322204 285588 322232
rect 284352 322192 284358 322204
rect 285582 322192 285588 322204
rect 285640 322232 285646 322244
rect 337746 322232 337752 322244
rect 285640 322204 337752 322232
rect 285640 322192 285646 322204
rect 337746 322192 337752 322204
rect 337804 322192 337810 322244
rect 282822 321512 282828 321564
rect 282880 321552 282886 321564
rect 284294 321552 284300 321564
rect 282880 321524 284300 321552
rect 282880 321512 282886 321524
rect 284294 321512 284300 321524
rect 284352 321512 284358 321564
rect 282822 320968 282828 321020
rect 282880 321008 282886 321020
rect 337378 321008 337384 321020
rect 282880 320980 337384 321008
rect 282880 320968 282886 320980
rect 337378 320968 337384 320980
rect 337436 321008 337442 321020
rect 338022 321008 338028 321020
rect 337436 320980 338028 321008
rect 337436 320968 337442 320980
rect 338022 320968 338028 320980
rect 338080 320968 338086 321020
rect 282178 320900 282184 320952
rect 282236 320940 282242 320952
rect 419534 320940 419540 320952
rect 282236 320912 419540 320940
rect 282236 320900 282242 320912
rect 419534 320900 419540 320912
rect 419592 320900 419598 320952
rect 282546 320832 282552 320884
rect 282604 320872 282610 320884
rect 419810 320872 419816 320884
rect 282604 320844 419816 320872
rect 282604 320832 282610 320844
rect 419810 320832 419816 320844
rect 419868 320832 419874 320884
rect 56594 320764 56600 320816
rect 56652 320804 56658 320816
rect 580902 320804 580908 320816
rect 56652 320776 580908 320804
rect 56652 320764 56658 320776
rect 580902 320764 580908 320776
rect 580960 320764 580966 320816
rect 57974 320696 57980 320748
rect 58032 320736 58038 320748
rect 580166 320736 580172 320748
rect 58032 320708 580172 320736
rect 58032 320696 58038 320708
rect 580166 320696 580172 320708
rect 580224 320696 580230 320748
rect 57514 320628 57520 320680
rect 57572 320668 57578 320680
rect 580718 320668 580724 320680
rect 57572 320640 580724 320668
rect 57572 320628 57578 320640
rect 580718 320628 580724 320640
rect 580776 320628 580782 320680
rect 57606 320560 57612 320612
rect 57664 320600 57670 320612
rect 280062 320600 280068 320612
rect 57664 320572 280068 320600
rect 57664 320560 57670 320572
rect 280062 320560 280068 320572
rect 280120 320560 280126 320612
rect 282362 320560 282368 320612
rect 282420 320600 282426 320612
rect 419718 320600 419724 320612
rect 282420 320572 419724 320600
rect 282420 320560 282426 320572
rect 419718 320560 419724 320572
rect 419776 320560 419782 320612
rect 59538 320492 59544 320544
rect 59596 320532 59602 320544
rect 279970 320532 279976 320544
rect 59596 320504 279976 320532
rect 59596 320492 59602 320504
rect 279970 320492 279976 320504
rect 280028 320492 280034 320544
rect 281994 320492 282000 320544
rect 282052 320532 282058 320544
rect 419626 320532 419632 320544
rect 282052 320504 419632 320532
rect 282052 320492 282058 320504
rect 419626 320492 419632 320504
rect 419684 320492 419690 320544
rect 59722 320424 59728 320476
rect 59780 320464 59786 320476
rect 280062 320464 280068 320476
rect 59780 320436 280068 320464
rect 59780 320424 59786 320436
rect 280062 320424 280068 320436
rect 280120 320424 280126 320476
rect 282454 320424 282460 320476
rect 282512 320464 282518 320476
rect 416406 320464 416412 320476
rect 282512 320436 416412 320464
rect 282512 320424 282518 320436
rect 416406 320424 416412 320436
rect 416464 320424 416470 320476
rect 282270 320356 282276 320408
rect 282328 320396 282334 320408
rect 420178 320396 420184 320408
rect 282328 320368 420184 320396
rect 282328 320356 282334 320368
rect 420178 320356 420184 320368
rect 420236 320356 420242 320408
rect 282730 320288 282736 320340
rect 282788 320328 282794 320340
rect 419902 320328 419908 320340
rect 282788 320300 419908 320328
rect 282788 320288 282794 320300
rect 419902 320288 419908 320300
rect 419960 320288 419966 320340
rect 282086 320220 282092 320272
rect 282144 320260 282150 320272
rect 419994 320260 420000 320272
rect 282144 320232 420000 320260
rect 282144 320220 282150 320232
rect 419994 320220 420000 320232
rect 420052 320220 420058 320272
rect 56870 320084 56876 320136
rect 56928 320124 56934 320136
rect 580810 320124 580816 320136
rect 56928 320096 580816 320124
rect 56928 320084 56934 320096
rect 580810 320084 580816 320096
rect 580868 320084 580874 320136
rect 59814 320016 59820 320068
rect 59872 320056 59878 320068
rect 580626 320056 580632 320068
rect 59872 320028 580632 320056
rect 59872 320016 59878 320028
rect 580626 320016 580632 320028
rect 580684 320016 580690 320068
rect 59630 319948 59636 320000
rect 59688 319988 59694 320000
rect 580442 319988 580448 320000
rect 59688 319960 580448 319988
rect 59688 319948 59694 319960
rect 580442 319948 580448 319960
rect 580500 319948 580506 320000
rect 59906 319880 59912 319932
rect 59964 319920 59970 319932
rect 580350 319920 580356 319932
rect 59964 319892 580356 319920
rect 59964 319880 59970 319892
rect 580350 319880 580356 319892
rect 580408 319880 580414 319932
rect 4062 318724 4068 318776
rect 4120 318764 4126 318776
rect 64782 318764 64788 318776
rect 4120 318736 64788 318764
rect 4120 318724 4126 318736
rect 64782 318724 64788 318736
rect 64840 318724 64846 318776
rect 82722 318724 82728 318776
rect 82780 318764 82786 318776
rect 193214 318764 193220 318776
rect 82780 318736 193220 318764
rect 82780 318724 82786 318736
rect 193214 318724 193220 318736
rect 193272 318724 193278 318776
rect 338022 318724 338028 318776
rect 338080 318764 338086 318776
rect 344002 318764 344008 318776
rect 338080 318736 344008 318764
rect 338080 318724 338086 318736
rect 344002 318724 344008 318736
rect 344060 318724 344066 318776
rect 50430 318656 50436 318708
rect 50488 318696 50494 318708
rect 88150 318696 88156 318708
rect 50488 318668 88156 318696
rect 50488 318656 50494 318668
rect 88150 318656 88156 318668
rect 88208 318656 88214 318708
rect 88242 318656 88248 318708
rect 88300 318696 88306 318708
rect 201034 318696 201040 318708
rect 88300 318668 201040 318696
rect 88300 318656 88306 318668
rect 201034 318656 201040 318668
rect 201092 318656 201098 318708
rect 8202 318588 8208 318640
rect 8260 318628 8266 318640
rect 72510 318628 72516 318640
rect 8260 318600 72516 318628
rect 8260 318588 8266 318600
rect 72510 318588 72516 318600
rect 72568 318588 72574 318640
rect 204898 318628 204904 318640
rect 75196 318600 84884 318628
rect 45462 318520 45468 318572
rect 45520 318560 45526 318572
rect 55214 318560 55220 318572
rect 45520 318532 55220 318560
rect 45520 318520 45526 318532
rect 55214 318520 55220 318532
rect 55272 318520 55278 318572
rect 64782 318520 64788 318572
rect 64840 318560 64846 318572
rect 75196 318560 75224 318600
rect 64840 318532 75224 318560
rect 84856 318560 84884 318600
rect 94516 318600 204904 318628
rect 94406 318560 94412 318572
rect 84856 318532 94412 318560
rect 64840 318520 64846 318532
rect 94406 318520 94412 318532
rect 94464 318520 94470 318572
rect 10962 318452 10968 318504
rect 11020 318492 11026 318504
rect 76466 318492 76472 318504
rect 11020 318464 76472 318492
rect 11020 318452 11026 318464
rect 76466 318452 76472 318464
rect 76524 318452 76530 318504
rect 86862 318452 86868 318504
rect 86920 318492 86926 318504
rect 88242 318492 88248 318504
rect 86920 318464 88248 318492
rect 86920 318452 86926 318464
rect 88242 318452 88248 318464
rect 88300 318452 88306 318504
rect 89530 318452 89536 318504
rect 89588 318492 89594 318504
rect 94516 318492 94544 318600
rect 204898 318588 204904 318600
rect 204956 318588 204962 318640
rect 94590 318520 94596 318572
rect 94648 318560 94654 318572
rect 212718 318560 212724 318572
rect 94648 318532 212724 318560
rect 94648 318520 94654 318532
rect 212718 318520 212724 318532
rect 212776 318520 212782 318572
rect 89588 318464 94544 318492
rect 89588 318452 89594 318464
rect 96522 318452 96528 318504
rect 96580 318492 96586 318504
rect 216582 318492 216588 318504
rect 96580 318464 216588 318492
rect 96580 318452 96586 318464
rect 216582 318452 216588 318464
rect 216640 318452 216646 318504
rect 42702 318384 42708 318436
rect 42760 318424 42766 318436
rect 128998 318424 129004 318436
rect 42760 318396 129004 318424
rect 42760 318384 42766 318396
rect 128998 318384 129004 318396
rect 129056 318384 129062 318436
rect 134518 318384 134524 318436
rect 134576 318424 134582 318436
rect 255498 318424 255504 318436
rect 134576 318396 255504 318424
rect 134576 318384 134582 318396
rect 255498 318384 255504 318396
rect 255556 318384 255562 318436
rect 16482 318316 16488 318368
rect 16540 318356 16546 318368
rect 86218 318356 86224 318368
rect 16540 318328 86224 318356
rect 16540 318316 16546 318328
rect 86218 318316 86224 318328
rect 86276 318316 86282 318368
rect 94406 318316 94412 318368
rect 94464 318356 94470 318368
rect 107562 318356 107568 318368
rect 94464 318328 107568 318356
rect 94464 318316 94470 318328
rect 107562 318316 107568 318328
rect 107620 318316 107626 318368
rect 107654 318316 107660 318368
rect 107712 318356 107718 318368
rect 224402 318356 224408 318368
rect 107712 318328 224408 318356
rect 107712 318316 107718 318328
rect 224402 318316 224408 318328
rect 224460 318316 224466 318368
rect 20622 318248 20628 318300
rect 20680 318288 20686 318300
rect 92014 318288 92020 318300
rect 20680 318260 92020 318288
rect 20680 318248 20686 318260
rect 92014 318248 92020 318260
rect 92072 318248 92078 318300
rect 93762 318248 93768 318300
rect 93820 318288 93826 318300
rect 94590 318288 94596 318300
rect 93820 318260 94596 318288
rect 93820 318248 93826 318260
rect 94590 318248 94596 318260
rect 94648 318248 94654 318300
rect 103422 318248 103428 318300
rect 103480 318288 103486 318300
rect 228266 318288 228272 318300
rect 103480 318260 228272 318288
rect 103480 318248 103486 318260
rect 228266 318248 228272 318260
rect 228324 318248 228330 318300
rect 21910 318180 21916 318232
rect 21968 318220 21974 318232
rect 93946 318220 93952 318232
rect 21968 318192 93952 318220
rect 21968 318180 21974 318192
rect 93946 318180 93952 318192
rect 94004 318180 94010 318232
rect 107562 318180 107568 318232
rect 107620 318220 107626 318232
rect 234154 318220 234160 318232
rect 107620 318192 234160 318220
rect 107620 318180 107626 318192
rect 234154 318180 234160 318192
rect 234212 318180 234218 318232
rect 24762 318112 24768 318164
rect 24820 318152 24826 318164
rect 99834 318152 99840 318164
rect 24820 318124 99840 318152
rect 24820 318112 24826 318124
rect 99834 318112 99840 318124
rect 99892 318112 99898 318164
rect 100662 318112 100668 318164
rect 100720 318152 100726 318164
rect 100720 318124 101996 318152
rect 100720 318112 100726 318124
rect 26142 318044 26148 318096
rect 26200 318084 26206 318096
rect 101766 318084 101772 318096
rect 26200 318056 101772 318084
rect 26200 318044 26206 318056
rect 101766 318044 101772 318056
rect 101824 318044 101830 318096
rect 101968 318084 101996 318124
rect 107470 318112 107476 318164
rect 107528 318152 107534 318164
rect 236086 318152 236092 318164
rect 107528 318124 236092 318152
rect 107528 318112 107534 318124
rect 236086 318112 236092 318124
rect 236144 318112 236150 318164
rect 107654 318084 107660 318096
rect 101968 318056 107660 318084
rect 107654 318044 107660 318056
rect 107712 318044 107718 318096
rect 114462 318044 114468 318096
rect 114520 318084 114526 318096
rect 245838 318084 245844 318096
rect 114520 318056 245844 318084
rect 114520 318044 114526 318056
rect 245838 318044 245844 318056
rect 245896 318044 245902 318096
rect 344002 318044 344008 318096
rect 344060 318084 344066 318096
rect 347774 318084 347780 318096
rect 344060 318056 347780 318084
rect 344060 318044 344066 318056
rect 347774 318044 347780 318056
rect 347832 318044 347838 318096
rect 32398 317976 32404 318028
rect 32456 318016 32462 318028
rect 78398 318016 78404 318028
rect 32456 317988 78404 318016
rect 32456 317976 32462 317988
rect 78398 317976 78404 317988
rect 78456 317976 78462 318028
rect 79962 317976 79968 318028
rect 80020 318016 80026 318028
rect 189350 318016 189356 318028
rect 80020 317988 189356 318016
rect 80020 317976 80026 317988
rect 189350 317976 189356 317988
rect 189408 317976 189414 318028
rect 39298 317908 39304 317960
rect 39356 317948 39362 317960
rect 68646 317948 68652 317960
rect 39356 317920 68652 317948
rect 39356 317908 39362 317920
rect 68646 317908 68652 317920
rect 68704 317908 68710 317960
rect 74442 317908 74448 317960
rect 74500 317948 74506 317960
rect 181530 317948 181536 317960
rect 74500 317920 181536 317948
rect 74500 317908 74506 317920
rect 181530 317908 181536 317920
rect 181588 317908 181594 317960
rect 2682 317840 2688 317892
rect 2740 317880 2746 317892
rect 62850 317880 62856 317892
rect 2740 317852 62856 317880
rect 2740 317840 2746 317852
rect 62850 317840 62856 317852
rect 62908 317840 62914 317892
rect 64782 317840 64788 317892
rect 64840 317840 64846 317892
rect 72970 317840 72976 317892
rect 73028 317880 73034 317892
rect 177666 317880 177672 317892
rect 73028 317852 177672 317880
rect 73028 317840 73034 317852
rect 177666 317840 177672 317852
rect 177724 317840 177730 317892
rect 42058 317772 42064 317824
rect 42116 317812 42122 317824
rect 45462 317812 45468 317824
rect 42116 317784 45468 317812
rect 42116 317772 42122 317784
rect 45462 317772 45468 317784
rect 45520 317772 45526 317824
rect 55214 317772 55220 317824
rect 55272 317812 55278 317824
rect 64800 317812 64828 317840
rect 55272 317784 64828 317812
rect 55272 317772 55278 317784
rect 67542 317772 67548 317824
rect 67600 317812 67606 317824
rect 169846 317812 169852 317824
rect 67600 317784 169852 317812
rect 67600 317772 67606 317784
rect 169846 317772 169852 317784
rect 169904 317772 169910 317824
rect 64782 317704 64788 317756
rect 64840 317744 64846 317756
rect 165982 317744 165988 317756
rect 64840 317716 165988 317744
rect 64840 317704 64846 317716
rect 165982 317704 165988 317716
rect 166040 317704 166046 317756
rect 62022 317636 62028 317688
rect 62080 317676 62086 317688
rect 160186 317676 160192 317688
rect 62080 317648 160192 317676
rect 62080 317636 62086 317648
rect 160186 317636 160192 317648
rect 160244 317636 160250 317688
rect 50982 317568 50988 317620
rect 51040 317608 51046 317620
rect 142614 317608 142620 317620
rect 51040 317580 142620 317608
rect 51040 317568 51046 317580
rect 142614 317568 142620 317580
rect 142672 317568 142678 317620
rect 48130 317500 48136 317552
rect 48188 317540 48194 317552
rect 136818 317540 136824 317552
rect 48188 317512 136824 317540
rect 48188 317500 48194 317512
rect 136818 317500 136824 317512
rect 136876 317500 136882 317552
rect 39942 317432 39948 317484
rect 40000 317472 40006 317484
rect 124766 317472 124772 317484
rect 40000 317444 124772 317472
rect 40000 317432 40006 317444
rect 124766 317432 124772 317444
rect 124824 317432 124830 317484
rect 124858 317432 124864 317484
rect 124916 317472 124922 317484
rect 146570 317472 146576 317484
rect 124916 317444 146576 317472
rect 124916 317432 124922 317444
rect 146570 317432 146576 317444
rect 146628 317432 146634 317484
rect 56686 311788 56692 311840
rect 56744 311828 56750 311840
rect 580166 311828 580172 311840
rect 56744 311800 580172 311828
rect 56744 311788 56750 311800
rect 580166 311788 580172 311800
rect 580224 311788 580230 311840
rect 3326 309068 3332 309120
rect 3384 309108 3390 309120
rect 20070 309108 20076 309120
rect 3384 309080 20076 309108
rect 3384 309068 3390 309080
rect 20070 309068 20076 309080
rect 20128 309068 20134 309120
rect 74442 299616 74448 299668
rect 74500 299616 74506 299668
rect 74460 299532 74488 299616
rect 74442 299480 74448 299532
rect 74500 299480 74506 299532
rect 56778 299412 56784 299464
rect 56836 299452 56842 299464
rect 579798 299452 579804 299464
rect 56836 299424 579804 299452
rect 56836 299412 56842 299424
rect 579798 299412 579804 299424
rect 579856 299412 579862 299464
rect 74258 298052 74264 298104
rect 74316 298092 74322 298104
rect 74442 298092 74448 298104
rect 74316 298064 74448 298092
rect 74316 298052 74322 298064
rect 74442 298052 74448 298064
rect 74500 298052 74506 298104
rect 3418 295264 3424 295316
rect 3476 295304 3482 295316
rect 57330 295304 57336 295316
rect 3476 295276 57336 295304
rect 3476 295264 3482 295276
rect 57330 295264 57336 295276
rect 57388 295264 57394 295316
rect 74258 288396 74264 288448
rect 74316 288436 74322 288448
rect 74350 288436 74356 288448
rect 74316 288408 74356 288436
rect 74316 288396 74322 288408
rect 74350 288396 74356 288408
rect 74408 288396 74414 288448
rect 3418 280100 3424 280152
rect 3476 280140 3482 280152
rect 37918 280140 37924 280152
rect 3476 280112 37924 280140
rect 3476 280100 3482 280112
rect 37918 280100 37924 280112
rect 37976 280100 37982 280152
rect 57146 275952 57152 276004
rect 57204 275992 57210 276004
rect 580166 275992 580172 276004
rect 57204 275964 580172 275992
rect 57204 275952 57210 275964
rect 580166 275952 580172 275964
rect 580224 275952 580230 276004
rect 74258 269084 74264 269136
rect 74316 269124 74322 269136
rect 74350 269124 74356 269136
rect 74316 269096 74356 269124
rect 74316 269084 74322 269096
rect 74350 269084 74356 269096
rect 74408 269084 74414 269136
rect 2866 266296 2872 266348
rect 2924 266336 2930 266348
rect 28350 266336 28356 266348
rect 2924 266308 28356 266336
rect 2924 266296 2930 266308
rect 28350 266296 28356 266308
rect 28408 266296 28414 266348
rect 147582 263780 147588 263832
rect 147640 263820 147646 263832
rect 154482 263820 154488 263832
rect 147640 263792 154488 263820
rect 147640 263780 147646 263792
rect 154482 263780 154488 263792
rect 154540 263780 154546 263832
rect 86862 263712 86868 263764
rect 86920 263712 86926 263764
rect 86880 263628 86908 263712
rect 115934 263644 115940 263696
rect 115992 263684 115998 263696
rect 118786 263684 118792 263696
rect 115992 263656 118792 263684
rect 115992 263644 115998 263656
rect 118786 263644 118792 263656
rect 118844 263644 118850 263696
rect 86862 263576 86868 263628
rect 86920 263576 86926 263628
rect 3418 252492 3424 252544
rect 3476 252532 3482 252544
rect 57238 252532 57244 252544
rect 3476 252504 57244 252532
rect 3476 252492 3482 252504
rect 57238 252492 57244 252504
rect 57296 252492 57302 252544
rect 59446 252492 59452 252544
rect 59504 252532 59510 252544
rect 579798 252532 579804 252544
rect 59504 252504 579804 252532
rect 59504 252492 59510 252504
rect 579798 252492 579804 252504
rect 579856 252492 579862 252544
rect 74258 249772 74264 249824
rect 74316 249812 74322 249824
rect 74442 249812 74448 249824
rect 74316 249784 74448 249812
rect 74316 249772 74322 249784
rect 74442 249772 74448 249784
rect 74500 249772 74506 249824
rect 74350 241476 74356 241528
rect 74408 241516 74414 241528
rect 74442 241516 74448 241528
rect 74408 241488 74448 241516
rect 74408 241476 74414 241488
rect 74442 241476 74448 241488
rect 74500 241476 74506 241528
rect 3418 237328 3424 237380
rect 3476 237368 3482 237380
rect 39390 237368 39396 237380
rect 3476 237340 39396 237368
rect 3476 237328 3482 237340
rect 39390 237328 39396 237340
rect 39448 237328 39454 237380
rect 74258 230460 74264 230512
rect 74316 230500 74322 230512
rect 74442 230500 74448 230512
rect 74316 230472 74448 230500
rect 74316 230460 74322 230472
rect 74442 230460 74448 230472
rect 74500 230460 74506 230512
rect 66254 227944 66260 227996
rect 66312 227984 66318 227996
rect 75822 227984 75828 227996
rect 66312 227956 75828 227984
rect 66312 227944 66318 227956
rect 75822 227944 75828 227956
rect 75880 227944 75886 227996
rect 147582 227876 147588 227928
rect 147640 227916 147646 227928
rect 154482 227916 154488 227928
rect 147640 227888 154488 227916
rect 147640 227876 147646 227888
rect 154482 227876 154488 227888
rect 154540 227876 154546 227928
rect 86862 227808 86868 227860
rect 86920 227808 86926 227860
rect 86880 227724 86908 227808
rect 115934 227740 115940 227792
rect 115992 227780 115998 227792
rect 118786 227780 118792 227792
rect 115992 227752 118792 227780
rect 115992 227740 115998 227752
rect 118786 227740 118792 227752
rect 118844 227740 118850 227792
rect 86862 227672 86868 227724
rect 86920 227672 86926 227724
rect 3142 223524 3148 223576
rect 3200 223564 3206 223576
rect 33870 223564 33876 223576
rect 3200 223536 33876 223564
rect 3200 223524 3206 223536
rect 33870 223524 33876 223536
rect 33928 223524 33934 223576
rect 69382 216928 69388 216980
rect 69440 216968 69446 216980
rect 77202 216968 77208 216980
rect 69440 216940 77208 216968
rect 69440 216928 69446 216940
rect 77202 216928 77208 216940
rect 77260 216928 77266 216980
rect 89530 216860 89536 216912
rect 89588 216900 89594 216912
rect 91738 216900 91744 216912
rect 89588 216872 91744 216900
rect 89588 216860 89594 216872
rect 91738 216860 91744 216872
rect 91796 216860 91802 216912
rect 147582 216860 147588 216912
rect 147640 216900 147646 216912
rect 154482 216900 154488 216912
rect 147640 216872 154488 216900
rect 147640 216860 147646 216872
rect 154482 216860 154488 216872
rect 154540 216860 154546 216912
rect 115934 216724 115940 216776
rect 115992 216764 115998 216776
rect 118786 216764 118792 216776
rect 115992 216736 118792 216764
rect 115992 216724 115998 216736
rect 118786 216724 118792 216736
rect 118844 216724 118850 216776
rect 2774 208156 2780 208208
rect 2832 208196 2838 208208
rect 5074 208196 5080 208208
rect 2832 208168 5080 208196
rect 2832 208156 2838 208168
rect 5074 208156 5080 208168
rect 5132 208156 5138 208208
rect 59354 205572 59360 205624
rect 59412 205612 59418 205624
rect 579798 205612 579804 205624
rect 59412 205584 579804 205612
rect 59412 205572 59418 205584
rect 579798 205572 579804 205584
rect 579856 205572 579862 205624
rect 89346 202852 89352 202904
rect 89404 202892 89410 202904
rect 89530 202892 89536 202904
rect 89404 202864 89536 202892
rect 89404 202852 89410 202864
rect 89530 202852 89536 202864
rect 89588 202852 89594 202904
rect 74258 201424 74264 201476
rect 74316 201464 74322 201476
rect 74442 201464 74448 201476
rect 74316 201436 74448 201464
rect 74316 201424 74322 201436
rect 74442 201424 74448 201436
rect 74500 201424 74506 201476
rect 89346 195984 89352 196036
rect 89404 195984 89410 196036
rect 89364 195888 89392 195984
rect 89438 195888 89444 195900
rect 89364 195860 89444 195888
rect 89438 195848 89444 195860
rect 89496 195848 89502 195900
rect 2866 194488 2872 194540
rect 2924 194528 2930 194540
rect 50338 194528 50344 194540
rect 2924 194500 50344 194528
rect 2924 194488 2930 194500
rect 50338 194488 50344 194500
rect 50396 194488 50402 194540
rect 74258 191836 74264 191888
rect 74316 191876 74322 191888
rect 74350 191876 74356 191888
rect 74316 191848 74356 191876
rect 74316 191836 74322 191848
rect 74350 191836 74356 191848
rect 74408 191836 74414 191888
rect 74350 183540 74356 183592
rect 74408 183580 74414 183592
rect 74442 183580 74448 183592
rect 74408 183552 74448 183580
rect 74408 183540 74414 183552
rect 74442 183540 74448 183552
rect 74500 183540 74506 183592
rect 74258 182112 74264 182164
rect 74316 182152 74322 182164
rect 74442 182152 74448 182164
rect 74316 182124 74448 182152
rect 74316 182112 74322 182124
rect 74442 182112 74448 182124
rect 74500 182112 74506 182164
rect 69382 181024 69388 181076
rect 69440 181064 69446 181076
rect 77202 181064 77208 181076
rect 69440 181036 77208 181064
rect 69440 181024 69446 181036
rect 77202 181024 77208 181036
rect 77260 181024 77266 181076
rect 86862 180888 86868 180940
rect 86920 180888 86926 180940
rect 86880 180804 86908 180888
rect 3234 180752 3240 180804
rect 3292 180792 3298 180804
rect 35158 180792 35164 180804
rect 3292 180764 35164 180792
rect 3292 180752 3298 180764
rect 35158 180752 35164 180764
rect 35216 180752 35222 180804
rect 86862 180752 86868 180804
rect 86920 180752 86926 180804
rect 89438 173884 89444 173936
rect 89496 173924 89502 173936
rect 89622 173924 89628 173936
rect 89496 173896 89628 173924
rect 89496 173884 89502 173896
rect 89622 173884 89628 173896
rect 89680 173884 89686 173936
rect 66254 170008 66260 170060
rect 66312 170048 66318 170060
rect 75822 170048 75828 170060
rect 66312 170020 75828 170048
rect 66312 170008 66318 170020
rect 75822 170008 75828 170020
rect 75880 170008 75886 170060
rect 147582 169940 147588 169992
rect 147640 169980 147646 169992
rect 154482 169980 154488 169992
rect 147640 169952 154488 169980
rect 147640 169940 147646 169952
rect 154482 169940 154488 169952
rect 154540 169940 154546 169992
rect 86862 169872 86868 169924
rect 86920 169872 86926 169924
rect 86880 169788 86908 169872
rect 115934 169804 115940 169856
rect 115992 169844 115998 169856
rect 118786 169844 118792 169856
rect 115992 169816 118792 169844
rect 115992 169804 115998 169816
rect 118786 169804 118792 169816
rect 118844 169804 118850 169856
rect 86862 169736 86868 169788
rect 86920 169736 86926 169788
rect 2774 165452 2780 165504
rect 2832 165492 2838 165504
rect 4982 165492 4988 165504
rect 2832 165464 4988 165492
rect 2832 165452 2838 165464
rect 4982 165452 4988 165464
rect 5040 165452 5046 165504
rect 74258 162800 74264 162852
rect 74316 162840 74322 162852
rect 74442 162840 74448 162852
rect 74316 162812 74448 162840
rect 74316 162800 74322 162812
rect 74442 162800 74448 162812
rect 74500 162800 74506 162852
rect 59078 158652 59084 158704
rect 59136 158692 59142 158704
rect 579798 158692 579804 158704
rect 59136 158664 579804 158692
rect 59136 158652 59142 158664
rect 579798 158652 579804 158664
rect 579856 158652 579862 158704
rect 89438 157428 89444 157480
rect 89496 157428 89502 157480
rect 89456 157344 89484 157428
rect 89438 157292 89444 157344
rect 89496 157292 89502 157344
rect 89254 154504 89260 154556
rect 89312 154544 89318 154556
rect 89530 154544 89536 154556
rect 89312 154516 89536 154544
rect 89312 154504 89318 154516
rect 89530 154504 89536 154516
rect 89588 154504 89594 154556
rect 3142 151716 3148 151768
rect 3200 151756 3206 151768
rect 51718 151756 51724 151768
rect 3200 151728 51724 151756
rect 3200 151716 3206 151728
rect 51718 151716 51724 151728
rect 51776 151716 51782 151768
rect 74442 143488 74448 143540
rect 74500 143528 74506 143540
rect 74626 143528 74632 143540
rect 74500 143500 74632 143528
rect 74500 143488 74506 143500
rect 74626 143488 74632 143500
rect 74684 143488 74690 143540
rect 89438 137980 89444 138032
rect 89496 137980 89502 138032
rect 89456 137884 89484 137980
rect 89530 137884 89536 137896
rect 89456 137856 89536 137884
rect 89530 137844 89536 137856
rect 89588 137844 89594 137896
rect 3234 136552 3240 136604
rect 3292 136592 3298 136604
rect 43438 136592 43444 136604
rect 3292 136564 43444 136592
rect 3292 136552 3298 136564
rect 43438 136552 43444 136564
rect 43496 136552 43502 136604
rect 57422 135192 57428 135244
rect 57480 135232 57486 135244
rect 580166 135232 580172 135244
rect 57480 135204 580172 135232
rect 57480 135192 57486 135204
rect 580166 135192 580172 135204
rect 580224 135192 580230 135244
rect 89530 128432 89536 128444
rect 89456 128404 89536 128432
rect 89456 128308 89484 128404
rect 89530 128392 89536 128404
rect 89588 128392 89594 128444
rect 89438 128256 89444 128308
rect 89496 128256 89502 128308
rect 56962 124108 56968 124160
rect 57020 124148 57026 124160
rect 580166 124148 580172 124160
rect 57020 124120 580172 124148
rect 57020 124108 57026 124120
rect 580166 124108 580172 124120
rect 580224 124108 580230 124160
rect 89438 124040 89444 124092
rect 89496 124080 89502 124092
rect 89622 124080 89628 124092
rect 89496 124052 89628 124080
rect 89496 124040 89502 124052
rect 89622 124040 89628 124052
rect 89680 124040 89686 124092
rect 2774 122340 2780 122392
rect 2832 122380 2838 122392
rect 4890 122380 4896 122392
rect 2832 122352 4896 122380
rect 2832 122340 2838 122352
rect 4890 122340 4896 122352
rect 4948 122340 4954 122392
rect 89622 118668 89628 118720
rect 89680 118668 89686 118720
rect 89530 118532 89536 118584
rect 89588 118572 89594 118584
rect 89640 118572 89668 118668
rect 89588 118544 89668 118572
rect 89588 118532 89594 118544
rect 74350 114520 74356 114572
rect 74408 114560 74414 114572
rect 74718 114560 74724 114572
rect 74408 114532 74724 114560
rect 74408 114520 74414 114532
rect 74718 114520 74724 114532
rect 74776 114520 74782 114572
rect 59170 111732 59176 111784
rect 59228 111772 59234 111784
rect 579798 111772 579804 111784
rect 59228 111744 579804 111772
rect 59228 111732 59234 111744
rect 579798 111732 579804 111744
rect 579856 111732 579862 111784
rect 89530 109120 89536 109132
rect 89456 109092 89536 109120
rect 89456 108996 89484 109092
rect 89530 109080 89536 109092
rect 89588 109080 89594 109132
rect 3234 108944 3240 108996
rect 3292 108984 3298 108996
rect 53098 108984 53104 108996
rect 3292 108956 53104 108984
rect 3292 108944 3298 108956
rect 53098 108944 53104 108956
rect 53156 108944 53162 108996
rect 89438 108944 89444 108996
rect 89496 108944 89502 108996
rect 74350 106360 74356 106412
rect 74408 106400 74414 106412
rect 74442 106400 74448 106412
rect 74408 106372 74448 106400
rect 74408 106360 74414 106372
rect 74442 106360 74448 106372
rect 74500 106360 74506 106412
rect 74258 104796 74264 104848
rect 74316 104836 74322 104848
rect 74442 104836 74448 104848
rect 74316 104808 74448 104836
rect 74316 104796 74322 104808
rect 74442 104796 74448 104808
rect 74500 104796 74506 104848
rect 89254 104796 89260 104848
rect 89312 104836 89318 104848
rect 89438 104836 89444 104848
rect 89312 104808 89444 104836
rect 89312 104796 89318 104808
rect 89438 104796 89444 104808
rect 89496 104796 89502 104848
rect 74258 95208 74264 95260
rect 74316 95248 74322 95260
rect 74350 95248 74356 95260
rect 74316 95220 74356 95248
rect 74316 95208 74322 95220
rect 74350 95208 74356 95220
rect 74408 95208 74414 95260
rect 89254 95208 89260 95260
rect 89312 95248 89318 95260
rect 89346 95248 89352 95260
rect 89312 95220 89352 95248
rect 89312 95208 89318 95220
rect 89346 95208 89352 95220
rect 89404 95208 89410 95260
rect 3418 93780 3424 93832
rect 3476 93820 3482 93832
rect 46198 93820 46204 93832
rect 3476 93792 46204 93820
rect 3476 93780 3482 93792
rect 46198 93780 46204 93792
rect 46256 93780 46262 93832
rect 57054 88272 57060 88324
rect 57112 88312 57118 88324
rect 580166 88312 580172 88324
rect 57112 88284 580172 88312
rect 57112 88272 57118 88284
rect 580166 88272 580172 88284
rect 580224 88272 580230 88324
rect 74350 87048 74356 87100
rect 74408 87088 74414 87100
rect 74442 87088 74448 87100
rect 74408 87060 74448 87088
rect 74408 87048 74414 87060
rect 74442 87048 74448 87060
rect 74500 87048 74506 87100
rect 74258 85484 74264 85536
rect 74316 85524 74322 85536
rect 74442 85524 74448 85536
rect 74316 85496 74448 85524
rect 74316 85484 74322 85496
rect 74442 85484 74448 85496
rect 74500 85484 74506 85536
rect 89530 80112 89536 80164
rect 89588 80112 89594 80164
rect 89548 80028 89576 80112
rect 89530 79976 89536 80028
rect 89588 79976 89594 80028
rect 2774 79024 2780 79076
rect 2832 79064 2838 79076
rect 4798 79064 4804 79076
rect 2832 79036 4804 79064
rect 2832 79024 2838 79036
rect 4798 79024 4804 79036
rect 4856 79024 4862 79076
rect 89622 76100 89628 76152
rect 89680 76140 89686 76152
rect 91738 76140 91744 76152
rect 89680 76112 91744 76140
rect 89680 76100 89686 76112
rect 91738 76100 91744 76112
rect 91796 76100 91802 76152
rect 147582 76100 147588 76152
rect 147640 76140 147646 76152
rect 154482 76140 154488 76152
rect 147640 76112 154488 76140
rect 147640 76100 147646 76112
rect 154482 76100 154488 76112
rect 154540 76100 154546 76152
rect 115934 75964 115940 76016
rect 115992 76004 115998 76016
rect 118786 76004 118792 76016
rect 115992 75976 118792 76004
rect 115992 75964 115998 75976
rect 118786 75964 118792 75976
rect 118844 75964 118850 76016
rect 74258 75896 74264 75948
rect 74316 75936 74322 75948
rect 74350 75936 74356 75948
rect 74316 75908 74356 75936
rect 74316 75896 74322 75908
rect 74350 75896 74356 75908
rect 74408 75896 74414 75948
rect 74350 67668 74356 67720
rect 74408 67708 74414 67720
rect 74442 67708 74448 67720
rect 74408 67680 74448 67708
rect 74408 67668 74414 67680
rect 74442 67668 74448 67680
rect 74500 67668 74506 67720
rect 74258 66172 74264 66224
rect 74316 66212 74322 66224
rect 74442 66212 74448 66224
rect 74316 66184 74448 66212
rect 74316 66172 74322 66184
rect 74442 66172 74448 66184
rect 74500 66172 74506 66224
rect 3326 64812 3332 64864
rect 3384 64852 3390 64864
rect 28258 64852 28264 64864
rect 3384 64824 28264 64852
rect 3384 64812 3390 64824
rect 28258 64812 28264 64824
rect 28316 64812 28322 64864
rect 59262 64812 59268 64864
rect 59320 64852 59326 64864
rect 579798 64852 579804 64864
rect 59320 64824 579804 64852
rect 59320 64812 59326 64824
rect 579798 64812 579804 64824
rect 579856 64812 579862 64864
rect 74258 56584 74264 56636
rect 74316 56624 74322 56636
rect 74442 56624 74448 56636
rect 74316 56596 74448 56624
rect 74316 56584 74322 56596
rect 74442 56584 74448 56596
rect 74500 56584 74506 56636
rect 3418 51008 3424 51060
rect 3476 51048 3482 51060
rect 48958 51048 48964 51060
rect 3476 51020 48964 51048
rect 3476 51008 3482 51020
rect 48958 51008 48964 51020
rect 49016 51008 49022 51060
rect 89438 51008 89444 51060
rect 89496 51048 89502 51060
rect 89622 51048 89628 51060
rect 89496 51020 89628 51048
rect 89496 51008 89502 51020
rect 89622 51008 89628 51020
rect 89680 51008 89686 51060
rect 89346 48220 89352 48272
rect 89404 48260 89410 48272
rect 89622 48260 89628 48272
rect 89404 48232 89628 48260
rect 89404 48220 89410 48232
rect 89622 48220 89628 48232
rect 89680 48220 89686 48272
rect 74258 46860 74264 46912
rect 74316 46900 74322 46912
rect 74442 46900 74448 46912
rect 74316 46872 74448 46900
rect 74316 46860 74322 46872
rect 74442 46860 74448 46872
rect 74500 46860 74506 46912
rect 57698 41352 57704 41404
rect 57756 41392 57762 41404
rect 580166 41392 580172 41404
rect 57756 41364 580172 41392
rect 57756 41352 57762 41364
rect 580166 41352 580172 41364
rect 580224 41352 580230 41404
rect 89346 38632 89352 38684
rect 89404 38672 89410 38684
rect 89530 38672 89536 38684
rect 89404 38644 89536 38672
rect 89404 38632 89410 38644
rect 89530 38632 89536 38644
rect 89588 38632 89594 38684
rect 74258 37272 74264 37324
rect 74316 37312 74322 37324
rect 74350 37312 74356 37324
rect 74316 37284 74356 37312
rect 74316 37272 74322 37284
rect 74350 37272 74356 37284
rect 74408 37272 74414 37324
rect 3418 35844 3424 35896
rect 3476 35884 3482 35896
rect 17218 35884 17224 35896
rect 3476 35856 17224 35884
rect 3476 35844 3482 35856
rect 17218 35844 17224 35856
rect 17276 35844 17282 35896
rect 57790 30268 57796 30320
rect 57848 30308 57854 30320
rect 580166 30308 580172 30320
rect 57848 30280 580172 30308
rect 57848 30268 57854 30280
rect 580166 30268 580172 30280
rect 580224 30268 580230 30320
rect 74258 27548 74264 27600
rect 74316 27588 74322 27600
rect 74442 27588 74448 27600
rect 74316 27560 74448 27588
rect 74316 27548 74322 27560
rect 74442 27548 74448 27560
rect 74500 27548 74506 27600
rect 89162 26188 89168 26240
rect 89220 26228 89226 26240
rect 89254 26228 89260 26240
rect 89220 26200 89260 26228
rect 89220 26188 89226 26200
rect 89254 26188 89260 26200
rect 89312 26188 89318 26240
rect 2866 22040 2872 22092
rect 2924 22080 2930 22092
rect 33778 22080 33784 22092
rect 2924 22052 33784 22080
rect 2924 22040 2930 22052
rect 33778 22040 33784 22052
rect 33836 22040 33842 22092
rect 89162 21360 89168 21412
rect 89220 21400 89226 21412
rect 89438 21400 89444 21412
rect 89220 21372 89444 21400
rect 89220 21360 89226 21372
rect 89438 21360 89444 21372
rect 89496 21360 89502 21412
rect 74074 17960 74080 18012
rect 74132 18000 74138 18012
rect 74258 18000 74264 18012
rect 74132 17972 74264 18000
rect 74132 17960 74138 17972
rect 74258 17960 74264 17972
rect 74316 17960 74322 18012
rect 57882 17892 57888 17944
rect 57940 17932 57946 17944
rect 579798 17932 579804 17944
rect 57940 17904 579804 17932
rect 57940 17892 57946 17904
rect 579798 17892 579804 17904
rect 579856 17892 579862 17944
rect 74074 9664 74080 9716
rect 74132 9704 74138 9716
rect 74258 9704 74264 9716
rect 74132 9676 74264 9704
rect 74132 9664 74138 9676
rect 74258 9664 74264 9676
rect 74316 9664 74322 9716
rect 89346 8304 89352 8356
rect 89404 8344 89410 8356
rect 89438 8344 89444 8356
rect 89404 8316 89444 8344
rect 89404 8304 89410 8316
rect 89438 8304 89444 8316
rect 89496 8304 89502 8356
rect 3418 8236 3424 8288
rect 3476 8276 3482 8288
rect 19978 8276 19984 8288
rect 3476 8248 19984 8276
rect 3476 8236 3482 8248
rect 19978 8236 19984 8248
rect 20036 8236 20042 8288
rect 59998 6400 60004 6452
rect 60056 6440 60062 6452
rect 157334 6440 157340 6452
rect 60056 6412 157340 6440
rect 60056 6400 60062 6412
rect 157334 6400 157340 6412
rect 157392 6400 157398 6452
rect 108758 6332 108764 6384
rect 108816 6372 108822 6384
rect 237374 6372 237380 6384
rect 108816 6344 237380 6372
rect 108816 6332 108822 6344
rect 237374 6332 237380 6344
rect 237432 6332 237438 6384
rect 112346 6264 112352 6316
rect 112404 6304 112410 6316
rect 242894 6304 242900 6316
rect 112404 6276 242900 6304
rect 112404 6264 112410 6276
rect 242894 6264 242900 6276
rect 242952 6264 242958 6316
rect 115934 6196 115940 6248
rect 115992 6236 115998 6248
rect 248414 6236 248420 6248
rect 115992 6208 248420 6236
rect 115992 6196 115998 6208
rect 248414 6196 248420 6208
rect 248472 6196 248478 6248
rect 123018 6128 123024 6180
rect 123076 6168 123082 6180
rect 260834 6168 260840 6180
rect 123076 6140 260840 6168
rect 123076 6128 123082 6140
rect 260834 6128 260840 6140
rect 260892 6128 260898 6180
rect 86126 5584 86132 5636
rect 86184 5624 86190 5636
rect 86862 5624 86868 5636
rect 86184 5596 86868 5624
rect 86184 5584 86190 5596
rect 86862 5584 86868 5596
rect 86920 5584 86926 5636
rect 93854 5516 93860 5568
rect 93912 5556 93918 5568
rect 103606 5556 103612 5568
rect 93912 5528 103612 5556
rect 93912 5516 93918 5528
rect 103606 5516 103612 5528
rect 103664 5516 103670 5568
rect 105078 5516 105084 5568
rect 105136 5556 105142 5568
rect 109034 5556 109040 5568
rect 105136 5528 109040 5556
rect 105136 5516 105142 5528
rect 109034 5516 109040 5528
rect 109092 5516 109098 5568
rect 80054 5488 80060 5500
rect 78692 5460 80060 5488
rect 60734 5380 60740 5432
rect 60792 5420 60798 5432
rect 78582 5420 78588 5432
rect 60792 5392 78588 5420
rect 60792 5380 60798 5392
rect 78582 5380 78588 5392
rect 78640 5380 78646 5432
rect 12434 5312 12440 5364
rect 12492 5352 12498 5364
rect 78692 5352 78720 5460
rect 80054 5448 80060 5460
rect 80112 5448 80118 5500
rect 80238 5448 80244 5500
rect 80296 5488 80302 5500
rect 190454 5488 190460 5500
rect 80296 5460 190460 5488
rect 80296 5448 80302 5460
rect 190454 5448 190460 5460
rect 190512 5448 190518 5500
rect 83826 5380 83832 5432
rect 83884 5420 83890 5432
rect 195974 5420 195980 5432
rect 83884 5392 195980 5420
rect 83884 5380 83890 5392
rect 195974 5380 195980 5392
rect 196032 5380 196038 5432
rect 12492 5324 78720 5352
rect 12492 5312 12498 5324
rect 87322 5312 87328 5364
rect 87380 5352 87386 5364
rect 202874 5352 202880 5364
rect 87380 5324 202880 5352
rect 87380 5312 87386 5324
rect 202874 5312 202880 5324
rect 202932 5312 202938 5364
rect 52822 5244 52828 5296
rect 52880 5284 52886 5296
rect 60734 5284 60740 5296
rect 52880 5256 60740 5284
rect 52880 5244 52886 5256
rect 60734 5244 60740 5256
rect 60792 5244 60798 5296
rect 78582 5244 78588 5296
rect 78640 5284 78646 5296
rect 93854 5284 93860 5296
rect 78640 5256 93860 5284
rect 78640 5244 78646 5256
rect 93854 5244 93860 5256
rect 93912 5244 93918 5296
rect 109034 5244 109040 5296
rect 109092 5284 109098 5296
rect 219434 5284 219440 5296
rect 109092 5256 219440 5284
rect 109092 5244 109098 5256
rect 219434 5244 219440 5256
rect 219492 5244 219498 5296
rect 22002 5176 22008 5228
rect 22060 5216 22066 5228
rect 95234 5216 95240 5228
rect 22060 5188 95240 5216
rect 22060 5176 22066 5188
rect 95234 5176 95240 5188
rect 95292 5176 95298 5228
rect 98086 5176 98092 5228
rect 98144 5216 98150 5228
rect 105078 5216 105084 5228
rect 98144 5188 105084 5216
rect 98144 5176 98150 5188
rect 105078 5176 105084 5188
rect 105136 5176 105142 5228
rect 105170 5176 105176 5228
rect 105228 5216 105234 5228
rect 231854 5216 231860 5228
rect 105228 5188 231860 5216
rect 105228 5176 105234 5188
rect 231854 5176 231860 5188
rect 231912 5176 231918 5228
rect 26694 5108 26700 5160
rect 26752 5148 26758 5160
rect 81894 5148 81900 5160
rect 26752 5120 81900 5148
rect 26752 5108 26758 5120
rect 81894 5108 81900 5120
rect 81952 5108 81958 5160
rect 82078 5108 82084 5160
rect 82136 5148 82142 5160
rect 103514 5148 103520 5160
rect 82136 5120 103520 5148
rect 82136 5108 82142 5120
rect 103514 5108 103520 5120
rect 103572 5108 103578 5160
rect 103606 5108 103612 5160
rect 103664 5148 103670 5160
rect 103664 5120 109264 5148
rect 103664 5108 103670 5120
rect 30282 5040 30288 5092
rect 30340 5080 30346 5092
rect 81986 5080 81992 5092
rect 30340 5052 81992 5080
rect 30340 5040 30346 5052
rect 81986 5040 81992 5052
rect 82044 5040 82050 5092
rect 82096 5052 86632 5080
rect 33870 4972 33876 5024
rect 33928 5012 33934 5024
rect 82096 5012 82124 5052
rect 33928 4984 82124 5012
rect 86604 5012 86632 5052
rect 86862 5040 86868 5092
rect 86920 5080 86926 5092
rect 109126 5080 109132 5092
rect 86920 5052 109132 5080
rect 86920 5040 86926 5052
rect 109126 5040 109132 5052
rect 109184 5040 109190 5092
rect 109236 5080 109264 5120
rect 127802 5108 127808 5160
rect 127860 5148 127866 5160
rect 127860 5120 137416 5148
rect 127860 5108 127866 5120
rect 124858 5080 124864 5092
rect 109236 5052 124864 5080
rect 124858 5040 124864 5052
rect 124916 5040 124922 5092
rect 130194 5040 130200 5092
rect 130252 5080 130258 5092
rect 137388 5080 137416 5120
rect 137462 5108 137468 5160
rect 137520 5148 137526 5160
rect 266354 5148 266360 5160
rect 137520 5120 266360 5148
rect 137520 5108 137526 5120
rect 266354 5108 266360 5120
rect 266412 5108 266418 5160
rect 269114 5080 269120 5092
rect 130252 5052 137324 5080
rect 137388 5052 269120 5080
rect 130252 5040 130258 5052
rect 114554 5012 114560 5024
rect 86604 4984 114560 5012
rect 33928 4972 33934 4984
rect 114554 4972 114560 4984
rect 114612 4972 114618 5024
rect 119430 4972 119436 5024
rect 119488 5012 119494 5024
rect 134518 5012 134524 5024
rect 119488 4984 134524 5012
rect 119488 4972 119494 4984
rect 134518 4972 134524 4984
rect 134576 4972 134582 5024
rect 134610 4972 134616 5024
rect 134668 5012 134674 5024
rect 137186 5012 137192 5024
rect 134668 4984 137192 5012
rect 134668 4972 134674 4984
rect 137186 4972 137192 4984
rect 137244 4972 137250 5024
rect 137296 5012 137324 5052
rect 269114 5040 269120 5052
rect 269172 5040 269178 5092
rect 271874 5012 271880 5024
rect 137296 4984 271880 5012
rect 271874 4972 271880 4984
rect 271932 4972 271938 5024
rect 37366 4904 37372 4956
rect 37424 4944 37430 4956
rect 81986 4944 81992 4956
rect 37424 4916 81992 4944
rect 37424 4904 37430 4916
rect 81986 4904 81992 4916
rect 82044 4904 82050 4956
rect 86770 4904 86776 4956
rect 86828 4944 86834 4956
rect 120074 4944 120080 4956
rect 86828 4916 120080 4944
rect 86828 4904 86834 4916
rect 120074 4904 120080 4916
rect 120132 4904 120138 4956
rect 128998 4904 129004 4956
rect 129056 4944 129062 4956
rect 270494 4944 270500 4956
rect 129056 4916 270500 4944
rect 129056 4904 129062 4916
rect 270494 4904 270500 4916
rect 270552 4904 270558 4956
rect 40954 4836 40960 4888
rect 41012 4876 41018 4888
rect 78858 4876 78864 4888
rect 41012 4848 78864 4876
rect 41012 4836 41018 4848
rect 78858 4836 78864 4848
rect 78916 4836 78922 4888
rect 86862 4836 86868 4888
rect 86920 4876 86926 4888
rect 126974 4876 126980 4888
rect 86920 4848 126980 4876
rect 86920 4836 86926 4848
rect 126974 4836 126980 4848
rect 127032 4836 127038 4888
rect 127066 4836 127072 4888
rect 127124 4876 127130 4888
rect 137462 4876 137468 4888
rect 127124 4848 137468 4876
rect 127124 4836 127130 4848
rect 137462 4836 137468 4848
rect 137520 4836 137526 4888
rect 137554 4836 137560 4888
rect 137612 4876 137618 4888
rect 276014 4876 276020 4888
rect 137612 4848 276020 4876
rect 137612 4836 137618 4848
rect 276014 4836 276020 4848
rect 276072 4836 276078 4888
rect 44542 4768 44548 4820
rect 44600 4808 44606 4820
rect 132494 4808 132500 4820
rect 44600 4780 132500 4808
rect 44600 4768 44606 4780
rect 132494 4768 132500 4780
rect 132552 4768 132558 4820
rect 132586 4768 132592 4820
rect 132644 4808 132650 4820
rect 134610 4808 134616 4820
rect 132644 4780 134616 4808
rect 132644 4768 132650 4780
rect 134610 4768 134616 4780
rect 134668 4768 134674 4820
rect 134886 4768 134892 4820
rect 134944 4808 134950 4820
rect 278774 4808 278780 4820
rect 134944 4780 278780 4808
rect 134944 4768 134950 4780
rect 278774 4768 278780 4780
rect 278832 4768 278838 4820
rect 67082 4700 67088 4752
rect 67140 4740 67146 4752
rect 67542 4740 67548 4752
rect 67140 4712 67548 4740
rect 67140 4700 67146 4712
rect 67542 4700 67548 4712
rect 67600 4700 67606 4752
rect 76650 4700 76656 4752
rect 76708 4740 76714 4752
rect 184934 4740 184940 4752
rect 76708 4712 184940 4740
rect 76708 4700 76714 4712
rect 184934 4700 184940 4712
rect 184992 4700 184998 4752
rect 73062 4632 73068 4684
rect 73120 4672 73126 4684
rect 179414 4672 179420 4684
rect 73120 4644 179420 4672
rect 73120 4632 73126 4644
rect 179414 4632 179420 4644
rect 179472 4632 179478 4684
rect 69474 4564 69480 4616
rect 69532 4604 69538 4616
rect 172514 4604 172520 4616
rect 69532 4576 172520 4604
rect 69532 4564 69538 4576
rect 172514 4564 172520 4576
rect 172572 4564 172578 4616
rect 65978 4496 65984 4548
rect 66036 4536 66042 4548
rect 166994 4536 167000 4548
rect 66036 4508 167000 4536
rect 66036 4496 66042 4508
rect 166994 4496 167000 4508
rect 167052 4496 167058 4548
rect 62390 4428 62396 4480
rect 62448 4468 62454 4480
rect 161474 4468 161480 4480
rect 62448 4440 161480 4468
rect 62448 4428 62454 4440
rect 161474 4428 161480 4440
rect 161532 4428 161538 4480
rect 58802 4360 58808 4412
rect 58860 4400 58866 4412
rect 155954 4400 155960 4412
rect 58860 4372 155960 4400
rect 58860 4360 58866 4372
rect 155954 4360 155960 4372
rect 156012 4360 156018 4412
rect 55214 4292 55220 4344
rect 55272 4332 55278 4344
rect 150434 4332 150440 4344
rect 55272 4304 150440 4332
rect 55272 4292 55278 4304
rect 150434 4292 150440 4304
rect 150492 4292 150498 4344
rect 51626 4224 51632 4276
rect 51684 4264 51690 4276
rect 143534 4264 143540 4276
rect 51684 4236 143540 4264
rect 51684 4224 51690 4236
rect 143534 4224 143540 4236
rect 143592 4224 143598 4276
rect 48222 4156 48228 4208
rect 48280 4196 48286 4208
rect 138014 4196 138020 4208
rect 48280 4168 138020 4196
rect 48280 4156 48286 4168
rect 138014 4156 138020 4168
rect 138072 4156 138078 4208
rect 8846 4088 8852 4140
rect 8904 4128 8910 4140
rect 71774 4128 71780 4140
rect 8904 4100 71780 4128
rect 8904 4088 8910 4100
rect 71774 4088 71780 4100
rect 71832 4088 71838 4140
rect 71866 4088 71872 4140
rect 71924 4128 71930 4140
rect 72970 4128 72976 4140
rect 71924 4100 72976 4128
rect 71924 4088 71930 4100
rect 72970 4088 72976 4100
rect 73028 4088 73034 4140
rect 73062 4088 73068 4140
rect 73120 4128 73126 4140
rect 74534 4128 74540 4140
rect 73120 4100 74540 4128
rect 73120 4088 73126 4100
rect 74534 4088 74540 4100
rect 74592 4088 74598 4140
rect 81342 4128 81348 4140
rect 75196 4100 81348 4128
rect 13630 4020 13636 4072
rect 13688 4060 13694 4072
rect 75196 4060 75224 4100
rect 81342 4088 81348 4100
rect 81400 4088 81406 4140
rect 81434 4088 81440 4140
rect 81492 4128 81498 4140
rect 82722 4128 82728 4140
rect 81492 4100 82728 4128
rect 81492 4088 81498 4100
rect 82722 4088 82728 4100
rect 82780 4088 82786 4140
rect 82814 4088 82820 4140
rect 82872 4128 82878 4140
rect 86034 4128 86040 4140
rect 82872 4100 86040 4128
rect 82872 4088 82878 4100
rect 86034 4088 86040 4100
rect 86092 4088 86098 4140
rect 186314 4128 186320 4140
rect 89456 4100 186320 4128
rect 13688 4032 75224 4060
rect 13688 4020 13694 4032
rect 79042 4020 79048 4072
rect 79100 4060 79106 4072
rect 79962 4060 79968 4072
rect 79100 4032 79968 4060
rect 79100 4020 79106 4032
rect 79962 4020 79968 4032
rect 80020 4020 80026 4072
rect 80054 4020 80060 4072
rect 80112 4060 80118 4072
rect 89456 4060 89484 4100
rect 186314 4088 186320 4100
rect 186372 4088 186378 4140
rect 80112 4032 89484 4060
rect 80112 4020 80118 4032
rect 89530 4020 89536 4072
rect 89588 4060 89594 4072
rect 194594 4060 194600 4072
rect 89588 4032 194600 4060
rect 89588 4020 89594 4032
rect 194594 4020 194600 4032
rect 194652 4020 194658 4072
rect 14826 3952 14832 4004
rect 14884 3992 14890 4004
rect 84194 3992 84200 4004
rect 14884 3964 84200 3992
rect 14884 3952 14890 3964
rect 84194 3952 84200 3964
rect 84252 3952 84258 4004
rect 84930 3952 84936 4004
rect 84988 3992 84994 4004
rect 89438 3992 89444 4004
rect 84988 3964 89444 3992
rect 84988 3952 84994 3964
rect 89438 3952 89444 3964
rect 89496 3952 89502 4004
rect 89714 3952 89720 4004
rect 89772 3992 89778 4004
rect 93210 3992 93216 4004
rect 89772 3964 93216 3992
rect 89772 3952 89778 3964
rect 93210 3952 93216 3964
rect 93268 3952 93274 4004
rect 198734 3992 198740 4004
rect 93320 3964 198740 3992
rect 18322 3884 18328 3936
rect 18380 3924 18386 3936
rect 89622 3924 89628 3936
rect 18380 3896 89628 3924
rect 18380 3884 18386 3896
rect 89622 3884 89628 3896
rect 89680 3884 89686 3936
rect 89898 3884 89904 3936
rect 89956 3924 89962 3936
rect 93320 3924 93348 3964
rect 198734 3952 198740 3964
rect 198792 3952 198798 4004
rect 89956 3896 93348 3924
rect 89956 3884 89962 3896
rect 93854 3884 93860 3936
rect 93912 3924 93918 3936
rect 205634 3924 205640 3936
rect 93912 3896 205640 3924
rect 93912 3884 93918 3896
rect 205634 3884 205640 3896
rect 205692 3884 205698 3936
rect 95510 3856 95516 3868
rect 27816 3828 95516 3856
rect 23106 3748 23112 3800
rect 23164 3788 23170 3800
rect 27816 3788 27844 3828
rect 95510 3816 95516 3828
rect 95568 3816 95574 3868
rect 95620 3828 96660 3856
rect 23164 3760 27844 3788
rect 23164 3748 23170 3760
rect 27890 3748 27896 3800
rect 27948 3788 27954 3800
rect 95620 3788 95648 3828
rect 27948 3760 95648 3788
rect 27948 3748 27954 3760
rect 95694 3748 95700 3800
rect 95752 3788 95758 3800
rect 96522 3788 96528 3800
rect 95752 3760 96528 3788
rect 95752 3748 95758 3760
rect 96522 3748 96528 3760
rect 96580 3748 96586 3800
rect 96632 3788 96660 3828
rect 96890 3816 96896 3868
rect 96948 3856 96954 3868
rect 96948 3828 102732 3856
rect 96948 3816 96954 3828
rect 102594 3788 102600 3800
rect 96632 3760 102600 3788
rect 102594 3748 102600 3760
rect 102652 3748 102658 3800
rect 102704 3788 102732 3828
rect 102778 3816 102784 3868
rect 102836 3856 102842 3868
rect 103422 3856 103428 3868
rect 102836 3828 103428 3856
rect 102836 3816 102842 3828
rect 103422 3816 103428 3828
rect 103480 3816 103486 3868
rect 103514 3816 103520 3868
rect 103572 3856 103578 3868
rect 104894 3856 104900 3868
rect 103572 3828 104900 3856
rect 103572 3816 103578 3828
rect 104894 3816 104900 3828
rect 104952 3816 104958 3868
rect 108206 3856 108212 3868
rect 106108 3828 108212 3856
rect 105998 3788 106004 3800
rect 102704 3760 106004 3788
rect 105998 3748 106004 3760
rect 106056 3748 106062 3800
rect 31478 3680 31484 3732
rect 31536 3720 31542 3732
rect 106108 3720 106136 3828
rect 108206 3816 108212 3828
rect 108264 3816 108270 3868
rect 218054 3856 218060 3868
rect 108316 3828 218060 3856
rect 106182 3748 106188 3800
rect 106240 3788 106246 3800
rect 108316 3788 108344 3828
rect 218054 3816 218060 3828
rect 218112 3816 218118 3868
rect 113174 3788 113180 3800
rect 106240 3760 108344 3788
rect 108408 3760 113180 3788
rect 106240 3748 106246 3760
rect 31536 3692 106136 3720
rect 31536 3680 31542 3692
rect 106274 3680 106280 3732
rect 106332 3720 106338 3732
rect 108408 3720 108436 3760
rect 113174 3748 113180 3760
rect 113232 3748 113238 3800
rect 113542 3748 113548 3800
rect 113600 3788 113606 3800
rect 114462 3788 114468 3800
rect 113600 3760 114468 3788
rect 113600 3748 113606 3760
rect 114462 3748 114468 3760
rect 114520 3748 114526 3800
rect 114738 3748 114744 3800
rect 114796 3788 114802 3800
rect 115842 3788 115848 3800
rect 114796 3760 115848 3788
rect 114796 3748 114802 3760
rect 115842 3748 115848 3760
rect 115900 3748 115906 3800
rect 116026 3748 116032 3800
rect 116084 3788 116090 3800
rect 238754 3788 238760 3800
rect 116084 3760 238760 3788
rect 116084 3748 116090 3760
rect 238754 3748 238760 3760
rect 238812 3748 238818 3800
rect 106332 3692 108436 3720
rect 106332 3680 106338 3692
rect 108482 3680 108488 3732
rect 108540 3720 108546 3732
rect 110414 3720 110420 3732
rect 108540 3692 110420 3720
rect 108540 3680 108546 3692
rect 110414 3680 110420 3692
rect 110472 3680 110478 3732
rect 111150 3680 111156 3732
rect 111208 3720 111214 3732
rect 241514 3720 241520 3732
rect 111208 3692 241520 3720
rect 111208 3680 111214 3692
rect 241514 3680 241520 3692
rect 241572 3680 241578 3732
rect 36170 3612 36176 3664
rect 36228 3652 36234 3664
rect 36228 3624 113864 3652
rect 36228 3612 36234 3624
rect 32674 3544 32680 3596
rect 32732 3584 32738 3596
rect 106274 3584 106280 3596
rect 32732 3556 106280 3584
rect 32732 3544 32738 3556
rect 106274 3544 106280 3556
rect 106332 3544 106338 3596
rect 106366 3544 106372 3596
rect 106424 3584 106430 3596
rect 107562 3584 107568 3596
rect 106424 3556 107568 3584
rect 106424 3544 106430 3556
rect 107562 3544 107568 3556
rect 107620 3544 107626 3596
rect 109954 3544 109960 3596
rect 110012 3584 110018 3596
rect 113726 3584 113732 3596
rect 110012 3556 113732 3584
rect 110012 3544 110018 3556
rect 113726 3544 113732 3556
rect 113784 3544 113790 3596
rect 1670 3476 1676 3528
rect 1728 3516 1734 3528
rect 2682 3516 2688 3528
rect 1728 3488 2688 3516
rect 1728 3476 1734 3488
rect 2682 3476 2688 3488
rect 2740 3476 2746 3528
rect 2866 3476 2872 3528
rect 2924 3516 2930 3528
rect 4062 3516 4068 3528
rect 2924 3488 4068 3516
rect 2924 3476 2930 3488
rect 4062 3476 4068 3488
rect 4120 3476 4126 3528
rect 7650 3476 7656 3528
rect 7708 3516 7714 3528
rect 8202 3516 8208 3528
rect 7708 3488 8208 3516
rect 7708 3476 7714 3488
rect 8202 3476 8208 3488
rect 8260 3476 8266 3528
rect 10042 3476 10048 3528
rect 10100 3516 10106 3528
rect 10962 3516 10968 3528
rect 10100 3488 10968 3516
rect 10100 3476 10106 3488
rect 10962 3476 10968 3488
rect 11020 3476 11026 3528
rect 16022 3476 16028 3528
rect 16080 3516 16086 3528
rect 16482 3516 16488 3528
rect 16080 3488 16488 3516
rect 16080 3476 16086 3488
rect 16482 3476 16488 3488
rect 16540 3476 16546 3528
rect 19518 3476 19524 3528
rect 19576 3516 19582 3528
rect 20622 3516 20628 3528
rect 19576 3488 20628 3516
rect 19576 3476 19582 3488
rect 20622 3476 20628 3488
rect 20680 3476 20686 3528
rect 20714 3476 20720 3528
rect 20772 3516 20778 3528
rect 21910 3516 21916 3528
rect 20772 3488 21916 3516
rect 20772 3476 20778 3488
rect 21910 3476 21916 3488
rect 21968 3476 21974 3528
rect 24302 3476 24308 3528
rect 24360 3516 24366 3528
rect 24762 3516 24768 3528
rect 24360 3488 24768 3516
rect 24360 3476 24366 3488
rect 24762 3476 24768 3488
rect 24820 3476 24826 3528
rect 25498 3476 25504 3528
rect 25556 3516 25562 3528
rect 26142 3516 26148 3528
rect 25556 3488 26148 3516
rect 25556 3476 25562 3488
rect 26142 3476 26148 3488
rect 26200 3476 26206 3528
rect 34974 3476 34980 3528
rect 35032 3516 35038 3528
rect 113634 3516 113640 3528
rect 35032 3488 113640 3516
rect 35032 3476 35038 3488
rect 113634 3476 113640 3488
rect 113692 3476 113698 3528
rect 113836 3516 113864 3624
rect 114002 3612 114008 3664
rect 114060 3652 114066 3664
rect 114060 3624 116164 3652
rect 114060 3612 114066 3624
rect 114094 3544 114100 3596
rect 114152 3584 114158 3596
rect 116026 3584 116032 3596
rect 114152 3556 116032 3584
rect 114152 3544 114158 3556
rect 116026 3544 116032 3556
rect 116084 3544 116090 3596
rect 116136 3584 116164 3624
rect 117130 3612 117136 3664
rect 117188 3652 117194 3664
rect 117188 3624 120580 3652
rect 117188 3612 117194 3624
rect 117314 3584 117320 3596
rect 116136 3556 117320 3584
rect 117314 3544 117320 3556
rect 117372 3544 117378 3596
rect 118234 3544 118240 3596
rect 118292 3584 118298 3596
rect 120552 3584 120580 3624
rect 120626 3612 120632 3664
rect 120684 3652 120690 3664
rect 121362 3652 121368 3664
rect 120684 3624 121368 3652
rect 120684 3612 120690 3624
rect 121362 3612 121368 3624
rect 121420 3612 121426 3664
rect 121822 3612 121828 3664
rect 121880 3652 121886 3664
rect 122742 3652 122748 3664
rect 121880 3624 122748 3652
rect 121880 3612 121886 3624
rect 122742 3612 122748 3624
rect 122800 3612 122806 3664
rect 122834 3612 122840 3664
rect 122892 3652 122898 3664
rect 252554 3652 252560 3664
rect 122892 3624 252560 3652
rect 122892 3612 122898 3624
rect 252554 3612 252560 3624
rect 252612 3612 252618 3664
rect 251174 3584 251180 3596
rect 118292 3556 120488 3584
rect 120552 3556 122788 3584
rect 118292 3544 118298 3556
rect 118694 3516 118700 3528
rect 113836 3488 118700 3516
rect 118694 3476 118700 3488
rect 118752 3476 118758 3528
rect 120460 3516 120488 3556
rect 122650 3516 122656 3528
rect 120460 3488 122656 3516
rect 122650 3476 122656 3488
rect 122708 3476 122714 3528
rect 122760 3516 122788 3556
rect 123036 3556 251180 3584
rect 123036 3516 123064 3556
rect 251174 3544 251180 3556
rect 251232 3544 251238 3596
rect 122760 3488 123064 3516
rect 124214 3476 124220 3528
rect 124272 3516 124278 3528
rect 262214 3516 262220 3528
rect 124272 3488 262220 3516
rect 124272 3476 124278 3488
rect 262214 3476 262220 3488
rect 262272 3476 262278 3528
rect 11238 3408 11244 3460
rect 11296 3448 11302 3460
rect 32398 3448 32404 3460
rect 11296 3420 32404 3448
rect 11296 3408 11302 3420
rect 32398 3408 32404 3420
rect 32456 3408 32462 3460
rect 42150 3408 42156 3460
rect 42208 3448 42214 3460
rect 42702 3448 42708 3460
rect 42208 3420 42708 3448
rect 42208 3408 42214 3420
rect 42702 3408 42708 3420
rect 42760 3408 42766 3460
rect 42794 3408 42800 3460
rect 42852 3448 42858 3460
rect 122926 3448 122932 3460
rect 42852 3420 122932 3448
rect 42852 3408 42858 3420
rect 122926 3408 122932 3420
rect 122984 3408 122990 3460
rect 125410 3408 125416 3460
rect 125468 3448 125474 3460
rect 264974 3448 264980 3460
rect 125468 3420 264980 3448
rect 125468 3408 125474 3420
rect 264974 3408 264980 3420
rect 265032 3408 265038 3460
rect 6454 3340 6460 3392
rect 6512 3380 6518 3392
rect 6512 3352 61148 3380
rect 6512 3340 6518 3352
rect 4062 3272 4068 3324
rect 4120 3312 4126 3324
rect 61010 3312 61016 3324
rect 4120 3284 61016 3312
rect 4120 3272 4126 3284
rect 61010 3272 61016 3284
rect 61068 3272 61074 3324
rect 61120 3312 61148 3352
rect 61194 3340 61200 3392
rect 61252 3380 61258 3392
rect 62022 3380 62028 3392
rect 61252 3352 62028 3380
rect 61252 3340 61258 3352
rect 62022 3340 62028 3352
rect 62080 3340 62086 3392
rect 62114 3340 62120 3392
rect 62172 3380 62178 3392
rect 66346 3380 66352 3392
rect 62172 3352 66352 3380
rect 62172 3340 62178 3352
rect 66346 3340 66352 3352
rect 66404 3340 66410 3392
rect 68278 3340 68284 3392
rect 68336 3380 68342 3392
rect 68336 3352 75224 3380
rect 68336 3340 68342 3352
rect 70394 3312 70400 3324
rect 61120 3284 70400 3312
rect 70394 3272 70400 3284
rect 70452 3272 70458 3324
rect 70670 3272 70676 3324
rect 70728 3312 70734 3324
rect 75086 3312 75092 3324
rect 70728 3284 75092 3312
rect 70728 3272 70734 3284
rect 75086 3272 75092 3284
rect 75144 3272 75150 3324
rect 75196 3312 75224 3352
rect 75270 3340 75276 3392
rect 75328 3380 75334 3392
rect 175274 3380 175280 3392
rect 75328 3352 175280 3380
rect 75328 3340 75334 3352
rect 175274 3340 175280 3352
rect 175332 3340 175338 3392
rect 171134 3312 171140 3324
rect 75196 3284 171140 3312
rect 171134 3272 171140 3284
rect 171192 3272 171198 3324
rect 566 3204 572 3256
rect 624 3244 630 3256
rect 61378 3244 61384 3256
rect 624 3216 61384 3244
rect 624 3204 630 3216
rect 61378 3204 61384 3216
rect 61436 3204 61442 3256
rect 63586 3204 63592 3256
rect 63644 3244 63650 3256
rect 162854 3244 162860 3256
rect 63644 3216 162860 3244
rect 63644 3204 63650 3216
rect 162854 3204 162860 3216
rect 162912 3204 162918 3256
rect 5258 3136 5264 3188
rect 5316 3176 5322 3188
rect 5316 3148 37780 3176
rect 5316 3136 5322 3148
rect 17218 3068 17224 3120
rect 17276 3108 17282 3120
rect 37752 3108 37780 3148
rect 38562 3136 38568 3188
rect 38620 3176 38626 3188
rect 42794 3176 42800 3188
rect 38620 3148 42800 3176
rect 38620 3136 38626 3148
rect 42794 3136 42800 3148
rect 42852 3136 42858 3188
rect 46934 3136 46940 3188
rect 46992 3176 46998 3188
rect 48130 3176 48136 3188
rect 46992 3148 48136 3176
rect 46992 3136 46998 3148
rect 48130 3136 48136 3148
rect 48188 3136 48194 3188
rect 50522 3136 50528 3188
rect 50580 3176 50586 3188
rect 50982 3176 50988 3188
rect 50580 3148 50988 3176
rect 50580 3136 50586 3148
rect 50982 3136 50988 3148
rect 51040 3136 51046 3188
rect 56410 3136 56416 3188
rect 56468 3176 56474 3188
rect 151814 3176 151820 3188
rect 56468 3148 151820 3176
rect 56468 3136 56474 3148
rect 151814 3136 151820 3148
rect 151872 3136 151878 3188
rect 39298 3108 39304 3120
rect 17276 3080 37596 3108
rect 37752 3080 39304 3108
rect 17276 3068 17282 3080
rect 29086 3000 29092 3052
rect 29144 3040 29150 3052
rect 29144 3012 37504 3040
rect 29144 3000 29150 3012
rect 37476 2904 37504 3012
rect 37568 2972 37596 3080
rect 39298 3068 39304 3080
rect 39356 3068 39362 3120
rect 50430 3108 50436 3120
rect 47964 3080 50436 3108
rect 47964 2972 47992 3080
rect 50430 3068 50436 3080
rect 50488 3068 50494 3120
rect 57606 3068 57612 3120
rect 57664 3108 57670 3120
rect 153194 3108 153200 3120
rect 57664 3080 153200 3108
rect 57664 3068 57670 3080
rect 153194 3068 153200 3080
rect 153252 3068 153258 3120
rect 54018 3000 54024 3052
rect 54076 3040 54082 3052
rect 147674 3040 147680 3052
rect 54076 3012 147680 3040
rect 54076 3000 54082 3012
rect 147674 3000 147680 3012
rect 147732 3000 147738 3052
rect 37568 2944 47992 2972
rect 49326 2932 49332 2984
rect 49384 2972 49390 2984
rect 139394 2972 139400 2984
rect 49384 2944 139400 2972
rect 49384 2932 49390 2944
rect 139394 2932 139400 2944
rect 139452 2932 139458 2984
rect 42058 2904 42064 2916
rect 37476 2876 42064 2904
rect 42058 2864 42064 2876
rect 42116 2864 42122 2916
rect 45738 2864 45744 2916
rect 45796 2904 45802 2916
rect 133966 2904 133972 2916
rect 45796 2876 133972 2904
rect 45796 2864 45802 2876
rect 133966 2864 133972 2876
rect 134024 2864 134030 2916
rect 43346 2796 43352 2848
rect 43404 2836 43410 2848
rect 129826 2836 129832 2848
rect 43404 2808 124168 2836
rect 43404 2796 43410 2808
rect 124140 2768 124168 2808
rect 127820 2808 129832 2836
rect 127820 2768 127848 2808
rect 129826 2796 129832 2808
rect 129884 2796 129890 2848
rect 124140 2740 127848 2768
rect 88518 1096 88524 1148
rect 88576 1136 88582 1148
rect 89346 1136 89352 1148
rect 88576 1108 89352 1136
rect 88576 1096 88582 1108
rect 89346 1096 89352 1108
rect 89404 1096 89410 1148
rect 67082 552 67088 604
rect 67140 592 67146 604
rect 67174 592 67180 604
rect 67140 564 67180 592
rect 67140 552 67146 564
rect 67174 552 67180 564
rect 67232 552 67238 604
<< via1 >>
rect 58624 700952 58676 701004
rect 137836 700952 137888 701004
rect 137928 700952 137980 701004
rect 235172 700952 235224 701004
rect 58716 700884 58768 700936
rect 202788 700884 202840 700936
rect 57796 700816 57848 700868
rect 218980 700816 219032 700868
rect 58900 700748 58952 700800
rect 267648 700748 267700 700800
rect 58808 700680 58860 700732
rect 283840 700680 283892 700732
rect 58992 700612 59044 700664
rect 332508 700612 332560 700664
rect 57888 700544 57940 700596
rect 348792 700544 348844 700596
rect 59176 700476 59228 700528
rect 397460 700476 397512 700528
rect 59084 700408 59136 700460
rect 413652 700408 413704 700460
rect 59268 700340 59320 700392
rect 478512 700340 478564 700392
rect 59360 700272 59412 700324
rect 527180 700272 527232 700324
rect 58532 700204 58584 700256
rect 154120 700204 154172 700256
rect 58348 700136 58400 700188
rect 89168 700136 89220 700188
rect 58440 700068 58492 700120
rect 72976 700068 73028 700120
rect 40500 699932 40552 699984
rect 42064 699932 42116 699984
rect 8116 699660 8168 699712
rect 10324 699660 10376 699712
rect 24308 699660 24360 699712
rect 24768 699660 24820 699712
rect 137284 699660 137336 699712
rect 137928 699660 137980 699712
rect 104992 698232 105044 698284
rect 105544 698232 105596 698284
rect 364432 698232 364484 698284
rect 365076 698232 365128 698284
rect 560300 697280 560352 697332
rect 565176 697280 565228 697332
rect 540980 697144 541032 697196
rect 548616 697144 548668 697196
rect 70308 697076 70360 697128
rect 77208 697076 77260 697128
rect 89628 697076 89680 697128
rect 96528 697076 96580 697128
rect 108948 697076 109000 697128
rect 115848 697076 115900 697128
rect 128268 697076 128320 697128
rect 135168 697076 135220 697128
rect 147588 697076 147640 697128
rect 154488 697076 154540 697128
rect 166908 697076 166960 697128
rect 173808 697076 173860 697128
rect 186228 697076 186280 697128
rect 193128 697076 193180 697128
rect 205548 697076 205600 697128
rect 212448 697076 212500 697128
rect 224868 697076 224920 697128
rect 231768 697076 231820 697128
rect 244188 697076 244240 697128
rect 251088 697076 251140 697128
rect 263508 697076 263560 697128
rect 270408 697076 270460 697128
rect 282828 697076 282880 697128
rect 289728 697076 289780 697128
rect 302148 697076 302200 697128
rect 309048 697076 309100 697128
rect 321468 697076 321520 697128
rect 328368 697076 328420 697128
rect 170128 695444 170180 695496
rect 170312 695444 170364 695496
rect 429200 692792 429252 692844
rect 429936 692792 429988 692844
rect 494060 692792 494112 692844
rect 494888 692792 494940 692844
rect 173900 686264 173952 686316
rect 178776 686264 178828 686316
rect 367100 686264 367152 686316
rect 371976 686264 372028 686316
rect 560300 686264 560352 686316
rect 565176 686264 565228 686316
rect 154580 686128 154632 686180
rect 162216 686128 162268 686180
rect 289820 686128 289872 686180
rect 294512 686128 294564 686180
rect 347780 686128 347832 686180
rect 355416 686128 355468 686180
rect 540980 686128 541032 686180
rect 548616 686128 548668 686180
rect 169852 685924 169904 685976
rect 170128 685924 170180 685976
rect 299572 685856 299624 685908
rect 300124 685856 300176 685908
rect 559012 684496 559064 684548
rect 559656 684496 559708 684548
rect 169852 684428 169904 684480
rect 170220 684428 170272 684480
rect 299572 684428 299624 684480
rect 299664 684428 299716 684480
rect 299664 678988 299716 679040
rect 299664 678852 299716 678904
rect 559012 674840 559064 674892
rect 559380 674840 559432 674892
rect 173900 673888 173952 673940
rect 178776 673888 178828 673940
rect 367100 673888 367152 673940
rect 371976 673888 372028 673940
rect 560300 673888 560352 673940
rect 565176 673888 565228 673940
rect 154580 673752 154632 673804
rect 162216 673752 162268 673804
rect 289820 673752 289872 673804
rect 292672 673752 292724 673804
rect 347780 673752 347832 673804
rect 355416 673752 355468 673804
rect 540980 673752 541032 673804
rect 548616 673752 548668 673804
rect 104900 673480 104952 673532
rect 105084 673480 105136 673532
rect 494060 673480 494112 673532
rect 494244 673480 494296 673532
rect 429200 673412 429252 673464
rect 429476 673412 429528 673464
rect 364432 669400 364484 669452
rect 364432 669264 364484 669316
rect 494060 669264 494112 669316
rect 494244 669264 494296 669316
rect 3516 667904 3568 667956
rect 21364 667904 21416 667956
rect 299664 666544 299716 666596
rect 299940 666544 299992 666596
rect 493968 666476 494020 666528
rect 494244 666476 494296 666528
rect 169944 661716 169996 661768
rect 170220 661716 170272 661768
rect 559104 661716 559156 661768
rect 559380 661716 559432 661768
rect 169944 656888 169996 656940
rect 170036 656888 170088 656940
rect 493968 656888 494020 656940
rect 494152 656888 494204 656940
rect 559104 656888 559156 656940
rect 559196 656888 559248 656940
rect 299480 656820 299532 656872
rect 299756 656820 299808 656872
rect 263508 653352 263560 653404
rect 378140 653352 378192 653404
rect 3056 652740 3108 652792
rect 13084 652740 13136 652792
rect 129280 652740 129332 652792
rect 133696 652740 133748 652792
rect 139400 652808 139452 652860
rect 378140 652808 378192 652860
rect 383476 652808 383528 652860
rect 387800 652808 387852 652860
rect 258632 652740 258684 652792
rect 263508 652740 263560 652792
rect 197360 650904 197412 650956
rect 206928 650904 206980 650956
rect 195244 650768 195296 650820
rect 197360 650768 197412 650820
rect 367100 650768 367152 650820
rect 370412 650768 370464 650820
rect 57704 650700 57756 650752
rect 105084 650700 105136 650752
rect 278780 650700 278832 650752
rect 288348 650700 288400 650752
rect 572628 650700 572680 650752
rect 579528 650700 579580 650752
rect 59452 650632 59504 650684
rect 364524 650632 364576 650684
rect 89628 650564 89680 650616
rect 96528 650564 96580 650616
rect 106740 650564 106792 650616
rect 115756 650564 115808 650616
rect 207020 650564 207072 650616
rect 115940 650496 115992 650548
rect 120724 650496 120776 650548
rect 137652 650428 137704 650480
rect 147588 650428 147640 650480
rect 147680 650360 147732 650412
rect 157248 650360 157300 650412
rect 157340 650360 157392 650412
rect 164148 650292 164200 650344
rect 164240 650292 164292 650344
rect 195244 650360 195296 650412
rect 237380 650496 237432 650548
rect 237564 650360 237616 650412
rect 340788 650564 340840 650616
rect 347688 650564 347740 650616
rect 560300 650564 560352 650616
rect 563152 650564 563204 650616
rect 289820 650496 289872 650548
rect 292672 650496 292724 650548
rect 405740 650496 405792 650548
rect 413376 650496 413428 650548
rect 533988 650496 534040 650548
rect 540888 650496 540940 650548
rect 266360 650428 266412 650480
rect 456708 650428 456760 650480
rect 463608 650428 463660 650480
rect 476028 650428 476080 650480
rect 482928 650428 482980 650480
rect 495348 650428 495400 650480
rect 502248 650428 502300 650480
rect 514668 650428 514720 650480
rect 521568 650428 521620 650480
rect 285588 650292 285640 650344
rect 386420 650292 386472 650344
rect 280068 650088 280120 650140
rect 285588 650156 285640 650208
rect 266360 650020 266412 650072
rect 270500 650020 270552 650072
rect 169944 647232 169996 647284
rect 170036 647232 170088 647284
rect 299480 647232 299532 647284
rect 299664 647232 299716 647284
rect 429384 647232 429436 647284
rect 429476 647232 429528 647284
rect 559104 647232 559156 647284
rect 559196 647232 559248 647284
rect 297364 645872 297416 645924
rect 307116 645872 307168 645924
rect 294604 644444 294656 644496
rect 307116 644444 307168 644496
rect 291844 643084 291896 643136
rect 307116 643084 307168 643136
rect 290464 641724 290516 641776
rect 307668 641724 307720 641776
rect 169944 640364 169996 640416
rect 170036 640364 170088 640416
rect 429384 640364 429436 640416
rect 429476 640364 429528 640416
rect 559104 640364 559156 640416
rect 559196 640364 559248 640416
rect 287704 640296 287756 640348
rect 307668 640296 307720 640348
rect 286324 638936 286376 638988
rect 306656 638936 306708 638988
rect 301504 637576 301556 637628
rect 306840 637576 306892 637628
rect 494060 634788 494112 634840
rect 494244 634788 494296 634840
rect 299664 630708 299716 630760
rect 299756 630708 299808 630760
rect 169852 630640 169904 630692
rect 170036 630640 170088 630692
rect 429292 630640 429344 630692
rect 429476 630640 429528 630692
rect 559012 630640 559064 630692
rect 559196 630640 559248 630692
rect 494060 615476 494112 615528
rect 494244 615476 494296 615528
rect 169852 611328 169904 611380
rect 170036 611328 170088 611380
rect 299572 611328 299624 611380
rect 299756 611328 299808 611380
rect 429292 611328 429344 611380
rect 429476 611328 429528 611380
rect 559012 611328 559064 611380
rect 559196 611328 559248 611380
rect 3608 609968 3660 610020
rect 31024 609968 31076 610020
rect 169852 608540 169904 608592
rect 169944 608540 169996 608592
rect 299572 608540 299624 608592
rect 299664 608540 299716 608592
rect 429292 608540 429344 608592
rect 429384 608540 429436 608592
rect 559012 608540 559064 608592
rect 559104 608540 559156 608592
rect 169852 601672 169904 601724
rect 170128 601672 170180 601724
rect 299572 601672 299624 601724
rect 299848 601672 299900 601724
rect 429292 601672 429344 601724
rect 429568 601672 429620 601724
rect 559012 601672 559064 601724
rect 559288 601672 559340 601724
rect 169944 598884 169996 598936
rect 170128 598884 170180 598936
rect 299664 598884 299716 598936
rect 299848 598884 299900 598936
rect 559104 598884 559156 598936
rect 559288 598884 559340 598936
rect 494060 596164 494112 596216
rect 494244 596164 494296 596216
rect 3332 594804 3384 594856
rect 14464 594804 14516 594856
rect 429568 592016 429620 592068
rect 429660 591880 429712 591932
rect 169944 589296 169996 589348
rect 170220 589296 170272 589348
rect 270408 589296 270460 589348
rect 309784 589296 309836 589348
rect 559104 589296 559156 589348
rect 559380 589296 559432 589348
rect 493876 589228 493928 589280
rect 494152 589228 494204 589280
rect 429292 583040 429344 583092
rect 429568 583040 429620 583092
rect 170220 582428 170272 582480
rect 299940 582428 299992 582480
rect 559380 582428 559432 582480
rect 170128 582292 170180 582344
rect 299848 582292 299900 582344
rect 559288 582292 559340 582344
rect 493876 579640 493928 579692
rect 494060 579640 494112 579692
rect 429292 578212 429344 578264
rect 429384 578212 429436 578264
rect 429384 572568 429436 572620
rect 429660 572568 429712 572620
rect 494152 569848 494204 569900
rect 494336 569848 494388 569900
rect 494336 563184 494388 563236
rect 494336 563048 494388 563100
rect 56876 560872 56928 560924
rect 188988 560872 189040 560924
rect 305644 560872 305696 560924
rect 429476 560260 429528 560312
rect 429660 560260 429712 560312
rect 559012 560260 559064 560312
rect 559104 560260 559156 560312
rect 309784 560192 309836 560244
rect 310428 560192 310480 560244
rect 389180 560192 389232 560244
rect 62028 558832 62080 558884
rect 197360 558832 197412 558884
rect 215300 558832 215352 558884
rect 224500 558832 224552 558884
rect 335452 558832 335504 558884
rect 344836 558832 344888 558884
rect 67456 558764 67508 558816
rect 201500 558764 201552 558816
rect 328460 558764 328512 558816
rect 338028 558764 338080 558816
rect 77392 558696 77444 558748
rect 86408 558696 86460 558748
rect 95792 558696 95844 558748
rect 105544 558696 105596 558748
rect 125508 558696 125560 558748
rect 208400 558696 208452 558748
rect 209688 558696 209740 558748
rect 223580 558696 223632 558748
rect 231860 558696 231912 558748
rect 328552 558696 328604 558748
rect 337936 558696 337988 558748
rect 76012 558628 76064 558680
rect 84292 558628 84344 558680
rect 93308 558628 93360 558680
rect 97816 558628 97868 558680
rect 133144 558628 133196 558680
rect 224500 558628 224552 558680
rect 233240 558628 233292 558680
rect 344836 558628 344888 558680
rect 353300 558628 353352 558680
rect 85212 558560 85264 558612
rect 94872 558560 94924 558612
rect 103888 558560 103940 558612
rect 104164 558560 104216 558612
rect 104808 558560 104860 558612
rect 137376 558560 137428 558612
rect 217784 558560 217836 558612
rect 225880 558560 225932 558612
rect 234896 558560 234948 558612
rect 336464 558560 336516 558612
rect 345756 558560 345808 558612
rect 354680 558560 354732 558612
rect 79600 558492 79652 558544
rect 88892 558492 88944 558544
rect 98092 558492 98144 558544
rect 99564 558492 99616 558544
rect 108304 558492 108356 558544
rect 209688 558492 209740 558544
rect 217968 558492 218020 558544
rect 78496 558424 78548 558476
rect 87880 558424 87932 558476
rect 96988 558424 97040 558476
rect 106924 558424 106976 558476
rect 108488 558424 108540 558476
rect 144184 558424 144236 558476
rect 213920 558424 213972 558476
rect 223580 558492 223632 558544
rect 330484 558492 330536 558544
rect 339868 558492 339920 558544
rect 349528 558492 349580 558544
rect 357716 558492 357768 558544
rect 80796 558356 80848 558408
rect 89812 558356 89864 558408
rect 99564 558356 99616 558408
rect 72608 558288 72660 558340
rect 81900 558288 81952 558340
rect 91100 558288 91152 558340
rect 92480 558288 92532 558340
rect 98000 558288 98052 558340
rect 98092 558288 98144 558340
rect 100576 558356 100628 558408
rect 101956 558356 102008 558408
rect 140044 558356 140096 558408
rect 208584 558356 208636 558408
rect 210608 558356 210660 558408
rect 100392 558288 100444 558340
rect 140136 558288 140188 558340
rect 211160 558288 211212 558340
rect 211804 558288 211856 558340
rect 215116 558288 215168 558340
rect 217968 558356 218020 558408
rect 227168 558424 227220 558476
rect 231860 558424 231912 558476
rect 337752 558424 337804 558476
rect 346860 558424 346912 558476
rect 356060 558424 356112 558476
rect 220084 558288 220136 558340
rect 220820 558288 220872 558340
rect 221096 558288 221148 558340
rect 229560 558356 229612 558408
rect 238760 558356 238812 558408
rect 329288 558356 329340 558408
rect 339040 558356 339092 558408
rect 348240 558356 348292 558408
rect 357440 558356 357492 558408
rect 221556 558288 221608 558340
rect 230480 558288 230532 558340
rect 332692 558288 332744 558340
rect 342536 558288 342588 558340
rect 348148 558288 348200 558340
rect 81256 558220 81308 558272
rect 145564 558220 145616 558272
rect 76840 558152 76892 558204
rect 141424 558152 141476 558204
rect 206928 558152 206980 558204
rect 215300 558152 215352 558204
rect 222384 558220 222436 558272
rect 231860 558220 231912 558272
rect 331312 558220 331364 558272
rect 331772 558220 331824 558272
rect 341248 558220 341300 558272
rect 350540 558220 350592 558272
rect 73804 558084 73856 558136
rect 82820 558084 82872 558136
rect 83832 558084 83884 558136
rect 152464 558084 152516 558136
rect 79416 558016 79468 558068
rect 148324 558016 148376 558068
rect 200120 558016 200172 558068
rect 213644 558016 213696 558068
rect 74264 557948 74316 558000
rect 135904 557948 135956 558000
rect 194416 557948 194468 558000
rect 200028 557948 200080 558000
rect 203524 557948 203576 558000
rect 213092 557948 213144 558000
rect 218980 558016 219032 558068
rect 228180 558152 228232 558204
rect 237380 558152 237432 558204
rect 288532 558152 288584 558204
rect 298008 558152 298060 558204
rect 302240 558152 302292 558204
rect 313372 558152 313424 558204
rect 334072 558152 334124 558204
rect 343640 558152 343692 558204
rect 351920 558152 351972 558204
rect 283748 558084 283800 558136
rect 354680 558084 354732 558136
rect 298008 557948 298060 558000
rect 302148 557948 302200 558000
rect 326344 557948 326396 558000
rect 335452 557948 335504 558000
rect 82820 557880 82872 557932
rect 92480 557880 92532 557932
rect 93768 557880 93820 557932
rect 127256 557880 127308 557932
rect 129648 557880 129700 557932
rect 208584 557880 208636 557932
rect 302884 557880 302936 557932
rect 317420 557880 317472 557932
rect 323584 557880 323636 557932
rect 332692 557880 332744 557932
rect 79968 557812 80020 557864
rect 102876 557812 102928 557864
rect 121368 557812 121420 557864
rect 206100 557812 206152 557864
rect 206928 557812 206980 557864
rect 209044 557812 209096 557864
rect 218980 557812 219032 557864
rect 288440 557812 288492 557864
rect 297456 557812 297508 557864
rect 320180 557812 320232 557864
rect 322204 557812 322256 557864
rect 331312 557812 331364 557864
rect 66168 557744 66220 557796
rect 200212 557744 200264 557796
rect 202144 557744 202196 557796
rect 211160 557744 211212 557796
rect 213644 557744 213696 557796
rect 222108 557744 222160 557796
rect 222200 557744 222252 557796
rect 229100 557744 229152 557796
rect 288348 557744 288400 557796
rect 302148 557744 302200 557796
rect 302240 557744 302292 557796
rect 324964 557744 325016 557796
rect 334072 557744 334124 557796
rect 75000 557676 75052 557728
rect 84200 557676 84252 557728
rect 93308 557676 93360 557728
rect 99840 557676 99892 557728
rect 107476 557676 107528 557728
rect 141516 557676 141568 557728
rect 204904 557676 204956 557728
rect 213920 557676 213972 557728
rect 63408 557608 63460 557660
rect 198740 557608 198792 557660
rect 207664 557608 207716 557660
rect 217784 557608 217836 557660
rect 238668 557608 238720 557660
rect 91100 557540 91152 557592
rect 100024 557540 100076 557592
rect 99840 557472 99892 557524
rect 102784 557540 102836 557592
rect 100576 557472 100628 557524
rect 107752 557540 107804 557592
rect 108488 557540 108540 557592
rect 127256 557540 127308 557592
rect 131764 557540 131816 557592
rect 200028 557540 200080 557592
rect 200120 557540 200172 557592
rect 241612 557676 241664 557728
rect 283656 557676 283708 557728
rect 351920 557676 351972 557728
rect 251088 557608 251140 557660
rect 253848 557608 253900 557660
rect 253940 557608 253992 557660
rect 270408 557608 270460 557660
rect 273168 557608 273220 557660
rect 273260 557608 273312 557660
rect 260840 557540 260892 557592
rect 283564 557608 283616 557660
rect 353300 557608 353352 557660
rect 282368 557540 282420 557592
rect 288348 557540 288400 557592
rect 327724 557540 327776 557592
rect 336464 557540 336516 557592
rect 58256 556180 58308 556232
rect 580172 556180 580224 556232
rect 282368 549244 282420 549296
rect 282460 549244 282512 549296
rect 77576 545708 77628 545760
rect 188804 545708 188856 545760
rect 560300 545504 560352 545556
rect 563152 545504 563204 545556
rect 302148 545436 302200 545488
rect 309048 545436 309100 545488
rect 572628 545436 572680 545488
rect 579528 545436 579580 545488
rect 115940 545368 115992 545420
rect 125416 545368 125468 545420
rect 135260 545368 135312 545420
rect 144828 545368 144880 545420
rect 195888 545368 195940 545420
rect 201408 545368 201460 545420
rect 212540 545368 212592 545420
rect 222016 545368 222068 545420
rect 231860 545368 231912 545420
rect 241428 545368 241480 545420
rect 251180 545368 251232 545420
rect 260748 545368 260800 545420
rect 483020 545368 483072 545420
rect 485872 545368 485924 545420
rect 540980 545368 541032 545420
rect 548616 545368 548668 545420
rect 85580 545300 85632 545352
rect 95056 545300 95108 545352
rect 166908 545300 166960 545352
rect 177304 545300 177356 545352
rect 321468 545300 321520 545352
rect 328368 545300 328420 545352
rect 96620 545232 96672 545284
rect 104808 545232 104860 545284
rect 57612 545028 57664 545080
rect 112812 545028 112864 545080
rect 114928 545028 114980 545080
rect 202144 545028 202196 545080
rect 89628 544960 89680 545012
rect 177212 544960 177264 545012
rect 92388 544892 92440 544944
rect 181352 544892 181404 544944
rect 96252 544824 96304 544876
rect 188344 544824 188396 544876
rect 91008 544756 91060 544808
rect 179236 544756 179288 544808
rect 96528 544688 96580 544740
rect 189632 544688 189684 544740
rect 94136 544620 94188 544672
rect 188436 544620 188488 544672
rect 89996 544552 90048 544604
rect 188620 544552 188672 544604
rect 57060 544484 57112 544536
rect 102508 544484 102560 544536
rect 103428 544484 103480 544536
rect 202052 544484 202104 544536
rect 57428 544416 57480 544468
rect 108672 544416 108724 544468
rect 110328 544416 110380 544468
rect 212172 544416 212224 544468
rect 81716 544348 81768 544400
rect 195980 544348 196032 544400
rect 86868 544280 86920 544332
rect 173072 544280 173124 544332
rect 88248 544212 88300 544264
rect 175096 544212 175148 544264
rect 86776 544144 86828 544196
rect 170956 544144 171008 544196
rect 85488 544076 85540 544128
rect 168840 544076 168892 544128
rect 73068 544008 73120 544060
rect 148140 544008 148192 544060
rect 102876 543940 102928 543992
rect 160560 543940 160612 543992
rect 57520 543872 57572 543924
rect 110788 543872 110840 543924
rect 57336 543804 57388 543856
rect 106648 543804 106700 543856
rect 57244 543736 57296 543788
rect 104532 543736 104584 543788
rect 429384 543736 429436 543788
rect 71688 543668 71740 543720
rect 75460 543668 75512 543720
rect 75828 543668 75880 543720
rect 152280 543668 152332 543720
rect 152464 543668 152516 543720
rect 166816 543668 166868 543720
rect 206928 543668 206980 543720
rect 220452 543668 220504 543720
rect 229008 543668 229060 543720
rect 260196 543668 260248 543720
rect 429476 543668 429528 543720
rect 78588 543600 78640 543652
rect 156420 543600 156472 543652
rect 205548 543600 205600 543652
rect 218704 543600 218756 543652
rect 227628 543600 227680 543652
rect 258080 543600 258132 543652
rect 61016 543532 61068 543584
rect 62028 543532 62080 543584
rect 70216 543532 70268 543584
rect 71320 543532 71372 543584
rect 82728 543532 82780 543584
rect 164700 543532 164752 543584
rect 208308 543532 208360 543584
rect 222844 543532 222896 543584
rect 230388 543532 230440 543584
rect 262220 543532 262272 543584
rect 127348 543464 127400 543516
rect 209044 543464 209096 543516
rect 209688 543464 209740 543516
rect 224500 543464 224552 543516
rect 231768 543464 231820 543516
rect 264336 543464 264388 543516
rect 123208 543396 123260 543448
rect 207664 543396 207716 543448
rect 211068 543396 211120 543448
rect 226984 543396 227036 543448
rect 233148 543396 233200 543448
rect 266452 543396 266504 543448
rect 119068 543328 119120 543380
rect 204904 543328 204956 543380
rect 212448 543328 212500 543380
rect 231124 543328 231176 543380
rect 233056 543328 233108 543380
rect 268476 543328 268528 543380
rect 117044 543260 117096 543312
rect 203524 543260 203576 543312
rect 215208 543260 215260 543312
rect 235264 543260 235316 543312
rect 235908 543260 235960 543312
rect 272616 543260 272668 543312
rect 93676 543192 93728 543244
rect 183376 543192 183428 543244
rect 210976 543192 211028 543244
rect 229100 543192 229152 543244
rect 234528 543192 234580 543244
rect 270592 543192 270644 543244
rect 56968 543124 57020 543176
rect 79692 543124 79744 543176
rect 95148 543124 95200 543176
rect 187516 543124 187568 543176
rect 204168 543124 204220 543176
rect 216220 543124 216272 543176
rect 216588 543124 216640 543176
rect 237380 543124 237432 543176
rect 238668 543124 238720 543176
rect 276756 543124 276808 543176
rect 67548 543056 67600 543108
rect 98368 543056 98420 543108
rect 99288 543056 99340 543108
rect 193772 543056 193824 543108
rect 213828 543056 213880 543108
rect 233240 543056 233292 543108
rect 237288 543056 237340 543108
rect 274732 543056 274784 543108
rect 57152 542988 57204 543040
rect 100392 542988 100444 543040
rect 102048 542988 102100 543040
rect 197912 542988 197964 543040
rect 202788 542988 202840 543040
rect 214564 542988 214616 543040
rect 217876 542988 217928 543040
rect 239404 542988 239456 543040
rect 240048 542988 240100 543040
rect 278872 542988 278924 543040
rect 104164 542920 104216 542972
rect 137744 542920 137796 542972
rect 70308 542852 70360 542904
rect 73436 542852 73488 542904
rect 105544 542852 105596 542904
rect 139860 542852 139912 542904
rect 100024 542784 100076 542836
rect 131488 542784 131540 542836
rect 133144 542784 133196 542836
rect 102784 542716 102836 542768
rect 135720 542716 135772 542768
rect 137376 542784 137428 542836
rect 204168 542920 204220 542972
rect 226248 542920 226300 542972
rect 256056 542920 256108 542972
rect 140044 542852 140096 542904
rect 200028 542852 200080 542904
rect 226156 542852 226208 542904
rect 253940 542852 253992 542904
rect 191748 542784 191800 542836
rect 223488 542784 223540 542836
rect 249800 542784 249852 542836
rect 140136 542716 140188 542768
rect 195888 542716 195940 542768
rect 224868 542716 224920 542768
rect 251916 542716 251968 542768
rect 131764 542648 131816 542700
rect 185492 542648 185544 542700
rect 222108 542648 222160 542700
rect 247776 542648 247828 542700
rect 108304 542580 108356 542632
rect 146024 542580 146076 542632
rect 65156 542512 65208 542564
rect 66168 542512 66220 542564
rect 108488 542512 108540 542564
rect 144000 542512 144052 542564
rect 145564 542512 145616 542564
rect 162676 542580 162728 542632
rect 220728 542580 220780 542632
rect 245660 542580 245712 542632
rect 148324 542512 148376 542564
rect 158536 542512 158588 542564
rect 217968 542512 218020 542564
rect 241520 542512 241572 542564
rect 106924 542444 106976 542496
rect 141884 542444 141936 542496
rect 101404 542376 101456 542428
rect 133604 542376 133656 542428
rect 135904 542376 135956 542428
rect 141424 542376 141476 542428
rect 154396 542444 154448 542496
rect 219348 542444 219400 542496
rect 243544 542444 243596 542496
rect 150164 542376 150216 542428
rect 429384 540948 429436 541000
rect 429476 540948 429528 541000
rect 56876 540812 56928 540864
rect 137284 540812 137336 540864
rect 56784 540744 56836 540796
rect 170036 540744 170088 540796
rect 56968 540676 57020 540728
rect 299756 540676 299808 540728
rect 59912 540608 59964 540660
rect 429384 540608 429436 540660
rect 57980 540540 58032 540592
rect 462320 540540 462372 540592
rect 59820 540472 59872 540524
rect 491760 540472 491812 540524
rect 59728 540404 59780 540456
rect 580356 540404 580408 540456
rect 59636 540336 59688 540388
rect 580724 540336 580776 540388
rect 58072 540268 58124 540320
rect 580264 540268 580316 540320
rect 58164 540200 58216 540252
rect 580448 540200 580500 540252
rect 59544 539724 59596 539776
rect 580908 539724 580960 539776
rect 57612 539656 57664 539708
rect 580540 539656 580592 539708
rect 57520 539588 57572 539640
rect 580816 539588 580868 539640
rect 57152 539180 57204 539232
rect 580264 539180 580316 539232
rect 33784 538228 33836 538280
rect 57428 538228 57480 538280
rect 19984 536800 20036 536852
rect 57428 536800 57480 536852
rect 17224 534080 17276 534132
rect 57428 534080 57480 534132
rect 28264 532720 28316 532772
rect 57428 532720 57480 532772
rect 48964 531360 49016 531412
rect 57428 531360 57480 531412
rect 4804 528572 4856 528624
rect 57428 528572 57480 528624
rect 53104 527144 53156 527196
rect 57428 527144 57480 527196
rect 46204 524424 46256 524476
rect 57428 524424 57480 524476
rect 282552 524424 282604 524476
rect 282644 524288 282696 524340
rect 4896 522996 4948 523048
rect 57428 522996 57480 523048
rect 51724 521704 51776 521756
rect 57428 521704 57480 521756
rect 43444 518916 43496 518968
rect 57428 518916 57480 518968
rect 4988 517488 5040 517540
rect 57428 517488 57480 517540
rect 50344 514768 50396 514820
rect 57428 514768 57480 514820
rect 282552 514768 282604 514820
rect 282644 514700 282696 514752
rect 35164 513340 35216 513392
rect 57428 513340 57480 513392
rect 5080 511980 5132 512032
rect 57428 511980 57480 512032
rect 282552 511980 282604 512032
rect 282644 511980 282696 512032
rect 39396 509260 39448 509312
rect 57428 509260 57480 509312
rect 33876 507832 33928 507884
rect 57428 507832 57480 507884
rect 282552 505112 282604 505164
rect 282644 504976 282696 505028
rect 37924 503684 37976 503736
rect 57428 503684 57480 503736
rect 28356 502324 28408 502376
rect 57428 502324 57480 502376
rect 32404 498176 32456 498228
rect 57428 498176 57480 498228
rect 282368 497496 282420 497548
rect 282552 497496 282604 497548
rect 3976 495456 4028 495508
rect 5172 495456 5224 495508
rect 20076 495456 20128 495508
rect 57428 495456 57480 495508
rect 15844 489880 15896 489932
rect 56692 489880 56744 489932
rect 3976 485800 4028 485852
rect 56692 485800 56744 485852
rect 282552 485800 282604 485852
rect 282644 485664 282696 485716
rect 3884 484372 3936 484424
rect 56692 484372 56744 484424
rect 282368 482944 282420 482996
rect 282644 482944 282696 482996
rect 56692 481720 56744 481772
rect 5172 481584 5224 481636
rect 56692 481584 56744 481636
rect 56692 481108 56744 481160
rect 2872 480156 2924 480208
rect 56508 480156 56560 480208
rect 4068 477436 4120 477488
rect 56508 477436 56560 477488
rect 3700 476008 3752 476060
rect 56508 476008 56560 476060
rect 3792 474648 3844 474700
rect 56508 474648 56560 474700
rect 3608 471928 3660 471980
rect 56508 471928 56560 471980
rect 31024 470500 31076 470552
rect 56508 470500 56560 470552
rect 14464 467780 14516 467832
rect 56508 467780 56560 467832
rect 282552 466420 282604 466472
rect 3516 466352 3568 466404
rect 56508 466352 56560 466404
rect 282644 466352 282696 466404
rect 21364 464992 21416 465044
rect 56508 464992 56560 465044
rect 282368 463632 282420 463684
rect 282644 463632 282696 463684
rect 13084 462272 13136 462324
rect 56508 462272 56560 462324
rect 3424 460844 3476 460896
rect 56600 460708 56652 460760
rect 24768 458124 24820 458176
rect 56600 458124 56652 458176
rect 10324 456696 10376 456748
rect 56600 456696 56652 456748
rect 42064 455336 42116 455388
rect 56600 455336 56652 455388
rect 3424 452548 3476 452600
rect 56600 452548 56652 452600
rect 282552 447108 282604 447160
rect 282644 447040 282696 447092
rect 282828 434664 282880 434716
rect 283012 434664 283064 434716
rect 281540 429156 281592 429208
rect 367100 429156 367152 429208
rect 281540 427796 281592 427848
rect 368480 427796 368532 427848
rect 281632 426504 281684 426556
rect 369860 426504 369912 426556
rect 281540 426436 281592 426488
rect 371240 426436 371292 426488
rect 281540 425076 281592 425128
rect 372620 425076 372672 425128
rect 281540 423648 281592 423700
rect 374000 423648 374052 423700
rect 281632 422356 281684 422408
rect 374092 422356 374144 422408
rect 281540 422288 281592 422340
rect 375380 422288 375432 422340
rect 281540 420928 281592 420980
rect 376760 420928 376812 420980
rect 281540 419500 281592 419552
rect 378140 419500 378192 419552
rect 59452 419432 59504 419484
rect 59912 419432 59964 419484
rect 281632 418208 281684 418260
rect 379520 418208 379572 418260
rect 281540 418140 281592 418192
rect 380900 418140 380952 418192
rect 282828 416780 282880 416832
rect 382280 416780 382332 416832
rect 282276 415420 282328 415472
rect 382372 415420 382424 415472
rect 281724 414060 281776 414112
rect 383844 414060 383896 414112
rect 282092 413992 282144 414044
rect 385040 413992 385092 414044
rect 282644 413924 282696 413976
rect 412640 413924 412692 413976
rect 383568 413856 383620 413908
rect 393136 413856 393188 413908
rect 325884 413788 325936 413840
rect 335176 413788 335228 413840
rect 345204 413788 345256 413840
rect 354496 413788 354548 413840
rect 378048 413788 378100 413840
rect 387340 413788 387392 413840
rect 396080 413788 396132 413840
rect 325792 413720 325844 413772
rect 335268 413720 335320 413772
rect 345112 413720 345164 413772
rect 354588 413720 354640 413772
rect 369768 413720 369820 413772
rect 378784 413720 378836 413772
rect 388352 413720 388404 413772
rect 397460 413720 397512 413772
rect 282644 413652 282696 413704
rect 368296 413652 368348 413704
rect 378048 413652 378100 413704
rect 386052 413652 386104 413704
rect 394700 413652 394752 413704
rect 281540 413584 281592 413636
rect 368756 413584 368808 413636
rect 368848 413584 368900 413636
rect 369860 413584 369912 413636
rect 379612 413584 379664 413636
rect 389640 413584 389692 413636
rect 318248 413516 318300 413568
rect 405740 413516 405792 413568
rect 281816 413448 281868 413500
rect 368848 413448 368900 413500
rect 368940 413448 368992 413500
rect 372988 413448 373040 413500
rect 382280 413448 382332 413500
rect 384948 413448 385000 413500
rect 393964 413448 394016 413500
rect 394700 413448 394752 413500
rect 395344 413448 395396 413500
rect 404360 413448 404412 413500
rect 287152 413380 287204 413432
rect 296536 413380 296588 413432
rect 306472 413380 306524 413432
rect 315856 413380 315908 413432
rect 318156 413380 318208 413432
rect 407120 413380 407172 413432
rect 282184 413312 282236 413364
rect 371976 413312 372028 413364
rect 381544 413312 381596 413364
rect 390928 413312 390980 413364
rect 391848 413312 391900 413364
rect 393136 413312 393188 413364
rect 401600 413312 401652 413364
rect 282828 413244 282880 413296
rect 386420 413244 386472 413296
rect 393964 413244 394016 413296
rect 403164 413244 403216 413296
rect 287060 413176 287112 413228
rect 296628 413176 296680 413228
rect 306380 413176 306432 413228
rect 315948 413176 316000 413228
rect 318064 413176 318116 413228
rect 408500 413176 408552 413228
rect 282368 413108 282420 413160
rect 368940 413108 368992 413160
rect 282000 413040 282052 413092
rect 287152 413040 287204 413092
rect 296536 413040 296588 413092
rect 306472 413040 306524 413092
rect 315856 413040 315908 413092
rect 325884 413040 325936 413092
rect 335176 413040 335228 413092
rect 345204 413040 345256 413092
rect 354496 413040 354548 413092
rect 368848 413040 368900 413092
rect 282460 412972 282512 413024
rect 287060 412972 287112 413024
rect 296628 412972 296680 413024
rect 306380 412972 306432 413024
rect 315948 412972 316000 413024
rect 325792 412972 325844 413024
rect 335268 412972 335320 413024
rect 345112 412972 345164 413024
rect 354588 412972 354640 413024
rect 382280 413108 382332 413160
rect 391756 413108 391808 413160
rect 391848 413108 391900 413160
rect 398840 413108 398892 413160
rect 375472 413040 375524 413092
rect 369308 412972 369360 413024
rect 374368 412972 374420 413024
rect 383476 412972 383528 413024
rect 400220 413040 400272 413092
rect 384948 412972 385000 413024
rect 282276 412904 282328 412956
rect 376576 412904 376628 412956
rect 386052 412904 386104 412956
rect 389640 412904 389692 412956
rect 397460 412904 397512 412956
rect 282736 412836 282788 412888
rect 393320 412836 393372 412888
rect 282092 412768 282144 412820
rect 394700 412768 394752 412820
rect 281540 412700 281592 412752
rect 281632 412700 281684 412752
rect 396080 412700 396132 412752
rect 405740 412632 405792 412684
rect 281540 412564 281592 412616
rect 281816 412496 281868 412548
rect 282736 412428 282788 412480
rect 281816 412360 281868 412412
rect 282092 412360 282144 412412
rect 284116 412360 284168 412412
rect 343732 412360 343784 412412
rect 281540 412292 281592 412344
rect 284024 412292 284076 412344
rect 343640 412292 343692 412344
rect 284208 412224 284260 412276
rect 345020 412224 345072 412276
rect 283472 412156 283524 412208
rect 346400 412156 346452 412208
rect 283380 412088 283432 412140
rect 347780 412088 347832 412140
rect 282920 412020 282972 412072
rect 349160 412020 349212 412072
rect 281908 411952 281960 412004
rect 350632 411952 350684 412004
rect 305644 411884 305696 411936
rect 419540 411884 419592 411936
rect 311164 411816 311216 411868
rect 397460 411816 397512 411868
rect 282092 411748 282144 411800
rect 388076 411748 388128 411800
rect 283012 411680 283064 411732
rect 391020 411680 391072 411732
rect 285036 411612 285088 411664
rect 399116 411612 399168 411664
rect 282092 411544 282144 411596
rect 398012 411544 398064 411596
rect 283104 411476 283156 411528
rect 400956 411476 401008 411528
rect 283288 411408 283340 411460
rect 401692 411408 401744 411460
rect 282460 411340 282512 411392
rect 282828 411340 282880 411392
rect 284944 411340 284996 411392
rect 404360 411340 404412 411392
rect 281908 411272 281960 411324
rect 283196 411272 283248 411324
rect 403256 411272 403308 411324
rect 282828 411204 282880 411256
rect 389272 411204 389324 411256
rect 281908 411136 281960 411188
rect 389732 411136 389784 411188
rect 298744 410728 298796 410780
rect 342260 410728 342312 410780
rect 283932 410660 283984 410712
rect 340880 410660 340932 410712
rect 282920 410592 282972 410644
rect 392308 410592 392360 410644
rect 283840 410524 283892 410576
rect 409972 410524 410024 410576
rect 281908 410116 281960 410168
rect 282092 407872 282144 407924
rect 282184 407872 282236 407924
rect 282644 407872 282696 407924
rect 281632 407804 281684 407856
rect 281632 407668 281684 407720
rect 281908 407668 281960 407720
rect 282000 407668 282052 407720
rect 281908 407532 281960 407584
rect 282000 407532 282052 407584
rect 282736 407532 282788 407584
rect 282828 404268 282880 404320
rect 311164 404268 311216 404320
rect 282276 402840 282328 402892
rect 282276 402636 282328 402688
rect 282184 402568 282236 402620
rect 285036 402568 285088 402620
rect 281632 401140 281684 401192
rect 283104 401140 283156 401192
rect 281632 400120 281684 400172
rect 283288 400120 283340 400172
rect 281632 399508 281684 399560
rect 283196 399508 283248 399560
rect 282184 398148 282236 398200
rect 284944 398148 284996 398200
rect 3148 395972 3200 396024
rect 56692 395972 56744 396024
rect 281632 394544 281684 394596
rect 283748 394544 283800 394596
rect 282184 393252 282236 393304
rect 282552 393252 282604 393304
rect 281816 393184 281868 393236
rect 282368 393184 282420 393236
rect 281632 393116 281684 393168
rect 283564 393116 283616 393168
rect 281632 392368 281684 392420
rect 283656 392368 283708 392420
rect 310428 389784 310480 389836
rect 338028 389784 338080 389836
rect 281632 388152 281684 388204
rect 283380 388152 283432 388204
rect 281632 386996 281684 387048
rect 283472 386996 283524 387048
rect 281724 386044 281776 386096
rect 284208 386044 284260 386096
rect 281632 385568 281684 385620
rect 284116 385568 284168 385620
rect 281632 384888 281684 384940
rect 284024 384888 284076 384940
rect 281724 383800 281776 383852
rect 281816 383732 281868 383784
rect 282368 383732 282420 383784
rect 282460 383732 282512 383784
rect 282184 383664 282236 383716
rect 282552 383664 282604 383716
rect 282828 383596 282880 383648
rect 298744 383596 298796 383648
rect 281724 382168 281776 382220
rect 339500 382168 339552 382220
rect 281632 381964 281684 382016
rect 283932 381964 283984 382016
rect 3240 380808 3292 380860
rect 57060 380808 57112 380860
rect 282828 380808 282880 380860
rect 338120 380808 338172 380860
rect 282828 379448 282880 379500
rect 336832 379448 336884 379500
rect 282828 378088 282880 378140
rect 336740 378088 336792 378140
rect 282184 378020 282236 378072
rect 335360 378020 335412 378072
rect 282828 376660 282880 376712
rect 333980 376660 334032 376712
rect 282828 375300 282880 375352
rect 332600 375300 332652 375352
rect 281908 373940 281960 373992
rect 282552 373940 282604 373992
rect 282828 373940 282880 373992
rect 331220 373940 331272 373992
rect 282184 373872 282236 373924
rect 329932 373872 329984 373924
rect 281816 373804 281868 373856
rect 282368 373804 282420 373856
rect 282460 373804 282512 373856
rect 281724 373736 281776 373788
rect 282828 372512 282880 372564
rect 329840 372512 329892 372564
rect 282828 371152 282880 371204
rect 328460 371152 328512 371204
rect 282184 371084 282236 371136
rect 327080 371084 327132 371136
rect 282828 369792 282880 369844
rect 325700 369792 325752 369844
rect 282828 368432 282880 368484
rect 324320 368432 324372 368484
rect 3148 367004 3200 367056
rect 15844 367004 15896 367056
rect 282828 367004 282880 367056
rect 322940 367004 322992 367056
rect 282184 366936 282236 366988
rect 321560 366936 321612 366988
rect 282828 365644 282880 365696
rect 330484 365644 330536 365696
rect 281724 364488 281776 364540
rect 281816 364420 281868 364472
rect 282368 364420 282420 364472
rect 282460 364420 282512 364472
rect 281908 364352 281960 364404
rect 282552 364352 282604 364404
rect 282828 364284 282880 364336
rect 329288 364284 329340 364336
rect 282184 362924 282236 362976
rect 282736 362924 282788 362976
rect 282828 362856 282880 362908
rect 329104 362856 329156 362908
rect 282736 362788 282788 362840
rect 327724 362788 327776 362840
rect 281724 361496 281776 361548
rect 326344 361496 326396 361548
rect 282828 360136 282880 360188
rect 324964 360136 325016 360188
rect 282736 360068 282788 360120
rect 323584 360068 323636 360120
rect 281908 358708 281960 358760
rect 322204 358708 322256 358760
rect 282092 354560 282144 354612
rect 282460 354560 282512 354612
rect 282828 349052 282880 349104
rect 297364 349052 297416 349104
rect 282828 347692 282880 347744
rect 294604 347692 294656 347744
rect 282276 347624 282328 347676
rect 291844 347624 291896 347676
rect 282092 346332 282144 346384
rect 290464 346332 290516 346384
rect 282828 344496 282880 344548
rect 287704 344496 287756 344548
rect 282552 343544 282604 343596
rect 301504 343544 301556 343596
rect 282736 343476 282788 343528
rect 286324 343476 286376 343528
rect 282828 342184 282880 342236
rect 316040 342184 316092 342236
rect 3424 338036 3476 338088
rect 57428 338036 57480 338088
rect 57796 336676 57848 336728
rect 59728 336676 59780 336728
rect 282184 333888 282236 333940
rect 307024 333888 307076 333940
rect 281632 333548 281684 333600
rect 283840 333548 283892 333600
rect 282000 331780 282052 331832
rect 282736 331780 282788 331832
rect 281632 331168 281684 331220
rect 320272 331168 320324 331220
rect 56968 330828 57020 330880
rect 59820 330828 59872 330880
rect 56600 330760 56652 330812
rect 56600 330624 56652 330676
rect 56876 330624 56928 330676
rect 57060 330420 57112 330472
rect 281632 329740 281684 329792
rect 318800 329740 318852 329792
rect 281540 329672 281592 329724
rect 297456 329672 297508 329724
rect 56968 329332 57020 329384
rect 57796 329332 57848 329384
rect 57060 329196 57112 329248
rect 57796 329196 57848 329248
rect 281540 328380 281592 328432
rect 302884 328380 302936 328432
rect 281540 327020 281592 327072
rect 318248 327020 318300 327072
rect 282092 326408 282144 326460
rect 282736 326408 282788 326460
rect 281908 326340 281960 326392
rect 282184 326340 282236 326392
rect 282276 326340 282328 326392
rect 282644 326340 282696 326392
rect 281816 326272 281868 326324
rect 282736 326272 282788 326324
rect 281540 325592 281592 325644
rect 318156 325592 318208 325644
rect 56600 325456 56652 325508
rect 57980 325456 58032 325508
rect 56600 325320 56652 325372
rect 56876 325320 56928 325372
rect 56876 325184 56928 325236
rect 57520 325184 57572 325236
rect 57888 325116 57940 325168
rect 59544 325116 59596 325168
rect 57704 325048 57756 325100
rect 59636 325048 59688 325100
rect 3240 324232 3292 324284
rect 32404 324232 32456 324284
rect 281540 324232 281592 324284
rect 318064 324232 318116 324284
rect 281540 322872 281592 322924
rect 305644 322872 305696 322924
rect 284300 322192 284352 322244
rect 285588 322192 285640 322244
rect 337752 322192 337804 322244
rect 282828 321512 282880 321564
rect 284300 321512 284352 321564
rect 282828 320968 282880 321020
rect 337384 320968 337436 321020
rect 338028 320968 338080 321020
rect 282184 320900 282236 320952
rect 419540 320900 419592 320952
rect 282552 320832 282604 320884
rect 419816 320832 419868 320884
rect 56600 320764 56652 320816
rect 580908 320764 580960 320816
rect 57980 320696 58032 320748
rect 580172 320696 580224 320748
rect 57520 320628 57572 320680
rect 580724 320628 580776 320680
rect 57612 320560 57664 320612
rect 280068 320560 280120 320612
rect 282368 320560 282420 320612
rect 419724 320560 419776 320612
rect 59544 320492 59596 320544
rect 279976 320492 280028 320544
rect 282000 320492 282052 320544
rect 419632 320492 419684 320544
rect 59728 320424 59780 320476
rect 280068 320424 280120 320476
rect 282460 320424 282512 320476
rect 416412 320424 416464 320476
rect 282276 320356 282328 320408
rect 420184 320356 420236 320408
rect 282736 320288 282788 320340
rect 419908 320288 419960 320340
rect 282092 320220 282144 320272
rect 420000 320220 420052 320272
rect 56876 320084 56928 320136
rect 580816 320084 580868 320136
rect 59820 320016 59872 320068
rect 580632 320016 580684 320068
rect 59636 319948 59688 320000
rect 580448 319948 580500 320000
rect 59912 319880 59964 319932
rect 580356 319880 580408 319932
rect 4068 318724 4120 318776
rect 64788 318724 64840 318776
rect 82728 318724 82780 318776
rect 193220 318724 193272 318776
rect 338028 318724 338080 318776
rect 344008 318724 344060 318776
rect 50436 318656 50488 318708
rect 88156 318656 88208 318708
rect 88248 318656 88300 318708
rect 201040 318656 201092 318708
rect 8208 318588 8260 318640
rect 72516 318588 72568 318640
rect 45468 318520 45520 318572
rect 55220 318520 55272 318572
rect 64788 318520 64840 318572
rect 94412 318520 94464 318572
rect 10968 318452 11020 318504
rect 76472 318452 76524 318504
rect 86868 318452 86920 318504
rect 88248 318452 88300 318504
rect 89536 318452 89588 318504
rect 204904 318588 204956 318640
rect 94596 318520 94648 318572
rect 212724 318520 212776 318572
rect 96528 318452 96580 318504
rect 216588 318452 216640 318504
rect 42708 318384 42760 318436
rect 129004 318384 129056 318436
rect 134524 318384 134576 318436
rect 255504 318384 255556 318436
rect 16488 318316 16540 318368
rect 86224 318316 86276 318368
rect 94412 318316 94464 318368
rect 107568 318316 107620 318368
rect 107660 318316 107712 318368
rect 224408 318316 224460 318368
rect 20628 318248 20680 318300
rect 92020 318248 92072 318300
rect 93768 318248 93820 318300
rect 94596 318248 94648 318300
rect 103428 318248 103480 318300
rect 228272 318248 228324 318300
rect 21916 318180 21968 318232
rect 93952 318180 94004 318232
rect 107568 318180 107620 318232
rect 234160 318180 234212 318232
rect 24768 318112 24820 318164
rect 99840 318112 99892 318164
rect 100668 318112 100720 318164
rect 26148 318044 26200 318096
rect 101772 318044 101824 318096
rect 107476 318112 107528 318164
rect 236092 318112 236144 318164
rect 107660 318044 107712 318096
rect 114468 318044 114520 318096
rect 245844 318044 245896 318096
rect 344008 318044 344060 318096
rect 347780 318044 347832 318096
rect 32404 317976 32456 318028
rect 78404 317976 78456 318028
rect 79968 317976 80020 318028
rect 189356 317976 189408 318028
rect 39304 317908 39356 317960
rect 68652 317908 68704 317960
rect 74448 317908 74500 317960
rect 181536 317908 181588 317960
rect 2688 317840 2740 317892
rect 62856 317840 62908 317892
rect 64788 317840 64840 317892
rect 72976 317840 73028 317892
rect 177672 317840 177724 317892
rect 42064 317772 42116 317824
rect 45468 317772 45520 317824
rect 55220 317772 55272 317824
rect 67548 317772 67600 317824
rect 169852 317772 169904 317824
rect 64788 317704 64840 317756
rect 165988 317704 166040 317756
rect 62028 317636 62080 317688
rect 160192 317636 160244 317688
rect 50988 317568 51040 317620
rect 142620 317568 142672 317620
rect 48136 317500 48188 317552
rect 136824 317500 136876 317552
rect 39948 317432 40000 317484
rect 124772 317432 124824 317484
rect 124864 317432 124916 317484
rect 146576 317432 146628 317484
rect 56692 311788 56744 311840
rect 580172 311788 580224 311840
rect 3332 309068 3384 309120
rect 20076 309068 20128 309120
rect 74448 299616 74500 299668
rect 74448 299480 74500 299532
rect 56784 299412 56836 299464
rect 579804 299412 579856 299464
rect 74264 298052 74316 298104
rect 74448 298052 74500 298104
rect 3424 295264 3476 295316
rect 57336 295264 57388 295316
rect 74264 288396 74316 288448
rect 74356 288396 74408 288448
rect 3424 280100 3476 280152
rect 37924 280100 37976 280152
rect 57152 275952 57204 276004
rect 580172 275952 580224 276004
rect 74264 269084 74316 269136
rect 74356 269084 74408 269136
rect 2872 266296 2924 266348
rect 28356 266296 28408 266348
rect 147588 263780 147640 263832
rect 154488 263780 154540 263832
rect 86868 263712 86920 263764
rect 115940 263644 115992 263696
rect 118792 263644 118844 263696
rect 86868 263576 86920 263628
rect 3424 252492 3476 252544
rect 57244 252492 57296 252544
rect 59452 252492 59504 252544
rect 579804 252492 579856 252544
rect 74264 249772 74316 249824
rect 74448 249772 74500 249824
rect 74356 241476 74408 241528
rect 74448 241476 74500 241528
rect 3424 237328 3476 237380
rect 39396 237328 39448 237380
rect 74264 230460 74316 230512
rect 74448 230460 74500 230512
rect 66260 227944 66312 227996
rect 75828 227944 75880 227996
rect 147588 227876 147640 227928
rect 154488 227876 154540 227928
rect 86868 227808 86920 227860
rect 115940 227740 115992 227792
rect 118792 227740 118844 227792
rect 86868 227672 86920 227724
rect 3148 223524 3200 223576
rect 33876 223524 33928 223576
rect 69388 216928 69440 216980
rect 77208 216928 77260 216980
rect 89536 216860 89588 216912
rect 91744 216860 91796 216912
rect 147588 216860 147640 216912
rect 154488 216860 154540 216912
rect 115940 216724 115992 216776
rect 118792 216724 118844 216776
rect 2780 208156 2832 208208
rect 5080 208156 5132 208208
rect 59360 205572 59412 205624
rect 579804 205572 579856 205624
rect 89352 202852 89404 202904
rect 89536 202852 89588 202904
rect 74264 201424 74316 201476
rect 74448 201424 74500 201476
rect 89352 195984 89404 196036
rect 89444 195848 89496 195900
rect 2872 194488 2924 194540
rect 50344 194488 50396 194540
rect 74264 191836 74316 191888
rect 74356 191836 74408 191888
rect 74356 183540 74408 183592
rect 74448 183540 74500 183592
rect 74264 182112 74316 182164
rect 74448 182112 74500 182164
rect 69388 181024 69440 181076
rect 77208 181024 77260 181076
rect 86868 180888 86920 180940
rect 3240 180752 3292 180804
rect 35164 180752 35216 180804
rect 86868 180752 86920 180804
rect 89444 173884 89496 173936
rect 89628 173884 89680 173936
rect 66260 170008 66312 170060
rect 75828 170008 75880 170060
rect 147588 169940 147640 169992
rect 154488 169940 154540 169992
rect 86868 169872 86920 169924
rect 115940 169804 115992 169856
rect 118792 169804 118844 169856
rect 86868 169736 86920 169788
rect 2780 165452 2832 165504
rect 4988 165452 5040 165504
rect 74264 162800 74316 162852
rect 74448 162800 74500 162852
rect 59084 158652 59136 158704
rect 579804 158652 579856 158704
rect 89444 157428 89496 157480
rect 89444 157292 89496 157344
rect 89260 154504 89312 154556
rect 89536 154504 89588 154556
rect 3148 151716 3200 151768
rect 51724 151716 51776 151768
rect 74448 143488 74500 143540
rect 74632 143488 74684 143540
rect 89444 137980 89496 138032
rect 89536 137844 89588 137896
rect 3240 136552 3292 136604
rect 43444 136552 43496 136604
rect 57428 135192 57480 135244
rect 580172 135192 580224 135244
rect 89536 128392 89588 128444
rect 89444 128256 89496 128308
rect 56968 124108 57020 124160
rect 580172 124108 580224 124160
rect 89444 124040 89496 124092
rect 89628 124040 89680 124092
rect 2780 122340 2832 122392
rect 4896 122340 4948 122392
rect 89628 118668 89680 118720
rect 89536 118532 89588 118584
rect 74356 114520 74408 114572
rect 74724 114520 74776 114572
rect 59176 111732 59228 111784
rect 579804 111732 579856 111784
rect 89536 109080 89588 109132
rect 3240 108944 3292 108996
rect 53104 108944 53156 108996
rect 89444 108944 89496 108996
rect 74356 106360 74408 106412
rect 74448 106360 74500 106412
rect 74264 104796 74316 104848
rect 74448 104796 74500 104848
rect 89260 104796 89312 104848
rect 89444 104796 89496 104848
rect 74264 95208 74316 95260
rect 74356 95208 74408 95260
rect 89260 95208 89312 95260
rect 89352 95208 89404 95260
rect 3424 93780 3476 93832
rect 46204 93780 46256 93832
rect 57060 88272 57112 88324
rect 580172 88272 580224 88324
rect 74356 87048 74408 87100
rect 74448 87048 74500 87100
rect 74264 85484 74316 85536
rect 74448 85484 74500 85536
rect 89536 80112 89588 80164
rect 89536 79976 89588 80028
rect 2780 79024 2832 79076
rect 4804 79024 4856 79076
rect 89628 76100 89680 76152
rect 91744 76100 91796 76152
rect 147588 76100 147640 76152
rect 154488 76100 154540 76152
rect 115940 75964 115992 76016
rect 118792 75964 118844 76016
rect 74264 75896 74316 75948
rect 74356 75896 74408 75948
rect 74356 67668 74408 67720
rect 74448 67668 74500 67720
rect 74264 66172 74316 66224
rect 74448 66172 74500 66224
rect 3332 64812 3384 64864
rect 28264 64812 28316 64864
rect 59268 64812 59320 64864
rect 579804 64812 579856 64864
rect 74264 56584 74316 56636
rect 74448 56584 74500 56636
rect 3424 51008 3476 51060
rect 48964 51008 49016 51060
rect 89444 51008 89496 51060
rect 89628 51008 89680 51060
rect 89352 48220 89404 48272
rect 89628 48220 89680 48272
rect 74264 46860 74316 46912
rect 74448 46860 74500 46912
rect 57704 41352 57756 41404
rect 580172 41352 580224 41404
rect 89352 38632 89404 38684
rect 89536 38632 89588 38684
rect 74264 37272 74316 37324
rect 74356 37272 74408 37324
rect 3424 35844 3476 35896
rect 17224 35844 17276 35896
rect 57796 30268 57848 30320
rect 580172 30268 580224 30320
rect 74264 27548 74316 27600
rect 74448 27548 74500 27600
rect 89168 26188 89220 26240
rect 89260 26188 89312 26240
rect 2872 22040 2924 22092
rect 33784 22040 33836 22092
rect 89168 21360 89220 21412
rect 89444 21360 89496 21412
rect 74080 17960 74132 18012
rect 74264 17960 74316 18012
rect 57888 17892 57940 17944
rect 579804 17892 579856 17944
rect 74080 9664 74132 9716
rect 74264 9664 74316 9716
rect 89352 8304 89404 8356
rect 89444 8304 89496 8356
rect 3424 8236 3476 8288
rect 19984 8236 20036 8288
rect 60004 6400 60056 6452
rect 157340 6400 157392 6452
rect 108764 6332 108816 6384
rect 237380 6332 237432 6384
rect 112352 6264 112404 6316
rect 242900 6264 242952 6316
rect 115940 6196 115992 6248
rect 248420 6196 248472 6248
rect 123024 6128 123076 6180
rect 260840 6128 260892 6180
rect 86132 5584 86184 5636
rect 86868 5584 86920 5636
rect 93860 5516 93912 5568
rect 103612 5516 103664 5568
rect 105084 5516 105136 5568
rect 109040 5516 109092 5568
rect 60740 5380 60792 5432
rect 78588 5380 78640 5432
rect 12440 5312 12492 5364
rect 80060 5448 80112 5500
rect 80244 5448 80296 5500
rect 190460 5448 190512 5500
rect 83832 5380 83884 5432
rect 195980 5380 196032 5432
rect 87328 5312 87380 5364
rect 202880 5312 202932 5364
rect 52828 5244 52880 5296
rect 60740 5244 60792 5296
rect 78588 5244 78640 5296
rect 93860 5244 93912 5296
rect 109040 5244 109092 5296
rect 219440 5244 219492 5296
rect 22008 5176 22060 5228
rect 95240 5176 95292 5228
rect 98092 5176 98144 5228
rect 105084 5176 105136 5228
rect 105176 5176 105228 5228
rect 231860 5176 231912 5228
rect 26700 5108 26752 5160
rect 81900 5108 81952 5160
rect 82084 5108 82136 5160
rect 103520 5108 103572 5160
rect 103612 5108 103664 5160
rect 30288 5040 30340 5092
rect 81992 5040 82044 5092
rect 33876 4972 33928 5024
rect 86868 5040 86920 5092
rect 109132 5040 109184 5092
rect 127808 5108 127860 5160
rect 124864 5040 124916 5092
rect 130200 5040 130252 5092
rect 137468 5108 137520 5160
rect 266360 5108 266412 5160
rect 114560 4972 114612 5024
rect 119436 4972 119488 5024
rect 134524 4972 134576 5024
rect 134616 4972 134668 5024
rect 137192 4972 137244 5024
rect 269120 5040 269172 5092
rect 271880 4972 271932 5024
rect 37372 4904 37424 4956
rect 81992 4904 82044 4956
rect 86776 4904 86828 4956
rect 120080 4904 120132 4956
rect 129004 4904 129056 4956
rect 270500 4904 270552 4956
rect 40960 4836 41012 4888
rect 78864 4836 78916 4888
rect 86868 4836 86920 4888
rect 126980 4836 127032 4888
rect 127072 4836 127124 4888
rect 137468 4836 137520 4888
rect 137560 4836 137612 4888
rect 276020 4836 276072 4888
rect 44548 4768 44600 4820
rect 132500 4768 132552 4820
rect 132592 4768 132644 4820
rect 134616 4768 134668 4820
rect 134892 4768 134944 4820
rect 278780 4768 278832 4820
rect 67088 4700 67140 4752
rect 67548 4700 67600 4752
rect 76656 4700 76708 4752
rect 184940 4700 184992 4752
rect 73068 4632 73120 4684
rect 179420 4632 179472 4684
rect 69480 4564 69532 4616
rect 172520 4564 172572 4616
rect 65984 4496 66036 4548
rect 167000 4496 167052 4548
rect 62396 4428 62448 4480
rect 161480 4428 161532 4480
rect 58808 4360 58860 4412
rect 155960 4360 156012 4412
rect 55220 4292 55272 4344
rect 150440 4292 150492 4344
rect 51632 4224 51684 4276
rect 143540 4224 143592 4276
rect 48228 4156 48280 4208
rect 138020 4156 138072 4208
rect 8852 4088 8904 4140
rect 71780 4088 71832 4140
rect 71872 4088 71924 4140
rect 72976 4088 73028 4140
rect 73068 4088 73120 4140
rect 74540 4088 74592 4140
rect 13636 4020 13688 4072
rect 81348 4088 81400 4140
rect 81440 4088 81492 4140
rect 82728 4088 82780 4140
rect 82820 4088 82872 4140
rect 86040 4088 86092 4140
rect 79048 4020 79100 4072
rect 79968 4020 80020 4072
rect 80060 4020 80112 4072
rect 186320 4088 186372 4140
rect 89536 4020 89588 4072
rect 194600 4020 194652 4072
rect 14832 3952 14884 4004
rect 84200 3952 84252 4004
rect 84936 3952 84988 4004
rect 89444 3952 89496 4004
rect 89720 3952 89772 4004
rect 93216 3952 93268 4004
rect 18328 3884 18380 3936
rect 89628 3884 89680 3936
rect 89904 3884 89956 3936
rect 198740 3952 198792 4004
rect 93860 3884 93912 3936
rect 205640 3884 205692 3936
rect 23112 3748 23164 3800
rect 95516 3816 95568 3868
rect 27896 3748 27948 3800
rect 95700 3748 95752 3800
rect 96528 3748 96580 3800
rect 96896 3816 96948 3868
rect 102600 3748 102652 3800
rect 102784 3816 102836 3868
rect 103428 3816 103480 3868
rect 103520 3816 103572 3868
rect 104900 3816 104952 3868
rect 106004 3748 106056 3800
rect 31484 3680 31536 3732
rect 108212 3816 108264 3868
rect 106188 3748 106240 3800
rect 218060 3816 218112 3868
rect 106280 3680 106332 3732
rect 113180 3748 113232 3800
rect 113548 3748 113600 3800
rect 114468 3748 114520 3800
rect 114744 3748 114796 3800
rect 115848 3748 115900 3800
rect 116032 3748 116084 3800
rect 238760 3748 238812 3800
rect 108488 3680 108540 3732
rect 110420 3680 110472 3732
rect 111156 3680 111208 3732
rect 241520 3680 241572 3732
rect 36176 3612 36228 3664
rect 32680 3544 32732 3596
rect 106280 3544 106332 3596
rect 106372 3544 106424 3596
rect 107568 3544 107620 3596
rect 109960 3544 110012 3596
rect 113732 3544 113784 3596
rect 1676 3476 1728 3528
rect 2688 3476 2740 3528
rect 2872 3476 2924 3528
rect 4068 3476 4120 3528
rect 7656 3476 7708 3528
rect 8208 3476 8260 3528
rect 10048 3476 10100 3528
rect 10968 3476 11020 3528
rect 16028 3476 16080 3528
rect 16488 3476 16540 3528
rect 19524 3476 19576 3528
rect 20628 3476 20680 3528
rect 20720 3476 20772 3528
rect 21916 3476 21968 3528
rect 24308 3476 24360 3528
rect 24768 3476 24820 3528
rect 25504 3476 25556 3528
rect 26148 3476 26200 3528
rect 34980 3476 35032 3528
rect 113640 3476 113692 3528
rect 114008 3612 114060 3664
rect 114100 3544 114152 3596
rect 116032 3544 116084 3596
rect 117136 3612 117188 3664
rect 117320 3544 117372 3596
rect 118240 3544 118292 3596
rect 120632 3612 120684 3664
rect 121368 3612 121420 3664
rect 121828 3612 121880 3664
rect 122748 3612 122800 3664
rect 122840 3612 122892 3664
rect 252560 3612 252612 3664
rect 118700 3476 118752 3528
rect 122656 3476 122708 3528
rect 251180 3544 251232 3596
rect 124220 3476 124272 3528
rect 262220 3476 262272 3528
rect 11244 3408 11296 3460
rect 32404 3408 32456 3460
rect 42156 3408 42208 3460
rect 42708 3408 42760 3460
rect 42800 3408 42852 3460
rect 122932 3408 122984 3460
rect 125416 3408 125468 3460
rect 264980 3408 265032 3460
rect 6460 3340 6512 3392
rect 4068 3272 4120 3324
rect 61016 3272 61068 3324
rect 61200 3340 61252 3392
rect 62028 3340 62080 3392
rect 62120 3340 62172 3392
rect 66352 3340 66404 3392
rect 68284 3340 68336 3392
rect 70400 3272 70452 3324
rect 70676 3272 70728 3324
rect 75092 3272 75144 3324
rect 75276 3340 75328 3392
rect 175280 3340 175332 3392
rect 171140 3272 171192 3324
rect 572 3204 624 3256
rect 61384 3204 61436 3256
rect 63592 3204 63644 3256
rect 162860 3204 162912 3256
rect 5264 3136 5316 3188
rect 17224 3068 17276 3120
rect 38568 3136 38620 3188
rect 42800 3136 42852 3188
rect 46940 3136 46992 3188
rect 48136 3136 48188 3188
rect 50528 3136 50580 3188
rect 50988 3136 51040 3188
rect 56416 3136 56468 3188
rect 151820 3136 151872 3188
rect 29092 3000 29144 3052
rect 39304 3068 39356 3120
rect 50436 3068 50488 3120
rect 57612 3068 57664 3120
rect 153200 3068 153252 3120
rect 54024 3000 54076 3052
rect 147680 3000 147732 3052
rect 49332 2932 49384 2984
rect 139400 2932 139452 2984
rect 42064 2864 42116 2916
rect 45744 2864 45796 2916
rect 133972 2864 134024 2916
rect 43352 2796 43404 2848
rect 129832 2796 129884 2848
rect 88524 1096 88576 1148
rect 89352 1096 89404 1148
rect 67088 552 67140 604
rect 67180 552 67232 604
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 699718 8156 703520
rect 24320 699718 24348 703520
rect 40512 699990 40540 703520
rect 58624 701004 58676 701010
rect 58624 700946 58676 700952
rect 57796 700868 57848 700874
rect 57796 700810 57848 700816
rect 40500 699984 40552 699990
rect 40500 699926 40552 699932
rect 42064 699984 42116 699990
rect 42064 699926 42116 699932
rect 8116 699712 8168 699718
rect 8116 699654 8168 699660
rect 10324 699712 10376 699718
rect 10324 699654 10376 699660
rect 24308 699712 24360 699718
rect 24308 699654 24360 699660
rect 24768 699712 24820 699718
rect 24768 699654 24820 699660
rect 3422 682272 3478 682281
rect 3422 682207 3478 682216
rect 3054 653576 3110 653585
rect 3054 653511 3110 653520
rect 3068 652798 3096 653511
rect 3056 652792 3108 652798
rect 3056 652734 3108 652740
rect 3330 596048 3386 596057
rect 3330 595983 3386 595992
rect 3344 594862 3372 595983
rect 3332 594856 3384 594862
rect 3332 594798 3384 594804
rect 2870 481128 2926 481137
rect 2870 481063 2926 481072
rect 2884 480214 2912 481063
rect 2872 480208 2924 480214
rect 2872 480150 2924 480156
rect 3436 460902 3464 682207
rect 3514 667992 3570 668001
rect 3514 667927 3516 667936
rect 3568 667927 3570 667936
rect 3516 667898 3568 667904
rect 3514 624880 3570 624889
rect 3514 624815 3570 624824
rect 3528 466410 3556 624815
rect 3606 610464 3662 610473
rect 3606 610399 3662 610408
rect 3620 610026 3648 610399
rect 3608 610020 3660 610026
rect 3608 609962 3660 609968
rect 3606 567352 3662 567361
rect 3606 567287 3662 567296
rect 3620 471986 3648 567287
rect 3698 553072 3754 553081
rect 3698 553007 3754 553016
rect 3712 476066 3740 553007
rect 3790 538656 3846 538665
rect 3790 538591 3846 538600
rect 3700 476060 3752 476066
rect 3700 476002 3752 476008
rect 3804 474706 3832 538591
rect 4804 528624 4856 528630
rect 4804 528566 4856 528572
rect 4066 509960 4122 509969
rect 4066 509895 4122 509904
rect 3974 495544 4030 495553
rect 3974 495479 3976 495488
rect 4028 495479 4030 495488
rect 3976 495450 4028 495456
rect 3976 485852 4028 485858
rect 3976 485794 4028 485800
rect 3884 484424 3936 484430
rect 3884 484366 3936 484372
rect 3792 474700 3844 474706
rect 3792 474642 3844 474648
rect 3608 471980 3660 471986
rect 3608 471922 3660 471928
rect 3516 466404 3568 466410
rect 3516 466346 3568 466352
rect 3424 460896 3476 460902
rect 3424 460838 3476 460844
rect 3424 452600 3476 452606
rect 3424 452542 3476 452548
rect 3436 452441 3464 452542
rect 3422 452432 3478 452441
rect 3422 452367 3478 452376
rect 3896 423745 3924 484366
rect 3988 438025 4016 485794
rect 4080 477494 4108 509895
rect 4068 477488 4120 477494
rect 4068 477430 4120 477436
rect 3974 438016 4030 438025
rect 3974 437951 4030 437960
rect 3882 423736 3938 423745
rect 3882 423671 3938 423680
rect 3148 396024 3200 396030
rect 3148 395966 3200 395972
rect 3160 395049 3188 395966
rect 3146 395040 3202 395049
rect 3146 394975 3202 394984
rect 3240 380860 3292 380866
rect 3240 380802 3292 380808
rect 3252 380633 3280 380802
rect 3238 380624 3294 380633
rect 3238 380559 3294 380568
rect 3148 367056 3200 367062
rect 3148 366998 3200 367004
rect 3160 366217 3188 366998
rect 3146 366208 3202 366217
rect 3146 366143 3202 366152
rect 3424 338088 3476 338094
rect 3424 338030 3476 338036
rect 3436 337521 3464 338030
rect 3422 337512 3478 337521
rect 3422 337447 3478 337456
rect 3240 324284 3292 324290
rect 3240 324226 3292 324232
rect 3252 323105 3280 324226
rect 3238 323096 3294 323105
rect 3238 323031 3294 323040
rect 4068 318776 4120 318782
rect 4068 318718 4120 318724
rect 2688 317892 2740 317898
rect 2688 317834 2740 317840
rect 2700 3534 2728 317834
rect 3332 309120 3384 309126
rect 3332 309062 3384 309068
rect 3344 308825 3372 309062
rect 3330 308816 3386 308825
rect 3330 308751 3386 308760
rect 3424 295316 3476 295322
rect 3424 295258 3476 295264
rect 3436 294409 3464 295258
rect 3422 294400 3478 294409
rect 3422 294335 3478 294344
rect 3424 280152 3476 280158
rect 3422 280120 3424 280129
rect 3476 280120 3478 280129
rect 3422 280055 3478 280064
rect 2872 266348 2924 266354
rect 2872 266290 2924 266296
rect 2884 265713 2912 266290
rect 2870 265704 2926 265713
rect 2870 265639 2926 265648
rect 3424 252544 3476 252550
rect 3424 252486 3476 252492
rect 3436 251297 3464 252486
rect 3422 251288 3478 251297
rect 3422 251223 3478 251232
rect 3424 237380 3476 237386
rect 3424 237322 3476 237328
rect 3436 237017 3464 237322
rect 3422 237008 3478 237017
rect 3422 236943 3478 236952
rect 3148 223576 3200 223582
rect 3148 223518 3200 223524
rect 3160 222601 3188 223518
rect 3146 222592 3202 222601
rect 3146 222527 3202 222536
rect 2780 208208 2832 208214
rect 2778 208176 2780 208185
rect 2832 208176 2834 208185
rect 2778 208111 2834 208120
rect 2872 194540 2924 194546
rect 2872 194482 2924 194488
rect 2884 193905 2912 194482
rect 2870 193896 2926 193905
rect 2870 193831 2926 193840
rect 3240 180804 3292 180810
rect 3240 180746 3292 180752
rect 3252 179489 3280 180746
rect 3238 179480 3294 179489
rect 3238 179415 3294 179424
rect 2780 165504 2832 165510
rect 2780 165446 2832 165452
rect 2792 165073 2820 165446
rect 2778 165064 2834 165073
rect 2778 164999 2834 165008
rect 3148 151768 3200 151774
rect 3148 151710 3200 151716
rect 3160 150793 3188 151710
rect 3146 150784 3202 150793
rect 3146 150719 3202 150728
rect 3240 136604 3292 136610
rect 3240 136546 3292 136552
rect 3252 136377 3280 136546
rect 3238 136368 3294 136377
rect 3238 136303 3294 136312
rect 2780 122392 2832 122398
rect 2780 122334 2832 122340
rect 2792 122097 2820 122334
rect 2778 122088 2834 122097
rect 2778 122023 2834 122032
rect 3240 108996 3292 109002
rect 3240 108938 3292 108944
rect 3252 107681 3280 108938
rect 3238 107672 3294 107681
rect 3238 107607 3294 107616
rect 3424 93832 3476 93838
rect 3424 93774 3476 93780
rect 3436 93265 3464 93774
rect 3422 93256 3478 93265
rect 3422 93191 3478 93200
rect 2780 79076 2832 79082
rect 2780 79018 2832 79024
rect 2792 78985 2820 79018
rect 2778 78976 2834 78985
rect 2778 78911 2834 78920
rect 3332 64864 3384 64870
rect 3332 64806 3384 64812
rect 3344 64569 3372 64806
rect 3330 64560 3386 64569
rect 3330 64495 3386 64504
rect 3424 51060 3476 51066
rect 3424 51002 3476 51008
rect 3436 50153 3464 51002
rect 3422 50144 3478 50153
rect 3422 50079 3478 50088
rect 3424 35896 3476 35902
rect 3422 35864 3424 35873
rect 3476 35864 3478 35873
rect 3422 35799 3478 35808
rect 2872 22092 2924 22098
rect 2872 22034 2924 22040
rect 2884 21457 2912 22034
rect 2870 21448 2926 21457
rect 2870 21383 2926 21392
rect 3424 8288 3476 8294
rect 3424 8230 3476 8236
rect 3436 7177 3464 8230
rect 3422 7168 3478 7177
rect 3422 7103 3478 7112
rect 4080 3534 4108 318718
rect 4816 79082 4844 528566
rect 4896 523048 4948 523054
rect 4896 522990 4948 522996
rect 4908 122398 4936 522990
rect 4988 517540 5040 517546
rect 4988 517482 5040 517488
rect 5000 165510 5028 517482
rect 5080 512032 5132 512038
rect 5080 511974 5132 511980
rect 5092 208214 5120 511974
rect 5172 495508 5224 495514
rect 5172 495450 5224 495456
rect 5184 481642 5212 495450
rect 5172 481636 5224 481642
rect 5172 481578 5224 481584
rect 10336 456754 10364 699654
rect 21364 667956 21416 667962
rect 21364 667898 21416 667904
rect 13084 652792 13136 652798
rect 13084 652734 13136 652740
rect 13096 462330 13124 652734
rect 14464 594856 14516 594862
rect 14464 594798 14516 594804
rect 14476 467838 14504 594798
rect 19984 536852 20036 536858
rect 19984 536794 20036 536800
rect 17224 534132 17276 534138
rect 17224 534074 17276 534080
rect 15844 489932 15896 489938
rect 15844 489874 15896 489880
rect 14464 467832 14516 467838
rect 14464 467774 14516 467780
rect 13084 462324 13136 462330
rect 13084 462266 13136 462272
rect 10324 456748 10376 456754
rect 10324 456690 10376 456696
rect 15856 367062 15884 489874
rect 15844 367056 15896 367062
rect 15844 366998 15896 367004
rect 8208 318640 8260 318646
rect 8208 318582 8260 318588
rect 5080 208208 5132 208214
rect 5080 208150 5132 208156
rect 4988 165504 5040 165510
rect 4988 165446 5040 165452
rect 4896 122392 4948 122398
rect 4896 122334 4948 122340
rect 4804 79076 4856 79082
rect 4804 79018 4856 79024
rect 8220 3534 8248 318582
rect 10968 318504 11020 318510
rect 10968 318446 11020 318452
rect 8852 4140 8904 4146
rect 8852 4082 8904 4088
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 2688 3528 2740 3534
rect 2688 3470 2740 3476
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 4068 3528 4120 3534
rect 4068 3470 4120 3476
rect 7656 3528 7708 3534
rect 7656 3470 7708 3476
rect 8208 3528 8260 3534
rect 8208 3470 8260 3476
rect 572 3256 624 3262
rect 572 3198 624 3204
rect 584 480 612 3198
rect 1688 480 1716 3470
rect 2884 480 2912 3470
rect 6460 3392 6512 3398
rect 6460 3334 6512 3340
rect 4068 3324 4120 3330
rect 4068 3266 4120 3272
rect 4080 480 4108 3266
rect 5264 3188 5316 3194
rect 5264 3130 5316 3136
rect 5276 480 5304 3130
rect 6472 480 6500 3334
rect 7668 480 7696 3470
rect 8864 480 8892 4082
rect 10980 3534 11008 318446
rect 16488 318368 16540 318374
rect 16488 318310 16540 318316
rect 12440 5364 12492 5370
rect 12440 5306 12492 5312
rect 10048 3528 10100 3534
rect 10048 3470 10100 3476
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 10060 480 10088 3470
rect 11244 3460 11296 3466
rect 11244 3402 11296 3408
rect 11256 480 11284 3402
rect 12452 480 12480 5306
rect 13636 4072 13688 4078
rect 13636 4014 13688 4020
rect 13648 480 13676 4014
rect 14832 4004 14884 4010
rect 14832 3946 14884 3952
rect 14844 480 14872 3946
rect 16500 3534 16528 318310
rect 17236 35902 17264 534074
rect 17224 35896 17276 35902
rect 17224 35838 17276 35844
rect 19996 8294 20024 536794
rect 20076 495508 20128 495514
rect 20076 495450 20128 495456
rect 20088 309126 20116 495450
rect 21376 465050 21404 667898
rect 21364 465044 21416 465050
rect 21364 464986 21416 464992
rect 24780 458182 24808 699654
rect 31024 610020 31076 610026
rect 31024 609962 31076 609968
rect 28264 532772 28316 532778
rect 28264 532714 28316 532720
rect 24768 458176 24820 458182
rect 24768 458118 24820 458124
rect 20628 318300 20680 318306
rect 20628 318242 20680 318248
rect 20076 309120 20128 309126
rect 20076 309062 20128 309068
rect 19984 8288 20036 8294
rect 19984 8230 20036 8236
rect 18328 3936 18380 3942
rect 18328 3878 18380 3884
rect 16028 3528 16080 3534
rect 16028 3470 16080 3476
rect 16488 3528 16540 3534
rect 16488 3470 16540 3476
rect 16040 480 16068 3470
rect 17224 3120 17276 3126
rect 17224 3062 17276 3068
rect 17236 480 17264 3062
rect 18340 480 18368 3878
rect 20640 3534 20668 318242
rect 21916 318232 21968 318238
rect 21916 318174 21968 318180
rect 21928 3534 21956 318174
rect 24768 318164 24820 318170
rect 24768 318106 24820 318112
rect 22008 5228 22060 5234
rect 22008 5170 22060 5176
rect 19524 3528 19576 3534
rect 19524 3470 19576 3476
rect 20628 3528 20680 3534
rect 20628 3470 20680 3476
rect 20720 3528 20772 3534
rect 20720 3470 20772 3476
rect 21916 3528 21968 3534
rect 21916 3470 21968 3476
rect 19536 480 19564 3470
rect 20732 480 20760 3470
rect 22020 2666 22048 5170
rect 23112 3800 23164 3806
rect 23112 3742 23164 3748
rect 21928 2638 22048 2666
rect 21928 480 21956 2638
rect 23124 480 23152 3742
rect 24780 3534 24808 318106
rect 26148 318096 26200 318102
rect 26148 318038 26200 318044
rect 26160 3534 26188 318038
rect 28276 64870 28304 532714
rect 28356 502376 28408 502382
rect 28356 502318 28408 502324
rect 28368 266354 28396 502318
rect 31036 470558 31064 609962
rect 33784 538280 33836 538286
rect 33784 538222 33836 538228
rect 32404 498228 32456 498234
rect 32404 498170 32456 498176
rect 31024 470552 31076 470558
rect 31024 470494 31076 470500
rect 32416 324290 32444 498170
rect 32404 324284 32456 324290
rect 32404 324226 32456 324232
rect 32404 318028 32456 318034
rect 32404 317970 32456 317976
rect 28356 266348 28408 266354
rect 28356 266290 28408 266296
rect 28264 64864 28316 64870
rect 28264 64806 28316 64812
rect 26700 5160 26752 5166
rect 26700 5102 26752 5108
rect 24308 3528 24360 3534
rect 24308 3470 24360 3476
rect 24768 3528 24820 3534
rect 24768 3470 24820 3476
rect 25504 3528 25556 3534
rect 25504 3470 25556 3476
rect 26148 3528 26200 3534
rect 26148 3470 26200 3476
rect 24320 480 24348 3470
rect 25516 480 25544 3470
rect 26712 480 26740 5102
rect 30288 5092 30340 5098
rect 30288 5034 30340 5040
rect 27896 3800 27948 3806
rect 27896 3742 27948 3748
rect 27908 480 27936 3742
rect 29092 3052 29144 3058
rect 29092 2994 29144 3000
rect 29104 480 29132 2994
rect 30300 480 30328 5034
rect 31484 3732 31536 3738
rect 31484 3674 31536 3680
rect 31496 480 31524 3674
rect 32416 3466 32444 317970
rect 33796 22098 33824 538222
rect 35164 513392 35216 513398
rect 35164 513334 35216 513340
rect 33876 507884 33928 507890
rect 33876 507826 33928 507832
rect 33888 223582 33916 507826
rect 33876 223576 33928 223582
rect 33876 223518 33928 223524
rect 35176 180810 35204 513334
rect 39396 509312 39448 509318
rect 39396 509254 39448 509260
rect 37924 503736 37976 503742
rect 37924 503678 37976 503684
rect 37936 280158 37964 503678
rect 39304 317960 39356 317966
rect 39304 317902 39356 317908
rect 37924 280152 37976 280158
rect 37924 280094 37976 280100
rect 35164 180804 35216 180810
rect 35164 180746 35216 180752
rect 33784 22092 33836 22098
rect 33784 22034 33836 22040
rect 33876 5024 33928 5030
rect 33876 4966 33928 4972
rect 32680 3596 32732 3602
rect 32680 3538 32732 3544
rect 32404 3460 32456 3466
rect 32404 3402 32456 3408
rect 32692 480 32720 3538
rect 33888 480 33916 4966
rect 37372 4956 37424 4962
rect 37372 4898 37424 4904
rect 36176 3664 36228 3670
rect 36176 3606 36228 3612
rect 34980 3528 35032 3534
rect 34980 3470 35032 3476
rect 34992 480 35020 3470
rect 36188 480 36216 3606
rect 37384 480 37412 4898
rect 38568 3188 38620 3194
rect 38568 3130 38620 3136
rect 38580 480 38608 3130
rect 39316 3126 39344 317902
rect 39408 237386 39436 509254
rect 42076 455394 42104 699926
rect 57704 650752 57756 650758
rect 57704 650694 57756 650700
rect 57610 646096 57666 646105
rect 57610 646031 57666 646040
rect 57518 645008 57574 645017
rect 57518 644943 57574 644952
rect 57426 643240 57482 643249
rect 57426 643175 57482 643184
rect 57334 642016 57390 642025
rect 57334 641951 57390 641960
rect 57242 640384 57298 640393
rect 57242 640319 57298 640328
rect 57058 639296 57114 639305
rect 57058 639231 57114 639240
rect 56966 579728 57022 579737
rect 56966 579663 57022 579672
rect 56874 578368 56930 578377
rect 56874 578303 56930 578312
rect 56888 560930 56916 578303
rect 56876 560924 56928 560930
rect 56876 560866 56928 560872
rect 56980 543182 57008 579663
rect 57072 544542 57100 639231
rect 57150 637664 57206 637673
rect 57150 637599 57206 637608
rect 57060 544536 57112 544542
rect 57060 544478 57112 544484
rect 56968 543176 57020 543182
rect 56968 543118 57020 543124
rect 57164 543046 57192 637599
rect 57256 543794 57284 640319
rect 57348 543862 57376 641951
rect 57440 544474 57468 643175
rect 57428 544468 57480 544474
rect 57428 544410 57480 544416
rect 57532 543930 57560 644943
rect 57624 545086 57652 646031
rect 57612 545080 57664 545086
rect 57612 545022 57664 545028
rect 57520 543924 57572 543930
rect 57520 543866 57572 543872
rect 57336 543856 57388 543862
rect 57336 543798 57388 543804
rect 57244 543788 57296 543794
rect 57244 543730 57296 543736
rect 57152 543040 57204 543046
rect 57152 542982 57204 542988
rect 56876 540864 56928 540870
rect 56876 540806 56928 540812
rect 56784 540796 56836 540802
rect 56784 540738 56836 540744
rect 48964 531412 49016 531418
rect 48964 531354 49016 531360
rect 46204 524476 46256 524482
rect 46204 524418 46256 524424
rect 43444 518968 43496 518974
rect 43444 518910 43496 518916
rect 42064 455388 42116 455394
rect 42064 455330 42116 455336
rect 42708 318436 42760 318442
rect 42708 318378 42760 318384
rect 42064 317824 42116 317830
rect 42064 317766 42116 317772
rect 39948 317484 40000 317490
rect 39948 317426 40000 317432
rect 39396 237380 39448 237386
rect 39396 237322 39448 237328
rect 39960 3346 39988 317426
rect 40960 4888 41012 4894
rect 40960 4830 41012 4836
rect 39776 3318 39988 3346
rect 39304 3120 39356 3126
rect 39304 3062 39356 3068
rect 39776 480 39804 3318
rect 40972 480 41000 4830
rect 42076 2922 42104 317766
rect 42720 3466 42748 318378
rect 43456 136610 43484 518910
rect 45468 318572 45520 318578
rect 45468 318514 45520 318520
rect 45480 317830 45508 318514
rect 45468 317824 45520 317830
rect 45468 317766 45520 317772
rect 43444 136604 43496 136610
rect 43444 136546 43496 136552
rect 46216 93838 46244 524418
rect 48136 317552 48188 317558
rect 48136 317494 48188 317500
rect 46204 93832 46256 93838
rect 46204 93774 46256 93780
rect 44548 4820 44600 4826
rect 44548 4762 44600 4768
rect 42156 3460 42208 3466
rect 42156 3402 42208 3408
rect 42708 3460 42760 3466
rect 42708 3402 42760 3408
rect 42800 3460 42852 3466
rect 42800 3402 42852 3408
rect 42064 2916 42116 2922
rect 42064 2858 42116 2864
rect 42168 480 42196 3402
rect 42812 3194 42840 3402
rect 42800 3188 42852 3194
rect 42800 3130 42852 3136
rect 43352 2848 43404 2854
rect 43352 2790 43404 2796
rect 43364 480 43392 2790
rect 44560 480 44588 4762
rect 48148 3194 48176 317494
rect 48976 51066 49004 531354
rect 53104 527196 53156 527202
rect 53104 527138 53156 527144
rect 51724 521756 51776 521762
rect 51724 521698 51776 521704
rect 50344 514820 50396 514826
rect 50344 514762 50396 514768
rect 50356 194546 50384 514762
rect 50436 318708 50488 318714
rect 50436 318650 50488 318656
rect 50344 194540 50396 194546
rect 50344 194482 50396 194488
rect 48964 51060 49016 51066
rect 48964 51002 49016 51008
rect 48228 4208 48280 4214
rect 48228 4150 48280 4156
rect 46940 3188 46992 3194
rect 46940 3130 46992 3136
rect 48136 3188 48188 3194
rect 48136 3130 48188 3136
rect 45744 2916 45796 2922
rect 45744 2858 45796 2864
rect 45756 480 45784 2858
rect 46952 480 46980 3130
rect 48240 2122 48268 4150
rect 50448 3126 50476 318650
rect 50988 317620 51040 317626
rect 50988 317562 51040 317568
rect 51000 3194 51028 317562
rect 51736 151774 51764 521698
rect 51724 151768 51776 151774
rect 51724 151710 51776 151716
rect 53116 109002 53144 527138
rect 56690 490784 56746 490793
rect 56690 490719 56746 490728
rect 56704 489938 56732 490719
rect 56692 489932 56744 489938
rect 56692 489874 56744 489880
rect 56598 488880 56654 488889
rect 56598 488815 56654 488824
rect 56612 484242 56640 488815
rect 56690 486976 56746 486985
rect 56690 486911 56746 486920
rect 56704 485858 56732 486911
rect 56692 485852 56744 485858
rect 56692 485794 56744 485800
rect 56690 485072 56746 485081
rect 56690 485007 56746 485016
rect 56704 484430 56732 485007
rect 56692 484424 56744 484430
rect 56692 484366 56744 484372
rect 56612 484214 56732 484242
rect 56598 483168 56654 483177
rect 56598 483103 56654 483112
rect 56508 480208 56560 480214
rect 56508 480150 56560 480156
rect 56520 479233 56548 480150
rect 56506 479224 56562 479233
rect 56506 479159 56562 479168
rect 56508 477488 56560 477494
rect 56508 477430 56560 477436
rect 56520 477329 56548 477430
rect 56506 477320 56562 477329
rect 56506 477255 56562 477264
rect 56508 476060 56560 476066
rect 56508 476002 56560 476008
rect 56520 475425 56548 476002
rect 56506 475416 56562 475425
rect 56506 475351 56562 475360
rect 56508 474700 56560 474706
rect 56508 474642 56560 474648
rect 56520 473521 56548 474642
rect 56506 473512 56562 473521
rect 56506 473447 56562 473456
rect 56508 471980 56560 471986
rect 56508 471922 56560 471928
rect 56520 471617 56548 471922
rect 56506 471608 56562 471617
rect 56506 471543 56562 471552
rect 56508 470552 56560 470558
rect 56508 470494 56560 470500
rect 56520 469577 56548 470494
rect 56506 469568 56562 469577
rect 56506 469503 56562 469512
rect 56508 467832 56560 467838
rect 56508 467774 56560 467780
rect 56520 467673 56548 467774
rect 56506 467664 56562 467673
rect 56506 467599 56562 467608
rect 56508 466404 56560 466410
rect 56508 466346 56560 466352
rect 56520 465769 56548 466346
rect 56506 465760 56562 465769
rect 56506 465695 56562 465704
rect 56508 465044 56560 465050
rect 56508 464986 56560 464992
rect 56520 463865 56548 464986
rect 56506 463856 56562 463865
rect 56506 463791 56562 463800
rect 56508 462324 56560 462330
rect 56508 462266 56560 462272
rect 56520 461961 56548 462266
rect 56506 461952 56562 461961
rect 56506 461887 56562 461896
rect 56612 460850 56640 483103
rect 56704 481778 56732 484214
rect 56692 481772 56744 481778
rect 56692 481714 56744 481720
rect 56692 481636 56744 481642
rect 56692 481578 56744 481584
rect 56704 481273 56732 481578
rect 56690 481264 56746 481273
rect 56690 481199 56746 481208
rect 56692 481160 56744 481166
rect 56692 481102 56744 481108
rect 56428 460822 56640 460850
rect 56428 459626 56456 460822
rect 56600 460760 56652 460766
rect 56600 460702 56652 460708
rect 56612 459921 56640 460702
rect 56598 459912 56654 459921
rect 56598 459847 56654 459856
rect 56428 459598 56640 459626
rect 56612 458266 56640 459598
rect 56520 458238 56640 458266
rect 56520 457858 56548 458238
rect 56600 458176 56652 458182
rect 56600 458118 56652 458124
rect 56612 458017 56640 458118
rect 56598 458008 56654 458017
rect 56598 457943 56654 457952
rect 56520 457830 56640 457858
rect 56612 456906 56640 457830
rect 56520 456878 56640 456906
rect 56520 454050 56548 456878
rect 56600 456748 56652 456754
rect 56600 456690 56652 456696
rect 56612 456113 56640 456690
rect 56598 456104 56654 456113
rect 56598 456039 56654 456048
rect 56600 455388 56652 455394
rect 56600 455330 56652 455336
rect 56612 454209 56640 455330
rect 56598 454200 56654 454209
rect 56598 454135 56654 454144
rect 56520 454022 56640 454050
rect 56612 452606 56640 454022
rect 56600 452600 56652 452606
rect 56600 452542 56652 452548
rect 56704 396030 56732 481102
rect 56796 442649 56824 540738
rect 56782 442640 56838 442649
rect 56782 442575 56838 442584
rect 56888 436801 56916 540806
rect 56968 540728 57020 540734
rect 56968 540670 57020 540676
rect 56874 436792 56930 436801
rect 56874 436727 56930 436736
rect 56980 431089 57008 540670
rect 57612 539708 57664 539714
rect 57612 539650 57664 539656
rect 57520 539640 57572 539646
rect 57520 539582 57572 539588
rect 57152 539232 57204 539238
rect 57152 539174 57204 539180
rect 57058 492824 57114 492833
rect 57058 492759 57114 492768
rect 56966 431080 57022 431089
rect 56966 431015 57022 431024
rect 56692 396024 56744 396030
rect 56692 395966 56744 395972
rect 57072 380866 57100 492759
rect 57164 382809 57192 539174
rect 57426 539064 57482 539073
rect 57426 538999 57482 539008
rect 57440 538286 57468 538999
rect 57428 538280 57480 538286
rect 57428 538222 57480 538228
rect 57426 537160 57482 537169
rect 57426 537095 57482 537104
rect 57440 536858 57468 537095
rect 57428 536852 57480 536858
rect 57428 536794 57480 536800
rect 57426 535256 57482 535265
rect 57426 535191 57482 535200
rect 57440 534138 57468 535191
rect 57428 534132 57480 534138
rect 57428 534074 57480 534080
rect 57426 533352 57482 533361
rect 57426 533287 57482 533296
rect 57440 532778 57468 533287
rect 57428 532772 57480 532778
rect 57428 532714 57480 532720
rect 57426 531448 57482 531457
rect 57426 531383 57428 531392
rect 57480 531383 57482 531392
rect 57428 531354 57480 531360
rect 57426 529408 57482 529417
rect 57426 529343 57482 529352
rect 57440 528630 57468 529343
rect 57428 528624 57480 528630
rect 57428 528566 57480 528572
rect 57426 527504 57482 527513
rect 57426 527439 57482 527448
rect 57440 527202 57468 527439
rect 57428 527196 57480 527202
rect 57428 527138 57480 527144
rect 57426 525600 57482 525609
rect 57426 525535 57482 525544
rect 57440 524482 57468 525535
rect 57428 524476 57480 524482
rect 57428 524418 57480 524424
rect 57426 523696 57482 523705
rect 57426 523631 57482 523640
rect 57440 523054 57468 523631
rect 57428 523048 57480 523054
rect 57428 522990 57480 522996
rect 57426 521792 57482 521801
rect 57426 521727 57428 521736
rect 57480 521727 57482 521736
rect 57428 521698 57480 521704
rect 57426 519752 57482 519761
rect 57426 519687 57482 519696
rect 57440 518974 57468 519687
rect 57428 518968 57480 518974
rect 57428 518910 57480 518916
rect 57426 517848 57482 517857
rect 57426 517783 57482 517792
rect 57440 517546 57468 517783
rect 57428 517540 57480 517546
rect 57428 517482 57480 517488
rect 57426 515944 57482 515953
rect 57426 515879 57482 515888
rect 57440 514826 57468 515879
rect 57428 514820 57480 514826
rect 57428 514762 57480 514768
rect 57426 514040 57482 514049
rect 57426 513975 57482 513984
rect 57440 513398 57468 513975
rect 57428 513392 57480 513398
rect 57428 513334 57480 513340
rect 57426 512136 57482 512145
rect 57426 512071 57482 512080
rect 57440 512038 57468 512071
rect 57428 512032 57480 512038
rect 57428 511974 57480 511980
rect 57426 510096 57482 510105
rect 57426 510031 57482 510040
rect 57440 509318 57468 510031
rect 57428 509312 57480 509318
rect 57428 509254 57480 509260
rect 57426 508192 57482 508201
rect 57426 508127 57482 508136
rect 57440 507890 57468 508127
rect 57428 507884 57480 507890
rect 57428 507826 57480 507832
rect 57242 506288 57298 506297
rect 57242 506223 57298 506232
rect 57150 382800 57206 382809
rect 57150 382735 57206 382744
rect 57060 380860 57112 380866
rect 57060 380802 57112 380808
rect 56966 371240 57022 371249
rect 56966 371175 57022 371184
rect 56874 361584 56930 361593
rect 56874 361519 56930 361528
rect 56690 359544 56746 359553
rect 56690 359479 56746 359488
rect 56598 357640 56654 357649
rect 56598 357575 56654 357584
rect 56612 330818 56640 357575
rect 56600 330812 56652 330818
rect 56600 330754 56652 330760
rect 56600 330676 56652 330682
rect 56600 330618 56652 330624
rect 56612 325514 56640 330618
rect 56600 325508 56652 325514
rect 56600 325450 56652 325456
rect 56600 325372 56652 325378
rect 56600 325314 56652 325320
rect 56612 320822 56640 325314
rect 56600 320816 56652 320822
rect 56600 320758 56652 320764
rect 55220 318572 55272 318578
rect 55220 318514 55272 318520
rect 55232 317830 55260 318514
rect 55220 317824 55272 317830
rect 55220 317766 55272 317772
rect 56704 311846 56732 359479
rect 56782 355736 56838 355745
rect 56782 355671 56838 355680
rect 56692 311840 56744 311846
rect 56692 311782 56744 311788
rect 56796 299470 56824 355671
rect 56888 330682 56916 361519
rect 56980 330886 57008 371175
rect 57058 365392 57114 365401
rect 57058 365327 57114 365336
rect 56968 330880 57020 330886
rect 56968 330822 57020 330828
rect 56876 330676 56928 330682
rect 56876 330618 56928 330624
rect 57072 330562 57100 365327
rect 57150 351928 57206 351937
rect 57150 351863 57206 351872
rect 56888 330534 57100 330562
rect 56888 325378 56916 330534
rect 57060 330472 57112 330478
rect 57060 330414 57112 330420
rect 56968 329384 57020 329390
rect 56968 329326 57020 329332
rect 56876 325372 56928 325378
rect 56876 325314 56928 325320
rect 56876 325236 56928 325242
rect 56876 325178 56928 325184
rect 56888 320142 56916 325178
rect 56876 320136 56928 320142
rect 56876 320078 56928 320084
rect 56784 299464 56836 299470
rect 56784 299406 56836 299412
rect 56980 124166 57008 329326
rect 57072 329254 57100 330414
rect 57060 329248 57112 329254
rect 57060 329190 57112 329196
rect 57058 328672 57114 328681
rect 57058 328607 57114 328616
rect 56968 124160 57020 124166
rect 56968 124102 57020 124108
rect 53104 108996 53156 109002
rect 53104 108938 53156 108944
rect 57072 88330 57100 328607
rect 57164 276010 57192 351863
rect 57152 276004 57204 276010
rect 57152 275946 57204 275952
rect 57256 252550 57284 506223
rect 57426 504384 57482 504393
rect 57426 504319 57482 504328
rect 57440 503742 57468 504319
rect 57428 503736 57480 503742
rect 57428 503678 57480 503684
rect 57426 502480 57482 502489
rect 57426 502415 57482 502424
rect 57440 502382 57468 502415
rect 57428 502376 57480 502382
rect 57428 502318 57480 502324
rect 57334 500440 57390 500449
rect 57334 500375 57390 500384
rect 57348 295322 57376 500375
rect 57426 498536 57482 498545
rect 57426 498471 57482 498480
rect 57440 498234 57468 498471
rect 57428 498228 57480 498234
rect 57428 498170 57480 498176
rect 57426 496632 57482 496641
rect 57426 496567 57482 496576
rect 57440 495514 57468 496567
rect 57428 495508 57480 495514
rect 57428 495450 57480 495456
rect 57426 494728 57482 494737
rect 57426 494663 57482 494672
rect 57440 338094 57468 494663
rect 57532 380769 57560 539582
rect 57518 380760 57574 380769
rect 57518 380695 57574 380704
rect 57624 378865 57652 539650
rect 57716 448361 57744 650694
rect 57702 448352 57758 448361
rect 57702 448287 57758 448296
rect 57808 440609 57836 700810
rect 57888 700596 57940 700602
rect 57888 700538 57940 700544
rect 57794 440600 57850 440609
rect 57794 440535 57850 440544
rect 57900 429049 57928 700538
rect 58532 700256 58584 700262
rect 58532 700198 58584 700204
rect 58348 700188 58400 700194
rect 58348 700130 58400 700136
rect 58256 556232 58308 556238
rect 58256 556174 58308 556180
rect 57980 540592 58032 540598
rect 57980 540534 58032 540540
rect 57886 429040 57942 429049
rect 57886 428975 57942 428984
rect 57992 415585 58020 540534
rect 58072 540320 58124 540326
rect 58072 540262 58124 540268
rect 57978 415576 58034 415585
rect 57978 415511 58034 415520
rect 58084 400081 58112 540262
rect 58164 540252 58216 540258
rect 58164 540194 58216 540200
rect 58070 400072 58126 400081
rect 58070 400007 58126 400016
rect 58176 392465 58204 540194
rect 58162 392456 58218 392465
rect 58162 392391 58218 392400
rect 58268 386617 58296 556174
rect 58360 452305 58388 700130
rect 58440 700120 58492 700126
rect 58440 700062 58492 700068
rect 58346 452296 58402 452305
rect 58346 452231 58402 452240
rect 58452 450265 58480 700062
rect 58438 450256 58494 450265
rect 58438 450191 58494 450200
rect 58544 446457 58572 700198
rect 58530 446448 58586 446457
rect 58530 446383 58586 446392
rect 58636 444553 58664 700946
rect 58716 700936 58768 700942
rect 58716 700878 58768 700884
rect 58622 444544 58678 444553
rect 58622 444479 58678 444488
rect 58728 438705 58756 700878
rect 58900 700800 58952 700806
rect 58900 700742 58952 700748
rect 58808 700732 58860 700738
rect 58808 700674 58860 700680
rect 58714 438696 58770 438705
rect 58714 438631 58770 438640
rect 58820 434897 58848 700674
rect 58806 434888 58862 434897
rect 58806 434823 58862 434832
rect 58912 432993 58940 700742
rect 58992 700664 59044 700670
rect 58992 700606 59044 700612
rect 58898 432984 58954 432993
rect 58898 432919 58954 432928
rect 59004 427145 59032 700606
rect 59176 700528 59228 700534
rect 59176 700470 59228 700476
rect 59084 700460 59136 700466
rect 59084 700402 59136 700408
rect 58990 427136 59046 427145
rect 58990 427071 59046 427080
rect 59096 423337 59124 700402
rect 59082 423328 59138 423337
rect 59082 423263 59138 423272
rect 59188 421433 59216 700470
rect 59268 700392 59320 700398
rect 59268 700334 59320 700340
rect 59174 421424 59230 421433
rect 59174 421359 59230 421368
rect 59280 417489 59308 700334
rect 59360 700324 59412 700330
rect 59360 700266 59412 700272
rect 59266 417480 59322 417489
rect 59266 417415 59322 417424
rect 59372 409737 59400 700266
rect 72988 700126 73016 703520
rect 89180 700194 89208 703520
rect 105464 703474 105492 703520
rect 105464 703446 105584 703474
rect 89168 700188 89220 700194
rect 89168 700130 89220 700136
rect 72976 700120 73028 700126
rect 72976 700062 73028 700068
rect 105556 698290 105584 703446
rect 137848 701010 137876 703520
rect 137836 701004 137888 701010
rect 137836 700946 137888 700952
rect 137928 701004 137980 701010
rect 137928 700946 137980 700952
rect 137940 699718 137968 700946
rect 154132 700262 154160 703520
rect 154120 700256 154172 700262
rect 154120 700198 154172 700204
rect 137284 699712 137336 699718
rect 137284 699654 137336 699660
rect 137928 699712 137980 699718
rect 137928 699654 137980 699660
rect 104992 698284 105044 698290
rect 104992 698226 105044 698232
rect 105544 698284 105596 698290
rect 105544 698226 105596 698232
rect 77206 697232 77262 697241
rect 77206 697167 77262 697176
rect 96526 697232 96582 697241
rect 96526 697167 96582 697176
rect 77220 697134 77248 697167
rect 96540 697134 96568 697167
rect 70308 697128 70360 697134
rect 70306 697096 70308 697105
rect 77208 697128 77260 697134
rect 70360 697096 70362 697105
rect 89628 697128 89680 697134
rect 77208 697070 77260 697076
rect 89626 697096 89628 697105
rect 96528 697128 96580 697134
rect 89680 697096 89682 697105
rect 70306 697031 70362 697040
rect 96528 697070 96580 697076
rect 89626 697031 89682 697040
rect 105004 688650 105032 698226
rect 115846 697232 115902 697241
rect 115846 697167 115902 697176
rect 135166 697232 135222 697241
rect 135166 697167 135222 697176
rect 115860 697134 115888 697167
rect 135180 697134 135208 697167
rect 108948 697128 109000 697134
rect 108946 697096 108948 697105
rect 115848 697128 115900 697134
rect 109000 697096 109002 697105
rect 128268 697128 128320 697134
rect 115848 697070 115900 697076
rect 128266 697096 128268 697105
rect 135168 697128 135220 697134
rect 128320 697096 128322 697105
rect 108946 697031 109002 697040
rect 135168 697070 135220 697076
rect 128266 697031 128322 697040
rect 104912 688622 105032 688650
rect 104912 683074 104940 688622
rect 104912 683046 105124 683074
rect 105096 673538 105124 683046
rect 104900 673532 104952 673538
rect 104900 673474 104952 673480
rect 105084 673532 105136 673538
rect 105084 673474 105136 673480
rect 104912 663762 104940 673474
rect 104912 663734 105124 663762
rect 105096 650758 105124 663734
rect 129278 652896 129334 652905
rect 129278 652831 129334 652840
rect 133694 652896 133750 652905
rect 133694 652831 133750 652840
rect 129292 652798 129320 652831
rect 133708 652798 133736 652831
rect 129280 652792 129332 652798
rect 129280 652734 129332 652740
rect 133696 652792 133748 652798
rect 133696 652734 133748 652740
rect 135166 650992 135222 651001
rect 135166 650927 135222 650936
rect 120722 650856 120778 650865
rect 120722 650791 120778 650800
rect 105084 650752 105136 650758
rect 89626 650720 89682 650729
rect 59452 650684 59504 650690
rect 105084 650694 105136 650700
rect 106738 650720 106794 650729
rect 89626 650655 89682 650664
rect 106738 650655 106794 650664
rect 59452 650626 59504 650632
rect 59464 425241 59492 650626
rect 89640 650622 89668 650655
rect 106752 650622 106780 650655
rect 89628 650616 89680 650622
rect 96528 650616 96580 650622
rect 89628 650558 89680 650564
rect 96526 650584 96528 650593
rect 106740 650616 106792 650622
rect 96580 650584 96582 650593
rect 115756 650616 115808 650622
rect 106740 650558 106792 650564
rect 115754 650584 115756 650593
rect 115808 650584 115810 650593
rect 96526 650519 96582 650528
rect 115754 650519 115810 650528
rect 115938 650584 115994 650593
rect 120736 650554 120764 650791
rect 135180 650593 135208 650927
rect 135166 650584 135222 650593
rect 115938 650519 115940 650528
rect 115992 650519 115994 650528
rect 120724 650548 120776 650554
rect 115940 650490 115992 650496
rect 135166 650519 135222 650528
rect 120724 650490 120776 650496
rect 67546 558920 67602 558929
rect 62028 558884 62080 558890
rect 67546 558855 67602 558864
rect 68926 558920 68982 558929
rect 68926 558855 68982 558864
rect 70306 558920 70362 558929
rect 70306 558855 70362 558864
rect 71686 558920 71742 558929
rect 71686 558855 71742 558864
rect 72606 558920 72662 558929
rect 72606 558855 72662 558864
rect 73066 558920 73122 558929
rect 73066 558855 73122 558864
rect 73802 558920 73858 558929
rect 73802 558855 73858 558864
rect 74262 558920 74318 558929
rect 74262 558855 74318 558864
rect 74998 558920 75054 558929
rect 74998 558855 75054 558864
rect 76010 558920 76066 558929
rect 76010 558855 76066 558864
rect 76838 558920 76894 558929
rect 76838 558855 76894 558864
rect 77390 558920 77446 558929
rect 77390 558855 77446 558864
rect 78494 558920 78550 558929
rect 78494 558855 78550 558864
rect 79414 558920 79470 558929
rect 79414 558855 79470 558864
rect 79966 558920 80022 558929
rect 79966 558855 80022 558864
rect 80794 558920 80850 558929
rect 80794 558855 80850 558864
rect 81254 558920 81310 558929
rect 81254 558855 81310 558864
rect 81898 558920 81954 558929
rect 81898 558855 81954 558864
rect 82726 558920 82782 558929
rect 82726 558855 82782 558864
rect 83830 558920 83886 558929
rect 83830 558855 83886 558864
rect 84198 558920 84254 558929
rect 84198 558855 84254 558864
rect 85486 558920 85542 558929
rect 85486 558855 85542 558864
rect 86406 558920 86462 558929
rect 86406 558855 86462 558864
rect 86866 558920 86922 558929
rect 86866 558855 86922 558864
rect 87878 558920 87934 558929
rect 87878 558855 87934 558864
rect 88246 558920 88302 558929
rect 88246 558855 88302 558864
rect 88890 558920 88946 558929
rect 88890 558855 88946 558864
rect 89626 558920 89682 558929
rect 89626 558855 89682 558864
rect 89810 558920 89866 558929
rect 89810 558855 89866 558864
rect 91006 558920 91062 558929
rect 91006 558855 91062 558864
rect 92478 558920 92534 558929
rect 92478 558855 92534 558864
rect 93674 558920 93730 558929
rect 93674 558855 93730 558864
rect 94870 558920 94926 558929
rect 94870 558855 94926 558864
rect 95146 558920 95202 558929
rect 95146 558855 95202 558864
rect 95790 558920 95846 558929
rect 95790 558855 95846 558864
rect 96526 558920 96582 558929
rect 96526 558855 96582 558864
rect 96986 558920 97042 558929
rect 96986 558855 97042 558864
rect 97814 558920 97870 558929
rect 97814 558855 97870 558864
rect 98090 558920 98146 558929
rect 98090 558855 98146 558864
rect 99286 558920 99342 558929
rect 99286 558855 99342 558864
rect 99562 558920 99618 558929
rect 99562 558855 99618 558864
rect 100390 558920 100446 558929
rect 100390 558855 100446 558864
rect 102046 558920 102102 558929
rect 102046 558855 102102 558864
rect 103426 558920 103482 558929
rect 103426 558855 103482 558864
rect 104806 558920 104862 558929
rect 104806 558855 104862 558864
rect 105542 558920 105598 558929
rect 105542 558855 105598 558864
rect 106186 558920 106242 558929
rect 106186 558855 106242 558864
rect 107474 558920 107530 558929
rect 107474 558855 107530 558864
rect 108486 558920 108542 558929
rect 108486 558855 108542 558864
rect 110326 558920 110382 558929
rect 110326 558855 110382 558864
rect 62028 558826 62080 558832
rect 62040 543590 62068 558826
rect 67456 558816 67508 558822
rect 67456 558758 67508 558764
rect 66168 557796 66220 557802
rect 66168 557738 66220 557744
rect 63408 557660 63460 557666
rect 63408 557602 63460 557608
rect 61016 543584 61068 543590
rect 61016 543526 61068 543532
rect 62028 543584 62080 543590
rect 62028 543526 62080 543532
rect 59912 540660 59964 540666
rect 59912 540602 59964 540608
rect 59820 540524 59872 540530
rect 59820 540466 59872 540472
rect 59728 540456 59780 540462
rect 59728 540398 59780 540404
rect 59636 540388 59688 540394
rect 59636 540330 59688 540336
rect 59544 539776 59596 539782
rect 59544 539718 59596 539724
rect 59450 425232 59506 425241
rect 59450 425167 59506 425176
rect 59452 419484 59504 419490
rect 59452 419426 59504 419432
rect 59464 419393 59492 419426
rect 59450 419384 59506 419393
rect 59450 419319 59506 419328
rect 59358 409728 59414 409737
rect 59358 409663 59414 409672
rect 58254 386608 58310 386617
rect 58254 386543 58310 386552
rect 59556 384713 59584 539718
rect 59648 390425 59676 540330
rect 59740 396273 59768 540398
rect 59832 413681 59860 540466
rect 59924 419490 59952 540602
rect 61028 539988 61056 543526
rect 63420 540002 63448 557602
rect 66180 542570 66208 557738
rect 65156 542564 65208 542570
rect 65156 542506 65208 542512
rect 66168 542564 66220 542570
rect 66168 542506 66220 542512
rect 63066 539974 63448 540002
rect 65168 539988 65196 542506
rect 67468 540002 67496 558758
rect 67560 543114 67588 558855
rect 67548 543108 67600 543114
rect 67548 543050 67600 543056
rect 68940 542450 68968 558855
rect 70214 558648 70270 558657
rect 70214 558583 70270 558592
rect 70228 543590 70256 558583
rect 70216 543584 70268 543590
rect 70216 543526 70268 543532
rect 70320 542910 70348 558855
rect 71700 543726 71728 558855
rect 72620 558346 72648 558855
rect 72608 558340 72660 558346
rect 72608 558282 72660 558288
rect 73080 544066 73108 558855
rect 73816 558142 73844 558855
rect 73804 558136 73856 558142
rect 73804 558078 73856 558084
rect 74276 558006 74304 558855
rect 74264 558000 74316 558006
rect 74264 557942 74316 557948
rect 75012 557734 75040 558855
rect 76024 558686 76052 558855
rect 76012 558680 76064 558686
rect 76012 558622 76064 558628
rect 75826 558240 75882 558249
rect 76852 558210 76880 558855
rect 77404 558754 77432 558855
rect 77392 558748 77444 558754
rect 77392 558690 77444 558696
rect 78508 558482 78536 558855
rect 78496 558476 78548 558482
rect 78496 558418 78548 558424
rect 78586 558376 78642 558385
rect 78586 558311 78642 558320
rect 75826 558175 75882 558184
rect 76840 558204 76892 558210
rect 75000 557728 75052 557734
rect 75000 557670 75052 557676
rect 73068 544060 73120 544066
rect 73068 544002 73120 544008
rect 75840 543726 75868 558175
rect 76840 558146 76892 558152
rect 77576 545760 77628 545766
rect 77576 545702 77628 545708
rect 71688 543720 71740 543726
rect 71688 543662 71740 543668
rect 75460 543720 75512 543726
rect 75460 543662 75512 543668
rect 75828 543720 75880 543726
rect 75828 543662 75880 543668
rect 71320 543584 71372 543590
rect 71320 543526 71372 543532
rect 70308 542904 70360 542910
rect 70308 542846 70360 542852
rect 68940 542422 69060 542450
rect 67206 539974 67496 540002
rect 69032 540002 69060 542422
rect 69032 539974 69322 540002
rect 71332 539988 71360 543526
rect 73436 542904 73488 542910
rect 73436 542846 73488 542852
rect 73448 539988 73476 542846
rect 75472 539988 75500 543662
rect 77588 539988 77616 545702
rect 78600 543658 78628 558311
rect 79428 558074 79456 558855
rect 79598 558648 79654 558657
rect 79598 558583 79654 558592
rect 79612 558550 79640 558583
rect 79600 558544 79652 558550
rect 79600 558486 79652 558492
rect 79416 558068 79468 558074
rect 79416 558010 79468 558016
rect 79980 557870 80008 558855
rect 80808 558414 80836 558855
rect 80796 558408 80848 558414
rect 80796 558350 80848 558356
rect 81268 558278 81296 558855
rect 81912 558346 81940 558855
rect 81900 558340 81952 558346
rect 81900 558282 81952 558288
rect 81256 558272 81308 558278
rect 81256 558214 81308 558220
rect 79968 557864 80020 557870
rect 79968 557806 80020 557812
rect 80702 545184 80758 545193
rect 80702 545119 80758 545128
rect 80716 544921 80744 545119
rect 80702 544912 80758 544921
rect 80702 544847 80758 544856
rect 81716 544400 81768 544406
rect 81716 544342 81768 544348
rect 78588 543652 78640 543658
rect 78588 543594 78640 543600
rect 79692 543176 79744 543182
rect 79692 543118 79744 543124
rect 79704 539988 79732 543118
rect 81728 539988 81756 544342
rect 82740 543590 82768 558855
rect 82818 558648 82874 558657
rect 82818 558583 82874 558592
rect 82832 558142 82860 558583
rect 83844 558142 83872 558855
rect 84212 558634 84240 558855
rect 84292 558680 84344 558686
rect 84212 558628 84292 558634
rect 84212 558622 84344 558628
rect 85210 558648 85266 558657
rect 84212 558606 84332 558622
rect 82820 558136 82872 558142
rect 82820 558078 82872 558084
rect 83832 558136 83884 558142
rect 83832 558078 83884 558084
rect 82832 557938 82860 558078
rect 82820 557932 82872 557938
rect 82820 557874 82872 557880
rect 84212 557734 84240 558606
rect 85210 558583 85212 558592
rect 85264 558583 85266 558592
rect 85212 558554 85264 558560
rect 84200 557728 84252 557734
rect 84200 557670 84252 557676
rect 83830 544368 83886 544377
rect 83830 544303 83886 544312
rect 82728 543584 82780 543590
rect 82728 543526 82780 543532
rect 83844 539988 83872 544303
rect 85500 544134 85528 558855
rect 86420 558754 86448 558855
rect 86408 558748 86460 558754
rect 86408 558690 86460 558696
rect 86774 558648 86830 558657
rect 86774 558583 86830 558592
rect 85580 545352 85632 545358
rect 85578 545320 85580 545329
rect 85632 545320 85634 545329
rect 85578 545255 85634 545264
rect 85854 544504 85910 544513
rect 85854 544439 85910 544448
rect 85488 544128 85540 544134
rect 85488 544070 85540 544076
rect 85868 539988 85896 544439
rect 86788 544202 86816 558583
rect 86880 544338 86908 558855
rect 87892 558482 87920 558855
rect 87880 558476 87932 558482
rect 87880 558418 87932 558424
rect 87970 544640 88026 544649
rect 87970 544575 88026 544584
rect 86868 544332 86920 544338
rect 86868 544274 86920 544280
rect 86776 544196 86828 544202
rect 86776 544138 86828 544144
rect 87984 539988 88012 544575
rect 88260 544270 88288 558855
rect 88904 558550 88932 558855
rect 88892 558544 88944 558550
rect 88892 558486 88944 558492
rect 89640 545018 89668 558855
rect 89824 558414 89852 558855
rect 89812 558408 89864 558414
rect 89812 558350 89864 558356
rect 89628 545012 89680 545018
rect 89628 544954 89680 544960
rect 91020 544814 91048 558855
rect 91098 558648 91154 558657
rect 91098 558583 91154 558592
rect 91112 558346 91140 558583
rect 92386 558376 92442 558385
rect 91100 558340 91152 558346
rect 92492 558346 92520 558855
rect 93308 558680 93360 558686
rect 93306 558648 93308 558657
rect 93360 558648 93362 558657
rect 93306 558583 93362 558592
rect 92386 558311 92442 558320
rect 92480 558340 92532 558346
rect 91100 558282 91152 558288
rect 91112 557598 91140 558282
rect 91100 557592 91152 557598
rect 91100 557534 91152 557540
rect 92400 544950 92428 558311
rect 92480 558282 92532 558288
rect 92492 557938 92520 558282
rect 92480 557932 92532 557938
rect 92480 557874 92532 557880
rect 93320 557734 93348 558583
rect 93308 557728 93360 557734
rect 93308 557670 93360 557676
rect 92388 544944 92440 544950
rect 92388 544886 92440 544892
rect 91008 544808 91060 544814
rect 91008 544750 91060 544756
rect 92110 544776 92166 544785
rect 92110 544711 92166 544720
rect 89996 544604 90048 544610
rect 89996 544546 90048 544552
rect 88248 544264 88300 544270
rect 88248 544206 88300 544212
rect 90008 539988 90036 544546
rect 92124 539988 92152 544711
rect 93688 543250 93716 558855
rect 93766 558648 93822 558657
rect 94884 558618 94912 558855
rect 93766 558583 93822 558592
rect 94872 558612 94924 558618
rect 93780 557938 93808 558583
rect 94872 558554 94924 558560
rect 93768 557932 93820 557938
rect 93768 557874 93820 557880
rect 95056 545352 95108 545358
rect 95054 545320 95056 545329
rect 95108 545320 95110 545329
rect 95054 545255 95110 545264
rect 94136 544672 94188 544678
rect 94136 544614 94188 544620
rect 93676 543244 93728 543250
rect 93676 543186 93728 543192
rect 94148 539988 94176 544614
rect 95160 543182 95188 558855
rect 95804 558754 95832 558855
rect 95792 558748 95844 558754
rect 95792 558690 95844 558696
rect 96252 544876 96304 544882
rect 96252 544818 96304 544824
rect 95148 543176 95200 543182
rect 95148 543118 95200 543124
rect 96264 539988 96292 544818
rect 96540 544746 96568 558855
rect 97000 558482 97028 558855
rect 97828 558686 97856 558855
rect 97816 558680 97868 558686
rect 97816 558622 97868 558628
rect 98104 558550 98132 558855
rect 98092 558544 98144 558550
rect 98092 558486 98144 558492
rect 96988 558476 97040 558482
rect 96988 558418 97040 558424
rect 97998 558376 98054 558385
rect 98104 558346 98132 558486
rect 97998 558311 98000 558320
rect 98052 558311 98054 558320
rect 98092 558340 98144 558346
rect 98000 558282 98052 558288
rect 98092 558282 98144 558288
rect 96618 545320 96674 545329
rect 96618 545255 96620 545264
rect 96672 545255 96674 545264
rect 96620 545226 96672 545232
rect 96528 544740 96580 544746
rect 96528 544682 96580 544688
rect 99300 543114 99328 558855
rect 99576 558550 99604 558855
rect 100022 558648 100078 558657
rect 100022 558583 100078 558592
rect 99564 558544 99616 558550
rect 99564 558486 99616 558492
rect 99576 558414 99604 558486
rect 99564 558408 99616 558414
rect 99564 558350 99616 558356
rect 99840 557728 99892 557734
rect 99840 557670 99892 557676
rect 99852 557530 99880 557670
rect 100036 557598 100064 558583
rect 100404 558346 100432 558855
rect 101954 558648 102010 558657
rect 101954 558583 102010 558592
rect 101968 558414 101996 558583
rect 100576 558408 100628 558414
rect 101956 558408 102008 558414
rect 100576 558350 100628 558356
rect 101402 558376 101458 558385
rect 100392 558340 100444 558346
rect 100392 558282 100444 558288
rect 100024 557592 100076 557598
rect 100024 557534 100076 557540
rect 99840 557524 99892 557530
rect 99840 557466 99892 557472
rect 98368 543108 98420 543114
rect 98368 543050 98420 543056
rect 99288 543108 99340 543114
rect 99288 543050 99340 543056
rect 98380 539988 98408 543050
rect 100036 542842 100064 557534
rect 100588 557530 100616 558350
rect 101956 558350 102008 558356
rect 101402 558311 101458 558320
rect 100576 557524 100628 557530
rect 100576 557466 100628 557472
rect 100392 543040 100444 543046
rect 100392 542982 100444 542988
rect 100024 542836 100076 542842
rect 100024 542778 100076 542784
rect 100404 539988 100432 542982
rect 101416 542434 101444 558311
rect 102060 543046 102088 558855
rect 102782 558648 102838 558657
rect 102782 558583 102838 558592
rect 102796 557598 102824 558583
rect 102876 557864 102928 557870
rect 102876 557806 102928 557812
rect 102784 557592 102836 557598
rect 102784 557534 102836 557540
rect 102508 544536 102560 544542
rect 102508 544478 102560 544484
rect 102048 543040 102100 543046
rect 102048 542982 102100 542988
rect 101404 542428 101456 542434
rect 101404 542370 101456 542376
rect 102520 539988 102548 544478
rect 102796 542774 102824 557534
rect 102888 543998 102916 557806
rect 103440 544542 103468 558855
rect 103886 558648 103942 558657
rect 104820 558618 104848 558855
rect 105556 558754 105584 558855
rect 105544 558748 105596 558754
rect 105544 558690 105596 558696
rect 103886 558583 103888 558592
rect 103940 558583 103942 558592
rect 104164 558612 104216 558618
rect 103888 558554 103940 558560
rect 104164 558554 104216 558560
rect 104808 558612 104860 558618
rect 104808 558554 104860 558560
rect 103428 544536 103480 544542
rect 103428 544478 103480 544484
rect 102876 543992 102928 543998
rect 102876 543934 102928 543940
rect 104176 542978 104204 558554
rect 104808 545284 104860 545290
rect 104808 545226 104860 545232
rect 104820 545193 104848 545226
rect 104806 545184 104862 545193
rect 104806 545119 104862 545128
rect 104532 543788 104584 543794
rect 104532 543730 104584 543736
rect 104164 542972 104216 542978
rect 104164 542914 104216 542920
rect 102784 542768 102836 542774
rect 102784 542710 102836 542716
rect 104544 539988 104572 543730
rect 105556 542910 105584 558690
rect 106200 543017 106228 558855
rect 106922 558648 106978 558657
rect 106922 558583 106978 558592
rect 106936 558482 106964 558583
rect 106924 558476 106976 558482
rect 106924 558418 106976 558424
rect 106648 543856 106700 543862
rect 106648 543798 106700 543804
rect 106186 543008 106242 543017
rect 106186 542943 106242 542952
rect 105544 542904 105596 542910
rect 105544 542846 105596 542852
rect 106660 539988 106688 543798
rect 106936 542502 106964 558418
rect 107488 557734 107516 558855
rect 107750 558648 107806 558657
rect 107750 558583 107806 558592
rect 108302 558648 108358 558657
rect 108302 558583 108358 558592
rect 107476 557728 107528 557734
rect 107476 557670 107528 557676
rect 107764 557598 107792 558583
rect 108316 558550 108344 558583
rect 108304 558544 108356 558550
rect 108304 558486 108356 558492
rect 107752 557592 107804 557598
rect 107752 557534 107804 557540
rect 108316 542638 108344 558486
rect 108500 558482 108528 558855
rect 108488 558476 108540 558482
rect 108488 558418 108540 558424
rect 108488 557592 108540 557598
rect 108488 557534 108540 557540
rect 108304 542632 108356 542638
rect 108304 542574 108356 542580
rect 108500 542570 108528 557534
rect 110340 544474 110368 558855
rect 125508 558748 125560 558754
rect 125508 558690 125560 558696
rect 121368 557864 121420 557870
rect 121368 557806 121420 557812
rect 115938 545456 115994 545465
rect 115938 545391 115940 545400
rect 115992 545391 115994 545400
rect 115940 545362 115992 545368
rect 112812 545080 112864 545086
rect 112812 545022 112864 545028
rect 114928 545080 114980 545086
rect 114928 545022 114980 545028
rect 108672 544468 108724 544474
rect 108672 544410 108724 544416
rect 110328 544468 110380 544474
rect 110328 544410 110380 544416
rect 108488 542564 108540 542570
rect 108488 542506 108540 542512
rect 106924 542496 106976 542502
rect 106924 542438 106976 542444
rect 108684 539988 108712 544410
rect 110788 543924 110840 543930
rect 110788 543866 110840 543872
rect 110800 539988 110828 543866
rect 112824 539988 112852 545022
rect 114940 539988 114968 545022
rect 119068 543380 119120 543386
rect 119068 543322 119120 543328
rect 117044 543312 117096 543318
rect 117044 543254 117096 543260
rect 117056 539988 117084 543254
rect 119080 539988 119108 543322
rect 121380 540002 121408 557806
rect 125416 545420 125468 545426
rect 125416 545362 125468 545368
rect 125428 545193 125456 545362
rect 125414 545184 125470 545193
rect 125414 545119 125470 545128
rect 123208 543448 123260 543454
rect 123208 543390 123260 543396
rect 121210 539974 121408 540002
rect 123220 539988 123248 543390
rect 125520 540002 125548 558690
rect 133144 558680 133196 558686
rect 133144 558622 133196 558628
rect 127256 557932 127308 557938
rect 127256 557874 127308 557880
rect 129648 557932 129700 557938
rect 129648 557874 129700 557880
rect 127268 557598 127296 557874
rect 127256 557592 127308 557598
rect 127256 557534 127308 557540
rect 127348 543516 127400 543522
rect 127348 543458 127400 543464
rect 125350 539974 125548 540002
rect 127360 539988 127388 543458
rect 129660 540002 129688 557874
rect 131764 557592 131816 557598
rect 131764 557534 131816 557540
rect 131488 542836 131540 542842
rect 131488 542778 131540 542784
rect 129490 539974 129688 540002
rect 131500 539988 131528 542778
rect 131776 542706 131804 557534
rect 133156 542842 133184 558622
rect 135904 558000 135956 558006
rect 135904 557942 135956 557948
rect 135258 545456 135314 545465
rect 135258 545391 135260 545400
rect 135312 545391 135314 545400
rect 135260 545362 135312 545368
rect 133144 542836 133196 542842
rect 133144 542778 133196 542784
rect 135720 542768 135772 542774
rect 135720 542710 135772 542716
rect 131764 542700 131816 542706
rect 131764 542642 131816 542648
rect 133604 542428 133656 542434
rect 133604 542370 133656 542376
rect 133616 539988 133644 542370
rect 135732 539988 135760 542710
rect 135916 542434 135944 557942
rect 135904 542428 135956 542434
rect 135904 542370 135956 542376
rect 137296 540870 137324 699654
rect 154486 697232 154542 697241
rect 154486 697167 154542 697176
rect 154500 697134 154528 697167
rect 147588 697128 147640 697134
rect 147586 697096 147588 697105
rect 154488 697128 154540 697134
rect 147640 697096 147642 697105
rect 166908 697128 166960 697134
rect 154488 697070 154540 697076
rect 166906 697096 166908 697105
rect 166960 697096 166962 697105
rect 147586 697031 147642 697040
rect 166906 697031 166962 697040
rect 170324 695502 170352 703520
rect 202800 700942 202828 703520
rect 202788 700936 202840 700942
rect 202788 700878 202840 700884
rect 218992 700874 219020 703520
rect 235184 701010 235212 703520
rect 235172 701004 235224 701010
rect 235172 700946 235224 700952
rect 218980 700868 219032 700874
rect 218980 700810 219032 700816
rect 267660 700806 267688 703520
rect 267648 700800 267700 700806
rect 267648 700742 267700 700748
rect 283852 700738 283880 703520
rect 283840 700732 283892 700738
rect 283840 700674 283892 700680
rect 173806 697232 173862 697241
rect 173806 697167 173862 697176
rect 193126 697232 193182 697241
rect 193126 697167 193182 697176
rect 212446 697232 212502 697241
rect 212446 697167 212502 697176
rect 231766 697232 231822 697241
rect 231766 697167 231822 697176
rect 251086 697232 251142 697241
rect 251086 697167 251142 697176
rect 270406 697232 270462 697241
rect 270406 697167 270462 697176
rect 289726 697232 289782 697241
rect 289726 697167 289782 697176
rect 173820 697134 173848 697167
rect 193140 697134 193168 697167
rect 212460 697134 212488 697167
rect 231780 697134 231808 697167
rect 251100 697134 251128 697167
rect 270420 697134 270448 697167
rect 289740 697134 289768 697167
rect 173808 697128 173860 697134
rect 186228 697128 186280 697134
rect 173808 697070 173860 697076
rect 186226 697096 186228 697105
rect 193128 697128 193180 697134
rect 186280 697096 186282 697105
rect 205548 697128 205600 697134
rect 193128 697070 193180 697076
rect 205546 697096 205548 697105
rect 212448 697128 212500 697134
rect 205600 697096 205602 697105
rect 186226 697031 186282 697040
rect 224868 697128 224920 697134
rect 212448 697070 212500 697076
rect 224866 697096 224868 697105
rect 231768 697128 231820 697134
rect 224920 697096 224922 697105
rect 205546 697031 205602 697040
rect 244188 697128 244240 697134
rect 231768 697070 231820 697076
rect 244186 697096 244188 697105
rect 251088 697128 251140 697134
rect 244240 697096 244242 697105
rect 224866 697031 224922 697040
rect 263508 697128 263560 697134
rect 251088 697070 251140 697076
rect 263506 697096 263508 697105
rect 270408 697128 270460 697134
rect 263560 697096 263562 697105
rect 244186 697031 244242 697040
rect 282828 697128 282880 697134
rect 270408 697070 270460 697076
rect 282826 697096 282828 697105
rect 289728 697128 289780 697134
rect 282880 697096 282882 697105
rect 263506 697031 263562 697040
rect 289728 697070 289780 697076
rect 282826 697031 282882 697040
rect 170128 695496 170180 695502
rect 170128 695438 170180 695444
rect 170312 695496 170364 695502
rect 170312 695438 170364 695444
rect 166906 686352 166962 686361
rect 167090 686352 167146 686361
rect 166962 686310 167090 686338
rect 166906 686287 166962 686296
rect 167090 686287 167146 686296
rect 154578 686216 154634 686225
rect 154578 686151 154580 686160
rect 154632 686151 154634 686160
rect 162216 686180 162268 686186
rect 154580 686122 154632 686128
rect 162216 686122 162268 686128
rect 162228 685953 162256 686122
rect 170140 685982 170168 695438
rect 188342 686488 188398 686497
rect 188342 686423 188398 686432
rect 173898 686352 173954 686361
rect 173898 686287 173900 686296
rect 173952 686287 173954 686296
rect 178776 686316 178828 686322
rect 173900 686258 173952 686264
rect 178776 686258 178828 686264
rect 178788 686225 178816 686258
rect 188356 686225 188384 686423
rect 178774 686216 178830 686225
rect 178774 686151 178830 686160
rect 188342 686216 188398 686225
rect 188342 686151 188398 686160
rect 289818 686216 289874 686225
rect 289818 686151 289820 686160
rect 289872 686151 289874 686160
rect 294512 686180 294564 686186
rect 289820 686122 289872 686128
rect 294512 686122 294564 686128
rect 169852 685976 169904 685982
rect 162214 685944 162270 685953
rect 169852 685918 169904 685924
rect 170128 685976 170180 685982
rect 294524 685953 294552 686122
rect 170128 685918 170180 685924
rect 294510 685944 294566 685953
rect 162214 685879 162270 685888
rect 169864 684486 169892 685918
rect 300136 685914 300164 703520
rect 332520 700670 332548 703520
rect 332508 700664 332560 700670
rect 332508 700606 332560 700612
rect 348804 700602 348832 703520
rect 364996 703474 365024 703520
rect 364996 703446 365116 703474
rect 348792 700596 348844 700602
rect 348792 700538 348844 700544
rect 365088 698290 365116 703446
rect 397472 700534 397500 703520
rect 397460 700528 397512 700534
rect 397460 700470 397512 700476
rect 413664 700466 413692 703520
rect 429856 703474 429884 703520
rect 429856 703446 429976 703474
rect 413652 700460 413704 700466
rect 413652 700402 413704 700408
rect 364432 698284 364484 698290
rect 364432 698226 364484 698232
rect 365076 698284 365128 698290
rect 365076 698226 365128 698232
rect 309046 697232 309102 697241
rect 309046 697167 309102 697176
rect 328366 697232 328422 697241
rect 328366 697167 328422 697176
rect 309060 697134 309088 697167
rect 328380 697134 328408 697167
rect 302148 697128 302200 697134
rect 302146 697096 302148 697105
rect 309048 697128 309100 697134
rect 302200 697096 302202 697105
rect 321468 697128 321520 697134
rect 309048 697070 309100 697076
rect 321466 697096 321468 697105
rect 328368 697128 328420 697134
rect 321520 697096 321522 697105
rect 302146 697031 302202 697040
rect 328368 697070 328420 697076
rect 321466 697031 321522 697040
rect 364444 688650 364472 698226
rect 429948 692850 429976 703446
rect 429200 692844 429252 692850
rect 429200 692786 429252 692792
rect 429936 692844 429988 692850
rect 429936 692786 429988 692792
rect 364352 688622 364472 688650
rect 364352 688514 364380 688622
rect 364352 688486 364472 688514
rect 360106 686352 360162 686361
rect 360290 686352 360346 686361
rect 360162 686310 360290 686338
rect 360106 686287 360162 686296
rect 360290 686287 360346 686296
rect 347778 686216 347834 686225
rect 347778 686151 347780 686160
rect 347832 686151 347834 686160
rect 355416 686180 355468 686186
rect 347780 686122 347832 686128
rect 355416 686122 355468 686128
rect 355428 685953 355456 686122
rect 355414 685944 355470 685953
rect 294510 685879 294566 685888
rect 299572 685908 299624 685914
rect 299572 685850 299624 685856
rect 300124 685908 300176 685914
rect 355414 685879 355470 685888
rect 300124 685850 300176 685856
rect 299584 684486 299612 685850
rect 169852 684480 169904 684486
rect 169852 684422 169904 684428
rect 170220 684480 170272 684486
rect 170220 684422 170272 684428
rect 299572 684480 299624 684486
rect 299572 684422 299624 684428
rect 299664 684480 299716 684486
rect 299664 684422 299716 684428
rect 166998 673976 167054 673985
rect 166998 673911 167054 673920
rect 154578 673840 154634 673849
rect 154578 673775 154580 673784
rect 154632 673775 154634 673784
rect 162216 673804 162268 673810
rect 154580 673746 154632 673752
rect 162216 673746 162268 673752
rect 162228 673577 162256 673746
rect 162214 673568 162270 673577
rect 162214 673503 162270 673512
rect 166906 673568 166962 673577
rect 167012 673554 167040 673911
rect 166962 673526 167040 673554
rect 166906 673503 166962 673512
rect 170232 661774 170260 684422
rect 299676 679046 299704 684422
rect 299664 679040 299716 679046
rect 299664 678982 299716 678988
rect 299664 678904 299716 678910
rect 299664 678846 299716 678852
rect 188342 674112 188398 674121
rect 188342 674047 188398 674056
rect 173898 673976 173954 673985
rect 173898 673911 173900 673920
rect 173952 673911 173954 673920
rect 178776 673940 178828 673946
rect 173900 673882 173952 673888
rect 178776 673882 178828 673888
rect 178788 673849 178816 673882
rect 188356 673849 188384 674047
rect 178774 673840 178830 673849
rect 178774 673775 178830 673784
rect 188342 673840 188398 673849
rect 188342 673775 188398 673784
rect 289818 673840 289874 673849
rect 289818 673775 289820 673784
rect 289872 673775 289874 673784
rect 292672 673804 292724 673810
rect 289820 673746 289872 673752
rect 292672 673746 292724 673752
rect 292684 673577 292712 673746
rect 292670 673568 292726 673577
rect 292670 673503 292726 673512
rect 299676 666602 299704 678846
rect 360106 673976 360162 673985
rect 360290 673976 360346 673985
rect 360162 673934 360290 673962
rect 360106 673911 360162 673920
rect 360290 673911 360346 673920
rect 347778 673840 347834 673849
rect 347778 673775 347780 673784
rect 347832 673775 347834 673784
rect 355416 673804 355468 673810
rect 347780 673746 347832 673752
rect 355416 673746 355468 673752
rect 355428 673577 355456 673746
rect 355414 673568 355470 673577
rect 355414 673503 355470 673512
rect 364444 669458 364472 688486
rect 379518 686488 379574 686497
rect 379518 686423 379574 686432
rect 367098 686352 367154 686361
rect 367098 686287 367100 686296
rect 367152 686287 367154 686296
rect 371976 686316 372028 686322
rect 367100 686258 367152 686264
rect 371976 686258 372028 686264
rect 371988 686225 372016 686258
rect 379532 686225 379560 686423
rect 371974 686216 372030 686225
rect 371974 686151 372030 686160
rect 379518 686216 379574 686225
rect 379518 686151 379574 686160
rect 427542 686216 427598 686225
rect 427726 686216 427782 686225
rect 427598 686174 427726 686202
rect 427542 686151 427598 686160
rect 427726 686151 427782 686160
rect 379518 674112 379574 674121
rect 379518 674047 379574 674056
rect 367098 673976 367154 673985
rect 367098 673911 367100 673920
rect 367152 673911 367154 673920
rect 371976 673940 372028 673946
rect 367100 673882 367152 673888
rect 371976 673882 372028 673888
rect 371988 673849 372016 673882
rect 379532 673849 379560 674047
rect 371974 673840 372030 673849
rect 371974 673775 372030 673784
rect 379518 673840 379574 673849
rect 379518 673775 379574 673784
rect 429212 673470 429240 692786
rect 441526 686488 441582 686497
rect 441526 686423 441582 686432
rect 441540 686225 441568 686423
rect 441526 686216 441582 686225
rect 441526 686151 441582 686160
rect 429200 673464 429252 673470
rect 429200 673406 429252 673412
rect 429476 673464 429528 673470
rect 429476 673406 429528 673412
rect 364432 669452 364484 669458
rect 364432 669394 364484 669400
rect 364432 669316 364484 669322
rect 364432 669258 364484 669264
rect 299664 666596 299716 666602
rect 299664 666538 299716 666544
rect 299940 666596 299992 666602
rect 299940 666538 299992 666544
rect 169944 661768 169996 661774
rect 169944 661710 169996 661716
rect 170220 661768 170272 661774
rect 170220 661710 170272 661716
rect 169956 656946 169984 661710
rect 299952 659682 299980 666538
rect 299768 659654 299980 659682
rect 364444 659682 364472 669258
rect 364444 659654 364564 659682
rect 169944 656940 169996 656946
rect 169944 656882 169996 656888
rect 170036 656940 170088 656946
rect 170036 656882 170088 656888
rect 139400 652860 139452 652866
rect 139400 652802 139452 652808
rect 137652 650480 137704 650486
rect 137652 650422 137704 650428
rect 137664 649720 137692 650422
rect 137650 649711 137706 649720
rect 137650 649646 137706 649655
rect 139412 589665 139440 652802
rect 140042 650992 140098 651001
rect 140098 650950 140176 650978
rect 140042 650927 140098 650936
rect 140148 650729 140176 650950
rect 140134 650720 140190 650729
rect 140134 650655 140190 650664
rect 147588 650480 147640 650486
rect 147640 650428 147720 650434
rect 147588 650422 147720 650428
rect 147600 650418 147720 650422
rect 157260 650418 157380 650434
rect 147600 650412 147732 650418
rect 147600 650406 147680 650412
rect 147680 650354 147732 650360
rect 157248 650412 157392 650418
rect 157300 650406 157340 650412
rect 157248 650354 157300 650360
rect 157340 650354 157392 650360
rect 164148 650344 164200 650350
rect 164240 650344 164292 650350
rect 164200 650292 164240 650298
rect 164148 650286 164292 650292
rect 164160 650270 164280 650286
rect 170048 647290 170076 656882
rect 299768 656878 299796 659654
rect 299480 656872 299532 656878
rect 299480 656814 299532 656820
rect 299756 656872 299808 656878
rect 299756 656814 299808 656820
rect 263508 653404 263560 653410
rect 263508 653346 263560 653352
rect 258630 652896 258686 652905
rect 258630 652831 258686 652840
rect 258644 652798 258672 652831
rect 263520 652798 263548 653346
rect 258632 652792 258684 652798
rect 258632 652734 258684 652740
rect 263508 652792 263560 652798
rect 263508 652734 263560 652740
rect 263520 651681 263548 652734
rect 263506 651672 263562 651681
rect 263506 651607 263562 651616
rect 197360 650956 197412 650962
rect 197360 650898 197412 650904
rect 206928 650956 206980 650962
rect 206928 650898 206980 650904
rect 197372 650826 197400 650898
rect 195244 650820 195296 650826
rect 195244 650762 195296 650768
rect 197360 650820 197412 650826
rect 206940 650808 206968 650898
rect 206940 650780 207060 650808
rect 197360 650762 197412 650768
rect 195256 650418 195284 650762
rect 207032 650622 207060 650780
rect 278780 650752 278832 650758
rect 278778 650720 278780 650729
rect 288348 650752 288400 650758
rect 278832 650720 278834 650729
rect 288348 650694 288400 650700
rect 292670 650720 292726 650729
rect 278778 650655 278834 650664
rect 207020 650616 207072 650622
rect 288360 650593 288388 650694
rect 292670 650655 292726 650664
rect 207020 650558 207072 650564
rect 237378 650584 237434 650593
rect 237378 650519 237380 650528
rect 237432 650519 237434 650528
rect 237562 650584 237618 650593
rect 237562 650519 237618 650528
rect 288346 650584 288402 650593
rect 288346 650519 288402 650528
rect 289818 650584 289874 650593
rect 292684 650554 292712 650655
rect 289818 650519 289820 650528
rect 237380 650490 237432 650496
rect 237576 650418 237604 650519
rect 289872 650519 289874 650528
rect 292672 650548 292724 650554
rect 289820 650490 289872 650496
rect 292672 650490 292724 650496
rect 266360 650480 266412 650486
rect 266360 650422 266412 650428
rect 195244 650412 195296 650418
rect 195244 650354 195296 650360
rect 237564 650412 237616 650418
rect 237564 650354 237616 650360
rect 266372 650078 266400 650422
rect 285588 650344 285640 650350
rect 285588 650286 285640 650292
rect 285600 650214 285628 650286
rect 285588 650208 285640 650214
rect 285588 650150 285640 650156
rect 280068 650140 280120 650146
rect 280068 650082 280120 650088
rect 266360 650072 266412 650078
rect 270500 650072 270552 650078
rect 266360 650014 266412 650020
rect 270498 650040 270500 650049
rect 280080 650049 280108 650082
rect 270552 650040 270554 650049
rect 266372 649890 266400 650014
rect 270498 649975 270554 649984
rect 280066 650040 280122 650049
rect 280066 649975 280122 649984
rect 266450 649904 266506 649913
rect 266372 649862 266450 649890
rect 266450 649839 266506 649848
rect 169944 647284 169996 647290
rect 169944 647226 169996 647232
rect 170036 647284 170088 647290
rect 170036 647226 170088 647232
rect 169956 640422 169984 647226
rect 188342 646096 188398 646105
rect 188342 646031 188398 646040
rect 169944 640416 169996 640422
rect 169944 640358 169996 640364
rect 170036 640416 170088 640422
rect 170036 640358 170088 640364
rect 170048 630698 170076 640358
rect 188250 637664 188306 637673
rect 188250 637599 188306 637608
rect 169852 630692 169904 630698
rect 169852 630634 169904 630640
rect 170036 630692 170088 630698
rect 170036 630634 170088 630640
rect 169864 630578 169892 630634
rect 169864 630550 169984 630578
rect 169956 621058 169984 630550
rect 169956 621030 170076 621058
rect 170048 611386 170076 621030
rect 169852 611380 169904 611386
rect 169852 611322 169904 611328
rect 170036 611380 170088 611386
rect 170036 611322 170088 611328
rect 169864 611266 169892 611322
rect 169864 611238 169984 611266
rect 169956 608598 169984 611238
rect 169852 608592 169904 608598
rect 169852 608534 169904 608540
rect 169944 608592 169996 608598
rect 169944 608534 169996 608540
rect 169864 601730 169892 608534
rect 169852 601724 169904 601730
rect 169852 601666 169904 601672
rect 170128 601724 170180 601730
rect 170128 601666 170180 601672
rect 170140 598942 170168 601666
rect 169944 598936 169996 598942
rect 169944 598878 169996 598884
rect 170128 598936 170180 598942
rect 170128 598878 170180 598884
rect 139398 589656 139454 589665
rect 139398 589591 139454 589600
rect 169956 589354 169984 598878
rect 169944 589348 169996 589354
rect 169944 589290 169996 589296
rect 170220 589348 170272 589354
rect 170220 589290 170272 589296
rect 170232 582486 170260 589290
rect 170220 582480 170272 582486
rect 170220 582422 170272 582428
rect 170128 582344 170180 582350
rect 170128 582286 170180 582292
rect 170140 572642 170168 582286
rect 169956 572614 170168 572642
rect 169956 563122 169984 572614
rect 169864 563094 169984 563122
rect 169864 562986 169892 563094
rect 169864 562958 169984 562986
rect 137376 558612 137428 558618
rect 137376 558554 137428 558560
rect 137388 542842 137416 558554
rect 144184 558476 144236 558482
rect 144184 558418 144236 558424
rect 140044 558408 140096 558414
rect 140044 558350 140096 558356
rect 137744 542972 137796 542978
rect 137744 542914 137796 542920
rect 137376 542836 137428 542842
rect 137376 542778 137428 542784
rect 137284 540864 137336 540870
rect 137284 540806 137336 540812
rect 137756 539988 137784 542914
rect 140056 542910 140084 558350
rect 140136 558340 140188 558346
rect 140136 558282 140188 558288
rect 139860 542904 139912 542910
rect 139860 542846 139912 542852
rect 140044 542904 140096 542910
rect 140044 542846 140096 542852
rect 139872 539988 139900 542846
rect 140148 542774 140176 558282
rect 141424 558204 141476 558210
rect 141424 558146 141476 558152
rect 140136 542768 140188 542774
rect 140136 542710 140188 542716
rect 141436 542434 141464 558146
rect 141516 557728 141568 557734
rect 141516 557670 141568 557676
rect 141528 543289 141556 557670
rect 141514 543280 141570 543289
rect 141514 543215 141570 543224
rect 144196 543153 144224 558418
rect 145564 558272 145616 558278
rect 145564 558214 145616 558220
rect 144828 545420 144880 545426
rect 144828 545362 144880 545368
rect 144840 545193 144868 545362
rect 144826 545184 144882 545193
rect 144826 545119 144882 545128
rect 144182 543144 144238 543153
rect 144182 543079 144238 543088
rect 145576 542570 145604 558214
rect 152464 558136 152516 558142
rect 152464 558078 152516 558084
rect 148324 558068 148376 558074
rect 148324 558010 148376 558016
rect 148140 544060 148192 544066
rect 148140 544002 148192 544008
rect 146024 542632 146076 542638
rect 146024 542574 146076 542580
rect 144000 542564 144052 542570
rect 144000 542506 144052 542512
rect 145564 542564 145616 542570
rect 145564 542506 145616 542512
rect 141884 542496 141936 542502
rect 141884 542438 141936 542444
rect 141424 542428 141476 542434
rect 141424 542370 141476 542376
rect 141896 539988 141924 542438
rect 144012 539988 144040 542506
rect 146036 539988 146064 542574
rect 148152 539988 148180 544002
rect 148336 542570 148364 558010
rect 152476 543726 152504 558078
rect 169956 553466 169984 562958
rect 169956 553438 170076 553466
rect 166908 545352 166960 545358
rect 166906 545320 166908 545329
rect 166960 545320 166962 545329
rect 166906 545255 166962 545264
rect 168840 544128 168892 544134
rect 168840 544070 168892 544076
rect 160560 543992 160612 543998
rect 160560 543934 160612 543940
rect 152280 543720 152332 543726
rect 152280 543662 152332 543668
rect 152464 543720 152516 543726
rect 152464 543662 152516 543668
rect 148324 542564 148376 542570
rect 148324 542506 148376 542512
rect 150164 542428 150216 542434
rect 150164 542370 150216 542376
rect 150176 539988 150204 542370
rect 152292 539988 152320 543662
rect 156420 543652 156472 543658
rect 156420 543594 156472 543600
rect 154396 542496 154448 542502
rect 154396 542438 154448 542444
rect 154408 539988 154436 542438
rect 156432 539988 156460 543594
rect 158536 542564 158588 542570
rect 158536 542506 158588 542512
rect 158548 539988 158576 542506
rect 160572 539988 160600 543934
rect 166816 543720 166868 543726
rect 166816 543662 166868 543668
rect 164700 543584 164752 543590
rect 164700 543526 164752 543532
rect 162676 542632 162728 542638
rect 162676 542574 162728 542580
rect 162688 539988 162716 542574
rect 164712 539988 164740 543526
rect 166828 539988 166856 543662
rect 168852 539988 168880 544070
rect 170048 540802 170076 553438
rect 177304 545352 177356 545358
rect 177302 545320 177304 545329
rect 177356 545320 177358 545329
rect 177302 545255 177358 545264
rect 177212 545012 177264 545018
rect 177212 544954 177264 544960
rect 173072 544332 173124 544338
rect 173072 544274 173124 544280
rect 170956 544196 171008 544202
rect 170956 544138 171008 544144
rect 170036 540796 170088 540802
rect 170036 540738 170088 540744
rect 170968 539988 170996 544138
rect 173084 539988 173112 544274
rect 175096 544264 175148 544270
rect 175096 544206 175148 544212
rect 175108 539988 175136 544206
rect 177224 539988 177252 544954
rect 181352 544944 181404 544950
rect 181352 544886 181404 544892
rect 179236 544808 179288 544814
rect 179236 544750 179288 544756
rect 179248 539988 179276 544750
rect 181364 539988 181392 544886
rect 188264 544377 188292 637599
rect 188356 544882 188384 646031
rect 188434 645008 188490 645017
rect 188434 644943 188490 644952
rect 188344 544876 188396 544882
rect 188344 544818 188396 544824
rect 188448 544678 188476 644943
rect 188526 643240 188582 643249
rect 188526 643175 188582 643184
rect 188540 544785 188568 643175
rect 188618 642016 188674 642025
rect 188618 641951 188674 641960
rect 188526 544776 188582 544785
rect 188526 544711 188582 544720
rect 188436 544672 188488 544678
rect 188436 544614 188488 544620
rect 188632 544610 188660 641951
rect 188710 640384 188766 640393
rect 188710 640319 188766 640328
rect 188724 544649 188752 640319
rect 188894 639296 188950 639305
rect 188894 639231 188950 639240
rect 188802 579728 188858 579737
rect 188802 579663 188858 579672
rect 188816 545766 188844 579663
rect 188804 545760 188856 545766
rect 188804 545702 188856 545708
rect 188710 544640 188766 544649
rect 188620 544604 188672 544610
rect 188710 544575 188766 544584
rect 188620 544546 188672 544552
rect 188908 544513 188936 639231
rect 269118 589384 269174 589393
rect 269118 589319 269174 589328
rect 270406 589384 270462 589393
rect 270406 589319 270408 589328
rect 269132 587761 269160 589319
rect 270460 589319 270462 589328
rect 270408 589290 270460 589296
rect 269118 587752 269174 587761
rect 269118 587687 269174 587696
rect 188986 578368 189042 578377
rect 188986 578303 189042 578312
rect 189000 560930 189028 578303
rect 188988 560924 189040 560930
rect 188988 560866 189040 560872
rect 210974 560008 211030 560017
rect 210974 559943 211030 559952
rect 195978 558920 196034 558929
rect 195978 558855 196034 558864
rect 197358 558920 197414 558929
rect 197358 558855 197360 558864
rect 194414 558784 194470 558793
rect 194414 558719 194470 558728
rect 194428 558006 194456 558719
rect 194416 558000 194468 558006
rect 194416 557942 194468 557948
rect 195886 545456 195942 545465
rect 195886 545391 195888 545400
rect 195940 545391 195942 545400
rect 195888 545362 195940 545368
rect 189632 544740 189684 544746
rect 189632 544682 189684 544688
rect 188894 544504 188950 544513
rect 188894 544439 188950 544448
rect 188250 544368 188306 544377
rect 188250 544303 188306 544312
rect 183376 543244 183428 543250
rect 183376 543186 183428 543192
rect 183388 539988 183416 543186
rect 187516 543176 187568 543182
rect 187516 543118 187568 543124
rect 185492 542700 185544 542706
rect 185492 542642 185544 542648
rect 185504 539988 185532 542642
rect 187528 539988 187556 543118
rect 189644 539988 189672 544682
rect 195992 544406 196020 558855
rect 197412 558855 197414 558864
rect 201498 558920 201554 558929
rect 201498 558855 201554 558864
rect 202786 558920 202842 558929
rect 202786 558855 202842 558864
rect 204166 558920 204222 558929
rect 204166 558855 204222 558864
rect 205546 558920 205602 558929
rect 205546 558855 205602 558864
rect 206098 558920 206154 558929
rect 206098 558855 206154 558864
rect 208398 558920 208454 558929
rect 208398 558855 208454 558864
rect 210606 558920 210662 558929
rect 210606 558855 210662 558864
rect 197360 558826 197412 558832
rect 201512 558822 201540 558855
rect 201500 558816 201552 558822
rect 201500 558758 201552 558764
rect 202142 558648 202198 558657
rect 202142 558583 202198 558592
rect 200120 558068 200172 558074
rect 200120 558010 200172 558016
rect 200028 558000 200080 558006
rect 200028 557942 200080 557948
rect 198738 557696 198794 557705
rect 198738 557631 198740 557640
rect 198792 557631 198794 557640
rect 198740 557602 198792 557608
rect 200040 557598 200068 557942
rect 200132 557598 200160 558010
rect 200210 557832 200266 557841
rect 202156 557802 202184 558583
rect 200210 557767 200212 557776
rect 200264 557767 200266 557776
rect 202144 557796 202196 557802
rect 200212 557738 200264 557744
rect 202144 557738 202196 557744
rect 200028 557592 200080 557598
rect 200028 557534 200080 557540
rect 200120 557592 200172 557598
rect 200120 557534 200172 557540
rect 201406 545456 201462 545465
rect 201406 545391 201408 545400
rect 201460 545391 201462 545400
rect 201408 545362 201460 545368
rect 202156 545086 202184 557738
rect 202144 545080 202196 545086
rect 202144 545022 202196 545028
rect 202052 544536 202104 544542
rect 202052 544478 202104 544484
rect 195980 544400 196032 544406
rect 195980 544342 196032 544348
rect 193772 543108 193824 543114
rect 193772 543050 193824 543056
rect 191748 542836 191800 542842
rect 191748 542778 191800 542784
rect 191760 539988 191788 542778
rect 193784 539988 193812 543050
rect 197912 543040 197964 543046
rect 197912 542982 197964 542988
rect 195888 542768 195940 542774
rect 195888 542710 195940 542716
rect 195900 539988 195928 542710
rect 197924 539988 197952 542982
rect 200028 542904 200080 542910
rect 200028 542846 200080 542852
rect 200040 539988 200068 542846
rect 202064 539988 202092 544478
rect 202800 543046 202828 558855
rect 203522 558784 203578 558793
rect 203522 558719 203578 558728
rect 203536 558006 203564 558719
rect 203524 558000 203576 558006
rect 203524 557942 203576 557948
rect 203536 543318 203564 557942
rect 203524 543312 203576 543318
rect 203524 543254 203576 543260
rect 204180 543182 204208 558855
rect 204902 558648 204958 558657
rect 204902 558583 204958 558592
rect 204916 557734 204944 558583
rect 204904 557728 204956 557734
rect 204904 557670 204956 557676
rect 204916 543386 204944 557670
rect 205560 543658 205588 558855
rect 206112 557870 206140 558855
rect 208412 558754 208440 558855
rect 208400 558748 208452 558754
rect 208400 558690 208452 558696
rect 209688 558748 209740 558754
rect 209688 558690 209740 558696
rect 209042 558648 209098 558657
rect 209042 558583 209098 558592
rect 208584 558408 208636 558414
rect 208584 558350 208636 558356
rect 206928 558204 206980 558210
rect 206928 558146 206980 558152
rect 206940 557870 206968 558146
rect 208596 557938 208624 558350
rect 208584 557932 208636 557938
rect 208584 557874 208636 557880
rect 209056 557870 209084 558583
rect 209700 558550 209728 558690
rect 209688 558544 209740 558550
rect 209688 558486 209740 558492
rect 210620 558414 210648 558855
rect 210608 558408 210660 558414
rect 210608 558350 210660 558356
rect 206100 557864 206152 557870
rect 206100 557806 206152 557812
rect 206928 557864 206980 557870
rect 206928 557806 206980 557812
rect 209044 557864 209096 557870
rect 209044 557806 209096 557812
rect 207662 557696 207718 557705
rect 207662 557631 207664 557640
rect 207716 557631 207718 557640
rect 207664 557602 207716 557608
rect 206926 557560 206982 557569
rect 206926 557495 206982 557504
rect 206940 543726 206968 557495
rect 207570 545728 207626 545737
rect 207570 545663 207626 545672
rect 207584 545465 207612 545663
rect 207570 545456 207626 545465
rect 207570 545391 207626 545400
rect 206928 543720 206980 543726
rect 206928 543662 206980 543668
rect 205548 543652 205600 543658
rect 205548 543594 205600 543600
rect 207676 543454 207704 557602
rect 208306 557560 208362 557569
rect 208306 557495 208362 557504
rect 208320 543590 208348 557495
rect 208308 543584 208360 543590
rect 208308 543526 208360 543532
rect 209056 543522 209084 557806
rect 209686 557560 209742 557569
rect 209686 557495 209742 557504
rect 209700 543522 209728 557495
rect 209044 543516 209096 543522
rect 209044 543458 209096 543464
rect 209688 543516 209740 543522
rect 209688 543458 209740 543464
rect 207664 543448 207716 543454
rect 207664 543390 207716 543396
rect 204904 543380 204956 543386
rect 204904 543322 204956 543328
rect 208306 543280 208362 543289
rect 210988 543250 211016 559943
rect 220082 559056 220138 559065
rect 220082 558991 220138 559000
rect 211802 558920 211858 558929
rect 211802 558855 211858 558864
rect 213090 558920 213146 558929
rect 213090 558855 213146 558864
rect 213918 558920 213974 558929
rect 213918 558855 213974 558864
rect 215298 558920 215354 558929
rect 215298 558855 215300 558864
rect 211816 558346 211844 558855
rect 211160 558340 211212 558346
rect 211160 558282 211212 558288
rect 211804 558340 211856 558346
rect 211804 558282 211856 558288
rect 211172 557802 211200 558282
rect 213104 558006 213132 558855
rect 213932 558482 213960 558855
rect 215352 558855 215354 558864
rect 217966 558920 218022 558929
rect 217966 558855 218022 558864
rect 218978 558920 219034 558929
rect 218978 558855 219034 558864
rect 215300 558826 215352 558832
rect 213920 558476 213972 558482
rect 213920 558418 213972 558424
rect 213644 558068 213696 558074
rect 213644 558010 213696 558016
rect 213092 558000 213144 558006
rect 213092 557942 213144 557948
rect 213656 557802 213684 558010
rect 211160 557796 211212 557802
rect 211160 557738 211212 557744
rect 213644 557796 213696 557802
rect 213644 557738 213696 557744
rect 213932 557734 213960 558418
rect 215114 558376 215170 558385
rect 215114 558311 215116 558320
rect 215168 558311 215170 558320
rect 215116 558282 215168 558288
rect 215312 558210 215340 558826
rect 217782 558784 217838 558793
rect 217782 558719 217838 558728
rect 217796 558618 217824 558719
rect 217784 558612 217836 558618
rect 217784 558554 217836 558560
rect 215300 558204 215352 558210
rect 215300 558146 215352 558152
rect 213920 557728 213972 557734
rect 211066 557696 211122 557705
rect 213920 557670 213972 557676
rect 217796 557666 217824 558554
rect 217980 558550 218008 558855
rect 217968 558544 218020 558550
rect 217968 558486 218020 558492
rect 217980 558414 218008 558486
rect 217968 558408 218020 558414
rect 217968 558350 218020 558356
rect 218992 558074 219020 558855
rect 220096 558346 220124 558991
rect 222382 558920 222438 558929
rect 222382 558855 222438 558864
rect 223578 558920 223634 558929
rect 223578 558855 223634 558864
rect 224498 558920 224554 558929
rect 224498 558855 224500 558864
rect 221554 558376 221610 558385
rect 220084 558340 220136 558346
rect 220084 558282 220136 558288
rect 220820 558340 220872 558346
rect 221096 558340 221148 558346
rect 220872 558300 221096 558328
rect 220820 558282 220872 558288
rect 221554 558311 221556 558320
rect 221096 558282 221148 558288
rect 221608 558311 221610 558320
rect 221556 558282 221608 558288
rect 222396 558278 222424 558855
rect 223592 558754 223620 558855
rect 224552 558855 224554 558864
rect 225878 558920 225934 558929
rect 225878 558855 225934 558864
rect 227166 558920 227222 558929
rect 227166 558855 227222 558864
rect 228178 558920 228234 558929
rect 228178 558855 228234 558864
rect 229558 558920 229614 558929
rect 229558 558855 229614 558864
rect 224500 558826 224552 558832
rect 223580 558748 223632 558754
rect 223580 558690 223632 558696
rect 223592 558550 223620 558690
rect 224512 558686 224540 558826
rect 224500 558680 224552 558686
rect 224500 558622 224552 558628
rect 225892 558618 225920 558855
rect 225880 558612 225932 558618
rect 225880 558554 225932 558560
rect 223580 558544 223632 558550
rect 223580 558486 223632 558492
rect 227180 558482 227208 558855
rect 227168 558476 227220 558482
rect 227168 558418 227220 558424
rect 222384 558272 222436 558278
rect 222384 558214 222436 558220
rect 228192 558210 228220 558855
rect 229572 558414 229600 558855
rect 231858 558784 231914 558793
rect 231858 558719 231860 558728
rect 231912 558719 231914 558728
rect 233238 558784 233294 558793
rect 233238 558719 233294 558728
rect 231860 558690 231912 558696
rect 233252 558686 233280 558719
rect 233240 558680 233292 558686
rect 233240 558622 233292 558628
rect 234894 558648 234950 558657
rect 234894 558583 234896 558592
rect 234948 558583 234950 558592
rect 237378 558648 237434 558657
rect 237378 558583 237434 558592
rect 234896 558554 234948 558560
rect 231950 558512 232006 558521
rect 231860 558476 231912 558482
rect 231912 558456 231950 558464
rect 231912 558447 232006 558456
rect 231912 558436 231992 558447
rect 231860 558418 231912 558424
rect 229560 558408 229612 558414
rect 229560 558350 229612 558356
rect 230478 558376 230534 558385
rect 230478 558311 230480 558320
rect 230532 558311 230534 558320
rect 231858 558376 231914 558385
rect 231858 558311 231914 558320
rect 230480 558282 230532 558288
rect 231872 558278 231900 558311
rect 231860 558272 231912 558278
rect 231860 558214 231912 558220
rect 237392 558210 237420 558583
rect 238758 558512 238814 558521
rect 238758 558447 238814 558456
rect 238772 558414 238800 558447
rect 238760 558408 238812 558414
rect 238760 558350 238812 558356
rect 228180 558204 228232 558210
rect 228180 558146 228232 558152
rect 237380 558204 237432 558210
rect 237380 558146 237432 558152
rect 283748 558136 283800 558142
rect 283748 558078 283800 558084
rect 218980 558068 219032 558074
rect 218980 558010 219032 558016
rect 218992 557870 219020 558010
rect 218980 557864 219032 557870
rect 229098 557832 229154 557841
rect 218980 557806 219032 557812
rect 222120 557802 222240 557818
rect 222108 557796 222252 557802
rect 222160 557790 222200 557796
rect 222108 557738 222160 557744
rect 229098 557767 229100 557776
rect 222200 557738 222252 557744
rect 229152 557767 229154 557776
rect 238666 557832 238722 557841
rect 238666 557767 238722 557776
rect 229100 557738 229152 557744
rect 217874 557696 217930 557705
rect 211066 557631 211122 557640
rect 217784 557660 217836 557666
rect 211080 543454 211108 557631
rect 217874 557631 217930 557640
rect 226154 557696 226210 557705
rect 226154 557631 226210 557640
rect 233146 557696 233202 557705
rect 238680 557666 238708 557767
rect 241612 557728 241664 557734
rect 283656 557728 283708 557734
rect 241612 557670 241664 557676
rect 233146 557631 233202 557640
rect 238668 557660 238720 557666
rect 217784 557602 217836 557608
rect 212446 557560 212502 557569
rect 212446 557495 212502 557504
rect 213826 557560 213882 557569
rect 213826 557495 213882 557504
rect 215206 557560 215262 557569
rect 215206 557495 215262 557504
rect 216586 557560 216642 557569
rect 216586 557495 216642 557504
rect 212172 544468 212224 544474
rect 212172 544410 212224 544416
rect 211068 543448 211120 543454
rect 211068 543390 211120 543396
rect 208306 543215 208362 543224
rect 210976 543244 211028 543250
rect 204168 543176 204220 543182
rect 204168 543118 204220 543124
rect 202788 543040 202840 543046
rect 202788 542982 202840 542988
rect 206190 543008 206246 543017
rect 204168 542972 204220 542978
rect 206190 542943 206246 542952
rect 204168 542914 204220 542920
rect 204180 539988 204208 542914
rect 206204 539988 206232 542943
rect 208320 539988 208348 543215
rect 210976 543186 211028 543192
rect 210422 543144 210478 543153
rect 210422 543079 210478 543088
rect 210436 539988 210464 543079
rect 212184 540002 212212 544410
rect 212460 543386 212488 557495
rect 212538 545456 212594 545465
rect 212538 545391 212540 545400
rect 212592 545391 212594 545400
rect 212540 545362 212592 545368
rect 212448 543380 212500 543386
rect 212448 543322 212500 543328
rect 213840 543114 213868 557495
rect 215220 543318 215248 557495
rect 215208 543312 215260 543318
rect 215208 543254 215260 543260
rect 216600 543182 216628 557495
rect 216220 543176 216272 543182
rect 216220 543118 216272 543124
rect 216588 543176 216640 543182
rect 216588 543118 216640 543124
rect 213828 543108 213880 543114
rect 213828 543050 213880 543056
rect 214564 543040 214616 543046
rect 214564 542982 214616 542988
rect 212184 539974 212474 540002
rect 214576 539988 214604 542982
rect 216232 540002 216260 543118
rect 217888 543046 217916 557631
rect 217966 557560 218022 557569
rect 217966 557495 218022 557504
rect 219346 557560 219402 557569
rect 219346 557495 219402 557504
rect 220726 557560 220782 557569
rect 220726 557495 220782 557504
rect 222106 557560 222162 557569
rect 222106 557495 222162 557504
rect 223486 557560 223542 557569
rect 223486 557495 223542 557504
rect 224866 557560 224922 557569
rect 224866 557495 224922 557504
rect 217876 543040 217928 543046
rect 217876 542982 217928 542988
rect 217980 542570 218008 557495
rect 218704 543652 218756 543658
rect 218704 543594 218756 543600
rect 217968 542564 218020 542570
rect 217968 542506 218020 542512
rect 216232 539974 216614 540002
rect 218716 539988 218744 543594
rect 219360 542502 219388 557495
rect 220452 543720 220504 543726
rect 220452 543662 220504 543668
rect 219348 542496 219400 542502
rect 219348 542438 219400 542444
rect 220464 540002 220492 543662
rect 220740 542638 220768 557495
rect 222016 545420 222068 545426
rect 222016 545362 222068 545368
rect 222028 545193 222056 545362
rect 222014 545184 222070 545193
rect 222014 545119 222070 545128
rect 222120 542706 222148 557495
rect 222844 543584 222896 543590
rect 222844 543526 222896 543532
rect 222108 542700 222160 542706
rect 222108 542642 222160 542648
rect 220728 542632 220780 542638
rect 220728 542574 220780 542580
rect 220464 539974 220754 540002
rect 222856 539988 222884 543526
rect 223500 542842 223528 557495
rect 224500 543516 224552 543522
rect 224500 543458 224552 543464
rect 223488 542836 223540 542842
rect 223488 542778 223540 542784
rect 224512 540002 224540 543458
rect 224880 542774 224908 557495
rect 226168 542910 226196 557631
rect 226246 557560 226302 557569
rect 226246 557495 226302 557504
rect 227626 557560 227682 557569
rect 227626 557495 227682 557504
rect 229006 557560 229062 557569
rect 229006 557495 229062 557504
rect 230386 557560 230442 557569
rect 230386 557495 230442 557504
rect 231766 557560 231822 557569
rect 231766 557495 231822 557504
rect 233054 557560 233110 557569
rect 233054 557495 233110 557504
rect 226260 542978 226288 557495
rect 227640 543658 227668 557495
rect 229020 543726 229048 557495
rect 229008 543720 229060 543726
rect 229008 543662 229060 543668
rect 227628 543652 227680 543658
rect 227628 543594 227680 543600
rect 230400 543590 230428 557495
rect 230388 543584 230440 543590
rect 230388 543526 230440 543532
rect 231780 543522 231808 557495
rect 231858 545456 231914 545465
rect 231858 545391 231860 545400
rect 231912 545391 231914 545400
rect 231860 545362 231912 545368
rect 231768 543516 231820 543522
rect 231768 543458 231820 543464
rect 226984 543448 227036 543454
rect 226984 543390 227036 543396
rect 226248 542972 226300 542978
rect 226248 542914 226300 542920
rect 226156 542904 226208 542910
rect 226156 542846 226208 542852
rect 224868 542768 224920 542774
rect 224868 542710 224920 542716
rect 224512 539974 224894 540002
rect 226996 539988 227024 543390
rect 233068 543386 233096 557495
rect 233160 543454 233188 557631
rect 238668 557602 238720 557608
rect 241624 557569 241652 557670
rect 253860 557666 253980 557682
rect 273180 557666 273300 557682
rect 283656 557670 283708 557676
rect 251088 557660 251140 557666
rect 251088 557602 251140 557608
rect 253848 557660 253992 557666
rect 253900 557654 253940 557660
rect 253848 557602 253900 557608
rect 253940 557602 253992 557608
rect 270408 557660 270460 557666
rect 270408 557602 270460 557608
rect 273168 557660 273312 557666
rect 273220 557654 273260 557660
rect 273168 557602 273220 557608
rect 273260 557602 273312 557608
rect 283564 557660 283616 557666
rect 283564 557602 283616 557608
rect 251100 557569 251128 557602
rect 260840 557592 260892 557598
rect 234526 557560 234582 557569
rect 234526 557495 234582 557504
rect 235906 557560 235962 557569
rect 235906 557495 235962 557504
rect 237286 557560 237342 557569
rect 237286 557495 237342 557504
rect 238666 557560 238722 557569
rect 238666 557495 238722 557504
rect 240046 557560 240102 557569
rect 240046 557495 240102 557504
rect 241610 557560 241666 557569
rect 241610 557495 241666 557504
rect 251086 557560 251142 557569
rect 251086 557495 251142 557504
rect 260838 557560 260840 557569
rect 270420 557569 270448 557602
rect 282368 557592 282420 557598
rect 260892 557560 260894 557569
rect 260838 557495 260894 557504
rect 270406 557560 270462 557569
rect 282368 557534 282420 557540
rect 270406 557495 270462 557504
rect 233148 543448 233200 543454
rect 233148 543390 233200 543396
rect 231124 543380 231176 543386
rect 231124 543322 231176 543328
rect 233056 543380 233108 543386
rect 233056 543322 233108 543328
rect 229100 543244 229152 543250
rect 229100 543186 229152 543192
rect 229112 539988 229140 543186
rect 231136 539988 231164 543322
rect 234540 543250 234568 557495
rect 235920 543318 235948 557495
rect 235264 543312 235316 543318
rect 235264 543254 235316 543260
rect 235908 543312 235960 543318
rect 235908 543254 235960 543260
rect 234528 543244 234580 543250
rect 234528 543186 234580 543192
rect 233240 543108 233292 543114
rect 233240 543050 233292 543056
rect 233252 539988 233280 543050
rect 235276 539988 235304 543254
rect 237300 543114 237328 557495
rect 238680 543182 238708 557495
rect 237380 543176 237432 543182
rect 237380 543118 237432 543124
rect 238668 543176 238720 543182
rect 238668 543118 238720 543124
rect 237288 543108 237340 543114
rect 237288 543050 237340 543056
rect 237392 539988 237420 543118
rect 240060 543046 240088 557495
rect 282380 549302 282408 557534
rect 282368 549296 282420 549302
rect 282368 549238 282420 549244
rect 282460 549296 282512 549302
rect 282460 549238 282512 549244
rect 251178 545456 251234 545465
rect 241428 545420 241480 545426
rect 251178 545391 251180 545400
rect 241428 545362 241480 545368
rect 251232 545391 251234 545400
rect 260748 545420 260800 545426
rect 251180 545362 251232 545368
rect 260748 545362 260800 545368
rect 241440 545193 241468 545362
rect 260760 545193 260788 545362
rect 241426 545184 241482 545193
rect 241426 545119 241482 545128
rect 260746 545184 260802 545193
rect 260746 545119 260802 545128
rect 260196 543720 260248 543726
rect 260196 543662 260248 543668
rect 258080 543652 258132 543658
rect 258080 543594 258132 543600
rect 239404 543040 239456 543046
rect 239404 542982 239456 542988
rect 240048 543040 240100 543046
rect 240048 542982 240100 542988
rect 239416 539988 239444 542982
rect 256056 542972 256108 542978
rect 256056 542914 256108 542920
rect 253940 542904 253992 542910
rect 253940 542846 253992 542852
rect 249800 542836 249852 542842
rect 249800 542778 249852 542784
rect 247776 542700 247828 542706
rect 247776 542642 247828 542648
rect 245660 542632 245712 542638
rect 245660 542574 245712 542580
rect 241520 542564 241572 542570
rect 241520 542506 241572 542512
rect 241532 539988 241560 542506
rect 243544 542496 243596 542502
rect 243544 542438 243596 542444
rect 243556 539988 243584 542438
rect 245672 539988 245700 542574
rect 247788 539988 247816 542642
rect 249812 539988 249840 542778
rect 251916 542768 251968 542774
rect 251916 542710 251968 542716
rect 251928 539988 251956 542710
rect 253952 539988 253980 542846
rect 256068 539988 256096 542914
rect 258092 539988 258120 543594
rect 260208 539988 260236 543662
rect 262220 543584 262272 543590
rect 262220 543526 262272 543532
rect 262232 539988 262260 543526
rect 264336 543516 264388 543522
rect 264336 543458 264388 543464
rect 264348 539988 264376 543458
rect 266452 543448 266504 543454
rect 266452 543390 266504 543396
rect 266464 539988 266492 543390
rect 268476 543380 268528 543386
rect 268476 543322 268528 543328
rect 268488 539988 268516 543322
rect 272616 543312 272668 543318
rect 272616 543254 272668 543260
rect 270592 543244 270644 543250
rect 270592 543186 270644 543192
rect 270604 539988 270632 543186
rect 272628 539988 272656 543254
rect 276756 543176 276808 543182
rect 276756 543118 276808 543124
rect 274732 543108 274784 543114
rect 274732 543050 274784 543056
rect 274744 539988 274772 543050
rect 276768 539988 276796 543118
rect 278872 543040 278924 543046
rect 278872 542982 278924 542988
rect 278884 539988 278912 542982
rect 282472 539594 282500 549238
rect 282472 539566 282592 539594
rect 282564 524482 282592 539566
rect 282552 524476 282604 524482
rect 282552 524418 282604 524424
rect 282644 524340 282696 524346
rect 282644 524282 282696 524288
rect 282656 521642 282684 524282
rect 282564 521614 282684 521642
rect 282564 514826 282592 521614
rect 282552 514820 282604 514826
rect 282552 514762 282604 514768
rect 282644 514752 282696 514758
rect 282644 514694 282696 514700
rect 282656 512038 282684 514694
rect 282552 512032 282604 512038
rect 282552 511974 282604 511980
rect 282644 512032 282696 512038
rect 282644 511974 282696 511980
rect 282564 505170 282592 511974
rect 282552 505164 282604 505170
rect 282552 505106 282604 505112
rect 282644 505028 282696 505034
rect 282644 504970 282696 504976
rect 282656 502330 282684 504970
rect 282564 502302 282684 502330
rect 282564 497554 282592 502302
rect 282368 497548 282420 497554
rect 282368 497490 282420 497496
rect 282552 497548 282604 497554
rect 282552 497490 282604 497496
rect 282380 492697 282408 497490
rect 282366 492688 282422 492697
rect 282366 492623 282422 492632
rect 282550 492688 282606 492697
rect 282550 492623 282606 492632
rect 282564 485858 282592 492623
rect 282552 485852 282604 485858
rect 282552 485794 282604 485800
rect 282644 485716 282696 485722
rect 282644 485658 282696 485664
rect 282656 483002 282684 485658
rect 282368 482996 282420 483002
rect 282368 482938 282420 482944
rect 282644 482996 282696 483002
rect 282644 482938 282696 482944
rect 282380 473385 282408 482938
rect 282366 473376 282422 473385
rect 282366 473311 282422 473320
rect 282550 473376 282606 473385
rect 282550 473311 282606 473320
rect 282564 466478 282592 473311
rect 282552 466472 282604 466478
rect 282552 466414 282604 466420
rect 282644 466404 282696 466410
rect 282644 466346 282696 466352
rect 282656 463690 282684 466346
rect 282368 463684 282420 463690
rect 282368 463626 282420 463632
rect 282644 463684 282696 463690
rect 282644 463626 282696 463632
rect 282380 454073 282408 463626
rect 282366 454064 282422 454073
rect 282366 453999 282422 454008
rect 282550 454064 282606 454073
rect 282550 453999 282606 454008
rect 282564 447166 282592 453999
rect 282552 447160 282604 447166
rect 282552 447102 282604 447108
rect 282644 447092 282696 447098
rect 282644 447034 282696 447040
rect 282656 437458 282684 447034
rect 282656 437430 282868 437458
rect 282840 434722 282868 437430
rect 282828 434716 282880 434722
rect 282828 434658 282880 434664
rect 283012 434716 283064 434722
rect 283012 434658 283064 434664
rect 281538 429448 281594 429457
rect 281538 429383 281594 429392
rect 281552 429214 281580 429383
rect 281540 429208 281592 429214
rect 281540 429150 281592 429156
rect 281538 428496 281594 428505
rect 281538 428431 281594 428440
rect 281552 427854 281580 428431
rect 281540 427848 281592 427854
rect 281540 427790 281592 427796
rect 281630 427408 281686 427417
rect 281630 427343 281686 427352
rect 281644 426562 281672 427343
rect 281632 426556 281684 426562
rect 281632 426498 281684 426504
rect 281540 426488 281592 426494
rect 281538 426456 281540 426465
rect 281592 426456 281594 426465
rect 281538 426391 281594 426400
rect 281538 425368 281594 425377
rect 281538 425303 281594 425312
rect 281552 425134 281580 425303
rect 281540 425128 281592 425134
rect 283024 425105 283052 434658
rect 281540 425070 281592 425076
rect 282642 425096 282698 425105
rect 282642 425031 282698 425040
rect 283010 425096 283066 425105
rect 283010 425031 283066 425040
rect 281538 424416 281594 424425
rect 281538 424351 281594 424360
rect 281552 423706 281580 424351
rect 281540 423700 281592 423706
rect 281540 423642 281592 423648
rect 281630 423464 281686 423473
rect 281630 423399 281686 423408
rect 281644 422414 281672 423399
rect 281632 422408 281684 422414
rect 281538 422376 281594 422385
rect 281632 422350 281684 422356
rect 281538 422311 281540 422320
rect 281592 422311 281594 422320
rect 281540 422282 281592 422288
rect 281538 421424 281594 421433
rect 281538 421359 281594 421368
rect 281552 420986 281580 421359
rect 281540 420980 281592 420986
rect 281540 420922 281592 420928
rect 281538 420336 281594 420345
rect 281538 420271 281594 420280
rect 281552 419558 281580 420271
rect 281540 419552 281592 419558
rect 281540 419494 281592 419500
rect 59912 419484 59964 419490
rect 59912 419426 59964 419432
rect 281630 419384 281686 419393
rect 281630 419319 281686 419328
rect 281538 418296 281594 418305
rect 281644 418266 281672 419319
rect 281538 418231 281594 418240
rect 281632 418260 281684 418266
rect 281552 418198 281580 418231
rect 281632 418202 281684 418208
rect 281540 418192 281592 418198
rect 281540 418134 281592 418140
rect 282274 416392 282330 416401
rect 282274 416327 282330 416336
rect 282288 415478 282316 416327
rect 282276 415472 282328 415478
rect 282276 415414 282328 415420
rect 281722 415304 281778 415313
rect 281722 415239 281778 415248
rect 281736 414118 281764 415239
rect 282090 414352 282146 414361
rect 282090 414287 282146 414296
rect 281724 414112 281776 414118
rect 281724 414054 281776 414060
rect 282104 414050 282132 414287
rect 282092 414044 282144 414050
rect 282092 413986 282144 413992
rect 282656 413982 282684 425031
rect 282826 417344 282882 417353
rect 282826 417279 282882 417288
rect 282840 416838 282868 417279
rect 282828 416832 282880 416838
rect 282828 416774 282880 416780
rect 282644 413976 282696 413982
rect 282642 413944 282644 413953
rect 282696 413944 282698 413953
rect 282642 413879 282698 413888
rect 282656 413853 282684 413879
rect 282644 413704 282696 413710
rect 59818 413672 59874 413681
rect 282644 413646 282696 413652
rect 59818 413607 59874 413616
rect 281540 413636 281592 413642
rect 281540 413578 281592 413584
rect 281552 412842 281580 413578
rect 281816 413500 281868 413506
rect 281816 413442 281868 413448
rect 281460 412814 281580 412842
rect 281460 412434 281488 412814
rect 281540 412752 281592 412758
rect 281540 412694 281592 412700
rect 281632 412752 281684 412758
rect 281632 412694 281684 412700
rect 281552 412622 281580 412694
rect 281540 412616 281592 412622
rect 281540 412558 281592 412564
rect 281644 412570 281672 412694
rect 281644 412542 281764 412570
rect 281828 412554 281856 413442
rect 282184 413364 282236 413370
rect 282184 413306 282236 413312
rect 282000 413092 282052 413098
rect 282000 413034 282052 413040
rect 281460 412406 281672 412434
rect 281540 412344 281592 412350
rect 281540 412286 281592 412292
rect 59726 396264 59782 396273
rect 59726 396199 59782 396208
rect 59634 390416 59690 390425
rect 59634 390351 59690 390360
rect 59542 384704 59598 384713
rect 59542 384639 59598 384648
rect 57610 378856 57666 378865
rect 57610 378791 57666 378800
rect 57794 376952 57850 376961
rect 57794 376887 57850 376896
rect 57702 373144 57758 373153
rect 57702 373079 57758 373088
rect 57610 367296 57666 367305
rect 57610 367231 57666 367240
rect 57518 363488 57574 363497
rect 57518 363423 57574 363432
rect 57428 338088 57480 338094
rect 57428 338030 57480 338036
rect 57426 334520 57482 334529
rect 57426 334455 57482 334464
rect 57336 295316 57388 295322
rect 57336 295258 57388 295264
rect 57244 252544 57296 252550
rect 57244 252486 57296 252492
rect 57440 135250 57468 334455
rect 57532 325242 57560 363423
rect 57520 325236 57572 325242
rect 57520 325178 57572 325184
rect 57624 325122 57652 367231
rect 57532 325094 57652 325122
rect 57716 325106 57744 373079
rect 57808 336734 57836 376887
rect 57886 369200 57942 369209
rect 57886 369135 57942 369144
rect 57796 336728 57848 336734
rect 57796 336670 57848 336676
rect 57794 336424 57850 336433
rect 57794 336359 57850 336368
rect 57808 329390 57836 336359
rect 57796 329384 57848 329390
rect 57796 329326 57848 329332
rect 57796 329248 57848 329254
rect 57796 329190 57848 329196
rect 57704 325100 57756 325106
rect 57532 320686 57560 325094
rect 57704 325042 57756 325048
rect 57808 324986 57836 329190
rect 57900 325174 57928 369135
rect 59450 349888 59506 349897
rect 59450 349823 59506 349832
rect 59358 344176 59414 344185
rect 59358 344111 59414 344120
rect 59082 338328 59138 338337
rect 59082 338263 59138 338272
rect 57980 325508 58032 325514
rect 57980 325450 58032 325456
rect 57888 325168 57940 325174
rect 57888 325110 57940 325116
rect 57992 324986 58020 325450
rect 57624 324958 57836 324986
rect 57900 324958 58020 324986
rect 57520 320680 57572 320686
rect 57520 320622 57572 320628
rect 57624 320618 57652 324958
rect 57794 324864 57850 324873
rect 57794 324799 57850 324808
rect 57702 322960 57758 322969
rect 57702 322895 57758 322904
rect 57612 320612 57664 320618
rect 57612 320554 57664 320560
rect 57428 135244 57480 135250
rect 57428 135186 57480 135192
rect 57060 88324 57112 88330
rect 57060 88266 57112 88272
rect 57716 41410 57744 322895
rect 57704 41404 57756 41410
rect 57704 41346 57756 41352
rect 57808 30326 57836 324799
rect 57900 321178 57928 324958
rect 57900 321150 58020 321178
rect 57886 321056 57942 321065
rect 57886 320991 57942 321000
rect 57796 30320 57848 30326
rect 57796 30262 57848 30268
rect 57900 17950 57928 320991
rect 57992 320754 58020 321150
rect 57980 320748 58032 320754
rect 57980 320690 58032 320696
rect 59096 158710 59124 338263
rect 59174 332616 59230 332625
rect 59174 332551 59230 332560
rect 59084 158704 59136 158710
rect 59084 158646 59136 158652
rect 59188 111790 59216 332551
rect 59266 326768 59322 326777
rect 59266 326703 59322 326712
rect 59176 111784 59228 111790
rect 59176 111726 59228 111732
rect 59280 64870 59308 326703
rect 59372 205630 59400 344111
rect 59464 252550 59492 349823
rect 59728 336728 59780 336734
rect 59780 336676 59952 336682
rect 59728 336670 59952 336676
rect 59740 336654 59952 336670
rect 59820 330880 59872 330886
rect 59820 330822 59872 330828
rect 59726 330712 59782 330721
rect 59726 330647 59782 330656
rect 59544 325168 59596 325174
rect 59544 325110 59596 325116
rect 59556 320550 59584 325110
rect 59636 325100 59688 325106
rect 59636 325042 59688 325048
rect 59544 320544 59596 320550
rect 59544 320486 59596 320492
rect 59648 320006 59676 325042
rect 59740 320482 59768 330647
rect 59728 320476 59780 320482
rect 59728 320418 59780 320424
rect 59832 320074 59860 330822
rect 59820 320068 59872 320074
rect 59820 320010 59872 320016
rect 59636 320000 59688 320006
rect 59636 319942 59688 319948
rect 59924 319938 59952 336654
rect 281552 330018 281580 412286
rect 281644 407862 281672 412406
rect 281632 407856 281684 407862
rect 281632 407798 281684 407804
rect 281632 407720 281684 407726
rect 281632 407662 281684 407668
rect 281644 403050 281672 407662
rect 281736 405249 281764 412542
rect 281816 412548 281868 412554
rect 281816 412490 281868 412496
rect 281816 412412 281868 412418
rect 281816 412354 281868 412360
rect 281828 406201 281856 412354
rect 281908 412004 281960 412010
rect 281908 411946 281960 411952
rect 281920 411330 281948 411946
rect 281908 411324 281960 411330
rect 281908 411266 281960 411272
rect 281908 411188 281960 411194
rect 281908 411130 281960 411136
rect 281920 410281 281948 411130
rect 281906 410272 281962 410281
rect 281906 410207 281962 410216
rect 281908 410168 281960 410174
rect 281908 410110 281960 410116
rect 281920 407726 281948 410110
rect 282012 407810 282040 413034
rect 282092 412820 282144 412826
rect 282092 412762 282144 412768
rect 282104 412418 282132 412762
rect 282092 412412 282144 412418
rect 282092 412354 282144 412360
rect 282090 412312 282146 412321
rect 282090 412247 282146 412256
rect 282104 411806 282132 412247
rect 282092 411800 282144 411806
rect 282092 411742 282144 411748
rect 282092 411596 282144 411602
rect 282092 411538 282144 411544
rect 282104 407930 282132 411538
rect 282196 407930 282224 413306
rect 282368 413160 282420 413166
rect 282368 413102 282420 413108
rect 282276 412956 282328 412962
rect 282276 412898 282328 412904
rect 282092 407924 282144 407930
rect 282092 407866 282144 407872
rect 282184 407924 282236 407930
rect 282184 407866 282236 407872
rect 282012 407782 282224 407810
rect 281908 407720 281960 407726
rect 281908 407662 281960 407668
rect 282000 407720 282052 407726
rect 282052 407668 282132 407674
rect 282000 407662 282132 407668
rect 282012 407646 282132 407662
rect 281908 407584 281960 407590
rect 281908 407526 281960 407532
rect 282000 407584 282052 407590
rect 282000 407526 282052 407532
rect 281814 406192 281870 406201
rect 281814 406127 281870 406136
rect 281722 405240 281778 405249
rect 281722 405175 281778 405184
rect 281920 403209 281948 407526
rect 281906 403200 281962 403209
rect 281906 403135 281962 403144
rect 281644 403022 281948 403050
rect 281632 401192 281684 401198
rect 281630 401160 281632 401169
rect 281684 401160 281686 401169
rect 281630 401095 281686 401104
rect 281630 400208 281686 400217
rect 281630 400143 281632 400152
rect 281684 400143 281686 400152
rect 281632 400114 281684 400120
rect 281632 399560 281684 399566
rect 281632 399502 281684 399508
rect 281644 399129 281672 399502
rect 281630 399120 281686 399129
rect 281630 399055 281686 399064
rect 281632 394596 281684 394602
rect 281632 394538 281684 394544
rect 281644 394097 281672 394538
rect 281630 394088 281686 394097
rect 281630 394023 281686 394032
rect 281722 393272 281778 393281
rect 281722 393207 281778 393216
rect 281816 393236 281868 393242
rect 281632 393168 281684 393174
rect 281630 393136 281632 393145
rect 281684 393136 281686 393145
rect 281630 393071 281686 393080
rect 281632 392420 281684 392426
rect 281632 392362 281684 392368
rect 281644 392057 281672 392362
rect 281630 392048 281686 392057
rect 281630 391983 281686 391992
rect 281632 388204 281684 388210
rect 281632 388146 281684 388152
rect 281644 388113 281672 388146
rect 281630 388104 281686 388113
rect 281630 388039 281686 388048
rect 281632 387048 281684 387054
rect 281630 387016 281632 387025
rect 281684 387016 281686 387025
rect 281630 386951 281686 386960
rect 281736 386186 281764 393207
rect 281816 393178 281868 393184
rect 281644 386158 281764 386186
rect 281644 385778 281672 386158
rect 281724 386096 281776 386102
rect 281722 386064 281724 386073
rect 281776 386064 281778 386073
rect 281722 385999 281778 386008
rect 281644 385750 281764 385778
rect 281632 385620 281684 385626
rect 281632 385562 281684 385568
rect 281644 385121 281672 385562
rect 281630 385112 281686 385121
rect 281630 385047 281686 385056
rect 281632 384940 281684 384946
rect 281632 384882 281684 384888
rect 281644 384033 281672 384882
rect 281630 384024 281686 384033
rect 281630 383959 281686 383968
rect 281736 383858 281764 385750
rect 281724 383852 281776 383858
rect 281724 383794 281776 383800
rect 281828 383790 281856 393178
rect 281920 390153 281948 403022
rect 281906 390144 281962 390153
rect 281906 390079 281962 390088
rect 281816 383784 281868 383790
rect 281816 383726 281868 383732
rect 281724 382220 281776 382226
rect 281724 382162 281776 382168
rect 281632 382016 281684 382022
rect 281630 381984 281632 381993
rect 281684 381984 281686 381993
rect 281630 381919 281686 381928
rect 281736 381041 281764 382162
rect 281722 381032 281778 381041
rect 281722 380967 281778 380976
rect 281908 373992 281960 373998
rect 281908 373934 281960 373940
rect 281816 373856 281868 373862
rect 281816 373798 281868 373804
rect 281724 373788 281776 373794
rect 281724 373730 281776 373736
rect 281736 364546 281764 373730
rect 281724 364540 281776 364546
rect 281724 364482 281776 364488
rect 281828 364478 281856 373798
rect 281816 364472 281868 364478
rect 281816 364414 281868 364420
rect 281920 364410 281948 373934
rect 281908 364404 281960 364410
rect 281908 364346 281960 364352
rect 281724 361548 281776 361554
rect 281724 361490 281776 361496
rect 281736 360777 281764 361490
rect 281722 360768 281778 360777
rect 281722 360703 281778 360712
rect 281908 358760 281960 358766
rect 281908 358702 281960 358708
rect 281920 357785 281948 358702
rect 281906 357776 281962 357785
rect 281906 357711 281962 357720
rect 282012 356833 282040 407526
rect 281998 356824 282054 356833
rect 281998 356759 282054 356768
rect 282104 355745 282132 407646
rect 282196 402778 282224 407782
rect 282288 402898 282316 412898
rect 282380 407810 282408 413102
rect 282460 413024 282512 413030
rect 282460 412966 282512 412972
rect 282472 411482 282500 412966
rect 282472 411454 282592 411482
rect 282460 411392 282512 411398
rect 282460 411334 282512 411340
rect 282472 407969 282500 411334
rect 282458 407960 282514 407969
rect 282458 407895 282514 407904
rect 282380 407782 282500 407810
rect 282276 402892 282328 402898
rect 282276 402834 282328 402840
rect 282196 402750 282408 402778
rect 282276 402688 282328 402694
rect 282276 402630 282328 402636
rect 282184 402620 282236 402626
rect 282184 402562 282236 402568
rect 282196 402257 282224 402562
rect 282182 402248 282238 402257
rect 282182 402183 282238 402192
rect 282184 398200 282236 398206
rect 282182 398168 282184 398177
rect 282236 398168 282238 398177
rect 282182 398103 282238 398112
rect 282184 393304 282236 393310
rect 282184 393246 282236 393252
rect 282196 383722 282224 393246
rect 282184 383716 282236 383722
rect 282184 383658 282236 383664
rect 282184 378072 282236 378078
rect 282184 378014 282236 378020
rect 282196 376961 282224 378014
rect 282182 376952 282238 376961
rect 282182 376887 282238 376896
rect 282184 373924 282236 373930
rect 282184 373866 282236 373872
rect 282196 372881 282224 373866
rect 282182 372872 282238 372881
rect 282182 372807 282238 372816
rect 282184 371136 282236 371142
rect 282184 371078 282236 371084
rect 282196 369889 282224 371078
rect 282182 369880 282238 369889
rect 282182 369815 282238 369824
rect 282184 366988 282236 366994
rect 282184 366930 282236 366936
rect 282196 365809 282224 366930
rect 282182 365800 282238 365809
rect 282182 365735 282238 365744
rect 282184 362976 282236 362982
rect 282184 362918 282236 362924
rect 282090 355736 282146 355745
rect 282090 355671 282146 355680
rect 282196 354793 282224 362918
rect 282182 354784 282238 354793
rect 282182 354719 282238 354728
rect 281998 354648 282054 354657
rect 281998 354583 282054 354592
rect 282092 354612 282144 354618
rect 282012 351801 282040 354583
rect 282092 354554 282144 354560
rect 282104 352753 282132 354554
rect 282090 352744 282146 352753
rect 282090 352679 282146 352688
rect 281998 351792 282054 351801
rect 281998 351727 282054 351736
rect 282288 349761 282316 402630
rect 282380 393242 282408 402750
rect 282472 393281 282500 407782
rect 282564 393310 282592 411454
rect 282656 408082 282684 413646
rect 282828 413296 282880 413302
rect 282826 413264 282828 413273
rect 282880 413264 282882 413273
rect 282826 413199 282882 413208
rect 282736 412888 282788 412894
rect 282736 412830 282788 412836
rect 282748 412570 282776 412830
rect 282748 412542 282868 412570
rect 282736 412480 282788 412486
rect 282736 412422 282788 412428
rect 282748 408218 282776 412422
rect 282840 411398 282868 412542
rect 283472 412208 283524 412214
rect 283472 412150 283524 412156
rect 283380 412140 283432 412146
rect 283380 412082 283432 412088
rect 282920 412072 282972 412078
rect 282920 412014 282972 412020
rect 282828 411392 282880 411398
rect 282828 411334 282880 411340
rect 282828 411256 282880 411262
rect 282826 411224 282828 411233
rect 282880 411224 282882 411233
rect 282826 411159 282882 411168
rect 282932 411074 282960 412014
rect 283012 411732 283064 411738
rect 283012 411674 283064 411680
rect 282840 411046 282960 411074
rect 282840 408354 282868 411046
rect 282920 410644 282972 410650
rect 282920 410586 282972 410592
rect 282932 408513 282960 410586
rect 283024 409329 283052 411674
rect 283104 411528 283156 411534
rect 283104 411470 283156 411476
rect 283010 409320 283066 409329
rect 283010 409255 283066 409264
rect 282918 408504 282974 408513
rect 282918 408439 282974 408448
rect 282840 408326 283052 408354
rect 282748 408190 282868 408218
rect 282656 408054 282776 408082
rect 282644 407924 282696 407930
rect 282644 407866 282696 407872
rect 282552 393304 282604 393310
rect 282458 393272 282514 393281
rect 282368 393236 282420 393242
rect 282552 393246 282604 393252
rect 282458 393207 282514 393216
rect 282368 393178 282420 393184
rect 282368 383784 282420 383790
rect 282368 383726 282420 383732
rect 282460 383784 282512 383790
rect 282460 383726 282512 383732
rect 282380 373862 282408 383726
rect 282472 373862 282500 383726
rect 282552 383716 282604 383722
rect 282552 383658 282604 383664
rect 282564 373998 282592 383658
rect 282552 373992 282604 373998
rect 282552 373934 282604 373940
rect 282368 373856 282420 373862
rect 282368 373798 282420 373804
rect 282460 373856 282512 373862
rect 282460 373798 282512 373804
rect 282368 364472 282420 364478
rect 282368 364414 282420 364420
rect 282460 364472 282512 364478
rect 282460 364414 282512 364420
rect 282380 354657 282408 364414
rect 282366 354648 282422 354657
rect 282472 354618 282500 364414
rect 282552 364404 282604 364410
rect 282552 364346 282604 364352
rect 282366 354583 282422 354592
rect 282460 354612 282512 354618
rect 282460 354554 282512 354560
rect 282564 350713 282592 364346
rect 282656 353705 282684 407866
rect 282748 407590 282776 408054
rect 282736 407584 282788 407590
rect 282736 407526 282788 407532
rect 282840 407402 282868 408190
rect 282748 407374 282868 407402
rect 282748 362982 282776 407374
rect 283024 407266 283052 408326
rect 282840 407238 283052 407266
rect 282840 404410 282868 407238
rect 282840 404382 282960 404410
rect 282828 404320 282880 404326
rect 282826 404288 282828 404297
rect 282880 404288 282882 404297
rect 282826 404223 282882 404232
rect 282932 404138 282960 404382
rect 282840 404110 282960 404138
rect 282840 389065 282868 404110
rect 283116 401198 283144 411470
rect 283288 411460 283340 411466
rect 283288 411402 283340 411408
rect 283196 411324 283248 411330
rect 283196 411266 283248 411272
rect 283104 401192 283156 401198
rect 283104 401134 283156 401140
rect 283208 399566 283236 411266
rect 283300 400178 283328 411402
rect 283288 400172 283340 400178
rect 283288 400114 283340 400120
rect 283196 399560 283248 399566
rect 283196 399502 283248 399508
rect 282826 389056 282882 389065
rect 282826 388991 282882 389000
rect 283392 388210 283420 412082
rect 283380 388204 283432 388210
rect 283380 388146 283432 388152
rect 283484 387054 283512 412150
rect 283576 393174 283604 557602
rect 283564 393168 283616 393174
rect 283564 393110 283616 393116
rect 283668 392426 283696 557670
rect 283760 394602 283788 558078
rect 284116 412412 284168 412418
rect 284116 412354 284168 412360
rect 284024 412344 284076 412350
rect 284024 412286 284076 412292
rect 283932 410712 283984 410718
rect 283932 410654 283984 410660
rect 283840 410576 283892 410582
rect 283840 410518 283892 410524
rect 283748 394596 283800 394602
rect 283748 394538 283800 394544
rect 283656 392420 283708 392426
rect 283656 392362 283708 392368
rect 283472 387048 283524 387054
rect 283472 386990 283524 386996
rect 282828 383648 282880 383654
rect 282828 383590 282880 383596
rect 282840 383081 282868 383590
rect 282826 383072 282882 383081
rect 282826 383007 282882 383016
rect 282828 380860 282880 380866
rect 282828 380802 282880 380808
rect 282840 379953 282868 380802
rect 282826 379944 282882 379953
rect 282826 379879 282882 379888
rect 282828 379500 282880 379506
rect 282828 379442 282880 379448
rect 282840 379001 282868 379442
rect 282826 378992 282882 379001
rect 282826 378927 282882 378936
rect 282828 378140 282880 378146
rect 282828 378082 282880 378088
rect 282840 378049 282868 378082
rect 282826 378040 282882 378049
rect 282826 377975 282882 377984
rect 282828 376712 282880 376718
rect 282828 376654 282880 376660
rect 282840 376009 282868 376654
rect 282826 376000 282882 376009
rect 282826 375935 282882 375944
rect 282828 375352 282880 375358
rect 282828 375294 282880 375300
rect 282840 374921 282868 375294
rect 282826 374912 282882 374921
rect 282826 374847 282882 374856
rect 282828 373992 282880 373998
rect 282826 373960 282828 373969
rect 282880 373960 282882 373969
rect 282826 373895 282882 373904
rect 282828 372564 282880 372570
rect 282828 372506 282880 372512
rect 282840 371929 282868 372506
rect 282826 371920 282882 371929
rect 282826 371855 282882 371864
rect 282828 371204 282880 371210
rect 282828 371146 282880 371152
rect 282840 370977 282868 371146
rect 282826 370968 282882 370977
rect 282826 370903 282882 370912
rect 282828 369844 282880 369850
rect 282828 369786 282880 369792
rect 282840 368937 282868 369786
rect 282826 368928 282882 368937
rect 282826 368863 282882 368872
rect 282828 368484 282880 368490
rect 282828 368426 282880 368432
rect 282840 367849 282868 368426
rect 282826 367840 282882 367849
rect 282826 367775 282882 367784
rect 282828 367056 282880 367062
rect 282828 366998 282880 367004
rect 282840 366897 282868 366998
rect 282826 366888 282882 366897
rect 282826 366823 282882 366832
rect 282828 365696 282880 365702
rect 282828 365638 282880 365644
rect 282840 364857 282868 365638
rect 282826 364848 282882 364857
rect 282826 364783 282882 364792
rect 282828 364336 282880 364342
rect 282828 364278 282880 364284
rect 282840 363905 282868 364278
rect 282826 363896 282882 363905
rect 282826 363831 282882 363840
rect 282736 362976 282788 362982
rect 282736 362918 282788 362924
rect 282828 362908 282880 362914
rect 282828 362850 282880 362856
rect 282736 362840 282788 362846
rect 282840 362817 282868 362850
rect 282736 362782 282788 362788
rect 282826 362808 282882 362817
rect 282748 361865 282776 362782
rect 282826 362743 282882 362752
rect 282734 361856 282790 361865
rect 282734 361791 282790 361800
rect 282828 360188 282880 360194
rect 282828 360130 282880 360136
rect 282736 360120 282788 360126
rect 282736 360062 282788 360068
rect 282748 358873 282776 360062
rect 282840 359825 282868 360130
rect 282826 359816 282882 359825
rect 282826 359751 282882 359760
rect 282734 358864 282790 358873
rect 282734 358799 282790 358808
rect 282642 353696 282698 353705
rect 282642 353631 282698 353640
rect 282550 350704 282606 350713
rect 282550 350639 282606 350648
rect 282274 349752 282330 349761
rect 282274 349687 282330 349696
rect 282828 349104 282880 349110
rect 282828 349046 282880 349052
rect 282840 348673 282868 349046
rect 282826 348664 282882 348673
rect 282826 348599 282882 348608
rect 282828 347744 282880 347750
rect 282826 347712 282828 347721
rect 282880 347712 282882 347721
rect 282276 347676 282328 347682
rect 282826 347647 282882 347656
rect 282276 347618 282328 347624
rect 282288 346633 282316 347618
rect 282274 346624 282330 346633
rect 282274 346559 282330 346568
rect 282092 346384 282144 346390
rect 282092 346326 282144 346332
rect 282104 345681 282132 346326
rect 282090 345672 282146 345681
rect 282090 345607 282146 345616
rect 282826 344720 282882 344729
rect 282826 344655 282882 344664
rect 282840 344554 282868 344655
rect 282828 344548 282880 344554
rect 282828 344490 282880 344496
rect 282734 343632 282790 343641
rect 282552 343596 282604 343602
rect 282734 343567 282790 343576
rect 282552 343538 282604 343544
rect 282564 342689 282592 343538
rect 282748 343534 282776 343567
rect 282736 343528 282788 343534
rect 282736 343470 282788 343476
rect 282550 342680 282606 342689
rect 282550 342615 282606 342624
rect 282828 342236 282880 342242
rect 282828 342178 282880 342184
rect 282840 341601 282868 342178
rect 282826 341592 282882 341601
rect 282826 341527 282882 341536
rect 282458 340640 282514 340649
rect 282458 340575 282514 340584
rect 282090 339688 282146 339697
rect 282090 339623 282146 339632
rect 281998 336560 282054 336569
rect 281998 336495 282054 336504
rect 281814 334520 281870 334529
rect 281814 334455 281870 334464
rect 281632 333600 281684 333606
rect 281630 333568 281632 333577
rect 281684 333568 281686 333577
rect 281630 333503 281686 333512
rect 281632 331220 281684 331226
rect 281632 331162 281684 331168
rect 281644 330585 281672 331162
rect 281630 330576 281686 330585
rect 281630 330511 281686 330520
rect 281552 329990 281764 330018
rect 281632 329792 281684 329798
rect 281632 329734 281684 329740
rect 281540 329724 281592 329730
rect 281540 329666 281592 329672
rect 281552 329497 281580 329666
rect 281538 329488 281594 329497
rect 281538 329423 281594 329432
rect 281644 328545 281672 329734
rect 281630 328536 281686 328545
rect 281630 328471 281686 328480
rect 281540 328432 281592 328438
rect 281540 328374 281592 328380
rect 281552 327457 281580 328374
rect 281538 327448 281594 327457
rect 281538 327383 281594 327392
rect 281540 327072 281592 327078
rect 281540 327014 281592 327020
rect 281552 326505 281580 327014
rect 281538 326496 281594 326505
rect 281538 326431 281594 326440
rect 281540 325644 281592 325650
rect 281540 325586 281592 325592
rect 281552 324465 281580 325586
rect 281736 325553 281764 329990
rect 281828 326330 281856 334455
rect 282012 331838 282040 336495
rect 282000 331832 282052 331838
rect 282000 331774 282052 331780
rect 281906 331528 281962 331537
rect 281906 331463 281962 331472
rect 281920 326398 281948 331463
rect 282104 326618 282132 339623
rect 282366 338600 282422 338609
rect 282366 338535 282422 338544
rect 282184 333940 282236 333946
rect 282184 333882 282236 333888
rect 282196 332625 282224 333882
rect 282182 332616 282238 332625
rect 282182 332551 282238 332560
rect 282012 326590 282132 326618
rect 281908 326392 281960 326398
rect 281908 326334 281960 326340
rect 281816 326324 281868 326330
rect 281816 326266 281868 326272
rect 281722 325544 281778 325553
rect 281722 325479 281778 325488
rect 281538 324456 281594 324465
rect 281538 324391 281594 324400
rect 281540 324284 281592 324290
rect 281540 324226 281592 324232
rect 281552 323513 281580 324226
rect 281538 323504 281594 323513
rect 281538 323439 281594 323448
rect 281540 322924 281592 322930
rect 281540 322866 281592 322872
rect 281552 322425 281580 322866
rect 281538 322416 281594 322425
rect 281538 322351 281594 322360
rect 279974 320920 280030 320929
rect 279974 320855 280030 320864
rect 279988 320550 280016 320855
rect 280066 320648 280122 320657
rect 280066 320583 280068 320592
rect 280120 320583 280122 320592
rect 280068 320554 280120 320560
rect 282012 320550 282040 326590
rect 282092 326460 282144 326466
rect 282092 326402 282144 326408
rect 279976 320544 280028 320550
rect 282000 320544 282052 320550
rect 279976 320486 280028 320492
rect 280066 320512 280122 320521
rect 282000 320486 282052 320492
rect 280066 320447 280068 320456
rect 280120 320447 280122 320456
rect 280068 320418 280120 320424
rect 282104 320278 282132 326402
rect 282184 326392 282236 326398
rect 282184 326334 282236 326340
rect 282276 326392 282328 326398
rect 282276 326334 282328 326340
rect 282196 320958 282224 326334
rect 282184 320952 282236 320958
rect 282184 320894 282236 320900
rect 282288 320414 282316 326334
rect 282380 320618 282408 338535
rect 282368 320612 282420 320618
rect 282368 320554 282420 320560
rect 282472 320482 282500 340575
rect 282550 337648 282606 337657
rect 282550 337583 282606 337592
rect 282564 320890 282592 337583
rect 282642 335608 282698 335617
rect 282642 335543 282698 335552
rect 282656 326398 282684 335543
rect 283852 333606 283880 410518
rect 283944 382022 283972 410654
rect 284036 384946 284064 412286
rect 284128 385626 284156 412354
rect 284208 412276 284260 412282
rect 284208 412218 284260 412224
rect 284220 386102 284248 412218
rect 285036 411664 285088 411670
rect 285036 411606 285088 411612
rect 284944 411392 284996 411398
rect 284944 411334 284996 411340
rect 284956 398206 284984 411334
rect 285048 402626 285076 411606
rect 285036 402620 285088 402626
rect 285036 402562 285088 402568
rect 284944 398200 284996 398206
rect 284944 398142 284996 398148
rect 284208 386096 284260 386102
rect 284208 386038 284260 386044
rect 284116 385620 284168 385626
rect 284116 385562 284168 385568
rect 284024 384940 284076 384946
rect 284024 384882 284076 384888
rect 283932 382016 283984 382022
rect 283932 381958 283984 381964
rect 283840 333600 283892 333606
rect 283840 333542 283892 333548
rect 282736 331832 282788 331838
rect 282736 331774 282788 331780
rect 282748 326466 282776 331774
rect 282736 326460 282788 326466
rect 282736 326402 282788 326408
rect 282644 326392 282696 326398
rect 282644 326334 282696 326340
rect 282736 326324 282788 326330
rect 282736 326266 282788 326272
rect 282552 320884 282604 320890
rect 282552 320826 282604 320832
rect 282460 320476 282512 320482
rect 282460 320418 282512 320424
rect 282276 320408 282328 320414
rect 282276 320350 282328 320356
rect 282748 320346 282776 326266
rect 285600 322250 285628 650150
rect 299492 647290 299520 656814
rect 311990 650992 312046 651001
rect 311820 650950 311990 650978
rect 311820 650865 311848 650950
rect 311990 650927 312046 650936
rect 309046 650856 309102 650865
rect 309046 650791 309102 650800
rect 311806 650856 311862 650865
rect 311806 650791 311862 650800
rect 309060 650457 309088 650791
rect 340786 650720 340842 650729
rect 364536 650690 364564 659654
rect 378140 653404 378192 653410
rect 378140 653346 378192 653352
rect 378152 652905 378180 653346
rect 378138 652896 378194 652905
rect 378138 652831 378140 652840
rect 378192 652831 378194 652840
rect 383474 652896 383530 652905
rect 383474 652831 383476 652840
rect 378140 652802 378192 652808
rect 383528 652831 383530 652840
rect 387800 652860 387852 652866
rect 383476 652802 383528 652808
rect 387800 652802 387852 652808
rect 378152 652771 378180 652802
rect 386326 651400 386382 651409
rect 386326 651335 386382 651344
rect 370410 651128 370466 651137
rect 370410 651063 370466 651072
rect 367098 650856 367154 650865
rect 370424 650826 370452 651063
rect 386340 651001 386368 651335
rect 386326 650992 386382 651001
rect 386326 650927 386382 650936
rect 367098 650791 367100 650800
rect 367152 650791 367154 650800
rect 370412 650820 370464 650826
rect 367100 650762 367152 650768
rect 370412 650762 370464 650768
rect 340786 650655 340842 650664
rect 364524 650684 364576 650690
rect 340800 650622 340828 650655
rect 364524 650626 364576 650632
rect 340788 650616 340840 650622
rect 321466 650584 321522 650593
rect 321650 650584 321706 650593
rect 321522 650542 321650 650570
rect 321466 650519 321522 650528
rect 347688 650616 347740 650622
rect 340788 650558 340840 650564
rect 347686 650584 347688 650593
rect 347740 650584 347742 650593
rect 321650 650519 321706 650528
rect 347686 650519 347742 650528
rect 309046 650448 309102 650457
rect 309046 650383 309102 650392
rect 386420 650344 386472 650350
rect 386420 650286 386472 650292
rect 386432 649913 386460 650286
rect 386418 649904 386474 649913
rect 386418 649839 386474 649848
rect 299480 647284 299532 647290
rect 299480 647226 299532 647232
rect 299664 647284 299716 647290
rect 299664 647226 299716 647232
rect 297364 645924 297416 645930
rect 297364 645866 297416 645872
rect 294604 644496 294656 644502
rect 294604 644438 294656 644444
rect 291844 643136 291896 643142
rect 291844 643078 291896 643084
rect 290464 641776 290516 641782
rect 290464 641718 290516 641724
rect 287704 640348 287756 640354
rect 287704 640290 287756 640296
rect 286324 638988 286376 638994
rect 286324 638930 286376 638936
rect 286336 343534 286364 638930
rect 287152 413432 287204 413438
rect 287152 413374 287204 413380
rect 287060 413228 287112 413234
rect 287060 413170 287112 413176
rect 287072 413030 287100 413170
rect 287164 413098 287192 413374
rect 287152 413092 287204 413098
rect 287152 413034 287204 413040
rect 287060 413024 287112 413030
rect 287060 412966 287112 412972
rect 287716 344554 287744 640290
rect 288532 558204 288584 558210
rect 288532 558146 288584 558152
rect 288440 557864 288492 557870
rect 288544 557818 288572 558146
rect 288492 557812 288572 557818
rect 288440 557806 288572 557812
rect 288348 557796 288400 557802
rect 288452 557790 288572 557806
rect 288348 557738 288400 557744
rect 288360 557598 288388 557738
rect 288348 557592 288400 557598
rect 288348 557534 288400 557540
rect 290476 346390 290504 641718
rect 291856 347682 291884 643078
rect 294616 347750 294644 644438
rect 296536 413432 296588 413438
rect 296536 413374 296588 413380
rect 296548 413098 296576 413374
rect 296628 413228 296680 413234
rect 296628 413170 296680 413176
rect 296536 413092 296588 413098
rect 296536 413034 296588 413040
rect 296640 413030 296668 413170
rect 296628 413024 296680 413030
rect 296628 412966 296680 412972
rect 297376 349110 297404 645866
rect 299676 630766 299704 647226
rect 307114 646368 307170 646377
rect 307114 646303 307170 646312
rect 307128 645930 307156 646303
rect 307116 645924 307168 645930
rect 307116 645866 307168 645872
rect 307114 645008 307170 645017
rect 307114 644943 307170 644952
rect 307128 644502 307156 644943
rect 307116 644496 307168 644502
rect 307116 644438 307168 644444
rect 307114 643512 307170 643521
rect 307114 643447 307170 643456
rect 307128 643142 307156 643447
rect 307116 643136 307168 643142
rect 307116 643078 307168 643084
rect 307666 642152 307722 642161
rect 307666 642087 307722 642096
rect 307680 641782 307708 642087
rect 307668 641776 307720 641782
rect 307668 641718 307720 641724
rect 307666 640520 307722 640529
rect 307666 640455 307722 640464
rect 307680 640354 307708 640455
rect 307668 640348 307720 640354
rect 307668 640290 307720 640296
rect 306654 639432 306710 639441
rect 306654 639367 306710 639376
rect 306668 638994 306696 639367
rect 306656 638988 306708 638994
rect 306656 638930 306708 638936
rect 306838 637936 306894 637945
rect 306838 637871 306894 637880
rect 306852 637634 306880 637871
rect 301504 637628 301556 637634
rect 301504 637570 301556 637576
rect 306840 637628 306892 637634
rect 306840 637570 306892 637576
rect 299664 630760 299716 630766
rect 299664 630702 299716 630708
rect 299756 630760 299808 630766
rect 299756 630702 299808 630708
rect 299768 611386 299796 630702
rect 299572 611380 299624 611386
rect 299572 611322 299624 611328
rect 299756 611380 299808 611386
rect 299756 611322 299808 611328
rect 299584 611266 299612 611322
rect 299584 611238 299704 611266
rect 299676 608598 299704 611238
rect 299572 608592 299624 608598
rect 299572 608534 299624 608540
rect 299664 608592 299716 608598
rect 299664 608534 299716 608540
rect 299584 601730 299612 608534
rect 299572 601724 299624 601730
rect 299572 601666 299624 601672
rect 299848 601724 299900 601730
rect 299848 601666 299900 601672
rect 299860 598942 299888 601666
rect 299664 598936 299716 598942
rect 299664 598878 299716 598884
rect 299848 598936 299900 598942
rect 299848 598878 299900 598884
rect 299676 589393 299704 598878
rect 299662 589384 299718 589393
rect 299662 589319 299718 589328
rect 299938 589384 299994 589393
rect 299938 589319 299994 589328
rect 299952 582486 299980 589319
rect 299940 582480 299992 582486
rect 299940 582422 299992 582428
rect 299848 582344 299900 582350
rect 299848 582286 299900 582292
rect 299860 572642 299888 582286
rect 299676 572614 299888 572642
rect 299676 563122 299704 572614
rect 299584 563094 299704 563122
rect 299584 562986 299612 563094
rect 299584 562958 299704 562986
rect 298008 558204 298060 558210
rect 298008 558146 298060 558152
rect 298020 558006 298048 558146
rect 298008 558000 298060 558006
rect 298008 557942 298060 557948
rect 297456 557864 297508 557870
rect 297456 557806 297508 557812
rect 297364 349104 297416 349110
rect 297364 349046 297416 349052
rect 294604 347744 294656 347750
rect 294604 347686 294656 347692
rect 291844 347676 291896 347682
rect 291844 347618 291896 347624
rect 290464 346384 290516 346390
rect 290464 346326 290516 346332
rect 287704 344548 287756 344554
rect 287704 344490 287756 344496
rect 286324 343528 286376 343534
rect 286324 343470 286376 343476
rect 297468 329730 297496 557806
rect 299676 553466 299704 562958
rect 299676 553438 299796 553466
rect 299768 540734 299796 553438
rect 299756 540728 299808 540734
rect 299756 540670 299808 540676
rect 298744 410780 298796 410786
rect 298744 410722 298796 410728
rect 298756 383654 298784 410722
rect 298744 383648 298796 383654
rect 298744 383590 298796 383596
rect 301516 343602 301544 637570
rect 387812 589665 387840 652802
rect 400862 651128 400918 651137
rect 400862 651063 400918 651072
rect 389178 650992 389234 651001
rect 389234 650950 389312 650978
rect 389178 650927 389234 650936
rect 389284 650865 389312 650950
rect 389270 650856 389326 650865
rect 389270 650791 389326 650800
rect 400876 650593 400904 651063
rect 400862 650584 400918 650593
rect 400862 650519 400918 650528
rect 405738 650584 405794 650593
rect 418250 650584 418306 650593
rect 405738 650519 405740 650528
rect 405792 650519 405794 650528
rect 413376 650548 413428 650554
rect 405740 650490 405792 650496
rect 413376 650490 413428 650496
rect 418080 650542 418250 650570
rect 413388 650185 413416 650490
rect 418080 650321 418108 650542
rect 418250 650519 418306 650528
rect 418066 650312 418122 650321
rect 418066 650247 418122 650256
rect 413374 650176 413430 650185
rect 413374 650111 413430 650120
rect 429488 647290 429516 673406
rect 444286 650856 444342 650865
rect 444286 650791 444342 650800
rect 444300 650593 444328 650791
rect 444286 650584 444342 650593
rect 444286 650519 444342 650528
rect 456708 650480 456760 650486
rect 456706 650448 456708 650457
rect 456760 650448 456762 650457
rect 456706 650383 456762 650392
rect 429384 647284 429436 647290
rect 429384 647226 429436 647232
rect 429476 647284 429528 647290
rect 429476 647226 429528 647232
rect 429396 640422 429424 647226
rect 429384 640416 429436 640422
rect 429384 640358 429436 640364
rect 429476 640416 429528 640422
rect 429476 640358 429528 640364
rect 429488 630698 429516 640358
rect 429292 630692 429344 630698
rect 429292 630634 429344 630640
rect 429476 630692 429528 630698
rect 429476 630634 429528 630640
rect 429304 630578 429332 630634
rect 429304 630550 429424 630578
rect 429396 621058 429424 630550
rect 429396 621030 429516 621058
rect 429488 611386 429516 621030
rect 429292 611380 429344 611386
rect 429292 611322 429344 611328
rect 429476 611380 429528 611386
rect 429476 611322 429528 611328
rect 429304 611266 429332 611322
rect 429304 611238 429424 611266
rect 429396 608598 429424 611238
rect 429292 608592 429344 608598
rect 429292 608534 429344 608540
rect 429384 608592 429436 608598
rect 429384 608534 429436 608540
rect 429304 601730 429332 608534
rect 429292 601724 429344 601730
rect 429292 601666 429344 601672
rect 429568 601724 429620 601730
rect 429568 601666 429620 601672
rect 429580 592074 429608 601666
rect 429568 592068 429620 592074
rect 429568 592010 429620 592016
rect 429660 591932 429712 591938
rect 429660 591874 429712 591880
rect 387798 589656 387854 589665
rect 387798 589591 387854 589600
rect 309784 589348 309836 589354
rect 309784 589290 309836 589296
rect 307022 579728 307078 579737
rect 307022 579663 307078 579672
rect 305642 578368 305698 578377
rect 305642 578303 305698 578312
rect 305656 560930 305684 578303
rect 305644 560924 305696 560930
rect 305644 560866 305696 560872
rect 302240 558204 302292 558210
rect 302240 558146 302292 558152
rect 302148 558000 302200 558006
rect 302148 557942 302200 557948
rect 302160 557802 302188 557942
rect 302252 557802 302280 558146
rect 302884 557932 302936 557938
rect 302884 557874 302936 557880
rect 302148 557796 302200 557802
rect 302148 557738 302200 557744
rect 302240 557796 302292 557802
rect 302240 557738 302292 557744
rect 302148 545488 302200 545494
rect 302146 545456 302148 545465
rect 302200 545456 302202 545465
rect 302146 545391 302202 545400
rect 301504 343596 301556 343602
rect 301504 343538 301556 343544
rect 297456 329724 297508 329730
rect 297456 329666 297508 329672
rect 302896 328438 302924 557874
rect 305656 411942 305684 560866
rect 306472 413432 306524 413438
rect 306472 413374 306524 413380
rect 306380 413228 306432 413234
rect 306380 413170 306432 413176
rect 306392 413030 306420 413170
rect 306484 413098 306512 413374
rect 306472 413092 306524 413098
rect 306472 413034 306524 413040
rect 306380 413024 306432 413030
rect 306380 412966 306432 412972
rect 305644 411936 305696 411942
rect 305644 411878 305696 411884
rect 302884 328432 302936 328438
rect 302884 328374 302936 328380
rect 305656 322930 305684 411878
rect 307036 333946 307064 579663
rect 309796 560250 309824 589290
rect 429672 587874 429700 591874
rect 429580 587846 429700 587874
rect 429580 583098 429608 587846
rect 429292 583092 429344 583098
rect 429292 583034 429344 583040
rect 429568 583092 429620 583098
rect 429568 583034 429620 583040
rect 389178 580952 389234 580961
rect 389178 580887 389234 580896
rect 389192 560250 389220 580887
rect 429304 578270 429332 583034
rect 429292 578264 429344 578270
rect 429292 578206 429344 578212
rect 429384 578264 429436 578270
rect 429384 578206 429436 578212
rect 429396 572626 429424 578206
rect 429384 572620 429436 572626
rect 429384 572562 429436 572568
rect 429660 572620 429712 572626
rect 429660 572562 429712 572568
rect 429672 560318 429700 572562
rect 429476 560312 429528 560318
rect 429476 560254 429528 560260
rect 429660 560312 429712 560318
rect 429660 560254 429712 560260
rect 309784 560244 309836 560250
rect 309784 560186 309836 560192
rect 310428 560244 310480 560250
rect 310428 560186 310480 560192
rect 389180 560244 389232 560250
rect 389180 560186 389232 560192
rect 309046 545592 309102 545601
rect 309046 545527 309102 545536
rect 309060 545494 309088 545527
rect 309048 545488 309100 545494
rect 309048 545430 309100 545436
rect 310440 389842 310468 560186
rect 329102 559872 329158 559881
rect 329102 559807 329158 559816
rect 337750 559872 337806 559881
rect 337750 559807 337806 559816
rect 357714 559872 357770 559881
rect 357714 559807 357770 559816
rect 313370 558920 313426 558929
rect 313370 558855 313426 558864
rect 321558 558920 321614 558929
rect 321558 558855 321614 558864
rect 322938 558920 322994 558929
rect 322938 558855 322994 558864
rect 324318 558920 324374 558929
rect 324318 558855 324374 558864
rect 325698 558920 325754 558929
rect 325698 558855 325754 558864
rect 327078 558920 327134 558929
rect 327078 558855 327134 558864
rect 313384 558210 313412 558855
rect 313372 558204 313424 558210
rect 313372 558146 313424 558152
rect 317418 557968 317474 557977
rect 317418 557903 317420 557912
rect 317472 557903 317474 557912
rect 320178 557968 320234 557977
rect 320178 557903 320234 557912
rect 317420 557874 317472 557880
rect 320192 557870 320220 557903
rect 320180 557864 320232 557870
rect 320180 557806 320232 557812
rect 316038 557560 316094 557569
rect 316038 557495 316094 557504
rect 318798 557560 318854 557569
rect 318798 557495 318854 557504
rect 320270 557560 320326 557569
rect 320270 557495 320326 557504
rect 315856 413432 315908 413438
rect 315856 413374 315908 413380
rect 315868 413098 315896 413374
rect 315948 413228 316000 413234
rect 315948 413170 316000 413176
rect 315856 413092 315908 413098
rect 315856 413034 315908 413040
rect 315960 413030 315988 413170
rect 315948 413024 316000 413030
rect 315948 412966 316000 412972
rect 311164 411868 311216 411874
rect 311164 411810 311216 411816
rect 311176 404326 311204 411810
rect 311164 404320 311216 404326
rect 311164 404262 311216 404268
rect 310428 389836 310480 389842
rect 310428 389778 310480 389784
rect 316052 342242 316080 557495
rect 318248 413568 318300 413574
rect 318248 413510 318300 413516
rect 318156 413432 318208 413438
rect 318156 413374 318208 413380
rect 318064 413228 318116 413234
rect 318064 413170 318116 413176
rect 316040 342236 316092 342242
rect 316040 342178 316092 342184
rect 307024 333940 307076 333946
rect 307024 333882 307076 333888
rect 318076 324290 318104 413170
rect 318168 325650 318196 413374
rect 318260 327078 318288 413510
rect 318812 329798 318840 557495
rect 320284 331226 320312 557495
rect 321468 545352 321520 545358
rect 321466 545320 321468 545329
rect 321520 545320 321522 545329
rect 321466 545255 321522 545264
rect 321572 366994 321600 558855
rect 322202 558784 322258 558793
rect 322202 558719 322258 558728
rect 322216 557870 322244 558719
rect 322204 557864 322256 557870
rect 322204 557806 322256 557812
rect 321560 366988 321612 366994
rect 321560 366930 321612 366936
rect 322216 358766 322244 557806
rect 322952 367062 322980 558855
rect 323582 558784 323638 558793
rect 323582 558719 323638 558728
rect 323596 557938 323624 558719
rect 323584 557932 323636 557938
rect 323584 557874 323636 557880
rect 322940 367056 322992 367062
rect 322940 366998 322992 367004
rect 323596 360126 323624 557874
rect 324332 368490 324360 558855
rect 324962 558784 325018 558793
rect 324962 558719 325018 558728
rect 324976 557802 325004 558719
rect 324964 557796 325016 557802
rect 324964 557738 325016 557744
rect 324320 368484 324372 368490
rect 324320 368426 324372 368432
rect 324976 360194 325004 557738
rect 325712 369850 325740 558855
rect 326342 558784 326398 558793
rect 326342 558719 326398 558728
rect 326356 558006 326384 558719
rect 326344 558000 326396 558006
rect 326344 557942 326396 557948
rect 325884 413840 325936 413846
rect 325884 413782 325936 413788
rect 325792 413772 325844 413778
rect 325792 413714 325844 413720
rect 325804 413030 325832 413714
rect 325896 413098 325924 413782
rect 325884 413092 325936 413098
rect 325884 413034 325936 413040
rect 325792 413024 325844 413030
rect 325792 412966 325844 412972
rect 325700 369844 325752 369850
rect 325700 369786 325752 369792
rect 326356 361554 326384 557942
rect 327092 371142 327120 558855
rect 328460 558816 328512 558822
rect 327722 558784 327778 558793
rect 327722 558719 327778 558728
rect 328458 558784 328460 558793
rect 328512 558784 328514 558793
rect 328458 558719 328514 558728
rect 328552 558748 328604 558754
rect 327736 557598 327764 558719
rect 328552 558690 328604 558696
rect 328564 558532 328592 558690
rect 328472 558521 328592 558532
rect 328458 558512 328592 558521
rect 328514 558504 328592 558512
rect 328458 558447 328514 558456
rect 327724 557592 327776 557598
rect 327724 557534 327776 557540
rect 327080 371136 327132 371142
rect 327080 371078 327132 371084
rect 327736 362846 327764 557534
rect 328458 557152 328514 557161
rect 328458 557087 328514 557096
rect 328366 545456 328422 545465
rect 328366 545391 328422 545400
rect 328380 545358 328408 545391
rect 328368 545352 328420 545358
rect 328368 545294 328420 545300
rect 328472 371210 328500 557087
rect 328460 371204 328512 371210
rect 328460 371146 328512 371152
rect 329116 362914 329144 559807
rect 329286 558920 329342 558929
rect 329286 558855 329342 558864
rect 329838 558920 329894 558929
rect 329838 558855 329894 558864
rect 330482 558920 330538 558929
rect 330482 558855 330538 558864
rect 331218 558920 331274 558929
rect 331218 558855 331274 558864
rect 332598 558920 332654 558929
rect 332598 558855 332654 558864
rect 333978 558920 334034 558929
rect 333978 558855 334034 558864
rect 335358 558920 335414 558929
rect 336738 558920 336794 558929
rect 335358 558855 335414 558864
rect 335452 558884 335504 558890
rect 329300 558414 329328 558855
rect 329288 558408 329340 558414
rect 329288 558350 329340 558356
rect 329300 364342 329328 558350
rect 329852 372570 329880 558855
rect 329930 558784 329986 558793
rect 329930 558719 329986 558728
rect 329944 373930 329972 558719
rect 330496 558550 330524 558855
rect 330484 558544 330536 558550
rect 330484 558486 330536 558492
rect 329932 373924 329984 373930
rect 329932 373866 329984 373872
rect 329840 372564 329892 372570
rect 329840 372506 329892 372512
rect 330496 365702 330524 558486
rect 331232 373998 331260 558855
rect 331770 558784 331826 558793
rect 331770 558719 331826 558728
rect 331784 558278 331812 558719
rect 331312 558272 331364 558278
rect 331312 558214 331364 558220
rect 331772 558272 331824 558278
rect 331772 558214 331824 558220
rect 331324 557870 331352 558214
rect 331312 557864 331364 557870
rect 331312 557806 331364 557812
rect 332612 375358 332640 558855
rect 332690 558784 332746 558793
rect 332690 558719 332746 558728
rect 332704 558346 332732 558719
rect 332692 558340 332744 558346
rect 332692 558282 332744 558288
rect 332704 557938 332732 558282
rect 332692 557932 332744 557938
rect 332692 557874 332744 557880
rect 333992 376718 334020 558855
rect 334070 558784 334126 558793
rect 334070 558719 334126 558728
rect 334084 558210 334112 558719
rect 334072 558204 334124 558210
rect 334072 558146 334124 558152
rect 334084 557802 334112 558146
rect 334072 557796 334124 557802
rect 334072 557738 334124 557744
rect 335176 413840 335228 413846
rect 335176 413782 335228 413788
rect 335188 413098 335216 413782
rect 335268 413772 335320 413778
rect 335268 413714 335320 413720
rect 335176 413092 335228 413098
rect 335176 413034 335228 413040
rect 335280 413030 335308 413714
rect 335268 413024 335320 413030
rect 335268 412966 335320 412972
rect 335372 378078 335400 558855
rect 336738 558855 336794 558864
rect 335452 558826 335504 558832
rect 335464 558793 335492 558826
rect 335450 558784 335506 558793
rect 335450 558719 335506 558728
rect 336462 558784 336518 558793
rect 336462 558719 336518 558728
rect 335464 558006 335492 558719
rect 336476 558618 336504 558719
rect 336464 558612 336516 558618
rect 336464 558554 336516 558560
rect 335452 558000 335504 558006
rect 335452 557942 335504 557948
rect 336476 557598 336504 558554
rect 336464 557592 336516 557598
rect 336464 557534 336516 557540
rect 336752 378146 336780 558855
rect 337764 558482 337792 559807
rect 348146 559328 348202 559337
rect 348146 559263 348202 559272
rect 348054 559192 348110 559201
rect 348054 559127 348110 559136
rect 338118 558920 338174 558929
rect 338118 558855 338174 558864
rect 339498 558920 339554 558929
rect 339498 558855 339554 558864
rect 341246 558920 341302 558929
rect 341246 558855 341302 558864
rect 342534 558920 342590 558929
rect 342534 558855 342590 558864
rect 343638 558920 343694 558929
rect 343638 558855 343694 558864
rect 344834 558920 344890 558929
rect 344834 558855 344836 558864
rect 338028 558816 338080 558822
rect 338026 558784 338028 558793
rect 338080 558784 338082 558793
rect 337936 558748 337988 558754
rect 338026 558719 338082 558728
rect 337936 558690 337988 558696
rect 337948 558532 337976 558690
rect 337948 558521 338068 558532
rect 337948 558512 338082 558521
rect 337948 558504 338026 558512
rect 337752 558476 337804 558482
rect 338026 558447 338082 558456
rect 337752 558418 337804 558424
rect 336830 557968 336886 557977
rect 336830 557903 336886 557912
rect 336844 379506 336872 557903
rect 338026 389872 338082 389881
rect 338026 389807 338028 389816
rect 338080 389807 338082 389816
rect 338028 389778 338080 389784
rect 337382 381304 337438 381313
rect 337382 381239 337438 381248
rect 336832 379500 336884 379506
rect 336832 379442 336884 379448
rect 336740 378140 336792 378146
rect 336740 378082 336792 378088
rect 335360 378072 335412 378078
rect 335360 378014 335412 378020
rect 333980 376712 334032 376718
rect 333980 376654 334032 376660
rect 332600 375352 332652 375358
rect 332600 375294 332652 375300
rect 331220 373992 331272 373998
rect 331220 373934 331272 373940
rect 330484 365696 330536 365702
rect 330484 365638 330536 365644
rect 329288 364336 329340 364342
rect 329288 364278 329340 364284
rect 329104 362908 329156 362914
rect 329104 362850 329156 362856
rect 327724 362840 327776 362846
rect 327724 362782 327776 362788
rect 326344 361548 326396 361554
rect 326344 361490 326396 361496
rect 324964 360188 325016 360194
rect 324964 360130 325016 360136
rect 323584 360120 323636 360126
rect 323584 360062 323636 360068
rect 322204 358760 322256 358766
rect 322204 358702 322256 358708
rect 320272 331220 320324 331226
rect 320272 331162 320324 331168
rect 318800 329792 318852 329798
rect 318800 329734 318852 329740
rect 318248 327072 318300 327078
rect 318248 327014 318300 327020
rect 318156 325644 318208 325650
rect 318156 325586 318208 325592
rect 318064 324284 318116 324290
rect 318064 324226 318116 324232
rect 305644 322924 305696 322930
rect 305644 322866 305696 322872
rect 284300 322244 284352 322250
rect 284300 322186 284352 322192
rect 285588 322244 285640 322250
rect 285588 322186 285640 322192
rect 284312 321570 284340 322186
rect 282828 321564 282880 321570
rect 282828 321506 282880 321512
rect 284300 321564 284352 321570
rect 284300 321506 284352 321512
rect 282840 321473 282868 321506
rect 282826 321464 282882 321473
rect 282826 321399 282882 321408
rect 337396 321026 337424 381239
rect 338132 380866 338160 558855
rect 339038 558784 339094 558793
rect 339038 558719 339094 558728
rect 339052 558414 339080 558719
rect 339040 558408 339092 558414
rect 339040 558350 339092 558356
rect 339512 382226 339540 558855
rect 339866 558784 339922 558793
rect 339866 558719 339922 558728
rect 339880 558550 339908 558719
rect 339868 558544 339920 558550
rect 339868 558486 339920 558492
rect 341260 558278 341288 558855
rect 342548 558346 342576 558855
rect 342536 558340 342588 558346
rect 342536 558282 342588 558288
rect 341248 558272 341300 558278
rect 341248 558214 341300 558220
rect 343652 558210 343680 558855
rect 344888 558855 344890 558864
rect 345754 558920 345810 558929
rect 345754 558855 345810 558864
rect 346858 558920 346914 558929
rect 346858 558855 346914 558864
rect 344836 558826 344888 558832
rect 344848 558686 344876 558826
rect 344836 558680 344888 558686
rect 344836 558622 344888 558628
rect 345768 558618 345796 558855
rect 345756 558612 345808 558618
rect 345756 558554 345808 558560
rect 345662 558512 345718 558521
rect 346872 558482 346900 558855
rect 348068 558657 348096 559127
rect 348054 558648 348110 558657
rect 348054 558583 348110 558592
rect 345662 558447 345718 558456
rect 346860 558476 346912 558482
rect 343640 558204 343692 558210
rect 343640 558146 343692 558152
rect 345676 558113 345704 558447
rect 346860 558418 346912 558424
rect 348160 558346 348188 559263
rect 348238 558920 348294 558929
rect 348238 558855 348294 558864
rect 349526 558920 349582 558929
rect 349526 558855 349582 558864
rect 351734 558920 351790 558929
rect 351734 558855 351790 558864
rect 348252 558414 348280 558855
rect 349540 558550 349568 558855
rect 349528 558544 349580 558550
rect 349528 558486 349580 558492
rect 350538 558512 350594 558521
rect 350538 558447 350594 558456
rect 348240 558408 348292 558414
rect 348240 558350 348292 558356
rect 348148 558340 348200 558346
rect 348148 558282 348200 558288
rect 350552 558278 350580 558447
rect 350540 558272 350592 558278
rect 351748 558249 351776 558855
rect 353298 558784 353354 558793
rect 353298 558719 353354 558728
rect 354678 558784 354734 558793
rect 354678 558719 354734 558728
rect 356058 558784 356114 558793
rect 356058 558719 356114 558728
rect 353312 558686 353340 558719
rect 353300 558680 353352 558686
rect 353300 558622 353352 558628
rect 354692 558618 354720 558719
rect 354680 558612 354732 558618
rect 354680 558554 354732 558560
rect 356072 558482 356100 558719
rect 357728 558550 357756 559807
rect 357716 558544 357768 558550
rect 357438 558512 357494 558521
rect 356060 558476 356112 558482
rect 357716 558486 357768 558492
rect 357438 558447 357494 558456
rect 356060 558418 356112 558424
rect 357452 558414 357480 558447
rect 357440 558408 357492 558414
rect 357440 558350 357492 558356
rect 350540 558214 350592 558220
rect 351734 558240 351790 558249
rect 351734 558175 351790 558184
rect 351918 558240 351974 558249
rect 351918 558175 351920 558184
rect 351972 558175 351974 558184
rect 354678 558240 354734 558249
rect 354678 558175 354734 558184
rect 351920 558146 351972 558152
rect 354692 558142 354720 558175
rect 354680 558136 354732 558142
rect 345662 558104 345718 558113
rect 345662 558039 345718 558048
rect 351918 558104 351974 558113
rect 354680 558078 354732 558084
rect 351918 558039 351974 558048
rect 351932 557734 351960 558039
rect 353298 557968 353354 557977
rect 353298 557903 353354 557912
rect 351920 557728 351972 557734
rect 343730 557696 343786 557705
rect 351920 557670 351972 557676
rect 353312 557666 353340 557903
rect 343730 557631 343786 557640
rect 353300 557660 353352 557666
rect 340878 557560 340934 557569
rect 340878 557495 340934 557504
rect 342258 557560 342314 557569
rect 342258 557495 342314 557504
rect 343638 557560 343694 557569
rect 343638 557495 343694 557504
rect 340892 410718 340920 557495
rect 342272 410786 342300 557495
rect 343652 412350 343680 557495
rect 343744 412418 343772 557631
rect 353300 557602 353352 557608
rect 345018 557560 345074 557569
rect 345018 557495 345074 557504
rect 346398 557560 346454 557569
rect 346398 557495 346454 557504
rect 347778 557560 347834 557569
rect 347778 557495 347834 557504
rect 349158 557560 349214 557569
rect 349158 557495 349214 557504
rect 350630 557560 350686 557569
rect 350630 557495 350686 557504
rect 343732 412412 343784 412418
rect 343732 412354 343784 412360
rect 343640 412344 343692 412350
rect 343640 412286 343692 412292
rect 345032 412282 345060 557495
rect 345204 413840 345256 413846
rect 345204 413782 345256 413788
rect 345112 413772 345164 413778
rect 345112 413714 345164 413720
rect 345124 413030 345152 413714
rect 345216 413098 345244 413782
rect 345204 413092 345256 413098
rect 345204 413034 345256 413040
rect 345112 413024 345164 413030
rect 345112 412966 345164 412972
rect 345020 412276 345072 412282
rect 345020 412218 345072 412224
rect 346412 412214 346440 557495
rect 347686 545456 347742 545465
rect 347686 545391 347742 545400
rect 347700 545329 347728 545391
rect 347686 545320 347742 545329
rect 347686 545255 347742 545264
rect 346400 412208 346452 412214
rect 346400 412150 346452 412156
rect 347792 412146 347820 557495
rect 347780 412140 347832 412146
rect 347780 412082 347832 412088
rect 349172 412078 349200 557495
rect 349160 412072 349212 412078
rect 349160 412014 349212 412020
rect 350644 412010 350672 557495
rect 429488 550610 429516 560254
rect 429396 550582 429516 550610
rect 371882 545592 371938 545601
rect 371882 545527 371938 545536
rect 367006 545320 367062 545329
rect 367006 545255 367062 545264
rect 367020 544921 367048 545255
rect 371896 545193 371924 545527
rect 371882 545184 371938 545193
rect 371882 545119 371938 545128
rect 367006 544912 367062 544921
rect 367006 544847 367062 544856
rect 429396 543794 429424 550582
rect 429384 543788 429436 543794
rect 429384 543730 429436 543736
rect 429476 543720 429528 543726
rect 429476 543662 429528 543668
rect 429488 541006 429516 543662
rect 429384 541000 429436 541006
rect 429384 540942 429436 540948
rect 429476 541000 429528 541006
rect 429476 540942 429528 540948
rect 429396 540666 429424 540942
rect 429384 540660 429436 540666
rect 429384 540602 429436 540608
rect 462332 540598 462360 703520
rect 478524 700398 478552 703520
rect 494808 703474 494836 703520
rect 494808 703446 494928 703474
rect 478512 700392 478564 700398
rect 478512 700334 478564 700340
rect 494900 692850 494928 703446
rect 527192 700330 527220 703520
rect 543476 700369 543504 703520
rect 543462 700360 543518 700369
rect 527180 700324 527232 700330
rect 543462 700295 543518 700304
rect 527180 700266 527232 700272
rect 553306 697368 553362 697377
rect 553490 697368 553546 697377
rect 553362 697326 553490 697354
rect 553306 697303 553362 697312
rect 553490 697303 553546 697312
rect 540978 697232 541034 697241
rect 540978 697167 540980 697176
rect 541032 697167 541034 697176
rect 548616 697196 548668 697202
rect 540980 697138 541032 697144
rect 548616 697138 548668 697144
rect 548628 696969 548656 697138
rect 548614 696960 548670 696969
rect 548614 696895 548670 696904
rect 494060 692844 494112 692850
rect 494060 692786 494112 692792
rect 494888 692844 494940 692850
rect 494888 692786 494940 692792
rect 494072 683074 494100 692786
rect 553306 686352 553362 686361
rect 553490 686352 553546 686361
rect 553362 686310 553490 686338
rect 553306 686287 553362 686296
rect 553490 686287 553546 686296
rect 540978 686216 541034 686225
rect 540978 686151 540980 686160
rect 541032 686151 541034 686160
rect 548616 686180 548668 686186
rect 540980 686122 541032 686128
rect 548616 686122 548668 686128
rect 548628 685953 548656 686122
rect 548614 685944 548670 685953
rect 548614 685879 548670 685888
rect 559668 684554 559696 703520
rect 560298 697368 560354 697377
rect 560298 697303 560300 697312
rect 560352 697303 560354 697312
rect 565176 697332 565228 697338
rect 560300 697274 560352 697280
rect 565176 697274 565228 697280
rect 565188 697241 565216 697274
rect 565174 697232 565230 697241
rect 572718 697232 572774 697241
rect 565174 697167 565230 697176
rect 572640 697190 572718 697218
rect 572640 697105 572668 697190
rect 572718 697167 572774 697176
rect 572626 697096 572682 697105
rect 572626 697031 572682 697040
rect 560298 686352 560354 686361
rect 560298 686287 560300 686296
rect 560352 686287 560354 686296
rect 565176 686316 565228 686322
rect 560300 686258 560352 686264
rect 565176 686258 565228 686264
rect 565188 686225 565216 686258
rect 565174 686216 565230 686225
rect 572718 686216 572774 686225
rect 565174 686151 565230 686160
rect 572640 686174 572718 686202
rect 572640 686089 572668 686174
rect 572718 686151 572774 686160
rect 572626 686080 572682 686089
rect 572626 686015 572682 686024
rect 559012 684548 559064 684554
rect 559012 684490 559064 684496
rect 559656 684548 559708 684554
rect 559656 684490 559708 684496
rect 559024 684457 559052 684490
rect 559010 684448 559066 684457
rect 559010 684383 559066 684392
rect 559010 684312 559066 684321
rect 559010 684247 559066 684256
rect 494072 683046 494284 683074
rect 494256 673538 494284 683046
rect 559024 674898 559052 684247
rect 559012 674892 559064 674898
rect 559012 674834 559064 674840
rect 559380 674892 559432 674898
rect 559380 674834 559432 674840
rect 553398 673976 553454 673985
rect 553398 673911 553454 673920
rect 540978 673840 541034 673849
rect 540978 673775 540980 673784
rect 541032 673775 541034 673784
rect 548616 673804 548668 673810
rect 540980 673746 541032 673752
rect 548616 673746 548668 673752
rect 548628 673577 548656 673746
rect 548614 673568 548670 673577
rect 494060 673532 494112 673538
rect 494060 673474 494112 673480
rect 494244 673532 494296 673538
rect 548614 673503 548670 673512
rect 553306 673568 553362 673577
rect 553412 673554 553440 673911
rect 553362 673526 553440 673554
rect 553306 673503 553362 673512
rect 494244 673474 494296 673480
rect 494072 669322 494100 673474
rect 494060 669316 494112 669322
rect 494060 669258 494112 669264
rect 494244 669316 494296 669322
rect 494244 669258 494296 669264
rect 494256 666534 494284 669258
rect 493968 666528 494020 666534
rect 493968 666470 494020 666476
rect 494244 666528 494296 666534
rect 494244 666470 494296 666476
rect 493980 656946 494008 666470
rect 559392 661774 559420 674834
rect 560298 673976 560354 673985
rect 560298 673911 560300 673920
rect 560352 673911 560354 673920
rect 565176 673940 565228 673946
rect 560300 673882 560352 673888
rect 565176 673882 565228 673888
rect 565188 673849 565216 673882
rect 565174 673840 565230 673849
rect 572718 673840 572774 673849
rect 565174 673775 565230 673784
rect 572640 673798 572718 673826
rect 572640 673713 572668 673798
rect 572718 673775 572774 673784
rect 572626 673704 572682 673713
rect 572626 673639 572682 673648
rect 559104 661768 559156 661774
rect 559104 661710 559156 661716
rect 559380 661768 559432 661774
rect 559380 661710 559432 661716
rect 559116 656946 559144 661710
rect 493968 656940 494020 656946
rect 493968 656882 494020 656888
rect 494152 656940 494204 656946
rect 494152 656882 494204 656888
rect 559104 656940 559156 656946
rect 559104 656882 559156 656888
rect 559196 656940 559248 656946
rect 559196 656882 559248 656888
rect 463606 650584 463662 650593
rect 463606 650519 463662 650528
rect 482926 650584 482982 650593
rect 482926 650519 482982 650528
rect 463620 650486 463648 650519
rect 482940 650486 482968 650519
rect 463608 650480 463660 650486
rect 476028 650480 476080 650486
rect 463608 650422 463660 650428
rect 476026 650448 476028 650457
rect 482928 650480 482980 650486
rect 476080 650448 476082 650457
rect 482928 650422 482980 650428
rect 476026 650383 476082 650392
rect 494164 650026 494192 656882
rect 502246 650584 502302 650593
rect 502246 650519 502302 650528
rect 521566 650584 521622 650593
rect 540886 650584 540942 650593
rect 521566 650519 521622 650528
rect 533988 650548 534040 650554
rect 502260 650486 502288 650519
rect 521580 650486 521608 650519
rect 540886 650519 540888 650528
rect 533988 650490 534040 650496
rect 540940 650519 540942 650528
rect 540888 650490 540940 650496
rect 495348 650480 495400 650486
rect 495346 650448 495348 650457
rect 502248 650480 502300 650486
rect 495400 650448 495402 650457
rect 514668 650480 514720 650486
rect 502248 650422 502300 650428
rect 514666 650448 514668 650457
rect 521568 650480 521620 650486
rect 514720 650448 514722 650457
rect 495346 650383 495402 650392
rect 534000 650457 534028 650490
rect 521568 650422 521620 650428
rect 533986 650448 534042 650457
rect 514666 650383 514722 650392
rect 533986 650383 534042 650392
rect 494072 649998 494192 650026
rect 494072 644450 494100 649998
rect 559208 647290 559236 656882
rect 583390 651128 583446 651137
rect 583390 651063 583446 651072
rect 583404 650865 583432 651063
rect 563150 650856 563206 650865
rect 563150 650791 563206 650800
rect 583390 650856 583446 650865
rect 583390 650791 583446 650800
rect 563164 650622 563192 650791
rect 572628 650752 572680 650758
rect 572626 650720 572628 650729
rect 579528 650752 579580 650758
rect 572680 650720 572682 650729
rect 572626 650655 572682 650664
rect 579526 650720 579528 650729
rect 579580 650720 579582 650729
rect 579526 650655 579582 650664
rect 560300 650616 560352 650622
rect 560298 650584 560300 650593
rect 563152 650616 563204 650622
rect 560352 650584 560354 650593
rect 563152 650558 563204 650564
rect 560298 650519 560354 650528
rect 559104 647284 559156 647290
rect 559104 647226 559156 647232
rect 559196 647284 559248 647290
rect 559196 647226 559248 647232
rect 494072 644422 494284 644450
rect 494256 634846 494284 644422
rect 559116 640422 559144 647226
rect 559104 640416 559156 640422
rect 559104 640358 559156 640364
rect 559196 640416 559248 640422
rect 559196 640358 559248 640364
rect 494060 634840 494112 634846
rect 494060 634782 494112 634788
rect 494244 634840 494296 634846
rect 494244 634782 494296 634788
rect 494072 625138 494100 634782
rect 559208 630698 559236 640358
rect 580262 639432 580318 639441
rect 580262 639367 580318 639376
rect 559012 630692 559064 630698
rect 559012 630634 559064 630640
rect 559196 630692 559248 630698
rect 559196 630634 559248 630640
rect 559024 630578 559052 630634
rect 559024 630550 559144 630578
rect 494072 625110 494284 625138
rect 494256 615534 494284 625110
rect 559116 621058 559144 630550
rect 559116 621030 559236 621058
rect 494060 615528 494112 615534
rect 494060 615470 494112 615476
rect 494244 615528 494296 615534
rect 494244 615470 494296 615476
rect 494072 605826 494100 615470
rect 559208 611386 559236 621030
rect 559012 611380 559064 611386
rect 559012 611322 559064 611328
rect 559196 611380 559248 611386
rect 559196 611322 559248 611328
rect 559024 611266 559052 611322
rect 559024 611238 559144 611266
rect 559116 608598 559144 611238
rect 559012 608592 559064 608598
rect 559012 608534 559064 608540
rect 559104 608592 559156 608598
rect 559104 608534 559156 608540
rect 494072 605798 494284 605826
rect 494256 596222 494284 605798
rect 559024 601730 559052 608534
rect 559012 601724 559064 601730
rect 559012 601666 559064 601672
rect 559288 601724 559340 601730
rect 559288 601666 559340 601672
rect 559300 598942 559328 601666
rect 559104 598936 559156 598942
rect 559104 598878 559156 598884
rect 559288 598936 559340 598942
rect 559288 598878 559340 598884
rect 494060 596216 494112 596222
rect 494244 596216 494296 596222
rect 494112 596164 494192 596170
rect 494060 596158 494192 596164
rect 494244 596158 494296 596164
rect 494072 596142 494192 596158
rect 494164 596034 494192 596142
rect 494164 596006 494284 596034
rect 494256 591954 494284 596006
rect 494164 591926 494284 591954
rect 494164 589286 494192 591926
rect 559116 589354 559144 598878
rect 559104 589348 559156 589354
rect 559104 589290 559156 589296
rect 559380 589348 559432 589354
rect 559380 589290 559432 589296
rect 493876 589280 493928 589286
rect 493876 589222 493928 589228
rect 494152 589280 494204 589286
rect 494152 589222 494204 589228
rect 493888 579698 493916 589222
rect 559392 582486 559420 589290
rect 559380 582480 559432 582486
rect 559380 582422 559432 582428
rect 559288 582344 559340 582350
rect 559288 582286 559340 582292
rect 493876 579692 493928 579698
rect 493876 579634 493928 579640
rect 494060 579692 494112 579698
rect 494060 579634 494112 579640
rect 494072 572642 494100 579634
rect 559300 572642 559328 582286
rect 494072 572614 494192 572642
rect 494164 569906 494192 572614
rect 559116 572614 559328 572642
rect 494152 569900 494204 569906
rect 494152 569842 494204 569848
rect 494336 569900 494388 569906
rect 494336 569842 494388 569848
rect 494348 563242 494376 569842
rect 494336 563236 494388 563242
rect 494336 563178 494388 563184
rect 494336 563100 494388 563106
rect 494336 563042 494388 563048
rect 494348 560266 494376 563042
rect 559116 560318 559144 572614
rect 559012 560312 559064 560318
rect 494348 560238 494560 560266
rect 559012 560254 559064 560260
rect 559104 560312 559156 560318
rect 559104 560254 559156 560260
rect 494532 553330 494560 560238
rect 494440 553302 494560 553330
rect 559024 553330 559052 560254
rect 580170 557288 580226 557297
rect 580170 557223 580226 557232
rect 580184 556238 580212 557223
rect 580172 556232 580224 556238
rect 580172 556174 580224 556180
rect 559024 553302 559144 553330
rect 494440 550610 494468 553302
rect 494440 550582 494652 550610
rect 494624 549273 494652 550582
rect 491758 549264 491814 549273
rect 491758 549199 491814 549208
rect 494610 549264 494666 549273
rect 494610 549199 494666 549208
rect 483018 545456 483074 545465
rect 483018 545391 483020 545400
rect 483072 545391 483074 545400
rect 485872 545420 485924 545426
rect 483020 545362 483072 545368
rect 485872 545362 485924 545368
rect 485884 545193 485912 545362
rect 485870 545184 485926 545193
rect 485870 545119 485926 545128
rect 462320 540592 462372 540598
rect 462320 540534 462372 540540
rect 491772 540530 491800 549199
rect 553306 545592 553362 545601
rect 553490 545592 553546 545601
rect 553362 545550 553490 545578
rect 553306 545527 553362 545536
rect 553490 545527 553546 545536
rect 540978 545456 541034 545465
rect 540978 545391 540980 545400
rect 541032 545391 541034 545400
rect 548616 545420 548668 545426
rect 540980 545362 541032 545368
rect 548616 545362 548668 545368
rect 548628 545193 548656 545362
rect 548614 545184 548670 545193
rect 548614 545119 548670 545128
rect 559116 543810 559144 553302
rect 560298 545592 560354 545601
rect 579526 545592 579582 545601
rect 560298 545527 560300 545536
rect 560352 545527 560354 545536
rect 563152 545556 563204 545562
rect 560300 545498 560352 545504
rect 579526 545527 579582 545536
rect 563152 545498 563204 545504
rect 563164 545329 563192 545498
rect 579540 545494 579568 545527
rect 572628 545488 572680 545494
rect 572626 545456 572628 545465
rect 579528 545488 579580 545494
rect 572680 545456 572682 545465
rect 579528 545430 579580 545436
rect 572626 545391 572682 545400
rect 563150 545320 563206 545329
rect 563150 545255 563206 545264
rect 559116 543782 559236 543810
rect 491760 540524 491812 540530
rect 491760 540466 491812 540472
rect 559208 540433 559236 543782
rect 559194 540424 559250 540433
rect 559194 540359 559250 540368
rect 580276 540326 580304 639367
rect 580354 627736 580410 627745
rect 580354 627671 580410 627680
rect 580368 540462 580396 627671
rect 580446 604208 580502 604217
rect 580446 604143 580502 604152
rect 580356 540456 580408 540462
rect 580356 540398 580408 540404
rect 580264 540320 580316 540326
rect 580264 540262 580316 540268
rect 580460 540258 580488 604143
rect 580630 592512 580686 592521
rect 580630 592447 580686 592456
rect 580644 540297 580672 592447
rect 580722 580816 580778 580825
rect 580722 580751 580778 580760
rect 580736 540394 580764 580751
rect 580724 540388 580776 540394
rect 580724 540330 580776 540336
rect 580630 540288 580686 540297
rect 580448 540252 580500 540258
rect 580630 540223 580686 540232
rect 580448 540194 580500 540200
rect 580908 539776 580960 539782
rect 580908 539718 580960 539724
rect 580540 539708 580592 539714
rect 580540 539650 580592 539656
rect 580264 539232 580316 539238
rect 580264 539174 580316 539180
rect 580276 498681 580304 539174
rect 580262 498672 580318 498681
rect 580262 498607 580318 498616
rect 580552 486849 580580 539650
rect 580816 539640 580868 539646
rect 580816 539582 580868 539588
rect 580828 510377 580856 539582
rect 580920 533905 580948 539718
rect 580906 533896 580962 533905
rect 580906 533831 580962 533840
rect 580814 510368 580870 510377
rect 580814 510303 580870 510312
rect 580538 486840 580594 486849
rect 580538 486775 580594 486784
rect 580262 463448 580318 463457
rect 580262 463383 580318 463392
rect 367100 429208 367152 429214
rect 367100 429150 367152 429156
rect 367112 413953 367140 429150
rect 368480 427848 368532 427854
rect 368480 427790 368532 427796
rect 368492 413953 368520 427790
rect 369860 426556 369912 426562
rect 369860 426498 369912 426504
rect 369872 413953 369900 426498
rect 371240 426488 371292 426494
rect 371240 426430 371292 426436
rect 371252 413953 371280 426430
rect 372620 425128 372672 425134
rect 372620 425070 372672 425076
rect 372632 413953 372660 425070
rect 374000 423700 374052 423706
rect 374000 423642 374052 423648
rect 374012 413953 374040 423642
rect 374092 422408 374144 422414
rect 374092 422350 374144 422356
rect 367098 413944 367154 413953
rect 367098 413879 367154 413888
rect 368478 413944 368534 413953
rect 368478 413879 368534 413888
rect 369858 413944 369914 413953
rect 369858 413879 369914 413888
rect 371238 413944 371294 413953
rect 371238 413879 371294 413888
rect 372618 413944 372674 413953
rect 372618 413879 372674 413888
rect 373998 413944 374054 413953
rect 373998 413879 374054 413888
rect 354496 413840 354548 413846
rect 374104 413817 374132 422350
rect 375380 422340 375432 422346
rect 375380 422282 375432 422288
rect 375392 413953 375420 422282
rect 376760 420980 376812 420986
rect 376760 420922 376812 420928
rect 376772 413953 376800 420922
rect 378140 419552 378192 419558
rect 378140 419494 378192 419500
rect 378152 413953 378180 419494
rect 379520 418260 379572 418266
rect 379520 418202 379572 418208
rect 379532 413953 379560 418202
rect 380900 418192 380952 418198
rect 380900 418134 380952 418140
rect 380912 413953 380940 418134
rect 382280 416832 382332 416838
rect 382280 416774 382332 416780
rect 382292 413953 382320 416774
rect 382372 415472 382424 415478
rect 382372 415414 382424 415420
rect 375378 413944 375434 413953
rect 375378 413879 375434 413888
rect 376758 413944 376814 413953
rect 376758 413879 376814 413888
rect 378138 413944 378194 413953
rect 378138 413879 378194 413888
rect 379518 413944 379574 413953
rect 379518 413879 379574 413888
rect 380898 413944 380954 413953
rect 380898 413879 380954 413888
rect 382278 413944 382334 413953
rect 382278 413879 382334 413888
rect 378048 413840 378100 413846
rect 354496 413782 354548 413788
rect 374090 413808 374146 413817
rect 354508 413098 354536 413782
rect 354588 413772 354640 413778
rect 354588 413714 354640 413720
rect 369768 413772 369820 413778
rect 382384 413817 382412 415414
rect 383844 414112 383896 414118
rect 383844 414054 383896 414060
rect 383568 413908 383620 413914
rect 383568 413850 383620 413856
rect 378048 413782 378100 413788
rect 382370 413808 382426 413817
rect 374090 413743 374146 413752
rect 369768 413714 369820 413720
rect 354496 413092 354548 413098
rect 354496 413034 354548 413040
rect 354600 413030 354628 413714
rect 368296 413704 368348 413710
rect 368296 413646 368348 413652
rect 368308 413409 368336 413646
rect 368756 413636 368808 413642
rect 368756 413578 368808 413584
rect 368848 413636 368900 413642
rect 368848 413578 368900 413584
rect 368768 413409 368796 413578
rect 368860 413506 368888 413578
rect 368848 413500 368900 413506
rect 368848 413442 368900 413448
rect 368940 413500 368992 413506
rect 368940 413442 368992 413448
rect 368294 413400 368350 413409
rect 368294 413335 368350 413344
rect 368754 413400 368810 413409
rect 368754 413335 368810 413344
rect 368952 413166 368980 413442
rect 369780 413409 369808 413714
rect 378060 413710 378088 413782
rect 378784 413772 378836 413778
rect 382370 413743 382426 413752
rect 378784 413714 378836 413720
rect 378048 413704 378100 413710
rect 378048 413646 378100 413652
rect 369860 413636 369912 413642
rect 369860 413578 369912 413584
rect 369766 413400 369822 413409
rect 369766 413335 369822 413344
rect 369872 413273 369900 413578
rect 372988 413500 373040 413506
rect 372988 413442 373040 413448
rect 371976 413364 372028 413370
rect 371976 413306 372028 413312
rect 369858 413264 369914 413273
rect 369858 413199 369914 413208
rect 368940 413160 368992 413166
rect 371988 413137 372016 413306
rect 373000 413137 373028 413442
rect 378060 413409 378088 413646
rect 378046 413400 378102 413409
rect 378046 413335 378102 413344
rect 378796 413137 378824 413714
rect 379612 413636 379664 413642
rect 379612 413578 379664 413584
rect 379624 413273 379652 413578
rect 382280 413500 382332 413506
rect 382280 413442 382332 413448
rect 381544 413364 381596 413370
rect 381544 413306 381596 413312
rect 379610 413264 379666 413273
rect 379610 413199 379666 413208
rect 381556 413137 381584 413306
rect 382292 413166 382320 413442
rect 382280 413160 382332 413166
rect 368940 413102 368992 413108
rect 371974 413128 372030 413137
rect 368848 413092 368900 413098
rect 371974 413063 372030 413072
rect 372986 413128 373042 413137
rect 378782 413128 378838 413137
rect 372986 413063 373042 413072
rect 375472 413092 375524 413098
rect 368848 413034 368900 413040
rect 378782 413063 378838 413072
rect 381542 413128 381598 413137
rect 381542 413063 381598 413072
rect 382278 413128 382280 413137
rect 382332 413128 382334 413137
rect 382278 413063 382334 413072
rect 375472 413034 375524 413040
rect 354588 413024 354640 413030
rect 354588 412966 354640 412972
rect 368860 412978 368888 413034
rect 369308 413024 369360 413030
rect 368860 412972 369308 412978
rect 374368 413024 374420 413030
rect 368860 412966 369360 412972
rect 374366 412992 374368 413001
rect 374420 412992 374422 413001
rect 368860 412950 369348 412966
rect 374366 412927 374422 412936
rect 375484 412865 375512 413034
rect 383476 413024 383528 413030
rect 383580 413001 383608 413850
rect 383856 413817 383884 414054
rect 385040 414044 385092 414050
rect 385040 413986 385092 413992
rect 385052 413953 385080 413986
rect 412640 413976 412692 413982
rect 385038 413944 385094 413953
rect 412640 413918 412692 413924
rect 385038 413879 385094 413888
rect 393136 413908 393188 413914
rect 393136 413850 393188 413856
rect 387340 413840 387392 413846
rect 383842 413808 383898 413817
rect 387340 413782 387392 413788
rect 383842 413743 383898 413752
rect 386052 413704 386104 413710
rect 386052 413646 386104 413652
rect 384948 413500 385000 413506
rect 384948 413442 385000 413448
rect 384960 413030 384988 413442
rect 384948 413024 385000 413030
rect 383566 412992 383622 413001
rect 383528 412972 383566 412978
rect 383476 412966 383566 412972
rect 376576 412956 376628 412962
rect 383488 412950 383566 412966
rect 383566 412927 383622 412936
rect 384946 412992 384948 413001
rect 386064 413001 386092 413646
rect 386420 413296 386472 413302
rect 386418 413264 386420 413273
rect 386472 413264 386474 413273
rect 386418 413199 386474 413208
rect 387352 413137 387380 413782
rect 388352 413772 388404 413778
rect 388352 413714 388404 413720
rect 388364 413409 388392 413714
rect 389640 413636 389692 413642
rect 389640 413578 389692 413584
rect 388350 413400 388406 413409
rect 388350 413335 388406 413344
rect 387338 413128 387394 413137
rect 387338 413063 387394 413072
rect 385000 412992 385002 413001
rect 384946 412927 385002 412936
rect 386050 412992 386106 413001
rect 389652 412962 389680 413578
rect 393148 413370 393176 413850
rect 396080 413840 396132 413846
rect 412652 413817 412680 413918
rect 396080 413782 396132 413788
rect 412638 413808 412694 413817
rect 394700 413704 394752 413710
rect 396092 413681 396120 413782
rect 397460 413772 397512 413778
rect 412638 413743 412694 413752
rect 397460 413714 397512 413720
rect 397472 413681 397500 413714
rect 394700 413646 394752 413652
rect 396078 413672 396134 413681
rect 394712 413506 394740 413646
rect 396078 413607 396134 413616
rect 397458 413672 397514 413681
rect 397458 413607 397514 413616
rect 405740 413568 405792 413574
rect 405738 413536 405740 413545
rect 405792 413536 405794 413545
rect 393964 413500 394016 413506
rect 393964 413442 394016 413448
rect 394700 413500 394752 413506
rect 394700 413442 394752 413448
rect 395344 413500 395396 413506
rect 395344 413442 395396 413448
rect 404360 413500 404412 413506
rect 405738 413471 405794 413480
rect 404360 413442 404412 413448
rect 390928 413364 390980 413370
rect 390928 413306 390980 413312
rect 391848 413364 391900 413370
rect 391848 413306 391900 413312
rect 393136 413364 393188 413370
rect 393136 413306 393188 413312
rect 386050 412927 386052 412936
rect 376576 412898 376628 412904
rect 386104 412927 386106 412936
rect 389640 412956 389692 412962
rect 386052 412898 386104 412904
rect 389640 412898 389692 412904
rect 376588 412865 376616 412898
rect 386064 412867 386092 412898
rect 375470 412856 375526 412865
rect 375470 412791 375526 412800
rect 376574 412856 376630 412865
rect 376574 412791 376630 412800
rect 389652 412729 389680 412898
rect 390940 412729 390968 413306
rect 391860 413166 391888 413306
rect 391756 413160 391808 413166
rect 391756 413102 391808 413108
rect 391848 413160 391900 413166
rect 391848 413102 391900 413108
rect 391768 412729 391796 413102
rect 393148 412729 393176 413306
rect 393976 413302 394004 413442
rect 393964 413296 394016 413302
rect 393964 413238 394016 413244
rect 393320 412888 393372 412894
rect 393318 412856 393320 412865
rect 393372 412856 393374 412865
rect 393318 412791 393374 412800
rect 393976 412729 394004 413238
rect 394700 412820 394752 412826
rect 394700 412762 394752 412768
rect 394712 412729 394740 412762
rect 395356 412729 395384 413442
rect 404372 413409 404400 413442
rect 407120 413432 407172 413438
rect 404358 413400 404414 413409
rect 401600 413364 401652 413370
rect 407120 413374 407172 413380
rect 404358 413335 404414 413344
rect 401600 413306 401652 413312
rect 401612 413273 401640 413306
rect 403164 413296 403216 413302
rect 401598 413264 401654 413273
rect 401598 413199 401654 413208
rect 403162 413264 403164 413273
rect 407132 413273 407160 413374
rect 403216 413264 403218 413273
rect 403162 413199 403218 413208
rect 407118 413264 407174 413273
rect 407118 413199 407174 413208
rect 408500 413228 408552 413234
rect 408500 413170 408552 413176
rect 398840 413160 398892 413166
rect 398838 413128 398840 413137
rect 408512 413137 408540 413170
rect 398892 413128 398894 413137
rect 408498 413128 408554 413137
rect 398838 413063 398894 413072
rect 400220 413092 400272 413098
rect 408498 413063 408554 413072
rect 400220 413034 400272 413040
rect 400232 413001 400260 413034
rect 400218 412992 400274 413001
rect 397460 412956 397512 412962
rect 400218 412927 400274 412936
rect 397460 412898 397512 412904
rect 397472 412865 397500 412898
rect 397458 412856 397514 412865
rect 397458 412791 397514 412800
rect 396080 412752 396132 412758
rect 389638 412720 389694 412729
rect 389638 412655 389694 412664
rect 390926 412720 390982 412729
rect 390926 412655 390982 412664
rect 391754 412720 391810 412729
rect 391754 412655 391810 412664
rect 393134 412720 393190 412729
rect 393134 412655 393190 412664
rect 393962 412720 394018 412729
rect 393962 412655 394018 412664
rect 394698 412720 394754 412729
rect 394698 412655 394754 412664
rect 395342 412720 395398 412729
rect 395342 412655 395398 412664
rect 396078 412720 396080 412729
rect 396132 412720 396134 412729
rect 396078 412655 396134 412664
rect 405738 412720 405794 412729
rect 405738 412655 405740 412664
rect 405792 412655 405794 412664
rect 405740 412626 405792 412632
rect 350632 412004 350684 412010
rect 350632 411946 350684 411952
rect 419540 411936 419592 411942
rect 419540 411878 419592 411884
rect 397460 411868 397512 411874
rect 397460 411810 397512 411816
rect 388076 411800 388128 411806
rect 388074 411768 388076 411777
rect 388128 411768 388130 411777
rect 388074 411703 388130 411712
rect 391020 411732 391072 411738
rect 391020 411674 391072 411680
rect 391032 411641 391060 411674
rect 397472 411641 397500 411810
rect 399116 411664 399168 411670
rect 391018 411632 391074 411641
rect 391018 411567 391074 411576
rect 397458 411632 397514 411641
rect 399114 411632 399116 411641
rect 399168 411632 399170 411641
rect 397458 411567 397514 411576
rect 398012 411596 398064 411602
rect 399114 411567 399170 411576
rect 398012 411538 398064 411544
rect 398024 411505 398052 411538
rect 400956 411528 401008 411534
rect 389270 411496 389326 411505
rect 389270 411431 389326 411440
rect 398010 411496 398066 411505
rect 398010 411431 398066 411440
rect 400954 411496 400956 411505
rect 401008 411496 401010 411505
rect 403254 411496 403310 411505
rect 400954 411431 401010 411440
rect 401692 411460 401744 411466
rect 389284 411262 389312 411431
rect 403254 411431 403310 411440
rect 401692 411402 401744 411408
rect 401704 411369 401732 411402
rect 401690 411360 401746 411369
rect 403268 411330 403296 411431
rect 404360 411392 404412 411398
rect 404358 411360 404360 411369
rect 404412 411360 404414 411369
rect 401690 411295 401746 411304
rect 403256 411324 403308 411330
rect 404358 411295 404414 411304
rect 403256 411266 403308 411272
rect 389272 411256 389324 411262
rect 389272 411198 389324 411204
rect 389732 411188 389784 411194
rect 389732 411130 389784 411136
rect 389744 411097 389772 411130
rect 389730 411088 389786 411097
rect 389730 411023 389786 411032
rect 342260 410780 342312 410786
rect 342260 410722 342312 410728
rect 340880 410712 340932 410718
rect 340880 410654 340932 410660
rect 392308 410644 392360 410650
rect 392308 410586 392360 410592
rect 392320 410417 392348 410586
rect 409972 410576 410024 410582
rect 409972 410518 410024 410524
rect 409984 410417 410012 410518
rect 392306 410408 392362 410417
rect 392306 410343 392362 410352
rect 409970 410408 410026 410417
rect 409970 410343 410026 410352
rect 419552 393009 419580 411878
rect 419538 393000 419594 393009
rect 419538 392935 419594 392944
rect 419538 390688 419594 390697
rect 419538 390623 419594 390632
rect 339500 382220 339552 382226
rect 339500 382162 339552 382168
rect 338120 380860 338172 380866
rect 338120 380802 338172 380808
rect 416410 324048 416466 324057
rect 416410 323983 416466 323992
rect 337752 322244 337804 322250
rect 337752 322186 337804 322192
rect 337764 322017 337792 322186
rect 337750 322008 337806 322017
rect 337750 321943 337806 321952
rect 282828 321020 282880 321026
rect 282828 320962 282880 320968
rect 337384 321020 337436 321026
rect 337384 320962 337436 320968
rect 338028 321020 338080 321026
rect 338028 320962 338080 320968
rect 282840 320793 282868 320962
rect 282826 320784 282882 320793
rect 282826 320719 282882 320728
rect 282736 320340 282788 320346
rect 282736 320282 282788 320288
rect 282092 320272 282144 320278
rect 282092 320214 282144 320220
rect 60950 320062 61424 320090
rect 59912 319932 59964 319938
rect 59912 319874 59964 319880
rect 61396 317393 61424 320062
rect 62868 317898 62896 320076
rect 64800 318782 64828 320076
rect 66364 320062 66746 320090
rect 64788 318776 64840 318782
rect 64788 318718 64840 318724
rect 64788 318572 64840 318578
rect 64788 318514 64840 318520
rect 64800 317898 64828 318514
rect 62856 317892 62908 317898
rect 62856 317834 62908 317840
rect 64788 317892 64840 317898
rect 64788 317834 64840 317840
rect 64788 317756 64840 317762
rect 64788 317698 64840 317704
rect 62028 317688 62080 317694
rect 62028 317630 62080 317636
rect 61382 317384 61438 317393
rect 61382 317319 61438 317328
rect 59452 252544 59504 252550
rect 59452 252486 59504 252492
rect 59360 205624 59412 205630
rect 59360 205566 59412 205572
rect 59268 64864 59320 64870
rect 59268 64806 59320 64812
rect 57888 17944 57940 17950
rect 57888 17886 57940 17892
rect 60004 6452 60056 6458
rect 60004 6394 60056 6400
rect 52828 5296 52880 5302
rect 52828 5238 52880 5244
rect 51632 4276 51684 4282
rect 51632 4218 51684 4224
rect 50528 3188 50580 3194
rect 50528 3130 50580 3136
rect 50988 3188 51040 3194
rect 50988 3130 51040 3136
rect 50436 3120 50488 3126
rect 50436 3062 50488 3068
rect 49332 2984 49384 2990
rect 49332 2926 49384 2932
rect 48148 2094 48268 2122
rect 48148 480 48176 2094
rect 49344 480 49372 2926
rect 50540 480 50568 3130
rect 51644 480 51672 4218
rect 52840 480 52868 5238
rect 58808 4412 58860 4418
rect 58808 4354 58860 4360
rect 55220 4344 55272 4350
rect 55220 4286 55272 4292
rect 54024 3052 54076 3058
rect 54024 2994 54076 3000
rect 54036 480 54064 2994
rect 55232 480 55260 4286
rect 56416 3188 56468 3194
rect 56416 3130 56468 3136
rect 56428 480 56456 3130
rect 57612 3120 57664 3126
rect 57612 3062 57664 3068
rect 57624 480 57652 3062
rect 58820 480 58848 4354
rect 60016 480 60044 6394
rect 60740 5432 60792 5438
rect 60740 5374 60792 5380
rect 60752 5302 60780 5374
rect 60740 5296 60792 5302
rect 60740 5238 60792 5244
rect 61200 3392 61252 3398
rect 61014 3360 61070 3369
rect 61200 3334 61252 3340
rect 61014 3295 61016 3304
rect 61068 3295 61070 3304
rect 61016 3266 61068 3272
rect 61212 480 61240 3334
rect 61396 3262 61424 317319
rect 62040 3398 62068 317630
rect 62396 4480 62448 4486
rect 62396 4422 62448 4428
rect 62028 3392 62080 3398
rect 62120 3392 62172 3398
rect 62028 3334 62080 3340
rect 62118 3360 62120 3369
rect 62172 3360 62174 3369
rect 62118 3295 62174 3304
rect 61384 3256 61436 3262
rect 61384 3198 61436 3204
rect 62408 480 62436 4422
rect 63592 3256 63644 3262
rect 63592 3198 63644 3204
rect 63604 480 63632 3198
rect 64800 480 64828 317698
rect 66260 227996 66312 228002
rect 66260 227938 66312 227944
rect 66272 227905 66300 227938
rect 66258 227896 66314 227905
rect 66258 227831 66314 227840
rect 66260 170060 66312 170066
rect 66260 170002 66312 170008
rect 66272 169969 66300 170002
rect 66258 169960 66314 169969
rect 66258 169895 66314 169904
rect 65984 4548 66036 4554
rect 65984 4490 66036 4496
rect 65996 480 66024 4490
rect 66364 3398 66392 320062
rect 68664 317966 68692 320076
rect 70412 320062 70610 320090
rect 68652 317960 68704 317966
rect 68652 317902 68704 317908
rect 67548 317824 67600 317830
rect 67548 317766 67600 317772
rect 67560 4758 67588 317766
rect 69388 216980 69440 216986
rect 69388 216922 69440 216928
rect 69400 216889 69428 216922
rect 69386 216880 69442 216889
rect 69386 216815 69442 216824
rect 69388 181076 69440 181082
rect 69388 181018 69440 181024
rect 69400 180985 69428 181018
rect 69386 180976 69442 180985
rect 69386 180911 69442 180920
rect 67088 4752 67140 4758
rect 67088 4694 67140 4700
rect 67548 4752 67600 4758
rect 67548 4694 67600 4700
rect 66352 3392 66404 3398
rect 66352 3334 66404 3340
rect 67100 610 67128 4694
rect 69480 4616 69532 4622
rect 69480 4558 69532 4564
rect 68284 3392 68336 3398
rect 68284 3334 68336 3340
rect 67088 604 67140 610
rect 67088 546 67140 552
rect 67180 604 67232 610
rect 67180 546 67232 552
rect 67192 480 67220 546
rect 68296 480 68324 3334
rect 69492 480 69520 4558
rect 70412 3330 70440 320062
rect 72528 318646 72556 320076
rect 72516 318640 72568 318646
rect 72516 318582 72568 318588
rect 74448 317960 74500 317966
rect 74448 317902 74500 317908
rect 72976 317892 73028 317898
rect 72976 317834 73028 317840
rect 71778 4176 71834 4185
rect 72988 4146 73016 317834
rect 74460 299674 74488 317902
rect 74448 299668 74500 299674
rect 74448 299610 74500 299616
rect 74448 299532 74500 299538
rect 74448 299474 74500 299480
rect 74460 298110 74488 299474
rect 74264 298104 74316 298110
rect 74264 298046 74316 298052
rect 74448 298104 74500 298110
rect 74448 298046 74500 298052
rect 74276 288454 74304 298046
rect 74264 288448 74316 288454
rect 74264 288390 74316 288396
rect 74356 288448 74408 288454
rect 74356 288390 74408 288396
rect 74368 280242 74396 288390
rect 74368 280214 74488 280242
rect 74460 278769 74488 280214
rect 74262 278760 74318 278769
rect 74262 278695 74318 278704
rect 74446 278760 74502 278769
rect 74446 278695 74502 278704
rect 74276 269142 74304 278695
rect 74264 269136 74316 269142
rect 74264 269078 74316 269084
rect 74356 269136 74408 269142
rect 74356 269078 74408 269084
rect 74368 260930 74396 269078
rect 74368 260902 74488 260930
rect 74460 259457 74488 260902
rect 74262 259448 74318 259457
rect 74262 259383 74318 259392
rect 74446 259448 74502 259457
rect 74446 259383 74502 259392
rect 74276 249830 74304 259383
rect 74264 249824 74316 249830
rect 74264 249766 74316 249772
rect 74448 249824 74500 249830
rect 74448 249766 74500 249772
rect 74460 241754 74488 249766
rect 74368 241726 74488 241754
rect 74368 241534 74396 241726
rect 74356 241528 74408 241534
rect 74356 241470 74408 241476
rect 74448 241528 74500 241534
rect 74448 241470 74500 241476
rect 74460 240145 74488 241470
rect 74262 240136 74318 240145
rect 74262 240071 74318 240080
rect 74446 240136 74502 240145
rect 74446 240071 74502 240080
rect 74276 230518 74304 240071
rect 74264 230512 74316 230518
rect 74264 230454 74316 230460
rect 74448 230512 74500 230518
rect 74448 230454 74500 230460
rect 74460 220833 74488 230454
rect 74262 220824 74318 220833
rect 74262 220759 74318 220768
rect 74446 220824 74502 220833
rect 74446 220759 74502 220768
rect 74276 211177 74304 220759
rect 74262 211168 74318 211177
rect 74262 211103 74318 211112
rect 74446 211168 74502 211177
rect 74446 211103 74502 211112
rect 74460 201482 74488 211103
rect 74264 201476 74316 201482
rect 74264 201418 74316 201424
rect 74448 201476 74500 201482
rect 74448 201418 74500 201424
rect 74276 191894 74304 201418
rect 74264 191888 74316 191894
rect 74264 191830 74316 191836
rect 74356 191888 74408 191894
rect 74356 191830 74408 191836
rect 74368 183598 74396 191830
rect 74356 183592 74408 183598
rect 74356 183534 74408 183540
rect 74448 183592 74500 183598
rect 74448 183534 74500 183540
rect 74460 182170 74488 183534
rect 74264 182164 74316 182170
rect 74264 182106 74316 182112
rect 74448 182164 74500 182170
rect 74448 182106 74500 182112
rect 74276 172553 74304 182106
rect 74262 172544 74318 172553
rect 74262 172479 74318 172488
rect 74446 172544 74502 172553
rect 74446 172479 74502 172488
rect 74460 162858 74488 172479
rect 74264 162852 74316 162858
rect 74264 162794 74316 162800
rect 74448 162852 74500 162858
rect 74448 162794 74500 162800
rect 74276 153241 74304 162794
rect 74262 153232 74318 153241
rect 74262 153167 74318 153176
rect 74446 153232 74502 153241
rect 74446 153167 74502 153176
rect 74460 143546 74488 153167
rect 74448 143540 74500 143546
rect 74448 143482 74500 143488
rect 74446 125624 74502 125633
rect 74446 125559 74502 125568
rect 74460 124137 74488 125559
rect 74446 124128 74502 124137
rect 74446 124063 74502 124072
rect 74356 114572 74408 114578
rect 74356 114514 74408 114520
rect 74368 106418 74396 114514
rect 74356 106412 74408 106418
rect 74356 106354 74408 106360
rect 74448 106412 74500 106418
rect 74448 106354 74500 106360
rect 74460 104854 74488 106354
rect 74264 104848 74316 104854
rect 74264 104790 74316 104796
rect 74448 104848 74500 104854
rect 74448 104790 74500 104796
rect 74276 95266 74304 104790
rect 74264 95260 74316 95266
rect 74264 95202 74316 95208
rect 74356 95260 74408 95266
rect 74356 95202 74408 95208
rect 74368 87106 74396 95202
rect 74356 87100 74408 87106
rect 74356 87042 74408 87048
rect 74448 87100 74500 87106
rect 74448 87042 74500 87048
rect 74460 85542 74488 87042
rect 74264 85536 74316 85542
rect 74264 85478 74316 85484
rect 74448 85536 74500 85542
rect 74448 85478 74500 85484
rect 74276 75954 74304 85478
rect 74264 75948 74316 75954
rect 74264 75890 74316 75896
rect 74356 75948 74408 75954
rect 74356 75890 74408 75896
rect 74368 67726 74396 75890
rect 74356 67720 74408 67726
rect 74356 67662 74408 67668
rect 74448 67720 74500 67726
rect 74448 67662 74500 67668
rect 74460 66230 74488 67662
rect 74264 66224 74316 66230
rect 74264 66166 74316 66172
rect 74448 66224 74500 66230
rect 74448 66166 74500 66172
rect 74276 56642 74304 66166
rect 74264 56636 74316 56642
rect 74264 56578 74316 56584
rect 74448 56636 74500 56642
rect 74448 56578 74500 56584
rect 74460 48498 74488 56578
rect 74368 48470 74488 48498
rect 74368 48362 74396 48470
rect 74368 48334 74488 48362
rect 74460 46918 74488 48334
rect 74264 46912 74316 46918
rect 74264 46854 74316 46860
rect 74448 46912 74500 46918
rect 74448 46854 74500 46860
rect 74276 37330 74304 46854
rect 74264 37324 74316 37330
rect 74264 37266 74316 37272
rect 74356 37324 74408 37330
rect 74356 37266 74408 37272
rect 74368 29050 74396 37266
rect 74368 29022 74488 29050
rect 74460 27606 74488 29022
rect 74264 27600 74316 27606
rect 74264 27542 74316 27548
rect 74448 27600 74500 27606
rect 74448 27542 74500 27548
rect 74276 18018 74304 27542
rect 74080 18012 74132 18018
rect 74080 17954 74132 17960
rect 74264 18012 74316 18018
rect 74264 17954 74316 17960
rect 74092 9722 74120 17954
rect 74080 9716 74132 9722
rect 74080 9658 74132 9664
rect 74264 9716 74316 9722
rect 74264 9658 74316 9664
rect 73068 4684 73120 4690
rect 73068 4626 73120 4632
rect 73080 4298 73108 4626
rect 73080 4270 73200 4298
rect 73066 4176 73122 4185
rect 71778 4111 71780 4120
rect 71832 4111 71834 4120
rect 71872 4140 71924 4146
rect 71780 4082 71832 4088
rect 71872 4082 71924 4088
rect 72976 4140 73028 4146
rect 73066 4111 73068 4120
rect 72976 4082 73028 4088
rect 73120 4111 73122 4120
rect 73068 4082 73120 4088
rect 70400 3324 70452 3330
rect 70400 3266 70452 3272
rect 70676 3324 70728 3330
rect 70676 3266 70728 3272
rect 70688 480 70716 3266
rect 71884 480 71912 4082
rect 73172 4026 73200 4270
rect 73080 3998 73200 4026
rect 73080 480 73108 3998
rect 74276 480 74304 9658
rect 74552 4146 74580 320076
rect 76484 318510 76512 320076
rect 76472 318504 76524 318510
rect 76472 318446 76524 318452
rect 78416 318034 78444 320076
rect 80072 320062 80362 320090
rect 81452 320062 82294 320090
rect 78404 318028 78456 318034
rect 78404 317970 78456 317976
rect 79968 318028 80020 318034
rect 79968 317970 80020 317976
rect 75826 228032 75882 228041
rect 75826 227967 75828 227976
rect 75880 227967 75882 227976
rect 75828 227938 75880 227944
rect 77206 217016 77262 217025
rect 77206 216951 77208 216960
rect 77260 216951 77262 216960
rect 77208 216922 77260 216928
rect 77206 181112 77262 181121
rect 77206 181047 77208 181056
rect 77260 181047 77262 181056
rect 77208 181018 77260 181024
rect 75826 170096 75882 170105
rect 75826 170031 75828 170040
rect 75880 170031 75882 170040
rect 75828 170002 75880 170008
rect 74632 143540 74684 143546
rect 74632 143482 74684 143488
rect 74644 125633 74672 143482
rect 74630 125624 74686 125633
rect 74630 125559 74686 125568
rect 74722 124128 74778 124137
rect 74722 124063 74778 124072
rect 74736 114578 74764 124063
rect 74724 114572 74776 114578
rect 74724 114514 74776 114520
rect 77206 76256 77262 76265
rect 77206 76191 77262 76200
rect 77220 76129 77248 76191
rect 77206 76120 77262 76129
rect 77206 76055 77262 76064
rect 78588 5432 78640 5438
rect 78588 5374 78640 5380
rect 78600 5302 78628 5374
rect 78588 5296 78640 5302
rect 78588 5238 78640 5244
rect 78864 4888 78916 4894
rect 78862 4856 78864 4865
rect 78916 4856 78918 4865
rect 78862 4791 78918 4800
rect 76656 4752 76708 4758
rect 76656 4694 76708 4700
rect 74540 4140 74592 4146
rect 74540 4082 74592 4088
rect 75458 3768 75514 3777
rect 75458 3703 75514 3712
rect 75276 3392 75328 3398
rect 75104 3340 75276 3346
rect 75104 3334 75328 3340
rect 75104 3330 75316 3334
rect 75092 3324 75316 3330
rect 75144 3318 75316 3324
rect 75092 3266 75144 3272
rect 75472 480 75500 3703
rect 76668 480 76696 4694
rect 79980 4078 80008 317970
rect 80072 5506 80100 320062
rect 80060 5500 80112 5506
rect 80060 5442 80112 5448
rect 80244 5500 80296 5506
rect 80244 5442 80296 5448
rect 79048 4072 79100 4078
rect 77850 4040 77906 4049
rect 79048 4014 79100 4020
rect 79968 4072 80020 4078
rect 80060 4072 80112 4078
rect 79968 4014 80020 4020
rect 80058 4040 80060 4049
rect 80112 4040 80114 4049
rect 77850 3975 77906 3984
rect 77864 480 77892 3975
rect 79060 480 79088 4014
rect 80058 3975 80114 3984
rect 80256 480 80284 5442
rect 81452 4298 81480 320062
rect 82728 318776 82780 318782
rect 82728 318718 82780 318724
rect 81912 5222 82124 5250
rect 81912 5166 81940 5222
rect 82096 5166 82124 5222
rect 81900 5160 81952 5166
rect 82084 5160 82136 5166
rect 81900 5102 81952 5108
rect 81990 5128 82046 5137
rect 82084 5102 82136 5108
rect 81990 5063 81992 5072
rect 82044 5063 82046 5072
rect 81992 5034 82044 5040
rect 81990 4992 82046 5001
rect 81990 4927 81992 4936
rect 82044 4927 82046 4936
rect 81992 4898 82044 4904
rect 81360 4270 81480 4298
rect 81360 4146 81388 4270
rect 82740 4146 82768 318718
rect 83832 5432 83884 5438
rect 83832 5374 83884 5380
rect 81348 4140 81400 4146
rect 81348 4082 81400 4088
rect 81440 4140 81492 4146
rect 81440 4082 81492 4088
rect 82728 4140 82780 4146
rect 82728 4082 82780 4088
rect 82820 4140 82872 4146
rect 82820 4082 82872 4088
rect 81452 480 81480 4082
rect 82832 4026 82860 4082
rect 82648 3998 82860 4026
rect 82648 480 82676 3998
rect 83844 480 83872 5374
rect 84212 4010 84240 320076
rect 86236 318374 86264 320076
rect 88168 318714 88196 320076
rect 89732 320062 90114 320090
rect 88156 318708 88208 318714
rect 88156 318650 88208 318656
rect 88248 318708 88300 318714
rect 88248 318650 88300 318656
rect 88260 318510 88288 318650
rect 86868 318504 86920 318510
rect 86868 318446 86920 318452
rect 88248 318504 88300 318510
rect 88248 318446 88300 318452
rect 89536 318504 89588 318510
rect 89536 318446 89588 318452
rect 86224 318368 86276 318374
rect 86224 318310 86276 318316
rect 86880 263770 86908 318446
rect 89548 302274 89576 318446
rect 89456 302246 89576 302274
rect 89456 302138 89484 302246
rect 89456 302110 89576 302138
rect 89548 292618 89576 302110
rect 89548 292590 89668 292618
rect 89640 292482 89668 292590
rect 89548 292454 89668 292482
rect 89548 282962 89576 292454
rect 89456 282934 89576 282962
rect 89456 282826 89484 282934
rect 89456 282798 89576 282826
rect 89548 273306 89576 282798
rect 89548 273278 89668 273306
rect 86868 263764 86920 263770
rect 86868 263706 86920 263712
rect 86868 263628 86920 263634
rect 86868 263570 86920 263576
rect 86880 227866 86908 263570
rect 89640 253858 89668 273278
rect 89548 253830 89668 253858
rect 89548 244338 89576 253830
rect 89456 244310 89576 244338
rect 89456 244202 89484 244310
rect 89456 244174 89576 244202
rect 89548 234682 89576 244174
rect 89548 234654 89668 234682
rect 86868 227860 86920 227866
rect 86868 227802 86920 227808
rect 86868 227724 86920 227730
rect 86868 227666 86920 227672
rect 86880 180946 86908 227666
rect 89536 216912 89588 216918
rect 89534 216880 89536 216889
rect 89588 216880 89590 216889
rect 89534 216815 89590 216824
rect 89640 215234 89668 234654
rect 89548 215206 89668 215234
rect 89548 202910 89576 215206
rect 89352 202904 89404 202910
rect 89352 202846 89404 202852
rect 89536 202904 89588 202910
rect 89536 202846 89588 202852
rect 89364 196042 89392 202846
rect 89352 196036 89404 196042
rect 89352 195978 89404 195984
rect 89444 195900 89496 195906
rect 89444 195842 89496 195848
rect 86868 180940 86920 180946
rect 86868 180882 86920 180888
rect 86868 180804 86920 180810
rect 86868 180746 86920 180752
rect 86880 169930 86908 180746
rect 89456 173942 89484 195842
rect 89444 173936 89496 173942
rect 89444 173878 89496 173884
rect 89628 173936 89680 173942
rect 89628 173878 89680 173884
rect 89534 170096 89590 170105
rect 89534 170031 89590 170040
rect 86868 169924 86920 169930
rect 86868 169866 86920 169872
rect 89548 169833 89576 170031
rect 89534 169824 89590 169833
rect 86868 169788 86920 169794
rect 89534 169759 89590 169768
rect 86868 169730 86920 169736
rect 86880 5642 86908 169730
rect 89640 167090 89668 173878
rect 89548 167062 89668 167090
rect 89548 166954 89576 167062
rect 89456 166926 89576 166954
rect 89456 157486 89484 166926
rect 89444 157480 89496 157486
rect 89444 157422 89496 157428
rect 89444 157344 89496 157350
rect 89444 157286 89496 157292
rect 89456 157162 89484 157286
rect 89456 157134 89576 157162
rect 89548 154562 89576 157134
rect 89260 154556 89312 154562
rect 89260 154498 89312 154504
rect 89536 154556 89588 154562
rect 89536 154498 89588 154504
rect 89272 144945 89300 154498
rect 89258 144936 89314 144945
rect 89258 144871 89314 144880
rect 89442 144936 89498 144945
rect 89442 144871 89498 144880
rect 89456 138038 89484 144871
rect 89444 138032 89496 138038
rect 89444 137974 89496 137980
rect 89536 137896 89588 137902
rect 89536 137838 89588 137844
rect 89548 128450 89576 137838
rect 89536 128444 89588 128450
rect 89536 128386 89588 128392
rect 89444 128308 89496 128314
rect 89444 128250 89496 128256
rect 89456 124098 89484 128250
rect 89444 124092 89496 124098
rect 89444 124034 89496 124040
rect 89628 124092 89680 124098
rect 89628 124034 89680 124040
rect 89640 118726 89668 124034
rect 89628 118720 89680 118726
rect 89628 118662 89680 118668
rect 89536 118584 89588 118590
rect 89536 118526 89588 118532
rect 89548 109138 89576 118526
rect 89536 109132 89588 109138
rect 89536 109074 89588 109080
rect 89444 108996 89496 109002
rect 89444 108938 89496 108944
rect 89456 104854 89484 108938
rect 89260 104848 89312 104854
rect 89260 104790 89312 104796
rect 89444 104848 89496 104854
rect 89444 104790 89496 104796
rect 89272 95266 89300 104790
rect 89260 95260 89312 95266
rect 89260 95202 89312 95208
rect 89352 95260 89404 95266
rect 89352 95202 89404 95208
rect 89364 89434 89392 95202
rect 89364 89406 89576 89434
rect 89548 80170 89576 89406
rect 89536 80164 89588 80170
rect 89536 80106 89588 80112
rect 89536 80028 89588 80034
rect 89536 79970 89588 79976
rect 89548 70394 89576 79970
rect 89628 76152 89680 76158
rect 89626 76120 89628 76129
rect 89680 76120 89682 76129
rect 89626 76055 89682 76064
rect 89456 70366 89576 70394
rect 89456 70258 89484 70366
rect 89456 70230 89576 70258
rect 89548 51082 89576 70230
rect 89456 51066 89576 51082
rect 89444 51060 89576 51066
rect 89496 51054 89576 51060
rect 89628 51060 89680 51066
rect 89444 51002 89496 51008
rect 89628 51002 89680 51008
rect 89456 50971 89484 51002
rect 89640 48278 89668 51002
rect 89352 48272 89404 48278
rect 89352 48214 89404 48220
rect 89628 48272 89680 48278
rect 89628 48214 89680 48220
rect 89364 38690 89392 48214
rect 89352 38684 89404 38690
rect 89352 38626 89404 38632
rect 89536 38684 89588 38690
rect 89536 38626 89588 38632
rect 89548 31793 89576 38626
rect 89534 31784 89590 31793
rect 89534 31719 89590 31728
rect 89258 26344 89314 26353
rect 89258 26279 89314 26288
rect 89272 26246 89300 26279
rect 89168 26240 89220 26246
rect 89168 26182 89220 26188
rect 89260 26240 89312 26246
rect 89260 26182 89312 26188
rect 89180 21418 89208 26182
rect 89168 21412 89220 21418
rect 89168 21354 89220 21360
rect 89444 21412 89496 21418
rect 89444 21354 89496 21360
rect 89456 8362 89484 21354
rect 89352 8356 89404 8362
rect 89352 8298 89404 8304
rect 89444 8356 89496 8362
rect 89444 8298 89496 8304
rect 86132 5636 86184 5642
rect 86132 5578 86184 5584
rect 86868 5636 86920 5642
rect 86868 5578 86920 5584
rect 86038 4176 86094 4185
rect 86038 4111 86040 4120
rect 86092 4111 86094 4120
rect 86040 4082 86092 4088
rect 84200 4004 84252 4010
rect 84200 3946 84252 3952
rect 84936 4004 84988 4010
rect 84936 3946 84988 3952
rect 84948 480 84976 3946
rect 86144 480 86172 5578
rect 87328 5364 87380 5370
rect 87328 5306 87380 5312
rect 86866 5128 86922 5137
rect 86866 5063 86868 5072
rect 86920 5063 86922 5072
rect 86868 5034 86920 5040
rect 86774 4992 86830 5001
rect 86774 4927 86776 4936
rect 86828 4927 86830 4936
rect 86776 4898 86828 4904
rect 86868 4888 86920 4894
rect 86866 4856 86868 4865
rect 86920 4856 86922 4865
rect 86866 4791 86922 4800
rect 87340 480 87368 5306
rect 89364 1154 89392 8298
rect 89534 4176 89590 4185
rect 89732 4162 89760 320062
rect 92032 318306 92060 320076
rect 92020 318300 92072 318306
rect 92020 318242 92072 318248
rect 93768 318300 93820 318306
rect 93768 318242 93820 318248
rect 91744 216912 91796 216918
rect 91742 216880 91744 216889
rect 91796 216880 91798 216889
rect 91742 216815 91798 216824
rect 91744 76152 91796 76158
rect 91742 76120 91744 76129
rect 91796 76120 91798 76129
rect 91742 76055 91798 76064
rect 90914 5264 90970 5273
rect 90914 5199 90970 5208
rect 89534 4111 89590 4120
rect 89640 4134 89760 4162
rect 89548 4078 89576 4111
rect 89536 4072 89588 4078
rect 89536 4014 89588 4020
rect 89444 4004 89496 4010
rect 89444 3946 89496 3952
rect 89456 3913 89484 3946
rect 89640 3942 89668 4134
rect 89720 4004 89772 4010
rect 89720 3946 89772 3952
rect 89628 3936 89680 3942
rect 89442 3904 89498 3913
rect 89628 3878 89680 3884
rect 89442 3839 89498 3848
rect 88524 1148 88576 1154
rect 88524 1090 88576 1096
rect 89352 1148 89404 1154
rect 89352 1090 89404 1096
rect 88536 480 88564 1090
rect 89732 480 89760 3946
rect 89904 3936 89956 3942
rect 89902 3904 89904 3913
rect 89956 3904 89958 3913
rect 89902 3839 89958 3848
rect 90928 480 90956 5199
rect 93216 4004 93268 4010
rect 93216 3946 93268 3952
rect 93228 3913 93256 3946
rect 93214 3904 93270 3913
rect 93214 3839 93270 3848
rect 92110 3632 92166 3641
rect 92110 3567 92166 3576
rect 92124 480 92152 3567
rect 93780 626 93808 318242
rect 93964 318238 93992 320076
rect 95252 320062 95910 320090
rect 96632 320062 97934 320090
rect 94412 318572 94464 318578
rect 94412 318514 94464 318520
rect 94596 318572 94648 318578
rect 94596 318514 94648 318520
rect 94424 318374 94452 318514
rect 94412 318368 94464 318374
rect 94412 318310 94464 318316
rect 94608 318306 94636 318514
rect 94596 318300 94648 318306
rect 94596 318242 94648 318248
rect 93952 318232 94004 318238
rect 93952 318174 94004 318180
rect 93860 5568 93912 5574
rect 93860 5510 93912 5516
rect 93872 5302 93900 5510
rect 93860 5296 93912 5302
rect 93860 5238 93912 5244
rect 95252 5234 95280 320062
rect 96528 318504 96580 318510
rect 96528 318446 96580 318452
rect 95240 5228 95292 5234
rect 95240 5170 95292 5176
rect 94502 5128 94558 5137
rect 94502 5063 94558 5072
rect 93860 3936 93912 3942
rect 93858 3904 93860 3913
rect 93912 3904 93914 3913
rect 93858 3839 93914 3848
rect 93320 598 93808 626
rect 93320 480 93348 598
rect 94516 480 94544 5063
rect 95514 3904 95570 3913
rect 95514 3839 95516 3848
rect 95568 3839 95570 3848
rect 95516 3810 95568 3816
rect 96540 3806 96568 318446
rect 96632 3913 96660 320062
rect 99852 318170 99880 320076
rect 99840 318164 99892 318170
rect 99840 318106 99892 318112
rect 100668 318164 100720 318170
rect 100668 318106 100720 318112
rect 98092 5228 98144 5234
rect 98092 5170 98144 5176
rect 96618 3904 96674 3913
rect 96618 3839 96674 3848
rect 96896 3868 96948 3874
rect 96896 3810 96948 3816
rect 95700 3800 95752 3806
rect 95700 3742 95752 3748
rect 96528 3800 96580 3806
rect 96528 3742 96580 3748
rect 95712 480 95740 3742
rect 96908 480 96936 3810
rect 98104 480 98132 5170
rect 99286 3496 99342 3505
rect 99286 3431 99342 3440
rect 99300 480 99328 3431
rect 100680 626 100708 318106
rect 101784 318102 101812 320076
rect 103532 320062 103730 320090
rect 104912 320062 105662 320090
rect 103428 318300 103480 318306
rect 103428 318242 103480 318248
rect 101772 318096 101824 318102
rect 101772 318038 101824 318044
rect 101586 4992 101642 5001
rect 101586 4927 101642 4936
rect 100496 598 100708 626
rect 100496 480 100524 598
rect 101600 480 101628 4927
rect 102598 3904 102654 3913
rect 103440 3874 103468 318242
rect 103532 5166 103560 320062
rect 103612 5568 103664 5574
rect 103612 5510 103664 5516
rect 103624 5166 103652 5510
rect 103520 5160 103572 5166
rect 103520 5102 103572 5108
rect 103612 5160 103664 5166
rect 103612 5102 103664 5108
rect 103518 3904 103574 3913
rect 102598 3839 102654 3848
rect 102784 3868 102836 3874
rect 102612 3806 102640 3839
rect 102784 3810 102836 3816
rect 103428 3868 103480 3874
rect 104912 3874 104940 320062
rect 107580 318374 107608 320076
rect 109052 320062 109526 320090
rect 110432 320062 111550 320090
rect 113192 320062 113482 320090
rect 114572 320062 115414 320090
rect 107568 318368 107620 318374
rect 107568 318310 107620 318316
rect 107660 318368 107712 318374
rect 107660 318310 107712 318316
rect 107568 318232 107620 318238
rect 107568 318174 107620 318180
rect 107476 318164 107528 318170
rect 107476 318106 107528 318112
rect 105084 5568 105136 5574
rect 105084 5510 105136 5516
rect 105096 5234 105124 5510
rect 105084 5228 105136 5234
rect 105084 5170 105136 5176
rect 105176 5228 105228 5234
rect 105176 5170 105228 5176
rect 103518 3839 103520 3848
rect 103428 3810 103480 3816
rect 103572 3839 103574 3848
rect 104900 3868 104952 3874
rect 103520 3810 103572 3816
rect 104900 3810 104952 3816
rect 102600 3800 102652 3806
rect 102600 3742 102652 3748
rect 102796 480 102824 3810
rect 103978 3360 104034 3369
rect 103978 3295 104034 3304
rect 103992 480 104020 3295
rect 105188 480 105216 5170
rect 106004 3800 106056 3806
rect 106188 3800 106240 3806
rect 106056 3760 106188 3788
rect 106004 3742 106056 3748
rect 106188 3742 106240 3748
rect 106280 3732 106332 3738
rect 106280 3674 106332 3680
rect 106292 3602 106320 3674
rect 106280 3596 106332 3602
rect 106280 3538 106332 3544
rect 106372 3596 106424 3602
rect 106372 3538 106424 3544
rect 106384 480 106412 3538
rect 107488 3482 107516 318106
rect 107580 3602 107608 318174
rect 107672 318102 107700 318310
rect 107660 318096 107712 318102
rect 107660 318038 107712 318044
rect 108764 6384 108816 6390
rect 108764 6326 108816 6332
rect 108212 3868 108264 3874
rect 108212 3810 108264 3816
rect 108224 3754 108252 3810
rect 108224 3738 108528 3754
rect 108224 3732 108540 3738
rect 108224 3726 108488 3732
rect 108488 3674 108540 3680
rect 107568 3596 107620 3602
rect 107568 3538 107620 3544
rect 107488 3454 107608 3482
rect 107580 480 107608 3454
rect 108776 480 108804 6326
rect 109052 5658 109080 320062
rect 109052 5630 109172 5658
rect 109040 5568 109092 5574
rect 109040 5510 109092 5516
rect 109052 5302 109080 5510
rect 109040 5296 109092 5302
rect 109040 5238 109092 5244
rect 109144 5098 109172 5630
rect 109132 5092 109184 5098
rect 109132 5034 109184 5040
rect 110432 3738 110460 320062
rect 111062 264344 111118 264353
rect 111062 264279 111118 264288
rect 111076 263673 111104 264279
rect 111062 263664 111118 263673
rect 111062 263599 111118 263608
rect 111062 228440 111118 228449
rect 111062 228375 111118 228384
rect 111076 227769 111104 228375
rect 111062 227760 111118 227769
rect 111062 227695 111118 227704
rect 111062 181520 111118 181529
rect 111062 181455 111118 181464
rect 111076 180849 111104 181455
rect 111062 180840 111118 180849
rect 111062 180775 111118 180784
rect 111062 170504 111118 170513
rect 111062 170439 111118 170448
rect 111076 169833 111104 170439
rect 111062 169824 111118 169833
rect 111062 169759 111118 169768
rect 112352 6316 112404 6322
rect 112352 6258 112404 6264
rect 110420 3732 110472 3738
rect 110420 3674 110472 3680
rect 111156 3732 111208 3738
rect 111156 3674 111208 3680
rect 109960 3596 110012 3602
rect 109960 3538 110012 3544
rect 109972 480 110000 3538
rect 111168 480 111196 3674
rect 112364 480 112392 6258
rect 113192 3806 113220 320062
rect 114468 318096 114520 318102
rect 114468 318038 114520 318044
rect 114480 3806 114508 318038
rect 114572 5030 114600 320062
rect 115846 318336 115902 318345
rect 115846 318271 115902 318280
rect 114560 5024 114612 5030
rect 114560 4966 114612 4972
rect 115860 3806 115888 318271
rect 115940 263696 115992 263702
rect 115938 263664 115940 263673
rect 115992 263664 115994 263673
rect 115938 263599 115994 263608
rect 115940 227792 115992 227798
rect 115938 227760 115940 227769
rect 115992 227760 115994 227769
rect 115938 227695 115994 227704
rect 115940 216776 115992 216782
rect 115938 216744 115940 216753
rect 115992 216744 115994 216753
rect 115938 216679 115994 216688
rect 115940 169856 115992 169862
rect 115938 169824 115940 169833
rect 115992 169824 115994 169833
rect 115938 169759 115994 169768
rect 115940 76016 115992 76022
rect 115938 75984 115940 75993
rect 115992 75984 115994 75993
rect 115938 75919 115994 75928
rect 115940 6248 115992 6254
rect 115940 6190 115992 6196
rect 113180 3800 113232 3806
rect 113180 3742 113232 3748
rect 113548 3800 113600 3806
rect 114468 3800 114520 3806
rect 113548 3742 113600 3748
rect 113560 480 113588 3742
rect 113744 3726 114140 3754
rect 114468 3742 114520 3748
rect 114744 3800 114796 3806
rect 114744 3742 114796 3748
rect 115848 3800 115900 3806
rect 115848 3742 115900 3748
rect 113744 3602 113772 3726
rect 114008 3664 114060 3670
rect 113836 3612 114008 3618
rect 113836 3606 114060 3612
rect 113732 3596 113784 3602
rect 113732 3538 113784 3544
rect 113836 3590 114048 3606
rect 114112 3602 114140 3726
rect 114100 3596 114152 3602
rect 113640 3528 113692 3534
rect 113836 3482 113864 3590
rect 114100 3538 114152 3544
rect 113692 3476 113864 3482
rect 113640 3470 113864 3476
rect 113652 3454 113864 3470
rect 114756 480 114784 3742
rect 115952 480 115980 6190
rect 116032 3800 116084 3806
rect 116032 3742 116084 3748
rect 116044 3602 116072 3742
rect 117136 3664 117188 3670
rect 117136 3606 117188 3612
rect 116032 3596 116084 3602
rect 116032 3538 116084 3544
rect 117148 480 117176 3606
rect 117332 3602 117360 320076
rect 118712 320062 119278 320090
rect 120092 320062 121210 320090
rect 122944 320062 123234 320090
rect 124784 320062 125166 320090
rect 126992 320062 127098 320090
rect 117320 3596 117372 3602
rect 117320 3538 117372 3544
rect 118240 3596 118292 3602
rect 118240 3538 118292 3544
rect 118252 480 118280 3538
rect 118712 3534 118740 320062
rect 118790 263936 118846 263945
rect 118790 263871 118846 263880
rect 118804 263702 118832 263871
rect 118792 263696 118844 263702
rect 118792 263638 118844 263644
rect 118790 228032 118846 228041
rect 118790 227967 118846 227976
rect 118804 227798 118832 227967
rect 118792 227792 118844 227798
rect 118792 227734 118844 227740
rect 118790 217016 118846 217025
rect 118790 216951 118846 216960
rect 118804 216782 118832 216951
rect 118792 216776 118844 216782
rect 118792 216718 118844 216724
rect 118790 170096 118846 170105
rect 118790 170031 118846 170040
rect 118804 169862 118832 170031
rect 118792 169856 118844 169862
rect 118792 169798 118844 169804
rect 118790 76256 118846 76265
rect 118790 76191 118846 76200
rect 118804 76022 118832 76191
rect 118792 76016 118844 76022
rect 118792 75958 118844 75964
rect 119436 5024 119488 5030
rect 119436 4966 119488 4972
rect 118700 3528 118752 3534
rect 118700 3470 118752 3476
rect 119448 480 119476 4966
rect 120092 4962 120120 320062
rect 121366 318200 121422 318209
rect 121366 318135 121422 318144
rect 120080 4956 120132 4962
rect 120080 4898 120132 4904
rect 121380 3670 121408 318135
rect 122746 318064 122802 318073
rect 122746 317999 122802 318008
rect 122760 3670 122788 317999
rect 120632 3664 120684 3670
rect 120632 3606 120684 3612
rect 121368 3664 121420 3670
rect 121368 3606 121420 3612
rect 121828 3664 121880 3670
rect 121828 3606 121880 3612
rect 122748 3664 122800 3670
rect 122748 3606 122800 3612
rect 122840 3664 122892 3670
rect 122840 3606 122892 3612
rect 120644 480 120672 3606
rect 121840 480 121868 3606
rect 122656 3528 122708 3534
rect 122852 3482 122880 3606
rect 122708 3476 122880 3482
rect 122656 3470 122880 3476
rect 122668 3454 122880 3470
rect 122944 3466 122972 320062
rect 124784 317490 124812 320062
rect 124772 317484 124824 317490
rect 124772 317426 124824 317432
rect 124864 317484 124916 317490
rect 124864 317426 124916 317432
rect 123024 6180 123076 6186
rect 123024 6122 123076 6128
rect 122932 3460 122984 3466
rect 122932 3402 122984 3408
rect 123036 480 123064 6122
rect 124876 5098 124904 317426
rect 124864 5092 124916 5098
rect 124864 5034 124916 5040
rect 126992 4894 127020 320062
rect 129016 318442 129044 320076
rect 129844 320062 130962 320090
rect 132512 320062 132894 320090
rect 133984 320062 134918 320090
rect 129004 318436 129056 318442
rect 129004 318378 129056 318384
rect 128266 180976 128322 180985
rect 128450 180976 128506 180985
rect 128322 180934 128450 180962
rect 128266 180911 128322 180920
rect 128450 180911 128506 180920
rect 127808 5160 127860 5166
rect 127808 5102 127860 5108
rect 126980 4888 127032 4894
rect 126980 4830 127032 4836
rect 127072 4888 127124 4894
rect 127072 4830 127124 4836
rect 127084 4706 127112 4830
rect 126624 4678 127112 4706
rect 124220 3528 124272 3534
rect 124220 3470 124272 3476
rect 124232 480 124260 3470
rect 125416 3460 125468 3466
rect 125416 3402 125468 3408
rect 125428 480 125456 3402
rect 126624 480 126652 4678
rect 127820 480 127848 5102
rect 129004 4956 129056 4962
rect 129004 4898 129056 4904
rect 129016 480 129044 4898
rect 129844 2854 129872 320062
rect 130200 5092 130252 5098
rect 130200 5034 130252 5040
rect 129832 2848 129884 2854
rect 129832 2790 129884 2796
rect 130212 480 130240 5034
rect 131394 4856 131450 4865
rect 132512 4826 132540 320062
rect 131394 4791 131450 4800
rect 132500 4820 132552 4826
rect 131408 480 131436 4791
rect 132500 4762 132552 4768
rect 132592 4820 132644 4826
rect 132592 4762 132644 4768
rect 132604 480 132632 4762
rect 133984 2922 134012 320062
rect 134524 318436 134576 318442
rect 134524 318378 134576 318384
rect 134536 5030 134564 318378
rect 136836 317558 136864 320076
rect 138032 320062 138782 320090
rect 139412 320062 140714 320090
rect 136824 317552 136876 317558
rect 136824 317494 136876 317500
rect 135166 264208 135222 264217
rect 135166 264143 135222 264152
rect 135180 263809 135208 264143
rect 135166 263800 135222 263809
rect 135166 263735 135222 263744
rect 135166 228304 135222 228313
rect 135166 228239 135222 228248
rect 135180 227905 135208 228239
rect 135166 227896 135222 227905
rect 135166 227831 135222 227840
rect 135166 217288 135222 217297
rect 135166 217223 135222 217232
rect 135180 216889 135208 217223
rect 135166 216880 135222 216889
rect 135166 216815 135222 216824
rect 135166 170368 135222 170377
rect 135166 170303 135222 170312
rect 135180 169969 135208 170303
rect 135166 169960 135222 169969
rect 135166 169895 135222 169904
rect 135166 76528 135222 76537
rect 135166 76463 135222 76472
rect 135180 76129 135208 76463
rect 135166 76120 135222 76129
rect 135166 76055 135222 76064
rect 137468 5160 137520 5166
rect 137468 5102 137520 5108
rect 134524 5024 134576 5030
rect 134524 4966 134576 4972
rect 134616 5024 134668 5030
rect 134616 4966 134668 4972
rect 137192 5024 137244 5030
rect 137192 4966 137244 4972
rect 134628 4826 134656 4966
rect 134616 4820 134668 4826
rect 134616 4762 134668 4768
rect 134892 4820 134944 4826
rect 134892 4762 134944 4768
rect 133972 2916 134024 2922
rect 133972 2858 134024 2864
rect 134904 480 134932 4762
rect 137204 4706 137232 4966
rect 137480 4894 137508 5102
rect 137468 4888 137520 4894
rect 137468 4830 137520 4836
rect 137560 4888 137612 4894
rect 137560 4830 137612 4836
rect 137572 4706 137600 4830
rect 137204 4678 137600 4706
rect 138032 4214 138060 320062
rect 138020 4208 138072 4214
rect 138020 4150 138072 4156
rect 139412 2990 139440 320062
rect 142632 317626 142660 320076
rect 143552 320062 144578 320090
rect 142620 317620 142672 317626
rect 142620 317562 142672 317568
rect 140042 264072 140098 264081
rect 140042 264007 140098 264016
rect 140056 263673 140084 264007
rect 140042 263664 140098 263673
rect 140042 263599 140098 263608
rect 140042 228168 140098 228177
rect 140042 228103 140098 228112
rect 140056 227769 140084 228103
rect 140042 227760 140098 227769
rect 140042 227695 140098 227704
rect 140042 217152 140098 217161
rect 140042 217087 140098 217096
rect 140056 216753 140084 217087
rect 140042 216744 140098 216753
rect 140042 216679 140098 216688
rect 140042 170232 140098 170241
rect 140042 170167 140098 170176
rect 140056 169833 140084 170167
rect 140042 169824 140098 169833
rect 140042 169759 140098 169768
rect 140042 76392 140098 76401
rect 140042 76327 140098 76336
rect 140056 75993 140084 76327
rect 140042 75984 140098 75993
rect 140042 75919 140098 75928
rect 143552 4282 143580 320062
rect 146588 317490 146616 320076
rect 147692 320062 148534 320090
rect 146576 317484 146628 317490
rect 146576 317426 146628 317432
rect 147588 263832 147640 263838
rect 147586 263800 147588 263809
rect 147640 263800 147642 263809
rect 147586 263735 147642 263744
rect 147588 227928 147640 227934
rect 147586 227896 147588 227905
rect 147640 227896 147642 227905
rect 147586 227831 147642 227840
rect 147588 216912 147640 216918
rect 147586 216880 147588 216889
rect 147640 216880 147642 216889
rect 147586 216815 147642 216824
rect 147588 169992 147640 169998
rect 147586 169960 147588 169969
rect 147640 169960 147642 169969
rect 147586 169895 147642 169904
rect 147588 76152 147640 76158
rect 147586 76120 147588 76129
rect 147640 76120 147642 76129
rect 147586 76055 147642 76064
rect 143540 4276 143592 4282
rect 143540 4218 143592 4224
rect 147692 3058 147720 320062
rect 150452 4350 150480 320076
rect 151832 320062 152398 320090
rect 153212 320062 154330 320090
rect 155972 320062 156262 320090
rect 157352 320062 158194 320090
rect 150440 4344 150492 4350
rect 150440 4286 150492 4292
rect 151832 3194 151860 320062
rect 151820 3188 151872 3194
rect 151820 3130 151872 3136
rect 153212 3126 153240 320062
rect 154486 263936 154542 263945
rect 154486 263871 154542 263880
rect 154500 263838 154528 263871
rect 154488 263832 154540 263838
rect 154488 263774 154540 263780
rect 154486 228032 154542 228041
rect 154486 227967 154542 227976
rect 154500 227934 154528 227967
rect 154488 227928 154540 227934
rect 154488 227870 154540 227876
rect 154486 217016 154542 217025
rect 154486 216951 154542 216960
rect 154500 216918 154528 216951
rect 154488 216912 154540 216918
rect 154488 216854 154540 216860
rect 154486 170096 154542 170105
rect 154486 170031 154542 170040
rect 154500 169998 154528 170031
rect 154488 169992 154540 169998
rect 154488 169934 154540 169940
rect 154486 76256 154542 76265
rect 154486 76191 154542 76200
rect 154500 76158 154528 76191
rect 154488 76152 154540 76158
rect 154488 76094 154540 76100
rect 155972 4418 156000 320062
rect 157352 6458 157380 320062
rect 160204 317694 160232 320076
rect 161492 320062 162150 320090
rect 162872 320062 164082 320090
rect 160192 317688 160244 317694
rect 160192 317630 160244 317636
rect 157340 6452 157392 6458
rect 157340 6394 157392 6400
rect 161492 4486 161520 320062
rect 161480 4480 161532 4486
rect 161480 4422 161532 4428
rect 155960 4412 156012 4418
rect 155960 4354 156012 4360
rect 162872 3262 162900 320062
rect 166000 317762 166028 320076
rect 167012 320062 167946 320090
rect 165988 317756 166040 317762
rect 165988 317698 166040 317704
rect 167012 4554 167040 320062
rect 169864 317830 169892 320076
rect 171152 320062 171902 320090
rect 172532 320062 173834 320090
rect 175292 320062 175766 320090
rect 169852 317824 169904 317830
rect 169852 317766 169904 317772
rect 167000 4548 167052 4554
rect 167000 4490 167052 4496
rect 171152 3330 171180 320062
rect 172532 4622 172560 320062
rect 172520 4616 172572 4622
rect 172520 4558 172572 4564
rect 175292 3398 175320 320062
rect 177684 317898 177712 320076
rect 179432 320062 179630 320090
rect 177672 317892 177724 317898
rect 177672 317834 177724 317840
rect 179432 4690 179460 320062
rect 181548 317966 181576 320076
rect 181536 317960 181588 317966
rect 181536 317902 181588 317908
rect 179420 4684 179472 4690
rect 179420 4626 179472 4632
rect 183572 3777 183600 320076
rect 184952 320062 185518 320090
rect 186332 320062 187450 320090
rect 184952 4758 184980 320062
rect 184940 4752 184992 4758
rect 184940 4694 184992 4700
rect 186332 4146 186360 320062
rect 189368 318034 189396 320076
rect 190472 320062 191314 320090
rect 189356 318028 189408 318034
rect 189356 317970 189408 317976
rect 190472 5506 190500 320062
rect 193232 318782 193260 320076
rect 194612 320062 195178 320090
rect 195992 320062 197202 320090
rect 198752 320062 199134 320090
rect 193220 318776 193272 318782
rect 193220 318718 193272 318724
rect 190460 5500 190512 5506
rect 190460 5442 190512 5448
rect 186320 4140 186372 4146
rect 186320 4082 186372 4088
rect 194612 4078 194640 320062
rect 195992 5438 196020 320062
rect 195980 5432 196032 5438
rect 195980 5374 196032 5380
rect 194600 4072 194652 4078
rect 194600 4014 194652 4020
rect 198752 4010 198780 320062
rect 201052 318714 201080 320076
rect 202892 320062 202998 320090
rect 201040 318708 201092 318714
rect 201040 318650 201092 318656
rect 202892 5370 202920 320062
rect 204916 318646 204944 320076
rect 205652 320062 206862 320090
rect 208412 320062 208886 320090
rect 209792 320062 210818 320090
rect 204904 318640 204956 318646
rect 204904 318582 204956 318588
rect 202880 5364 202932 5370
rect 202880 5306 202932 5312
rect 198740 4004 198792 4010
rect 198740 3946 198792 3952
rect 205652 3942 205680 320062
rect 208412 5273 208440 320062
rect 208398 5264 208454 5273
rect 208398 5199 208454 5208
rect 205640 3936 205692 3942
rect 205640 3878 205692 3884
rect 183558 3768 183614 3777
rect 183558 3703 183614 3712
rect 209792 3641 209820 320062
rect 212736 318578 212764 320076
rect 213932 320062 214682 320090
rect 212724 318572 212776 318578
rect 212724 318514 212776 318520
rect 213932 5137 213960 320062
rect 216600 318510 216628 320076
rect 218072 320062 218546 320090
rect 219452 320062 220570 320090
rect 222212 320062 222502 320090
rect 216588 318504 216640 318510
rect 216588 318446 216640 318452
rect 213918 5128 213974 5137
rect 213918 5063 213974 5072
rect 218072 3874 218100 320062
rect 219452 5302 219480 320062
rect 219440 5296 219492 5302
rect 219440 5238 219492 5244
rect 218060 3868 218112 3874
rect 218060 3810 218112 3816
rect 209778 3632 209834 3641
rect 209778 3567 209834 3576
rect 222212 3505 222240 320062
rect 224420 318374 224448 320076
rect 224408 318368 224460 318374
rect 224408 318310 224460 318316
rect 226352 5001 226380 320076
rect 228284 318306 228312 320076
rect 229112 320062 230230 320090
rect 231872 320062 232254 320090
rect 228272 318300 228324 318306
rect 228272 318242 228324 318248
rect 226338 4992 226394 5001
rect 226338 4927 226394 4936
rect 222198 3496 222254 3505
rect 222198 3431 222254 3440
rect 175280 3392 175332 3398
rect 229112 3369 229140 320062
rect 231872 5234 231900 320062
rect 234172 318238 234200 320076
rect 234160 318232 234212 318238
rect 234160 318174 234212 318180
rect 236104 318170 236132 320076
rect 237392 320062 238050 320090
rect 238772 320062 239982 320090
rect 241532 320062 241914 320090
rect 242912 320062 243846 320090
rect 236092 318164 236144 318170
rect 236092 318106 236144 318112
rect 237392 6390 237420 320062
rect 237380 6384 237432 6390
rect 237380 6326 237432 6332
rect 231860 5228 231912 5234
rect 231860 5170 231912 5176
rect 238772 3806 238800 320062
rect 238760 3800 238812 3806
rect 238760 3742 238812 3748
rect 241532 3738 241560 320062
rect 242912 6322 242940 320062
rect 245856 318102 245884 320076
rect 247788 318345 247816 320076
rect 248432 320062 249734 320090
rect 251192 320062 251666 320090
rect 252572 320062 253598 320090
rect 247774 318336 247830 318345
rect 247774 318271 247830 318280
rect 245844 318096 245896 318102
rect 245844 318038 245896 318044
rect 242900 6316 242952 6322
rect 242900 6258 242952 6264
rect 248432 6254 248460 320062
rect 248420 6248 248472 6254
rect 248420 6190 248472 6196
rect 241520 3732 241572 3738
rect 241520 3674 241572 3680
rect 251192 3602 251220 320062
rect 252572 3670 252600 320062
rect 255516 318442 255544 320076
rect 255504 318436 255556 318442
rect 255504 318378 255556 318384
rect 257540 318209 257568 320076
rect 257526 318200 257582 318209
rect 257526 318135 257582 318144
rect 259472 318073 259500 320076
rect 260852 320062 261418 320090
rect 262232 320062 263350 320090
rect 264992 320062 265282 320090
rect 266372 320062 267214 320090
rect 269132 320062 269238 320090
rect 270512 320062 271170 320090
rect 271892 320062 273102 320090
rect 274652 320062 275034 320090
rect 276032 320062 276966 320090
rect 278792 320062 278898 320090
rect 259458 318064 259514 318073
rect 259458 317999 259514 318008
rect 260852 6186 260880 320062
rect 260840 6180 260892 6186
rect 260840 6122 260892 6128
rect 252560 3664 252612 3670
rect 252560 3606 252612 3612
rect 251180 3596 251232 3602
rect 251180 3538 251232 3544
rect 262232 3534 262260 320062
rect 262220 3528 262272 3534
rect 262220 3470 262272 3476
rect 264992 3466 265020 320062
rect 266372 5166 266400 320062
rect 266360 5160 266412 5166
rect 266360 5102 266412 5108
rect 269132 5098 269160 320062
rect 269120 5092 269172 5098
rect 269120 5034 269172 5040
rect 270512 4962 270540 320062
rect 271892 5030 271920 320062
rect 271880 5024 271932 5030
rect 271880 4966 271932 4972
rect 270500 4956 270552 4962
rect 270500 4898 270552 4904
rect 274652 4865 274680 320062
rect 276032 4894 276060 320062
rect 276020 4888 276072 4894
rect 274638 4856 274694 4865
rect 276020 4830 276072 4836
rect 278792 4826 278820 320062
rect 338040 318782 338068 320962
rect 339774 320648 339830 320657
rect 339774 320583 339830 320592
rect 349986 320648 350042 320657
rect 349986 320583 350042 320592
rect 339788 320385 339816 320583
rect 350000 320385 350028 320583
rect 416424 320482 416452 323983
rect 419552 320958 419580 390623
rect 580170 346080 580226 346089
rect 580170 346015 580226 346024
rect 419906 332616 419962 332625
rect 419906 332551 419962 332560
rect 419814 328672 419870 328681
rect 419814 328607 419870 328616
rect 419722 327176 419778 327185
rect 419722 327111 419778 327120
rect 419630 325816 419686 325825
rect 419630 325751 419686 325760
rect 419540 320952 419592 320958
rect 419540 320894 419592 320900
rect 419644 320550 419672 325751
rect 419736 320618 419764 327111
rect 419828 320890 419856 328607
rect 419816 320884 419868 320890
rect 419816 320826 419868 320832
rect 419724 320612 419776 320618
rect 419724 320554 419776 320560
rect 419632 320544 419684 320550
rect 419632 320486 419684 320492
rect 416412 320476 416464 320482
rect 416412 320418 416464 320424
rect 339774 320376 339830 320385
rect 339774 320311 339830 320320
rect 349986 320376 350042 320385
rect 419920 320346 419948 332551
rect 420182 331256 420238 331265
rect 420182 331191 420238 331200
rect 419998 329896 420054 329905
rect 419998 329831 420054 329840
rect 349986 320311 350042 320320
rect 419908 320340 419960 320346
rect 419908 320282 419960 320288
rect 420012 320278 420040 329831
rect 420196 320414 420224 331191
rect 579986 322688 580042 322697
rect 579986 322623 580042 322632
rect 580000 320657 580028 322623
rect 580184 320754 580212 346015
rect 580172 320748 580224 320754
rect 580172 320690 580224 320696
rect 579986 320648 580042 320657
rect 579986 320583 580042 320592
rect 580276 320521 580304 463383
rect 580354 451752 580410 451761
rect 580354 451687 580410 451696
rect 580262 320512 580318 320521
rect 580262 320447 580318 320456
rect 420184 320408 420236 320414
rect 420184 320350 420236 320356
rect 420000 320272 420052 320278
rect 420000 320214 420052 320220
rect 580368 319938 580396 451687
rect 580446 439920 580502 439929
rect 580446 439855 580502 439864
rect 580460 320006 580488 439855
rect 580538 416528 580594 416537
rect 580538 416463 580594 416472
rect 580552 320929 580580 416463
rect 580630 404832 580686 404841
rect 580630 404767 580686 404776
rect 580538 320920 580594 320929
rect 580538 320855 580594 320864
rect 580644 320074 580672 404767
rect 580722 393000 580778 393009
rect 580722 392935 580778 392944
rect 580736 320686 580764 392935
rect 580814 369608 580870 369617
rect 580814 369543 580870 369552
rect 580724 320680 580776 320686
rect 580724 320622 580776 320628
rect 580828 320142 580856 369543
rect 580906 357912 580962 357921
rect 580906 357847 580962 357856
rect 580920 320822 580948 357847
rect 580908 320816 580960 320822
rect 580908 320758 580960 320764
rect 580816 320136 580868 320142
rect 580816 320078 580868 320084
rect 580632 320068 580684 320074
rect 580632 320010 580684 320016
rect 580448 320000 580500 320006
rect 580448 319942 580500 319948
rect 580356 319932 580408 319938
rect 580356 319874 580408 319880
rect 344020 318782 344048 318813
rect 338028 318776 338080 318782
rect 344008 318776 344060 318782
rect 338028 318718 338080 318724
rect 344006 318744 344008 318753
rect 344060 318744 344062 318753
rect 344006 318679 344062 318688
rect 344020 318102 344048 318679
rect 347778 318472 347834 318481
rect 347778 318407 347834 318416
rect 347792 318102 347820 318407
rect 344008 318096 344060 318102
rect 344008 318038 344060 318044
rect 347780 318096 347832 318102
rect 347780 318038 347832 318044
rect 580172 311840 580224 311846
rect 580172 311782 580224 311788
rect 580184 310865 580212 311782
rect 580170 310856 580226 310865
rect 580170 310791 580226 310800
rect 579804 299464 579856 299470
rect 579804 299406 579856 299412
rect 579816 299169 579844 299406
rect 579802 299160 579858 299169
rect 579802 299095 579858 299104
rect 580172 276004 580224 276010
rect 580172 275946 580224 275952
rect 580184 275777 580212 275946
rect 580170 275768 580226 275777
rect 580170 275703 580226 275712
rect 579804 252544 579856 252550
rect 579804 252486 579856 252492
rect 579816 252249 579844 252486
rect 579802 252240 579858 252249
rect 579802 252175 579858 252184
rect 579804 205624 579856 205630
rect 579804 205566 579856 205572
rect 579816 205329 579844 205566
rect 579802 205320 579858 205329
rect 579802 205255 579858 205264
rect 579804 158704 579856 158710
rect 579804 158646 579856 158652
rect 579816 158409 579844 158646
rect 579802 158400 579858 158409
rect 579802 158335 579858 158344
rect 580172 135244 580224 135250
rect 580172 135186 580224 135192
rect 580184 134881 580212 135186
rect 580170 134872 580226 134881
rect 580170 134807 580226 134816
rect 580172 124160 580224 124166
rect 580172 124102 580224 124108
rect 580184 123185 580212 124102
rect 580170 123176 580226 123185
rect 580170 123111 580226 123120
rect 579804 111784 579856 111790
rect 579804 111726 579856 111732
rect 579816 111489 579844 111726
rect 579802 111480 579858 111489
rect 579802 111415 579858 111424
rect 580172 88324 580224 88330
rect 580172 88266 580224 88272
rect 580184 87961 580212 88266
rect 580170 87952 580226 87961
rect 580170 87887 580226 87896
rect 579804 64864 579856 64870
rect 579804 64806 579856 64812
rect 579816 64569 579844 64806
rect 579802 64560 579858 64569
rect 579802 64495 579858 64504
rect 580172 41404 580224 41410
rect 580172 41346 580224 41352
rect 580184 41041 580212 41346
rect 580170 41032 580226 41041
rect 580170 40967 580226 40976
rect 580172 30320 580224 30326
rect 580172 30262 580224 30268
rect 580184 29345 580212 30262
rect 580170 29336 580226 29345
rect 580170 29271 580226 29280
rect 579804 17944 579856 17950
rect 579804 17886 579856 17892
rect 579816 17649 579844 17886
rect 579802 17640 579858 17649
rect 579802 17575 579858 17584
rect 274638 4791 274694 4800
rect 278780 4820 278832 4826
rect 278780 4762 278832 4768
rect 264980 3460 265032 3466
rect 264980 3402 265032 3408
rect 175280 3334 175332 3340
rect 229098 3360 229154 3369
rect 171140 3324 171192 3330
rect 229098 3295 229154 3304
rect 171140 3266 171192 3272
rect 162860 3256 162912 3262
rect 162860 3198 162912 3204
rect 153200 3120 153252 3126
rect 153200 3062 153252 3068
rect 147680 3052 147732 3058
rect 147680 2994 147732 3000
rect 139400 2984 139452 2990
rect 139400 2926 139452 2932
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 13606 -960 13718 480
rect 14802 -960 14914 480
rect 15998 -960 16110 480
rect 17194 -960 17306 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 27866 -960 27978 480
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44518 -960 44630 480
rect 45714 -960 45826 480
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49302 -960 49414 480
rect 50498 -960 50610 480
rect 51602 -960 51714 480
rect 52798 -960 52910 480
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 56386 -960 56498 480
rect 57582 -960 57694 480
rect 58778 -960 58890 480
rect 59974 -960 60086 480
rect 61170 -960 61282 480
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64758 -960 64870 480
rect 65954 -960 66066 480
rect 67150 -960 67262 480
rect 68254 -960 68366 480
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 73038 -960 73150 480
rect 74234 -960 74346 480
rect 75430 -960 75542 480
rect 76626 -960 76738 480
rect 77822 -960 77934 480
rect 79018 -960 79130 480
rect 80214 -960 80326 480
rect 81410 -960 81522 480
rect 82606 -960 82718 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 88494 -960 88606 480
rect 89690 -960 89802 480
rect 90886 -960 90998 480
rect 92082 -960 92194 480
rect 93278 -960 93390 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 107538 -960 107650 480
rect 108734 -960 108846 480
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 151514 -960 151626 480
rect 152710 -960 152822 480
rect 153906 -960 154018 480
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157494 -960 157606 480
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 162278 -960 162390 480
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 189602 -960 189714 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197974 -960 198086 480
rect 199170 -960 199282 480
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246734 -960 246846 480
rect 247930 -960 248042 480
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 252622 -960 252734 480
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259798 -960 259910 480
rect 260994 -960 261106 480
rect 262190 -960 262302 480
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 268078 -960 268190 480
rect 269274 -960 269386 480
rect 270470 -960 270582 480
rect 271666 -960 271778 480
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 280038 -960 280150 480
rect 281234 -960 281346 480
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 289514 -960 289626 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436990 -960 437102 480
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441774 -960 441886 480
rect 442970 -960 443082 480
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 459622 -960 459734 480
rect 460818 -960 460930 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509578 -960 509690 480
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528622 -960 528734 480
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 569010 -960 569122 480
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 682216 3478 682272
rect 3054 653520 3110 653576
rect 3330 595992 3386 596048
rect 2870 481072 2926 481128
rect 3514 667956 3570 667992
rect 3514 667936 3516 667956
rect 3516 667936 3568 667956
rect 3568 667936 3570 667956
rect 3514 624824 3570 624880
rect 3606 610408 3662 610464
rect 3606 567296 3662 567352
rect 3698 553016 3754 553072
rect 3790 538600 3846 538656
rect 4066 509904 4122 509960
rect 3974 495508 4030 495544
rect 3974 495488 3976 495508
rect 3976 495488 4028 495508
rect 4028 495488 4030 495508
rect 3422 452376 3478 452432
rect 3974 437960 4030 438016
rect 3882 423680 3938 423736
rect 3146 394984 3202 395040
rect 3238 380568 3294 380624
rect 3146 366152 3202 366208
rect 3422 337456 3478 337512
rect 3238 323040 3294 323096
rect 3330 308760 3386 308816
rect 3422 294344 3478 294400
rect 3422 280100 3424 280120
rect 3424 280100 3476 280120
rect 3476 280100 3478 280120
rect 3422 280064 3478 280100
rect 2870 265648 2926 265704
rect 3422 251232 3478 251288
rect 3422 236952 3478 237008
rect 3146 222536 3202 222592
rect 2778 208156 2780 208176
rect 2780 208156 2832 208176
rect 2832 208156 2834 208176
rect 2778 208120 2834 208156
rect 2870 193840 2926 193896
rect 3238 179424 3294 179480
rect 2778 165008 2834 165064
rect 3146 150728 3202 150784
rect 3238 136312 3294 136368
rect 2778 122032 2834 122088
rect 3238 107616 3294 107672
rect 3422 93200 3478 93256
rect 2778 78920 2834 78976
rect 3330 64504 3386 64560
rect 3422 50088 3478 50144
rect 3422 35844 3424 35864
rect 3424 35844 3476 35864
rect 3476 35844 3478 35864
rect 3422 35808 3478 35844
rect 2870 21392 2926 21448
rect 3422 7112 3478 7168
rect 57610 646040 57666 646096
rect 57518 644952 57574 645008
rect 57426 643184 57482 643240
rect 57334 641960 57390 642016
rect 57242 640328 57298 640384
rect 57058 639240 57114 639296
rect 56966 579672 57022 579728
rect 56874 578312 56930 578368
rect 57150 637608 57206 637664
rect 56690 490728 56746 490784
rect 56598 488824 56654 488880
rect 56690 486920 56746 486976
rect 56690 485016 56746 485072
rect 56598 483112 56654 483168
rect 56506 479168 56562 479224
rect 56506 477264 56562 477320
rect 56506 475360 56562 475416
rect 56506 473456 56562 473512
rect 56506 471552 56562 471608
rect 56506 469512 56562 469568
rect 56506 467608 56562 467664
rect 56506 465704 56562 465760
rect 56506 463800 56562 463856
rect 56506 461896 56562 461952
rect 56690 481208 56746 481264
rect 56598 459856 56654 459912
rect 56598 457952 56654 458008
rect 56598 456048 56654 456104
rect 56598 454144 56654 454200
rect 56782 442584 56838 442640
rect 56874 436736 56930 436792
rect 57058 492768 57114 492824
rect 56966 431024 57022 431080
rect 57426 539008 57482 539064
rect 57426 537104 57482 537160
rect 57426 535200 57482 535256
rect 57426 533296 57482 533352
rect 57426 531412 57482 531448
rect 57426 531392 57428 531412
rect 57428 531392 57480 531412
rect 57480 531392 57482 531412
rect 57426 529352 57482 529408
rect 57426 527448 57482 527504
rect 57426 525544 57482 525600
rect 57426 523640 57482 523696
rect 57426 521756 57482 521792
rect 57426 521736 57428 521756
rect 57428 521736 57480 521756
rect 57480 521736 57482 521756
rect 57426 519696 57482 519752
rect 57426 517792 57482 517848
rect 57426 515888 57482 515944
rect 57426 513984 57482 514040
rect 57426 512080 57482 512136
rect 57426 510040 57482 510096
rect 57426 508136 57482 508192
rect 57242 506232 57298 506288
rect 57150 382744 57206 382800
rect 56966 371184 57022 371240
rect 56874 361528 56930 361584
rect 56690 359488 56746 359544
rect 56598 357584 56654 357640
rect 56782 355680 56838 355736
rect 57058 365336 57114 365392
rect 57150 351872 57206 351928
rect 57058 328616 57114 328672
rect 57426 504328 57482 504384
rect 57426 502424 57482 502480
rect 57334 500384 57390 500440
rect 57426 498480 57482 498536
rect 57426 496576 57482 496632
rect 57426 494672 57482 494728
rect 57518 380704 57574 380760
rect 57702 448296 57758 448352
rect 57794 440544 57850 440600
rect 57886 428984 57942 429040
rect 57978 415520 58034 415576
rect 58070 400016 58126 400072
rect 58162 392400 58218 392456
rect 58346 452240 58402 452296
rect 58438 450200 58494 450256
rect 58530 446392 58586 446448
rect 58622 444488 58678 444544
rect 58714 438640 58770 438696
rect 58806 434832 58862 434888
rect 58898 432928 58954 432984
rect 58990 427080 59046 427136
rect 59082 423272 59138 423328
rect 59174 421368 59230 421424
rect 59266 417424 59322 417480
rect 77206 697176 77262 697232
rect 96526 697176 96582 697232
rect 70306 697076 70308 697096
rect 70308 697076 70360 697096
rect 70360 697076 70362 697096
rect 70306 697040 70362 697076
rect 89626 697076 89628 697096
rect 89628 697076 89680 697096
rect 89680 697076 89682 697096
rect 89626 697040 89682 697076
rect 115846 697176 115902 697232
rect 135166 697176 135222 697232
rect 108946 697076 108948 697096
rect 108948 697076 109000 697096
rect 109000 697076 109002 697096
rect 108946 697040 109002 697076
rect 128266 697076 128268 697096
rect 128268 697076 128320 697096
rect 128320 697076 128322 697096
rect 128266 697040 128322 697076
rect 129278 652840 129334 652896
rect 133694 652840 133750 652896
rect 135166 650936 135222 650992
rect 120722 650800 120778 650856
rect 89626 650664 89682 650720
rect 106738 650664 106794 650720
rect 96526 650564 96528 650584
rect 96528 650564 96580 650584
rect 96580 650564 96582 650584
rect 96526 650528 96582 650564
rect 115754 650564 115756 650584
rect 115756 650564 115808 650584
rect 115808 650564 115810 650584
rect 115754 650528 115810 650564
rect 115938 650548 115994 650584
rect 115938 650528 115940 650548
rect 115940 650528 115992 650548
rect 115992 650528 115994 650548
rect 135166 650528 135222 650584
rect 67546 558864 67602 558920
rect 68926 558864 68982 558920
rect 70306 558864 70362 558920
rect 71686 558864 71742 558920
rect 72606 558864 72662 558920
rect 73066 558864 73122 558920
rect 73802 558864 73858 558920
rect 74262 558864 74318 558920
rect 74998 558864 75054 558920
rect 76010 558864 76066 558920
rect 76838 558864 76894 558920
rect 77390 558864 77446 558920
rect 78494 558864 78550 558920
rect 79414 558864 79470 558920
rect 79966 558864 80022 558920
rect 80794 558864 80850 558920
rect 81254 558864 81310 558920
rect 81898 558864 81954 558920
rect 82726 558864 82782 558920
rect 83830 558864 83886 558920
rect 84198 558864 84254 558920
rect 85486 558864 85542 558920
rect 86406 558864 86462 558920
rect 86866 558864 86922 558920
rect 87878 558864 87934 558920
rect 88246 558864 88302 558920
rect 88890 558864 88946 558920
rect 89626 558864 89682 558920
rect 89810 558864 89866 558920
rect 91006 558864 91062 558920
rect 92478 558864 92534 558920
rect 93674 558864 93730 558920
rect 94870 558864 94926 558920
rect 95146 558864 95202 558920
rect 95790 558864 95846 558920
rect 96526 558864 96582 558920
rect 96986 558864 97042 558920
rect 97814 558864 97870 558920
rect 98090 558864 98146 558920
rect 99286 558864 99342 558920
rect 99562 558864 99618 558920
rect 100390 558864 100446 558920
rect 102046 558864 102102 558920
rect 103426 558864 103482 558920
rect 104806 558864 104862 558920
rect 105542 558864 105598 558920
rect 106186 558864 106242 558920
rect 107474 558864 107530 558920
rect 108486 558864 108542 558920
rect 110326 558864 110382 558920
rect 59450 425176 59506 425232
rect 59450 419328 59506 419384
rect 59358 409672 59414 409728
rect 58254 386552 58310 386608
rect 70214 558592 70270 558648
rect 75826 558184 75882 558240
rect 78586 558320 78642 558376
rect 79598 558592 79654 558648
rect 80702 545128 80758 545184
rect 80702 544856 80758 544912
rect 82818 558592 82874 558648
rect 85210 558612 85266 558648
rect 85210 558592 85212 558612
rect 85212 558592 85264 558612
rect 85264 558592 85266 558612
rect 83830 544312 83886 544368
rect 86774 558592 86830 558648
rect 85578 545300 85580 545320
rect 85580 545300 85632 545320
rect 85632 545300 85634 545320
rect 85578 545264 85634 545300
rect 85854 544448 85910 544504
rect 87970 544584 88026 544640
rect 91098 558592 91154 558648
rect 92386 558320 92442 558376
rect 93306 558628 93308 558648
rect 93308 558628 93360 558648
rect 93360 558628 93362 558648
rect 93306 558592 93362 558628
rect 92110 544720 92166 544776
rect 93766 558592 93822 558648
rect 95054 545300 95056 545320
rect 95056 545300 95108 545320
rect 95108 545300 95110 545320
rect 95054 545264 95110 545300
rect 97998 558340 98054 558376
rect 97998 558320 98000 558340
rect 98000 558320 98052 558340
rect 98052 558320 98054 558340
rect 96618 545284 96674 545320
rect 96618 545264 96620 545284
rect 96620 545264 96672 545284
rect 96672 545264 96674 545284
rect 100022 558592 100078 558648
rect 101954 558592 102010 558648
rect 101402 558320 101458 558376
rect 102782 558592 102838 558648
rect 103886 558612 103942 558648
rect 103886 558592 103888 558612
rect 103888 558592 103940 558612
rect 103940 558592 103942 558612
rect 104806 545128 104862 545184
rect 106922 558592 106978 558648
rect 106186 542952 106242 543008
rect 107750 558592 107806 558648
rect 108302 558592 108358 558648
rect 115938 545420 115994 545456
rect 115938 545400 115940 545420
rect 115940 545400 115992 545420
rect 115992 545400 115994 545420
rect 125414 545128 125470 545184
rect 135258 545420 135314 545456
rect 135258 545400 135260 545420
rect 135260 545400 135312 545420
rect 135312 545400 135314 545420
rect 154486 697176 154542 697232
rect 147586 697076 147588 697096
rect 147588 697076 147640 697096
rect 147640 697076 147642 697096
rect 147586 697040 147642 697076
rect 166906 697076 166908 697096
rect 166908 697076 166960 697096
rect 166960 697076 166962 697096
rect 166906 697040 166962 697076
rect 173806 697176 173862 697232
rect 193126 697176 193182 697232
rect 212446 697176 212502 697232
rect 231766 697176 231822 697232
rect 251086 697176 251142 697232
rect 270406 697176 270462 697232
rect 289726 697176 289782 697232
rect 186226 697076 186228 697096
rect 186228 697076 186280 697096
rect 186280 697076 186282 697096
rect 186226 697040 186282 697076
rect 205546 697076 205548 697096
rect 205548 697076 205600 697096
rect 205600 697076 205602 697096
rect 205546 697040 205602 697076
rect 224866 697076 224868 697096
rect 224868 697076 224920 697096
rect 224920 697076 224922 697096
rect 224866 697040 224922 697076
rect 244186 697076 244188 697096
rect 244188 697076 244240 697096
rect 244240 697076 244242 697096
rect 244186 697040 244242 697076
rect 263506 697076 263508 697096
rect 263508 697076 263560 697096
rect 263560 697076 263562 697096
rect 263506 697040 263562 697076
rect 282826 697076 282828 697096
rect 282828 697076 282880 697096
rect 282880 697076 282882 697096
rect 282826 697040 282882 697076
rect 166906 686296 166962 686352
rect 167090 686296 167146 686352
rect 154578 686180 154634 686216
rect 154578 686160 154580 686180
rect 154580 686160 154632 686180
rect 154632 686160 154634 686180
rect 188342 686432 188398 686488
rect 173898 686316 173954 686352
rect 173898 686296 173900 686316
rect 173900 686296 173952 686316
rect 173952 686296 173954 686316
rect 178774 686160 178830 686216
rect 188342 686160 188398 686216
rect 289818 686180 289874 686216
rect 289818 686160 289820 686180
rect 289820 686160 289872 686180
rect 289872 686160 289874 686180
rect 162214 685888 162270 685944
rect 294510 685888 294566 685944
rect 309046 697176 309102 697232
rect 328366 697176 328422 697232
rect 302146 697076 302148 697096
rect 302148 697076 302200 697096
rect 302200 697076 302202 697096
rect 302146 697040 302202 697076
rect 321466 697076 321468 697096
rect 321468 697076 321520 697096
rect 321520 697076 321522 697096
rect 321466 697040 321522 697076
rect 360106 686296 360162 686352
rect 360290 686296 360346 686352
rect 347778 686180 347834 686216
rect 347778 686160 347780 686180
rect 347780 686160 347832 686180
rect 347832 686160 347834 686180
rect 355414 685888 355470 685944
rect 166998 673920 167054 673976
rect 154578 673804 154634 673840
rect 154578 673784 154580 673804
rect 154580 673784 154632 673804
rect 154632 673784 154634 673804
rect 162214 673512 162270 673568
rect 166906 673512 166962 673568
rect 188342 674056 188398 674112
rect 173898 673940 173954 673976
rect 173898 673920 173900 673940
rect 173900 673920 173952 673940
rect 173952 673920 173954 673940
rect 178774 673784 178830 673840
rect 188342 673784 188398 673840
rect 289818 673804 289874 673840
rect 289818 673784 289820 673804
rect 289820 673784 289872 673804
rect 289872 673784 289874 673804
rect 292670 673512 292726 673568
rect 360106 673920 360162 673976
rect 360290 673920 360346 673976
rect 347778 673804 347834 673840
rect 347778 673784 347780 673804
rect 347780 673784 347832 673804
rect 347832 673784 347834 673804
rect 355414 673512 355470 673568
rect 379518 686432 379574 686488
rect 367098 686316 367154 686352
rect 367098 686296 367100 686316
rect 367100 686296 367152 686316
rect 367152 686296 367154 686316
rect 371974 686160 372030 686216
rect 379518 686160 379574 686216
rect 427542 686160 427598 686216
rect 427726 686160 427782 686216
rect 379518 674056 379574 674112
rect 367098 673940 367154 673976
rect 367098 673920 367100 673940
rect 367100 673920 367152 673940
rect 367152 673920 367154 673940
rect 371974 673784 372030 673840
rect 379518 673784 379574 673840
rect 441526 686432 441582 686488
rect 441526 686160 441582 686216
rect 137650 649655 137706 649711
rect 140042 650936 140098 650992
rect 140134 650664 140190 650720
rect 258630 652840 258686 652896
rect 263506 651616 263562 651672
rect 278778 650700 278780 650720
rect 278780 650700 278832 650720
rect 278832 650700 278834 650720
rect 278778 650664 278834 650700
rect 292670 650664 292726 650720
rect 237378 650548 237434 650584
rect 237378 650528 237380 650548
rect 237380 650528 237432 650548
rect 237432 650528 237434 650548
rect 237562 650528 237618 650584
rect 288346 650528 288402 650584
rect 289818 650548 289874 650584
rect 289818 650528 289820 650548
rect 289820 650528 289872 650548
rect 289872 650528 289874 650548
rect 270498 650020 270500 650040
rect 270500 650020 270552 650040
rect 270552 650020 270554 650040
rect 270498 649984 270554 650020
rect 280066 649984 280122 650040
rect 266450 649848 266506 649904
rect 188342 646040 188398 646096
rect 188250 637608 188306 637664
rect 139398 589600 139454 589656
rect 141514 543224 141570 543280
rect 144826 545128 144882 545184
rect 144182 543088 144238 543144
rect 166906 545300 166908 545320
rect 166908 545300 166960 545320
rect 166960 545300 166962 545320
rect 166906 545264 166962 545300
rect 177302 545300 177304 545320
rect 177304 545300 177356 545320
rect 177356 545300 177358 545320
rect 177302 545264 177358 545300
rect 188434 644952 188490 645008
rect 188526 643184 188582 643240
rect 188618 641960 188674 642016
rect 188526 544720 188582 544776
rect 188710 640328 188766 640384
rect 188894 639240 188950 639296
rect 188802 579672 188858 579728
rect 188710 544584 188766 544640
rect 269118 589328 269174 589384
rect 270406 589348 270462 589384
rect 270406 589328 270408 589348
rect 270408 589328 270460 589348
rect 270460 589328 270462 589348
rect 269118 587696 269174 587752
rect 188986 578312 189042 578368
rect 210974 559952 211030 560008
rect 195978 558864 196034 558920
rect 197358 558884 197414 558920
rect 197358 558864 197360 558884
rect 197360 558864 197412 558884
rect 197412 558864 197414 558884
rect 194414 558728 194470 558784
rect 195886 545420 195942 545456
rect 195886 545400 195888 545420
rect 195888 545400 195940 545420
rect 195940 545400 195942 545420
rect 188894 544448 188950 544504
rect 188250 544312 188306 544368
rect 201498 558864 201554 558920
rect 202786 558864 202842 558920
rect 204166 558864 204222 558920
rect 205546 558864 205602 558920
rect 206098 558864 206154 558920
rect 208398 558864 208454 558920
rect 210606 558864 210662 558920
rect 202142 558592 202198 558648
rect 198738 557660 198794 557696
rect 198738 557640 198740 557660
rect 198740 557640 198792 557660
rect 198792 557640 198794 557660
rect 200210 557796 200266 557832
rect 200210 557776 200212 557796
rect 200212 557776 200264 557796
rect 200264 557776 200266 557796
rect 201406 545420 201462 545456
rect 201406 545400 201408 545420
rect 201408 545400 201460 545420
rect 201460 545400 201462 545420
rect 203522 558728 203578 558784
rect 204902 558592 204958 558648
rect 209042 558592 209098 558648
rect 207662 557660 207718 557696
rect 207662 557640 207664 557660
rect 207664 557640 207716 557660
rect 207716 557640 207718 557660
rect 206926 557504 206982 557560
rect 207570 545672 207626 545728
rect 207570 545400 207626 545456
rect 208306 557504 208362 557560
rect 209686 557504 209742 557560
rect 208306 543224 208362 543280
rect 220082 559000 220138 559056
rect 211802 558864 211858 558920
rect 213090 558864 213146 558920
rect 213918 558864 213974 558920
rect 215298 558884 215354 558920
rect 215298 558864 215300 558884
rect 215300 558864 215352 558884
rect 215352 558864 215354 558884
rect 217966 558864 218022 558920
rect 218978 558864 219034 558920
rect 215114 558340 215170 558376
rect 215114 558320 215116 558340
rect 215116 558320 215168 558340
rect 215168 558320 215170 558340
rect 217782 558728 217838 558784
rect 211066 557640 211122 557696
rect 222382 558864 222438 558920
rect 223578 558864 223634 558920
rect 224498 558884 224554 558920
rect 224498 558864 224500 558884
rect 224500 558864 224552 558884
rect 224552 558864 224554 558884
rect 221554 558340 221610 558376
rect 221554 558320 221556 558340
rect 221556 558320 221608 558340
rect 221608 558320 221610 558340
rect 225878 558864 225934 558920
rect 227166 558864 227222 558920
rect 228178 558864 228234 558920
rect 229558 558864 229614 558920
rect 231858 558748 231914 558784
rect 231858 558728 231860 558748
rect 231860 558728 231912 558748
rect 231912 558728 231914 558748
rect 233238 558728 233294 558784
rect 234894 558612 234950 558648
rect 234894 558592 234896 558612
rect 234896 558592 234948 558612
rect 234948 558592 234950 558612
rect 237378 558592 237434 558648
rect 231950 558456 232006 558512
rect 230478 558340 230534 558376
rect 230478 558320 230480 558340
rect 230480 558320 230532 558340
rect 230532 558320 230534 558340
rect 231858 558320 231914 558376
rect 238758 558456 238814 558512
rect 229098 557796 229154 557832
rect 229098 557776 229100 557796
rect 229100 557776 229152 557796
rect 229152 557776 229154 557796
rect 238666 557776 238722 557832
rect 217874 557640 217930 557696
rect 226154 557640 226210 557696
rect 233146 557640 233202 557696
rect 212446 557504 212502 557560
rect 213826 557504 213882 557560
rect 215206 557504 215262 557560
rect 216586 557504 216642 557560
rect 206190 542952 206246 543008
rect 210422 543088 210478 543144
rect 212538 545420 212594 545456
rect 212538 545400 212540 545420
rect 212540 545400 212592 545420
rect 212592 545400 212594 545420
rect 217966 557504 218022 557560
rect 219346 557504 219402 557560
rect 220726 557504 220782 557560
rect 222106 557504 222162 557560
rect 223486 557504 223542 557560
rect 224866 557504 224922 557560
rect 222014 545128 222070 545184
rect 226246 557504 226302 557560
rect 227626 557504 227682 557560
rect 229006 557504 229062 557560
rect 230386 557504 230442 557560
rect 231766 557504 231822 557560
rect 233054 557504 233110 557560
rect 231858 545420 231914 545456
rect 231858 545400 231860 545420
rect 231860 545400 231912 545420
rect 231912 545400 231914 545420
rect 234526 557504 234582 557560
rect 235906 557504 235962 557560
rect 237286 557504 237342 557560
rect 238666 557504 238722 557560
rect 240046 557504 240102 557560
rect 241610 557504 241666 557560
rect 251086 557504 251142 557560
rect 260838 557540 260840 557560
rect 260840 557540 260892 557560
rect 260892 557540 260894 557560
rect 260838 557504 260894 557540
rect 270406 557504 270462 557560
rect 251178 545420 251234 545456
rect 251178 545400 251180 545420
rect 251180 545400 251232 545420
rect 251232 545400 251234 545420
rect 241426 545128 241482 545184
rect 260746 545128 260802 545184
rect 282366 492632 282422 492688
rect 282550 492632 282606 492688
rect 282366 473320 282422 473376
rect 282550 473320 282606 473376
rect 282366 454008 282422 454064
rect 282550 454008 282606 454064
rect 281538 429392 281594 429448
rect 281538 428440 281594 428496
rect 281630 427352 281686 427408
rect 281538 426436 281540 426456
rect 281540 426436 281592 426456
rect 281592 426436 281594 426456
rect 281538 426400 281594 426436
rect 281538 425312 281594 425368
rect 282642 425040 282698 425096
rect 283010 425040 283066 425096
rect 281538 424360 281594 424416
rect 281630 423408 281686 423464
rect 281538 422340 281594 422376
rect 281538 422320 281540 422340
rect 281540 422320 281592 422340
rect 281592 422320 281594 422340
rect 281538 421368 281594 421424
rect 281538 420280 281594 420336
rect 281630 419328 281686 419384
rect 281538 418240 281594 418296
rect 282274 416336 282330 416392
rect 281722 415248 281778 415304
rect 282090 414296 282146 414352
rect 282826 417288 282882 417344
rect 282642 413924 282644 413944
rect 282644 413924 282696 413944
rect 282696 413924 282698 413944
rect 282642 413888 282698 413924
rect 59818 413616 59874 413672
rect 59726 396208 59782 396264
rect 59634 390360 59690 390416
rect 59542 384648 59598 384704
rect 57610 378800 57666 378856
rect 57794 376896 57850 376952
rect 57702 373088 57758 373144
rect 57610 367240 57666 367296
rect 57518 363432 57574 363488
rect 57426 334464 57482 334520
rect 57886 369144 57942 369200
rect 57794 336368 57850 336424
rect 59450 349832 59506 349888
rect 59358 344120 59414 344176
rect 59082 338272 59138 338328
rect 57794 324808 57850 324864
rect 57702 322904 57758 322960
rect 57886 321000 57942 321056
rect 59174 332560 59230 332616
rect 59266 326712 59322 326768
rect 59726 330656 59782 330712
rect 281906 410216 281962 410272
rect 282090 412256 282146 412312
rect 281814 406136 281870 406192
rect 281722 405184 281778 405240
rect 281906 403144 281962 403200
rect 281630 401140 281632 401160
rect 281632 401140 281684 401160
rect 281684 401140 281686 401160
rect 281630 401104 281686 401140
rect 281630 400172 281686 400208
rect 281630 400152 281632 400172
rect 281632 400152 281684 400172
rect 281684 400152 281686 400172
rect 281630 399064 281686 399120
rect 281630 394032 281686 394088
rect 281722 393216 281778 393272
rect 281630 393116 281632 393136
rect 281632 393116 281684 393136
rect 281684 393116 281686 393136
rect 281630 393080 281686 393116
rect 281630 391992 281686 392048
rect 281630 388048 281686 388104
rect 281630 386996 281632 387016
rect 281632 386996 281684 387016
rect 281684 386996 281686 387016
rect 281630 386960 281686 386996
rect 281722 386044 281724 386064
rect 281724 386044 281776 386064
rect 281776 386044 281778 386064
rect 281722 386008 281778 386044
rect 281630 385056 281686 385112
rect 281630 383968 281686 384024
rect 281906 390088 281962 390144
rect 281630 381964 281632 381984
rect 281632 381964 281684 381984
rect 281684 381964 281686 381984
rect 281630 381928 281686 381964
rect 281722 380976 281778 381032
rect 281722 360712 281778 360768
rect 281906 357720 281962 357776
rect 281998 356768 282054 356824
rect 282458 407904 282514 407960
rect 282182 402192 282238 402248
rect 282182 398148 282184 398168
rect 282184 398148 282236 398168
rect 282236 398148 282238 398168
rect 282182 398112 282238 398148
rect 282182 376896 282238 376952
rect 282182 372816 282238 372872
rect 282182 369824 282238 369880
rect 282182 365744 282238 365800
rect 282090 355680 282146 355736
rect 282182 354728 282238 354784
rect 281998 354592 282054 354648
rect 282090 352688 282146 352744
rect 281998 351736 282054 351792
rect 282826 413244 282828 413264
rect 282828 413244 282880 413264
rect 282880 413244 282882 413264
rect 282826 413208 282882 413244
rect 282826 411204 282828 411224
rect 282828 411204 282880 411224
rect 282880 411204 282882 411224
rect 282826 411168 282882 411204
rect 283010 409264 283066 409320
rect 282918 408448 282974 408504
rect 282458 393216 282514 393272
rect 282366 354592 282422 354648
rect 282826 404268 282828 404288
rect 282828 404268 282880 404288
rect 282880 404268 282882 404288
rect 282826 404232 282882 404268
rect 282826 389000 282882 389056
rect 282826 383016 282882 383072
rect 282826 379888 282882 379944
rect 282826 378936 282882 378992
rect 282826 377984 282882 378040
rect 282826 375944 282882 376000
rect 282826 374856 282882 374912
rect 282826 373940 282828 373960
rect 282828 373940 282880 373960
rect 282880 373940 282882 373960
rect 282826 373904 282882 373940
rect 282826 371864 282882 371920
rect 282826 370912 282882 370968
rect 282826 368872 282882 368928
rect 282826 367784 282882 367840
rect 282826 366832 282882 366888
rect 282826 364792 282882 364848
rect 282826 363840 282882 363896
rect 282826 362752 282882 362808
rect 282734 361800 282790 361856
rect 282826 359760 282882 359816
rect 282734 358808 282790 358864
rect 282642 353640 282698 353696
rect 282550 350648 282606 350704
rect 282274 349696 282330 349752
rect 282826 348608 282882 348664
rect 282826 347692 282828 347712
rect 282828 347692 282880 347712
rect 282880 347692 282882 347712
rect 282826 347656 282882 347692
rect 282274 346568 282330 346624
rect 282090 345616 282146 345672
rect 282826 344664 282882 344720
rect 282734 343576 282790 343632
rect 282550 342624 282606 342680
rect 282826 341536 282882 341592
rect 282458 340584 282514 340640
rect 282090 339632 282146 339688
rect 281998 336504 282054 336560
rect 281814 334464 281870 334520
rect 281630 333548 281632 333568
rect 281632 333548 281684 333568
rect 281684 333548 281686 333568
rect 281630 333512 281686 333548
rect 281630 330520 281686 330576
rect 281538 329432 281594 329488
rect 281630 328480 281686 328536
rect 281538 327392 281594 327448
rect 281538 326440 281594 326496
rect 281906 331472 281962 331528
rect 282366 338544 282422 338600
rect 282182 332560 282238 332616
rect 281722 325488 281778 325544
rect 281538 324400 281594 324456
rect 281538 323448 281594 323504
rect 281538 322360 281594 322416
rect 279974 320864 280030 320920
rect 280066 320612 280122 320648
rect 280066 320592 280068 320612
rect 280068 320592 280120 320612
rect 280120 320592 280122 320612
rect 280066 320476 280122 320512
rect 280066 320456 280068 320476
rect 280068 320456 280120 320476
rect 280120 320456 280122 320476
rect 282550 337592 282606 337648
rect 282642 335552 282698 335608
rect 311990 650936 312046 650992
rect 309046 650800 309102 650856
rect 311806 650800 311862 650856
rect 340786 650664 340842 650720
rect 378138 652860 378194 652896
rect 378138 652840 378140 652860
rect 378140 652840 378192 652860
rect 378192 652840 378194 652860
rect 383474 652860 383530 652896
rect 383474 652840 383476 652860
rect 383476 652840 383528 652860
rect 383528 652840 383530 652860
rect 386326 651344 386382 651400
rect 370410 651072 370466 651128
rect 367098 650820 367154 650856
rect 386326 650936 386382 650992
rect 367098 650800 367100 650820
rect 367100 650800 367152 650820
rect 367152 650800 367154 650820
rect 321466 650528 321522 650584
rect 321650 650528 321706 650584
rect 347686 650564 347688 650584
rect 347688 650564 347740 650584
rect 347740 650564 347742 650584
rect 347686 650528 347742 650564
rect 309046 650392 309102 650448
rect 386418 649848 386474 649904
rect 307114 646312 307170 646368
rect 307114 644952 307170 645008
rect 307114 643456 307170 643512
rect 307666 642096 307722 642152
rect 307666 640464 307722 640520
rect 306654 639376 306710 639432
rect 306838 637880 306894 637936
rect 299662 589328 299718 589384
rect 299938 589328 299994 589384
rect 400862 651072 400918 651128
rect 389178 650936 389234 650992
rect 389270 650800 389326 650856
rect 400862 650528 400918 650584
rect 405738 650548 405794 650584
rect 405738 650528 405740 650548
rect 405740 650528 405792 650548
rect 405792 650528 405794 650548
rect 418250 650528 418306 650584
rect 418066 650256 418122 650312
rect 413374 650120 413430 650176
rect 444286 650800 444342 650856
rect 444286 650528 444342 650584
rect 456706 650428 456708 650448
rect 456708 650428 456760 650448
rect 456760 650428 456762 650448
rect 456706 650392 456762 650428
rect 387798 589600 387854 589656
rect 307022 579672 307078 579728
rect 305642 578312 305698 578368
rect 302146 545436 302148 545456
rect 302148 545436 302200 545456
rect 302200 545436 302202 545456
rect 302146 545400 302202 545436
rect 389178 580896 389234 580952
rect 309046 545536 309102 545592
rect 329102 559816 329158 559872
rect 337750 559816 337806 559872
rect 357714 559816 357770 559872
rect 313370 558864 313426 558920
rect 321558 558864 321614 558920
rect 322938 558864 322994 558920
rect 324318 558864 324374 558920
rect 325698 558864 325754 558920
rect 327078 558864 327134 558920
rect 317418 557932 317474 557968
rect 317418 557912 317420 557932
rect 317420 557912 317472 557932
rect 317472 557912 317474 557932
rect 320178 557912 320234 557968
rect 316038 557504 316094 557560
rect 318798 557504 318854 557560
rect 320270 557504 320326 557560
rect 321466 545300 321468 545320
rect 321468 545300 321520 545320
rect 321520 545300 321522 545320
rect 321466 545264 321522 545300
rect 322202 558728 322258 558784
rect 323582 558728 323638 558784
rect 324962 558728 325018 558784
rect 326342 558728 326398 558784
rect 327722 558728 327778 558784
rect 328458 558764 328460 558784
rect 328460 558764 328512 558784
rect 328512 558764 328514 558784
rect 328458 558728 328514 558764
rect 328458 558456 328514 558512
rect 328458 557096 328514 557152
rect 328366 545400 328422 545456
rect 329286 558864 329342 558920
rect 329838 558864 329894 558920
rect 330482 558864 330538 558920
rect 331218 558864 331274 558920
rect 332598 558864 332654 558920
rect 333978 558864 334034 558920
rect 335358 558864 335414 558920
rect 329930 558728 329986 558784
rect 331770 558728 331826 558784
rect 332690 558728 332746 558784
rect 334070 558728 334126 558784
rect 336738 558864 336794 558920
rect 335450 558728 335506 558784
rect 336462 558728 336518 558784
rect 348146 559272 348202 559328
rect 348054 559136 348110 559192
rect 338118 558864 338174 558920
rect 339498 558864 339554 558920
rect 341246 558864 341302 558920
rect 342534 558864 342590 558920
rect 343638 558864 343694 558920
rect 344834 558884 344890 558920
rect 344834 558864 344836 558884
rect 344836 558864 344888 558884
rect 344888 558864 344890 558884
rect 338026 558764 338028 558784
rect 338028 558764 338080 558784
rect 338080 558764 338082 558784
rect 338026 558728 338082 558764
rect 338026 558456 338082 558512
rect 336830 557912 336886 557968
rect 338026 389836 338082 389872
rect 338026 389816 338028 389836
rect 338028 389816 338080 389836
rect 338080 389816 338082 389836
rect 337382 381248 337438 381304
rect 282826 321408 282882 321464
rect 339038 558728 339094 558784
rect 339866 558728 339922 558784
rect 345754 558864 345810 558920
rect 346858 558864 346914 558920
rect 345662 558456 345718 558512
rect 348054 558592 348110 558648
rect 348238 558864 348294 558920
rect 349526 558864 349582 558920
rect 351734 558864 351790 558920
rect 350538 558456 350594 558512
rect 353298 558728 353354 558784
rect 354678 558728 354734 558784
rect 356058 558728 356114 558784
rect 357438 558456 357494 558512
rect 351734 558184 351790 558240
rect 351918 558204 351974 558240
rect 351918 558184 351920 558204
rect 351920 558184 351972 558204
rect 351972 558184 351974 558204
rect 354678 558184 354734 558240
rect 345662 558048 345718 558104
rect 351918 558048 351974 558104
rect 353298 557912 353354 557968
rect 343730 557640 343786 557696
rect 340878 557504 340934 557560
rect 342258 557504 342314 557560
rect 343638 557504 343694 557560
rect 345018 557504 345074 557560
rect 346398 557504 346454 557560
rect 347778 557504 347834 557560
rect 349158 557504 349214 557560
rect 350630 557504 350686 557560
rect 347686 545400 347742 545456
rect 347686 545264 347742 545320
rect 371882 545536 371938 545592
rect 367006 545264 367062 545320
rect 371882 545128 371938 545184
rect 367006 544856 367062 544912
rect 543462 700304 543518 700360
rect 553306 697312 553362 697368
rect 553490 697312 553546 697368
rect 540978 697196 541034 697232
rect 540978 697176 540980 697196
rect 540980 697176 541032 697196
rect 541032 697176 541034 697196
rect 548614 696904 548670 696960
rect 553306 686296 553362 686352
rect 553490 686296 553546 686352
rect 540978 686180 541034 686216
rect 540978 686160 540980 686180
rect 540980 686160 541032 686180
rect 541032 686160 541034 686180
rect 548614 685888 548670 685944
rect 560298 697332 560354 697368
rect 560298 697312 560300 697332
rect 560300 697312 560352 697332
rect 560352 697312 560354 697332
rect 565174 697176 565230 697232
rect 572718 697176 572774 697232
rect 572626 697040 572682 697096
rect 560298 686316 560354 686352
rect 560298 686296 560300 686316
rect 560300 686296 560352 686316
rect 560352 686296 560354 686316
rect 565174 686160 565230 686216
rect 572718 686160 572774 686216
rect 572626 686024 572682 686080
rect 559010 684392 559066 684448
rect 559010 684256 559066 684312
rect 553398 673920 553454 673976
rect 540978 673804 541034 673840
rect 540978 673784 540980 673804
rect 540980 673784 541032 673804
rect 541032 673784 541034 673804
rect 548614 673512 548670 673568
rect 553306 673512 553362 673568
rect 560298 673940 560354 673976
rect 560298 673920 560300 673940
rect 560300 673920 560352 673940
rect 560352 673920 560354 673940
rect 565174 673784 565230 673840
rect 572718 673784 572774 673840
rect 572626 673648 572682 673704
rect 463606 650528 463662 650584
rect 482926 650528 482982 650584
rect 476026 650428 476028 650448
rect 476028 650428 476080 650448
rect 476080 650428 476082 650448
rect 476026 650392 476082 650428
rect 502246 650528 502302 650584
rect 521566 650528 521622 650584
rect 540886 650548 540942 650584
rect 540886 650528 540888 650548
rect 540888 650528 540940 650548
rect 540940 650528 540942 650548
rect 495346 650428 495348 650448
rect 495348 650428 495400 650448
rect 495400 650428 495402 650448
rect 495346 650392 495402 650428
rect 514666 650428 514668 650448
rect 514668 650428 514720 650448
rect 514720 650428 514722 650448
rect 514666 650392 514722 650428
rect 533986 650392 534042 650448
rect 583390 651072 583446 651128
rect 563150 650800 563206 650856
rect 583390 650800 583446 650856
rect 572626 650700 572628 650720
rect 572628 650700 572680 650720
rect 572680 650700 572682 650720
rect 572626 650664 572682 650700
rect 579526 650700 579528 650720
rect 579528 650700 579580 650720
rect 579580 650700 579582 650720
rect 579526 650664 579582 650700
rect 560298 650564 560300 650584
rect 560300 650564 560352 650584
rect 560352 650564 560354 650584
rect 560298 650528 560354 650564
rect 580262 639376 580318 639432
rect 580170 557232 580226 557288
rect 491758 549208 491814 549264
rect 494610 549208 494666 549264
rect 483018 545420 483074 545456
rect 483018 545400 483020 545420
rect 483020 545400 483072 545420
rect 483072 545400 483074 545420
rect 485870 545128 485926 545184
rect 553306 545536 553362 545592
rect 553490 545536 553546 545592
rect 540978 545420 541034 545456
rect 540978 545400 540980 545420
rect 540980 545400 541032 545420
rect 541032 545400 541034 545420
rect 548614 545128 548670 545184
rect 560298 545556 560354 545592
rect 560298 545536 560300 545556
rect 560300 545536 560352 545556
rect 560352 545536 560354 545556
rect 579526 545536 579582 545592
rect 572626 545436 572628 545456
rect 572628 545436 572680 545456
rect 572680 545436 572682 545456
rect 572626 545400 572682 545436
rect 563150 545264 563206 545320
rect 559194 540368 559250 540424
rect 580354 627680 580410 627736
rect 580446 604152 580502 604208
rect 580630 592456 580686 592512
rect 580722 580760 580778 580816
rect 580630 540232 580686 540288
rect 580262 498616 580318 498672
rect 580906 533840 580962 533896
rect 580814 510312 580870 510368
rect 580538 486784 580594 486840
rect 580262 463392 580318 463448
rect 367098 413888 367154 413944
rect 368478 413888 368534 413944
rect 369858 413888 369914 413944
rect 371238 413888 371294 413944
rect 372618 413888 372674 413944
rect 373998 413888 374054 413944
rect 375378 413888 375434 413944
rect 376758 413888 376814 413944
rect 378138 413888 378194 413944
rect 379518 413888 379574 413944
rect 380898 413888 380954 413944
rect 382278 413888 382334 413944
rect 374090 413752 374146 413808
rect 368294 413344 368350 413400
rect 368754 413344 368810 413400
rect 382370 413752 382426 413808
rect 369766 413344 369822 413400
rect 369858 413208 369914 413264
rect 378046 413344 378102 413400
rect 379610 413208 379666 413264
rect 371974 413072 372030 413128
rect 372986 413072 373042 413128
rect 378782 413072 378838 413128
rect 381542 413072 381598 413128
rect 382278 413108 382280 413128
rect 382280 413108 382332 413128
rect 382332 413108 382334 413128
rect 382278 413072 382334 413108
rect 374366 412972 374368 412992
rect 374368 412972 374420 412992
rect 374420 412972 374422 412992
rect 374366 412936 374422 412972
rect 385038 413888 385094 413944
rect 383842 413752 383898 413808
rect 383566 412936 383622 412992
rect 386418 413244 386420 413264
rect 386420 413244 386472 413264
rect 386472 413244 386474 413264
rect 386418 413208 386474 413244
rect 388350 413344 388406 413400
rect 387338 413072 387394 413128
rect 384946 412972 384948 412992
rect 384948 412972 385000 412992
rect 385000 412972 385002 412992
rect 384946 412936 385002 412972
rect 386050 412956 386106 412992
rect 412638 413752 412694 413808
rect 396078 413616 396134 413672
rect 397458 413616 397514 413672
rect 405738 413516 405740 413536
rect 405740 413516 405792 413536
rect 405792 413516 405794 413536
rect 405738 413480 405794 413516
rect 386050 412936 386052 412956
rect 386052 412936 386104 412956
rect 386104 412936 386106 412956
rect 375470 412800 375526 412856
rect 376574 412800 376630 412856
rect 393318 412836 393320 412856
rect 393320 412836 393372 412856
rect 393372 412836 393374 412856
rect 393318 412800 393374 412836
rect 404358 413344 404414 413400
rect 401598 413208 401654 413264
rect 403162 413244 403164 413264
rect 403164 413244 403216 413264
rect 403216 413244 403218 413264
rect 403162 413208 403218 413244
rect 407118 413208 407174 413264
rect 398838 413108 398840 413128
rect 398840 413108 398892 413128
rect 398892 413108 398894 413128
rect 398838 413072 398894 413108
rect 408498 413072 408554 413128
rect 400218 412936 400274 412992
rect 397458 412800 397514 412856
rect 389638 412664 389694 412720
rect 390926 412664 390982 412720
rect 391754 412664 391810 412720
rect 393134 412664 393190 412720
rect 393962 412664 394018 412720
rect 394698 412664 394754 412720
rect 395342 412664 395398 412720
rect 396078 412700 396080 412720
rect 396080 412700 396132 412720
rect 396132 412700 396134 412720
rect 396078 412664 396134 412700
rect 405738 412684 405794 412720
rect 405738 412664 405740 412684
rect 405740 412664 405792 412684
rect 405792 412664 405794 412684
rect 388074 411748 388076 411768
rect 388076 411748 388128 411768
rect 388128 411748 388130 411768
rect 388074 411712 388130 411748
rect 391018 411576 391074 411632
rect 397458 411576 397514 411632
rect 399114 411612 399116 411632
rect 399116 411612 399168 411632
rect 399168 411612 399170 411632
rect 399114 411576 399170 411612
rect 389270 411440 389326 411496
rect 398010 411440 398066 411496
rect 400954 411476 400956 411496
rect 400956 411476 401008 411496
rect 401008 411476 401010 411496
rect 400954 411440 401010 411476
rect 403254 411440 403310 411496
rect 401690 411304 401746 411360
rect 404358 411340 404360 411360
rect 404360 411340 404412 411360
rect 404412 411340 404414 411360
rect 404358 411304 404414 411340
rect 389730 411032 389786 411088
rect 392306 410352 392362 410408
rect 409970 410352 410026 410408
rect 419538 392944 419594 393000
rect 419538 390632 419594 390688
rect 416410 323992 416466 324048
rect 337750 321952 337806 322008
rect 282826 320728 282882 320784
rect 61382 317328 61438 317384
rect 61014 3324 61070 3360
rect 61014 3304 61016 3324
rect 61016 3304 61068 3324
rect 61068 3304 61070 3324
rect 62118 3340 62120 3360
rect 62120 3340 62172 3360
rect 62172 3340 62174 3360
rect 62118 3304 62174 3340
rect 66258 227840 66314 227896
rect 66258 169904 66314 169960
rect 69386 216824 69442 216880
rect 69386 180920 69442 180976
rect 71778 4140 71834 4176
rect 74262 278704 74318 278760
rect 74446 278704 74502 278760
rect 74262 259392 74318 259448
rect 74446 259392 74502 259448
rect 74262 240080 74318 240136
rect 74446 240080 74502 240136
rect 74262 220768 74318 220824
rect 74446 220768 74502 220824
rect 74262 211112 74318 211168
rect 74446 211112 74502 211168
rect 74262 172488 74318 172544
rect 74446 172488 74502 172544
rect 74262 153176 74318 153232
rect 74446 153176 74502 153232
rect 74446 125568 74502 125624
rect 74446 124072 74502 124128
rect 71778 4120 71780 4140
rect 71780 4120 71832 4140
rect 71832 4120 71834 4140
rect 73066 4140 73122 4176
rect 73066 4120 73068 4140
rect 73068 4120 73120 4140
rect 73120 4120 73122 4140
rect 75826 227996 75882 228032
rect 75826 227976 75828 227996
rect 75828 227976 75880 227996
rect 75880 227976 75882 227996
rect 77206 216980 77262 217016
rect 77206 216960 77208 216980
rect 77208 216960 77260 216980
rect 77260 216960 77262 216980
rect 77206 181076 77262 181112
rect 77206 181056 77208 181076
rect 77208 181056 77260 181076
rect 77260 181056 77262 181076
rect 75826 170060 75882 170096
rect 75826 170040 75828 170060
rect 75828 170040 75880 170060
rect 75880 170040 75882 170060
rect 74630 125568 74686 125624
rect 74722 124072 74778 124128
rect 77206 76200 77262 76256
rect 77206 76064 77262 76120
rect 78862 4836 78864 4856
rect 78864 4836 78916 4856
rect 78916 4836 78918 4856
rect 78862 4800 78918 4836
rect 75458 3712 75514 3768
rect 77850 3984 77906 4040
rect 80058 4020 80060 4040
rect 80060 4020 80112 4040
rect 80112 4020 80114 4040
rect 80058 3984 80114 4020
rect 81990 5092 82046 5128
rect 81990 5072 81992 5092
rect 81992 5072 82044 5092
rect 82044 5072 82046 5092
rect 81990 4956 82046 4992
rect 81990 4936 81992 4956
rect 81992 4936 82044 4956
rect 82044 4936 82046 4956
rect 89534 216860 89536 216880
rect 89536 216860 89588 216880
rect 89588 216860 89590 216880
rect 89534 216824 89590 216860
rect 89534 170040 89590 170096
rect 89534 169768 89590 169824
rect 89258 144880 89314 144936
rect 89442 144880 89498 144936
rect 89626 76100 89628 76120
rect 89628 76100 89680 76120
rect 89680 76100 89682 76120
rect 89626 76064 89682 76100
rect 89534 31728 89590 31784
rect 89258 26288 89314 26344
rect 86038 4140 86094 4176
rect 86038 4120 86040 4140
rect 86040 4120 86092 4140
rect 86092 4120 86094 4140
rect 86866 5092 86922 5128
rect 86866 5072 86868 5092
rect 86868 5072 86920 5092
rect 86920 5072 86922 5092
rect 86774 4956 86830 4992
rect 86774 4936 86776 4956
rect 86776 4936 86828 4956
rect 86828 4936 86830 4956
rect 86866 4836 86868 4856
rect 86868 4836 86920 4856
rect 86920 4836 86922 4856
rect 86866 4800 86922 4836
rect 89534 4120 89590 4176
rect 91742 216860 91744 216880
rect 91744 216860 91796 216880
rect 91796 216860 91798 216880
rect 91742 216824 91798 216860
rect 91742 76100 91744 76120
rect 91744 76100 91796 76120
rect 91796 76100 91798 76120
rect 91742 76064 91798 76100
rect 90914 5208 90970 5264
rect 89442 3848 89498 3904
rect 89902 3884 89904 3904
rect 89904 3884 89956 3904
rect 89956 3884 89958 3904
rect 89902 3848 89958 3884
rect 93214 3848 93270 3904
rect 92110 3576 92166 3632
rect 94502 5072 94558 5128
rect 93858 3884 93860 3904
rect 93860 3884 93912 3904
rect 93912 3884 93914 3904
rect 93858 3848 93914 3884
rect 95514 3868 95570 3904
rect 95514 3848 95516 3868
rect 95516 3848 95568 3868
rect 95568 3848 95570 3868
rect 96618 3848 96674 3904
rect 99286 3440 99342 3496
rect 101586 4936 101642 4992
rect 102598 3848 102654 3904
rect 103518 3868 103574 3904
rect 103518 3848 103520 3868
rect 103520 3848 103572 3868
rect 103572 3848 103574 3868
rect 103978 3304 104034 3360
rect 111062 264288 111118 264344
rect 111062 263608 111118 263664
rect 111062 228384 111118 228440
rect 111062 227704 111118 227760
rect 111062 181464 111118 181520
rect 111062 180784 111118 180840
rect 111062 170448 111118 170504
rect 111062 169768 111118 169824
rect 115846 318280 115902 318336
rect 115938 263644 115940 263664
rect 115940 263644 115992 263664
rect 115992 263644 115994 263664
rect 115938 263608 115994 263644
rect 115938 227740 115940 227760
rect 115940 227740 115992 227760
rect 115992 227740 115994 227760
rect 115938 227704 115994 227740
rect 115938 216724 115940 216744
rect 115940 216724 115992 216744
rect 115992 216724 115994 216744
rect 115938 216688 115994 216724
rect 115938 169804 115940 169824
rect 115940 169804 115992 169824
rect 115992 169804 115994 169824
rect 115938 169768 115994 169804
rect 115938 75964 115940 75984
rect 115940 75964 115992 75984
rect 115992 75964 115994 75984
rect 115938 75928 115994 75964
rect 118790 263880 118846 263936
rect 118790 227976 118846 228032
rect 118790 216960 118846 217016
rect 118790 170040 118846 170096
rect 118790 76200 118846 76256
rect 121366 318144 121422 318200
rect 122746 318008 122802 318064
rect 128266 180920 128322 180976
rect 128450 180920 128506 180976
rect 131394 4800 131450 4856
rect 135166 264152 135222 264208
rect 135166 263744 135222 263800
rect 135166 228248 135222 228304
rect 135166 227840 135222 227896
rect 135166 217232 135222 217288
rect 135166 216824 135222 216880
rect 135166 170312 135222 170368
rect 135166 169904 135222 169960
rect 135166 76472 135222 76528
rect 135166 76064 135222 76120
rect 140042 264016 140098 264072
rect 140042 263608 140098 263664
rect 140042 228112 140098 228168
rect 140042 227704 140098 227760
rect 140042 217096 140098 217152
rect 140042 216688 140098 216744
rect 140042 170176 140098 170232
rect 140042 169768 140098 169824
rect 140042 76336 140098 76392
rect 140042 75928 140098 75984
rect 147586 263780 147588 263800
rect 147588 263780 147640 263800
rect 147640 263780 147642 263800
rect 147586 263744 147642 263780
rect 147586 227876 147588 227896
rect 147588 227876 147640 227896
rect 147640 227876 147642 227896
rect 147586 227840 147642 227876
rect 147586 216860 147588 216880
rect 147588 216860 147640 216880
rect 147640 216860 147642 216880
rect 147586 216824 147642 216860
rect 147586 169940 147588 169960
rect 147588 169940 147640 169960
rect 147640 169940 147642 169960
rect 147586 169904 147642 169940
rect 147586 76100 147588 76120
rect 147588 76100 147640 76120
rect 147640 76100 147642 76120
rect 147586 76064 147642 76100
rect 154486 263880 154542 263936
rect 154486 227976 154542 228032
rect 154486 216960 154542 217016
rect 154486 170040 154542 170096
rect 154486 76200 154542 76256
rect 208398 5208 208454 5264
rect 183558 3712 183614 3768
rect 213918 5072 213974 5128
rect 209778 3576 209834 3632
rect 226338 4936 226394 4992
rect 222198 3440 222254 3496
rect 247774 318280 247830 318336
rect 257526 318144 257582 318200
rect 259458 318008 259514 318064
rect 274638 4800 274694 4856
rect 339774 320592 339830 320648
rect 349986 320592 350042 320648
rect 580170 346024 580226 346080
rect 419906 332560 419962 332616
rect 419814 328616 419870 328672
rect 419722 327120 419778 327176
rect 419630 325760 419686 325816
rect 339774 320320 339830 320376
rect 349986 320320 350042 320376
rect 420182 331200 420238 331256
rect 419998 329840 420054 329896
rect 579986 322632 580042 322688
rect 579986 320592 580042 320648
rect 580354 451696 580410 451752
rect 580262 320456 580318 320512
rect 580446 439864 580502 439920
rect 580538 416472 580594 416528
rect 580630 404776 580686 404832
rect 580538 320864 580594 320920
rect 580722 392944 580778 393000
rect 580814 369552 580870 369608
rect 580906 357856 580962 357912
rect 344006 318724 344008 318744
rect 344008 318724 344060 318744
rect 344060 318724 344062 318744
rect 344006 318688 344062 318724
rect 347778 318416 347834 318472
rect 580170 310800 580226 310856
rect 579802 299104 579858 299160
rect 580170 275712 580226 275768
rect 579802 252184 579858 252240
rect 579802 205264 579858 205320
rect 579802 158344 579858 158400
rect 580170 134816 580226 134872
rect 580170 123120 580226 123176
rect 579802 111424 579858 111480
rect 580170 87896 580226 87952
rect 579802 64504 579858 64560
rect 580170 40976 580226 41032
rect 580170 29280 580226 29336
rect 579802 17584 579858 17640
rect 229098 3304 229154 3360
<< metal3 >>
rect 57830 700300 57836 700364
rect 57900 700362 57906 700364
rect 543457 700362 543523 700365
rect 57900 700360 543523 700362
rect 57900 700304 543462 700360
rect 543518 700304 543523 700360
rect 57900 700302 543523 700304
rect 57900 700300 57906 700302
rect 543457 700299 543523 700302
rect 583520 698050 584960 698140
rect 583342 697990 584960 698050
rect 550582 697308 550588 697372
rect 550652 697370 550658 697372
rect 553301 697370 553367 697373
rect 550652 697368 553367 697370
rect 550652 697312 553306 697368
rect 553362 697312 553367 697368
rect 550652 697310 553367 697312
rect 550652 697308 550658 697310
rect 553301 697307 553367 697310
rect 553485 697370 553551 697373
rect 560293 697370 560359 697373
rect 553485 697368 560359 697370
rect 553485 697312 553490 697368
rect 553546 697312 560298 697368
rect 560354 697312 560359 697368
rect 553485 697310 560359 697312
rect 553485 697307 553551 697310
rect 560293 697307 560359 697310
rect 59118 697172 59124 697236
rect 59188 697234 59194 697236
rect 77201 697234 77267 697237
rect 96521 697234 96587 697237
rect 115841 697234 115907 697237
rect 135161 697234 135227 697237
rect 154481 697234 154547 697237
rect 173801 697234 173867 697237
rect 193121 697234 193187 697237
rect 212441 697234 212507 697237
rect 231761 697234 231827 697237
rect 251081 697234 251147 697237
rect 270401 697234 270467 697237
rect 289721 697234 289787 697237
rect 309041 697234 309107 697237
rect 328361 697234 328427 697237
rect 540973 697234 541039 697237
rect 59188 697174 60842 697234
rect 59188 697172 59194 697174
rect 60782 697098 60842 697174
rect 77201 697232 80162 697234
rect 77201 697176 77206 697232
rect 77262 697176 80162 697232
rect 77201 697174 80162 697176
rect 77201 697171 77267 697174
rect 70301 697098 70367 697101
rect 60782 697096 70367 697098
rect 60782 697040 70306 697096
rect 70362 697040 70367 697096
rect 60782 697038 70367 697040
rect 80102 697098 80162 697174
rect 96521 697232 99482 697234
rect 96521 697176 96526 697232
rect 96582 697176 99482 697232
rect 96521 697174 99482 697176
rect 96521 697171 96587 697174
rect 89621 697098 89687 697101
rect 80102 697096 89687 697098
rect 80102 697040 89626 697096
rect 89682 697040 89687 697096
rect 80102 697038 89687 697040
rect 99422 697098 99482 697174
rect 115841 697232 118802 697234
rect 115841 697176 115846 697232
rect 115902 697176 118802 697232
rect 115841 697174 118802 697176
rect 115841 697171 115907 697174
rect 108941 697098 109007 697101
rect 99422 697096 109007 697098
rect 99422 697040 108946 697096
rect 109002 697040 109007 697096
rect 99422 697038 109007 697040
rect 118742 697098 118802 697174
rect 135161 697232 138122 697234
rect 135161 697176 135166 697232
rect 135222 697176 138122 697232
rect 135161 697174 138122 697176
rect 135161 697171 135227 697174
rect 128261 697098 128327 697101
rect 118742 697096 128327 697098
rect 118742 697040 128266 697096
rect 128322 697040 128327 697096
rect 118742 697038 128327 697040
rect 138062 697098 138122 697174
rect 154481 697232 157442 697234
rect 154481 697176 154486 697232
rect 154542 697176 157442 697232
rect 154481 697174 157442 697176
rect 154481 697171 154547 697174
rect 147581 697098 147647 697101
rect 138062 697096 147647 697098
rect 138062 697040 147586 697096
rect 147642 697040 147647 697096
rect 138062 697038 147647 697040
rect 157382 697098 157442 697174
rect 173801 697232 176762 697234
rect 173801 697176 173806 697232
rect 173862 697176 176762 697232
rect 173801 697174 176762 697176
rect 173801 697171 173867 697174
rect 166901 697098 166967 697101
rect 157382 697096 166967 697098
rect 157382 697040 166906 697096
rect 166962 697040 166967 697096
rect 157382 697038 166967 697040
rect 176702 697098 176762 697174
rect 193121 697232 196082 697234
rect 193121 697176 193126 697232
rect 193182 697176 196082 697232
rect 193121 697174 196082 697176
rect 193121 697171 193187 697174
rect 186221 697098 186287 697101
rect 176702 697096 186287 697098
rect 176702 697040 186226 697096
rect 186282 697040 186287 697096
rect 176702 697038 186287 697040
rect 196022 697098 196082 697174
rect 212441 697232 215402 697234
rect 212441 697176 212446 697232
rect 212502 697176 215402 697232
rect 212441 697174 215402 697176
rect 212441 697171 212507 697174
rect 205541 697098 205607 697101
rect 196022 697096 205607 697098
rect 196022 697040 205546 697096
rect 205602 697040 205607 697096
rect 196022 697038 205607 697040
rect 215342 697098 215402 697174
rect 231761 697232 234722 697234
rect 231761 697176 231766 697232
rect 231822 697176 234722 697232
rect 231761 697174 234722 697176
rect 231761 697171 231827 697174
rect 224861 697098 224927 697101
rect 215342 697096 224927 697098
rect 215342 697040 224866 697096
rect 224922 697040 224927 697096
rect 215342 697038 224927 697040
rect 234662 697098 234722 697174
rect 251081 697232 254042 697234
rect 251081 697176 251086 697232
rect 251142 697176 254042 697232
rect 251081 697174 254042 697176
rect 251081 697171 251147 697174
rect 244181 697098 244247 697101
rect 234662 697096 244247 697098
rect 234662 697040 244186 697096
rect 244242 697040 244247 697096
rect 234662 697038 244247 697040
rect 253982 697098 254042 697174
rect 270401 697232 273362 697234
rect 270401 697176 270406 697232
rect 270462 697176 273362 697232
rect 270401 697174 273362 697176
rect 270401 697171 270467 697174
rect 263501 697098 263567 697101
rect 253982 697096 263567 697098
rect 253982 697040 263506 697096
rect 263562 697040 263567 697096
rect 253982 697038 263567 697040
rect 273302 697098 273362 697174
rect 289721 697232 292682 697234
rect 289721 697176 289726 697232
rect 289782 697176 292682 697232
rect 289721 697174 292682 697176
rect 289721 697171 289787 697174
rect 282821 697098 282887 697101
rect 273302 697096 282887 697098
rect 273302 697040 282826 697096
rect 282882 697040 282887 697096
rect 273302 697038 282887 697040
rect 292622 697098 292682 697174
rect 309041 697232 312002 697234
rect 309041 697176 309046 697232
rect 309102 697176 312002 697232
rect 309041 697174 312002 697176
rect 309041 697171 309107 697174
rect 302141 697098 302207 697101
rect 292622 697096 302207 697098
rect 292622 697040 302146 697096
rect 302202 697040 302207 697096
rect 292622 697038 302207 697040
rect 311942 697098 312002 697174
rect 328361 697232 340890 697234
rect 328361 697176 328366 697232
rect 328422 697176 340890 697232
rect 328361 697174 340890 697176
rect 328361 697171 328427 697174
rect 321461 697098 321527 697101
rect 311942 697096 321527 697098
rect 311942 697040 321466 697096
rect 321522 697040 321527 697096
rect 311942 697038 321527 697040
rect 340830 697098 340890 697174
rect 373950 697174 383578 697234
rect 340830 697038 350458 697098
rect 70301 697035 70367 697038
rect 89621 697035 89687 697038
rect 108941 697035 109007 697038
rect 128261 697035 128327 697038
rect 147581 697035 147647 697038
rect 166901 697035 166967 697038
rect 186221 697035 186287 697038
rect 205541 697035 205607 697038
rect 224861 697035 224927 697038
rect 244181 697035 244247 697038
rect 263501 697035 263567 697038
rect 282821 697035 282887 697038
rect 302141 697035 302207 697038
rect 321461 697035 321527 697038
rect 350398 696962 350458 697038
rect 373950 696962 374010 697174
rect 350398 696902 374010 696962
rect 383518 696962 383578 697174
rect 383702 697174 393330 697234
rect 383702 696962 383762 697174
rect 393270 697098 393330 697174
rect 403022 697174 412650 697234
rect 393270 697038 402898 697098
rect 383518 696902 383762 696962
rect 402838 696962 402898 697038
rect 403022 696962 403082 697174
rect 412590 697098 412650 697174
rect 422342 697174 431970 697234
rect 412590 697038 422218 697098
rect 402838 696902 403082 696962
rect 422158 696962 422218 697038
rect 422342 696962 422402 697174
rect 431910 697098 431970 697174
rect 441662 697174 451290 697234
rect 431910 697038 441538 697098
rect 422158 696902 422402 696962
rect 441478 696962 441538 697038
rect 441662 696962 441722 697174
rect 451230 697098 451290 697174
rect 460982 697174 470610 697234
rect 451230 697038 460858 697098
rect 441478 696902 441722 696962
rect 460798 696962 460858 697038
rect 460982 696962 461042 697174
rect 470550 697098 470610 697174
rect 480302 697174 489930 697234
rect 470550 697038 480178 697098
rect 460798 696902 461042 696962
rect 480118 696962 480178 697038
rect 480302 696962 480362 697174
rect 489870 697098 489930 697174
rect 499622 697174 509250 697234
rect 489870 697038 499498 697098
rect 480118 696902 480362 696962
rect 499438 696962 499498 697038
rect 499622 696962 499682 697174
rect 509190 697098 509250 697174
rect 518942 697174 528570 697234
rect 509190 697038 518818 697098
rect 499438 696902 499682 696962
rect 518758 696962 518818 697038
rect 518942 696962 519002 697174
rect 528510 697098 528570 697174
rect 538262 697232 541039 697234
rect 538262 697176 540978 697232
rect 541034 697176 541039 697232
rect 538262 697174 541039 697176
rect 528510 697038 538138 697098
rect 518758 696902 519002 696962
rect 538078 696962 538138 697038
rect 538262 696962 538322 697174
rect 540973 697171 541039 697174
rect 565169 697234 565235 697237
rect 572713 697234 572779 697237
rect 565169 697232 569970 697234
rect 565169 697176 565174 697232
rect 565230 697176 569970 697232
rect 565169 697174 569970 697176
rect 565169 697171 565235 697174
rect 569910 697098 569970 697174
rect 572713 697232 576962 697234
rect 572713 697176 572718 697232
rect 572774 697176 576962 697232
rect 572713 697174 576962 697176
rect 572713 697171 572779 697174
rect 572621 697098 572687 697101
rect 569910 697096 572687 697098
rect 569910 697040 572626 697096
rect 572682 697040 572687 697096
rect 569910 697038 572687 697040
rect 576902 697098 576962 697174
rect 583342 697098 583402 697990
rect 583520 697900 584960 697990
rect 576902 697038 583402 697098
rect 572621 697035 572687 697038
rect 538078 696902 538322 696962
rect 548609 696962 548675 696965
rect 550582 696962 550588 696964
rect 548609 696960 550588 696962
rect 548609 696904 548614 696960
rect 548670 696904 550588 696960
rect 548609 696902 550588 696904
rect 548609 696899 548675 696902
rect 550582 696900 550588 696902
rect 550652 696900 550658 696964
rect -960 696540 480 696780
rect 183502 686428 183508 686492
rect 183572 686490 183578 686492
rect 188337 686490 188403 686493
rect 183572 686488 188403 686490
rect 183572 686432 188342 686488
rect 188398 686432 188403 686488
rect 183572 686430 188403 686432
rect 183572 686428 183578 686430
rect 188337 686427 188403 686430
rect 376702 686428 376708 686492
rect 376772 686490 376778 686492
rect 379513 686490 379579 686493
rect 376772 686488 379579 686490
rect 376772 686432 379518 686488
rect 379574 686432 379579 686488
rect 376772 686430 379579 686432
rect 376772 686428 376778 686430
rect 379513 686427 379579 686430
rect 434662 686428 434668 686492
rect 434732 686490 434738 686492
rect 441521 686490 441587 686493
rect 434732 686488 441587 686490
rect 434732 686432 441526 686488
rect 441582 686432 441587 686488
rect 434732 686430 441587 686432
rect 434732 686428 434738 686430
rect 441521 686427 441587 686430
rect 164182 686292 164188 686356
rect 164252 686354 164258 686356
rect 166901 686354 166967 686357
rect 164252 686352 166967 686354
rect 164252 686296 166906 686352
rect 166962 686296 166967 686352
rect 164252 686294 166967 686296
rect 164252 686292 164258 686294
rect 166901 686291 166967 686294
rect 167085 686354 167151 686357
rect 173893 686354 173959 686357
rect 167085 686352 173959 686354
rect 167085 686296 167090 686352
rect 167146 686296 173898 686352
rect 173954 686296 173959 686352
rect 167085 686294 173959 686296
rect 167085 686291 167151 686294
rect 173893 686291 173959 686294
rect 357382 686292 357388 686356
rect 357452 686354 357458 686356
rect 360101 686354 360167 686357
rect 357452 686352 360167 686354
rect 357452 686296 360106 686352
rect 360162 686296 360167 686352
rect 357452 686294 360167 686296
rect 357452 686292 357458 686294
rect 360101 686291 360167 686294
rect 360285 686354 360351 686357
rect 367093 686354 367159 686357
rect 360285 686352 367159 686354
rect 360285 686296 360290 686352
rect 360346 686296 367098 686352
rect 367154 686296 367159 686352
rect 360285 686294 367159 686296
rect 360285 686291 360351 686294
rect 367093 686291 367159 686294
rect 550582 686292 550588 686356
rect 550652 686354 550658 686356
rect 553301 686354 553367 686357
rect 550652 686352 553367 686354
rect 550652 686296 553306 686352
rect 553362 686296 553367 686352
rect 550652 686294 553367 686296
rect 550652 686292 550658 686294
rect 553301 686291 553367 686294
rect 553485 686354 553551 686357
rect 560293 686354 560359 686357
rect 583520 686354 584960 686444
rect 553485 686352 560359 686354
rect 553485 686296 553490 686352
rect 553546 686296 560298 686352
rect 560354 686296 560359 686352
rect 553485 686294 560359 686296
rect 553485 686291 553551 686294
rect 560293 686291 560359 686294
rect 583342 686294 584960 686354
rect 57646 686156 57652 686220
rect 57716 686218 57722 686220
rect 154573 686218 154639 686221
rect 57716 686158 64890 686218
rect 57716 686156 57722 686158
rect 64830 686082 64890 686158
rect 74582 686158 84210 686218
rect 64830 686022 74458 686082
rect 74398 685946 74458 686022
rect 74582 685946 74642 686158
rect 84150 686082 84210 686158
rect 93902 686158 103530 686218
rect 84150 686022 93778 686082
rect 74398 685886 74642 685946
rect 93718 685946 93778 686022
rect 93902 685946 93962 686158
rect 103470 686082 103530 686158
rect 113222 686158 122850 686218
rect 103470 686022 113098 686082
rect 93718 685886 93962 685946
rect 113038 685946 113098 686022
rect 113222 685946 113282 686158
rect 122790 686082 122850 686158
rect 132542 686158 142170 686218
rect 122790 686022 132418 686082
rect 113038 685886 113282 685946
rect 132358 685946 132418 686022
rect 132542 685946 132602 686158
rect 142110 686082 142170 686158
rect 151862 686216 154639 686218
rect 151862 686160 154578 686216
rect 154634 686160 154639 686216
rect 151862 686158 154639 686160
rect 142110 686022 151738 686082
rect 132358 685886 132602 685946
rect 151678 685946 151738 686022
rect 151862 685946 151922 686158
rect 154573 686155 154639 686158
rect 178769 686218 178835 686221
rect 183502 686218 183508 686220
rect 178769 686216 183508 686218
rect 178769 686160 178774 686216
rect 178830 686160 183508 686216
rect 178769 686158 183508 686160
rect 178769 686155 178835 686158
rect 183502 686156 183508 686158
rect 183572 686156 183578 686220
rect 188337 686218 188403 686221
rect 289813 686218 289879 686221
rect 188337 686216 200130 686218
rect 188337 686160 188342 686216
rect 188398 686160 200130 686216
rect 188337 686158 200130 686160
rect 188337 686155 188403 686158
rect 200070 686082 200130 686158
rect 209822 686158 219450 686218
rect 200070 686022 209698 686082
rect 151678 685886 151922 685946
rect 162209 685946 162275 685949
rect 164182 685946 164188 685948
rect 162209 685944 164188 685946
rect 162209 685888 162214 685944
rect 162270 685888 164188 685944
rect 162209 685886 164188 685888
rect 162209 685883 162275 685886
rect 164182 685884 164188 685886
rect 164252 685884 164258 685948
rect 209638 685946 209698 686022
rect 209822 685946 209882 686158
rect 219390 686082 219450 686158
rect 229142 686158 238770 686218
rect 219390 686022 229018 686082
rect 209638 685886 209882 685946
rect 228958 685946 229018 686022
rect 229142 685946 229202 686158
rect 238710 686082 238770 686158
rect 248462 686158 258090 686218
rect 238710 686022 248338 686082
rect 228958 685886 229202 685946
rect 248278 685946 248338 686022
rect 248462 685946 248522 686158
rect 258030 686082 258090 686158
rect 267782 686158 277410 686218
rect 258030 686022 267658 686082
rect 248278 685886 248522 685946
rect 267598 685946 267658 686022
rect 267782 685946 267842 686158
rect 277350 686082 277410 686158
rect 287102 686216 289879 686218
rect 287102 686160 289818 686216
rect 289874 686160 289879 686216
rect 287102 686158 289879 686160
rect 277350 686022 286978 686082
rect 267598 685886 267842 685946
rect 286918 685946 286978 686022
rect 287102 685946 287162 686158
rect 289813 686155 289879 686158
rect 299422 686156 299428 686220
rect 299492 686218 299498 686220
rect 347773 686218 347839 686221
rect 299492 686158 316050 686218
rect 299492 686156 299498 686158
rect 315990 686082 316050 686158
rect 325742 686158 335370 686218
rect 315990 686022 325618 686082
rect 286918 685886 287162 685946
rect 294505 685946 294571 685949
rect 299422 685946 299428 685948
rect 294505 685944 299428 685946
rect 294505 685888 294510 685944
rect 294566 685888 299428 685944
rect 294505 685886 299428 685888
rect 294505 685883 294571 685886
rect 299422 685884 299428 685886
rect 299492 685884 299498 685948
rect 325558 685946 325618 686022
rect 325742 685946 325802 686158
rect 335310 686082 335370 686158
rect 345062 686216 347839 686218
rect 345062 686160 347778 686216
rect 347834 686160 347839 686216
rect 345062 686158 347839 686160
rect 335310 686022 344938 686082
rect 325558 685886 325802 685946
rect 344878 685946 344938 686022
rect 345062 685946 345122 686158
rect 347773 686155 347839 686158
rect 371969 686218 372035 686221
rect 376702 686218 376708 686220
rect 371969 686216 376708 686218
rect 371969 686160 371974 686216
rect 372030 686160 376708 686216
rect 371969 686158 376708 686160
rect 371969 686155 372035 686158
rect 376702 686156 376708 686158
rect 376772 686156 376778 686220
rect 379513 686218 379579 686221
rect 427537 686218 427603 686221
rect 379513 686216 393330 686218
rect 379513 686160 379518 686216
rect 379574 686160 393330 686216
rect 379513 686158 393330 686160
rect 379513 686155 379579 686158
rect 393270 686082 393330 686158
rect 403022 686216 427603 686218
rect 403022 686160 427542 686216
rect 427598 686160 427603 686216
rect 403022 686158 427603 686160
rect 393270 686022 402898 686082
rect 344878 685886 345122 685946
rect 355409 685946 355475 685949
rect 357382 685946 357388 685948
rect 355409 685944 357388 685946
rect 355409 685888 355414 685944
rect 355470 685888 357388 685944
rect 355409 685886 357388 685888
rect 355409 685883 355475 685886
rect 357382 685884 357388 685886
rect 357452 685884 357458 685948
rect 402838 685946 402898 686022
rect 403022 685946 403082 686158
rect 427537 686155 427603 686158
rect 427721 686218 427787 686221
rect 441521 686218 441587 686221
rect 540973 686218 541039 686221
rect 427721 686216 429762 686218
rect 427721 686160 427726 686216
rect 427782 686160 429762 686216
rect 427721 686158 429762 686160
rect 427721 686155 427787 686158
rect 429702 686082 429762 686158
rect 441521 686216 451290 686218
rect 441521 686160 441526 686216
rect 441582 686160 451290 686216
rect 441521 686158 451290 686160
rect 441521 686155 441587 686158
rect 434662 686082 434668 686084
rect 429702 686022 434668 686082
rect 434662 686020 434668 686022
rect 434732 686020 434738 686084
rect 451230 686082 451290 686158
rect 460982 686158 470610 686218
rect 451230 686022 460858 686082
rect 402838 685886 403082 685946
rect 460798 685946 460858 686022
rect 460982 685946 461042 686158
rect 470550 686082 470610 686158
rect 480302 686158 489930 686218
rect 470550 686022 480178 686082
rect 460798 685886 461042 685946
rect 480118 685946 480178 686022
rect 480302 685946 480362 686158
rect 489870 686082 489930 686158
rect 499622 686158 509250 686218
rect 489870 686022 499498 686082
rect 480118 685886 480362 685946
rect 499438 685946 499498 686022
rect 499622 685946 499682 686158
rect 509190 686082 509250 686158
rect 518942 686158 528570 686218
rect 509190 686022 518818 686082
rect 499438 685886 499682 685946
rect 518758 685946 518818 686022
rect 518942 685946 519002 686158
rect 528510 686082 528570 686158
rect 538262 686216 541039 686218
rect 538262 686160 540978 686216
rect 541034 686160 541039 686216
rect 538262 686158 541039 686160
rect 528510 686022 538138 686082
rect 518758 685886 519002 685946
rect 538078 685946 538138 686022
rect 538262 685946 538322 686158
rect 540973 686155 541039 686158
rect 565169 686218 565235 686221
rect 572713 686218 572779 686221
rect 565169 686216 569970 686218
rect 565169 686160 565174 686216
rect 565230 686160 569970 686216
rect 565169 686158 569970 686160
rect 565169 686155 565235 686158
rect 569910 686082 569970 686158
rect 572713 686216 576962 686218
rect 572713 686160 572718 686216
rect 572774 686160 576962 686216
rect 572713 686158 576962 686160
rect 572713 686155 572779 686158
rect 572621 686082 572687 686085
rect 569910 686080 572687 686082
rect 569910 686024 572626 686080
rect 572682 686024 572687 686080
rect 569910 686022 572687 686024
rect 576902 686082 576962 686158
rect 583342 686082 583402 686294
rect 583520 686204 584960 686294
rect 576902 686022 583402 686082
rect 572621 686019 572687 686022
rect 538078 685886 538322 685946
rect 548609 685946 548675 685949
rect 550582 685946 550588 685948
rect 548609 685944 550588 685946
rect 548609 685888 548614 685944
rect 548670 685888 550588 685944
rect 548609 685886 550588 685888
rect 548609 685883 548675 685886
rect 550582 685884 550588 685886
rect 550652 685884 550658 685948
rect 559005 684448 559071 684453
rect 559005 684392 559010 684448
rect 559066 684392 559071 684448
rect 559005 684387 559071 684392
rect 559008 684317 559068 684387
rect 559005 684312 559071 684317
rect 559005 684256 559010 684312
rect 559066 684256 559071 684312
rect 559005 684251 559071 684256
rect -960 682274 480 682364
rect 3417 682274 3483 682277
rect -960 682272 3483 682274
rect -960 682216 3422 682272
rect 3478 682216 3483 682272
rect -960 682214 3483 682216
rect -960 682124 480 682214
rect 3417 682211 3483 682214
rect 583520 674658 584960 674748
rect 583342 674598 584960 674658
rect 183502 674052 183508 674116
rect 183572 674114 183578 674116
rect 188337 674114 188403 674117
rect 183572 674112 188403 674114
rect 183572 674056 188342 674112
rect 188398 674056 188403 674112
rect 183572 674054 188403 674056
rect 183572 674052 183578 674054
rect 188337 674051 188403 674054
rect 376702 674052 376708 674116
rect 376772 674114 376778 674116
rect 379513 674114 379579 674117
rect 376772 674112 379579 674114
rect 376772 674056 379518 674112
rect 379574 674056 379579 674112
rect 376772 674054 379579 674056
rect 376772 674052 376778 674054
rect 379513 674051 379579 674054
rect 166993 673978 167059 673981
rect 173893 673978 173959 673981
rect 166993 673976 173959 673978
rect 166993 673920 166998 673976
rect 167054 673920 173898 673976
rect 173954 673920 173959 673976
rect 166993 673918 173959 673920
rect 166993 673915 167059 673918
rect 173893 673915 173959 673918
rect 357382 673916 357388 673980
rect 357452 673978 357458 673980
rect 360101 673978 360167 673981
rect 357452 673976 360167 673978
rect 357452 673920 360106 673976
rect 360162 673920 360167 673976
rect 357452 673918 360167 673920
rect 357452 673916 357458 673918
rect 360101 673915 360167 673918
rect 360285 673978 360351 673981
rect 367093 673978 367159 673981
rect 360285 673976 367159 673978
rect 360285 673920 360290 673976
rect 360346 673920 367098 673976
rect 367154 673920 367159 673976
rect 360285 673918 367159 673920
rect 360285 673915 360351 673918
rect 367093 673915 367159 673918
rect 553393 673978 553459 673981
rect 560293 673978 560359 673981
rect 553393 673976 560359 673978
rect 553393 673920 553398 673976
rect 553454 673920 560298 673976
rect 560354 673920 560359 673976
rect 553393 673918 560359 673920
rect 553393 673915 553459 673918
rect 560293 673915 560359 673918
rect 59302 673780 59308 673844
rect 59372 673842 59378 673844
rect 154573 673842 154639 673845
rect 59372 673782 64890 673842
rect 59372 673780 59378 673782
rect 64830 673706 64890 673782
rect 74582 673782 84210 673842
rect 64830 673646 74458 673706
rect 74398 673570 74458 673646
rect 74582 673570 74642 673782
rect 84150 673706 84210 673782
rect 93902 673782 103530 673842
rect 84150 673646 93778 673706
rect 74398 673510 74642 673570
rect 93718 673570 93778 673646
rect 93902 673570 93962 673782
rect 103470 673706 103530 673782
rect 113222 673782 122850 673842
rect 103470 673646 113098 673706
rect 93718 673510 93962 673570
rect 113038 673570 113098 673646
rect 113222 673570 113282 673782
rect 122790 673706 122850 673782
rect 132542 673782 142170 673842
rect 122790 673646 132418 673706
rect 113038 673510 113282 673570
rect 132358 673570 132418 673646
rect 132542 673570 132602 673782
rect 142110 673706 142170 673782
rect 151862 673840 154639 673842
rect 151862 673784 154578 673840
rect 154634 673784 154639 673840
rect 151862 673782 154639 673784
rect 142110 673646 151738 673706
rect 132358 673510 132602 673570
rect 151678 673570 151738 673646
rect 151862 673570 151922 673782
rect 154573 673779 154639 673782
rect 178769 673842 178835 673845
rect 183502 673842 183508 673844
rect 178769 673840 183508 673842
rect 178769 673784 178774 673840
rect 178830 673784 183508 673840
rect 178769 673782 183508 673784
rect 178769 673779 178835 673782
rect 183502 673780 183508 673782
rect 183572 673780 183578 673844
rect 188337 673842 188403 673845
rect 289813 673842 289879 673845
rect 188337 673840 200130 673842
rect 188337 673784 188342 673840
rect 188398 673784 200130 673840
rect 188337 673782 200130 673784
rect 188337 673779 188403 673782
rect 200070 673706 200130 673782
rect 209822 673782 219450 673842
rect 200070 673646 209698 673706
rect 151678 673510 151922 673570
rect 162209 673570 162275 673573
rect 166901 673570 166967 673573
rect 162209 673568 166967 673570
rect 162209 673512 162214 673568
rect 162270 673512 166906 673568
rect 166962 673512 166967 673568
rect 162209 673510 166967 673512
rect 209638 673570 209698 673646
rect 209822 673570 209882 673782
rect 219390 673706 219450 673782
rect 229142 673782 238770 673842
rect 219390 673646 229018 673706
rect 209638 673510 209882 673570
rect 228958 673570 229018 673646
rect 229142 673570 229202 673782
rect 238710 673706 238770 673782
rect 248462 673782 258090 673842
rect 238710 673646 248338 673706
rect 228958 673510 229202 673570
rect 248278 673570 248338 673646
rect 248462 673570 248522 673782
rect 258030 673706 258090 673782
rect 267782 673782 277410 673842
rect 258030 673646 267658 673706
rect 248278 673510 248522 673570
rect 267598 673570 267658 673646
rect 267782 673570 267842 673782
rect 277350 673706 277410 673782
rect 287102 673840 289879 673842
rect 287102 673784 289818 673840
rect 289874 673784 289879 673840
rect 287102 673782 289879 673784
rect 277350 673646 286978 673706
rect 267598 673510 267842 673570
rect 286918 673570 286978 673646
rect 287102 673570 287162 673782
rect 289813 673779 289879 673782
rect 299422 673780 299428 673844
rect 299492 673842 299498 673844
rect 347773 673842 347839 673845
rect 299492 673782 316050 673842
rect 299492 673780 299498 673782
rect 315990 673706 316050 673782
rect 325742 673782 335370 673842
rect 315990 673646 325618 673706
rect 286918 673510 287162 673570
rect 292665 673570 292731 673573
rect 299422 673570 299428 673572
rect 292665 673568 299428 673570
rect 292665 673512 292670 673568
rect 292726 673512 299428 673568
rect 292665 673510 299428 673512
rect 162209 673507 162275 673510
rect 166901 673507 166967 673510
rect 292665 673507 292731 673510
rect 299422 673508 299428 673510
rect 299492 673508 299498 673572
rect 325558 673570 325618 673646
rect 325742 673570 325802 673782
rect 335310 673706 335370 673782
rect 345062 673840 347839 673842
rect 345062 673784 347778 673840
rect 347834 673784 347839 673840
rect 345062 673782 347839 673784
rect 335310 673646 344938 673706
rect 325558 673510 325802 673570
rect 344878 673570 344938 673646
rect 345062 673570 345122 673782
rect 347773 673779 347839 673782
rect 371969 673842 372035 673845
rect 376702 673842 376708 673844
rect 371969 673840 376708 673842
rect 371969 673784 371974 673840
rect 372030 673784 376708 673840
rect 371969 673782 376708 673784
rect 371969 673779 372035 673782
rect 376702 673780 376708 673782
rect 376772 673780 376778 673844
rect 379513 673842 379579 673845
rect 540973 673842 541039 673845
rect 379513 673840 393330 673842
rect 379513 673784 379518 673840
rect 379574 673784 393330 673840
rect 379513 673782 393330 673784
rect 379513 673779 379579 673782
rect 393270 673706 393330 673782
rect 403022 673782 412650 673842
rect 393270 673646 402898 673706
rect 344878 673510 345122 673570
rect 355409 673570 355475 673573
rect 357382 673570 357388 673572
rect 355409 673568 357388 673570
rect 355409 673512 355414 673568
rect 355470 673512 357388 673568
rect 355409 673510 357388 673512
rect 355409 673507 355475 673510
rect 357382 673508 357388 673510
rect 357452 673508 357458 673572
rect 402838 673570 402898 673646
rect 403022 673570 403082 673782
rect 412590 673706 412650 673782
rect 431910 673782 441538 673842
rect 412590 673646 422218 673706
rect 402838 673510 403082 673570
rect 422158 673570 422218 673646
rect 431910 673570 431970 673782
rect 422158 673510 431970 673570
rect 441478 673570 441538 673782
rect 441662 673782 451290 673842
rect 441662 673570 441722 673782
rect 451230 673706 451290 673782
rect 460982 673782 470610 673842
rect 451230 673646 460858 673706
rect 441478 673510 441722 673570
rect 460798 673570 460858 673646
rect 460982 673570 461042 673782
rect 470550 673706 470610 673782
rect 480302 673782 489930 673842
rect 470550 673646 480178 673706
rect 460798 673510 461042 673570
rect 480118 673570 480178 673646
rect 480302 673570 480362 673782
rect 489870 673706 489930 673782
rect 499622 673782 509250 673842
rect 489870 673646 499498 673706
rect 480118 673510 480362 673570
rect 499438 673570 499498 673646
rect 499622 673570 499682 673782
rect 509190 673706 509250 673782
rect 518942 673782 528570 673842
rect 509190 673646 518818 673706
rect 499438 673510 499682 673570
rect 518758 673570 518818 673646
rect 518942 673570 519002 673782
rect 528510 673706 528570 673782
rect 538262 673840 541039 673842
rect 538262 673784 540978 673840
rect 541034 673784 541039 673840
rect 538262 673782 541039 673784
rect 528510 673646 538138 673706
rect 518758 673510 519002 673570
rect 538078 673570 538138 673646
rect 538262 673570 538322 673782
rect 540973 673779 541039 673782
rect 565169 673842 565235 673845
rect 572713 673842 572779 673845
rect 565169 673840 569970 673842
rect 565169 673784 565174 673840
rect 565230 673784 569970 673840
rect 565169 673782 569970 673784
rect 565169 673779 565235 673782
rect 569910 673706 569970 673782
rect 572713 673840 576962 673842
rect 572713 673784 572718 673840
rect 572774 673784 576962 673840
rect 572713 673782 576962 673784
rect 572713 673779 572779 673782
rect 572621 673706 572687 673709
rect 569910 673704 572687 673706
rect 569910 673648 572626 673704
rect 572682 673648 572687 673704
rect 569910 673646 572687 673648
rect 576902 673706 576962 673782
rect 583342 673706 583402 674598
rect 583520 674508 584960 674598
rect 576902 673646 583402 673706
rect 572621 673643 572687 673646
rect 538078 673510 538322 673570
rect 548609 673570 548675 673573
rect 553301 673570 553367 673573
rect 548609 673568 553367 673570
rect 548609 673512 548614 673568
rect 548670 673512 553306 673568
rect 553362 673512 553367 673568
rect 548609 673510 553367 673512
rect 548609 673507 548675 673510
rect 553301 673507 553367 673510
rect -960 667994 480 668084
rect 3509 667994 3575 667997
rect -960 667992 3575 667994
rect -960 667936 3514 667992
rect 3570 667936 3575 667992
rect -960 667934 3575 667936
rect -960 667844 480 667934
rect 3509 667931 3575 667934
rect 583520 662676 584960 662916
rect -960 653578 480 653668
rect 3049 653578 3115 653581
rect -960 653576 3115 653578
rect -960 653520 3054 653576
rect 3110 653520 3115 653576
rect -960 653518 3115 653520
rect -960 653428 480 653518
rect 3049 653515 3115 653518
rect 129273 652900 129339 652901
rect 133689 652900 133755 652901
rect 258625 652900 258691 652901
rect 129222 652898 129228 652900
rect 129182 652838 129228 652898
rect 129292 652896 129339 652900
rect 133638 652898 133644 652900
rect 129334 652840 129339 652896
rect 129222 652836 129228 652838
rect 129292 652836 129339 652840
rect 133598 652838 133644 652898
rect 133708 652896 133755 652900
rect 258574 652898 258580 652900
rect 133750 652840 133755 652896
rect 133638 652836 133644 652838
rect 133708 652836 133755 652840
rect 258534 652838 258580 652898
rect 258644 652896 258691 652900
rect 258686 652840 258691 652896
rect 258574 652836 258580 652838
rect 258644 652836 258691 652840
rect 129273 652835 129339 652836
rect 133689 652835 133755 652836
rect 258625 652835 258691 652836
rect 378133 652900 378199 652901
rect 383469 652900 383535 652901
rect 378133 652896 378180 652900
rect 378244 652898 378250 652900
rect 378133 652840 378138 652896
rect 378133 652836 378180 652840
rect 378244 652838 378290 652898
rect 383469 652896 383516 652900
rect 383580 652898 383586 652900
rect 383469 652840 383474 652896
rect 378244 652836 378250 652838
rect 383469 652836 383516 652840
rect 383580 652838 383626 652898
rect 383580 652836 383586 652838
rect 378133 652835 378199 652836
rect 383469 652835 383535 652836
rect 263501 651676 263567 651677
rect 263501 651672 263571 651676
rect 263501 651616 263506 651672
rect 263562 651616 263571 651672
rect 263501 651612 263571 651616
rect 263635 651674 263641 651676
rect 263635 651614 263658 651674
rect 263635 651612 263641 651614
rect 263501 651611 263567 651612
rect 376702 651340 376708 651404
rect 376772 651402 376778 651404
rect 386321 651402 386387 651405
rect 376772 651400 386387 651402
rect 376772 651344 386326 651400
rect 386382 651344 386387 651400
rect 376772 651342 386387 651344
rect 376772 651340 376778 651342
rect 386321 651339 386387 651342
rect 370405 651130 370471 651133
rect 376702 651130 376708 651132
rect 370405 651128 376708 651130
rect 370405 651072 370410 651128
rect 370466 651072 376708 651128
rect 370405 651070 376708 651072
rect 370405 651067 370471 651070
rect 376702 651068 376708 651070
rect 376772 651068 376778 651132
rect 396022 651068 396028 651132
rect 396092 651130 396098 651132
rect 400857 651130 400923 651133
rect 396092 651128 400923 651130
rect 396092 651072 400862 651128
rect 400918 651072 400923 651128
rect 396092 651070 400923 651072
rect 396092 651068 396098 651070
rect 400857 651067 400923 651070
rect 583385 651130 583451 651133
rect 583520 651130 584960 651220
rect 583385 651128 584960 651130
rect 583385 651072 583390 651128
rect 583446 651072 584960 651128
rect 583385 651070 584960 651072
rect 583385 651067 583451 651070
rect 135161 650994 135227 650997
rect 140037 650994 140103 650997
rect 135161 650992 140103 650994
rect 135161 650936 135166 650992
rect 135222 650936 140042 650992
rect 140098 650936 140103 650992
rect 135161 650934 140103 650936
rect 135161 650931 135227 650934
rect 140037 650931 140103 650934
rect 311985 650994 312051 650997
rect 318742 650994 318748 650996
rect 311985 650992 318748 650994
rect 311985 650936 311990 650992
rect 312046 650936 318748 650992
rect 311985 650934 318748 650936
rect 311985 650931 312051 650934
rect 318742 650932 318748 650934
rect 318812 650932 318818 650996
rect 386321 650994 386387 650997
rect 389173 650994 389239 650997
rect 386321 650992 389239 650994
rect 386321 650936 386326 650992
rect 386382 650936 389178 650992
rect 389234 650936 389239 650992
rect 583520 650980 584960 651070
rect 386321 650934 389239 650936
rect 386321 650931 386387 650934
rect 389173 650931 389239 650934
rect 58198 650796 58204 650860
rect 58268 650858 58274 650860
rect 120717 650858 120783 650861
rect 125542 650858 125548 650860
rect 58268 650798 70410 650858
rect 58268 650796 58274 650798
rect 70350 650586 70410 650798
rect 120717 650856 125548 650858
rect 120717 650800 120722 650856
rect 120778 650800 125548 650856
rect 120717 650798 125548 650800
rect 120717 650795 120783 650798
rect 125542 650796 125548 650798
rect 125612 650796 125618 650860
rect 309041 650858 309107 650861
rect 311801 650858 311867 650861
rect 367093 650858 367159 650861
rect 146894 650798 167010 650858
rect 89621 650722 89687 650725
rect 106733 650722 106799 650725
rect 80102 650720 89687 650722
rect 80102 650664 89626 650720
rect 89682 650664 89687 650720
rect 80102 650662 89687 650664
rect 80102 650586 80162 650662
rect 89621 650659 89687 650662
rect 99422 650720 106799 650722
rect 99422 650664 106738 650720
rect 106794 650664 106799 650720
rect 99422 650662 106799 650664
rect 70350 650526 80162 650586
rect 96521 650586 96587 650589
rect 99422 650586 99482 650662
rect 106733 650659 106799 650662
rect 140129 650722 140195 650725
rect 146894 650722 146954 650798
rect 140129 650720 146954 650722
rect 140129 650664 140134 650720
rect 140190 650664 146954 650720
rect 140129 650662 146954 650664
rect 140129 650659 140195 650662
rect 96521 650584 99482 650586
rect 96521 650528 96526 650584
rect 96582 650528 99482 650584
rect 96521 650526 99482 650528
rect 115749 650586 115815 650589
rect 115933 650586 115999 650589
rect 115749 650584 115999 650586
rect 115749 650528 115754 650584
rect 115810 650528 115938 650584
rect 115994 650528 115999 650584
rect 115749 650526 115999 650528
rect 96521 650523 96587 650526
rect 115749 650523 115815 650526
rect 115933 650523 115999 650526
rect 125542 650524 125548 650588
rect 125612 650586 125618 650588
rect 135161 650586 135227 650589
rect 125612 650584 135227 650586
rect 125612 650528 135166 650584
rect 135222 650528 135227 650584
rect 125612 650526 135227 650528
rect 166950 650586 167010 650798
rect 309041 650856 311867 650858
rect 309041 650800 309046 650856
rect 309102 650800 311806 650856
rect 311862 650800 311867 650856
rect 309041 650798 311867 650800
rect 309041 650795 309107 650798
rect 311801 650795 311867 650798
rect 360150 650856 367159 650858
rect 360150 650800 367098 650856
rect 367154 650800 367159 650856
rect 360150 650798 367159 650800
rect 278773 650722 278839 650725
rect 176702 650662 186146 650722
rect 176702 650586 176762 650662
rect 166950 650526 176762 650586
rect 186086 650586 186146 650662
rect 196022 650662 203626 650722
rect 196022 650586 196082 650662
rect 186086 650526 196082 650586
rect 203566 650586 203626 650662
rect 215342 650662 221474 650722
rect 215342 650586 215402 650662
rect 203566 650526 215402 650586
rect 221414 650586 221474 650662
rect 234662 650662 242266 650722
rect 234662 650586 234722 650662
rect 221414 650526 234722 650586
rect 237373 650586 237439 650589
rect 237557 650586 237623 650589
rect 237373 650584 237623 650586
rect 237373 650528 237378 650584
rect 237434 650528 237562 650584
rect 237618 650528 237623 650584
rect 237373 650526 237623 650528
rect 242206 650586 242266 650662
rect 253982 650662 263633 650722
rect 253982 650586 254042 650662
rect 242206 650526 254042 650586
rect 263573 650586 263633 650662
rect 273302 650720 278839 650722
rect 273302 650664 278778 650720
rect 278834 650664 278839 650720
rect 273302 650662 278839 650664
rect 273302 650586 273362 650662
rect 278773 650659 278839 650662
rect 292665 650722 292731 650725
rect 299422 650722 299428 650724
rect 292665 650720 299428 650722
rect 292665 650664 292670 650720
rect 292726 650664 299428 650720
rect 292665 650662 299428 650664
rect 292665 650659 292731 650662
rect 299422 650660 299428 650662
rect 299492 650660 299498 650724
rect 340781 650722 340847 650725
rect 331262 650720 340847 650722
rect 331262 650664 340786 650720
rect 340842 650664 340847 650720
rect 331262 650662 340847 650664
rect 263573 650526 273362 650586
rect 288341 650586 288407 650589
rect 289813 650586 289879 650589
rect 288341 650584 289879 650586
rect 288341 650528 288346 650584
rect 288402 650528 289818 650584
rect 289874 650528 289879 650584
rect 288341 650526 289879 650528
rect 125612 650524 125618 650526
rect 135161 650523 135227 650526
rect 237373 650523 237439 650526
rect 237557 650523 237623 650526
rect 288341 650523 288407 650526
rect 289813 650523 289879 650526
rect 318742 650524 318748 650588
rect 318812 650586 318818 650588
rect 321461 650586 321527 650589
rect 318812 650584 321527 650586
rect 318812 650528 321466 650584
rect 321522 650528 321527 650584
rect 318812 650526 321527 650528
rect 318812 650524 318818 650526
rect 321461 650523 321527 650526
rect 321645 650586 321711 650589
rect 331262 650586 331322 650662
rect 340781 650659 340847 650662
rect 321645 650584 331322 650586
rect 321645 650528 321650 650584
rect 321706 650528 331322 650584
rect 321645 650526 331322 650528
rect 347681 650586 347747 650589
rect 360150 650586 360210 650798
rect 367093 650795 367159 650798
rect 389265 650858 389331 650861
rect 396022 650858 396028 650860
rect 389265 650856 396028 650858
rect 389265 650800 389270 650856
rect 389326 650800 396028 650856
rect 389265 650798 396028 650800
rect 389265 650795 389331 650798
rect 396022 650796 396028 650798
rect 396092 650796 396098 650860
rect 434662 650796 434668 650860
rect 434732 650858 434738 650860
rect 444281 650858 444347 650861
rect 434732 650856 444347 650858
rect 434732 650800 444286 650856
rect 444342 650800 444347 650856
rect 434732 650798 444347 650800
rect 434732 650796 434738 650798
rect 444281 650795 444347 650798
rect 563145 650858 563211 650861
rect 563145 650856 569970 650858
rect 563145 650800 563150 650856
rect 563206 650800 569970 650856
rect 563145 650798 569970 650800
rect 563145 650795 563211 650798
rect 569910 650722 569970 650798
rect 579654 650796 579660 650860
rect 579724 650858 579730 650860
rect 583385 650858 583451 650861
rect 579724 650856 583451 650858
rect 579724 650800 583390 650856
rect 583446 650800 583451 650856
rect 579724 650798 583451 650800
rect 579724 650796 579730 650798
rect 583385 650795 583451 650798
rect 572621 650722 572687 650725
rect 569910 650720 572687 650722
rect 569910 650664 572626 650720
rect 572682 650664 572687 650720
rect 569910 650662 572687 650664
rect 572621 650659 572687 650662
rect 579521 650722 579587 650725
rect 579521 650720 579722 650722
rect 579521 650664 579526 650720
rect 579582 650664 579722 650720
rect 579521 650662 579722 650664
rect 579521 650659 579587 650662
rect 347681 650584 360210 650586
rect 347681 650528 347686 650584
rect 347742 650528 360210 650584
rect 347681 650526 360210 650528
rect 400857 650586 400923 650589
rect 405733 650586 405799 650589
rect 400857 650584 405799 650586
rect 400857 650528 400862 650584
rect 400918 650528 405738 650584
rect 405794 650528 405799 650584
rect 400857 650526 405799 650528
rect 321645 650523 321711 650526
rect 347681 650523 347747 650526
rect 400857 650523 400923 650526
rect 405733 650523 405799 650526
rect 418245 650586 418311 650589
rect 444281 650586 444347 650589
rect 463601 650586 463667 650589
rect 482921 650586 482987 650589
rect 502241 650586 502307 650589
rect 521561 650586 521627 650589
rect 540881 650586 540947 650589
rect 560293 650586 560359 650589
rect 579662 650588 579722 650662
rect 418245 650584 427922 650586
rect 418245 650528 418250 650584
rect 418306 650528 427922 650584
rect 418245 650526 427922 650528
rect 418245 650523 418311 650526
rect 299422 650388 299428 650452
rect 299492 650450 299498 650452
rect 309041 650450 309107 650453
rect 299492 650448 309107 650450
rect 299492 650392 309046 650448
rect 309102 650392 309107 650448
rect 299492 650390 309107 650392
rect 427862 650450 427922 650526
rect 444281 650584 447242 650586
rect 444281 650528 444286 650584
rect 444342 650528 447242 650584
rect 444281 650526 447242 650528
rect 444281 650523 444347 650526
rect 434662 650450 434668 650452
rect 427862 650390 434668 650450
rect 299492 650388 299498 650390
rect 309041 650387 309107 650390
rect 434662 650388 434668 650390
rect 434732 650388 434738 650452
rect 447182 650450 447242 650526
rect 463601 650584 466562 650586
rect 463601 650528 463606 650584
rect 463662 650528 466562 650584
rect 463601 650526 466562 650528
rect 463601 650523 463667 650526
rect 456701 650450 456767 650453
rect 447182 650448 456767 650450
rect 447182 650392 456706 650448
rect 456762 650392 456767 650448
rect 447182 650390 456767 650392
rect 466502 650450 466562 650526
rect 482921 650584 485882 650586
rect 482921 650528 482926 650584
rect 482982 650528 485882 650584
rect 482921 650526 485882 650528
rect 482921 650523 482987 650526
rect 476021 650450 476087 650453
rect 466502 650448 476087 650450
rect 466502 650392 476026 650448
rect 476082 650392 476087 650448
rect 466502 650390 476087 650392
rect 485822 650450 485882 650526
rect 502241 650584 505202 650586
rect 502241 650528 502246 650584
rect 502302 650528 505202 650584
rect 502241 650526 505202 650528
rect 502241 650523 502307 650526
rect 495341 650450 495407 650453
rect 485822 650448 495407 650450
rect 485822 650392 495346 650448
rect 495402 650392 495407 650448
rect 485822 650390 495407 650392
rect 505142 650450 505202 650526
rect 521561 650584 524522 650586
rect 521561 650528 521566 650584
rect 521622 650528 524522 650584
rect 521561 650526 524522 650528
rect 521561 650523 521627 650526
rect 514661 650450 514727 650453
rect 505142 650448 514727 650450
rect 505142 650392 514666 650448
rect 514722 650392 514727 650448
rect 505142 650390 514727 650392
rect 524462 650450 524522 650526
rect 540881 650584 543842 650586
rect 540881 650528 540886 650584
rect 540942 650528 543842 650584
rect 540881 650526 543842 650528
rect 540881 650523 540947 650526
rect 533981 650450 534047 650453
rect 524462 650448 534047 650450
rect 524462 650392 533986 650448
rect 534042 650392 534047 650448
rect 524462 650390 534047 650392
rect 543782 650450 543842 650526
rect 560158 650584 560359 650586
rect 560158 650528 560298 650584
rect 560354 650528 560359 650584
rect 560158 650526 560359 650528
rect 543782 650390 550650 650450
rect 456701 650387 456767 650390
rect 476021 650387 476087 650390
rect 495341 650387 495407 650390
rect 514661 650387 514727 650390
rect 533981 650387 534047 650390
rect 418061 650314 418127 650317
rect 415350 650312 418127 650314
rect 415350 650256 418066 650312
rect 418122 650256 418127 650312
rect 415350 650254 418127 650256
rect 413369 650178 413435 650181
rect 415350 650178 415410 650254
rect 418061 650251 418127 650254
rect 413369 650176 415410 650178
rect 413369 650120 413374 650176
rect 413430 650120 415410 650176
rect 413369 650118 415410 650120
rect 550590 650178 550650 650390
rect 560158 650178 560218 650526
rect 560293 650523 560359 650526
rect 579654 650524 579660 650588
rect 579724 650524 579730 650588
rect 550590 650118 560218 650178
rect 413369 650115 413435 650118
rect 270493 650042 270559 650045
rect 280061 650042 280127 650045
rect 270493 650040 280127 650042
rect 270493 649984 270498 650040
rect 270554 649984 280066 650040
rect 280122 649984 280127 650040
rect 270493 649982 280127 649984
rect 270493 649979 270559 649982
rect 280061 649979 280127 649982
rect 266445 649906 266511 649909
rect 386413 649906 386479 649909
rect 266445 649904 266554 649906
rect 266445 649848 266450 649904
rect 266506 649848 266554 649904
rect 266445 649843 266554 649848
rect 386413 649904 386522 649906
rect 386413 649848 386418 649904
rect 386474 649848 386522 649904
rect 386413 649843 386522 649848
rect 137645 649713 137711 649716
rect 137172 649711 137711 649713
rect 137172 649655 137650 649711
rect 137706 649655 137711 649711
rect 266494 649683 266554 649843
rect 386462 649683 386522 649843
rect 137172 649653 137711 649655
rect 137645 649650 137711 649653
rect 57605 646098 57671 646101
rect 60046 646098 60106 646587
rect 57605 646096 60106 646098
rect 57605 646040 57610 646096
rect 57666 646040 60106 646096
rect 57605 646038 60106 646040
rect 188337 646098 188403 646101
rect 190134 646098 190194 646587
rect 307109 646370 307175 646373
rect 310102 646370 310162 646587
rect 307109 646368 310162 646370
rect 307109 646312 307114 646368
rect 307170 646312 310162 646368
rect 307109 646310 310162 646312
rect 307109 646307 307175 646310
rect 188337 646096 190194 646098
rect 188337 646040 188342 646096
rect 188398 646040 190194 646096
rect 188337 646038 190194 646040
rect 57605 646035 57671 646038
rect 188337 646035 188403 646038
rect 57513 645010 57579 645013
rect 60046 645010 60106 645459
rect 57513 645008 60106 645010
rect 57513 644952 57518 645008
rect 57574 644952 60106 645008
rect 57513 644950 60106 644952
rect 188429 645010 188495 645013
rect 190134 645010 190194 645459
rect 188429 645008 190194 645010
rect 188429 644952 188434 645008
rect 188490 644952 190194 645008
rect 188429 644950 190194 644952
rect 307109 645010 307175 645013
rect 310102 645010 310162 645459
rect 307109 645008 310162 645010
rect 307109 644952 307114 645008
rect 307170 644952 310162 645008
rect 307109 644950 310162 644952
rect 57513 644947 57579 644950
rect 188429 644947 188495 644950
rect 307109 644947 307175 644950
rect 57421 643242 57487 643245
rect 60046 643242 60106 643759
rect 57421 643240 60106 643242
rect 57421 643184 57426 643240
rect 57482 643184 60106 643240
rect 57421 643182 60106 643184
rect 188521 643242 188587 643245
rect 190134 643242 190194 643759
rect 307109 643514 307175 643517
rect 310102 643514 310162 643759
rect 307109 643512 310162 643514
rect 307109 643456 307114 643512
rect 307170 643456 310162 643512
rect 307109 643454 310162 643456
rect 307109 643451 307175 643454
rect 188521 643240 190194 643242
rect 188521 643184 188526 643240
rect 188582 643184 190194 643240
rect 188521 643182 190194 643184
rect 57421 643179 57487 643182
rect 188521 643179 188587 643182
rect 57329 642018 57395 642021
rect 60046 642018 60106 642631
rect 57329 642016 60106 642018
rect 57329 641960 57334 642016
rect 57390 641960 60106 642016
rect 57329 641958 60106 641960
rect 188613 642018 188679 642021
rect 190134 642018 190194 642631
rect 307661 642154 307727 642157
rect 310102 642154 310162 642631
rect 307661 642152 310162 642154
rect 307661 642096 307666 642152
rect 307722 642096 310162 642152
rect 307661 642094 310162 642096
rect 307661 642091 307727 642094
rect 188613 642016 190194 642018
rect 188613 641960 188618 642016
rect 188674 641960 190194 642016
rect 188613 641958 190194 641960
rect 57329 641955 57395 641958
rect 188613 641955 188679 641958
rect 57237 640386 57303 640389
rect 60046 640386 60106 640931
rect 57237 640384 60106 640386
rect 57237 640328 57242 640384
rect 57298 640328 60106 640384
rect 57237 640326 60106 640328
rect 188705 640386 188771 640389
rect 190134 640386 190194 640931
rect 307661 640522 307727 640525
rect 310102 640522 310162 640931
rect 307661 640520 310162 640522
rect 307661 640464 307666 640520
rect 307722 640464 310162 640520
rect 307661 640462 310162 640464
rect 307661 640459 307727 640462
rect 188705 640384 190194 640386
rect 188705 640328 188710 640384
rect 188766 640328 190194 640384
rect 188705 640326 190194 640328
rect 57237 640323 57303 640326
rect 188705 640323 188771 640326
rect 57053 639298 57119 639301
rect 60046 639298 60106 639803
rect 57053 639296 60106 639298
rect -960 639012 480 639252
rect 57053 639240 57058 639296
rect 57114 639240 60106 639296
rect 57053 639238 60106 639240
rect 188889 639298 188955 639301
rect 190134 639298 190194 639803
rect 306649 639434 306715 639437
rect 310102 639434 310162 639803
rect 306649 639432 310162 639434
rect 306649 639376 306654 639432
rect 306710 639376 310162 639432
rect 306649 639374 310162 639376
rect 580257 639434 580323 639437
rect 583520 639434 584960 639524
rect 580257 639432 584960 639434
rect 580257 639376 580262 639432
rect 580318 639376 584960 639432
rect 580257 639374 584960 639376
rect 306649 639371 306715 639374
rect 580257 639371 580323 639374
rect 188889 639296 190194 639298
rect 188889 639240 188894 639296
rect 188950 639240 190194 639296
rect 583520 639284 584960 639374
rect 188889 639238 190194 639240
rect 57053 639235 57119 639238
rect 188889 639235 188955 639238
rect 57145 637666 57211 637669
rect 60046 637666 60106 638103
rect 57145 637664 60106 637666
rect 57145 637608 57150 637664
rect 57206 637608 60106 637664
rect 57145 637606 60106 637608
rect 188245 637666 188311 637669
rect 190134 637666 190194 638103
rect 306833 637938 306899 637941
rect 310102 637938 310162 638103
rect 306833 637936 310162 637938
rect 306833 637880 306838 637936
rect 306894 637880 310162 637936
rect 306833 637878 310162 637880
rect 306833 637875 306899 637878
rect 188245 637664 190194 637666
rect 188245 637608 188250 637664
rect 188306 637608 190194 637664
rect 188245 637606 190194 637608
rect 57145 637603 57211 637606
rect 188245 637603 188311 637606
rect 580349 627738 580415 627741
rect 583520 627738 584960 627828
rect 580349 627736 584960 627738
rect 580349 627680 580354 627736
rect 580410 627680 584960 627736
rect 580349 627678 584960 627680
rect 580349 627675 580415 627678
rect 583520 627588 584960 627678
rect -960 624882 480 624972
rect 3509 624882 3575 624885
rect -960 624880 3575 624882
rect -960 624824 3514 624880
rect 3570 624824 3575 624880
rect -960 624822 3575 624824
rect -960 624732 480 624822
rect 3509 624819 3575 624822
rect 583520 615756 584960 615996
rect -960 610466 480 610556
rect 3601 610466 3667 610469
rect -960 610464 3667 610466
rect -960 610408 3606 610464
rect 3662 610408 3667 610464
rect -960 610406 3667 610408
rect -960 610316 480 610406
rect 3601 610403 3667 610406
rect 580441 604210 580507 604213
rect 583520 604210 584960 604300
rect 580441 604208 584960 604210
rect 580441 604152 580446 604208
rect 580502 604152 584960 604208
rect 580441 604150 584960 604152
rect 580441 604147 580507 604150
rect 583520 604060 584960 604150
rect -960 596050 480 596140
rect 3325 596050 3391 596053
rect -960 596048 3391 596050
rect -960 595992 3330 596048
rect 3386 595992 3391 596048
rect -960 595990 3391 595992
rect -960 595900 480 595990
rect 3325 595987 3391 595990
rect 580625 592514 580691 592517
rect 583520 592514 584960 592604
rect 580625 592512 584960 592514
rect 580625 592456 580630 592512
rect 580686 592456 584960 592512
rect 580625 592454 584960 592456
rect 580625 592451 580691 592454
rect 583520 592364 584960 592454
rect 139393 589658 139459 589661
rect 387793 589658 387859 589661
rect 136958 589656 139459 589658
rect 136958 589600 139398 589656
rect 139454 589600 139459 589656
rect 136958 589598 139459 589600
rect 136958 586614 137018 589598
rect 139393 589595 139459 589598
rect 387014 589656 387859 589658
rect 387014 589600 387798 589656
rect 387854 589600 387859 589656
rect 387014 589598 387859 589600
rect 267230 589386 267290 589412
rect 269113 589386 269179 589389
rect 270401 589386 270467 589389
rect 267230 589384 270467 589386
rect 267230 589328 269118 589384
rect 269174 589328 270406 589384
rect 270462 589328 270467 589384
rect 267230 589326 270467 589328
rect 269113 589323 269179 589326
rect 270401 589323 270467 589326
rect 299657 589386 299723 589389
rect 299933 589386 299999 589389
rect 299657 589384 299999 589386
rect 299657 589328 299662 589384
rect 299718 589328 299938 589384
rect 299994 589328 299999 589384
rect 299657 589326 299999 589328
rect 299657 589323 299723 589326
rect 299933 589323 299999 589326
rect 269113 587754 269179 587757
rect 267230 587752 269179 587754
rect 267230 587696 269118 587752
rect 269174 587696 269179 587752
rect 267230 587694 269179 587696
rect 136958 586584 137172 586614
rect 136988 586554 137202 586584
rect -960 581620 480 581860
rect 137142 580928 137202 586554
rect 267230 580928 267290 587694
rect 269113 587691 269179 587694
rect 387014 586614 387074 589598
rect 387793 589595 387859 589598
rect 387014 586584 387228 586614
rect 387044 586554 387258 586584
rect 387198 580954 387258 586554
rect 389173 580954 389239 580957
rect 387198 580952 389239 580954
rect 387198 580896 389178 580952
rect 389234 580896 389239 580952
rect 387198 580894 389239 580896
rect 389173 580891 389239 580894
rect 580717 580818 580783 580821
rect 583520 580818 584960 580908
rect 580717 580816 584960 580818
rect 580717 580760 580722 580816
rect 580778 580760 584960 580816
rect 580717 580758 584960 580760
rect 580717 580755 580783 580758
rect 583520 580668 584960 580758
rect 56961 579730 57027 579733
rect 60046 579730 60106 580255
rect 56961 579728 60106 579730
rect 56961 579672 56966 579728
rect 57022 579672 60106 579728
rect 56961 579670 60106 579672
rect 188797 579730 188863 579733
rect 190134 579730 190194 580255
rect 188797 579728 190194 579730
rect 188797 579672 188802 579728
rect 188858 579672 190194 579728
rect 188797 579670 190194 579672
rect 307017 579730 307083 579733
rect 310102 579730 310162 580255
rect 307017 579728 310162 579730
rect 307017 579672 307022 579728
rect 307078 579672 310162 579728
rect 307017 579670 310162 579672
rect 56961 579667 57027 579670
rect 188797 579667 188863 579670
rect 307017 579667 307083 579670
rect 56869 578370 56935 578373
rect 60046 578370 60106 578555
rect 56869 578368 60106 578370
rect 56869 578312 56874 578368
rect 56930 578312 60106 578368
rect 56869 578310 60106 578312
rect 188981 578370 189047 578373
rect 190134 578370 190194 578555
rect 188981 578368 190194 578370
rect 188981 578312 188986 578368
rect 189042 578312 190194 578368
rect 188981 578310 190194 578312
rect 305637 578370 305703 578373
rect 310102 578370 310162 578555
rect 305637 578368 310162 578370
rect 305637 578312 305642 578368
rect 305698 578312 310162 578368
rect 305637 578310 310162 578312
rect 56869 578307 56935 578310
rect 188981 578307 189047 578310
rect 305637 578307 305703 578310
rect 583520 568836 584960 569076
rect -960 567354 480 567444
rect 3601 567354 3667 567357
rect -960 567352 3667 567354
rect -960 567296 3606 567352
rect 3662 567296 3667 567352
rect -960 567294 3667 567296
rect -960 567204 480 567294
rect 3601 567291 3667 567294
rect 210969 560010 211035 560013
rect 211102 560010 211108 560012
rect 210969 560008 211108 560010
rect 210969 559952 210974 560008
rect 211030 559952 211108 560008
rect 210969 559950 211108 559952
rect 210969 559947 211035 559950
rect 211102 559948 211108 559950
rect 211172 559948 211178 560012
rect 328474 559812 328480 559876
rect 328544 559874 328550 559876
rect 329097 559874 329163 559877
rect 337745 559876 337811 559877
rect 337694 559874 337700 559876
rect 328544 559872 337700 559874
rect 337764 559874 337811 559876
rect 357709 559874 357775 559877
rect 358842 559874 358848 559876
rect 337764 559872 337892 559874
rect 328544 559816 329102 559872
rect 329158 559816 337700 559872
rect 337806 559816 337892 559872
rect 328544 559814 337700 559816
rect 328544 559812 328550 559814
rect 329097 559811 329163 559814
rect 337694 559812 337700 559814
rect 337764 559814 337892 559816
rect 357709 559872 358848 559874
rect 357709 559816 357714 559872
rect 357770 559816 358848 559872
rect 357709 559814 358848 559816
rect 337764 559812 337811 559814
rect 337745 559811 337811 559812
rect 357709 559811 357775 559814
rect 358842 559812 358848 559814
rect 358912 559812 358918 559876
rect 358854 559676 358860 559740
rect 358924 559738 358930 559740
rect 359406 559738 359412 559740
rect 358924 559678 359412 559738
rect 358924 559676 358930 559678
rect 359406 559676 359412 559678
rect 359476 559676 359482 559740
rect 348141 559330 348207 559333
rect 351862 559330 351868 559332
rect 348141 559328 351868 559330
rect 348141 559272 348146 559328
rect 348202 559272 351868 559328
rect 348141 559270 351868 559272
rect 348141 559267 348207 559270
rect 351862 559268 351868 559270
rect 351932 559268 351938 559332
rect 348049 559194 348115 559197
rect 352230 559194 352236 559196
rect 348049 559192 352236 559194
rect 348049 559136 348054 559192
rect 348110 559136 352236 559192
rect 348049 559134 352236 559136
rect 348049 559131 348115 559134
rect 352230 559132 352236 559134
rect 352300 559132 352306 559196
rect 220077 559060 220143 559061
rect 220077 559056 220124 559060
rect 220188 559058 220194 559060
rect 220077 559000 220082 559056
rect 220077 558996 220124 559000
rect 220188 558998 220234 559058
rect 220188 558996 220194 558998
rect 220077 558995 220143 558996
rect 67398 558860 67404 558924
rect 67468 558922 67474 558924
rect 67541 558922 67607 558925
rect 67468 558920 67607 558922
rect 67468 558864 67546 558920
rect 67602 558864 67607 558920
rect 67468 558862 67607 558864
rect 67468 558860 67474 558862
rect 67541 558859 67607 558862
rect 68502 558860 68508 558924
rect 68572 558922 68578 558924
rect 68921 558922 68987 558925
rect 68572 558920 68987 558922
rect 68572 558864 68926 558920
rect 68982 558864 68987 558920
rect 68572 558862 68987 558864
rect 68572 558860 68578 558862
rect 68921 558859 68987 558862
rect 70158 558860 70164 558924
rect 70228 558922 70234 558924
rect 70301 558922 70367 558925
rect 71681 558924 71747 558925
rect 70228 558920 70367 558922
rect 70228 558864 70306 558920
rect 70362 558864 70367 558920
rect 70228 558862 70367 558864
rect 70228 558860 70234 558862
rect 70301 558859 70367 558862
rect 71630 558860 71636 558924
rect 71700 558922 71747 558924
rect 71700 558920 71792 558922
rect 71742 558864 71792 558920
rect 71700 558862 71792 558864
rect 71700 558860 71747 558862
rect 72366 558860 72372 558924
rect 72436 558922 72442 558924
rect 72601 558922 72667 558925
rect 72436 558920 72667 558922
rect 72436 558864 72606 558920
rect 72662 558864 72667 558920
rect 72436 558862 72667 558864
rect 72436 558860 72442 558862
rect 71681 558859 71747 558860
rect 72601 558859 72667 558862
rect 72918 558860 72924 558924
rect 72988 558922 72994 558924
rect 73061 558922 73127 558925
rect 72988 558920 73127 558922
rect 72988 558864 73066 558920
rect 73122 558864 73127 558920
rect 72988 558862 73127 558864
rect 72988 558860 72994 558862
rect 73061 558859 73127 558862
rect 73654 558860 73660 558924
rect 73724 558922 73730 558924
rect 73797 558922 73863 558925
rect 74257 558924 74323 558925
rect 74993 558924 75059 558925
rect 74206 558922 74212 558924
rect 73724 558920 73863 558922
rect 73724 558864 73802 558920
rect 73858 558864 73863 558920
rect 73724 558862 73863 558864
rect 74166 558862 74212 558922
rect 74276 558920 74323 558924
rect 74942 558922 74948 558924
rect 74318 558864 74323 558920
rect 73724 558860 73730 558862
rect 73797 558859 73863 558862
rect 74206 558860 74212 558862
rect 74276 558860 74323 558864
rect 74902 558862 74948 558922
rect 75012 558920 75059 558924
rect 75054 558864 75059 558920
rect 74942 558860 74948 558862
rect 75012 558860 75059 558864
rect 75862 558860 75868 558924
rect 75932 558922 75938 558924
rect 76005 558922 76071 558925
rect 76833 558924 76899 558925
rect 77385 558924 77451 558925
rect 78489 558924 78555 558925
rect 76782 558922 76788 558924
rect 75932 558920 76071 558922
rect 75932 558864 76010 558920
rect 76066 558864 76071 558920
rect 75932 558862 76071 558864
rect 76742 558862 76788 558922
rect 76852 558920 76899 558924
rect 77334 558922 77340 558924
rect 76894 558864 76899 558920
rect 75932 558860 75938 558862
rect 74257 558859 74323 558860
rect 74993 558859 75059 558860
rect 76005 558859 76071 558862
rect 76782 558860 76788 558862
rect 76852 558860 76899 558864
rect 77294 558862 77340 558922
rect 77404 558920 77451 558924
rect 78438 558922 78444 558924
rect 77446 558864 77451 558920
rect 77334 558860 77340 558862
rect 77404 558860 77451 558864
rect 78398 558862 78444 558922
rect 78508 558920 78555 558924
rect 78550 558864 78555 558920
rect 78438 558860 78444 558862
rect 78508 558860 78555 558864
rect 79174 558860 79180 558924
rect 79244 558922 79250 558924
rect 79409 558922 79475 558925
rect 79961 558924 80027 558925
rect 79910 558922 79916 558924
rect 79244 558920 79475 558922
rect 79244 558864 79414 558920
rect 79470 558864 79475 558920
rect 79244 558862 79475 558864
rect 79870 558862 79916 558922
rect 79980 558920 80027 558924
rect 80022 558864 80027 558920
rect 79244 558860 79250 558862
rect 76833 558859 76899 558860
rect 77385 558859 77451 558860
rect 78489 558859 78555 558860
rect 79409 558859 79475 558862
rect 79910 558860 79916 558862
rect 79980 558860 80027 558864
rect 80646 558860 80652 558924
rect 80716 558922 80722 558924
rect 80789 558922 80855 558925
rect 81249 558924 81315 558925
rect 81198 558922 81204 558924
rect 80716 558920 80855 558922
rect 80716 558864 80794 558920
rect 80850 558864 80855 558920
rect 80716 558862 80855 558864
rect 81158 558862 81204 558922
rect 81268 558920 81315 558924
rect 81310 558864 81315 558920
rect 80716 558860 80722 558862
rect 79961 558859 80027 558860
rect 80789 558859 80855 558862
rect 81198 558860 81204 558862
rect 81268 558860 81315 558864
rect 81249 558859 81315 558860
rect 81893 558924 81959 558925
rect 82721 558924 82787 558925
rect 83825 558924 83891 558925
rect 84193 558924 84259 558925
rect 81893 558920 81940 558924
rect 82004 558922 82010 558924
rect 81893 558864 81898 558920
rect 81893 558860 81940 558864
rect 82004 558862 82050 558922
rect 82004 558860 82010 558862
rect 82670 558860 82676 558924
rect 82740 558922 82787 558924
rect 83774 558922 83780 558924
rect 82740 558920 82832 558922
rect 82782 558864 82832 558920
rect 82740 558862 82832 558864
rect 83734 558862 83780 558922
rect 83844 558920 83891 558924
rect 83886 558864 83891 558920
rect 82740 558860 82787 558862
rect 83774 558860 83780 558862
rect 83844 558860 83891 558864
rect 84142 558860 84148 558924
rect 84212 558922 84259 558924
rect 84212 558920 84304 558922
rect 84254 558864 84304 558920
rect 84212 558862 84304 558864
rect 84212 558860 84259 558862
rect 85062 558860 85068 558924
rect 85132 558922 85138 558924
rect 85481 558922 85547 558925
rect 86401 558924 86467 558925
rect 86350 558922 86356 558924
rect 85132 558920 85547 558922
rect 85132 558864 85486 558920
rect 85542 558864 85547 558920
rect 85132 558862 85547 558864
rect 86310 558862 86356 558922
rect 86420 558920 86467 558924
rect 86462 558864 86467 558920
rect 85132 558860 85138 558862
rect 81893 558859 81959 558860
rect 82721 558859 82787 558860
rect 83825 558859 83891 558860
rect 84193 558859 84259 558860
rect 85481 558859 85547 558862
rect 86350 558860 86356 558862
rect 86420 558860 86467 558864
rect 86718 558860 86724 558924
rect 86788 558922 86794 558924
rect 86861 558922 86927 558925
rect 87873 558924 87939 558925
rect 88241 558924 88307 558925
rect 87822 558922 87828 558924
rect 86788 558920 86927 558922
rect 86788 558864 86866 558920
rect 86922 558864 86927 558920
rect 86788 558862 86927 558864
rect 87782 558862 87828 558922
rect 87892 558920 87939 558924
rect 87934 558864 87939 558920
rect 86788 558860 86794 558862
rect 86401 558859 86467 558860
rect 86861 558859 86927 558862
rect 87822 558860 87828 558862
rect 87892 558860 87939 558864
rect 88190 558860 88196 558924
rect 88260 558922 88307 558924
rect 88885 558924 88951 558925
rect 88885 558922 88932 558924
rect 88260 558920 88352 558922
rect 88302 558864 88352 558920
rect 88260 558862 88352 558864
rect 88840 558920 88932 558922
rect 88840 558864 88890 558920
rect 88840 558862 88932 558864
rect 88260 558860 88307 558862
rect 87873 558859 87939 558860
rect 88241 558859 88307 558860
rect 88885 558860 88932 558862
rect 88996 558860 89002 558924
rect 89110 558860 89116 558924
rect 89180 558922 89186 558924
rect 89621 558922 89687 558925
rect 89180 558920 89687 558922
rect 89180 558864 89626 558920
rect 89682 558864 89687 558920
rect 89180 558862 89687 558864
rect 89180 558860 89186 558862
rect 88885 558859 88951 558860
rect 89621 558859 89687 558862
rect 89805 558924 89871 558925
rect 91001 558924 91067 558925
rect 92473 558924 92539 558925
rect 89805 558920 89852 558924
rect 89916 558922 89922 558924
rect 89805 558864 89810 558920
rect 89805 558860 89852 558864
rect 89916 558862 89962 558922
rect 89916 558860 89922 558862
rect 90950 558860 90956 558924
rect 91020 558922 91067 558924
rect 92422 558922 92428 558924
rect 91020 558920 91112 558922
rect 91062 558864 91112 558920
rect 91020 558862 91112 558864
rect 92382 558862 92428 558922
rect 92492 558920 92539 558924
rect 92534 558864 92539 558920
rect 91020 558860 91067 558862
rect 92422 558860 92428 558862
rect 92492 558860 92539 558864
rect 93158 558860 93164 558924
rect 93228 558922 93234 558924
rect 93669 558922 93735 558925
rect 94865 558924 94931 558925
rect 94814 558922 94820 558924
rect 93228 558920 93735 558922
rect 93228 558864 93674 558920
rect 93730 558864 93735 558920
rect 93228 558862 93735 558864
rect 94774 558862 94820 558922
rect 94884 558920 94931 558924
rect 94926 558864 94931 558920
rect 93228 558860 93234 558862
rect 89805 558859 89871 558860
rect 91001 558859 91067 558860
rect 92473 558859 92539 558860
rect 93669 558859 93735 558862
rect 94814 558860 94820 558862
rect 94884 558860 94931 558864
rect 94998 558860 95004 558924
rect 95068 558922 95074 558924
rect 95141 558922 95207 558925
rect 95785 558924 95851 558925
rect 96521 558924 96587 558925
rect 95734 558922 95740 558924
rect 95068 558920 95207 558922
rect 95068 558864 95146 558920
rect 95202 558864 95207 558920
rect 95068 558862 95207 558864
rect 95694 558862 95740 558922
rect 95804 558920 95851 558924
rect 95846 558864 95851 558920
rect 95068 558860 95074 558862
rect 94865 558859 94931 558860
rect 95141 558859 95207 558862
rect 95734 558860 95740 558862
rect 95804 558860 95851 558864
rect 96470 558860 96476 558924
rect 96540 558922 96587 558924
rect 96981 558924 97047 558925
rect 97809 558924 97875 558925
rect 96540 558920 96632 558922
rect 96582 558864 96632 558920
rect 96540 558862 96632 558864
rect 96981 558920 97028 558924
rect 97092 558922 97098 558924
rect 97758 558922 97764 558924
rect 96981 558864 96986 558920
rect 96540 558860 96587 558862
rect 95785 558859 95851 558860
rect 96521 558859 96587 558860
rect 96981 558860 97028 558864
rect 97092 558862 97138 558922
rect 97718 558862 97764 558922
rect 97828 558920 97875 558924
rect 97870 558864 97875 558920
rect 97092 558860 97098 558862
rect 97758 558860 97764 558862
rect 97828 558860 97875 558864
rect 96981 558859 97047 558860
rect 97809 558859 97875 558860
rect 98085 558924 98151 558925
rect 98085 558920 98132 558924
rect 98196 558922 98202 558924
rect 98085 558864 98090 558920
rect 98085 558860 98132 558864
rect 98196 558862 98242 558922
rect 98196 558860 98202 558862
rect 99046 558860 99052 558924
rect 99116 558922 99122 558924
rect 99281 558922 99347 558925
rect 99116 558920 99347 558922
rect 99116 558864 99286 558920
rect 99342 558864 99347 558920
rect 99116 558862 99347 558864
rect 99116 558860 99122 558862
rect 98085 558859 98151 558860
rect 99281 558859 99347 558862
rect 99557 558924 99623 558925
rect 99557 558920 99604 558924
rect 99668 558922 99674 558924
rect 99557 558864 99562 558920
rect 99557 558860 99604 558864
rect 99668 558862 99714 558922
rect 99668 558860 99674 558862
rect 100150 558860 100156 558924
rect 100220 558922 100226 558924
rect 100385 558922 100451 558925
rect 100220 558920 100451 558922
rect 100220 558864 100390 558920
rect 100446 558864 100451 558920
rect 100220 558862 100451 558864
rect 100220 558860 100226 558862
rect 99557 558859 99623 558860
rect 100385 558859 100451 558862
rect 101438 558860 101444 558924
rect 101508 558922 101514 558924
rect 102041 558922 102107 558925
rect 101508 558920 102107 558922
rect 101508 558864 102046 558920
rect 102102 558864 102107 558920
rect 101508 558862 102107 558864
rect 101508 558860 101514 558862
rect 102041 558859 102107 558862
rect 103278 558860 103284 558924
rect 103348 558922 103354 558924
rect 103421 558922 103487 558925
rect 104801 558924 104867 558925
rect 104750 558922 104756 558924
rect 103348 558920 103487 558922
rect 103348 558864 103426 558920
rect 103482 558864 103487 558920
rect 103348 558862 103487 558864
rect 104710 558862 104756 558922
rect 104820 558920 104867 558924
rect 104862 558864 104867 558920
rect 103348 558860 103354 558862
rect 103421 558859 103487 558862
rect 104750 558860 104756 558862
rect 104820 558860 104867 558864
rect 105302 558860 105308 558924
rect 105372 558922 105378 558924
rect 105537 558922 105603 558925
rect 105372 558920 105603 558922
rect 105372 558864 105542 558920
rect 105598 558864 105603 558920
rect 105372 558862 105603 558864
rect 105372 558860 105378 558862
rect 104801 558859 104867 558860
rect 105537 558859 105603 558862
rect 106038 558860 106044 558924
rect 106108 558922 106114 558924
rect 106181 558922 106247 558925
rect 106108 558920 106247 558922
rect 106108 558864 106186 558920
rect 106242 558864 106247 558920
rect 106108 558862 106247 558864
rect 106108 558860 106114 558862
rect 106181 558859 106247 558862
rect 107142 558860 107148 558924
rect 107212 558922 107218 558924
rect 107469 558922 107535 558925
rect 108481 558924 108547 558925
rect 108430 558922 108436 558924
rect 107212 558920 107535 558922
rect 107212 558864 107474 558920
rect 107530 558864 107535 558920
rect 107212 558862 107535 558864
rect 108390 558862 108436 558922
rect 108500 558920 108547 558924
rect 108542 558864 108547 558920
rect 107212 558860 107218 558862
rect 107469 558859 107535 558862
rect 108430 558860 108436 558862
rect 108500 558860 108547 558864
rect 109534 558860 109540 558924
rect 109604 558922 109610 558924
rect 110321 558922 110387 558925
rect 109604 558920 110387 558922
rect 109604 558864 110326 558920
rect 110382 558864 110387 558920
rect 109604 558862 110387 558864
rect 109604 558860 109610 558862
rect 108481 558859 108547 558860
rect 110321 558859 110387 558862
rect 195973 558922 196039 558925
rect 196198 558922 196204 558924
rect 195973 558920 196204 558922
rect 195973 558864 195978 558920
rect 196034 558864 196204 558920
rect 195973 558862 196204 558864
rect 195973 558859 196039 558862
rect 196198 558860 196204 558862
rect 196268 558860 196274 558924
rect 197353 558922 197419 558925
rect 197486 558922 197492 558924
rect 197353 558920 197492 558922
rect 197353 558864 197358 558920
rect 197414 558864 197492 558920
rect 197353 558862 197492 558864
rect 197353 558859 197419 558862
rect 197486 558860 197492 558862
rect 197556 558860 197562 558924
rect 201493 558922 201559 558925
rect 201718 558922 201724 558924
rect 201493 558920 201724 558922
rect 201493 558864 201498 558920
rect 201554 558864 201724 558920
rect 201493 558862 201724 558864
rect 201493 558859 201559 558862
rect 201718 558860 201724 558862
rect 201788 558860 201794 558924
rect 202638 558860 202644 558924
rect 202708 558922 202714 558924
rect 202781 558922 202847 558925
rect 202708 558920 202847 558922
rect 202708 558864 202786 558920
rect 202842 558864 202847 558920
rect 202708 558862 202847 558864
rect 202708 558860 202714 558862
rect 202781 558859 202847 558862
rect 203926 558860 203932 558924
rect 203996 558922 204002 558924
rect 204161 558922 204227 558925
rect 203996 558920 204227 558922
rect 203996 558864 204166 558920
rect 204222 558864 204227 558920
rect 203996 558862 204227 558864
rect 203996 558860 204002 558862
rect 204161 558859 204227 558862
rect 205398 558860 205404 558924
rect 205468 558922 205474 558924
rect 205541 558922 205607 558925
rect 205468 558920 205607 558922
rect 205468 558864 205546 558920
rect 205602 558864 205607 558920
rect 205468 558862 205607 558864
rect 205468 558860 205474 558862
rect 205541 558859 205607 558862
rect 206093 558924 206159 558925
rect 208393 558924 208459 558925
rect 210601 558924 210667 558925
rect 206093 558920 206140 558924
rect 206204 558922 206210 558924
rect 208342 558922 208348 558924
rect 206093 558864 206098 558920
rect 206093 558860 206140 558864
rect 206204 558862 206250 558922
rect 208302 558862 208348 558922
rect 208412 558920 208459 558924
rect 210550 558922 210556 558924
rect 208454 558864 208459 558920
rect 206204 558860 206210 558862
rect 208342 558860 208348 558862
rect 208412 558860 208459 558864
rect 210510 558862 210556 558922
rect 210620 558920 210667 558924
rect 210662 558864 210667 558920
rect 210550 558860 210556 558862
rect 210620 558860 210667 558864
rect 206093 558859 206159 558860
rect 208393 558859 208459 558860
rect 210601 558859 210667 558860
rect 211797 558924 211863 558925
rect 213085 558924 213151 558925
rect 211797 558920 211844 558924
rect 211908 558922 211914 558924
rect 211797 558864 211802 558920
rect 211797 558860 211844 558864
rect 211908 558862 211954 558922
rect 213085 558920 213132 558924
rect 213196 558922 213202 558924
rect 213913 558922 213979 558925
rect 215293 558924 215359 558925
rect 214046 558922 214052 558924
rect 213085 558864 213090 558920
rect 211908 558860 211914 558862
rect 213085 558860 213132 558864
rect 213196 558862 213242 558922
rect 213913 558920 214052 558922
rect 213913 558864 213918 558920
rect 213974 558864 214052 558920
rect 213913 558862 214052 558864
rect 213196 558860 213202 558862
rect 211797 558859 211863 558860
rect 213085 558859 213151 558860
rect 213913 558859 213979 558862
rect 214046 558860 214052 558862
rect 214116 558860 214122 558924
rect 215293 558920 215340 558924
rect 215404 558922 215410 558924
rect 215293 558864 215298 558920
rect 215293 558860 215340 558864
rect 215404 558862 215450 558922
rect 215404 558860 215410 558862
rect 217542 558860 217548 558924
rect 217612 558922 217618 558924
rect 217961 558922 218027 558925
rect 217612 558920 218027 558922
rect 217612 558864 217966 558920
rect 218022 558864 218027 558920
rect 217612 558862 218027 558864
rect 217612 558860 217618 558862
rect 215293 558859 215359 558860
rect 217961 558859 218027 558862
rect 218830 558860 218836 558924
rect 218900 558922 218906 558924
rect 218973 558922 219039 558925
rect 222377 558924 222443 558925
rect 222326 558922 222332 558924
rect 218900 558920 219039 558922
rect 218900 558864 218978 558920
rect 219034 558864 219039 558920
rect 218900 558862 219039 558864
rect 222286 558862 222332 558922
rect 222396 558920 222443 558924
rect 222438 558864 222443 558920
rect 218900 558860 218906 558862
rect 218973 558859 219039 558862
rect 222326 558860 222332 558862
rect 222396 558860 222443 558864
rect 222377 558859 222443 558860
rect 223573 558924 223639 558925
rect 224493 558924 224559 558925
rect 225873 558924 225939 558925
rect 227161 558924 227227 558925
rect 223573 558920 223620 558924
rect 223684 558922 223690 558924
rect 223573 558864 223578 558920
rect 223573 558860 223620 558864
rect 223684 558862 223730 558922
rect 224493 558920 224540 558924
rect 224604 558922 224610 558924
rect 225822 558922 225828 558924
rect 224493 558864 224498 558920
rect 223684 558860 223690 558862
rect 224493 558860 224540 558864
rect 224604 558862 224650 558922
rect 225782 558862 225828 558922
rect 225892 558920 225939 558924
rect 227110 558922 227116 558924
rect 225934 558864 225939 558920
rect 224604 558860 224610 558862
rect 225822 558860 225828 558862
rect 225892 558860 225939 558864
rect 227070 558862 227116 558922
rect 227180 558920 227227 558924
rect 227222 558864 227227 558920
rect 227110 558860 227116 558862
rect 227180 558860 227227 558864
rect 223573 558859 223639 558860
rect 224493 558859 224559 558860
rect 225873 558859 225939 558860
rect 227161 558859 227227 558860
rect 228173 558924 228239 558925
rect 229553 558924 229619 558925
rect 228173 558920 228220 558924
rect 228284 558922 228290 558924
rect 229502 558922 229508 558924
rect 228173 558864 228178 558920
rect 228173 558860 228220 558864
rect 228284 558862 228330 558922
rect 229462 558862 229508 558922
rect 229572 558920 229619 558924
rect 229614 558864 229619 558920
rect 228284 558860 228290 558862
rect 229502 558860 229508 558862
rect 229572 558860 229619 558864
rect 228173 558859 228239 558860
rect 229553 558859 229619 558860
rect 313365 558924 313431 558925
rect 313365 558920 313412 558924
rect 313476 558922 313482 558924
rect 321553 558922 321619 558925
rect 322790 558922 322796 558924
rect 313365 558864 313370 558920
rect 313365 558860 313412 558864
rect 313476 558862 313522 558922
rect 321553 558920 322796 558922
rect 321553 558864 321558 558920
rect 321614 558864 322796 558920
rect 321553 558862 322796 558864
rect 313476 558860 313482 558862
rect 313365 558859 313431 558860
rect 321553 558859 321619 558862
rect 322790 558860 322796 558862
rect 322860 558860 322866 558924
rect 322933 558922 322999 558925
rect 324078 558922 324084 558924
rect 322933 558920 324084 558922
rect 322933 558864 322938 558920
rect 322994 558864 324084 558920
rect 322933 558862 324084 558864
rect 322933 558859 322999 558862
rect 324078 558860 324084 558862
rect 324148 558860 324154 558924
rect 324313 558922 324379 558925
rect 325182 558922 325188 558924
rect 324313 558920 325188 558922
rect 324313 558864 324318 558920
rect 324374 558864 325188 558920
rect 324313 558862 325188 558864
rect 324313 558859 324379 558862
rect 325182 558860 325188 558862
rect 325252 558860 325258 558924
rect 325693 558922 325759 558925
rect 326286 558922 326292 558924
rect 325693 558920 326292 558922
rect 325693 558864 325698 558920
rect 325754 558864 326292 558920
rect 325693 558862 326292 558864
rect 325693 558859 325759 558862
rect 326286 558860 326292 558862
rect 326356 558860 326362 558924
rect 327073 558922 327139 558925
rect 327574 558922 327580 558924
rect 327073 558920 327580 558922
rect 327073 558864 327078 558920
rect 327134 558864 327580 558920
rect 327073 558862 327580 558864
rect 327073 558859 327139 558862
rect 327574 558860 327580 558862
rect 327644 558860 327650 558924
rect 329281 558922 329347 558925
rect 329833 558924 329899 558925
rect 329598 558922 329604 558924
rect 329281 558920 329604 558922
rect 329281 558864 329286 558920
rect 329342 558864 329604 558920
rect 329281 558862 329604 558864
rect 329281 558859 329347 558862
rect 329598 558860 329604 558862
rect 329668 558860 329674 558924
rect 329782 558860 329788 558924
rect 329852 558922 329899 558924
rect 330477 558924 330543 558925
rect 329852 558920 329944 558922
rect 329894 558864 329944 558920
rect 329852 558862 329944 558864
rect 330477 558920 330524 558924
rect 330588 558922 330594 558924
rect 331213 558922 331279 558925
rect 332358 558922 332364 558924
rect 330477 558864 330482 558920
rect 329852 558860 329899 558862
rect 329833 558859 329899 558860
rect 330477 558860 330524 558864
rect 330588 558862 330634 558922
rect 331213 558920 332364 558922
rect 331213 558864 331218 558920
rect 331274 558864 332364 558920
rect 331213 558862 332364 558864
rect 330588 558860 330594 558862
rect 330477 558859 330543 558860
rect 331213 558859 331279 558862
rect 332358 558860 332364 558862
rect 332428 558860 332434 558924
rect 332593 558922 332659 558925
rect 333278 558922 333284 558924
rect 332593 558920 333284 558922
rect 332593 558864 332598 558920
rect 332654 558864 333284 558920
rect 332593 558862 333284 558864
rect 332593 558859 332659 558862
rect 333278 558860 333284 558862
rect 333348 558860 333354 558924
rect 333973 558922 334039 558925
rect 334566 558922 334572 558924
rect 333973 558920 334572 558922
rect 333973 558864 333978 558920
rect 334034 558864 334572 558920
rect 333973 558862 334572 558864
rect 333973 558859 334039 558862
rect 334566 558860 334572 558862
rect 334636 558860 334642 558924
rect 335353 558922 335419 558925
rect 336733 558924 336799 558925
rect 335854 558922 335860 558924
rect 335353 558920 335860 558922
rect 335353 558864 335358 558920
rect 335414 558864 335860 558920
rect 335353 558862 335860 558864
rect 335353 558859 335419 558862
rect 335854 558860 335860 558862
rect 335924 558860 335930 558924
rect 336733 558922 336780 558924
rect 336688 558920 336780 558922
rect 336688 558864 336738 558920
rect 336688 558862 336780 558864
rect 336733 558860 336780 558862
rect 336844 558860 336850 558924
rect 338113 558922 338179 558925
rect 339166 558922 339172 558924
rect 338113 558920 339172 558922
rect 338113 558864 338118 558920
rect 338174 558864 339172 558920
rect 338113 558862 339172 558864
rect 336733 558859 336799 558860
rect 338113 558859 338179 558862
rect 339166 558860 339172 558862
rect 339236 558860 339242 558924
rect 339493 558922 339559 558925
rect 341241 558924 341307 558925
rect 342529 558924 342595 558925
rect 343633 558924 343699 558925
rect 340454 558922 340460 558924
rect 339493 558920 340460 558922
rect 339493 558864 339498 558920
rect 339554 558864 340460 558920
rect 339493 558862 340460 558864
rect 339493 558859 339559 558862
rect 340454 558860 340460 558862
rect 340524 558860 340530 558924
rect 341190 558922 341196 558924
rect 341150 558862 341196 558922
rect 341260 558920 341307 558924
rect 342478 558922 342484 558924
rect 341302 558864 341307 558920
rect 341190 558860 341196 558862
rect 341260 558860 341307 558864
rect 342438 558862 342484 558922
rect 342548 558920 342595 558924
rect 343582 558922 343588 558924
rect 342590 558864 342595 558920
rect 342478 558860 342484 558862
rect 342548 558860 342595 558864
rect 343542 558862 343588 558922
rect 343652 558920 343699 558924
rect 343694 558864 343699 558920
rect 343582 558860 343588 558862
rect 343652 558860 343699 558864
rect 344686 558860 344692 558924
rect 344756 558922 344762 558924
rect 344829 558922 344895 558925
rect 344756 558920 344895 558922
rect 344756 558864 344834 558920
rect 344890 558864 344895 558920
rect 344756 558862 344895 558864
rect 344756 558860 344762 558862
rect 341241 558859 341307 558860
rect 342529 558859 342595 558860
rect 343633 558859 343699 558860
rect 344829 558859 344895 558862
rect 345749 558924 345815 558925
rect 346853 558924 346919 558925
rect 348233 558924 348299 558925
rect 349521 558924 349587 558925
rect 345749 558920 345796 558924
rect 345860 558922 345866 558924
rect 345749 558864 345754 558920
rect 345749 558860 345796 558864
rect 345860 558862 345906 558922
rect 346853 558920 346900 558924
rect 346964 558922 346970 558924
rect 348182 558922 348188 558924
rect 346853 558864 346858 558920
rect 345860 558860 345866 558862
rect 346853 558860 346900 558864
rect 346964 558862 347010 558922
rect 348142 558862 348188 558922
rect 348252 558920 348299 558924
rect 349470 558922 349476 558924
rect 348294 558864 348299 558920
rect 346964 558860 346970 558862
rect 348182 558860 348188 558862
rect 348252 558860 348299 558864
rect 349430 558862 349476 558922
rect 349540 558920 349587 558924
rect 349582 558864 349587 558920
rect 349470 558860 349476 558862
rect 349540 558860 349587 558864
rect 345749 558859 345815 558860
rect 346853 558859 346919 558860
rect 348233 558859 348299 558860
rect 349521 558859 349587 558860
rect 351729 558922 351795 558925
rect 358854 558922 358860 558924
rect 351729 558920 358860 558922
rect 351729 558864 351734 558920
rect 351790 558864 358860 558920
rect 351729 558862 358860 558864
rect 351729 558859 351795 558862
rect 358854 558860 358860 558862
rect 358924 558860 358930 558924
rect 194409 558788 194475 558789
rect 64270 558724 64276 558788
rect 64340 558786 64346 558788
rect 194358 558786 194364 558788
rect 64340 558726 194364 558786
rect 194428 558784 194475 558788
rect 194470 558728 194475 558784
rect 64340 558724 64346 558726
rect 194358 558724 194364 558726
rect 194428 558724 194475 558728
rect 194409 558723 194475 558724
rect 203517 558786 203583 558789
rect 203742 558786 203748 558788
rect 203517 558784 203748 558786
rect 203517 558728 203522 558784
rect 203578 558728 203748 558784
rect 203517 558726 203748 558728
rect 203517 558723 203583 558726
rect 203742 558724 203748 558726
rect 203812 558724 203818 558788
rect 216622 558724 216628 558788
rect 216692 558786 216698 558788
rect 217777 558786 217843 558789
rect 216692 558784 217843 558786
rect 216692 558728 217782 558784
rect 217838 558728 217843 558784
rect 216692 558726 217843 558728
rect 216692 558724 216698 558726
rect 217777 558723 217843 558726
rect 231853 558786 231919 558789
rect 232814 558786 232820 558788
rect 231853 558784 232820 558786
rect 231853 558728 231858 558784
rect 231914 558728 232820 558784
rect 231853 558726 232820 558728
rect 231853 558723 231919 558726
rect 232814 558724 232820 558726
rect 232884 558724 232890 558788
rect 233233 558786 233299 558789
rect 322197 558788 322263 558789
rect 323577 558788 323643 558789
rect 233550 558786 233556 558788
rect 233233 558784 233556 558786
rect 233233 558728 233238 558784
rect 233294 558728 233556 558784
rect 233233 558726 233556 558728
rect 233233 558723 233299 558726
rect 233550 558724 233556 558726
rect 233620 558724 233626 558788
rect 322197 558786 322244 558788
rect 322152 558784 322244 558786
rect 322152 558728 322202 558784
rect 322152 558726 322244 558728
rect 322197 558724 322244 558726
rect 322308 558724 322314 558788
rect 323526 558724 323532 558788
rect 323596 558786 323643 558788
rect 323596 558784 323688 558786
rect 323638 558728 323688 558784
rect 323596 558726 323688 558728
rect 323596 558724 323643 558726
rect 324814 558724 324820 558788
rect 324884 558786 324890 558788
rect 324957 558786 325023 558789
rect 324884 558784 325023 558786
rect 324884 558728 324962 558784
rect 325018 558728 325023 558784
rect 324884 558726 325023 558728
rect 324884 558724 324890 558726
rect 322197 558723 322263 558724
rect 323577 558723 323643 558724
rect 324957 558723 325023 558726
rect 326102 558724 326108 558788
rect 326172 558786 326178 558788
rect 326337 558786 326403 558789
rect 326172 558784 326403 558786
rect 326172 558728 326342 558784
rect 326398 558728 326403 558784
rect 326172 558726 326403 558728
rect 326172 558724 326178 558726
rect 326337 558723 326403 558726
rect 327022 558724 327028 558788
rect 327092 558786 327098 558788
rect 327717 558786 327783 558789
rect 327092 558784 327783 558786
rect 327092 558728 327722 558784
rect 327778 558728 327783 558784
rect 327092 558726 327783 558728
rect 327092 558724 327098 558726
rect 327717 558723 327783 558726
rect 328453 558784 328519 558789
rect 328453 558728 328458 558784
rect 328514 558728 328519 558784
rect 328453 558723 328519 558728
rect 329925 558786 329991 558789
rect 331765 558788 331831 558789
rect 332685 558788 332751 558789
rect 334065 558788 334131 558789
rect 331070 558786 331076 558788
rect 329925 558784 331076 558786
rect 329925 558728 329930 558784
rect 329986 558728 331076 558784
rect 329925 558726 331076 558728
rect 329925 558723 329991 558726
rect 331070 558724 331076 558726
rect 331140 558724 331146 558788
rect 331765 558784 331812 558788
rect 331876 558786 331882 558788
rect 331765 558728 331770 558784
rect 331765 558724 331812 558728
rect 331876 558726 331922 558786
rect 332685 558784 332732 558788
rect 332796 558786 332802 558788
rect 334014 558786 334020 558788
rect 332685 558728 332690 558784
rect 331876 558724 331882 558726
rect 332685 558724 332732 558728
rect 332796 558726 332842 558786
rect 333974 558726 334020 558786
rect 334084 558784 334131 558788
rect 334126 558728 334131 558784
rect 332796 558724 332802 558726
rect 334014 558724 334020 558726
rect 334084 558724 334131 558728
rect 331765 558723 331831 558724
rect 332685 558723 332751 558724
rect 334065 558723 334131 558724
rect 335445 558788 335511 558789
rect 335445 558784 335492 558788
rect 335556 558786 335562 558788
rect 336457 558786 336523 558789
rect 336590 558786 336596 558788
rect 335445 558728 335450 558784
rect 335445 558724 335492 558728
rect 335556 558726 335602 558786
rect 336457 558784 336596 558786
rect 336457 558728 336462 558784
rect 336518 558728 336596 558784
rect 336457 558726 336596 558728
rect 335556 558724 335562 558726
rect 335445 558723 335511 558724
rect 336457 558723 336523 558726
rect 336590 558724 336596 558726
rect 336660 558724 336666 558788
rect 338021 558784 338087 558789
rect 339033 558788 339099 558789
rect 338982 558786 338988 558788
rect 338021 558728 338026 558784
rect 338082 558728 338087 558784
rect 338021 558723 338087 558728
rect 338942 558726 338988 558786
rect 339052 558784 339099 558788
rect 339094 558728 339099 558784
rect 338982 558724 338988 558726
rect 339052 558724 339099 558728
rect 339033 558723 339099 558724
rect 339861 558788 339927 558789
rect 339861 558784 339908 558788
rect 339972 558786 339978 558788
rect 353293 558786 353359 558789
rect 353518 558786 353524 558788
rect 339861 558728 339866 558784
rect 339861 558724 339908 558728
rect 339972 558726 340018 558786
rect 353293 558784 353524 558786
rect 353293 558728 353298 558784
rect 353354 558728 353524 558784
rect 353293 558726 353524 558728
rect 339972 558724 339978 558726
rect 339861 558723 339927 558724
rect 353293 558723 353359 558726
rect 353518 558724 353524 558726
rect 353588 558724 353594 558788
rect 354673 558786 354739 558789
rect 356053 558788 356119 558789
rect 354806 558786 354812 558788
rect 354673 558784 354812 558786
rect 354673 558728 354678 558784
rect 354734 558728 354812 558784
rect 354673 558726 354812 558728
rect 354673 558723 354739 558726
rect 354806 558724 354812 558726
rect 354876 558724 354882 558788
rect 356053 558786 356100 558788
rect 356008 558784 356100 558786
rect 356008 558728 356058 558784
rect 356008 558726 356100 558728
rect 356053 558724 356100 558726
rect 356164 558724 356170 558788
rect 356053 558723 356119 558724
rect 69790 558588 69796 558652
rect 69860 558650 69866 558652
rect 70209 558650 70275 558653
rect 69860 558648 70275 558650
rect 69860 558592 70214 558648
rect 70270 558592 70275 558648
rect 69860 558590 70275 558592
rect 69860 558588 69866 558590
rect 70209 558587 70275 558590
rect 79358 558588 79364 558652
rect 79428 558650 79434 558652
rect 79593 558650 79659 558653
rect 79428 558648 79659 558650
rect 79428 558592 79598 558648
rect 79654 558592 79659 558648
rect 79428 558590 79659 558592
rect 79428 558588 79434 558590
rect 79593 558587 79659 558590
rect 82813 558652 82879 558653
rect 82813 558648 82860 558652
rect 82924 558650 82930 558652
rect 85205 558650 85271 558653
rect 85430 558650 85436 558652
rect 82813 558592 82818 558648
rect 82813 558588 82860 558592
rect 82924 558590 82970 558650
rect 85205 558648 85436 558650
rect 85205 558592 85210 558648
rect 85266 558592 85436 558648
rect 85205 558590 85436 558592
rect 82924 558588 82930 558590
rect 82813 558587 82879 558588
rect 85205 558587 85271 558590
rect 85430 558588 85436 558590
rect 85500 558588 85506 558652
rect 86166 558588 86172 558652
rect 86236 558650 86242 558652
rect 86769 558650 86835 558653
rect 86236 558648 86835 558650
rect 86236 558592 86774 558648
rect 86830 558592 86835 558648
rect 86236 558590 86835 558592
rect 86236 558588 86242 558590
rect 86769 558587 86835 558590
rect 91093 558652 91159 558653
rect 93301 558652 93367 558653
rect 93761 558652 93827 558653
rect 91093 558648 91140 558652
rect 91204 558650 91210 558652
rect 91093 558592 91098 558648
rect 91093 558588 91140 558592
rect 91204 558590 91250 558650
rect 93301 558648 93348 558652
rect 93412 558650 93418 558652
rect 93710 558650 93716 558652
rect 93301 558592 93306 558648
rect 91204 558588 91210 558590
rect 93301 558588 93348 558592
rect 93412 558590 93458 558650
rect 93670 558590 93716 558650
rect 93780 558648 93827 558652
rect 93822 558592 93827 558648
rect 93412 558588 93418 558590
rect 93710 558588 93716 558590
rect 93780 558588 93827 558592
rect 91093 558587 91159 558588
rect 93301 558587 93367 558588
rect 93761 558587 93827 558588
rect 100017 558650 100083 558653
rect 101949 558652 102015 558653
rect 102777 558652 102843 558653
rect 100334 558650 100340 558652
rect 100017 558648 100340 558650
rect 100017 558592 100022 558648
rect 100078 558592 100340 558648
rect 100017 558590 100340 558592
rect 100017 558587 100083 558590
rect 100334 558588 100340 558590
rect 100404 558588 100410 558652
rect 101949 558648 101996 558652
rect 102060 558650 102066 558652
rect 101949 558592 101954 558648
rect 101949 558588 101996 558592
rect 102060 558590 102106 558650
rect 102060 558588 102066 558590
rect 102726 558588 102732 558652
rect 102796 558650 102843 558652
rect 103881 558650 103947 558653
rect 104014 558650 104020 558652
rect 102796 558648 102888 558650
rect 102838 558592 102888 558648
rect 102796 558590 102888 558592
rect 103881 558648 104020 558650
rect 103881 558592 103886 558648
rect 103942 558592 104020 558648
rect 103881 558590 104020 558592
rect 102796 558588 102843 558590
rect 101949 558587 102015 558588
rect 102777 558587 102843 558588
rect 103881 558587 103947 558590
rect 104014 558588 104020 558590
rect 104084 558588 104090 558652
rect 106222 558588 106228 558652
rect 106292 558650 106298 558652
rect 106917 558650 106983 558653
rect 107745 558652 107811 558653
rect 107694 558650 107700 558652
rect 106292 558648 106983 558650
rect 106292 558592 106922 558648
rect 106978 558592 106983 558648
rect 106292 558590 106983 558592
rect 107654 558590 107700 558650
rect 107764 558648 107811 558652
rect 107806 558592 107811 558648
rect 106292 558588 106298 558590
rect 106917 558587 106983 558590
rect 107694 558588 107700 558590
rect 107764 558588 107811 558592
rect 107745 558587 107811 558588
rect 108297 558650 108363 558653
rect 108614 558650 108620 558652
rect 108297 558648 108620 558650
rect 108297 558592 108302 558648
rect 108358 558592 108620 558648
rect 108297 558590 108620 558592
rect 108297 558587 108363 558590
rect 108614 558588 108620 558590
rect 108684 558588 108690 558652
rect 202137 558650 202203 558653
rect 204897 558652 204963 558653
rect 202454 558650 202460 558652
rect 202137 558648 202460 558650
rect 202137 558592 202142 558648
rect 202198 558592 202460 558648
rect 202137 558590 202460 558592
rect 202137 558587 202203 558590
rect 202454 558588 202460 558590
rect 202524 558588 202530 558652
rect 204846 558650 204852 558652
rect 204806 558590 204852 558650
rect 204916 558648 204963 558652
rect 204958 558592 204963 558648
rect 204846 558588 204852 558590
rect 204916 558588 204963 558592
rect 204897 558587 204963 558588
rect 209037 558650 209103 558653
rect 209630 558650 209636 558652
rect 209037 558648 209636 558650
rect 209037 558592 209042 558648
rect 209098 558592 209636 558648
rect 209037 558590 209636 558592
rect 209037 558587 209103 558590
rect 209630 558588 209636 558590
rect 209700 558588 209706 558652
rect 234889 558650 234955 558653
rect 237373 558652 237439 558653
rect 235022 558650 235028 558652
rect 234889 558648 235028 558650
rect 234889 558592 234894 558648
rect 234950 558592 235028 558648
rect 234889 558590 235028 558592
rect 234889 558587 234955 558590
rect 235022 558588 235028 558590
rect 235092 558588 235098 558652
rect 237373 558650 237420 558652
rect 237328 558648 237420 558650
rect 237328 558592 237378 558648
rect 237328 558590 237420 558592
rect 237373 558588 237420 558590
rect 237484 558588 237490 558652
rect 282310 558588 282316 558652
rect 282380 558650 282386 558652
rect 328456 558650 328516 558723
rect 282380 558590 328516 558650
rect 338024 558650 338084 558723
rect 348049 558650 348115 558653
rect 357934 558650 357940 558652
rect 338024 558648 348115 558650
rect 338024 558592 348054 558648
rect 348110 558592 348115 558648
rect 338024 558590 348115 558592
rect 282380 558588 282386 558590
rect 237373 558587 237439 558588
rect 348049 558587 348115 558590
rect 352238 558590 357940 558650
rect 231945 558514 232011 558517
rect 238753 558516 238819 558517
rect 236126 558514 236132 558516
rect 231945 558512 236132 558514
rect 231945 558456 231950 558512
rect 232006 558456 236132 558512
rect 231945 558454 236132 558456
rect 231945 558451 232011 558454
rect 236126 558452 236132 558454
rect 236196 558452 236202 558516
rect 238702 558452 238708 558516
rect 238772 558514 238819 558516
rect 238772 558512 238864 558514
rect 238814 558456 238864 558512
rect 238772 558454 238864 558456
rect 238772 558452 238819 558454
rect 283414 558452 283420 558516
rect 283484 558514 283490 558516
rect 328453 558514 328519 558517
rect 283484 558512 328519 558514
rect 283484 558456 328458 558512
rect 328514 558456 328519 558512
rect 283484 558454 328519 558456
rect 283484 558452 283490 558454
rect 238753 558451 238819 558452
rect 328453 558451 328519 558454
rect 338021 558514 338087 558517
rect 345657 558514 345723 558517
rect 338021 558512 345723 558514
rect 338021 558456 338026 558512
rect 338082 558456 345662 558512
rect 345718 558456 345723 558512
rect 338021 558454 345723 558456
rect 338021 558451 338087 558454
rect 345657 558451 345723 558454
rect 350533 558516 350599 558517
rect 350533 558512 350580 558516
rect 350644 558514 350650 558516
rect 352238 558514 352298 558590
rect 357934 558588 357940 558590
rect 358004 558588 358010 558652
rect 350533 558456 350538 558512
rect 350533 558452 350580 558456
rect 350644 558454 350690 558514
rect 351686 558454 352298 558514
rect 357433 558514 357499 558517
rect 357566 558514 357572 558516
rect 357433 558512 357572 558514
rect 357433 558456 357438 558512
rect 357494 558456 357572 558512
rect 357433 558454 357572 558456
rect 350644 558452 350650 558454
rect 350533 558451 350599 558452
rect 78070 558316 78076 558380
rect 78140 558378 78146 558380
rect 78581 558378 78647 558381
rect 78140 558376 78647 558378
rect 78140 558320 78586 558376
rect 78642 558320 78647 558376
rect 78140 558318 78647 558320
rect 78140 558316 78146 558318
rect 78581 558315 78647 558318
rect 92054 558316 92060 558380
rect 92124 558378 92130 558380
rect 92381 558378 92447 558381
rect 92124 558376 92447 558378
rect 92124 558320 92386 558376
rect 92442 558320 92447 558376
rect 92124 558318 92447 558320
rect 92124 558316 92130 558318
rect 92381 558315 92447 558318
rect 97993 558378 98059 558381
rect 101397 558378 101463 558381
rect 101622 558378 101628 558380
rect 97993 558376 101628 558378
rect 97993 558320 97998 558376
rect 98054 558320 101402 558376
rect 101458 558320 101628 558376
rect 97993 558318 101628 558320
rect 97993 558315 98059 558318
rect 101397 558315 101463 558318
rect 101622 558316 101628 558318
rect 101692 558316 101698 558380
rect 215109 558378 215175 558381
rect 221038 558378 221044 558380
rect 215109 558376 221044 558378
rect 215109 558320 215114 558376
rect 215170 558320 221044 558376
rect 215109 558318 221044 558320
rect 215109 558315 215175 558318
rect 221038 558316 221044 558318
rect 221108 558378 221114 558380
rect 221549 558378 221615 558381
rect 221108 558376 221615 558378
rect 221108 558320 221554 558376
rect 221610 558320 221615 558376
rect 221108 558318 221615 558320
rect 221108 558316 221114 558318
rect 221549 558315 221615 558318
rect 230473 558378 230539 558381
rect 231853 558380 231919 558381
rect 230606 558378 230612 558380
rect 230473 558376 230612 558378
rect 230473 558320 230478 558376
rect 230534 558320 230612 558376
rect 230473 558318 230612 558320
rect 230473 558315 230539 558318
rect 230606 558316 230612 558318
rect 230676 558316 230682 558380
rect 231853 558378 231900 558380
rect 231808 558376 231900 558378
rect 231808 558320 231858 558376
rect 231808 558318 231900 558320
rect 231853 558316 231900 558318
rect 231964 558316 231970 558380
rect 283782 558316 283788 558380
rect 283852 558378 283858 558380
rect 351686 558378 351746 558454
rect 357433 558451 357499 558454
rect 357566 558452 357572 558454
rect 357636 558452 357642 558516
rect 283852 558318 351746 558378
rect 283852 558316 283858 558318
rect 231853 558315 231919 558316
rect 75678 558180 75684 558244
rect 75748 558242 75754 558244
rect 75821 558242 75887 558245
rect 75748 558240 75887 558242
rect 75748 558184 75826 558240
rect 75882 558184 75887 558240
rect 75748 558182 75887 558184
rect 75748 558180 75754 558182
rect 75821 558179 75887 558182
rect 283598 558180 283604 558244
rect 283668 558242 283674 558244
rect 351729 558242 351795 558245
rect 283668 558240 351795 558242
rect 283668 558184 351734 558240
rect 351790 558184 351795 558240
rect 283668 558182 351795 558184
rect 283668 558180 283674 558182
rect 351729 558179 351795 558182
rect 351913 558242 351979 558245
rect 352414 558242 352420 558244
rect 351913 558240 352420 558242
rect 351913 558184 351918 558240
rect 351974 558184 352420 558240
rect 351913 558182 352420 558184
rect 351913 558179 351979 558182
rect 352414 558180 352420 558182
rect 352484 558180 352490 558244
rect 354673 558242 354739 558245
rect 355726 558242 355732 558244
rect 354673 558240 355732 558242
rect 354673 558184 354678 558240
rect 354734 558184 355732 558240
rect 354673 558182 355732 558184
rect 354673 558179 354739 558182
rect 355726 558180 355732 558182
rect 355796 558180 355802 558244
rect 345657 558106 345723 558109
rect 351913 558106 351979 558109
rect 353150 558106 353156 558108
rect 345657 558104 351746 558106
rect 345657 558048 345662 558104
rect 345718 558048 351746 558104
rect 345657 558046 351746 558048
rect 345657 558043 345723 558046
rect 317413 557972 317479 557973
rect 317413 557970 317460 557972
rect 317368 557968 317460 557970
rect 317368 557912 317418 557968
rect 317368 557910 317460 557912
rect 317413 557908 317460 557910
rect 317524 557908 317530 557972
rect 320173 557970 320239 557973
rect 320582 557970 320588 557972
rect 320173 557968 320588 557970
rect 320173 557912 320178 557968
rect 320234 557912 320588 557968
rect 320173 557910 320588 557912
rect 317413 557907 317479 557908
rect 320173 557907 320239 557910
rect 320582 557908 320588 557910
rect 320652 557908 320658 557972
rect 336825 557970 336891 557973
rect 337878 557970 337884 557972
rect 336825 557968 337884 557970
rect 336825 557912 336830 557968
rect 336886 557912 337884 557968
rect 336825 557910 337884 557912
rect 336825 557907 336891 557910
rect 337878 557908 337884 557910
rect 337948 557908 337954 557972
rect 200205 557836 200271 557837
rect 200205 557834 200252 557836
rect 200160 557832 200252 557834
rect 200160 557776 200210 557832
rect 200160 557774 200252 557776
rect 200205 557772 200252 557774
rect 200316 557772 200322 557836
rect 229093 557834 229159 557837
rect 238661 557834 238727 557837
rect 229093 557832 238727 557834
rect 229093 557776 229098 557832
rect 229154 557776 238666 557832
rect 238722 557776 238727 557832
rect 229093 557774 238727 557776
rect 200205 557771 200271 557772
rect 229093 557771 229159 557774
rect 238661 557771 238727 557774
rect 198733 557700 198799 557701
rect 198733 557698 198780 557700
rect 198688 557696 198780 557698
rect 198688 557640 198738 557696
rect 198688 557638 198780 557640
rect 198733 557636 198780 557638
rect 198844 557636 198850 557700
rect 207054 557636 207060 557700
rect 207124 557698 207130 557700
rect 207657 557698 207723 557701
rect 207124 557696 207723 557698
rect 207124 557640 207662 557696
rect 207718 557640 207723 557696
rect 207124 557638 207723 557640
rect 207124 557636 207130 557638
rect 198733 557635 198799 557636
rect 207657 557635 207723 557638
rect 210366 557636 210372 557700
rect 210436 557698 210442 557700
rect 211061 557698 211127 557701
rect 210436 557696 211127 557698
rect 210436 557640 211066 557696
rect 211122 557640 211127 557696
rect 210436 557638 211127 557640
rect 210436 557636 210442 557638
rect 211061 557635 211127 557638
rect 217358 557636 217364 557700
rect 217428 557698 217434 557700
rect 217869 557698 217935 557701
rect 217428 557696 217935 557698
rect 217428 557640 217874 557696
rect 217930 557640 217935 557696
rect 217428 557638 217935 557640
rect 217428 557636 217434 557638
rect 217869 557635 217935 557638
rect 225638 557636 225644 557700
rect 225708 557698 225714 557700
rect 226149 557698 226215 557701
rect 225708 557696 226215 557698
rect 225708 557640 226154 557696
rect 226210 557640 226215 557696
rect 225708 557638 226215 557640
rect 225708 557636 225714 557638
rect 226149 557635 226215 557638
rect 232630 557636 232636 557700
rect 232700 557698 232706 557700
rect 233141 557698 233207 557701
rect 232700 557696 233207 557698
rect 232700 557640 233146 557696
rect 233202 557640 233207 557696
rect 232700 557638 233207 557640
rect 232700 557636 232706 557638
rect 233141 557635 233207 557638
rect 343725 557698 343791 557701
rect 344870 557698 344876 557700
rect 343725 557696 344876 557698
rect 343725 557640 343730 557696
rect 343786 557640 344876 557696
rect 343725 557638 344876 557640
rect 343725 557635 343791 557638
rect 344870 557636 344876 557638
rect 344940 557636 344946 557700
rect 351686 557698 351746 558046
rect 351913 558104 353156 558106
rect 351913 558048 351918 558104
rect 351974 558048 353156 558104
rect 351913 558046 353156 558048
rect 351913 558043 351979 558046
rect 353150 558044 353156 558046
rect 353220 558044 353226 558108
rect 353293 557970 353359 557973
rect 354438 557970 354444 557972
rect 353293 557968 354444 557970
rect 353293 557912 353298 557968
rect 353354 557912 354444 557968
rect 353293 557910 354444 557912
rect 353293 557907 353359 557910
rect 354438 557908 354444 557910
rect 354508 557908 354514 557972
rect 356646 557698 356652 557700
rect 351686 557638 356652 557698
rect 356646 557636 356652 557638
rect 356716 557636 356722 557700
rect 206921 557564 206987 557565
rect 206870 557500 206876 557564
rect 206940 557562 206987 557564
rect 206940 557560 207032 557562
rect 206982 557504 207032 557560
rect 206940 557502 207032 557504
rect 206940 557500 206987 557502
rect 207974 557500 207980 557564
rect 208044 557562 208050 557564
rect 208301 557562 208367 557565
rect 208044 557560 208367 557562
rect 208044 557504 208306 557560
rect 208362 557504 208367 557560
rect 208044 557502 208367 557504
rect 208044 557500 208050 557502
rect 206921 557499 206987 557500
rect 208301 557499 208367 557502
rect 209262 557500 209268 557564
rect 209332 557562 209338 557564
rect 209681 557562 209747 557565
rect 212441 557564 212507 557565
rect 209332 557560 209747 557562
rect 209332 557504 209686 557560
rect 209742 557504 209747 557560
rect 209332 557502 209747 557504
rect 209332 557500 209338 557502
rect 209681 557499 209747 557502
rect 212390 557500 212396 557564
rect 212460 557562 212507 557564
rect 212460 557560 212552 557562
rect 212502 557504 212552 557560
rect 212460 557502 212552 557504
rect 212460 557500 212507 557502
rect 213494 557500 213500 557564
rect 213564 557562 213570 557564
rect 213821 557562 213887 557565
rect 213564 557560 213887 557562
rect 213564 557504 213826 557560
rect 213882 557504 213887 557560
rect 213564 557502 213887 557504
rect 213564 557500 213570 557502
rect 212441 557499 212507 557500
rect 213821 557499 213887 557502
rect 214782 557500 214788 557564
rect 214852 557562 214858 557564
rect 215201 557562 215267 557565
rect 214852 557560 215267 557562
rect 214852 557504 215206 557560
rect 215262 557504 215267 557560
rect 214852 557502 215267 557504
rect 214852 557500 214858 557502
rect 215201 557499 215267 557502
rect 216254 557500 216260 557564
rect 216324 557562 216330 557564
rect 216581 557562 216647 557565
rect 217961 557564 218027 557565
rect 216324 557560 216647 557562
rect 216324 557504 216586 557560
rect 216642 557504 216647 557560
rect 216324 557502 216647 557504
rect 216324 557500 216330 557502
rect 216581 557499 216647 557502
rect 217910 557500 217916 557564
rect 217980 557562 218027 557564
rect 217980 557560 218072 557562
rect 218022 557504 218072 557560
rect 217980 557502 218072 557504
rect 217980 557500 218027 557502
rect 219198 557500 219204 557564
rect 219268 557562 219274 557564
rect 219341 557562 219407 557565
rect 220721 557564 220787 557565
rect 219268 557560 219407 557562
rect 219268 557504 219346 557560
rect 219402 557504 219407 557560
rect 219268 557502 219407 557504
rect 219268 557500 219274 557502
rect 217961 557499 218027 557500
rect 219341 557499 219407 557502
rect 220670 557500 220676 557564
rect 220740 557562 220787 557564
rect 220740 557560 220832 557562
rect 220782 557504 220832 557560
rect 220740 557502 220832 557504
rect 220740 557500 220787 557502
rect 221958 557500 221964 557564
rect 222028 557562 222034 557564
rect 222101 557562 222167 557565
rect 222028 557560 222167 557562
rect 222028 557504 222106 557560
rect 222162 557504 222167 557560
rect 222028 557502 222167 557504
rect 222028 557500 222034 557502
rect 220721 557499 220787 557500
rect 222101 557499 222167 557502
rect 223246 557500 223252 557564
rect 223316 557562 223322 557564
rect 223481 557562 223547 557565
rect 223316 557560 223547 557562
rect 223316 557504 223486 557560
rect 223542 557504 223547 557560
rect 223316 557502 223547 557504
rect 223316 557500 223322 557502
rect 223481 557499 223547 557502
rect 224350 557500 224356 557564
rect 224420 557562 224426 557564
rect 224861 557562 224927 557565
rect 226241 557564 226307 557565
rect 224420 557560 224927 557562
rect 224420 557504 224866 557560
rect 224922 557504 224927 557560
rect 224420 557502 224927 557504
rect 224420 557500 224426 557502
rect 224861 557499 224927 557502
rect 226190 557500 226196 557564
rect 226260 557562 226307 557564
rect 226260 557560 226352 557562
rect 226302 557504 226352 557560
rect 226260 557502 226352 557504
rect 226260 557500 226307 557502
rect 227478 557500 227484 557564
rect 227548 557562 227554 557564
rect 227621 557562 227687 557565
rect 227548 557560 227687 557562
rect 227548 557504 227626 557560
rect 227682 557504 227687 557560
rect 227548 557502 227687 557504
rect 227548 557500 227554 557502
rect 226241 557499 226307 557500
rect 227621 557499 227687 557502
rect 228766 557500 228772 557564
rect 228836 557562 228842 557564
rect 229001 557562 229067 557565
rect 228836 557560 229067 557562
rect 228836 557504 229006 557560
rect 229062 557504 229067 557560
rect 228836 557502 229067 557504
rect 228836 557500 228842 557502
rect 229001 557499 229067 557502
rect 230238 557500 230244 557564
rect 230308 557562 230314 557564
rect 230381 557562 230447 557565
rect 230308 557560 230447 557562
rect 230308 557504 230386 557560
rect 230442 557504 230447 557560
rect 230308 557502 230447 557504
rect 230308 557500 230314 557502
rect 230381 557499 230447 557502
rect 230790 557500 230796 557564
rect 230860 557562 230866 557564
rect 231761 557562 231827 557565
rect 233049 557564 233115 557565
rect 234521 557564 234587 557565
rect 230860 557560 231827 557562
rect 230860 557504 231766 557560
rect 231822 557504 231827 557560
rect 230860 557502 231827 557504
rect 230860 557500 230866 557502
rect 231761 557499 231827 557502
rect 232998 557500 233004 557564
rect 233068 557562 233115 557564
rect 234470 557562 234476 557564
rect 233068 557560 233160 557562
rect 233110 557504 233160 557560
rect 233068 557502 233160 557504
rect 234430 557502 234476 557562
rect 234540 557560 234587 557564
rect 234582 557504 234587 557560
rect 233068 557500 233115 557502
rect 234470 557500 234476 557502
rect 234540 557500 234587 557504
rect 235758 557500 235764 557564
rect 235828 557562 235834 557564
rect 235901 557562 235967 557565
rect 237281 557564 237347 557565
rect 235828 557560 235967 557562
rect 235828 557504 235906 557560
rect 235962 557504 235967 557560
rect 235828 557502 235967 557504
rect 235828 557500 235834 557502
rect 233049 557499 233115 557500
rect 234521 557499 234587 557500
rect 235901 557499 235967 557502
rect 237230 557500 237236 557564
rect 237300 557562 237347 557564
rect 237300 557560 237392 557562
rect 237342 557504 237392 557560
rect 237300 557502 237392 557504
rect 237300 557500 237347 557502
rect 238334 557500 238340 557564
rect 238404 557562 238410 557564
rect 238661 557562 238727 557565
rect 238404 557560 238727 557562
rect 238404 557504 238666 557560
rect 238722 557504 238727 557560
rect 238404 557502 238727 557504
rect 238404 557500 238410 557502
rect 237281 557499 237347 557500
rect 238661 557499 238727 557502
rect 239622 557500 239628 557564
rect 239692 557562 239698 557564
rect 240041 557562 240107 557565
rect 239692 557560 240107 557562
rect 239692 557504 240046 557560
rect 240102 557504 240107 557560
rect 239692 557502 240107 557504
rect 239692 557500 239698 557502
rect 240041 557499 240107 557502
rect 241605 557562 241671 557565
rect 251081 557562 251147 557565
rect 241605 557560 251147 557562
rect 241605 557504 241610 557560
rect 241666 557504 251086 557560
rect 251142 557504 251147 557560
rect 241605 557502 251147 557504
rect 241605 557499 241671 557502
rect 251081 557499 251147 557502
rect 260833 557562 260899 557565
rect 270401 557562 270467 557565
rect 260833 557560 270467 557562
rect 260833 557504 260838 557560
rect 260894 557504 270406 557560
rect 270462 557504 270467 557560
rect 260833 557502 270467 557504
rect 260833 557499 260899 557502
rect 270401 557499 270467 557502
rect 316033 557562 316099 557565
rect 316350 557562 316356 557564
rect 316033 557560 316356 557562
rect 316033 557504 316038 557560
rect 316094 557504 316356 557560
rect 316033 557502 316356 557504
rect 316033 557499 316099 557502
rect 316350 557500 316356 557502
rect 316420 557500 316426 557564
rect 318793 557562 318859 557565
rect 318926 557562 318932 557564
rect 318793 557560 318932 557562
rect 318793 557504 318798 557560
rect 318854 557504 318932 557560
rect 318793 557502 318932 557504
rect 318793 557499 318859 557502
rect 318926 557500 318932 557502
rect 318996 557500 319002 557564
rect 320265 557562 320331 557565
rect 320950 557562 320956 557564
rect 320265 557560 320956 557562
rect 320265 557504 320270 557560
rect 320326 557504 320956 557560
rect 320265 557502 320956 557504
rect 320265 557499 320331 557502
rect 320950 557500 320956 557502
rect 321020 557500 321026 557564
rect 340873 557562 340939 557565
rect 341742 557562 341748 557564
rect 340873 557560 341748 557562
rect 340873 557504 340878 557560
rect 340934 557504 341748 557560
rect 340873 557502 341748 557504
rect 340873 557499 340939 557502
rect 341742 557500 341748 557502
rect 341812 557500 341818 557564
rect 342253 557562 342319 557565
rect 342662 557562 342668 557564
rect 342253 557560 342668 557562
rect 342253 557504 342258 557560
rect 342314 557504 342668 557560
rect 342253 557502 342668 557504
rect 342253 557499 342319 557502
rect 342662 557500 342668 557502
rect 342732 557500 342738 557564
rect 343633 557562 343699 557565
rect 343950 557562 343956 557564
rect 343633 557560 343956 557562
rect 343633 557504 343638 557560
rect 343694 557504 343956 557560
rect 343633 557502 343956 557504
rect 343633 557499 343699 557502
rect 343950 557500 343956 557502
rect 344020 557500 344026 557564
rect 345013 557562 345079 557565
rect 346158 557562 346164 557564
rect 345013 557560 346164 557562
rect 345013 557504 345018 557560
rect 345074 557504 346164 557560
rect 345013 557502 346164 557504
rect 345013 557499 345079 557502
rect 346158 557500 346164 557502
rect 346228 557500 346234 557564
rect 346393 557562 346459 557565
rect 347446 557562 347452 557564
rect 346393 557560 347452 557562
rect 346393 557504 346398 557560
rect 346454 557504 347452 557560
rect 346393 557502 347452 557504
rect 346393 557499 346459 557502
rect 347446 557500 347452 557502
rect 347516 557500 347522 557564
rect 347773 557562 347839 557565
rect 348734 557562 348740 557564
rect 347773 557560 348740 557562
rect 347773 557504 347778 557560
rect 347834 557504 348740 557560
rect 347773 557502 348740 557504
rect 347773 557499 347839 557502
rect 348734 557500 348740 557502
rect 348804 557500 348810 557564
rect 349153 557562 349219 557565
rect 349654 557562 349660 557564
rect 349153 557560 349660 557562
rect 349153 557504 349158 557560
rect 349214 557504 349660 557560
rect 349153 557502 349660 557504
rect 349153 557499 349219 557502
rect 349654 557500 349660 557502
rect 349724 557500 349730 557564
rect 350625 557562 350691 557565
rect 350942 557562 350948 557564
rect 350625 557560 350948 557562
rect 350625 557504 350630 557560
rect 350686 557504 350948 557560
rect 350625 557502 350948 557504
rect 350625 557499 350691 557502
rect 350942 557500 350948 557502
rect 351012 557500 351018 557564
rect 580165 557290 580231 557293
rect 583520 557290 584960 557380
rect 580165 557288 584960 557290
rect 580165 557232 580170 557288
rect 580226 557232 584960 557288
rect 580165 557230 584960 557232
rect 580165 557227 580231 557230
rect 328453 557154 328519 557157
rect 328862 557154 328868 557156
rect 328453 557152 328868 557154
rect 328453 557096 328458 557152
rect 328514 557096 328868 557152
rect 328453 557094 328868 557096
rect 328453 557091 328519 557094
rect 328862 557092 328868 557094
rect 328932 557092 328938 557156
rect 583520 557140 584960 557230
rect -960 553074 480 553164
rect 3693 553074 3759 553077
rect -960 553072 3759 553074
rect -960 553016 3698 553072
rect 3754 553016 3759 553072
rect -960 553014 3759 553016
rect -960 552924 480 553014
rect 3693 553011 3759 553014
rect 491753 549266 491819 549269
rect 494605 549266 494671 549269
rect 491753 549264 494671 549266
rect 491753 549208 491758 549264
rect 491814 549208 494610 549264
rect 494666 549208 494671 549264
rect 491753 549206 494671 549208
rect 491753 549203 491819 549206
rect 494605 549203 494671 549206
rect 207565 545730 207631 545733
rect 202830 545728 207631 545730
rect 202830 545672 207570 545728
rect 207626 545672 207631 545728
rect 202830 545670 207631 545672
rect 57462 545532 57468 545596
rect 57532 545594 57538 545596
rect 57532 545534 60842 545594
rect 57532 545532 57538 545534
rect 60782 545322 60842 545534
rect 115933 545458 115999 545461
rect 135253 545458 135319 545461
rect 195881 545458 195947 545461
rect 108990 545456 115999 545458
rect 108990 545400 115938 545456
rect 115994 545400 115999 545456
rect 108990 545398 115999 545400
rect 85573 545322 85639 545325
rect 60782 545262 72434 545322
rect 72374 545186 72434 545262
rect 85438 545320 85639 545322
rect 85438 545264 85578 545320
rect 85634 545264 85639 545320
rect 85438 545262 85639 545264
rect 75862 545186 75868 545188
rect 72374 545126 75868 545186
rect 75862 545124 75868 545126
rect 75932 545124 75938 545188
rect 80697 545186 80763 545189
rect 85438 545186 85498 545262
rect 85573 545259 85639 545262
rect 95049 545322 95115 545325
rect 96613 545322 96679 545325
rect 95049 545320 96679 545322
rect 95049 545264 95054 545320
rect 95110 545264 96618 545320
rect 96674 545264 96679 545320
rect 95049 545262 96679 545264
rect 95049 545259 95115 545262
rect 96613 545259 96679 545262
rect 80697 545184 85498 545186
rect 80697 545128 80702 545184
rect 80758 545128 85498 545184
rect 80697 545126 85498 545128
rect 104801 545186 104867 545189
rect 108990 545186 109050 545398
rect 115933 545395 115999 545398
rect 128310 545456 135319 545458
rect 128310 545400 135258 545456
rect 135314 545400 135319 545456
rect 128310 545398 135319 545400
rect 104801 545184 109050 545186
rect 104801 545128 104806 545184
rect 104862 545128 109050 545184
rect 104801 545126 109050 545128
rect 125409 545186 125475 545189
rect 128310 545186 128370 545398
rect 135253 545395 135319 545398
rect 147630 545398 157442 545458
rect 125409 545184 128370 545186
rect 125409 545128 125414 545184
rect 125470 545128 128370 545184
rect 125409 545126 128370 545128
rect 144821 545186 144887 545189
rect 147630 545186 147690 545398
rect 157382 545322 157442 545398
rect 191790 545456 195947 545458
rect 191790 545400 195886 545456
rect 195942 545400 195947 545456
rect 191790 545398 195947 545400
rect 166901 545322 166967 545325
rect 157382 545320 166967 545322
rect 157382 545264 166906 545320
rect 166962 545264 166967 545320
rect 157382 545262 166967 545264
rect 166901 545259 166967 545262
rect 177297 545322 177363 545325
rect 191790 545322 191850 545398
rect 195881 545395 195947 545398
rect 201401 545458 201467 545461
rect 202830 545458 202890 545670
rect 207565 545667 207631 545670
rect 309041 545594 309107 545597
rect 371877 545594 371943 545597
rect 309041 545592 312002 545594
rect 309041 545536 309046 545592
rect 309102 545536 312002 545592
rect 309041 545534 312002 545536
rect 309041 545531 309107 545534
rect 201401 545456 202890 545458
rect 201401 545400 201406 545456
rect 201462 545400 202890 545456
rect 201401 545398 202890 545400
rect 207565 545458 207631 545461
rect 212533 545458 212599 545461
rect 231853 545458 231919 545461
rect 251173 545458 251239 545461
rect 302141 545458 302207 545461
rect 207565 545456 212599 545458
rect 207565 545400 207570 545456
rect 207626 545400 212538 545456
rect 212594 545400 212599 545456
rect 207565 545398 212599 545400
rect 201401 545395 201467 545398
rect 207565 545395 207631 545398
rect 212533 545395 212599 545398
rect 224910 545456 231919 545458
rect 224910 545400 231858 545456
rect 231914 545400 231919 545456
rect 224910 545398 231919 545400
rect 177297 545320 191850 545322
rect 177297 545264 177302 545320
rect 177358 545264 191850 545320
rect 177297 545262 191850 545264
rect 177297 545259 177363 545262
rect 144821 545184 147690 545186
rect 144821 545128 144826 545184
rect 144882 545128 147690 545184
rect 144821 545126 147690 545128
rect 222009 545186 222075 545189
rect 224910 545186 224970 545398
rect 231853 545395 231919 545398
rect 244230 545456 251239 545458
rect 244230 545400 251178 545456
rect 251234 545400 251239 545456
rect 244230 545398 251239 545400
rect 222009 545184 224970 545186
rect 222009 545128 222014 545184
rect 222070 545128 224970 545184
rect 222009 545126 224970 545128
rect 241421 545186 241487 545189
rect 244230 545186 244290 545398
rect 251173 545395 251239 545398
rect 263550 545398 282930 545458
rect 241421 545184 244290 545186
rect 241421 545128 241426 545184
rect 241482 545128 244290 545184
rect 241421 545126 244290 545128
rect 260741 545186 260807 545189
rect 263550 545186 263610 545398
rect 282870 545322 282930 545398
rect 292622 545456 302207 545458
rect 292622 545400 302146 545456
rect 302202 545400 302207 545456
rect 292622 545398 302207 545400
rect 282870 545262 292498 545322
rect 260741 545184 263610 545186
rect 260741 545128 260746 545184
rect 260802 545128 263610 545184
rect 260741 545126 263610 545128
rect 292438 545186 292498 545262
rect 292622 545186 292682 545398
rect 302141 545395 302207 545398
rect 311942 545322 312002 545534
rect 367142 545592 371943 545594
rect 367142 545536 371882 545592
rect 371938 545536 371943 545592
rect 367142 545534 371943 545536
rect 328361 545458 328427 545461
rect 347681 545458 347747 545461
rect 347814 545458 347820 545460
rect 328361 545456 331322 545458
rect 328361 545400 328366 545456
rect 328422 545400 331322 545456
rect 328361 545398 331322 545400
rect 328361 545395 328427 545398
rect 321461 545322 321527 545325
rect 311942 545320 321527 545322
rect 311942 545264 321466 545320
rect 321522 545264 321527 545320
rect 311942 545262 321527 545264
rect 331262 545322 331322 545398
rect 347681 545456 347820 545458
rect 347681 545400 347686 545456
rect 347742 545400 347820 545456
rect 347681 545398 347820 545400
rect 347681 545395 347747 545398
rect 347814 545396 347820 545398
rect 347884 545396 347890 545460
rect 347681 545322 347747 545325
rect 331262 545320 347747 545322
rect 331262 545264 347686 545320
rect 347742 545264 347747 545320
rect 331262 545262 347747 545264
rect 321461 545259 321527 545262
rect 347681 545259 347747 545262
rect 367001 545322 367067 545325
rect 367142 545322 367202 545534
rect 371877 545531 371943 545534
rect 550582 545532 550588 545596
rect 550652 545594 550658 545596
rect 553301 545594 553367 545597
rect 550652 545592 553367 545594
rect 550652 545536 553306 545592
rect 553362 545536 553367 545592
rect 550652 545534 553367 545536
rect 550652 545532 550658 545534
rect 553301 545531 553367 545534
rect 553485 545594 553551 545597
rect 560293 545594 560359 545597
rect 553485 545592 560359 545594
rect 553485 545536 553490 545592
rect 553546 545536 560298 545592
rect 560354 545536 560359 545592
rect 553485 545534 560359 545536
rect 553485 545531 553551 545534
rect 560293 545531 560359 545534
rect 579521 545594 579587 545597
rect 583520 545594 584960 545684
rect 579521 545592 584960 545594
rect 579521 545536 579526 545592
rect 579582 545536 584960 545592
rect 579521 545534 584960 545536
rect 579521 545531 579587 545534
rect 376702 545396 376708 545460
rect 376772 545458 376778 545460
rect 483013 545458 483079 545461
rect 376772 545398 393330 545458
rect 376772 545396 376778 545398
rect 367001 545320 367202 545322
rect 367001 545264 367006 545320
rect 367062 545264 367202 545320
rect 367001 545262 367202 545264
rect 393270 545322 393330 545398
rect 403022 545398 427738 545458
rect 393270 545262 402898 545322
rect 367001 545259 367067 545262
rect 292438 545126 292682 545186
rect 80697 545123 80763 545126
rect 104801 545123 104867 545126
rect 125409 545123 125475 545126
rect 144821 545123 144887 545126
rect 222009 545123 222075 545126
rect 241421 545123 241487 545126
rect 260741 545123 260807 545126
rect 347814 545124 347820 545188
rect 347884 545186 347890 545188
rect 357382 545186 357388 545188
rect 347884 545126 357388 545186
rect 347884 545124 347890 545126
rect 357382 545124 357388 545126
rect 357452 545124 357458 545188
rect 371877 545186 371943 545189
rect 376702 545186 376708 545188
rect 371877 545184 376708 545186
rect 371877 545128 371882 545184
rect 371938 545128 376708 545184
rect 371877 545126 376708 545128
rect 371877 545123 371943 545126
rect 376702 545124 376708 545126
rect 376772 545124 376778 545188
rect 402838 545186 402898 545262
rect 403022 545186 403082 545398
rect 402838 545126 403082 545186
rect 427678 545050 427738 545398
rect 441662 545398 451290 545458
rect 441662 545186 441722 545398
rect 451230 545322 451290 545398
rect 460982 545398 470610 545458
rect 451230 545262 460858 545322
rect 434670 545126 441722 545186
rect 460798 545186 460858 545262
rect 460982 545186 461042 545398
rect 470550 545322 470610 545398
rect 480302 545456 483079 545458
rect 480302 545400 483018 545456
rect 483074 545400 483079 545456
rect 480302 545398 483079 545400
rect 470550 545262 480178 545322
rect 460798 545126 461042 545186
rect 480118 545186 480178 545262
rect 480302 545186 480362 545398
rect 483013 545395 483079 545398
rect 492622 545396 492628 545460
rect 492692 545458 492698 545460
rect 540973 545458 541039 545461
rect 572621 545458 572687 545461
rect 492692 545398 509250 545458
rect 492692 545396 492698 545398
rect 509190 545322 509250 545398
rect 518942 545398 528570 545458
rect 509190 545262 518818 545322
rect 480118 545126 480362 545186
rect 485865 545186 485931 545189
rect 492622 545186 492628 545188
rect 485865 545184 492628 545186
rect 485865 545128 485870 545184
rect 485926 545128 492628 545184
rect 485865 545126 492628 545128
rect 434670 545050 434730 545126
rect 485865 545123 485931 545126
rect 492622 545124 492628 545126
rect 492692 545124 492698 545188
rect 518758 545186 518818 545262
rect 518942 545186 519002 545398
rect 528510 545322 528570 545398
rect 538262 545456 541039 545458
rect 538262 545400 540978 545456
rect 541034 545400 541039 545456
rect 538262 545398 541039 545400
rect 528510 545262 538138 545322
rect 518758 545126 519002 545186
rect 538078 545186 538138 545262
rect 538262 545186 538322 545398
rect 540973 545395 541039 545398
rect 569910 545456 572687 545458
rect 569910 545400 572626 545456
rect 572682 545400 572687 545456
rect 583520 545444 584960 545534
rect 569910 545398 572687 545400
rect 563145 545322 563211 545325
rect 569910 545322 569970 545398
rect 572621 545395 572687 545398
rect 563145 545320 569970 545322
rect 563145 545264 563150 545320
rect 563206 545264 569970 545320
rect 563145 545262 569970 545264
rect 563145 545259 563211 545262
rect 538078 545126 538322 545186
rect 548609 545186 548675 545189
rect 550582 545186 550588 545188
rect 548609 545184 550588 545186
rect 548609 545128 548614 545184
rect 548670 545128 550588 545184
rect 548609 545126 550588 545128
rect 548609 545123 548675 545126
rect 550582 545124 550588 545126
rect 550652 545124 550658 545188
rect 427678 544990 434730 545050
rect 75862 544852 75868 544916
rect 75932 544914 75938 544916
rect 80697 544914 80763 544917
rect 75932 544912 80763 544914
rect 75932 544856 80702 544912
rect 80758 544856 80763 544912
rect 75932 544854 80763 544856
rect 75932 544852 75938 544854
rect 80697 544851 80763 544854
rect 357382 544852 357388 544916
rect 357452 544914 357458 544916
rect 367001 544914 367067 544917
rect 357452 544912 367067 544914
rect 357452 544856 367006 544912
rect 367062 544856 367067 544912
rect 357452 544854 367067 544856
rect 357452 544852 357458 544854
rect 367001 544851 367067 544854
rect 92105 544778 92171 544781
rect 188521 544778 188587 544781
rect 92105 544776 188587 544778
rect 92105 544720 92110 544776
rect 92166 544720 188526 544776
rect 188582 544720 188587 544776
rect 92105 544718 188587 544720
rect 92105 544715 92171 544718
rect 188521 544715 188587 544718
rect 87965 544642 88031 544645
rect 188705 544642 188771 544645
rect 87965 544640 188771 544642
rect 87965 544584 87970 544640
rect 88026 544584 188710 544640
rect 188766 544584 188771 544640
rect 87965 544582 188771 544584
rect 87965 544579 88031 544582
rect 188705 544579 188771 544582
rect 85849 544506 85915 544509
rect 188889 544506 188955 544509
rect 85849 544504 188955 544506
rect 85849 544448 85854 544504
rect 85910 544448 188894 544504
rect 188950 544448 188955 544504
rect 85849 544446 188955 544448
rect 85849 544443 85915 544446
rect 188889 544443 188955 544446
rect 83825 544370 83891 544373
rect 188245 544370 188311 544373
rect 83825 544368 188311 544370
rect 83825 544312 83830 544368
rect 83886 544312 188250 544368
rect 188306 544312 188311 544368
rect 83825 544310 188311 544312
rect 83825 544307 83891 544310
rect 188245 544307 188311 544310
rect 141509 543282 141575 543285
rect 208301 543282 208367 543285
rect 141509 543280 208367 543282
rect 141509 543224 141514 543280
rect 141570 543224 208306 543280
rect 208362 543224 208367 543280
rect 141509 543222 208367 543224
rect 141509 543219 141575 543222
rect 208301 543219 208367 543222
rect 144177 543146 144243 543149
rect 210417 543146 210483 543149
rect 144177 543144 210483 543146
rect 144177 543088 144182 543144
rect 144238 543088 210422 543144
rect 210478 543088 210483 543144
rect 144177 543086 210483 543088
rect 144177 543083 144243 543086
rect 210417 543083 210483 543086
rect 106181 543010 106247 543013
rect 206185 543010 206251 543013
rect 106181 543008 206251 543010
rect 106181 542952 106186 543008
rect 106242 542952 206190 543008
rect 206246 542952 206251 543008
rect 106181 542950 206251 542952
rect 106181 542947 106247 542950
rect 206185 542947 206251 542950
rect 59486 540364 59492 540428
rect 59556 540426 59562 540428
rect 559189 540426 559255 540429
rect 59556 540424 559255 540426
rect 59556 540368 559194 540424
rect 559250 540368 559255 540424
rect 59556 540366 559255 540368
rect 59556 540364 59562 540366
rect 559189 540363 559255 540366
rect 57278 540228 57284 540292
rect 57348 540290 57354 540292
rect 580625 540290 580691 540293
rect 57348 540288 580691 540290
rect 57348 540232 580630 540288
rect 580686 540232 580691 540288
rect 57348 540230 580691 540232
rect 57348 540228 57354 540230
rect 580625 540227 580691 540230
rect 57421 539066 57487 539069
rect 57421 539064 60076 539066
rect 57421 539008 57426 539064
rect 57482 539008 60076 539064
rect 57421 539006 60076 539008
rect 57421 539003 57487 539006
rect -960 538658 480 538748
rect 3785 538658 3851 538661
rect -960 538656 3851 538658
rect -960 538600 3790 538656
rect 3846 538600 3851 538656
rect -960 538598 3851 538600
rect -960 538508 480 538598
rect 3785 538595 3851 538598
rect 57421 537162 57487 537165
rect 57421 537160 60076 537162
rect 57421 537104 57426 537160
rect 57482 537104 60076 537160
rect 57421 537102 60076 537104
rect 57421 537099 57487 537102
rect 57421 535258 57487 535261
rect 57421 535256 60076 535258
rect 57421 535200 57426 535256
rect 57482 535200 60076 535256
rect 57421 535198 60076 535200
rect 57421 535195 57487 535198
rect 580901 533898 580967 533901
rect 583520 533898 584960 533988
rect 580901 533896 584960 533898
rect 580901 533840 580906 533896
rect 580962 533840 584960 533896
rect 580901 533838 584960 533840
rect 580901 533835 580967 533838
rect 583520 533748 584960 533838
rect 57421 533354 57487 533357
rect 57421 533352 60076 533354
rect 57421 533296 57426 533352
rect 57482 533296 60076 533352
rect 57421 533294 60076 533296
rect 57421 533291 57487 533294
rect 57421 531450 57487 531453
rect 57421 531448 60076 531450
rect 57421 531392 57426 531448
rect 57482 531392 60076 531448
rect 57421 531390 60076 531392
rect 57421 531387 57487 531390
rect 57421 529410 57487 529413
rect 57421 529408 60076 529410
rect 57421 529352 57426 529408
rect 57482 529352 60076 529408
rect 57421 529350 60076 529352
rect 57421 529347 57487 529350
rect 57421 527506 57487 527509
rect 57421 527504 60076 527506
rect 57421 527448 57426 527504
rect 57482 527448 60076 527504
rect 57421 527446 60076 527448
rect 57421 527443 57487 527446
rect 57421 525602 57487 525605
rect 57421 525600 60076 525602
rect 57421 525544 57426 525600
rect 57482 525544 60076 525600
rect 57421 525542 60076 525544
rect 57421 525539 57487 525542
rect -960 524092 480 524332
rect 57421 523698 57487 523701
rect 57421 523696 60076 523698
rect 57421 523640 57426 523696
rect 57482 523640 60076 523696
rect 57421 523638 60076 523640
rect 57421 523635 57487 523638
rect 583520 521916 584960 522156
rect 57421 521794 57487 521797
rect 57421 521792 60076 521794
rect 57421 521736 57426 521792
rect 57482 521736 60076 521792
rect 57421 521734 60076 521736
rect 57421 521731 57487 521734
rect 57421 519754 57487 519757
rect 57421 519752 60076 519754
rect 57421 519696 57426 519752
rect 57482 519696 60076 519752
rect 57421 519694 60076 519696
rect 57421 519691 57487 519694
rect 57421 517850 57487 517853
rect 57421 517848 60076 517850
rect 57421 517792 57426 517848
rect 57482 517792 60076 517848
rect 57421 517790 60076 517792
rect 57421 517787 57487 517790
rect 57421 515946 57487 515949
rect 57421 515944 60076 515946
rect 57421 515888 57426 515944
rect 57482 515888 60076 515944
rect 57421 515886 60076 515888
rect 57421 515883 57487 515886
rect 57421 514042 57487 514045
rect 57421 514040 60076 514042
rect 57421 513984 57426 514040
rect 57482 513984 60076 514040
rect 57421 513982 60076 513984
rect 57421 513979 57487 513982
rect 57421 512138 57487 512141
rect 57421 512136 60076 512138
rect 57421 512080 57426 512136
rect 57482 512080 60076 512136
rect 57421 512078 60076 512080
rect 57421 512075 57487 512078
rect 580809 510370 580875 510373
rect 583520 510370 584960 510460
rect 580809 510368 584960 510370
rect 580809 510312 580814 510368
rect 580870 510312 584960 510368
rect 580809 510310 584960 510312
rect 580809 510307 580875 510310
rect 583520 510220 584960 510310
rect 57421 510098 57487 510101
rect 57421 510096 60076 510098
rect -960 509962 480 510052
rect 57421 510040 57426 510096
rect 57482 510040 60076 510096
rect 57421 510038 60076 510040
rect 57421 510035 57487 510038
rect 4061 509962 4127 509965
rect -960 509960 4127 509962
rect -960 509904 4066 509960
rect 4122 509904 4127 509960
rect -960 509902 4127 509904
rect -960 509812 480 509902
rect 4061 509899 4127 509902
rect 57421 508194 57487 508197
rect 57421 508192 60076 508194
rect 57421 508136 57426 508192
rect 57482 508136 60076 508192
rect 57421 508134 60076 508136
rect 57421 508131 57487 508134
rect 57237 506290 57303 506293
rect 57237 506288 60076 506290
rect 57237 506232 57242 506288
rect 57298 506232 60076 506288
rect 57237 506230 60076 506232
rect 57237 506227 57303 506230
rect 57421 504386 57487 504389
rect 57421 504384 60076 504386
rect 57421 504328 57426 504384
rect 57482 504328 60076 504384
rect 57421 504326 60076 504328
rect 57421 504323 57487 504326
rect 57421 502482 57487 502485
rect 57421 502480 60076 502482
rect 57421 502424 57426 502480
rect 57482 502424 60076 502480
rect 57421 502422 60076 502424
rect 57421 502419 57487 502422
rect 57329 500442 57395 500445
rect 57329 500440 60076 500442
rect 57329 500384 57334 500440
rect 57390 500384 60076 500440
rect 57329 500382 60076 500384
rect 57329 500379 57395 500382
rect 580257 498674 580323 498677
rect 583520 498674 584960 498764
rect 580257 498672 584960 498674
rect 580257 498616 580262 498672
rect 580318 498616 584960 498672
rect 580257 498614 584960 498616
rect 580257 498611 580323 498614
rect 57421 498538 57487 498541
rect 57421 498536 60076 498538
rect 57421 498480 57426 498536
rect 57482 498480 60076 498536
rect 583520 498524 584960 498614
rect 57421 498478 60076 498480
rect 57421 498475 57487 498478
rect 57421 496634 57487 496637
rect 57421 496632 60076 496634
rect 57421 496576 57426 496632
rect 57482 496576 60076 496632
rect 57421 496574 60076 496576
rect 57421 496571 57487 496574
rect -960 495546 480 495636
rect 3969 495546 4035 495549
rect -960 495544 4035 495546
rect -960 495488 3974 495544
rect 4030 495488 4035 495544
rect -960 495486 4035 495488
rect -960 495396 480 495486
rect 3969 495483 4035 495486
rect 57421 494730 57487 494733
rect 57421 494728 60076 494730
rect 57421 494672 57426 494728
rect 57482 494672 60076 494728
rect 57421 494670 60076 494672
rect 57421 494667 57487 494670
rect 57053 492826 57119 492829
rect 57053 492824 60076 492826
rect 57053 492768 57058 492824
rect 57114 492768 60076 492824
rect 57053 492766 60076 492768
rect 57053 492763 57119 492766
rect 282361 492690 282427 492693
rect 282545 492690 282611 492693
rect 282361 492688 282611 492690
rect 282361 492632 282366 492688
rect 282422 492632 282550 492688
rect 282606 492632 282611 492688
rect 282361 492630 282611 492632
rect 282361 492627 282427 492630
rect 282545 492627 282611 492630
rect 56685 490786 56751 490789
rect 56685 490784 60076 490786
rect 56685 490728 56690 490784
rect 56746 490728 60076 490784
rect 56685 490726 60076 490728
rect 56685 490723 56751 490726
rect 56593 488882 56659 488885
rect 56593 488880 60076 488882
rect 56593 488824 56598 488880
rect 56654 488824 60076 488880
rect 56593 488822 60076 488824
rect 56593 488819 56659 488822
rect 56685 486978 56751 486981
rect 56685 486976 60076 486978
rect 56685 486920 56690 486976
rect 56746 486920 60076 486976
rect 56685 486918 60076 486920
rect 56685 486915 56751 486918
rect 580533 486842 580599 486845
rect 583520 486842 584960 486932
rect 580533 486840 584960 486842
rect 580533 486784 580538 486840
rect 580594 486784 584960 486840
rect 580533 486782 584960 486784
rect 580533 486779 580599 486782
rect 583520 486692 584960 486782
rect 56685 485074 56751 485077
rect 56685 485072 60076 485074
rect 56685 485016 56690 485072
rect 56746 485016 60076 485072
rect 56685 485014 60076 485016
rect 56685 485011 56751 485014
rect 56593 483170 56659 483173
rect 56593 483168 60076 483170
rect 56593 483112 56598 483168
rect 56654 483112 60076 483168
rect 56593 483110 60076 483112
rect 56593 483107 56659 483110
rect 56685 481266 56751 481269
rect 56685 481264 60076 481266
rect -960 481130 480 481220
rect 56685 481208 56690 481264
rect 56746 481208 60076 481264
rect 56685 481206 60076 481208
rect 56685 481203 56751 481206
rect 2865 481130 2931 481133
rect -960 481128 2931 481130
rect -960 481072 2870 481128
rect 2926 481072 2931 481128
rect -960 481070 2931 481072
rect -960 480980 480 481070
rect 2865 481067 2931 481070
rect 56501 479226 56567 479229
rect 56501 479224 60076 479226
rect 56501 479168 56506 479224
rect 56562 479168 60076 479224
rect 56501 479166 60076 479168
rect 56501 479163 56567 479166
rect 56501 477322 56567 477325
rect 56501 477320 60076 477322
rect 56501 477264 56506 477320
rect 56562 477264 60076 477320
rect 56501 477262 60076 477264
rect 56501 477259 56567 477262
rect 56501 475418 56567 475421
rect 56501 475416 60076 475418
rect 56501 475360 56506 475416
rect 56562 475360 60076 475416
rect 56501 475358 60076 475360
rect 56501 475355 56567 475358
rect 583520 474996 584960 475236
rect 56501 473514 56567 473517
rect 56501 473512 60076 473514
rect 56501 473456 56506 473512
rect 56562 473456 60076 473512
rect 56501 473454 60076 473456
rect 56501 473451 56567 473454
rect 282361 473378 282427 473381
rect 282545 473378 282611 473381
rect 282361 473376 282611 473378
rect 282361 473320 282366 473376
rect 282422 473320 282550 473376
rect 282606 473320 282611 473376
rect 282361 473318 282611 473320
rect 282361 473315 282427 473318
rect 282545 473315 282611 473318
rect 56501 471610 56567 471613
rect 56501 471608 60076 471610
rect 56501 471552 56506 471608
rect 56562 471552 60076 471608
rect 56501 471550 60076 471552
rect 56501 471547 56567 471550
rect 56501 469570 56567 469573
rect 56501 469568 60076 469570
rect 56501 469512 56506 469568
rect 56562 469512 60076 469568
rect 56501 469510 60076 469512
rect 56501 469507 56567 469510
rect 56501 467666 56567 467669
rect 56501 467664 60076 467666
rect 56501 467608 56506 467664
rect 56562 467608 60076 467664
rect 56501 467606 60076 467608
rect 56501 467603 56567 467606
rect -960 466700 480 466940
rect 56501 465762 56567 465765
rect 56501 465760 60076 465762
rect 56501 465704 56506 465760
rect 56562 465704 60076 465760
rect 56501 465702 60076 465704
rect 56501 465699 56567 465702
rect 56501 463858 56567 463861
rect 56501 463856 60076 463858
rect 56501 463800 56506 463856
rect 56562 463800 60076 463856
rect 56501 463798 60076 463800
rect 56501 463795 56567 463798
rect 580257 463450 580323 463453
rect 583520 463450 584960 463540
rect 580257 463448 584960 463450
rect 580257 463392 580262 463448
rect 580318 463392 584960 463448
rect 580257 463390 584960 463392
rect 580257 463387 580323 463390
rect 583520 463300 584960 463390
rect 56501 461954 56567 461957
rect 56501 461952 60076 461954
rect 56501 461896 56506 461952
rect 56562 461896 60076 461952
rect 56501 461894 60076 461896
rect 56501 461891 56567 461894
rect 56593 459914 56659 459917
rect 56593 459912 60076 459914
rect 56593 459856 56598 459912
rect 56654 459856 60076 459912
rect 56593 459854 60076 459856
rect 56593 459851 56659 459854
rect 56593 458010 56659 458013
rect 56593 458008 60076 458010
rect 56593 457952 56598 458008
rect 56654 457952 60076 458008
rect 56593 457950 60076 457952
rect 56593 457947 56659 457950
rect 56593 456106 56659 456109
rect 56593 456104 60076 456106
rect 56593 456048 56598 456104
rect 56654 456048 60076 456104
rect 56593 456046 60076 456048
rect 56593 456043 56659 456046
rect 56593 454202 56659 454205
rect 56593 454200 60076 454202
rect 56593 454144 56598 454200
rect 56654 454144 60076 454200
rect 56593 454142 60076 454144
rect 56593 454139 56659 454142
rect 282361 454066 282427 454069
rect 282545 454066 282611 454069
rect 282361 454064 282611 454066
rect 282361 454008 282366 454064
rect 282422 454008 282550 454064
rect 282606 454008 282611 454064
rect 282361 454006 282611 454008
rect 282361 454003 282427 454006
rect 282545 454003 282611 454006
rect -960 452434 480 452524
rect 3417 452434 3483 452437
rect -960 452432 3483 452434
rect -960 452376 3422 452432
rect 3478 452376 3483 452432
rect -960 452374 3483 452376
rect -960 452284 480 452374
rect 3417 452371 3483 452374
rect 58341 452298 58407 452301
rect 58341 452296 60076 452298
rect 58341 452240 58346 452296
rect 58402 452240 60076 452296
rect 58341 452238 60076 452240
rect 58341 452235 58407 452238
rect 580349 451754 580415 451757
rect 583520 451754 584960 451844
rect 580349 451752 584960 451754
rect 580349 451696 580354 451752
rect 580410 451696 584960 451752
rect 580349 451694 584960 451696
rect 580349 451691 580415 451694
rect 583520 451604 584960 451694
rect 58433 450258 58499 450261
rect 58433 450256 60076 450258
rect 58433 450200 58438 450256
rect 58494 450200 60076 450256
rect 58433 450198 60076 450200
rect 58433 450195 58499 450198
rect 57697 448354 57763 448357
rect 57697 448352 60076 448354
rect 57697 448296 57702 448352
rect 57758 448296 60076 448352
rect 57697 448294 60076 448296
rect 57697 448291 57763 448294
rect 58525 446450 58591 446453
rect 58525 446448 60076 446450
rect 58525 446392 58530 446448
rect 58586 446392 60076 446448
rect 58525 446390 60076 446392
rect 58525 446387 58591 446390
rect 58617 444546 58683 444549
rect 58617 444544 60076 444546
rect 58617 444488 58622 444544
rect 58678 444488 60076 444544
rect 58617 444486 60076 444488
rect 58617 444483 58683 444486
rect 56777 442642 56843 442645
rect 56777 442640 60076 442642
rect 56777 442584 56782 442640
rect 56838 442584 60076 442640
rect 56777 442582 60076 442584
rect 56777 442579 56843 442582
rect 57789 440602 57855 440605
rect 57789 440600 60076 440602
rect 57789 440544 57794 440600
rect 57850 440544 60076 440600
rect 57789 440542 60076 440544
rect 57789 440539 57855 440542
rect 580441 439922 580507 439925
rect 583520 439922 584960 440012
rect 580441 439920 584960 439922
rect 580441 439864 580446 439920
rect 580502 439864 584960 439920
rect 580441 439862 584960 439864
rect 580441 439859 580507 439862
rect 583520 439772 584960 439862
rect 58709 438698 58775 438701
rect 58709 438696 60076 438698
rect 58709 438640 58714 438696
rect 58770 438640 60076 438696
rect 58709 438638 60076 438640
rect 58709 438635 58775 438638
rect -960 438018 480 438108
rect 3969 438018 4035 438021
rect -960 438016 4035 438018
rect -960 437960 3974 438016
rect 4030 437960 4035 438016
rect -960 437958 4035 437960
rect -960 437868 480 437958
rect 3969 437955 4035 437958
rect 56869 436794 56935 436797
rect 56869 436792 60076 436794
rect 56869 436736 56874 436792
rect 56930 436736 60076 436792
rect 56869 436734 60076 436736
rect 56869 436731 56935 436734
rect 58801 434890 58867 434893
rect 58801 434888 60076 434890
rect 58801 434832 58806 434888
rect 58862 434832 60076 434888
rect 58801 434830 60076 434832
rect 58801 434827 58867 434830
rect 58893 432986 58959 432989
rect 58893 432984 60076 432986
rect 58893 432928 58898 432984
rect 58954 432928 60076 432984
rect 58893 432926 60076 432928
rect 58893 432923 58959 432926
rect 56961 431082 57027 431085
rect 56961 431080 60076 431082
rect 56961 431024 56966 431080
rect 57022 431024 60076 431080
rect 56961 431022 60076 431024
rect 56961 431019 57027 431022
rect 281533 429450 281599 429453
rect 279956 429448 281599 429450
rect 279956 429392 281538 429448
rect 281594 429392 281599 429448
rect 279956 429390 281599 429392
rect 281533 429387 281599 429390
rect 57881 429042 57947 429045
rect 57881 429040 60076 429042
rect 57881 428984 57886 429040
rect 57942 428984 60076 429040
rect 57881 428982 60076 428984
rect 57881 428979 57947 428982
rect 281533 428498 281599 428501
rect 279956 428496 281599 428498
rect 279956 428440 281538 428496
rect 281594 428440 281599 428496
rect 279956 428438 281599 428440
rect 281533 428435 281599 428438
rect 583520 428076 584960 428316
rect 281625 427410 281691 427413
rect 279956 427408 281691 427410
rect 279956 427352 281630 427408
rect 281686 427352 281691 427408
rect 279956 427350 281691 427352
rect 281625 427347 281691 427350
rect 58985 427138 59051 427141
rect 58985 427136 60076 427138
rect 58985 427080 58990 427136
rect 59046 427080 60076 427136
rect 58985 427078 60076 427080
rect 58985 427075 59051 427078
rect 281533 426458 281599 426461
rect 279956 426456 281599 426458
rect 279956 426400 281538 426456
rect 281594 426400 281599 426456
rect 279956 426398 281599 426400
rect 281533 426395 281599 426398
rect 281533 425370 281599 425373
rect 279956 425368 281599 425370
rect 279956 425312 281538 425368
rect 281594 425312 281599 425368
rect 279956 425310 281599 425312
rect 281533 425307 281599 425310
rect 59445 425234 59511 425237
rect 59445 425232 60076 425234
rect 59445 425176 59450 425232
rect 59506 425176 60076 425232
rect 59445 425174 60076 425176
rect 59445 425171 59511 425174
rect 282637 425098 282703 425101
rect 283005 425098 283071 425101
rect 282637 425096 283071 425098
rect 282637 425040 282642 425096
rect 282698 425040 283010 425096
rect 283066 425040 283071 425096
rect 282637 425038 283071 425040
rect 282637 425035 282703 425038
rect 283005 425035 283071 425038
rect 281533 424418 281599 424421
rect 279956 424416 281599 424418
rect 279956 424360 281538 424416
rect 281594 424360 281599 424416
rect 279956 424358 281599 424360
rect 281533 424355 281599 424358
rect -960 423738 480 423828
rect 3877 423738 3943 423741
rect -960 423736 3943 423738
rect -960 423680 3882 423736
rect 3938 423680 3943 423736
rect -960 423678 3943 423680
rect -960 423588 480 423678
rect 3877 423675 3943 423678
rect 281625 423466 281691 423469
rect 279956 423464 281691 423466
rect 279956 423408 281630 423464
rect 281686 423408 281691 423464
rect 279956 423406 281691 423408
rect 281625 423403 281691 423406
rect 59077 423330 59143 423333
rect 59077 423328 60076 423330
rect 59077 423272 59082 423328
rect 59138 423272 60076 423328
rect 59077 423270 60076 423272
rect 59077 423267 59143 423270
rect 281533 422378 281599 422381
rect 279956 422376 281599 422378
rect 279956 422320 281538 422376
rect 281594 422320 281599 422376
rect 279956 422318 281599 422320
rect 281533 422315 281599 422318
rect 59169 421426 59235 421429
rect 281533 421426 281599 421429
rect 59169 421424 60076 421426
rect 59169 421368 59174 421424
rect 59230 421368 60076 421424
rect 59169 421366 60076 421368
rect 279956 421424 281599 421426
rect 279956 421368 281538 421424
rect 281594 421368 281599 421424
rect 279956 421366 281599 421368
rect 59169 421363 59235 421366
rect 281533 421363 281599 421366
rect 281533 420338 281599 420341
rect 279956 420336 281599 420338
rect 279956 420280 281538 420336
rect 281594 420280 281599 420336
rect 279956 420278 281599 420280
rect 281533 420275 281599 420278
rect 59445 419386 59511 419389
rect 281625 419386 281691 419389
rect 59445 419384 60076 419386
rect 59445 419328 59450 419384
rect 59506 419328 60076 419384
rect 59445 419326 60076 419328
rect 279956 419384 281691 419386
rect 279956 419328 281630 419384
rect 281686 419328 281691 419384
rect 279956 419326 281691 419328
rect 59445 419323 59511 419326
rect 281625 419323 281691 419326
rect 281533 418298 281599 418301
rect 279956 418296 281599 418298
rect 279956 418240 281538 418296
rect 281594 418240 281599 418296
rect 279956 418238 281599 418240
rect 281533 418235 281599 418238
rect 59261 417482 59327 417485
rect 59261 417480 60076 417482
rect 59261 417424 59266 417480
rect 59322 417424 60076 417480
rect 59261 417422 60076 417424
rect 59261 417419 59327 417422
rect 282821 417346 282887 417349
rect 279956 417344 282887 417346
rect 279956 417288 282826 417344
rect 282882 417288 282887 417344
rect 279956 417286 282887 417288
rect 282821 417283 282887 417286
rect 580533 416530 580599 416533
rect 583520 416530 584960 416620
rect 580533 416528 584960 416530
rect 580533 416472 580538 416528
rect 580594 416472 584960 416528
rect 580533 416470 584960 416472
rect 580533 416467 580599 416470
rect 282269 416394 282335 416397
rect 279956 416392 282335 416394
rect 279956 416336 282274 416392
rect 282330 416336 282335 416392
rect 583520 416380 584960 416470
rect 279956 416334 282335 416336
rect 282269 416331 282335 416334
rect 57973 415578 58039 415581
rect 57973 415576 60076 415578
rect 57973 415520 57978 415576
rect 58034 415520 60076 415576
rect 57973 415518 60076 415520
rect 57973 415515 58039 415518
rect 281717 415306 281783 415309
rect 279956 415304 281783 415306
rect 279956 415248 281722 415304
rect 281778 415248 281783 415304
rect 279956 415246 281783 415248
rect 281717 415243 281783 415246
rect 282085 414354 282151 414357
rect 279956 414352 282151 414354
rect 279956 414296 282090 414352
rect 282146 414296 282151 414352
rect 279956 414294 282151 414296
rect 282085 414291 282151 414294
rect 281574 413884 281580 413948
rect 281644 413946 281650 413948
rect 282637 413946 282703 413949
rect 281644 413944 282703 413946
rect 281644 413888 282642 413944
rect 282698 413888 282703 413944
rect 281644 413886 282703 413888
rect 281644 413884 281650 413886
rect 282637 413883 282703 413886
rect 367093 413946 367159 413949
rect 367686 413946 367692 413948
rect 367093 413944 367692 413946
rect 367093 413888 367098 413944
rect 367154 413888 367692 413944
rect 367093 413886 367692 413888
rect 367093 413883 367159 413886
rect 367686 413884 367692 413886
rect 367756 413884 367762 413948
rect 368473 413946 368539 413949
rect 368974 413946 368980 413948
rect 368473 413944 368980 413946
rect 368473 413888 368478 413944
rect 368534 413888 368980 413944
rect 368473 413886 368980 413888
rect 368473 413883 368539 413886
rect 368974 413884 368980 413886
rect 369044 413884 369050 413948
rect 369853 413946 369919 413949
rect 370262 413946 370268 413948
rect 369853 413944 370268 413946
rect 369853 413888 369858 413944
rect 369914 413888 370268 413944
rect 369853 413886 370268 413888
rect 369853 413883 369919 413886
rect 370262 413884 370268 413886
rect 370332 413884 370338 413948
rect 371233 413946 371299 413949
rect 372613 413948 372679 413949
rect 373993 413948 374059 413949
rect 371550 413946 371556 413948
rect 371233 413944 371556 413946
rect 371233 413888 371238 413944
rect 371294 413888 371556 413944
rect 371233 413886 371556 413888
rect 371233 413883 371299 413886
rect 371550 413884 371556 413886
rect 371620 413884 371626 413948
rect 372613 413946 372660 413948
rect 372568 413944 372660 413946
rect 372568 413888 372618 413944
rect 372568 413886 372660 413888
rect 372613 413884 372660 413886
rect 372724 413884 372730 413948
rect 373942 413884 373948 413948
rect 374012 413946 374059 413948
rect 375373 413946 375439 413949
rect 375966 413946 375972 413948
rect 374012 413944 374104 413946
rect 374054 413888 374104 413944
rect 374012 413886 374104 413888
rect 375373 413944 375972 413946
rect 375373 413888 375378 413944
rect 375434 413888 375972 413944
rect 375373 413886 375972 413888
rect 374012 413884 374059 413886
rect 372613 413883 372679 413884
rect 373993 413883 374059 413884
rect 375373 413883 375439 413886
rect 375966 413884 375972 413886
rect 376036 413884 376042 413948
rect 376753 413946 376819 413949
rect 377254 413946 377260 413948
rect 376753 413944 377260 413946
rect 376753 413888 376758 413944
rect 376814 413888 377260 413944
rect 376753 413886 377260 413888
rect 376753 413883 376819 413886
rect 377254 413884 377260 413886
rect 377324 413884 377330 413948
rect 378133 413946 378199 413949
rect 378358 413946 378364 413948
rect 378133 413944 378364 413946
rect 378133 413888 378138 413944
rect 378194 413888 378364 413944
rect 378133 413886 378364 413888
rect 378133 413883 378199 413886
rect 378358 413884 378364 413886
rect 378428 413884 378434 413948
rect 379513 413946 379579 413949
rect 380893 413948 380959 413949
rect 382273 413948 382339 413949
rect 379646 413946 379652 413948
rect 379513 413944 379652 413946
rect 379513 413888 379518 413944
rect 379574 413888 379652 413944
rect 379513 413886 379652 413888
rect 379513 413883 379579 413886
rect 379646 413884 379652 413886
rect 379716 413884 379722 413948
rect 380893 413946 380940 413948
rect 380848 413944 380940 413946
rect 380848 413888 380898 413944
rect 380848 413886 380940 413888
rect 380893 413884 380940 413886
rect 381004 413884 381010 413948
rect 382222 413884 382228 413948
rect 382292 413946 382339 413948
rect 385033 413946 385099 413949
rect 385166 413946 385172 413948
rect 382292 413944 382384 413946
rect 382334 413888 382384 413944
rect 382292 413886 382384 413888
rect 385033 413944 385172 413946
rect 385033 413888 385038 413944
rect 385094 413888 385172 413944
rect 385033 413886 385172 413888
rect 382292 413884 382339 413886
rect 380893 413883 380959 413884
rect 382273 413883 382339 413884
rect 385033 413883 385099 413886
rect 385166 413884 385172 413886
rect 385236 413884 385242 413948
rect 374085 413810 374151 413813
rect 374678 413810 374684 413812
rect 374085 413808 374684 413810
rect 374085 413752 374090 413808
rect 374146 413752 374684 413808
rect 374085 413750 374684 413752
rect 374085 413747 374151 413750
rect 374678 413748 374684 413750
rect 374748 413748 374754 413812
rect 382365 413810 382431 413813
rect 382958 413810 382964 413812
rect 382365 413808 382964 413810
rect 382365 413752 382370 413808
rect 382426 413752 382964 413808
rect 382365 413750 382964 413752
rect 382365 413747 382431 413750
rect 382958 413748 382964 413750
rect 383028 413748 383034 413812
rect 383837 413810 383903 413813
rect 384062 413810 384068 413812
rect 383837 413808 384068 413810
rect 383837 413752 383842 413808
rect 383898 413752 384068 413808
rect 383837 413750 384068 413752
rect 383837 413747 383903 413750
rect 384062 413748 384068 413750
rect 384132 413748 384138 413812
rect 412633 413810 412699 413813
rect 412766 413810 412772 413812
rect 412633 413808 412772 413810
rect 412633 413752 412638 413808
rect 412694 413752 412772 413808
rect 412633 413750 412772 413752
rect 412633 413747 412699 413750
rect 412766 413748 412772 413750
rect 412836 413748 412842 413812
rect 59813 413674 59879 413677
rect 396073 413674 396139 413677
rect 397453 413676 397519 413677
rect 396390 413674 396396 413676
rect 59813 413672 60076 413674
rect 59813 413616 59818 413672
rect 59874 413616 60076 413672
rect 59813 413614 60076 413616
rect 396073 413672 396396 413674
rect 396073 413616 396078 413672
rect 396134 413616 396396 413672
rect 396073 413614 396396 413616
rect 59813 413611 59879 413614
rect 396073 413611 396139 413614
rect 396390 413612 396396 413614
rect 396460 413612 396466 413676
rect 397453 413674 397500 413676
rect 397408 413672 397500 413674
rect 397408 413616 397458 413672
rect 397408 413614 397500 413616
rect 397453 413612 397500 413614
rect 397564 413612 397570 413676
rect 397453 413611 397519 413612
rect 405733 413540 405799 413541
rect 405733 413538 405780 413540
rect 405688 413536 405780 413538
rect 405688 413480 405738 413536
rect 405688 413478 405780 413480
rect 405733 413476 405780 413478
rect 405844 413476 405850 413540
rect 405733 413475 405799 413476
rect 368289 413404 368355 413405
rect 368238 413402 368244 413404
rect 368198 413342 368244 413402
rect 368308 413400 368355 413404
rect 368350 413344 368355 413400
rect 368238 413340 368244 413342
rect 368308 413340 368355 413344
rect 368289 413339 368355 413340
rect 368749 413402 368815 413405
rect 369761 413404 369827 413405
rect 378041 413404 378107 413405
rect 388345 413404 388411 413405
rect 369710 413402 369716 413404
rect 368749 413400 369716 413402
rect 369780 413402 369827 413404
rect 377990 413402 377996 413404
rect 369780 413400 369908 413402
rect 368749 413344 368754 413400
rect 368810 413344 369716 413400
rect 369822 413344 369908 413400
rect 368749 413342 369716 413344
rect 368749 413339 368815 413342
rect 369710 413340 369716 413342
rect 369780 413342 369908 413344
rect 377950 413342 377996 413402
rect 378060 413400 378107 413404
rect 388294 413402 388300 413404
rect 378102 413344 378107 413400
rect 369780 413340 369827 413342
rect 377990 413340 377996 413342
rect 378060 413340 378107 413344
rect 388254 413342 388300 413402
rect 388364 413400 388411 413404
rect 388406 413344 388411 413400
rect 388294 413340 388300 413342
rect 388364 413340 388411 413344
rect 369761 413339 369827 413340
rect 378041 413339 378107 413340
rect 388345 413339 388411 413340
rect 404353 413402 404419 413405
rect 404670 413402 404676 413404
rect 404353 413400 404676 413402
rect 404353 413344 404358 413400
rect 404414 413344 404676 413400
rect 404353 413342 404676 413344
rect 404353 413339 404419 413342
rect 404670 413340 404676 413342
rect 404740 413340 404746 413404
rect 282821 413266 282887 413269
rect 279956 413264 282887 413266
rect 279956 413208 282826 413264
rect 282882 413208 282887 413264
rect 279956 413206 282887 413208
rect 282821 413203 282887 413206
rect 369853 413266 369919 413269
rect 370998 413266 371004 413268
rect 369853 413264 371004 413266
rect 369853 413208 369858 413264
rect 369914 413208 371004 413264
rect 369853 413206 371004 413208
rect 369853 413203 369919 413206
rect 370998 413204 371004 413206
rect 371068 413204 371074 413268
rect 379605 413266 379671 413269
rect 380198 413266 380204 413268
rect 379605 413264 380204 413266
rect 379605 413208 379610 413264
rect 379666 413208 380204 413264
rect 379605 413206 380204 413208
rect 379605 413203 379671 413206
rect 380198 413204 380204 413206
rect 380268 413204 380274 413268
rect 386413 413266 386479 413269
rect 386822 413266 386828 413268
rect 386413 413264 386828 413266
rect 386413 413208 386418 413264
rect 386474 413208 386828 413264
rect 386413 413206 386828 413208
rect 386413 413203 386479 413206
rect 386822 413204 386828 413206
rect 386892 413204 386898 413268
rect 401593 413266 401659 413269
rect 402278 413266 402284 413268
rect 401593 413264 402284 413266
rect 401593 413208 401598 413264
rect 401654 413208 402284 413264
rect 401593 413206 402284 413208
rect 401593 413203 401659 413206
rect 402278 413204 402284 413206
rect 402348 413204 402354 413268
rect 403157 413266 403223 413269
rect 403382 413266 403388 413268
rect 403157 413264 403388 413266
rect 403157 413208 403162 413264
rect 403218 413208 403388 413264
rect 403157 413206 403388 413208
rect 403157 413203 403223 413206
rect 403382 413204 403388 413206
rect 403452 413204 403458 413268
rect 407113 413266 407179 413269
rect 407430 413266 407436 413268
rect 407113 413264 407436 413266
rect 407113 413208 407118 413264
rect 407174 413208 407436 413264
rect 407113 413206 407436 413208
rect 407113 413203 407179 413206
rect 407430 413204 407436 413206
rect 407500 413204 407506 413268
rect 371969 413132 372035 413133
rect 371918 413130 371924 413132
rect 371878 413070 371924 413130
rect 371988 413128 372035 413132
rect 372030 413072 372035 413128
rect 371918 413068 371924 413070
rect 371988 413068 372035 413072
rect 371969 413067 372035 413068
rect 372981 413132 373047 413133
rect 372981 413128 373028 413132
rect 373092 413130 373098 413132
rect 378777 413130 378843 413133
rect 381537 413132 381603 413133
rect 378910 413130 378916 413132
rect 372981 413072 372986 413128
rect 372981 413068 373028 413072
rect 373092 413070 373138 413130
rect 378777 413128 378916 413130
rect 378777 413072 378782 413128
rect 378838 413072 378916 413128
rect 378777 413070 378916 413072
rect 373092 413068 373098 413070
rect 372981 413067 373047 413068
rect 378777 413067 378843 413070
rect 378910 413068 378916 413070
rect 378980 413068 378986 413132
rect 381486 413130 381492 413132
rect 381446 413070 381492 413130
rect 381556 413128 381603 413132
rect 381598 413072 381603 413128
rect 381486 413068 381492 413070
rect 381556 413068 381603 413072
rect 381537 413067 381603 413068
rect 382273 413130 382339 413133
rect 382406 413130 382412 413132
rect 382273 413128 382412 413130
rect 382273 413072 382278 413128
rect 382334 413072 382412 413128
rect 382273 413070 382412 413072
rect 382273 413067 382339 413070
rect 382406 413068 382412 413070
rect 382476 413068 382482 413132
rect 387190 413068 387196 413132
rect 387260 413130 387266 413132
rect 387333 413130 387399 413133
rect 387260 413128 387399 413130
rect 387260 413072 387338 413128
rect 387394 413072 387399 413128
rect 387260 413070 387399 413072
rect 387260 413068 387266 413070
rect 387333 413067 387399 413070
rect 398833 413130 398899 413133
rect 399886 413130 399892 413132
rect 398833 413128 399892 413130
rect 398833 413072 398838 413128
rect 398894 413072 399892 413128
rect 398833 413070 399892 413072
rect 398833 413067 398899 413070
rect 399886 413068 399892 413070
rect 399956 413068 399962 413132
rect 408493 413130 408559 413133
rect 408718 413130 408724 413132
rect 408493 413128 408724 413130
rect 408493 413072 408498 413128
rect 408554 413072 408724 413128
rect 408493 413070 408724 413072
rect 408493 413067 408559 413070
rect 408718 413068 408724 413070
rect 408788 413068 408794 413132
rect 374361 412996 374427 412997
rect 383561 412996 383627 412997
rect 374310 412994 374316 412996
rect 374270 412934 374316 412994
rect 374380 412992 374427 412996
rect 383510 412994 383516 412996
rect 374422 412936 374427 412992
rect 374310 412932 374316 412934
rect 374380 412932 374427 412936
rect 383470 412934 383516 412994
rect 383580 412992 383627 412996
rect 383622 412936 383627 412992
rect 383510 412932 383516 412934
rect 383580 412932 383627 412936
rect 384798 412932 384804 412996
rect 384868 412994 384874 412996
rect 384941 412994 385007 412997
rect 384868 412992 385007 412994
rect 384868 412936 384946 412992
rect 385002 412936 385007 412992
rect 384868 412934 385007 412936
rect 384868 412932 384874 412934
rect 374361 412931 374427 412932
rect 383561 412931 383627 412932
rect 384941 412931 385007 412934
rect 385902 412932 385908 412996
rect 385972 412994 385978 412996
rect 386045 412994 386111 412997
rect 385972 412992 386111 412994
rect 385972 412936 386050 412992
rect 386106 412936 386111 412992
rect 385972 412934 386111 412936
rect 385972 412932 385978 412934
rect 386045 412931 386111 412934
rect 400213 412994 400279 412997
rect 401174 412994 401180 412996
rect 400213 412992 401180 412994
rect 400213 412936 400218 412992
rect 400274 412936 401180 412992
rect 400213 412934 401180 412936
rect 400213 412931 400279 412934
rect 401174 412932 401180 412934
rect 401244 412932 401250 412996
rect 375465 412860 375531 412861
rect 376569 412860 376635 412861
rect 375414 412858 375420 412860
rect 375374 412798 375420 412858
rect 375484 412856 375531 412860
rect 376518 412858 376524 412860
rect 375526 412800 375531 412856
rect 375414 412796 375420 412798
rect 375484 412796 375531 412800
rect 376478 412798 376524 412858
rect 376588 412856 376635 412860
rect 376630 412800 376635 412856
rect 376518 412796 376524 412798
rect 376588 412796 376635 412800
rect 375465 412795 375531 412796
rect 376569 412795 376635 412796
rect 393313 412858 393379 412861
rect 393446 412858 393452 412860
rect 393313 412856 393452 412858
rect 393313 412800 393318 412856
rect 393374 412800 393452 412856
rect 393313 412798 393452 412800
rect 393313 412795 393379 412798
rect 393446 412796 393452 412798
rect 393516 412796 393522 412860
rect 397453 412858 397519 412861
rect 398598 412858 398604 412860
rect 397453 412856 398604 412858
rect 397453 412800 397458 412856
rect 397514 412800 398604 412856
rect 397453 412798 398604 412800
rect 397453 412795 397519 412798
rect 398598 412796 398604 412798
rect 398668 412796 398674 412860
rect 389633 412724 389699 412725
rect 390921 412724 390987 412725
rect 389582 412722 389588 412724
rect 389542 412662 389588 412722
rect 389652 412720 389699 412724
rect 390870 412722 390876 412724
rect 389694 412664 389699 412720
rect 389582 412660 389588 412662
rect 389652 412660 389699 412664
rect 390830 412662 390876 412722
rect 390940 412720 390987 412724
rect 390982 412664 390987 412720
rect 390870 412660 390876 412662
rect 390940 412660 390987 412664
rect 389633 412659 389699 412660
rect 390921 412659 390987 412660
rect 391749 412724 391815 412725
rect 393129 412724 393195 412725
rect 391749 412720 391796 412724
rect 391860 412722 391866 412724
rect 393078 412722 393084 412724
rect 391749 412664 391754 412720
rect 391749 412660 391796 412664
rect 391860 412662 391906 412722
rect 393038 412662 393084 412722
rect 393148 412720 393195 412724
rect 393190 412664 393195 412720
rect 391860 412660 391866 412662
rect 393078 412660 393084 412662
rect 393148 412660 393195 412664
rect 391749 412659 391815 412660
rect 393129 412659 393195 412660
rect 393957 412724 394023 412725
rect 394693 412724 394759 412725
rect 395337 412724 395403 412725
rect 396073 412724 396139 412725
rect 393957 412720 394004 412724
rect 394068 412722 394074 412724
rect 394693 412722 394740 412724
rect 393957 412664 393962 412720
rect 393957 412660 394004 412664
rect 394068 412662 394114 412722
rect 394648 412720 394740 412722
rect 394648 412664 394698 412720
rect 394648 412662 394740 412664
rect 394068 412660 394074 412662
rect 394693 412660 394740 412662
rect 394804 412660 394810 412724
rect 395286 412722 395292 412724
rect 395246 412662 395292 412722
rect 395356 412720 395403 412724
rect 395398 412664 395403 412720
rect 395286 412660 395292 412662
rect 395356 412660 395403 412664
rect 396022 412660 396028 412724
rect 396092 412722 396139 412724
rect 405733 412722 405799 412725
rect 406326 412722 406332 412724
rect 396092 412720 396184 412722
rect 396134 412664 396184 412720
rect 396092 412662 396184 412664
rect 405733 412720 406332 412722
rect 405733 412664 405738 412720
rect 405794 412664 406332 412720
rect 405733 412662 406332 412664
rect 396092 412660 396139 412662
rect 393957 412659 394023 412660
rect 394693 412659 394759 412660
rect 395337 412659 395403 412660
rect 396073 412659 396139 412660
rect 405733 412659 405799 412662
rect 406326 412660 406332 412662
rect 406396 412660 406402 412724
rect 282085 412314 282151 412317
rect 279956 412312 282151 412314
rect 279956 412256 282090 412312
rect 282146 412256 282151 412312
rect 279956 412254 282151 412256
rect 282085 412251 282151 412254
rect 388069 411772 388135 411773
rect 57830 411708 57836 411772
rect 57900 411770 57906 411772
rect 388069 411770 388116 411772
rect 57900 411710 60076 411770
rect 388024 411768 388116 411770
rect 388024 411712 388074 411768
rect 388024 411710 388116 411712
rect 57900 411708 57906 411710
rect 388069 411708 388116 411710
rect 388180 411708 388186 411772
rect 388069 411707 388135 411708
rect 391013 411636 391079 411637
rect 397453 411636 397519 411637
rect 399109 411636 399175 411637
rect 391013 411634 391060 411636
rect 390968 411632 391060 411634
rect 390968 411576 391018 411632
rect 390968 411574 391060 411576
rect 391013 411572 391060 411574
rect 391124 411572 391130 411636
rect 397453 411634 397460 411636
rect 397368 411632 397460 411634
rect 397368 411576 397458 411632
rect 397368 411574 397460 411576
rect 397453 411572 397460 411574
rect 397524 411572 397530 411636
rect 399109 411634 399156 411636
rect 399064 411632 399156 411634
rect 399064 411576 399114 411632
rect 399064 411574 399156 411576
rect 399109 411572 399156 411574
rect 399220 411572 399226 411636
rect 391013 411571 391079 411572
rect 397453 411571 397519 411572
rect 399109 411571 399175 411572
rect 389265 411500 389331 411501
rect 398005 411500 398071 411501
rect 400949 411500 401015 411501
rect 403249 411500 403315 411501
rect 389265 411498 389284 411500
rect 389192 411496 389284 411498
rect 389192 411440 389270 411496
rect 389192 411438 389284 411440
rect 389265 411436 389284 411438
rect 389348 411436 389354 411500
rect 398005 411498 398052 411500
rect 397960 411496 398052 411498
rect 397960 411440 398010 411496
rect 397960 411438 398052 411440
rect 398005 411436 398052 411438
rect 398116 411436 398122 411500
rect 400949 411498 400964 411500
rect 400872 411496 400964 411498
rect 400872 411440 400954 411496
rect 400872 411438 400964 411440
rect 400949 411436 400964 411438
rect 401028 411436 401034 411500
rect 403249 411498 403300 411500
rect 403208 411496 403300 411498
rect 403208 411440 403254 411496
rect 403208 411438 403300 411440
rect 403249 411436 403300 411438
rect 403364 411436 403370 411500
rect 389265 411435 389331 411436
rect 398005 411435 398071 411436
rect 400949 411435 401015 411436
rect 403249 411435 403315 411436
rect 401685 411364 401751 411365
rect 404353 411364 404419 411365
rect 401685 411362 401732 411364
rect 401640 411360 401732 411362
rect 401640 411304 401690 411360
rect 401640 411302 401732 411304
rect 401685 411300 401732 411302
rect 401796 411300 401802 411364
rect 404302 411300 404308 411364
rect 404372 411362 404419 411364
rect 404372 411360 404464 411362
rect 404414 411304 404464 411360
rect 404372 411302 404464 411304
rect 404372 411300 404419 411302
rect 401685 411299 401751 411300
rect 404353 411299 404419 411300
rect 282821 411226 282887 411229
rect 279956 411224 282887 411226
rect 279956 411168 282826 411224
rect 282882 411168 282887 411224
rect 279956 411166 282887 411168
rect 282821 411163 282887 411166
rect 389725 411092 389791 411093
rect 389725 411090 389772 411092
rect 389680 411088 389772 411090
rect 389680 411032 389730 411088
rect 389680 411030 389772 411032
rect 389725 411028 389772 411030
rect 389836 411028 389842 411092
rect 389725 411027 389791 411028
rect 392301 410412 392367 410413
rect 409965 410412 410031 410413
rect 392296 410410 392302 410412
rect 392210 410350 392302 410410
rect 392296 410348 392302 410350
rect 392366 410348 392372 410412
rect 409965 410410 410012 410412
rect 409920 410408 410012 410410
rect 409920 410352 409970 410408
rect 409920 410350 410012 410352
rect 409965 410348 410012 410350
rect 410076 410348 410082 410412
rect 392301 410347 392367 410348
rect 409965 410347 410031 410348
rect 281901 410274 281967 410277
rect 279956 410272 281967 410274
rect 279956 410216 281906 410272
rect 281962 410216 281967 410272
rect 279956 410214 281967 410216
rect 281901 410211 281967 410214
rect 59353 409730 59419 409733
rect 59353 409728 60076 409730
rect 59353 409672 59358 409728
rect 59414 409672 60076 409728
rect 59353 409670 60076 409672
rect 59353 409667 59419 409670
rect -960 409172 480 409412
rect 283005 409322 283071 409325
rect 279956 409320 283071 409322
rect 279956 409264 283010 409320
rect 283066 409264 283071 409320
rect 279956 409262 283071 409264
rect 283005 409259 283071 409262
rect 282913 408506 282979 408509
rect 279926 408504 282979 408506
rect 279926 408448 282918 408504
rect 282974 408448 282979 408504
rect 279926 408446 282979 408448
rect 279926 408204 279986 408446
rect 282913 408443 282979 408446
rect 282453 407962 282519 407965
rect 279926 407960 282519 407962
rect 279926 407904 282458 407960
rect 282514 407904 282519 407960
rect 279926 407902 282519 407904
rect 59486 407764 59492 407828
rect 59556 407826 59562 407828
rect 59556 407766 60076 407826
rect 59556 407764 59562 407766
rect 279926 407252 279986 407902
rect 282453 407899 282519 407902
rect 281809 406194 281875 406197
rect 279956 406192 281875 406194
rect 279956 406136 281814 406192
rect 281870 406136 281875 406192
rect 279956 406134 281875 406136
rect 281809 406131 281875 406134
rect 57646 405860 57652 405924
rect 57716 405922 57722 405924
rect 57716 405862 60076 405922
rect 57716 405860 57722 405862
rect 281717 405242 281783 405245
rect 279956 405240 281783 405242
rect 279956 405184 281722 405240
rect 281778 405184 281783 405240
rect 279956 405182 281783 405184
rect 281717 405179 281783 405182
rect 580625 404834 580691 404837
rect 583520 404834 584960 404924
rect 580625 404832 584960 404834
rect 580625 404776 580630 404832
rect 580686 404776 584960 404832
rect 580625 404774 584960 404776
rect 580625 404771 580691 404774
rect 583520 404684 584960 404774
rect 282821 404290 282887 404293
rect 279956 404288 282887 404290
rect 279956 404232 282826 404288
rect 282882 404232 282887 404288
rect 279956 404230 282887 404232
rect 282821 404227 282887 404230
rect 59118 403956 59124 404020
rect 59188 404018 59194 404020
rect 59188 403958 60076 404018
rect 59188 403956 59194 403958
rect 281901 403202 281967 403205
rect 279956 403200 281967 403202
rect 279956 403144 281906 403200
rect 281962 403144 281967 403200
rect 279956 403142 281967 403144
rect 281901 403139 281967 403142
rect 282177 402250 282243 402253
rect 279956 402248 282243 402250
rect 279956 402192 282182 402248
rect 282238 402192 282243 402248
rect 279956 402190 282243 402192
rect 282177 402187 282243 402190
rect 59302 402052 59308 402116
rect 59372 402114 59378 402116
rect 59372 402054 60076 402114
rect 59372 402052 59378 402054
rect 281625 401162 281691 401165
rect 279956 401160 281691 401162
rect 279956 401104 281630 401160
rect 281686 401104 281691 401160
rect 279956 401102 281691 401104
rect 281625 401099 281691 401102
rect 281625 400210 281691 400213
rect 279956 400208 281691 400210
rect 279956 400152 281630 400208
rect 281686 400152 281691 400208
rect 279956 400150 281691 400152
rect 281625 400147 281691 400150
rect 58065 400074 58131 400077
rect 58065 400072 60076 400074
rect 58065 400016 58070 400072
rect 58126 400016 60076 400072
rect 58065 400014 60076 400016
rect 58065 400011 58131 400014
rect 281625 399122 281691 399125
rect 279956 399120 281691 399122
rect 279956 399064 281630 399120
rect 281686 399064 281691 399120
rect 279956 399062 281691 399064
rect 281625 399059 281691 399062
rect 58198 398108 58204 398172
rect 58268 398170 58274 398172
rect 282177 398170 282243 398173
rect 58268 398110 60076 398170
rect 279956 398168 282243 398170
rect 279956 398112 282182 398168
rect 282238 398112 282243 398168
rect 279956 398110 282243 398112
rect 58268 398108 58274 398110
rect 282177 398107 282243 398110
rect 283598 397218 283604 397220
rect 279956 397158 283604 397218
rect 283598 397156 283604 397158
rect 283668 397156 283674 397220
rect 59721 396266 59787 396269
rect 59721 396264 60076 396266
rect 59721 396208 59726 396264
rect 59782 396208 60076 396264
rect 59721 396206 60076 396208
rect 59721 396203 59787 396206
rect 283782 396130 283788 396132
rect 279956 396070 283788 396130
rect 283782 396068 283788 396070
rect 283852 396068 283858 396132
rect 283414 395178 283420 395180
rect -960 395042 480 395132
rect 279956 395118 283420 395178
rect 283414 395116 283420 395118
rect 283484 395116 283490 395180
rect 3141 395042 3207 395045
rect -960 395040 3207 395042
rect -960 394984 3146 395040
rect 3202 394984 3207 395040
rect -960 394982 3207 394984
rect -960 394892 480 394982
rect 3141 394979 3207 394982
rect 57278 394300 57284 394364
rect 57348 394362 57354 394364
rect 57348 394302 60076 394362
rect 57348 394300 57354 394302
rect 281625 394090 281691 394093
rect 279956 394088 281691 394090
rect 279956 394032 281630 394088
rect 281686 394032 281691 394088
rect 279956 394030 281691 394032
rect 281625 394027 281691 394030
rect 281717 393274 281783 393277
rect 282453 393274 282519 393277
rect 281717 393272 282519 393274
rect 281717 393216 281722 393272
rect 281778 393216 282458 393272
rect 282514 393216 282519 393272
rect 281717 393214 282519 393216
rect 281717 393211 281783 393214
rect 282453 393211 282519 393214
rect 281625 393138 281691 393141
rect 279956 393136 281691 393138
rect 279956 393080 281630 393136
rect 281686 393080 281691 393136
rect 279956 393078 281691 393080
rect 281625 393075 281691 393078
rect 419533 393002 419599 393005
rect 417190 393000 419599 393002
rect 417190 392944 419538 393000
rect 419594 392944 419599 393000
rect 417190 392942 419599 392944
rect 417190 392692 417250 392942
rect 419533 392939 419599 392942
rect 580717 393002 580783 393005
rect 583520 393002 584960 393092
rect 580717 393000 584960 393002
rect 580717 392944 580722 393000
rect 580778 392944 584960 393000
rect 580717 392942 584960 392944
rect 580717 392939 580783 392942
rect 583520 392852 584960 392942
rect 58157 392458 58223 392461
rect 58157 392456 60076 392458
rect 58157 392400 58162 392456
rect 58218 392400 60076 392456
rect 58157 392398 60076 392400
rect 58157 392395 58223 392398
rect 281625 392050 281691 392053
rect 279956 392048 281691 392050
rect 279956 391992 281630 392048
rect 281686 391992 281691 392048
rect 279956 391990 281691 391992
rect 281625 391987 281691 391990
rect 282310 391098 282316 391100
rect 279956 391038 282316 391098
rect 282310 391036 282316 391038
rect 282380 391036 282386 391100
rect 417190 390690 417250 390992
rect 419533 390690 419599 390693
rect 417190 390688 419599 390690
rect 417190 390632 419538 390688
rect 419594 390632 419599 390688
rect 417190 390630 419599 390632
rect 419533 390627 419599 390630
rect 59629 390418 59695 390421
rect 59629 390416 60076 390418
rect 59629 390360 59634 390416
rect 59690 390360 60076 390416
rect 59629 390358 60076 390360
rect 59629 390355 59695 390358
rect 281901 390146 281967 390149
rect 279956 390144 281967 390146
rect 279956 390088 281906 390144
rect 281962 390088 281967 390144
rect 279956 390086 281967 390088
rect 281901 390083 281967 390086
rect 338021 389874 338087 389877
rect 340094 389874 340154 390319
rect 338021 389872 340154 389874
rect 338021 389816 338026 389872
rect 338082 389816 340154 389872
rect 338021 389814 340154 389816
rect 338021 389811 338087 389814
rect 282821 389058 282887 389061
rect 279956 389056 282887 389058
rect 279956 389000 282826 389056
rect 282882 389000 282887 389056
rect 279956 388998 282887 389000
rect 282821 388995 282887 388998
rect 57462 388452 57468 388516
rect 57532 388514 57538 388516
rect 57532 388454 60076 388514
rect 57532 388452 57538 388454
rect 281625 388106 281691 388109
rect 279956 388104 281691 388106
rect 279956 388048 281630 388104
rect 281686 388048 281691 388104
rect 279956 388046 281691 388048
rect 281625 388043 281691 388046
rect 281625 387018 281691 387021
rect 279956 387016 281691 387018
rect 279956 386960 281630 387016
rect 281686 386960 281691 387016
rect 279956 386958 281691 386960
rect 281625 386955 281691 386958
rect 58249 386610 58315 386613
rect 58249 386608 60076 386610
rect 58249 386552 58254 386608
rect 58310 386552 60076 386608
rect 58249 386550 60076 386552
rect 58249 386547 58315 386550
rect 281717 386066 281783 386069
rect 279956 386064 281783 386066
rect 279956 386008 281722 386064
rect 281778 386008 281783 386064
rect 279956 386006 281783 386008
rect 281717 386003 281783 386006
rect 281625 385114 281691 385117
rect 279956 385112 281691 385114
rect 279956 385056 281630 385112
rect 281686 385056 281691 385112
rect 279956 385054 281691 385056
rect 281625 385051 281691 385054
rect 59537 384706 59603 384709
rect 59537 384704 60076 384706
rect 59537 384648 59542 384704
rect 59598 384648 60076 384704
rect 59537 384646 60076 384648
rect 59537 384643 59603 384646
rect 281625 384026 281691 384029
rect 279956 384024 281691 384026
rect 279956 383968 281630 384024
rect 281686 383968 281691 384024
rect 279956 383966 281691 383968
rect 281625 383963 281691 383966
rect 282821 383074 282887 383077
rect 279956 383072 282887 383074
rect 279956 383016 282826 383072
rect 282882 383016 282887 383072
rect 279956 383014 282887 383016
rect 282821 383011 282887 383014
rect 57145 382802 57211 382805
rect 57145 382800 60076 382802
rect 57145 382744 57150 382800
rect 57206 382744 60076 382800
rect 57145 382742 60076 382744
rect 57145 382739 57211 382742
rect 281625 381986 281691 381989
rect 279956 381984 281691 381986
rect 279956 381928 281630 381984
rect 281686 381928 281691 381984
rect 279956 381926 281691 381928
rect 281625 381923 281691 381926
rect 337377 381306 337443 381309
rect 340094 381306 340154 389814
rect 337377 381304 340154 381306
rect 337377 381248 337382 381304
rect 337438 381248 340154 381304
rect 337377 381246 340154 381248
rect 337377 381243 337443 381246
rect 583520 381156 584960 381396
rect 281717 381034 281783 381037
rect 279956 381032 281783 381034
rect 279956 380976 281722 381032
rect 281778 380976 281783 381032
rect 279956 380974 281783 380976
rect 281717 380971 281783 380974
rect 57513 380762 57579 380765
rect 57513 380760 60076 380762
rect -960 380626 480 380716
rect 57513 380704 57518 380760
rect 57574 380704 60076 380760
rect 57513 380702 60076 380704
rect 57513 380699 57579 380702
rect 3233 380626 3299 380629
rect -960 380624 3299 380626
rect -960 380568 3238 380624
rect 3294 380568 3299 380624
rect -960 380566 3299 380568
rect -960 380476 480 380566
rect 3233 380563 3299 380566
rect 282821 379946 282887 379949
rect 279956 379944 282887 379946
rect 279956 379888 282826 379944
rect 282882 379888 282887 379944
rect 279956 379886 282887 379888
rect 282821 379883 282887 379886
rect 282821 378994 282887 378997
rect 279956 378992 282887 378994
rect 279956 378936 282826 378992
rect 282882 378936 282887 378992
rect 279956 378934 282887 378936
rect 282821 378931 282887 378934
rect 57605 378858 57671 378861
rect 57605 378856 60076 378858
rect 57605 378800 57610 378856
rect 57666 378800 60076 378856
rect 57605 378798 60076 378800
rect 57605 378795 57671 378798
rect 282821 378042 282887 378045
rect 279956 378040 282887 378042
rect 279956 377984 282826 378040
rect 282882 377984 282887 378040
rect 279956 377982 282887 377984
rect 282821 377979 282887 377982
rect 57789 376954 57855 376957
rect 282177 376954 282243 376957
rect 57789 376952 60076 376954
rect 57789 376896 57794 376952
rect 57850 376896 60076 376952
rect 57789 376894 60076 376896
rect 279956 376952 282243 376954
rect 279956 376896 282182 376952
rect 282238 376896 282243 376952
rect 279956 376894 282243 376896
rect 57789 376891 57855 376894
rect 282177 376891 282243 376894
rect 282821 376002 282887 376005
rect 279956 376000 282887 376002
rect 279956 375944 282826 376000
rect 282882 375944 282887 376000
rect 279956 375942 282887 375944
rect 282821 375939 282887 375942
rect 57830 374988 57836 375052
rect 57900 375050 57906 375052
rect 57900 374990 60076 375050
rect 57900 374988 57906 374990
rect 282821 374914 282887 374917
rect 279956 374912 282887 374914
rect 279956 374856 282826 374912
rect 282882 374856 282887 374912
rect 279956 374854 282887 374856
rect 282821 374851 282887 374854
rect 282821 373962 282887 373965
rect 279956 373960 282887 373962
rect 279956 373904 282826 373960
rect 282882 373904 282887 373960
rect 279956 373902 282887 373904
rect 282821 373899 282887 373902
rect 57697 373146 57763 373149
rect 57697 373144 60076 373146
rect 57697 373088 57702 373144
rect 57758 373088 60076 373144
rect 57697 373086 60076 373088
rect 57697 373083 57763 373086
rect 282177 372874 282243 372877
rect 279956 372872 282243 372874
rect 279956 372816 282182 372872
rect 282238 372816 282243 372872
rect 279956 372814 282243 372816
rect 282177 372811 282243 372814
rect 282821 371922 282887 371925
rect 279956 371920 282887 371922
rect 279956 371864 282826 371920
rect 282882 371864 282887 371920
rect 279956 371862 282887 371864
rect 282821 371859 282887 371862
rect 56961 371242 57027 371245
rect 56961 371240 60076 371242
rect 56961 371184 56966 371240
rect 57022 371184 60076 371240
rect 56961 371182 60076 371184
rect 56961 371179 57027 371182
rect 282821 370970 282887 370973
rect 279956 370968 282887 370970
rect 279956 370912 282826 370968
rect 282882 370912 282887 370968
rect 279956 370910 282887 370912
rect 282821 370907 282887 370910
rect 282177 369882 282243 369885
rect 279956 369880 282243 369882
rect 279956 369824 282182 369880
rect 282238 369824 282243 369880
rect 279956 369822 282243 369824
rect 282177 369819 282243 369822
rect 580809 369610 580875 369613
rect 583520 369610 584960 369700
rect 580809 369608 584960 369610
rect 580809 369552 580814 369608
rect 580870 369552 584960 369608
rect 580809 369550 584960 369552
rect 580809 369547 580875 369550
rect 583520 369460 584960 369550
rect 57881 369202 57947 369205
rect 57881 369200 60076 369202
rect 57881 369144 57886 369200
rect 57942 369144 60076 369200
rect 57881 369142 60076 369144
rect 57881 369139 57947 369142
rect 282821 368930 282887 368933
rect 279956 368928 282887 368930
rect 279956 368872 282826 368928
rect 282882 368872 282887 368928
rect 279956 368870 282887 368872
rect 282821 368867 282887 368870
rect 282821 367842 282887 367845
rect 279956 367840 282887 367842
rect 279956 367784 282826 367840
rect 282882 367784 282887 367840
rect 279956 367782 282887 367784
rect 282821 367779 282887 367782
rect 57605 367298 57671 367301
rect 57605 367296 60076 367298
rect 57605 367240 57610 367296
rect 57666 367240 60076 367296
rect 57605 367238 60076 367240
rect 57605 367235 57671 367238
rect 282821 366890 282887 366893
rect 279956 366888 282887 366890
rect 279956 366832 282826 366888
rect 282882 366832 282887 366888
rect 279956 366830 282887 366832
rect 282821 366827 282887 366830
rect -960 366210 480 366300
rect 3141 366210 3207 366213
rect -960 366208 3207 366210
rect -960 366152 3146 366208
rect 3202 366152 3207 366208
rect -960 366150 3207 366152
rect -960 366060 480 366150
rect 3141 366147 3207 366150
rect 282177 365802 282243 365805
rect 279956 365800 282243 365802
rect 279956 365744 282182 365800
rect 282238 365744 282243 365800
rect 279956 365742 282243 365744
rect 282177 365739 282243 365742
rect 57053 365394 57119 365397
rect 57053 365392 60076 365394
rect 57053 365336 57058 365392
rect 57114 365336 60076 365392
rect 57053 365334 60076 365336
rect 57053 365331 57119 365334
rect 282821 364850 282887 364853
rect 279956 364848 282887 364850
rect 279956 364792 282826 364848
rect 282882 364792 282887 364848
rect 279956 364790 282887 364792
rect 282821 364787 282887 364790
rect 282821 363898 282887 363901
rect 279956 363896 282887 363898
rect 279956 363840 282826 363896
rect 282882 363840 282887 363896
rect 279956 363838 282887 363840
rect 282821 363835 282887 363838
rect 57513 363490 57579 363493
rect 57513 363488 60076 363490
rect 57513 363432 57518 363488
rect 57574 363432 60076 363488
rect 57513 363430 60076 363432
rect 57513 363427 57579 363430
rect 282821 362810 282887 362813
rect 279956 362808 282887 362810
rect 279956 362752 282826 362808
rect 282882 362752 282887 362808
rect 279956 362750 282887 362752
rect 282821 362747 282887 362750
rect 282729 361858 282795 361861
rect 279956 361856 282795 361858
rect 279956 361800 282734 361856
rect 282790 361800 282795 361856
rect 279956 361798 282795 361800
rect 282729 361795 282795 361798
rect 56869 361586 56935 361589
rect 56869 361584 60076 361586
rect 56869 361528 56874 361584
rect 56930 361528 60076 361584
rect 56869 361526 60076 361528
rect 56869 361523 56935 361526
rect 281717 360770 281783 360773
rect 279956 360768 281783 360770
rect 279956 360712 281722 360768
rect 281778 360712 281783 360768
rect 279956 360710 281783 360712
rect 281717 360707 281783 360710
rect 282821 359818 282887 359821
rect 279956 359816 282887 359818
rect 279956 359760 282826 359816
rect 282882 359760 282887 359816
rect 279956 359758 282887 359760
rect 282821 359755 282887 359758
rect 56685 359546 56751 359549
rect 56685 359544 60076 359546
rect 56685 359488 56690 359544
rect 56746 359488 60076 359544
rect 56685 359486 60076 359488
rect 56685 359483 56751 359486
rect 282729 358866 282795 358869
rect 279956 358864 282795 358866
rect 279956 358808 282734 358864
rect 282790 358808 282795 358864
rect 279956 358806 282795 358808
rect 282729 358803 282795 358806
rect 580901 357914 580967 357917
rect 583520 357914 584960 358004
rect 580901 357912 584960 357914
rect 580901 357856 580906 357912
rect 580962 357856 584960 357912
rect 580901 357854 584960 357856
rect 580901 357851 580967 357854
rect 281901 357778 281967 357781
rect 279956 357776 281967 357778
rect 279956 357720 281906 357776
rect 281962 357720 281967 357776
rect 583520 357764 584960 357854
rect 279956 357718 281967 357720
rect 281901 357715 281967 357718
rect 56593 357642 56659 357645
rect 56593 357640 60076 357642
rect 56593 357584 56598 357640
rect 56654 357584 60076 357640
rect 56593 357582 60076 357584
rect 56593 357579 56659 357582
rect 281993 356826 282059 356829
rect 279956 356824 282059 356826
rect 279956 356768 281998 356824
rect 282054 356768 282059 356824
rect 279956 356766 282059 356768
rect 281993 356763 282059 356766
rect 56777 355738 56843 355741
rect 282085 355738 282151 355741
rect 56777 355736 60076 355738
rect 56777 355680 56782 355736
rect 56838 355680 60076 355736
rect 56777 355678 60076 355680
rect 279956 355736 282151 355738
rect 279956 355680 282090 355736
rect 282146 355680 282151 355736
rect 279956 355678 282151 355680
rect 56777 355675 56843 355678
rect 282085 355675 282151 355678
rect 282177 354786 282243 354789
rect 279956 354784 282243 354786
rect 279956 354728 282182 354784
rect 282238 354728 282243 354784
rect 279956 354726 282243 354728
rect 282177 354723 282243 354726
rect 281993 354650 282059 354653
rect 282361 354650 282427 354653
rect 281993 354648 282427 354650
rect 281993 354592 281998 354648
rect 282054 354592 282366 354648
rect 282422 354592 282427 354648
rect 281993 354590 282427 354592
rect 281993 354587 282059 354590
rect 282361 354587 282427 354590
rect 56910 353772 56916 353836
rect 56980 353834 56986 353836
rect 56980 353774 60076 353834
rect 56980 353772 56986 353774
rect 282637 353698 282703 353701
rect 279956 353696 282703 353698
rect 279956 353640 282642 353696
rect 282698 353640 282703 353696
rect 279956 353638 282703 353640
rect 282637 353635 282703 353638
rect 282085 352746 282151 352749
rect 279956 352744 282151 352746
rect 279956 352688 282090 352744
rect 282146 352688 282151 352744
rect 279956 352686 282151 352688
rect 282085 352683 282151 352686
rect -960 351780 480 352020
rect 57145 351930 57211 351933
rect 57145 351928 60076 351930
rect 57145 351872 57150 351928
rect 57206 351872 60076 351928
rect 57145 351870 60076 351872
rect 57145 351867 57211 351870
rect 281993 351794 282059 351797
rect 279956 351792 282059 351794
rect 279956 351736 281998 351792
rect 282054 351736 282059 351792
rect 279956 351734 282059 351736
rect 281993 351731 282059 351734
rect 282545 350706 282611 350709
rect 279956 350704 282611 350706
rect 279956 350648 282550 350704
rect 282606 350648 282611 350704
rect 279956 350646 282611 350648
rect 282545 350643 282611 350646
rect 59445 349890 59511 349893
rect 59445 349888 60076 349890
rect 59445 349832 59450 349888
rect 59506 349832 60076 349888
rect 59445 349830 60076 349832
rect 59445 349827 59511 349830
rect 282269 349754 282335 349757
rect 279956 349752 282335 349754
rect 279956 349696 282274 349752
rect 282330 349696 282335 349752
rect 279956 349694 282335 349696
rect 282269 349691 282335 349694
rect 282821 348666 282887 348669
rect 279956 348664 282887 348666
rect 279956 348608 282826 348664
rect 282882 348608 282887 348664
rect 279956 348606 282887 348608
rect 282821 348603 282887 348606
rect 57278 347924 57284 347988
rect 57348 347986 57354 347988
rect 57348 347926 60076 347986
rect 57348 347924 57354 347926
rect 282821 347714 282887 347717
rect 279956 347712 282887 347714
rect 279956 347656 282826 347712
rect 282882 347656 282887 347712
rect 279956 347654 282887 347656
rect 282821 347651 282887 347654
rect 282269 346626 282335 346629
rect 279956 346624 282335 346626
rect 279956 346568 282274 346624
rect 282330 346568 282335 346624
rect 279956 346566 282335 346568
rect 282269 346563 282335 346566
rect 57094 346020 57100 346084
rect 57164 346082 57170 346084
rect 580165 346082 580231 346085
rect 583520 346082 584960 346172
rect 57164 346022 60076 346082
rect 580165 346080 584960 346082
rect 580165 346024 580170 346080
rect 580226 346024 584960 346080
rect 580165 346022 584960 346024
rect 57164 346020 57170 346022
rect 580165 346019 580231 346022
rect 583520 345932 584960 346022
rect 282085 345674 282151 345677
rect 279956 345672 282151 345674
rect 279956 345616 282090 345672
rect 282146 345616 282151 345672
rect 279956 345614 282151 345616
rect 282085 345611 282151 345614
rect 282821 344722 282887 344725
rect 279956 344720 282887 344722
rect 279956 344664 282826 344720
rect 282882 344664 282887 344720
rect 279956 344662 282887 344664
rect 282821 344659 282887 344662
rect 59353 344178 59419 344181
rect 59353 344176 60076 344178
rect 59353 344120 59358 344176
rect 59414 344120 60076 344176
rect 59353 344118 60076 344120
rect 59353 344115 59419 344118
rect 282729 343634 282795 343637
rect 279956 343632 282795 343634
rect 279956 343576 282734 343632
rect 282790 343576 282795 343632
rect 279956 343574 282795 343576
rect 282729 343571 282795 343574
rect 282545 342682 282611 342685
rect 279956 342680 282611 342682
rect 279956 342624 282550 342680
rect 282606 342624 282611 342680
rect 279956 342622 282611 342624
rect 282545 342619 282611 342622
rect 57646 342212 57652 342276
rect 57716 342274 57722 342276
rect 57716 342214 60076 342274
rect 57716 342212 57722 342214
rect 282821 341594 282887 341597
rect 279956 341592 282887 341594
rect 279956 341536 282826 341592
rect 282882 341536 282887 341592
rect 279956 341534 282887 341536
rect 282821 341531 282887 341534
rect 282453 340642 282519 340645
rect 279956 340640 282519 340642
rect 279956 340584 282458 340640
rect 282514 340584 282519 340640
rect 279956 340582 282519 340584
rect 282453 340579 282519 340582
rect 57462 340172 57468 340236
rect 57532 340234 57538 340236
rect 57532 340174 60076 340234
rect 57532 340172 57538 340174
rect 282085 339690 282151 339693
rect 279956 339688 282151 339690
rect 279956 339632 282090 339688
rect 282146 339632 282151 339688
rect 279956 339630 282151 339632
rect 282085 339627 282151 339630
rect 282361 338602 282427 338605
rect 279956 338600 282427 338602
rect 279956 338544 282366 338600
rect 282422 338544 282427 338600
rect 279956 338542 282427 338544
rect 282361 338539 282427 338542
rect 59077 338330 59143 338333
rect 59077 338328 60076 338330
rect 59077 338272 59082 338328
rect 59138 338272 60076 338328
rect 59077 338270 60076 338272
rect 59077 338267 59143 338270
rect 282545 337650 282611 337653
rect 279956 337648 282611 337650
rect -960 337514 480 337604
rect 279956 337592 282550 337648
rect 282606 337592 282611 337648
rect 279956 337590 282611 337592
rect 282545 337587 282611 337590
rect 3417 337514 3483 337517
rect -960 337512 3483 337514
rect -960 337456 3422 337512
rect 3478 337456 3483 337512
rect -960 337454 3483 337456
rect -960 337364 480 337454
rect 3417 337451 3483 337454
rect 281993 336562 282059 336565
rect 279956 336560 282059 336562
rect 279956 336504 281998 336560
rect 282054 336504 282059 336560
rect 279956 336502 282059 336504
rect 281993 336499 282059 336502
rect 57789 336426 57855 336429
rect 57789 336424 60076 336426
rect 57789 336368 57794 336424
rect 57850 336368 60076 336424
rect 57789 336366 60076 336368
rect 57789 336363 57855 336366
rect 282637 335610 282703 335613
rect 279956 335608 282703 335610
rect 279956 335552 282642 335608
rect 282698 335552 282703 335608
rect 279956 335550 282703 335552
rect 282637 335547 282703 335550
rect 57421 334522 57487 334525
rect 281809 334522 281875 334525
rect 57421 334520 60076 334522
rect 57421 334464 57426 334520
rect 57482 334464 60076 334520
rect 57421 334462 60076 334464
rect 279956 334520 281875 334522
rect 279956 334464 281814 334520
rect 281870 334464 281875 334520
rect 279956 334462 281875 334464
rect 57421 334459 57487 334462
rect 281809 334459 281875 334462
rect 583520 334236 584960 334476
rect 281625 333570 281691 333573
rect 279956 333568 281691 333570
rect 279956 333512 281630 333568
rect 281686 333512 281691 333568
rect 279956 333510 281691 333512
rect 281625 333507 281691 333510
rect 59169 332618 59235 332621
rect 282177 332618 282243 332621
rect 59169 332616 60076 332618
rect 59169 332560 59174 332616
rect 59230 332560 60076 332616
rect 59169 332558 60076 332560
rect 279956 332616 282243 332618
rect 279956 332560 282182 332616
rect 282238 332560 282243 332616
rect 279956 332558 282243 332560
rect 417190 332618 417250 333144
rect 419901 332618 419967 332621
rect 417190 332616 419967 332618
rect 417190 332560 419906 332616
rect 419962 332560 419967 332616
rect 417190 332558 419967 332560
rect 59169 332555 59235 332558
rect 282177 332555 282243 332558
rect 419901 332555 419967 332558
rect 281901 331530 281967 331533
rect 279956 331528 281967 331530
rect 279956 331472 281906 331528
rect 281962 331472 281967 331528
rect 279956 331470 281967 331472
rect 281901 331467 281967 331470
rect 417190 331258 417250 331444
rect 420177 331258 420243 331261
rect 417190 331256 420243 331258
rect 417190 331200 420182 331256
rect 420238 331200 420243 331256
rect 417190 331198 420243 331200
rect 420177 331195 420243 331198
rect 57830 330652 57836 330716
rect 57900 330714 57906 330716
rect 59721 330714 59787 330717
rect 57900 330712 59787 330714
rect 57900 330656 59726 330712
rect 59782 330656 59787 330712
rect 57900 330654 59787 330656
rect 57900 330652 57906 330654
rect 59721 330651 59787 330654
rect 57830 330516 57836 330580
rect 57900 330578 57906 330580
rect 281625 330578 281691 330581
rect 57900 330518 60076 330578
rect 279956 330576 281691 330578
rect 279956 330520 281630 330576
rect 281686 330520 281691 330576
rect 279956 330518 281691 330520
rect 57900 330516 57906 330518
rect 281625 330515 281691 330518
rect 417190 329898 417250 330316
rect 419993 329898 420059 329901
rect 417190 329896 420059 329898
rect 417190 329840 419998 329896
rect 420054 329840 420059 329896
rect 417190 329838 420059 329840
rect 419993 329835 420059 329838
rect 281533 329490 281599 329493
rect 279956 329488 281599 329490
rect 279956 329432 281538 329488
rect 281594 329432 281599 329488
rect 279956 329430 281599 329432
rect 281533 329427 281599 329430
rect 57053 328674 57119 328677
rect 419809 328674 419875 328677
rect 57053 328672 60076 328674
rect 57053 328616 57058 328672
rect 57114 328616 60076 328672
rect 57053 328614 60076 328616
rect 417190 328672 419875 328674
rect 417190 328616 419814 328672
rect 419870 328616 419875 328672
rect 417190 328614 419875 328616
rect 57053 328611 57119 328614
rect 419809 328611 419875 328614
rect 281625 328538 281691 328541
rect 279956 328536 281691 328538
rect 279956 328480 281630 328536
rect 281686 328480 281691 328536
rect 279956 328478 281691 328480
rect 281625 328475 281691 328478
rect 281533 327450 281599 327453
rect 279956 327448 281599 327450
rect 279956 327392 281538 327448
rect 281594 327392 281599 327448
rect 279956 327390 281599 327392
rect 281533 327387 281599 327390
rect 417190 327178 417250 327488
rect 419717 327178 419783 327181
rect 417190 327176 419783 327178
rect 417190 327120 419722 327176
rect 419778 327120 419783 327176
rect 417190 327118 419783 327120
rect 419717 327115 419783 327118
rect 59261 326770 59327 326773
rect 59261 326768 60076 326770
rect 59261 326712 59266 326768
rect 59322 326712 60076 326768
rect 59261 326710 60076 326712
rect 59261 326707 59327 326710
rect 281533 326498 281599 326501
rect 279956 326496 281599 326498
rect 279956 326440 281538 326496
rect 281594 326440 281599 326496
rect 279956 326438 281599 326440
rect 281533 326435 281599 326438
rect 419625 325818 419691 325821
rect 417220 325816 419691 325818
rect 417220 325760 419630 325816
rect 419686 325760 419691 325816
rect 417220 325758 419691 325760
rect 419625 325755 419691 325758
rect 281717 325546 281783 325549
rect 279956 325544 281783 325546
rect 279956 325488 281722 325544
rect 281778 325488 281783 325544
rect 279956 325486 281783 325488
rect 281717 325483 281783 325486
rect 57789 324866 57855 324869
rect 57789 324864 60076 324866
rect 57789 324808 57794 324864
rect 57850 324808 60076 324864
rect 57789 324806 60076 324808
rect 57789 324803 57855 324806
rect 281533 324458 281599 324461
rect 279956 324456 281599 324458
rect 279956 324400 281538 324456
rect 281594 324400 281599 324456
rect 279956 324398 281599 324400
rect 281533 324395 281599 324398
rect 416454 324053 416514 324660
rect 416405 324048 416514 324053
rect 416405 323992 416410 324048
rect 416466 323992 416514 324048
rect 416405 323990 416514 323992
rect 416405 323987 416471 323990
rect 281533 323506 281599 323509
rect 279956 323504 281599 323506
rect 279956 323448 281538 323504
rect 281594 323448 281599 323504
rect 279956 323446 281599 323448
rect 281533 323443 281599 323446
rect -960 323098 480 323188
rect 3233 323098 3299 323101
rect -960 323096 3299 323098
rect -960 323040 3238 323096
rect 3294 323040 3299 323096
rect -960 323038 3299 323040
rect -960 322948 480 323038
rect 3233 323035 3299 323038
rect 57697 322962 57763 322965
rect 57697 322960 60076 322962
rect 57697 322904 57702 322960
rect 57758 322904 60076 322960
rect 57697 322902 60076 322904
rect 57697 322899 57763 322902
rect 579981 322690 580047 322693
rect 583520 322690 584960 322780
rect 579981 322688 584960 322690
rect 579981 322632 579986 322688
rect 580042 322632 584960 322688
rect 579981 322630 584960 322632
rect 579981 322627 580047 322630
rect 583520 322540 584960 322630
rect 281533 322418 281599 322421
rect 279956 322416 281599 322418
rect 279956 322360 281538 322416
rect 281594 322360 281599 322416
rect 279956 322358 281599 322360
rect 281533 322355 281599 322358
rect 337745 322010 337811 322013
rect 337745 322008 340154 322010
rect 337745 321952 337750 322008
rect 337806 321952 340154 322008
rect 337745 321950 340154 321952
rect 337745 321947 337811 321950
rect 340094 321564 340154 321950
rect 282821 321466 282887 321469
rect 279956 321464 282887 321466
rect 279956 321408 282826 321464
rect 282882 321408 282887 321464
rect 279956 321406 282887 321408
rect 282821 321403 282887 321406
rect 57881 321058 57947 321061
rect 57881 321056 60076 321058
rect 57881 321000 57886 321056
rect 57942 321000 60076 321056
rect 57881 320998 60076 321000
rect 57881 320995 57947 320998
rect 279969 320922 280035 320925
rect 580533 320922 580599 320925
rect 279969 320920 339970 320922
rect 279969 320864 279974 320920
rect 280030 320864 339970 320920
rect 279969 320862 339970 320864
rect 279969 320859 280035 320862
rect 282821 320786 282887 320789
rect 279926 320784 282887 320786
rect 279926 320728 282826 320784
rect 282882 320728 282887 320784
rect 279926 320726 282887 320728
rect 279926 320484 279986 320726
rect 282821 320723 282887 320726
rect 280061 320650 280127 320653
rect 339769 320650 339835 320653
rect 280061 320648 339835 320650
rect 280061 320592 280066 320648
rect 280122 320592 339774 320648
rect 339830 320592 339835 320648
rect 280061 320590 339835 320592
rect 339910 320650 339970 320862
rect 349662 320920 580599 320922
rect 349662 320864 580538 320920
rect 580594 320864 580599 320920
rect 349662 320862 580599 320864
rect 349662 320650 349722 320862
rect 580533 320859 580599 320862
rect 339910 320590 349722 320650
rect 349981 320650 350047 320653
rect 579981 320650 580047 320653
rect 349981 320648 580047 320650
rect 349981 320592 349986 320648
rect 350042 320592 579986 320648
rect 580042 320592 580047 320648
rect 349981 320590 580047 320592
rect 280061 320587 280127 320590
rect 339769 320587 339835 320590
rect 349981 320587 350047 320590
rect 579981 320587 580047 320590
rect 280061 320514 280127 320517
rect 580257 320514 580323 320517
rect 280061 320512 580323 320514
rect 280061 320456 280066 320512
rect 280122 320456 580262 320512
rect 580318 320456 580323 320512
rect 280061 320454 580323 320456
rect 280061 320451 280127 320454
rect 580257 320451 580323 320454
rect 339769 320378 339835 320381
rect 349981 320378 350047 320381
rect 339769 320376 350047 320378
rect 339769 320320 339774 320376
rect 339830 320320 349986 320376
rect 350042 320320 350047 320376
rect 339769 320318 350047 320320
rect 339769 320315 339835 320318
rect 349981 320315 350047 320318
rect 344001 318748 344067 318749
rect 343950 318746 343956 318748
rect 343910 318686 343956 318746
rect 344020 318744 344067 318748
rect 344062 318688 344067 318744
rect 343950 318684 343956 318686
rect 344020 318684 344067 318688
rect 344001 318683 344067 318684
rect 347773 318474 347839 318477
rect 347998 318474 348004 318476
rect 347773 318472 348004 318474
rect 347773 318416 347778 318472
rect 347834 318416 348004 318472
rect 347773 318414 348004 318416
rect 347773 318411 347839 318414
rect 347998 318412 348004 318414
rect 348068 318412 348074 318476
rect 115841 318338 115907 318341
rect 247769 318338 247835 318341
rect 115841 318336 247835 318338
rect 115841 318280 115846 318336
rect 115902 318280 247774 318336
rect 247830 318280 247835 318336
rect 115841 318278 247835 318280
rect 115841 318275 115907 318278
rect 247769 318275 247835 318278
rect 121361 318202 121427 318205
rect 257521 318202 257587 318205
rect 121361 318200 257587 318202
rect 121361 318144 121366 318200
rect 121422 318144 257526 318200
rect 257582 318144 257587 318200
rect 121361 318142 257587 318144
rect 121361 318139 121427 318142
rect 257521 318139 257587 318142
rect 122741 318066 122807 318069
rect 259453 318066 259519 318069
rect 122741 318064 259519 318066
rect 122741 318008 122746 318064
rect 122802 318008 259458 318064
rect 259514 318008 259519 318064
rect 122741 318006 259519 318008
rect 122741 318003 122807 318006
rect 259453 318003 259519 318006
rect 61377 317386 61443 317389
rect 281574 317386 281580 317388
rect 61377 317384 281580 317386
rect 61377 317328 61382 317384
rect 61438 317328 281580 317384
rect 61377 317326 281580 317328
rect 61377 317323 61443 317326
rect 281574 317324 281580 317326
rect 281644 317324 281650 317388
rect 580165 310858 580231 310861
rect 583520 310858 584960 310948
rect 580165 310856 584960 310858
rect 580165 310800 580170 310856
rect 580226 310800 584960 310856
rect 580165 310798 584960 310800
rect 580165 310795 580231 310798
rect 583520 310708 584960 310798
rect -960 308818 480 308908
rect 3325 308818 3391 308821
rect -960 308816 3391 308818
rect -960 308760 3330 308816
rect 3386 308760 3391 308816
rect -960 308758 3391 308760
rect -960 308668 480 308758
rect 3325 308755 3391 308758
rect 579797 299162 579863 299165
rect 583520 299162 584960 299252
rect 579797 299160 584960 299162
rect 579797 299104 579802 299160
rect 579858 299104 584960 299160
rect 579797 299102 584960 299104
rect 579797 299099 579863 299102
rect 583520 299012 584960 299102
rect -960 294402 480 294492
rect 3417 294402 3483 294405
rect -960 294400 3483 294402
rect -960 294344 3422 294400
rect 3478 294344 3483 294400
rect -960 294342 3483 294344
rect -960 294252 480 294342
rect 3417 294339 3483 294342
rect 583520 287316 584960 287556
rect -960 280122 480 280212
rect 3417 280122 3483 280125
rect -960 280120 3483 280122
rect -960 280064 3422 280120
rect 3478 280064 3483 280120
rect -960 280062 3483 280064
rect -960 279972 480 280062
rect 3417 280059 3483 280062
rect 74257 278762 74323 278765
rect 74441 278762 74507 278765
rect 74257 278760 74507 278762
rect 74257 278704 74262 278760
rect 74318 278704 74446 278760
rect 74502 278704 74507 278760
rect 74257 278702 74507 278704
rect 74257 278699 74323 278702
rect 74441 278699 74507 278702
rect 580165 275770 580231 275773
rect 583520 275770 584960 275860
rect 580165 275768 584960 275770
rect 580165 275712 580170 275768
rect 580226 275712 584960 275768
rect 580165 275710 584960 275712
rect 580165 275707 580231 275710
rect 583520 275620 584960 275710
rect -960 265706 480 265796
rect 2865 265706 2931 265709
rect -960 265704 2931 265706
rect -960 265648 2870 265704
rect 2926 265648 2931 265704
rect -960 265646 2931 265648
rect -960 265556 480 265646
rect 2865 265643 2931 265646
rect 106222 264284 106228 264348
rect 106292 264346 106298 264348
rect 111057 264346 111123 264349
rect 106292 264344 111123 264346
rect 106292 264288 111062 264344
rect 111118 264288 111123 264344
rect 106292 264286 111123 264288
rect 106292 264284 106298 264286
rect 111057 264283 111123 264286
rect 125542 264148 125548 264212
rect 125612 264210 125618 264212
rect 135161 264210 135227 264213
rect 125612 264208 135227 264210
rect 125612 264152 135166 264208
rect 135222 264152 135227 264208
rect 125612 264150 135227 264152
rect 125612 264148 125618 264150
rect 135161 264147 135227 264150
rect 86902 264012 86908 264076
rect 86972 264074 86978 264076
rect 96470 264074 96476 264076
rect 86972 264014 96476 264074
rect 86972 264012 86978 264014
rect 96470 264012 96476 264014
rect 96540 264012 96546 264076
rect 106222 264074 106228 264076
rect 99422 264014 106228 264074
rect 56910 263876 56916 263940
rect 56980 263938 56986 263940
rect 56980 263878 64890 263938
rect 56980 263876 56986 263878
rect 64830 263666 64890 263878
rect 70350 263878 82186 263938
rect 70350 263666 70410 263878
rect 64830 263606 70410 263666
rect 82126 263666 82186 263878
rect 96470 263740 96476 263804
rect 96540 263802 96546 263804
rect 99422 263802 99482 264014
rect 106222 264012 106228 264014
rect 106292 264012 106298 264076
rect 140037 264074 140103 264077
rect 135302 264072 140103 264074
rect 135302 264016 140042 264072
rect 140098 264016 140103 264072
rect 135302 264014 140103 264016
rect 118785 263938 118851 263941
rect 125542 263938 125548 263940
rect 118785 263936 125548 263938
rect 118785 263880 118790 263936
rect 118846 263880 125548 263936
rect 118785 263878 125548 263880
rect 118785 263875 118851 263878
rect 125542 263876 125548 263878
rect 125612 263876 125618 263940
rect 96540 263742 99482 263802
rect 135161 263802 135227 263805
rect 135302 263802 135362 264014
rect 140037 264011 140103 264014
rect 154481 263938 154547 263941
rect 583520 263938 584960 264028
rect 154481 263936 161490 263938
rect 154481 263880 154486 263936
rect 154542 263880 161490 263936
rect 154481 263878 161490 263880
rect 154481 263875 154547 263878
rect 147581 263802 147647 263805
rect 135161 263800 135362 263802
rect 135161 263744 135166 263800
rect 135222 263744 135362 263800
rect 135161 263742 135362 263744
rect 144870 263800 147647 263802
rect 144870 263744 147586 263800
rect 147642 263744 147647 263800
rect 144870 263742 147647 263744
rect 161430 263802 161490 263878
rect 171182 263878 180810 263938
rect 161430 263742 171058 263802
rect 96540 263740 96546 263742
rect 135161 263739 135227 263742
rect 86902 263666 86908 263668
rect 82126 263606 86908 263666
rect 86902 263604 86908 263606
rect 86972 263604 86978 263668
rect 111057 263666 111123 263669
rect 115933 263666 115999 263669
rect 111057 263664 115999 263666
rect 111057 263608 111062 263664
rect 111118 263608 115938 263664
rect 115994 263608 115999 263664
rect 111057 263606 115999 263608
rect 111057 263603 111123 263606
rect 115933 263603 115999 263606
rect 140037 263666 140103 263669
rect 144870 263666 144930 263742
rect 147581 263739 147647 263742
rect 140037 263664 144930 263666
rect 140037 263608 140042 263664
rect 140098 263608 144930 263664
rect 140037 263606 144930 263608
rect 170998 263666 171058 263742
rect 171182 263666 171242 263878
rect 180750 263802 180810 263878
rect 190502 263878 200130 263938
rect 180750 263742 190378 263802
rect 170998 263606 171242 263666
rect 190318 263666 190378 263742
rect 190502 263666 190562 263878
rect 200070 263802 200130 263878
rect 209822 263878 219450 263938
rect 200070 263742 209698 263802
rect 190318 263606 190562 263666
rect 209638 263666 209698 263742
rect 209822 263666 209882 263878
rect 219390 263802 219450 263878
rect 229142 263878 238770 263938
rect 219390 263742 229018 263802
rect 209638 263606 209882 263666
rect 228958 263666 229018 263742
rect 229142 263666 229202 263878
rect 238710 263802 238770 263878
rect 248462 263878 258090 263938
rect 238710 263742 248338 263802
rect 228958 263606 229202 263666
rect 248278 263666 248338 263742
rect 248462 263666 248522 263878
rect 258030 263802 258090 263878
rect 267782 263878 277410 263938
rect 258030 263742 267658 263802
rect 248278 263606 248522 263666
rect 267598 263666 267658 263742
rect 267782 263666 267842 263878
rect 277350 263802 277410 263878
rect 287102 263878 296730 263938
rect 277350 263742 286978 263802
rect 267598 263606 267842 263666
rect 286918 263666 286978 263742
rect 287102 263666 287162 263878
rect 296670 263802 296730 263878
rect 306422 263878 316050 263938
rect 296670 263742 306298 263802
rect 286918 263606 287162 263666
rect 306238 263666 306298 263742
rect 306422 263666 306482 263878
rect 315990 263802 316050 263878
rect 325742 263878 335370 263938
rect 315990 263742 325618 263802
rect 306238 263606 306482 263666
rect 325558 263666 325618 263742
rect 325742 263666 325802 263878
rect 335310 263802 335370 263878
rect 345062 263878 354690 263938
rect 335310 263742 344938 263802
rect 325558 263606 325802 263666
rect 344878 263666 344938 263742
rect 345062 263666 345122 263878
rect 354630 263802 354690 263878
rect 364382 263878 374010 263938
rect 354630 263742 364258 263802
rect 344878 263606 345122 263666
rect 364198 263666 364258 263742
rect 364382 263666 364442 263878
rect 373950 263802 374010 263878
rect 383702 263878 393330 263938
rect 373950 263742 383578 263802
rect 364198 263606 364442 263666
rect 383518 263666 383578 263742
rect 383702 263666 383762 263878
rect 393270 263802 393330 263878
rect 403022 263878 412650 263938
rect 393270 263742 402898 263802
rect 383518 263606 383762 263666
rect 402838 263666 402898 263742
rect 403022 263666 403082 263878
rect 412590 263802 412650 263878
rect 422342 263878 431970 263938
rect 412590 263742 422218 263802
rect 402838 263606 403082 263666
rect 422158 263666 422218 263742
rect 422342 263666 422402 263878
rect 431910 263802 431970 263878
rect 441662 263878 451290 263938
rect 431910 263742 441538 263802
rect 422158 263606 422402 263666
rect 441478 263666 441538 263742
rect 441662 263666 441722 263878
rect 451230 263802 451290 263878
rect 460982 263878 470610 263938
rect 451230 263742 460858 263802
rect 441478 263606 441722 263666
rect 460798 263666 460858 263742
rect 460982 263666 461042 263878
rect 470550 263802 470610 263878
rect 480302 263878 489930 263938
rect 470550 263742 480178 263802
rect 460798 263606 461042 263666
rect 480118 263666 480178 263742
rect 480302 263666 480362 263878
rect 489870 263802 489930 263878
rect 499622 263878 509250 263938
rect 489870 263742 499498 263802
rect 480118 263606 480362 263666
rect 499438 263666 499498 263742
rect 499622 263666 499682 263878
rect 509190 263802 509250 263878
rect 518942 263878 528570 263938
rect 509190 263742 518818 263802
rect 499438 263606 499682 263666
rect 518758 263666 518818 263742
rect 518942 263666 519002 263878
rect 528510 263802 528570 263878
rect 538262 263878 547890 263938
rect 528510 263742 538138 263802
rect 518758 263606 519002 263666
rect 538078 263666 538138 263742
rect 538262 263666 538322 263878
rect 547830 263802 547890 263878
rect 557582 263878 567210 263938
rect 547830 263742 557458 263802
rect 538078 263606 538322 263666
rect 557398 263666 557458 263742
rect 557582 263666 557642 263878
rect 567150 263802 567210 263878
rect 583342 263878 584960 263938
rect 583342 263802 583402 263878
rect 567150 263742 576778 263802
rect 557398 263606 557642 263666
rect 576718 263666 576778 263742
rect 576902 263742 583402 263802
rect 583520 263788 584960 263878
rect 576902 263666 576962 263742
rect 576718 263606 576962 263666
rect 140037 263603 140103 263606
rect 74257 259450 74323 259453
rect 74441 259450 74507 259453
rect 74257 259448 74507 259450
rect 74257 259392 74262 259448
rect 74318 259392 74446 259448
rect 74502 259392 74507 259448
rect 74257 259390 74507 259392
rect 74257 259387 74323 259390
rect 74441 259387 74507 259390
rect 579797 252242 579863 252245
rect 583520 252242 584960 252332
rect 579797 252240 584960 252242
rect 579797 252184 579802 252240
rect 579858 252184 584960 252240
rect 579797 252182 584960 252184
rect 579797 252179 579863 252182
rect 583520 252092 584960 252182
rect -960 251290 480 251380
rect 3417 251290 3483 251293
rect -960 251288 3483 251290
rect -960 251232 3422 251288
rect 3478 251232 3483 251288
rect -960 251230 3483 251232
rect -960 251140 480 251230
rect 3417 251227 3483 251230
rect 583520 240396 584960 240636
rect 74257 240138 74323 240141
rect 74441 240138 74507 240141
rect 74257 240136 74507 240138
rect 74257 240080 74262 240136
rect 74318 240080 74446 240136
rect 74502 240080 74507 240136
rect 74257 240078 74507 240080
rect 74257 240075 74323 240078
rect 74441 240075 74507 240078
rect -960 237010 480 237100
rect 3417 237010 3483 237013
rect -960 237008 3483 237010
rect -960 236952 3422 237008
rect 3478 236952 3483 237008
rect -960 236950 3483 236952
rect -960 236860 480 236950
rect 3417 236947 3483 236950
rect 583520 228850 584960 228940
rect 583342 228790 584960 228850
rect 106222 228380 106228 228444
rect 106292 228442 106298 228444
rect 111057 228442 111123 228445
rect 106292 228440 111123 228442
rect 106292 228384 111062 228440
rect 111118 228384 111123 228440
rect 106292 228382 111123 228384
rect 106292 228380 106298 228382
rect 111057 228379 111123 228382
rect 125542 228244 125548 228308
rect 125612 228306 125618 228308
rect 135161 228306 135227 228309
rect 125612 228304 135227 228306
rect 125612 228248 135166 228304
rect 135222 228248 135227 228304
rect 125612 228246 135227 228248
rect 125612 228244 125618 228246
rect 135161 228243 135227 228246
rect 106222 228170 106228 228172
rect 99422 228110 106228 228170
rect 57094 227972 57100 228036
rect 57164 228034 57170 228036
rect 75821 228034 75887 228037
rect 57164 227974 60842 228034
rect 57164 227972 57170 227974
rect 60782 227898 60842 227974
rect 75821 228032 82186 228034
rect 75821 227976 75826 228032
rect 75882 227976 82186 228032
rect 75821 227974 82186 227976
rect 75821 227971 75887 227974
rect 66253 227898 66319 227901
rect 60782 227896 66319 227898
rect 60782 227840 66258 227896
rect 66314 227840 66319 227896
rect 60782 227838 66319 227840
rect 66253 227835 66319 227838
rect 82126 227762 82186 227974
rect 96470 227836 96476 227900
rect 96540 227898 96546 227900
rect 99422 227898 99482 228110
rect 106222 228108 106228 228110
rect 106292 228108 106298 228172
rect 140037 228170 140103 228173
rect 135302 228168 140103 228170
rect 135302 228112 140042 228168
rect 140098 228112 140103 228168
rect 135302 228110 140103 228112
rect 118785 228034 118851 228037
rect 125542 228034 125548 228036
rect 118785 228032 125548 228034
rect 118785 227976 118790 228032
rect 118846 227976 125548 228032
rect 118785 227974 125548 227976
rect 118785 227971 118851 227974
rect 125542 227972 125548 227974
rect 125612 227972 125618 228036
rect 96540 227838 99482 227898
rect 135161 227898 135227 227901
rect 135302 227898 135362 228110
rect 140037 228107 140103 228110
rect 154481 228034 154547 228037
rect 154481 228032 161490 228034
rect 154481 227976 154486 228032
rect 154542 227976 161490 228032
rect 154481 227974 161490 227976
rect 154481 227971 154547 227974
rect 147581 227898 147647 227901
rect 135161 227896 135362 227898
rect 135161 227840 135166 227896
rect 135222 227840 135362 227896
rect 135161 227838 135362 227840
rect 144870 227896 147647 227898
rect 144870 227840 147586 227896
rect 147642 227840 147647 227896
rect 144870 227838 147647 227840
rect 161430 227898 161490 227974
rect 171182 227974 180810 228034
rect 161430 227838 171058 227898
rect 96540 227836 96546 227838
rect 135161 227835 135227 227838
rect 86902 227762 86908 227764
rect 82126 227702 86908 227762
rect 86902 227700 86908 227702
rect 86972 227700 86978 227764
rect 111057 227762 111123 227765
rect 115933 227762 115999 227765
rect 111057 227760 115999 227762
rect 111057 227704 111062 227760
rect 111118 227704 115938 227760
rect 115994 227704 115999 227760
rect 111057 227702 115999 227704
rect 111057 227699 111123 227702
rect 115933 227699 115999 227702
rect 140037 227762 140103 227765
rect 144870 227762 144930 227838
rect 147581 227835 147647 227838
rect 140037 227760 144930 227762
rect 140037 227704 140042 227760
rect 140098 227704 144930 227760
rect 140037 227702 144930 227704
rect 170998 227762 171058 227838
rect 171182 227762 171242 227974
rect 180750 227898 180810 227974
rect 190502 227974 200130 228034
rect 180750 227838 190378 227898
rect 170998 227702 171242 227762
rect 190318 227762 190378 227838
rect 190502 227762 190562 227974
rect 200070 227898 200130 227974
rect 209822 227974 219450 228034
rect 200070 227838 209698 227898
rect 190318 227702 190562 227762
rect 209638 227762 209698 227838
rect 209822 227762 209882 227974
rect 219390 227898 219450 227974
rect 229142 227974 238770 228034
rect 219390 227838 229018 227898
rect 209638 227702 209882 227762
rect 228958 227762 229018 227838
rect 229142 227762 229202 227974
rect 238710 227898 238770 227974
rect 248462 227974 258090 228034
rect 238710 227838 248338 227898
rect 228958 227702 229202 227762
rect 248278 227762 248338 227838
rect 248462 227762 248522 227974
rect 258030 227898 258090 227974
rect 267782 227974 277410 228034
rect 258030 227838 267658 227898
rect 248278 227702 248522 227762
rect 267598 227762 267658 227838
rect 267782 227762 267842 227974
rect 277350 227898 277410 227974
rect 287102 227974 296730 228034
rect 277350 227838 286978 227898
rect 267598 227702 267842 227762
rect 286918 227762 286978 227838
rect 287102 227762 287162 227974
rect 296670 227898 296730 227974
rect 306422 227974 316050 228034
rect 296670 227838 306298 227898
rect 286918 227702 287162 227762
rect 306238 227762 306298 227838
rect 306422 227762 306482 227974
rect 315990 227898 316050 227974
rect 325742 227974 335370 228034
rect 315990 227838 325618 227898
rect 306238 227702 306482 227762
rect 325558 227762 325618 227838
rect 325742 227762 325802 227974
rect 335310 227898 335370 227974
rect 345062 227974 354690 228034
rect 335310 227838 344938 227898
rect 325558 227702 325802 227762
rect 344878 227762 344938 227838
rect 345062 227762 345122 227974
rect 354630 227898 354690 227974
rect 364382 227974 374010 228034
rect 354630 227838 364258 227898
rect 344878 227702 345122 227762
rect 364198 227762 364258 227838
rect 364382 227762 364442 227974
rect 373950 227898 374010 227974
rect 383702 227974 393330 228034
rect 373950 227838 383578 227898
rect 364198 227702 364442 227762
rect 383518 227762 383578 227838
rect 383702 227762 383762 227974
rect 393270 227898 393330 227974
rect 403022 227974 412650 228034
rect 393270 227838 402898 227898
rect 383518 227702 383762 227762
rect 402838 227762 402898 227838
rect 403022 227762 403082 227974
rect 412590 227898 412650 227974
rect 422342 227974 431970 228034
rect 412590 227838 422218 227898
rect 402838 227702 403082 227762
rect 422158 227762 422218 227838
rect 422342 227762 422402 227974
rect 431910 227898 431970 227974
rect 441662 227974 451290 228034
rect 431910 227838 441538 227898
rect 422158 227702 422402 227762
rect 441478 227762 441538 227838
rect 441662 227762 441722 227974
rect 451230 227898 451290 227974
rect 460982 227974 470610 228034
rect 451230 227838 460858 227898
rect 441478 227702 441722 227762
rect 460798 227762 460858 227838
rect 460982 227762 461042 227974
rect 470550 227898 470610 227974
rect 480302 227974 489930 228034
rect 470550 227838 480178 227898
rect 460798 227702 461042 227762
rect 480118 227762 480178 227838
rect 480302 227762 480362 227974
rect 489870 227898 489930 227974
rect 499622 227974 509250 228034
rect 489870 227838 499498 227898
rect 480118 227702 480362 227762
rect 499438 227762 499498 227838
rect 499622 227762 499682 227974
rect 509190 227898 509250 227974
rect 518942 227974 528570 228034
rect 509190 227838 518818 227898
rect 499438 227702 499682 227762
rect 518758 227762 518818 227838
rect 518942 227762 519002 227974
rect 528510 227898 528570 227974
rect 538262 227974 547890 228034
rect 528510 227838 538138 227898
rect 518758 227702 519002 227762
rect 538078 227762 538138 227838
rect 538262 227762 538322 227974
rect 547830 227898 547890 227974
rect 557582 227974 567210 228034
rect 547830 227838 557458 227898
rect 538078 227702 538322 227762
rect 557398 227762 557458 227838
rect 557582 227762 557642 227974
rect 567150 227898 567210 227974
rect 583342 227898 583402 228790
rect 583520 228700 584960 228790
rect 567150 227838 576778 227898
rect 557398 227702 557642 227762
rect 576718 227762 576778 227838
rect 576902 227838 583402 227898
rect 576902 227762 576962 227838
rect 576718 227702 576962 227762
rect 140037 227699 140103 227702
rect 86902 227428 86908 227492
rect 86972 227490 86978 227492
rect 96470 227490 96476 227492
rect 86972 227430 96476 227490
rect 86972 227428 86978 227430
rect 96470 227428 96476 227430
rect 96540 227428 96546 227492
rect -960 222594 480 222684
rect 3141 222594 3207 222597
rect -960 222592 3207 222594
rect -960 222536 3146 222592
rect 3202 222536 3207 222592
rect -960 222534 3207 222536
rect -960 222444 480 222534
rect 3141 222531 3207 222534
rect 74257 220826 74323 220829
rect 74441 220826 74507 220829
rect 74257 220824 74507 220826
rect 74257 220768 74262 220824
rect 74318 220768 74446 220824
rect 74502 220768 74507 220824
rect 74257 220766 74507 220768
rect 74257 220763 74323 220766
rect 74441 220763 74507 220766
rect 125542 217228 125548 217292
rect 125612 217290 125618 217292
rect 135161 217290 135227 217293
rect 125612 217288 135227 217290
rect 125612 217232 135166 217288
rect 135222 217232 135227 217288
rect 125612 217230 135227 217232
rect 125612 217228 125618 217230
rect 135161 217227 135227 217230
rect 140037 217154 140103 217157
rect 135302 217152 140103 217154
rect 135302 217096 140042 217152
rect 140098 217096 140103 217152
rect 135302 217094 140103 217096
rect 57278 216956 57284 217020
rect 57348 217018 57354 217020
rect 77201 217018 77267 217021
rect 118785 217018 118851 217021
rect 125542 217018 125548 217020
rect 57348 216958 60842 217018
rect 57348 216956 57354 216958
rect 60782 216882 60842 216958
rect 77201 217016 80162 217018
rect 77201 216960 77206 217016
rect 77262 216960 80162 217016
rect 77201 216958 80162 216960
rect 77201 216955 77267 216958
rect 69381 216882 69447 216885
rect 60782 216880 69447 216882
rect 60782 216824 69386 216880
rect 69442 216824 69447 216880
rect 60782 216822 69447 216824
rect 80102 216882 80162 216958
rect 96478 216958 109050 217018
rect 89529 216882 89595 216885
rect 80102 216880 89595 216882
rect 80102 216824 89534 216880
rect 89590 216824 89595 216880
rect 80102 216822 89595 216824
rect 69381 216819 69447 216822
rect 89529 216819 89595 216822
rect 91737 216882 91803 216885
rect 96478 216882 96538 216958
rect 91737 216880 96538 216882
rect 91737 216824 91742 216880
rect 91798 216824 96538 216880
rect 91737 216822 96538 216824
rect 91737 216819 91803 216822
rect 108990 216746 109050 216958
rect 118785 217016 125548 217018
rect 118785 216960 118790 217016
rect 118846 216960 125548 217016
rect 118785 216958 125548 216960
rect 118785 216955 118851 216958
rect 125542 216956 125548 216958
rect 125612 216956 125618 217020
rect 135161 216882 135227 216885
rect 135302 216882 135362 217094
rect 140037 217091 140103 217094
rect 154481 217018 154547 217021
rect 583520 217018 584960 217108
rect 154481 217016 161490 217018
rect 154481 216960 154486 217016
rect 154542 216960 161490 217016
rect 154481 216958 161490 216960
rect 154481 216955 154547 216958
rect 147581 216882 147647 216885
rect 135161 216880 135362 216882
rect 135161 216824 135166 216880
rect 135222 216824 135362 216880
rect 135161 216822 135362 216824
rect 144870 216880 147647 216882
rect 144870 216824 147586 216880
rect 147642 216824 147647 216880
rect 144870 216822 147647 216824
rect 161430 216882 161490 216958
rect 171182 216958 180810 217018
rect 161430 216822 171058 216882
rect 135161 216819 135227 216822
rect 115933 216746 115999 216749
rect 108990 216744 115999 216746
rect 108990 216688 115938 216744
rect 115994 216688 115999 216744
rect 108990 216686 115999 216688
rect 115933 216683 115999 216686
rect 140037 216746 140103 216749
rect 144870 216746 144930 216822
rect 147581 216819 147647 216822
rect 140037 216744 144930 216746
rect 140037 216688 140042 216744
rect 140098 216688 144930 216744
rect 140037 216686 144930 216688
rect 170998 216746 171058 216822
rect 171182 216746 171242 216958
rect 180750 216882 180810 216958
rect 190502 216958 200130 217018
rect 180750 216822 190378 216882
rect 170998 216686 171242 216746
rect 190318 216746 190378 216822
rect 190502 216746 190562 216958
rect 200070 216882 200130 216958
rect 209822 216958 219450 217018
rect 200070 216822 209698 216882
rect 190318 216686 190562 216746
rect 209638 216746 209698 216822
rect 209822 216746 209882 216958
rect 219390 216882 219450 216958
rect 229142 216958 238770 217018
rect 219390 216822 229018 216882
rect 209638 216686 209882 216746
rect 228958 216746 229018 216822
rect 229142 216746 229202 216958
rect 238710 216882 238770 216958
rect 248462 216958 258090 217018
rect 238710 216822 248338 216882
rect 228958 216686 229202 216746
rect 248278 216746 248338 216822
rect 248462 216746 248522 216958
rect 258030 216882 258090 216958
rect 267782 216958 277410 217018
rect 258030 216822 267658 216882
rect 248278 216686 248522 216746
rect 267598 216746 267658 216822
rect 267782 216746 267842 216958
rect 277350 216882 277410 216958
rect 287102 216958 296730 217018
rect 277350 216822 286978 216882
rect 267598 216686 267842 216746
rect 286918 216746 286978 216822
rect 287102 216746 287162 216958
rect 296670 216882 296730 216958
rect 306422 216958 316050 217018
rect 296670 216822 306298 216882
rect 286918 216686 287162 216746
rect 306238 216746 306298 216822
rect 306422 216746 306482 216958
rect 315990 216882 316050 216958
rect 325742 216958 335370 217018
rect 315990 216822 325618 216882
rect 306238 216686 306482 216746
rect 325558 216746 325618 216822
rect 325742 216746 325802 216958
rect 335310 216882 335370 216958
rect 345062 216958 354690 217018
rect 335310 216822 344938 216882
rect 325558 216686 325802 216746
rect 344878 216746 344938 216822
rect 345062 216746 345122 216958
rect 354630 216882 354690 216958
rect 364382 216958 374010 217018
rect 354630 216822 364258 216882
rect 344878 216686 345122 216746
rect 364198 216746 364258 216822
rect 364382 216746 364442 216958
rect 373950 216882 374010 216958
rect 383702 216958 393330 217018
rect 373950 216822 383578 216882
rect 364198 216686 364442 216746
rect 383518 216746 383578 216822
rect 383702 216746 383762 216958
rect 393270 216882 393330 216958
rect 403022 216958 412650 217018
rect 393270 216822 402898 216882
rect 383518 216686 383762 216746
rect 402838 216746 402898 216822
rect 403022 216746 403082 216958
rect 412590 216882 412650 216958
rect 422342 216958 431970 217018
rect 412590 216822 422218 216882
rect 402838 216686 403082 216746
rect 422158 216746 422218 216822
rect 422342 216746 422402 216958
rect 431910 216882 431970 216958
rect 441662 216958 451290 217018
rect 431910 216822 441538 216882
rect 422158 216686 422402 216746
rect 441478 216746 441538 216822
rect 441662 216746 441722 216958
rect 451230 216882 451290 216958
rect 460982 216958 470610 217018
rect 451230 216822 460858 216882
rect 441478 216686 441722 216746
rect 460798 216746 460858 216822
rect 460982 216746 461042 216958
rect 470550 216882 470610 216958
rect 480302 216958 489930 217018
rect 470550 216822 480178 216882
rect 460798 216686 461042 216746
rect 480118 216746 480178 216822
rect 480302 216746 480362 216958
rect 489870 216882 489930 216958
rect 499622 216958 509250 217018
rect 489870 216822 499498 216882
rect 480118 216686 480362 216746
rect 499438 216746 499498 216822
rect 499622 216746 499682 216958
rect 509190 216882 509250 216958
rect 518942 216958 528570 217018
rect 509190 216822 518818 216882
rect 499438 216686 499682 216746
rect 518758 216746 518818 216822
rect 518942 216746 519002 216958
rect 528510 216882 528570 216958
rect 538262 216958 547890 217018
rect 528510 216822 538138 216882
rect 518758 216686 519002 216746
rect 538078 216746 538138 216822
rect 538262 216746 538322 216958
rect 547830 216882 547890 216958
rect 557582 216958 567210 217018
rect 547830 216822 557458 216882
rect 538078 216686 538322 216746
rect 557398 216746 557458 216822
rect 557582 216746 557642 216958
rect 567150 216882 567210 216958
rect 583342 216958 584960 217018
rect 583342 216882 583402 216958
rect 567150 216822 576778 216882
rect 557398 216686 557642 216746
rect 576718 216746 576778 216822
rect 576902 216822 583402 216882
rect 583520 216868 584960 216958
rect 576902 216746 576962 216822
rect 576718 216686 576962 216746
rect 140037 216683 140103 216686
rect 74257 211170 74323 211173
rect 74441 211170 74507 211173
rect 74257 211168 74507 211170
rect 74257 211112 74262 211168
rect 74318 211112 74446 211168
rect 74502 211112 74507 211168
rect 74257 211110 74507 211112
rect 74257 211107 74323 211110
rect 74441 211107 74507 211110
rect -960 208178 480 208268
rect 2773 208178 2839 208181
rect -960 208176 2839 208178
rect -960 208120 2778 208176
rect 2834 208120 2839 208176
rect -960 208118 2839 208120
rect -960 208028 480 208118
rect 2773 208115 2839 208118
rect 579797 205322 579863 205325
rect 583520 205322 584960 205412
rect 579797 205320 584960 205322
rect 579797 205264 579802 205320
rect 579858 205264 584960 205320
rect 579797 205262 584960 205264
rect 579797 205259 579863 205262
rect 583520 205172 584960 205262
rect -960 193898 480 193988
rect 2865 193898 2931 193901
rect -960 193896 2931 193898
rect -960 193840 2870 193896
rect 2926 193840 2931 193896
rect -960 193838 2931 193840
rect -960 193748 480 193838
rect 2865 193835 2931 193838
rect 583520 193476 584960 193716
rect 583520 181930 584960 182020
rect 583342 181870 584960 181930
rect 106222 181460 106228 181524
rect 106292 181522 106298 181524
rect 111057 181522 111123 181525
rect 106292 181520 111123 181522
rect 106292 181464 111062 181520
rect 111118 181464 111123 181520
rect 106292 181462 111123 181464
rect 106292 181460 106298 181462
rect 111057 181459 111123 181462
rect 106222 181250 106228 181252
rect 99422 181190 106228 181250
rect 57462 181052 57468 181116
rect 57532 181114 57538 181116
rect 77201 181114 77267 181117
rect 57532 181054 60842 181114
rect 57532 181052 57538 181054
rect 60782 180978 60842 181054
rect 77201 181112 82186 181114
rect 77201 181056 77206 181112
rect 77262 181056 82186 181112
rect 77201 181054 82186 181056
rect 77201 181051 77267 181054
rect 69381 180978 69447 180981
rect 60782 180976 69447 180978
rect 60782 180920 69386 180976
rect 69442 180920 69447 180976
rect 60782 180918 69447 180920
rect 69381 180915 69447 180918
rect 82126 180842 82186 181054
rect 96470 180916 96476 180980
rect 96540 180978 96546 180980
rect 99422 180978 99482 181190
rect 106222 181188 106228 181190
rect 106292 181188 106298 181252
rect 166950 181054 176578 181114
rect 128261 180978 128327 180981
rect 96540 180918 99482 180978
rect 118742 180976 128327 180978
rect 118742 180920 128266 180976
rect 128322 180920 128327 180976
rect 118742 180918 128327 180920
rect 96540 180916 96546 180918
rect 96470 180842 96476 180844
rect 82126 180782 96476 180842
rect 96470 180780 96476 180782
rect 96540 180780 96546 180844
rect 111057 180842 111123 180845
rect 118742 180842 118802 180918
rect 128261 180915 128327 180918
rect 128445 180978 128511 180981
rect 128445 180976 137938 180978
rect 128445 180920 128450 180976
rect 128506 180920 137938 180976
rect 128445 180918 137938 180920
rect 128445 180915 128511 180918
rect 111057 180840 118802 180842
rect 111057 180784 111062 180840
rect 111118 180784 118802 180840
rect 111057 180782 118802 180784
rect 137878 180842 137938 180918
rect 166950 180842 167010 181054
rect 137878 180782 167010 180842
rect 176518 180842 176578 181054
rect 186270 181054 195898 181114
rect 186270 180842 186330 181054
rect 176518 180782 186330 180842
rect 195838 180842 195898 181054
rect 205590 181054 215218 181114
rect 205590 180842 205650 181054
rect 195838 180782 205650 180842
rect 215158 180842 215218 181054
rect 224910 181054 234538 181114
rect 224910 180842 224970 181054
rect 215158 180782 224970 180842
rect 234478 180842 234538 181054
rect 244230 181054 253858 181114
rect 244230 180842 244290 181054
rect 234478 180782 244290 180842
rect 253798 180842 253858 181054
rect 263550 181054 273178 181114
rect 263550 180842 263610 181054
rect 253798 180782 263610 180842
rect 273118 180842 273178 181054
rect 277350 181054 296730 181114
rect 277350 180842 277410 181054
rect 296670 180978 296730 181054
rect 306422 181054 316050 181114
rect 296670 180918 306298 180978
rect 273118 180782 277410 180842
rect 306238 180842 306298 180918
rect 306422 180842 306482 181054
rect 315990 180978 316050 181054
rect 325742 181054 335370 181114
rect 315990 180918 325618 180978
rect 306238 180782 306482 180842
rect 325558 180842 325618 180918
rect 325742 180842 325802 181054
rect 335310 180978 335370 181054
rect 345062 181054 354690 181114
rect 335310 180918 344938 180978
rect 325558 180782 325802 180842
rect 344878 180842 344938 180918
rect 345062 180842 345122 181054
rect 354630 180978 354690 181054
rect 364382 181054 374010 181114
rect 354630 180918 364258 180978
rect 344878 180782 345122 180842
rect 364198 180842 364258 180918
rect 364382 180842 364442 181054
rect 373950 180978 374010 181054
rect 383702 181054 393330 181114
rect 373950 180918 383578 180978
rect 364198 180782 364442 180842
rect 383518 180842 383578 180918
rect 383702 180842 383762 181054
rect 393270 180978 393330 181054
rect 403022 181054 412650 181114
rect 393270 180918 402898 180978
rect 383518 180782 383762 180842
rect 402838 180842 402898 180918
rect 403022 180842 403082 181054
rect 412590 180978 412650 181054
rect 422342 181054 431970 181114
rect 412590 180918 422218 180978
rect 402838 180782 403082 180842
rect 422158 180842 422218 180918
rect 422342 180842 422402 181054
rect 431910 180978 431970 181054
rect 441662 181054 451290 181114
rect 431910 180918 441538 180978
rect 422158 180782 422402 180842
rect 441478 180842 441538 180918
rect 441662 180842 441722 181054
rect 451230 180978 451290 181054
rect 460982 181054 470610 181114
rect 451230 180918 460858 180978
rect 441478 180782 441722 180842
rect 460798 180842 460858 180918
rect 460982 180842 461042 181054
rect 470550 180978 470610 181054
rect 480302 181054 489930 181114
rect 470550 180918 480178 180978
rect 460798 180782 461042 180842
rect 480118 180842 480178 180918
rect 480302 180842 480362 181054
rect 489870 180978 489930 181054
rect 499622 181054 509250 181114
rect 489870 180918 499498 180978
rect 480118 180782 480362 180842
rect 499438 180842 499498 180918
rect 499622 180842 499682 181054
rect 509190 180978 509250 181054
rect 518942 181054 528570 181114
rect 509190 180918 518818 180978
rect 499438 180782 499682 180842
rect 518758 180842 518818 180918
rect 518942 180842 519002 181054
rect 528510 180978 528570 181054
rect 538262 181054 547890 181114
rect 528510 180918 538138 180978
rect 518758 180782 519002 180842
rect 538078 180842 538138 180918
rect 538262 180842 538322 181054
rect 547830 180978 547890 181054
rect 557582 181054 567210 181114
rect 547830 180918 557458 180978
rect 538078 180782 538322 180842
rect 557398 180842 557458 180918
rect 557582 180842 557642 181054
rect 567150 180978 567210 181054
rect 583342 180978 583402 181870
rect 583520 181780 584960 181870
rect 567150 180918 576778 180978
rect 557398 180782 557642 180842
rect 576718 180842 576778 180918
rect 576902 180918 583402 180978
rect 576902 180842 576962 180918
rect 576718 180782 576962 180842
rect 111057 180779 111123 180782
rect -960 179482 480 179572
rect 3233 179482 3299 179485
rect -960 179480 3299 179482
rect -960 179424 3238 179480
rect 3294 179424 3299 179480
rect -960 179422 3299 179424
rect -960 179332 480 179422
rect 3233 179419 3299 179422
rect 74257 172546 74323 172549
rect 74441 172546 74507 172549
rect 74257 172544 74507 172546
rect 74257 172488 74262 172544
rect 74318 172488 74446 172544
rect 74502 172488 74507 172544
rect 74257 172486 74507 172488
rect 74257 172483 74323 172486
rect 74441 172483 74507 172486
rect 106222 170444 106228 170508
rect 106292 170506 106298 170508
rect 111057 170506 111123 170509
rect 106292 170504 111123 170506
rect 106292 170448 111062 170504
rect 111118 170448 111123 170504
rect 106292 170446 111123 170448
rect 106292 170444 106298 170446
rect 111057 170443 111123 170446
rect 125542 170308 125548 170372
rect 125612 170370 125618 170372
rect 135161 170370 135227 170373
rect 125612 170368 135227 170370
rect 125612 170312 135166 170368
rect 135222 170312 135227 170368
rect 125612 170310 135227 170312
rect 125612 170308 125618 170310
rect 135161 170307 135227 170310
rect 106222 170234 106228 170236
rect 99422 170174 106228 170234
rect 57646 170036 57652 170100
rect 57716 170098 57722 170100
rect 75821 170098 75887 170101
rect 89529 170098 89595 170101
rect 57716 170038 60842 170098
rect 57716 170036 57722 170038
rect 60782 169962 60842 170038
rect 75821 170096 82186 170098
rect 75821 170040 75826 170096
rect 75882 170040 82186 170096
rect 75821 170038 82186 170040
rect 75821 170035 75887 170038
rect 66253 169962 66319 169965
rect 60782 169960 66319 169962
rect 60782 169904 66258 169960
rect 66314 169904 66319 169960
rect 60782 169902 66319 169904
rect 66253 169899 66319 169902
rect 82126 169826 82186 170038
rect 89529 170096 96538 170098
rect 89529 170040 89534 170096
rect 89590 170040 96538 170096
rect 89529 170038 96538 170040
rect 89529 170035 89595 170038
rect 96478 169962 96538 170038
rect 99422 169962 99482 170174
rect 106222 170172 106228 170174
rect 106292 170172 106298 170236
rect 140037 170234 140103 170237
rect 135302 170232 140103 170234
rect 135302 170176 140042 170232
rect 140098 170176 140103 170232
rect 135302 170174 140103 170176
rect 118785 170098 118851 170101
rect 125542 170098 125548 170100
rect 118785 170096 125548 170098
rect 118785 170040 118790 170096
rect 118846 170040 125548 170096
rect 118785 170038 125548 170040
rect 118785 170035 118851 170038
rect 125542 170036 125548 170038
rect 125612 170036 125618 170100
rect 96478 169902 99482 169962
rect 135161 169962 135227 169965
rect 135302 169962 135362 170174
rect 140037 170171 140103 170174
rect 154481 170098 154547 170101
rect 583520 170098 584960 170188
rect 154481 170096 161490 170098
rect 154481 170040 154486 170096
rect 154542 170040 161490 170096
rect 154481 170038 161490 170040
rect 154481 170035 154547 170038
rect 147581 169962 147647 169965
rect 135161 169960 135362 169962
rect 135161 169904 135166 169960
rect 135222 169904 135362 169960
rect 135161 169902 135362 169904
rect 144870 169960 147647 169962
rect 144870 169904 147586 169960
rect 147642 169904 147647 169960
rect 144870 169902 147647 169904
rect 161430 169962 161490 170038
rect 171182 170038 180810 170098
rect 161430 169902 171058 169962
rect 135161 169899 135227 169902
rect 89529 169826 89595 169829
rect 82126 169824 89595 169826
rect 82126 169768 89534 169824
rect 89590 169768 89595 169824
rect 82126 169766 89595 169768
rect 89529 169763 89595 169766
rect 111057 169826 111123 169829
rect 115933 169826 115999 169829
rect 111057 169824 115999 169826
rect 111057 169768 111062 169824
rect 111118 169768 115938 169824
rect 115994 169768 115999 169824
rect 111057 169766 115999 169768
rect 111057 169763 111123 169766
rect 115933 169763 115999 169766
rect 140037 169826 140103 169829
rect 144870 169826 144930 169902
rect 147581 169899 147647 169902
rect 140037 169824 144930 169826
rect 140037 169768 140042 169824
rect 140098 169768 144930 169824
rect 140037 169766 144930 169768
rect 170998 169826 171058 169902
rect 171182 169826 171242 170038
rect 180750 169962 180810 170038
rect 190502 170038 200130 170098
rect 180750 169902 190378 169962
rect 170998 169766 171242 169826
rect 190318 169826 190378 169902
rect 190502 169826 190562 170038
rect 200070 169962 200130 170038
rect 209822 170038 219450 170098
rect 200070 169902 209698 169962
rect 190318 169766 190562 169826
rect 209638 169826 209698 169902
rect 209822 169826 209882 170038
rect 219390 169962 219450 170038
rect 229142 170038 238770 170098
rect 219390 169902 229018 169962
rect 209638 169766 209882 169826
rect 228958 169826 229018 169902
rect 229142 169826 229202 170038
rect 238710 169962 238770 170038
rect 248462 170038 258090 170098
rect 238710 169902 248338 169962
rect 228958 169766 229202 169826
rect 248278 169826 248338 169902
rect 248462 169826 248522 170038
rect 258030 169962 258090 170038
rect 267782 170038 277410 170098
rect 258030 169902 267658 169962
rect 248278 169766 248522 169826
rect 267598 169826 267658 169902
rect 267782 169826 267842 170038
rect 277350 169962 277410 170038
rect 287102 170038 296730 170098
rect 277350 169902 286978 169962
rect 267598 169766 267842 169826
rect 286918 169826 286978 169902
rect 287102 169826 287162 170038
rect 296670 169962 296730 170038
rect 306422 170038 316050 170098
rect 296670 169902 306298 169962
rect 286918 169766 287162 169826
rect 306238 169826 306298 169902
rect 306422 169826 306482 170038
rect 315990 169962 316050 170038
rect 325742 170038 335370 170098
rect 315990 169902 325618 169962
rect 306238 169766 306482 169826
rect 325558 169826 325618 169902
rect 325742 169826 325802 170038
rect 335310 169962 335370 170038
rect 345062 170038 354690 170098
rect 335310 169902 344938 169962
rect 325558 169766 325802 169826
rect 344878 169826 344938 169902
rect 345062 169826 345122 170038
rect 354630 169962 354690 170038
rect 364382 170038 374010 170098
rect 354630 169902 364258 169962
rect 344878 169766 345122 169826
rect 364198 169826 364258 169902
rect 364382 169826 364442 170038
rect 373950 169962 374010 170038
rect 383702 170038 393330 170098
rect 373950 169902 383578 169962
rect 364198 169766 364442 169826
rect 383518 169826 383578 169902
rect 383702 169826 383762 170038
rect 393270 169962 393330 170038
rect 403022 170038 412650 170098
rect 393270 169902 402898 169962
rect 383518 169766 383762 169826
rect 402838 169826 402898 169902
rect 403022 169826 403082 170038
rect 412590 169962 412650 170038
rect 422342 170038 431970 170098
rect 412590 169902 422218 169962
rect 402838 169766 403082 169826
rect 422158 169826 422218 169902
rect 422342 169826 422402 170038
rect 431910 169962 431970 170038
rect 441662 170038 451290 170098
rect 431910 169902 441538 169962
rect 422158 169766 422402 169826
rect 441478 169826 441538 169902
rect 441662 169826 441722 170038
rect 451230 169962 451290 170038
rect 460982 170038 470610 170098
rect 451230 169902 460858 169962
rect 441478 169766 441722 169826
rect 460798 169826 460858 169902
rect 460982 169826 461042 170038
rect 470550 169962 470610 170038
rect 480302 170038 489930 170098
rect 470550 169902 480178 169962
rect 460798 169766 461042 169826
rect 480118 169826 480178 169902
rect 480302 169826 480362 170038
rect 489870 169962 489930 170038
rect 499622 170038 509250 170098
rect 489870 169902 499498 169962
rect 480118 169766 480362 169826
rect 499438 169826 499498 169902
rect 499622 169826 499682 170038
rect 509190 169962 509250 170038
rect 518942 170038 528570 170098
rect 509190 169902 518818 169962
rect 499438 169766 499682 169826
rect 518758 169826 518818 169902
rect 518942 169826 519002 170038
rect 528510 169962 528570 170038
rect 538262 170038 547890 170098
rect 528510 169902 538138 169962
rect 518758 169766 519002 169826
rect 538078 169826 538138 169902
rect 538262 169826 538322 170038
rect 547830 169962 547890 170038
rect 557582 170038 567210 170098
rect 547830 169902 557458 169962
rect 538078 169766 538322 169826
rect 557398 169826 557458 169902
rect 557582 169826 557642 170038
rect 567150 169962 567210 170038
rect 583342 170038 584960 170098
rect 583342 169962 583402 170038
rect 567150 169902 576778 169962
rect 557398 169766 557642 169826
rect 576718 169826 576778 169902
rect 576902 169902 583402 169962
rect 583520 169948 584960 170038
rect 576902 169826 576962 169902
rect 576718 169766 576962 169826
rect 140037 169763 140103 169766
rect -960 165066 480 165156
rect 2773 165066 2839 165069
rect -960 165064 2839 165066
rect -960 165008 2778 165064
rect 2834 165008 2839 165064
rect -960 165006 2839 165008
rect -960 164916 480 165006
rect 2773 165003 2839 165006
rect 579797 158402 579863 158405
rect 583520 158402 584960 158492
rect 579797 158400 584960 158402
rect 579797 158344 579802 158400
rect 579858 158344 584960 158400
rect 579797 158342 584960 158344
rect 579797 158339 579863 158342
rect 583520 158252 584960 158342
rect 74257 153234 74323 153237
rect 74441 153234 74507 153237
rect 74257 153232 74507 153234
rect 74257 153176 74262 153232
rect 74318 153176 74446 153232
rect 74502 153176 74507 153232
rect 74257 153174 74507 153176
rect 74257 153171 74323 153174
rect 74441 153171 74507 153174
rect -960 150786 480 150876
rect 3141 150786 3207 150789
rect -960 150784 3207 150786
rect -960 150728 3146 150784
rect 3202 150728 3207 150784
rect -960 150726 3207 150728
rect -960 150636 480 150726
rect 3141 150723 3207 150726
rect 583520 146556 584960 146796
rect 89253 144938 89319 144941
rect 89437 144938 89503 144941
rect 89253 144936 89503 144938
rect 89253 144880 89258 144936
rect 89314 144880 89442 144936
rect 89498 144880 89503 144936
rect 89253 144878 89503 144880
rect 89253 144875 89319 144878
rect 89437 144875 89503 144878
rect -960 136370 480 136460
rect 3233 136370 3299 136373
rect -960 136368 3299 136370
rect -960 136312 3238 136368
rect 3294 136312 3299 136368
rect -960 136310 3299 136312
rect -960 136220 480 136310
rect 3233 136307 3299 136310
rect 580165 134874 580231 134877
rect 583520 134874 584960 134964
rect 580165 134872 584960 134874
rect 580165 134816 580170 134872
rect 580226 134816 584960 134872
rect 580165 134814 584960 134816
rect 580165 134811 580231 134814
rect 583520 134724 584960 134814
rect 74441 125626 74507 125629
rect 74625 125626 74691 125629
rect 74441 125624 74691 125626
rect 74441 125568 74446 125624
rect 74502 125568 74630 125624
rect 74686 125568 74691 125624
rect 74441 125566 74691 125568
rect 74441 125563 74507 125566
rect 74625 125563 74691 125566
rect 74441 124130 74507 124133
rect 74717 124130 74783 124133
rect 74441 124128 74783 124130
rect 74441 124072 74446 124128
rect 74502 124072 74722 124128
rect 74778 124072 74783 124128
rect 74441 124070 74783 124072
rect 74441 124067 74507 124070
rect 74717 124067 74783 124070
rect 580165 123178 580231 123181
rect 583520 123178 584960 123268
rect 580165 123176 584960 123178
rect 580165 123120 580170 123176
rect 580226 123120 584960 123176
rect 580165 123118 584960 123120
rect 580165 123115 580231 123118
rect 583520 123028 584960 123118
rect -960 122090 480 122180
rect 2773 122090 2839 122093
rect -960 122088 2839 122090
rect -960 122032 2778 122088
rect 2834 122032 2839 122088
rect -960 122030 2839 122032
rect -960 121940 480 122030
rect 2773 122027 2839 122030
rect 579797 111482 579863 111485
rect 583520 111482 584960 111572
rect 579797 111480 584960 111482
rect 579797 111424 579802 111480
rect 579858 111424 584960 111480
rect 579797 111422 584960 111424
rect 579797 111419 579863 111422
rect 583520 111332 584960 111422
rect -960 107674 480 107764
rect 3233 107674 3299 107677
rect -960 107672 3299 107674
rect -960 107616 3238 107672
rect 3294 107616 3299 107672
rect -960 107614 3299 107616
rect -960 107524 480 107614
rect 3233 107611 3299 107614
rect 583520 99636 584960 99876
rect -960 93258 480 93348
rect 3417 93258 3483 93261
rect -960 93256 3483 93258
rect -960 93200 3422 93256
rect 3478 93200 3483 93256
rect -960 93198 3483 93200
rect -960 93108 480 93198
rect 3417 93195 3483 93198
rect 580165 87954 580231 87957
rect 583520 87954 584960 88044
rect 580165 87952 584960 87954
rect 580165 87896 580170 87952
rect 580226 87896 584960 87952
rect 580165 87894 584960 87896
rect 580165 87891 580231 87894
rect 583520 87804 584960 87894
rect -960 78978 480 79068
rect 2773 78978 2839 78981
rect -960 78976 2839 78978
rect -960 78920 2778 78976
rect 2834 78920 2839 78976
rect -960 78918 2839 78920
rect -960 78828 480 78918
rect 2773 78915 2839 78918
rect 125542 76468 125548 76532
rect 125612 76530 125618 76532
rect 135161 76530 135227 76533
rect 125612 76528 135227 76530
rect 125612 76472 135166 76528
rect 135222 76472 135227 76528
rect 125612 76470 135227 76472
rect 125612 76468 125618 76470
rect 135161 76467 135227 76470
rect 140037 76394 140103 76397
rect 135302 76392 140103 76394
rect 135302 76336 140042 76392
rect 140098 76336 140103 76392
rect 135302 76334 140103 76336
rect 57830 76196 57836 76260
rect 57900 76258 57906 76260
rect 77201 76258 77267 76261
rect 118785 76258 118851 76261
rect 125542 76258 125548 76260
rect 57900 76198 60842 76258
rect 57900 76196 57906 76198
rect 60782 76122 60842 76198
rect 77201 76256 80162 76258
rect 77201 76200 77206 76256
rect 77262 76200 80162 76256
rect 77201 76198 80162 76200
rect 77201 76195 77267 76198
rect 77201 76122 77267 76125
rect 60782 76120 77267 76122
rect 60782 76064 77206 76120
rect 77262 76064 77267 76120
rect 60782 76062 77267 76064
rect 80102 76122 80162 76198
rect 96478 76198 109050 76258
rect 89621 76122 89687 76125
rect 80102 76120 89687 76122
rect 80102 76064 89626 76120
rect 89682 76064 89687 76120
rect 80102 76062 89687 76064
rect 77201 76059 77267 76062
rect 89621 76059 89687 76062
rect 91737 76122 91803 76125
rect 96478 76122 96538 76198
rect 91737 76120 96538 76122
rect 91737 76064 91742 76120
rect 91798 76064 96538 76120
rect 91737 76062 96538 76064
rect 91737 76059 91803 76062
rect 108990 75986 109050 76198
rect 118785 76256 125548 76258
rect 118785 76200 118790 76256
rect 118846 76200 125548 76256
rect 118785 76198 125548 76200
rect 118785 76195 118851 76198
rect 125542 76196 125548 76198
rect 125612 76196 125618 76260
rect 135161 76122 135227 76125
rect 135302 76122 135362 76334
rect 140037 76331 140103 76334
rect 154481 76258 154547 76261
rect 583520 76258 584960 76348
rect 154481 76256 161490 76258
rect 154481 76200 154486 76256
rect 154542 76200 161490 76256
rect 154481 76198 161490 76200
rect 154481 76195 154547 76198
rect 147581 76122 147647 76125
rect 135161 76120 135362 76122
rect 135161 76064 135166 76120
rect 135222 76064 135362 76120
rect 135161 76062 135362 76064
rect 144870 76120 147647 76122
rect 144870 76064 147586 76120
rect 147642 76064 147647 76120
rect 144870 76062 147647 76064
rect 161430 76122 161490 76198
rect 171182 76198 180810 76258
rect 161430 76062 171058 76122
rect 135161 76059 135227 76062
rect 115933 75986 115999 75989
rect 108990 75984 115999 75986
rect 108990 75928 115938 75984
rect 115994 75928 115999 75984
rect 108990 75926 115999 75928
rect 115933 75923 115999 75926
rect 140037 75986 140103 75989
rect 144870 75986 144930 76062
rect 147581 76059 147647 76062
rect 140037 75984 144930 75986
rect 140037 75928 140042 75984
rect 140098 75928 144930 75984
rect 140037 75926 144930 75928
rect 170998 75986 171058 76062
rect 171182 75986 171242 76198
rect 180750 76122 180810 76198
rect 190502 76198 200130 76258
rect 180750 76062 190378 76122
rect 170998 75926 171242 75986
rect 190318 75986 190378 76062
rect 190502 75986 190562 76198
rect 200070 76122 200130 76198
rect 209822 76198 219450 76258
rect 200070 76062 209698 76122
rect 190318 75926 190562 75986
rect 209638 75986 209698 76062
rect 209822 75986 209882 76198
rect 219390 76122 219450 76198
rect 229142 76198 238770 76258
rect 219390 76062 229018 76122
rect 209638 75926 209882 75986
rect 228958 75986 229018 76062
rect 229142 75986 229202 76198
rect 238710 76122 238770 76198
rect 248462 76198 258090 76258
rect 238710 76062 248338 76122
rect 228958 75926 229202 75986
rect 248278 75986 248338 76062
rect 248462 75986 248522 76198
rect 258030 76122 258090 76198
rect 267782 76198 277410 76258
rect 258030 76062 267658 76122
rect 248278 75926 248522 75986
rect 267598 75986 267658 76062
rect 267782 75986 267842 76198
rect 277350 76122 277410 76198
rect 287102 76198 296730 76258
rect 277350 76062 286978 76122
rect 267598 75926 267842 75986
rect 286918 75986 286978 76062
rect 287102 75986 287162 76198
rect 296670 76122 296730 76198
rect 306422 76198 316050 76258
rect 296670 76062 306298 76122
rect 286918 75926 287162 75986
rect 306238 75986 306298 76062
rect 306422 75986 306482 76198
rect 315990 76122 316050 76198
rect 325742 76198 335370 76258
rect 315990 76062 325618 76122
rect 306238 75926 306482 75986
rect 325558 75986 325618 76062
rect 325742 75986 325802 76198
rect 335310 76122 335370 76198
rect 345062 76198 354690 76258
rect 335310 76062 344938 76122
rect 325558 75926 325802 75986
rect 344878 75986 344938 76062
rect 345062 75986 345122 76198
rect 354630 76122 354690 76198
rect 364382 76198 374010 76258
rect 354630 76062 364258 76122
rect 344878 75926 345122 75986
rect 364198 75986 364258 76062
rect 364382 75986 364442 76198
rect 373950 76122 374010 76198
rect 383702 76198 393330 76258
rect 373950 76062 383578 76122
rect 364198 75926 364442 75986
rect 383518 75986 383578 76062
rect 383702 75986 383762 76198
rect 393270 76122 393330 76198
rect 403022 76198 412650 76258
rect 393270 76062 402898 76122
rect 383518 75926 383762 75986
rect 402838 75986 402898 76062
rect 403022 75986 403082 76198
rect 412590 76122 412650 76198
rect 422342 76198 431970 76258
rect 412590 76062 422218 76122
rect 402838 75926 403082 75986
rect 422158 75986 422218 76062
rect 422342 75986 422402 76198
rect 431910 76122 431970 76198
rect 441662 76198 451290 76258
rect 431910 76062 441538 76122
rect 422158 75926 422402 75986
rect 441478 75986 441538 76062
rect 441662 75986 441722 76198
rect 451230 76122 451290 76198
rect 460982 76198 470610 76258
rect 451230 76062 460858 76122
rect 441478 75926 441722 75986
rect 460798 75986 460858 76062
rect 460982 75986 461042 76198
rect 470550 76122 470610 76198
rect 480302 76198 489930 76258
rect 470550 76062 480178 76122
rect 460798 75926 461042 75986
rect 480118 75986 480178 76062
rect 480302 75986 480362 76198
rect 489870 76122 489930 76198
rect 499622 76198 509250 76258
rect 489870 76062 499498 76122
rect 480118 75926 480362 75986
rect 499438 75986 499498 76062
rect 499622 75986 499682 76198
rect 509190 76122 509250 76198
rect 518942 76198 528570 76258
rect 509190 76062 518818 76122
rect 499438 75926 499682 75986
rect 518758 75986 518818 76062
rect 518942 75986 519002 76198
rect 528510 76122 528570 76198
rect 538262 76198 547890 76258
rect 528510 76062 538138 76122
rect 518758 75926 519002 75986
rect 538078 75986 538138 76062
rect 538262 75986 538322 76198
rect 547830 76122 547890 76198
rect 557582 76198 567210 76258
rect 547830 76062 557458 76122
rect 538078 75926 538322 75986
rect 557398 75986 557458 76062
rect 557582 75986 557642 76198
rect 567150 76122 567210 76198
rect 583342 76198 584960 76258
rect 583342 76122 583402 76198
rect 567150 76062 576778 76122
rect 557398 75926 557642 75986
rect 576718 75986 576778 76062
rect 576902 76062 583402 76122
rect 583520 76108 584960 76198
rect 576902 75986 576962 76062
rect 576718 75926 576962 75986
rect 140037 75923 140103 75926
rect -960 64562 480 64652
rect 3325 64562 3391 64565
rect -960 64560 3391 64562
rect -960 64504 3330 64560
rect 3386 64504 3391 64560
rect -960 64502 3391 64504
rect -960 64412 480 64502
rect 3325 64499 3391 64502
rect 579797 64562 579863 64565
rect 583520 64562 584960 64652
rect 579797 64560 584960 64562
rect 579797 64504 579802 64560
rect 579858 64504 584960 64560
rect 579797 64502 584960 64504
rect 579797 64499 579863 64502
rect 583520 64412 584960 64502
rect 583520 52716 584960 52956
rect -960 50146 480 50236
rect 3417 50146 3483 50149
rect -960 50144 3483 50146
rect -960 50088 3422 50144
rect 3478 50088 3483 50144
rect -960 50086 3483 50088
rect -960 49996 480 50086
rect 3417 50083 3483 50086
rect 580165 41034 580231 41037
rect 583520 41034 584960 41124
rect 580165 41032 584960 41034
rect 580165 40976 580170 41032
rect 580226 40976 584960 41032
rect 580165 40974 584960 40976
rect 580165 40971 580231 40974
rect 583520 40884 584960 40974
rect -960 35866 480 35956
rect 3417 35866 3483 35869
rect -960 35864 3483 35866
rect -960 35808 3422 35864
rect 3478 35808 3483 35864
rect -960 35806 3483 35808
rect -960 35716 480 35806
rect 3417 35803 3483 35806
rect 89294 31724 89300 31788
rect 89364 31786 89370 31788
rect 89529 31786 89595 31789
rect 89364 31784 89595 31786
rect 89364 31728 89534 31784
rect 89590 31728 89595 31784
rect 89364 31726 89595 31728
rect 89364 31724 89370 31726
rect 89529 31723 89595 31726
rect 580165 29338 580231 29341
rect 583520 29338 584960 29428
rect 580165 29336 584960 29338
rect 580165 29280 580170 29336
rect 580226 29280 584960 29336
rect 580165 29278 584960 29280
rect 580165 29275 580231 29278
rect 583520 29188 584960 29278
rect 89253 26348 89319 26349
rect 89253 26346 89300 26348
rect 89208 26344 89300 26346
rect 89208 26288 89258 26344
rect 89208 26286 89300 26288
rect 89253 26284 89300 26286
rect 89364 26284 89370 26348
rect 89253 26283 89319 26284
rect -960 21450 480 21540
rect 2865 21450 2931 21453
rect -960 21448 2931 21450
rect -960 21392 2870 21448
rect 2926 21392 2931 21448
rect -960 21390 2931 21392
rect -960 21300 480 21390
rect 2865 21387 2931 21390
rect 579797 17642 579863 17645
rect 583520 17642 584960 17732
rect 579797 17640 584960 17642
rect 579797 17584 579802 17640
rect 579858 17584 584960 17640
rect 579797 17582 584960 17584
rect 579797 17579 579863 17582
rect 583520 17492 584960 17582
rect -960 7170 480 7260
rect 3417 7170 3483 7173
rect -960 7168 3483 7170
rect -960 7112 3422 7168
rect 3478 7112 3483 7168
rect -960 7110 3483 7112
rect -960 7020 480 7110
rect 3417 7107 3483 7110
rect 583520 5796 584960 6036
rect 90909 5266 90975 5269
rect 208393 5266 208459 5269
rect 90909 5264 208459 5266
rect 90909 5208 90914 5264
rect 90970 5208 208398 5264
rect 208454 5208 208459 5264
rect 90909 5206 208459 5208
rect 90909 5203 90975 5206
rect 208393 5203 208459 5206
rect 81985 5130 82051 5133
rect 86861 5130 86927 5133
rect 81985 5128 86927 5130
rect 81985 5072 81990 5128
rect 82046 5072 86866 5128
rect 86922 5072 86927 5128
rect 81985 5070 86927 5072
rect 81985 5067 82051 5070
rect 86861 5067 86927 5070
rect 94497 5130 94563 5133
rect 213913 5130 213979 5133
rect 94497 5128 213979 5130
rect 94497 5072 94502 5128
rect 94558 5072 213918 5128
rect 213974 5072 213979 5128
rect 94497 5070 213979 5072
rect 94497 5067 94563 5070
rect 213913 5067 213979 5070
rect 81985 4994 82051 4997
rect 86769 4994 86835 4997
rect 81985 4992 86835 4994
rect 81985 4936 81990 4992
rect 82046 4936 86774 4992
rect 86830 4936 86835 4992
rect 81985 4934 86835 4936
rect 81985 4931 82051 4934
rect 86769 4931 86835 4934
rect 101581 4994 101647 4997
rect 226333 4994 226399 4997
rect 101581 4992 226399 4994
rect 101581 4936 101586 4992
rect 101642 4936 226338 4992
rect 226394 4936 226399 4992
rect 101581 4934 226399 4936
rect 101581 4931 101647 4934
rect 226333 4931 226399 4934
rect 78857 4858 78923 4861
rect 86861 4858 86927 4861
rect 78857 4856 86927 4858
rect 78857 4800 78862 4856
rect 78918 4800 86866 4856
rect 86922 4800 86927 4856
rect 78857 4798 86927 4800
rect 78857 4795 78923 4798
rect 86861 4795 86927 4798
rect 131389 4858 131455 4861
rect 274633 4858 274699 4861
rect 131389 4856 274699 4858
rect 131389 4800 131394 4856
rect 131450 4800 274638 4856
rect 274694 4800 274699 4856
rect 131389 4798 274699 4800
rect 131389 4795 131455 4798
rect 274633 4795 274699 4798
rect 71773 4178 71839 4181
rect 73061 4178 73127 4181
rect 71773 4176 73127 4178
rect 71773 4120 71778 4176
rect 71834 4120 73066 4176
rect 73122 4120 73127 4176
rect 71773 4118 73127 4120
rect 71773 4115 71839 4118
rect 73061 4115 73127 4118
rect 86033 4178 86099 4181
rect 89529 4178 89595 4181
rect 86033 4176 89595 4178
rect 86033 4120 86038 4176
rect 86094 4120 89534 4176
rect 89590 4120 89595 4176
rect 86033 4118 89595 4120
rect 86033 4115 86099 4118
rect 89529 4115 89595 4118
rect 77845 4042 77911 4045
rect 80053 4042 80119 4045
rect 77845 4040 80119 4042
rect 77845 3984 77850 4040
rect 77906 3984 80058 4040
rect 80114 3984 80119 4040
rect 77845 3982 80119 3984
rect 77845 3979 77911 3982
rect 80053 3979 80119 3982
rect 89437 3906 89503 3909
rect 89897 3906 89963 3909
rect 89437 3904 89963 3906
rect 89437 3848 89442 3904
rect 89498 3848 89902 3904
rect 89958 3848 89963 3904
rect 89437 3846 89963 3848
rect 89437 3843 89503 3846
rect 89897 3843 89963 3846
rect 93209 3906 93275 3909
rect 93853 3906 93919 3909
rect 93209 3904 93919 3906
rect 93209 3848 93214 3904
rect 93270 3848 93858 3904
rect 93914 3848 93919 3904
rect 93209 3846 93919 3848
rect 93209 3843 93275 3846
rect 93853 3843 93919 3846
rect 95509 3906 95575 3909
rect 96613 3906 96679 3909
rect 95509 3904 96679 3906
rect 95509 3848 95514 3904
rect 95570 3848 96618 3904
rect 96674 3848 96679 3904
rect 95509 3846 96679 3848
rect 95509 3843 95575 3846
rect 96613 3843 96679 3846
rect 102593 3906 102659 3909
rect 103513 3906 103579 3909
rect 102593 3904 103579 3906
rect 102593 3848 102598 3904
rect 102654 3848 103518 3904
rect 103574 3848 103579 3904
rect 102593 3846 103579 3848
rect 102593 3843 102659 3846
rect 103513 3843 103579 3846
rect 75453 3770 75519 3773
rect 183553 3770 183619 3773
rect 75453 3768 183619 3770
rect 75453 3712 75458 3768
rect 75514 3712 183558 3768
rect 183614 3712 183619 3768
rect 75453 3710 183619 3712
rect 75453 3707 75519 3710
rect 183553 3707 183619 3710
rect 92105 3634 92171 3637
rect 209773 3634 209839 3637
rect 92105 3632 209839 3634
rect 92105 3576 92110 3632
rect 92166 3576 209778 3632
rect 209834 3576 209839 3632
rect 92105 3574 209839 3576
rect 92105 3571 92171 3574
rect 209773 3571 209839 3574
rect 99281 3498 99347 3501
rect 222193 3498 222259 3501
rect 99281 3496 222259 3498
rect 99281 3440 99286 3496
rect 99342 3440 222198 3496
rect 222254 3440 222259 3496
rect 99281 3438 222259 3440
rect 99281 3435 99347 3438
rect 222193 3435 222259 3438
rect 61009 3362 61075 3365
rect 62113 3362 62179 3365
rect 61009 3360 62179 3362
rect 61009 3304 61014 3360
rect 61070 3304 62118 3360
rect 62174 3304 62179 3360
rect 61009 3302 62179 3304
rect 61009 3299 61075 3302
rect 62113 3299 62179 3302
rect 103973 3362 104039 3365
rect 229093 3362 229159 3365
rect 103973 3360 229159 3362
rect 103973 3304 103978 3360
rect 104034 3304 229098 3360
rect 229154 3304 229159 3360
rect 103973 3302 229159 3304
rect 103973 3299 104039 3302
rect 229093 3299 229159 3302
<< via3 >>
rect 57836 700300 57900 700364
rect 550588 697308 550652 697372
rect 59124 697172 59188 697236
rect 550588 696900 550652 696964
rect 183508 686428 183572 686492
rect 376708 686428 376772 686492
rect 434668 686428 434732 686492
rect 164188 686292 164252 686356
rect 357388 686292 357452 686356
rect 550588 686292 550652 686356
rect 57652 686156 57716 686220
rect 183508 686156 183572 686220
rect 164188 685884 164252 685948
rect 299428 686156 299492 686220
rect 299428 685884 299492 685948
rect 376708 686156 376772 686220
rect 357388 685884 357452 685948
rect 434668 686020 434732 686084
rect 550588 685884 550652 685948
rect 183508 674052 183572 674116
rect 376708 674052 376772 674116
rect 357388 673916 357452 673980
rect 59308 673780 59372 673844
rect 183508 673780 183572 673844
rect 299428 673780 299492 673844
rect 299428 673508 299492 673572
rect 376708 673780 376772 673844
rect 357388 673508 357452 673572
rect 129228 652896 129292 652900
rect 129228 652840 129278 652896
rect 129278 652840 129292 652896
rect 129228 652836 129292 652840
rect 133644 652896 133708 652900
rect 133644 652840 133694 652896
rect 133694 652840 133708 652896
rect 133644 652836 133708 652840
rect 258580 652896 258644 652900
rect 258580 652840 258630 652896
rect 258630 652840 258644 652896
rect 258580 652836 258644 652840
rect 378180 652896 378244 652900
rect 378180 652840 378194 652896
rect 378194 652840 378244 652896
rect 378180 652836 378244 652840
rect 383516 652896 383580 652900
rect 383516 652840 383530 652896
rect 383530 652840 383580 652896
rect 383516 652836 383580 652840
rect 263571 651612 263635 651676
rect 376708 651340 376772 651404
rect 376708 651068 376772 651132
rect 396028 651068 396092 651132
rect 318748 650932 318812 650996
rect 58204 650796 58268 650860
rect 125548 650796 125612 650860
rect 125548 650524 125612 650588
rect 299428 650660 299492 650724
rect 318748 650524 318812 650588
rect 396028 650796 396092 650860
rect 434668 650796 434732 650860
rect 579660 650796 579724 650860
rect 299428 650388 299492 650452
rect 434668 650388 434732 650452
rect 579660 650524 579724 650588
rect 211108 559948 211172 560012
rect 328480 559812 328544 559876
rect 337700 559872 337764 559876
rect 337700 559816 337750 559872
rect 337750 559816 337764 559872
rect 337700 559812 337764 559816
rect 358848 559812 358912 559876
rect 358860 559676 358924 559740
rect 359412 559676 359476 559740
rect 351868 559268 351932 559332
rect 352236 559132 352300 559196
rect 220124 559056 220188 559060
rect 220124 559000 220138 559056
rect 220138 559000 220188 559056
rect 220124 558996 220188 559000
rect 67404 558860 67468 558924
rect 68508 558860 68572 558924
rect 70164 558860 70228 558924
rect 71636 558920 71700 558924
rect 71636 558864 71686 558920
rect 71686 558864 71700 558920
rect 71636 558860 71700 558864
rect 72372 558860 72436 558924
rect 72924 558860 72988 558924
rect 73660 558860 73724 558924
rect 74212 558920 74276 558924
rect 74212 558864 74262 558920
rect 74262 558864 74276 558920
rect 74212 558860 74276 558864
rect 74948 558920 75012 558924
rect 74948 558864 74998 558920
rect 74998 558864 75012 558920
rect 74948 558860 75012 558864
rect 75868 558860 75932 558924
rect 76788 558920 76852 558924
rect 76788 558864 76838 558920
rect 76838 558864 76852 558920
rect 76788 558860 76852 558864
rect 77340 558920 77404 558924
rect 77340 558864 77390 558920
rect 77390 558864 77404 558920
rect 77340 558860 77404 558864
rect 78444 558920 78508 558924
rect 78444 558864 78494 558920
rect 78494 558864 78508 558920
rect 78444 558860 78508 558864
rect 79180 558860 79244 558924
rect 79916 558920 79980 558924
rect 79916 558864 79966 558920
rect 79966 558864 79980 558920
rect 79916 558860 79980 558864
rect 80652 558860 80716 558924
rect 81204 558920 81268 558924
rect 81204 558864 81254 558920
rect 81254 558864 81268 558920
rect 81204 558860 81268 558864
rect 81940 558920 82004 558924
rect 81940 558864 81954 558920
rect 81954 558864 82004 558920
rect 81940 558860 82004 558864
rect 82676 558920 82740 558924
rect 82676 558864 82726 558920
rect 82726 558864 82740 558920
rect 82676 558860 82740 558864
rect 83780 558920 83844 558924
rect 83780 558864 83830 558920
rect 83830 558864 83844 558920
rect 83780 558860 83844 558864
rect 84148 558920 84212 558924
rect 84148 558864 84198 558920
rect 84198 558864 84212 558920
rect 84148 558860 84212 558864
rect 85068 558860 85132 558924
rect 86356 558920 86420 558924
rect 86356 558864 86406 558920
rect 86406 558864 86420 558920
rect 86356 558860 86420 558864
rect 86724 558860 86788 558924
rect 87828 558920 87892 558924
rect 87828 558864 87878 558920
rect 87878 558864 87892 558920
rect 87828 558860 87892 558864
rect 88196 558920 88260 558924
rect 88196 558864 88246 558920
rect 88246 558864 88260 558920
rect 88196 558860 88260 558864
rect 88932 558920 88996 558924
rect 88932 558864 88946 558920
rect 88946 558864 88996 558920
rect 88932 558860 88996 558864
rect 89116 558860 89180 558924
rect 89852 558920 89916 558924
rect 89852 558864 89866 558920
rect 89866 558864 89916 558920
rect 89852 558860 89916 558864
rect 90956 558920 91020 558924
rect 90956 558864 91006 558920
rect 91006 558864 91020 558920
rect 90956 558860 91020 558864
rect 92428 558920 92492 558924
rect 92428 558864 92478 558920
rect 92478 558864 92492 558920
rect 92428 558860 92492 558864
rect 93164 558860 93228 558924
rect 94820 558920 94884 558924
rect 94820 558864 94870 558920
rect 94870 558864 94884 558920
rect 94820 558860 94884 558864
rect 95004 558860 95068 558924
rect 95740 558920 95804 558924
rect 95740 558864 95790 558920
rect 95790 558864 95804 558920
rect 95740 558860 95804 558864
rect 96476 558920 96540 558924
rect 96476 558864 96526 558920
rect 96526 558864 96540 558920
rect 96476 558860 96540 558864
rect 97028 558920 97092 558924
rect 97028 558864 97042 558920
rect 97042 558864 97092 558920
rect 97028 558860 97092 558864
rect 97764 558920 97828 558924
rect 97764 558864 97814 558920
rect 97814 558864 97828 558920
rect 97764 558860 97828 558864
rect 98132 558920 98196 558924
rect 98132 558864 98146 558920
rect 98146 558864 98196 558920
rect 98132 558860 98196 558864
rect 99052 558860 99116 558924
rect 99604 558920 99668 558924
rect 99604 558864 99618 558920
rect 99618 558864 99668 558920
rect 99604 558860 99668 558864
rect 100156 558860 100220 558924
rect 101444 558860 101508 558924
rect 103284 558860 103348 558924
rect 104756 558920 104820 558924
rect 104756 558864 104806 558920
rect 104806 558864 104820 558920
rect 104756 558860 104820 558864
rect 105308 558860 105372 558924
rect 106044 558860 106108 558924
rect 107148 558860 107212 558924
rect 108436 558920 108500 558924
rect 108436 558864 108486 558920
rect 108486 558864 108500 558920
rect 108436 558860 108500 558864
rect 109540 558860 109604 558924
rect 196204 558860 196268 558924
rect 197492 558860 197556 558924
rect 201724 558860 201788 558924
rect 202644 558860 202708 558924
rect 203932 558860 203996 558924
rect 205404 558860 205468 558924
rect 206140 558920 206204 558924
rect 206140 558864 206154 558920
rect 206154 558864 206204 558920
rect 206140 558860 206204 558864
rect 208348 558920 208412 558924
rect 208348 558864 208398 558920
rect 208398 558864 208412 558920
rect 208348 558860 208412 558864
rect 210556 558920 210620 558924
rect 210556 558864 210606 558920
rect 210606 558864 210620 558920
rect 210556 558860 210620 558864
rect 211844 558920 211908 558924
rect 211844 558864 211858 558920
rect 211858 558864 211908 558920
rect 211844 558860 211908 558864
rect 213132 558920 213196 558924
rect 213132 558864 213146 558920
rect 213146 558864 213196 558920
rect 213132 558860 213196 558864
rect 214052 558860 214116 558924
rect 215340 558920 215404 558924
rect 215340 558864 215354 558920
rect 215354 558864 215404 558920
rect 215340 558860 215404 558864
rect 217548 558860 217612 558924
rect 218836 558860 218900 558924
rect 222332 558920 222396 558924
rect 222332 558864 222382 558920
rect 222382 558864 222396 558920
rect 222332 558860 222396 558864
rect 223620 558920 223684 558924
rect 223620 558864 223634 558920
rect 223634 558864 223684 558920
rect 223620 558860 223684 558864
rect 224540 558920 224604 558924
rect 224540 558864 224554 558920
rect 224554 558864 224604 558920
rect 224540 558860 224604 558864
rect 225828 558920 225892 558924
rect 225828 558864 225878 558920
rect 225878 558864 225892 558920
rect 225828 558860 225892 558864
rect 227116 558920 227180 558924
rect 227116 558864 227166 558920
rect 227166 558864 227180 558920
rect 227116 558860 227180 558864
rect 228220 558920 228284 558924
rect 228220 558864 228234 558920
rect 228234 558864 228284 558920
rect 228220 558860 228284 558864
rect 229508 558920 229572 558924
rect 229508 558864 229558 558920
rect 229558 558864 229572 558920
rect 229508 558860 229572 558864
rect 313412 558920 313476 558924
rect 313412 558864 313426 558920
rect 313426 558864 313476 558920
rect 313412 558860 313476 558864
rect 322796 558860 322860 558924
rect 324084 558860 324148 558924
rect 325188 558860 325252 558924
rect 326292 558860 326356 558924
rect 327580 558860 327644 558924
rect 329604 558860 329668 558924
rect 329788 558920 329852 558924
rect 329788 558864 329838 558920
rect 329838 558864 329852 558920
rect 329788 558860 329852 558864
rect 330524 558920 330588 558924
rect 330524 558864 330538 558920
rect 330538 558864 330588 558920
rect 330524 558860 330588 558864
rect 332364 558860 332428 558924
rect 333284 558860 333348 558924
rect 334572 558860 334636 558924
rect 335860 558860 335924 558924
rect 336780 558920 336844 558924
rect 336780 558864 336794 558920
rect 336794 558864 336844 558920
rect 336780 558860 336844 558864
rect 339172 558860 339236 558924
rect 340460 558860 340524 558924
rect 341196 558920 341260 558924
rect 341196 558864 341246 558920
rect 341246 558864 341260 558920
rect 341196 558860 341260 558864
rect 342484 558920 342548 558924
rect 342484 558864 342534 558920
rect 342534 558864 342548 558920
rect 342484 558860 342548 558864
rect 343588 558920 343652 558924
rect 343588 558864 343638 558920
rect 343638 558864 343652 558920
rect 343588 558860 343652 558864
rect 344692 558860 344756 558924
rect 345796 558920 345860 558924
rect 345796 558864 345810 558920
rect 345810 558864 345860 558920
rect 345796 558860 345860 558864
rect 346900 558920 346964 558924
rect 346900 558864 346914 558920
rect 346914 558864 346964 558920
rect 346900 558860 346964 558864
rect 348188 558920 348252 558924
rect 348188 558864 348238 558920
rect 348238 558864 348252 558920
rect 348188 558860 348252 558864
rect 349476 558920 349540 558924
rect 349476 558864 349526 558920
rect 349526 558864 349540 558920
rect 349476 558860 349540 558864
rect 358860 558860 358924 558924
rect 64276 558724 64340 558788
rect 194364 558784 194428 558788
rect 194364 558728 194414 558784
rect 194414 558728 194428 558784
rect 194364 558724 194428 558728
rect 203748 558724 203812 558788
rect 216628 558724 216692 558788
rect 232820 558724 232884 558788
rect 233556 558724 233620 558788
rect 322244 558784 322308 558788
rect 322244 558728 322258 558784
rect 322258 558728 322308 558784
rect 322244 558724 322308 558728
rect 323532 558784 323596 558788
rect 323532 558728 323582 558784
rect 323582 558728 323596 558784
rect 323532 558724 323596 558728
rect 324820 558724 324884 558788
rect 326108 558724 326172 558788
rect 327028 558724 327092 558788
rect 331076 558724 331140 558788
rect 331812 558784 331876 558788
rect 331812 558728 331826 558784
rect 331826 558728 331876 558784
rect 331812 558724 331876 558728
rect 332732 558784 332796 558788
rect 332732 558728 332746 558784
rect 332746 558728 332796 558784
rect 332732 558724 332796 558728
rect 334020 558784 334084 558788
rect 334020 558728 334070 558784
rect 334070 558728 334084 558784
rect 334020 558724 334084 558728
rect 335492 558784 335556 558788
rect 335492 558728 335506 558784
rect 335506 558728 335556 558784
rect 335492 558724 335556 558728
rect 336596 558724 336660 558788
rect 338988 558784 339052 558788
rect 338988 558728 339038 558784
rect 339038 558728 339052 558784
rect 338988 558724 339052 558728
rect 339908 558784 339972 558788
rect 339908 558728 339922 558784
rect 339922 558728 339972 558784
rect 339908 558724 339972 558728
rect 353524 558724 353588 558788
rect 354812 558724 354876 558788
rect 356100 558784 356164 558788
rect 356100 558728 356114 558784
rect 356114 558728 356164 558784
rect 356100 558724 356164 558728
rect 69796 558588 69860 558652
rect 79364 558588 79428 558652
rect 82860 558648 82924 558652
rect 82860 558592 82874 558648
rect 82874 558592 82924 558648
rect 82860 558588 82924 558592
rect 85436 558588 85500 558652
rect 86172 558588 86236 558652
rect 91140 558648 91204 558652
rect 91140 558592 91154 558648
rect 91154 558592 91204 558648
rect 91140 558588 91204 558592
rect 93348 558648 93412 558652
rect 93348 558592 93362 558648
rect 93362 558592 93412 558648
rect 93348 558588 93412 558592
rect 93716 558648 93780 558652
rect 93716 558592 93766 558648
rect 93766 558592 93780 558648
rect 93716 558588 93780 558592
rect 100340 558588 100404 558652
rect 101996 558648 102060 558652
rect 101996 558592 102010 558648
rect 102010 558592 102060 558648
rect 101996 558588 102060 558592
rect 102732 558648 102796 558652
rect 102732 558592 102782 558648
rect 102782 558592 102796 558648
rect 102732 558588 102796 558592
rect 104020 558588 104084 558652
rect 106228 558588 106292 558652
rect 107700 558648 107764 558652
rect 107700 558592 107750 558648
rect 107750 558592 107764 558648
rect 107700 558588 107764 558592
rect 108620 558588 108684 558652
rect 202460 558588 202524 558652
rect 204852 558648 204916 558652
rect 204852 558592 204902 558648
rect 204902 558592 204916 558648
rect 204852 558588 204916 558592
rect 209636 558588 209700 558652
rect 235028 558588 235092 558652
rect 237420 558648 237484 558652
rect 237420 558592 237434 558648
rect 237434 558592 237484 558648
rect 237420 558588 237484 558592
rect 282316 558588 282380 558652
rect 236132 558452 236196 558516
rect 238708 558512 238772 558516
rect 238708 558456 238758 558512
rect 238758 558456 238772 558512
rect 238708 558452 238772 558456
rect 283420 558452 283484 558516
rect 350580 558512 350644 558516
rect 357940 558588 358004 558652
rect 350580 558456 350594 558512
rect 350594 558456 350644 558512
rect 350580 558452 350644 558456
rect 78076 558316 78140 558380
rect 92060 558316 92124 558380
rect 101628 558316 101692 558380
rect 221044 558316 221108 558380
rect 230612 558316 230676 558380
rect 231900 558376 231964 558380
rect 231900 558320 231914 558376
rect 231914 558320 231964 558376
rect 231900 558316 231964 558320
rect 283788 558316 283852 558380
rect 357572 558452 357636 558516
rect 75684 558180 75748 558244
rect 283604 558180 283668 558244
rect 352420 558180 352484 558244
rect 355732 558180 355796 558244
rect 317460 557968 317524 557972
rect 317460 557912 317474 557968
rect 317474 557912 317524 557968
rect 317460 557908 317524 557912
rect 320588 557908 320652 557972
rect 337884 557908 337948 557972
rect 200252 557832 200316 557836
rect 200252 557776 200266 557832
rect 200266 557776 200316 557832
rect 200252 557772 200316 557776
rect 198780 557696 198844 557700
rect 198780 557640 198794 557696
rect 198794 557640 198844 557696
rect 198780 557636 198844 557640
rect 207060 557636 207124 557700
rect 210372 557636 210436 557700
rect 217364 557636 217428 557700
rect 225644 557636 225708 557700
rect 232636 557636 232700 557700
rect 344876 557636 344940 557700
rect 353156 558044 353220 558108
rect 354444 557908 354508 557972
rect 356652 557636 356716 557700
rect 206876 557560 206940 557564
rect 206876 557504 206926 557560
rect 206926 557504 206940 557560
rect 206876 557500 206940 557504
rect 207980 557500 208044 557564
rect 209268 557500 209332 557564
rect 212396 557560 212460 557564
rect 212396 557504 212446 557560
rect 212446 557504 212460 557560
rect 212396 557500 212460 557504
rect 213500 557500 213564 557564
rect 214788 557500 214852 557564
rect 216260 557500 216324 557564
rect 217916 557560 217980 557564
rect 217916 557504 217966 557560
rect 217966 557504 217980 557560
rect 217916 557500 217980 557504
rect 219204 557500 219268 557564
rect 220676 557560 220740 557564
rect 220676 557504 220726 557560
rect 220726 557504 220740 557560
rect 220676 557500 220740 557504
rect 221964 557500 222028 557564
rect 223252 557500 223316 557564
rect 224356 557500 224420 557564
rect 226196 557560 226260 557564
rect 226196 557504 226246 557560
rect 226246 557504 226260 557560
rect 226196 557500 226260 557504
rect 227484 557500 227548 557564
rect 228772 557500 228836 557564
rect 230244 557500 230308 557564
rect 230796 557500 230860 557564
rect 233004 557560 233068 557564
rect 233004 557504 233054 557560
rect 233054 557504 233068 557560
rect 233004 557500 233068 557504
rect 234476 557560 234540 557564
rect 234476 557504 234526 557560
rect 234526 557504 234540 557560
rect 234476 557500 234540 557504
rect 235764 557500 235828 557564
rect 237236 557560 237300 557564
rect 237236 557504 237286 557560
rect 237286 557504 237300 557560
rect 237236 557500 237300 557504
rect 238340 557500 238404 557564
rect 239628 557500 239692 557564
rect 316356 557500 316420 557564
rect 318932 557500 318996 557564
rect 320956 557500 321020 557564
rect 341748 557500 341812 557564
rect 342668 557500 342732 557564
rect 343956 557500 344020 557564
rect 346164 557500 346228 557564
rect 347452 557500 347516 557564
rect 348740 557500 348804 557564
rect 349660 557500 349724 557564
rect 350948 557500 351012 557564
rect 328868 557092 328932 557156
rect 57468 545532 57532 545596
rect 75868 545124 75932 545188
rect 347820 545396 347884 545460
rect 550588 545532 550652 545596
rect 376708 545396 376772 545460
rect 347820 545124 347884 545188
rect 357388 545124 357452 545188
rect 376708 545124 376772 545188
rect 492628 545396 492692 545460
rect 492628 545124 492692 545188
rect 550588 545124 550652 545188
rect 75868 544852 75932 544916
rect 357388 544852 357452 544916
rect 59492 540364 59556 540428
rect 57284 540228 57348 540292
rect 281580 413884 281644 413948
rect 367692 413884 367756 413948
rect 368980 413884 369044 413948
rect 370268 413884 370332 413948
rect 371556 413884 371620 413948
rect 372660 413944 372724 413948
rect 372660 413888 372674 413944
rect 372674 413888 372724 413944
rect 372660 413884 372724 413888
rect 373948 413944 374012 413948
rect 373948 413888 373998 413944
rect 373998 413888 374012 413944
rect 373948 413884 374012 413888
rect 375972 413884 376036 413948
rect 377260 413884 377324 413948
rect 378364 413884 378428 413948
rect 379652 413884 379716 413948
rect 380940 413944 381004 413948
rect 380940 413888 380954 413944
rect 380954 413888 381004 413944
rect 380940 413884 381004 413888
rect 382228 413944 382292 413948
rect 382228 413888 382278 413944
rect 382278 413888 382292 413944
rect 382228 413884 382292 413888
rect 385172 413884 385236 413948
rect 374684 413748 374748 413812
rect 382964 413748 383028 413812
rect 384068 413748 384132 413812
rect 412772 413748 412836 413812
rect 396396 413612 396460 413676
rect 397500 413672 397564 413676
rect 397500 413616 397514 413672
rect 397514 413616 397564 413672
rect 397500 413612 397564 413616
rect 405780 413536 405844 413540
rect 405780 413480 405794 413536
rect 405794 413480 405844 413536
rect 405780 413476 405844 413480
rect 368244 413400 368308 413404
rect 368244 413344 368294 413400
rect 368294 413344 368308 413400
rect 368244 413340 368308 413344
rect 369716 413400 369780 413404
rect 369716 413344 369766 413400
rect 369766 413344 369780 413400
rect 369716 413340 369780 413344
rect 377996 413400 378060 413404
rect 377996 413344 378046 413400
rect 378046 413344 378060 413400
rect 377996 413340 378060 413344
rect 388300 413400 388364 413404
rect 388300 413344 388350 413400
rect 388350 413344 388364 413400
rect 388300 413340 388364 413344
rect 404676 413340 404740 413404
rect 371004 413204 371068 413268
rect 380204 413204 380268 413268
rect 386828 413204 386892 413268
rect 402284 413204 402348 413268
rect 403388 413204 403452 413268
rect 407436 413204 407500 413268
rect 371924 413128 371988 413132
rect 371924 413072 371974 413128
rect 371974 413072 371988 413128
rect 371924 413068 371988 413072
rect 373028 413128 373092 413132
rect 373028 413072 373042 413128
rect 373042 413072 373092 413128
rect 373028 413068 373092 413072
rect 378916 413068 378980 413132
rect 381492 413128 381556 413132
rect 381492 413072 381542 413128
rect 381542 413072 381556 413128
rect 381492 413068 381556 413072
rect 382412 413068 382476 413132
rect 387196 413068 387260 413132
rect 399892 413068 399956 413132
rect 408724 413068 408788 413132
rect 374316 412992 374380 412996
rect 374316 412936 374366 412992
rect 374366 412936 374380 412992
rect 374316 412932 374380 412936
rect 383516 412992 383580 412996
rect 383516 412936 383566 412992
rect 383566 412936 383580 412992
rect 383516 412932 383580 412936
rect 384804 412932 384868 412996
rect 385908 412932 385972 412996
rect 401180 412932 401244 412996
rect 375420 412856 375484 412860
rect 375420 412800 375470 412856
rect 375470 412800 375484 412856
rect 375420 412796 375484 412800
rect 376524 412856 376588 412860
rect 376524 412800 376574 412856
rect 376574 412800 376588 412856
rect 376524 412796 376588 412800
rect 393452 412796 393516 412860
rect 398604 412796 398668 412860
rect 389588 412720 389652 412724
rect 389588 412664 389638 412720
rect 389638 412664 389652 412720
rect 389588 412660 389652 412664
rect 390876 412720 390940 412724
rect 390876 412664 390926 412720
rect 390926 412664 390940 412720
rect 390876 412660 390940 412664
rect 391796 412720 391860 412724
rect 391796 412664 391810 412720
rect 391810 412664 391860 412720
rect 391796 412660 391860 412664
rect 393084 412720 393148 412724
rect 393084 412664 393134 412720
rect 393134 412664 393148 412720
rect 393084 412660 393148 412664
rect 394004 412720 394068 412724
rect 394004 412664 394018 412720
rect 394018 412664 394068 412720
rect 394004 412660 394068 412664
rect 394740 412720 394804 412724
rect 394740 412664 394754 412720
rect 394754 412664 394804 412720
rect 394740 412660 394804 412664
rect 395292 412720 395356 412724
rect 395292 412664 395342 412720
rect 395342 412664 395356 412720
rect 395292 412660 395356 412664
rect 396028 412720 396092 412724
rect 396028 412664 396078 412720
rect 396078 412664 396092 412720
rect 396028 412660 396092 412664
rect 406332 412660 406396 412724
rect 57836 411708 57900 411772
rect 388116 411768 388180 411772
rect 388116 411712 388130 411768
rect 388130 411712 388180 411768
rect 388116 411708 388180 411712
rect 391060 411632 391124 411636
rect 391060 411576 391074 411632
rect 391074 411576 391124 411632
rect 391060 411572 391124 411576
rect 397460 411632 397524 411636
rect 397460 411576 397514 411632
rect 397514 411576 397524 411632
rect 397460 411572 397524 411576
rect 399156 411632 399220 411636
rect 399156 411576 399170 411632
rect 399170 411576 399220 411632
rect 399156 411572 399220 411576
rect 389284 411496 389348 411500
rect 389284 411440 389326 411496
rect 389326 411440 389348 411496
rect 389284 411436 389348 411440
rect 398052 411496 398116 411500
rect 398052 411440 398066 411496
rect 398066 411440 398116 411496
rect 398052 411436 398116 411440
rect 400964 411496 401028 411500
rect 400964 411440 401010 411496
rect 401010 411440 401028 411496
rect 400964 411436 401028 411440
rect 403300 411496 403364 411500
rect 403300 411440 403310 411496
rect 403310 411440 403364 411496
rect 403300 411436 403364 411440
rect 401732 411360 401796 411364
rect 401732 411304 401746 411360
rect 401746 411304 401796 411360
rect 401732 411300 401796 411304
rect 404308 411360 404372 411364
rect 404308 411304 404358 411360
rect 404358 411304 404372 411360
rect 404308 411300 404372 411304
rect 389772 411088 389836 411092
rect 389772 411032 389786 411088
rect 389786 411032 389836 411088
rect 389772 411028 389836 411032
rect 392302 410408 392366 410412
rect 392302 410352 392306 410408
rect 392306 410352 392362 410408
rect 392362 410352 392366 410408
rect 392302 410348 392366 410352
rect 410012 410408 410076 410412
rect 410012 410352 410026 410408
rect 410026 410352 410076 410408
rect 410012 410348 410076 410352
rect 59492 407764 59556 407828
rect 57652 405860 57716 405924
rect 59124 403956 59188 404020
rect 59308 402052 59372 402116
rect 58204 398108 58268 398172
rect 283604 397156 283668 397220
rect 283788 396068 283852 396132
rect 283420 395116 283484 395180
rect 57284 394300 57348 394364
rect 282316 391036 282380 391100
rect 57468 388452 57532 388516
rect 57836 374988 57900 375052
rect 56916 353772 56980 353836
rect 57284 347924 57348 347988
rect 57100 346020 57164 346084
rect 57652 342212 57716 342276
rect 57468 340172 57532 340236
rect 57836 330652 57900 330716
rect 57836 330516 57900 330580
rect 343956 318744 344020 318748
rect 343956 318688 344006 318744
rect 344006 318688 344020 318744
rect 343956 318684 344020 318688
rect 348004 318412 348068 318476
rect 281580 317324 281644 317388
rect 106228 264284 106292 264348
rect 125548 264148 125612 264212
rect 86908 264012 86972 264076
rect 96476 264012 96540 264076
rect 56916 263876 56980 263940
rect 96476 263740 96540 263804
rect 106228 264012 106292 264076
rect 125548 263876 125612 263940
rect 86908 263604 86972 263668
rect 106228 228380 106292 228444
rect 125548 228244 125612 228308
rect 57100 227972 57164 228036
rect 96476 227836 96540 227900
rect 106228 228108 106292 228172
rect 125548 227972 125612 228036
rect 86908 227700 86972 227764
rect 86908 227428 86972 227492
rect 96476 227428 96540 227492
rect 125548 217228 125612 217292
rect 57284 216956 57348 217020
rect 125548 216956 125612 217020
rect 106228 181460 106292 181524
rect 57468 181052 57532 181116
rect 96476 180916 96540 180980
rect 106228 181188 106292 181252
rect 96476 180780 96540 180844
rect 106228 170444 106292 170508
rect 125548 170308 125612 170372
rect 57652 170036 57716 170100
rect 106228 170172 106292 170236
rect 125548 170036 125612 170100
rect 125548 76468 125612 76532
rect 57836 76196 57900 76260
rect 125548 76196 125612 76260
rect 89300 31724 89364 31788
rect 89300 26344 89364 26348
rect 89300 26288 89314 26344
rect 89314 26288 89364 26344
rect 89300 26284 89364 26288
<< metal4 >>
rect -8576 711418 -7976 711440
rect -8576 711182 -8394 711418
rect -8158 711182 -7976 711418
rect -8576 711098 -7976 711182
rect -8576 710862 -8394 711098
rect -8158 710862 -7976 711098
rect -8576 679254 -7976 710862
rect -8576 679018 -8394 679254
rect -8158 679018 -7976 679254
rect -8576 678934 -7976 679018
rect -8576 678698 -8394 678934
rect -8158 678698 -7976 678934
rect -8576 643254 -7976 678698
rect -8576 643018 -8394 643254
rect -8158 643018 -7976 643254
rect -8576 642934 -7976 643018
rect -8576 642698 -8394 642934
rect -8158 642698 -7976 642934
rect -8576 607254 -7976 642698
rect -8576 607018 -8394 607254
rect -8158 607018 -7976 607254
rect -8576 606934 -7976 607018
rect -8576 606698 -8394 606934
rect -8158 606698 -7976 606934
rect -8576 571254 -7976 606698
rect -8576 571018 -8394 571254
rect -8158 571018 -7976 571254
rect -8576 570934 -7976 571018
rect -8576 570698 -8394 570934
rect -8158 570698 -7976 570934
rect -8576 535254 -7976 570698
rect -8576 535018 -8394 535254
rect -8158 535018 -7976 535254
rect -8576 534934 -7976 535018
rect -8576 534698 -8394 534934
rect -8158 534698 -7976 534934
rect -8576 499254 -7976 534698
rect -8576 499018 -8394 499254
rect -8158 499018 -7976 499254
rect -8576 498934 -7976 499018
rect -8576 498698 -8394 498934
rect -8158 498698 -7976 498934
rect -8576 463254 -7976 498698
rect -8576 463018 -8394 463254
rect -8158 463018 -7976 463254
rect -8576 462934 -7976 463018
rect -8576 462698 -8394 462934
rect -8158 462698 -7976 462934
rect -8576 427254 -7976 462698
rect -8576 427018 -8394 427254
rect -8158 427018 -7976 427254
rect -8576 426934 -7976 427018
rect -8576 426698 -8394 426934
rect -8158 426698 -7976 426934
rect -8576 391254 -7976 426698
rect -8576 391018 -8394 391254
rect -8158 391018 -7976 391254
rect -8576 390934 -7976 391018
rect -8576 390698 -8394 390934
rect -8158 390698 -7976 390934
rect -8576 355254 -7976 390698
rect -8576 355018 -8394 355254
rect -8158 355018 -7976 355254
rect -8576 354934 -7976 355018
rect -8576 354698 -8394 354934
rect -8158 354698 -7976 354934
rect -8576 319254 -7976 354698
rect -8576 319018 -8394 319254
rect -8158 319018 -7976 319254
rect -8576 318934 -7976 319018
rect -8576 318698 -8394 318934
rect -8158 318698 -7976 318934
rect -8576 283254 -7976 318698
rect -8576 283018 -8394 283254
rect -8158 283018 -7976 283254
rect -8576 282934 -7976 283018
rect -8576 282698 -8394 282934
rect -8158 282698 -7976 282934
rect -8576 247254 -7976 282698
rect -8576 247018 -8394 247254
rect -8158 247018 -7976 247254
rect -8576 246934 -7976 247018
rect -8576 246698 -8394 246934
rect -8158 246698 -7976 246934
rect -8576 211254 -7976 246698
rect -8576 211018 -8394 211254
rect -8158 211018 -7976 211254
rect -8576 210934 -7976 211018
rect -8576 210698 -8394 210934
rect -8158 210698 -7976 210934
rect -8576 175254 -7976 210698
rect -8576 175018 -8394 175254
rect -8158 175018 -7976 175254
rect -8576 174934 -7976 175018
rect -8576 174698 -8394 174934
rect -8158 174698 -7976 174934
rect -8576 139254 -7976 174698
rect -8576 139018 -8394 139254
rect -8158 139018 -7976 139254
rect -8576 138934 -7976 139018
rect -8576 138698 -8394 138934
rect -8158 138698 -7976 138934
rect -8576 103254 -7976 138698
rect -8576 103018 -8394 103254
rect -8158 103018 -7976 103254
rect -8576 102934 -7976 103018
rect -8576 102698 -8394 102934
rect -8158 102698 -7976 102934
rect -8576 67254 -7976 102698
rect -8576 67018 -8394 67254
rect -8158 67018 -7976 67254
rect -8576 66934 -7976 67018
rect -8576 66698 -8394 66934
rect -8158 66698 -7976 66934
rect -8576 31254 -7976 66698
rect -8576 31018 -8394 31254
rect -8158 31018 -7976 31254
rect -8576 30934 -7976 31018
rect -8576 30698 -8394 30934
rect -8158 30698 -7976 30934
rect -8576 -6926 -7976 30698
rect -7636 710478 -7036 710500
rect -7636 710242 -7454 710478
rect -7218 710242 -7036 710478
rect -7636 710158 -7036 710242
rect -7636 709922 -7454 710158
rect -7218 709922 -7036 710158
rect -7636 697254 -7036 709922
rect 11604 710478 12204 711440
rect 11604 710242 11786 710478
rect 12022 710242 12204 710478
rect 11604 710158 12204 710242
rect 11604 709922 11786 710158
rect 12022 709922 12204 710158
rect -7636 697018 -7454 697254
rect -7218 697018 -7036 697254
rect -7636 696934 -7036 697018
rect -7636 696698 -7454 696934
rect -7218 696698 -7036 696934
rect -7636 661254 -7036 696698
rect -7636 661018 -7454 661254
rect -7218 661018 -7036 661254
rect -7636 660934 -7036 661018
rect -7636 660698 -7454 660934
rect -7218 660698 -7036 660934
rect -7636 625254 -7036 660698
rect -7636 625018 -7454 625254
rect -7218 625018 -7036 625254
rect -7636 624934 -7036 625018
rect -7636 624698 -7454 624934
rect -7218 624698 -7036 624934
rect -7636 589254 -7036 624698
rect -7636 589018 -7454 589254
rect -7218 589018 -7036 589254
rect -7636 588934 -7036 589018
rect -7636 588698 -7454 588934
rect -7218 588698 -7036 588934
rect -7636 553254 -7036 588698
rect -7636 553018 -7454 553254
rect -7218 553018 -7036 553254
rect -7636 552934 -7036 553018
rect -7636 552698 -7454 552934
rect -7218 552698 -7036 552934
rect -7636 517254 -7036 552698
rect -7636 517018 -7454 517254
rect -7218 517018 -7036 517254
rect -7636 516934 -7036 517018
rect -7636 516698 -7454 516934
rect -7218 516698 -7036 516934
rect -7636 481254 -7036 516698
rect -7636 481018 -7454 481254
rect -7218 481018 -7036 481254
rect -7636 480934 -7036 481018
rect -7636 480698 -7454 480934
rect -7218 480698 -7036 480934
rect -7636 445254 -7036 480698
rect -7636 445018 -7454 445254
rect -7218 445018 -7036 445254
rect -7636 444934 -7036 445018
rect -7636 444698 -7454 444934
rect -7218 444698 -7036 444934
rect -7636 409254 -7036 444698
rect -7636 409018 -7454 409254
rect -7218 409018 -7036 409254
rect -7636 408934 -7036 409018
rect -7636 408698 -7454 408934
rect -7218 408698 -7036 408934
rect -7636 373254 -7036 408698
rect -7636 373018 -7454 373254
rect -7218 373018 -7036 373254
rect -7636 372934 -7036 373018
rect -7636 372698 -7454 372934
rect -7218 372698 -7036 372934
rect -7636 337254 -7036 372698
rect -7636 337018 -7454 337254
rect -7218 337018 -7036 337254
rect -7636 336934 -7036 337018
rect -7636 336698 -7454 336934
rect -7218 336698 -7036 336934
rect -7636 301254 -7036 336698
rect -7636 301018 -7454 301254
rect -7218 301018 -7036 301254
rect -7636 300934 -7036 301018
rect -7636 300698 -7454 300934
rect -7218 300698 -7036 300934
rect -7636 265254 -7036 300698
rect -7636 265018 -7454 265254
rect -7218 265018 -7036 265254
rect -7636 264934 -7036 265018
rect -7636 264698 -7454 264934
rect -7218 264698 -7036 264934
rect -7636 229254 -7036 264698
rect -7636 229018 -7454 229254
rect -7218 229018 -7036 229254
rect -7636 228934 -7036 229018
rect -7636 228698 -7454 228934
rect -7218 228698 -7036 228934
rect -7636 193254 -7036 228698
rect -7636 193018 -7454 193254
rect -7218 193018 -7036 193254
rect -7636 192934 -7036 193018
rect -7636 192698 -7454 192934
rect -7218 192698 -7036 192934
rect -7636 157254 -7036 192698
rect -7636 157018 -7454 157254
rect -7218 157018 -7036 157254
rect -7636 156934 -7036 157018
rect -7636 156698 -7454 156934
rect -7218 156698 -7036 156934
rect -7636 121254 -7036 156698
rect -7636 121018 -7454 121254
rect -7218 121018 -7036 121254
rect -7636 120934 -7036 121018
rect -7636 120698 -7454 120934
rect -7218 120698 -7036 120934
rect -7636 85254 -7036 120698
rect -7636 85018 -7454 85254
rect -7218 85018 -7036 85254
rect -7636 84934 -7036 85018
rect -7636 84698 -7454 84934
rect -7218 84698 -7036 84934
rect -7636 49254 -7036 84698
rect -7636 49018 -7454 49254
rect -7218 49018 -7036 49254
rect -7636 48934 -7036 49018
rect -7636 48698 -7454 48934
rect -7218 48698 -7036 48934
rect -7636 13254 -7036 48698
rect -7636 13018 -7454 13254
rect -7218 13018 -7036 13254
rect -7636 12934 -7036 13018
rect -7636 12698 -7454 12934
rect -7218 12698 -7036 12934
rect -7636 -5986 -7036 12698
rect -6696 709538 -6096 709560
rect -6696 709302 -6514 709538
rect -6278 709302 -6096 709538
rect -6696 709218 -6096 709302
rect -6696 708982 -6514 709218
rect -6278 708982 -6096 709218
rect -6696 675654 -6096 708982
rect -6696 675418 -6514 675654
rect -6278 675418 -6096 675654
rect -6696 675334 -6096 675418
rect -6696 675098 -6514 675334
rect -6278 675098 -6096 675334
rect -6696 639654 -6096 675098
rect -6696 639418 -6514 639654
rect -6278 639418 -6096 639654
rect -6696 639334 -6096 639418
rect -6696 639098 -6514 639334
rect -6278 639098 -6096 639334
rect -6696 603654 -6096 639098
rect -6696 603418 -6514 603654
rect -6278 603418 -6096 603654
rect -6696 603334 -6096 603418
rect -6696 603098 -6514 603334
rect -6278 603098 -6096 603334
rect -6696 567654 -6096 603098
rect -6696 567418 -6514 567654
rect -6278 567418 -6096 567654
rect -6696 567334 -6096 567418
rect -6696 567098 -6514 567334
rect -6278 567098 -6096 567334
rect -6696 531654 -6096 567098
rect -6696 531418 -6514 531654
rect -6278 531418 -6096 531654
rect -6696 531334 -6096 531418
rect -6696 531098 -6514 531334
rect -6278 531098 -6096 531334
rect -6696 495654 -6096 531098
rect -6696 495418 -6514 495654
rect -6278 495418 -6096 495654
rect -6696 495334 -6096 495418
rect -6696 495098 -6514 495334
rect -6278 495098 -6096 495334
rect -6696 459654 -6096 495098
rect -6696 459418 -6514 459654
rect -6278 459418 -6096 459654
rect -6696 459334 -6096 459418
rect -6696 459098 -6514 459334
rect -6278 459098 -6096 459334
rect -6696 423654 -6096 459098
rect -6696 423418 -6514 423654
rect -6278 423418 -6096 423654
rect -6696 423334 -6096 423418
rect -6696 423098 -6514 423334
rect -6278 423098 -6096 423334
rect -6696 387654 -6096 423098
rect -6696 387418 -6514 387654
rect -6278 387418 -6096 387654
rect -6696 387334 -6096 387418
rect -6696 387098 -6514 387334
rect -6278 387098 -6096 387334
rect -6696 351654 -6096 387098
rect -6696 351418 -6514 351654
rect -6278 351418 -6096 351654
rect -6696 351334 -6096 351418
rect -6696 351098 -6514 351334
rect -6278 351098 -6096 351334
rect -6696 315654 -6096 351098
rect -6696 315418 -6514 315654
rect -6278 315418 -6096 315654
rect -6696 315334 -6096 315418
rect -6696 315098 -6514 315334
rect -6278 315098 -6096 315334
rect -6696 279654 -6096 315098
rect -6696 279418 -6514 279654
rect -6278 279418 -6096 279654
rect -6696 279334 -6096 279418
rect -6696 279098 -6514 279334
rect -6278 279098 -6096 279334
rect -6696 243654 -6096 279098
rect -6696 243418 -6514 243654
rect -6278 243418 -6096 243654
rect -6696 243334 -6096 243418
rect -6696 243098 -6514 243334
rect -6278 243098 -6096 243334
rect -6696 207654 -6096 243098
rect -6696 207418 -6514 207654
rect -6278 207418 -6096 207654
rect -6696 207334 -6096 207418
rect -6696 207098 -6514 207334
rect -6278 207098 -6096 207334
rect -6696 171654 -6096 207098
rect -6696 171418 -6514 171654
rect -6278 171418 -6096 171654
rect -6696 171334 -6096 171418
rect -6696 171098 -6514 171334
rect -6278 171098 -6096 171334
rect -6696 135654 -6096 171098
rect -6696 135418 -6514 135654
rect -6278 135418 -6096 135654
rect -6696 135334 -6096 135418
rect -6696 135098 -6514 135334
rect -6278 135098 -6096 135334
rect -6696 99654 -6096 135098
rect -6696 99418 -6514 99654
rect -6278 99418 -6096 99654
rect -6696 99334 -6096 99418
rect -6696 99098 -6514 99334
rect -6278 99098 -6096 99334
rect -6696 63654 -6096 99098
rect -6696 63418 -6514 63654
rect -6278 63418 -6096 63654
rect -6696 63334 -6096 63418
rect -6696 63098 -6514 63334
rect -6278 63098 -6096 63334
rect -6696 27654 -6096 63098
rect -6696 27418 -6514 27654
rect -6278 27418 -6096 27654
rect -6696 27334 -6096 27418
rect -6696 27098 -6514 27334
rect -6278 27098 -6096 27334
rect -6696 -5046 -6096 27098
rect -5756 708598 -5156 708620
rect -5756 708362 -5574 708598
rect -5338 708362 -5156 708598
rect -5756 708278 -5156 708362
rect -5756 708042 -5574 708278
rect -5338 708042 -5156 708278
rect -5756 693654 -5156 708042
rect 8004 708598 8604 709560
rect 8004 708362 8186 708598
rect 8422 708362 8604 708598
rect 8004 708278 8604 708362
rect 8004 708042 8186 708278
rect 8422 708042 8604 708278
rect -5756 693418 -5574 693654
rect -5338 693418 -5156 693654
rect -5756 693334 -5156 693418
rect -5756 693098 -5574 693334
rect -5338 693098 -5156 693334
rect -5756 657654 -5156 693098
rect -5756 657418 -5574 657654
rect -5338 657418 -5156 657654
rect -5756 657334 -5156 657418
rect -5756 657098 -5574 657334
rect -5338 657098 -5156 657334
rect -5756 621654 -5156 657098
rect -5756 621418 -5574 621654
rect -5338 621418 -5156 621654
rect -5756 621334 -5156 621418
rect -5756 621098 -5574 621334
rect -5338 621098 -5156 621334
rect -5756 585654 -5156 621098
rect -5756 585418 -5574 585654
rect -5338 585418 -5156 585654
rect -5756 585334 -5156 585418
rect -5756 585098 -5574 585334
rect -5338 585098 -5156 585334
rect -5756 549654 -5156 585098
rect -5756 549418 -5574 549654
rect -5338 549418 -5156 549654
rect -5756 549334 -5156 549418
rect -5756 549098 -5574 549334
rect -5338 549098 -5156 549334
rect -5756 513654 -5156 549098
rect -5756 513418 -5574 513654
rect -5338 513418 -5156 513654
rect -5756 513334 -5156 513418
rect -5756 513098 -5574 513334
rect -5338 513098 -5156 513334
rect -5756 477654 -5156 513098
rect -5756 477418 -5574 477654
rect -5338 477418 -5156 477654
rect -5756 477334 -5156 477418
rect -5756 477098 -5574 477334
rect -5338 477098 -5156 477334
rect -5756 441654 -5156 477098
rect -5756 441418 -5574 441654
rect -5338 441418 -5156 441654
rect -5756 441334 -5156 441418
rect -5756 441098 -5574 441334
rect -5338 441098 -5156 441334
rect -5756 405654 -5156 441098
rect -5756 405418 -5574 405654
rect -5338 405418 -5156 405654
rect -5756 405334 -5156 405418
rect -5756 405098 -5574 405334
rect -5338 405098 -5156 405334
rect -5756 369654 -5156 405098
rect -5756 369418 -5574 369654
rect -5338 369418 -5156 369654
rect -5756 369334 -5156 369418
rect -5756 369098 -5574 369334
rect -5338 369098 -5156 369334
rect -5756 333654 -5156 369098
rect -5756 333418 -5574 333654
rect -5338 333418 -5156 333654
rect -5756 333334 -5156 333418
rect -5756 333098 -5574 333334
rect -5338 333098 -5156 333334
rect -5756 297654 -5156 333098
rect -5756 297418 -5574 297654
rect -5338 297418 -5156 297654
rect -5756 297334 -5156 297418
rect -5756 297098 -5574 297334
rect -5338 297098 -5156 297334
rect -5756 261654 -5156 297098
rect -5756 261418 -5574 261654
rect -5338 261418 -5156 261654
rect -5756 261334 -5156 261418
rect -5756 261098 -5574 261334
rect -5338 261098 -5156 261334
rect -5756 225654 -5156 261098
rect -5756 225418 -5574 225654
rect -5338 225418 -5156 225654
rect -5756 225334 -5156 225418
rect -5756 225098 -5574 225334
rect -5338 225098 -5156 225334
rect -5756 189654 -5156 225098
rect -5756 189418 -5574 189654
rect -5338 189418 -5156 189654
rect -5756 189334 -5156 189418
rect -5756 189098 -5574 189334
rect -5338 189098 -5156 189334
rect -5756 153654 -5156 189098
rect -5756 153418 -5574 153654
rect -5338 153418 -5156 153654
rect -5756 153334 -5156 153418
rect -5756 153098 -5574 153334
rect -5338 153098 -5156 153334
rect -5756 117654 -5156 153098
rect -5756 117418 -5574 117654
rect -5338 117418 -5156 117654
rect -5756 117334 -5156 117418
rect -5756 117098 -5574 117334
rect -5338 117098 -5156 117334
rect -5756 81654 -5156 117098
rect -5756 81418 -5574 81654
rect -5338 81418 -5156 81654
rect -5756 81334 -5156 81418
rect -5756 81098 -5574 81334
rect -5338 81098 -5156 81334
rect -5756 45654 -5156 81098
rect -5756 45418 -5574 45654
rect -5338 45418 -5156 45654
rect -5756 45334 -5156 45418
rect -5756 45098 -5574 45334
rect -5338 45098 -5156 45334
rect -5756 9654 -5156 45098
rect -5756 9418 -5574 9654
rect -5338 9418 -5156 9654
rect -5756 9334 -5156 9418
rect -5756 9098 -5574 9334
rect -5338 9098 -5156 9334
rect -5756 -4106 -5156 9098
rect -4816 707658 -4216 707680
rect -4816 707422 -4634 707658
rect -4398 707422 -4216 707658
rect -4816 707338 -4216 707422
rect -4816 707102 -4634 707338
rect -4398 707102 -4216 707338
rect -4816 672054 -4216 707102
rect -4816 671818 -4634 672054
rect -4398 671818 -4216 672054
rect -4816 671734 -4216 671818
rect -4816 671498 -4634 671734
rect -4398 671498 -4216 671734
rect -4816 636054 -4216 671498
rect -4816 635818 -4634 636054
rect -4398 635818 -4216 636054
rect -4816 635734 -4216 635818
rect -4816 635498 -4634 635734
rect -4398 635498 -4216 635734
rect -4816 600054 -4216 635498
rect -4816 599818 -4634 600054
rect -4398 599818 -4216 600054
rect -4816 599734 -4216 599818
rect -4816 599498 -4634 599734
rect -4398 599498 -4216 599734
rect -4816 564054 -4216 599498
rect -4816 563818 -4634 564054
rect -4398 563818 -4216 564054
rect -4816 563734 -4216 563818
rect -4816 563498 -4634 563734
rect -4398 563498 -4216 563734
rect -4816 528054 -4216 563498
rect -4816 527818 -4634 528054
rect -4398 527818 -4216 528054
rect -4816 527734 -4216 527818
rect -4816 527498 -4634 527734
rect -4398 527498 -4216 527734
rect -4816 492054 -4216 527498
rect -4816 491818 -4634 492054
rect -4398 491818 -4216 492054
rect -4816 491734 -4216 491818
rect -4816 491498 -4634 491734
rect -4398 491498 -4216 491734
rect -4816 456054 -4216 491498
rect -4816 455818 -4634 456054
rect -4398 455818 -4216 456054
rect -4816 455734 -4216 455818
rect -4816 455498 -4634 455734
rect -4398 455498 -4216 455734
rect -4816 420054 -4216 455498
rect -4816 419818 -4634 420054
rect -4398 419818 -4216 420054
rect -4816 419734 -4216 419818
rect -4816 419498 -4634 419734
rect -4398 419498 -4216 419734
rect -4816 384054 -4216 419498
rect -4816 383818 -4634 384054
rect -4398 383818 -4216 384054
rect -4816 383734 -4216 383818
rect -4816 383498 -4634 383734
rect -4398 383498 -4216 383734
rect -4816 348054 -4216 383498
rect -4816 347818 -4634 348054
rect -4398 347818 -4216 348054
rect -4816 347734 -4216 347818
rect -4816 347498 -4634 347734
rect -4398 347498 -4216 347734
rect -4816 312054 -4216 347498
rect -4816 311818 -4634 312054
rect -4398 311818 -4216 312054
rect -4816 311734 -4216 311818
rect -4816 311498 -4634 311734
rect -4398 311498 -4216 311734
rect -4816 276054 -4216 311498
rect -4816 275818 -4634 276054
rect -4398 275818 -4216 276054
rect -4816 275734 -4216 275818
rect -4816 275498 -4634 275734
rect -4398 275498 -4216 275734
rect -4816 240054 -4216 275498
rect -4816 239818 -4634 240054
rect -4398 239818 -4216 240054
rect -4816 239734 -4216 239818
rect -4816 239498 -4634 239734
rect -4398 239498 -4216 239734
rect -4816 204054 -4216 239498
rect -4816 203818 -4634 204054
rect -4398 203818 -4216 204054
rect -4816 203734 -4216 203818
rect -4816 203498 -4634 203734
rect -4398 203498 -4216 203734
rect -4816 168054 -4216 203498
rect -4816 167818 -4634 168054
rect -4398 167818 -4216 168054
rect -4816 167734 -4216 167818
rect -4816 167498 -4634 167734
rect -4398 167498 -4216 167734
rect -4816 132054 -4216 167498
rect -4816 131818 -4634 132054
rect -4398 131818 -4216 132054
rect -4816 131734 -4216 131818
rect -4816 131498 -4634 131734
rect -4398 131498 -4216 131734
rect -4816 96054 -4216 131498
rect -4816 95818 -4634 96054
rect -4398 95818 -4216 96054
rect -4816 95734 -4216 95818
rect -4816 95498 -4634 95734
rect -4398 95498 -4216 95734
rect -4816 60054 -4216 95498
rect -4816 59818 -4634 60054
rect -4398 59818 -4216 60054
rect -4816 59734 -4216 59818
rect -4816 59498 -4634 59734
rect -4398 59498 -4216 59734
rect -4816 24054 -4216 59498
rect -4816 23818 -4634 24054
rect -4398 23818 -4216 24054
rect -4816 23734 -4216 23818
rect -4816 23498 -4634 23734
rect -4398 23498 -4216 23734
rect -4816 -3166 -4216 23498
rect -3876 706718 -3276 706740
rect -3876 706482 -3694 706718
rect -3458 706482 -3276 706718
rect -3876 706398 -3276 706482
rect -3876 706162 -3694 706398
rect -3458 706162 -3276 706398
rect -3876 690054 -3276 706162
rect 4404 706718 5004 707680
rect 4404 706482 4586 706718
rect 4822 706482 5004 706718
rect 4404 706398 5004 706482
rect 4404 706162 4586 706398
rect 4822 706162 5004 706398
rect -3876 689818 -3694 690054
rect -3458 689818 -3276 690054
rect -3876 689734 -3276 689818
rect -3876 689498 -3694 689734
rect -3458 689498 -3276 689734
rect -3876 654054 -3276 689498
rect -3876 653818 -3694 654054
rect -3458 653818 -3276 654054
rect -3876 653734 -3276 653818
rect -3876 653498 -3694 653734
rect -3458 653498 -3276 653734
rect -3876 618054 -3276 653498
rect -3876 617818 -3694 618054
rect -3458 617818 -3276 618054
rect -3876 617734 -3276 617818
rect -3876 617498 -3694 617734
rect -3458 617498 -3276 617734
rect -3876 582054 -3276 617498
rect -3876 581818 -3694 582054
rect -3458 581818 -3276 582054
rect -3876 581734 -3276 581818
rect -3876 581498 -3694 581734
rect -3458 581498 -3276 581734
rect -3876 546054 -3276 581498
rect -3876 545818 -3694 546054
rect -3458 545818 -3276 546054
rect -3876 545734 -3276 545818
rect -3876 545498 -3694 545734
rect -3458 545498 -3276 545734
rect -3876 510054 -3276 545498
rect -3876 509818 -3694 510054
rect -3458 509818 -3276 510054
rect -3876 509734 -3276 509818
rect -3876 509498 -3694 509734
rect -3458 509498 -3276 509734
rect -3876 474054 -3276 509498
rect -3876 473818 -3694 474054
rect -3458 473818 -3276 474054
rect -3876 473734 -3276 473818
rect -3876 473498 -3694 473734
rect -3458 473498 -3276 473734
rect -3876 438054 -3276 473498
rect -3876 437818 -3694 438054
rect -3458 437818 -3276 438054
rect -3876 437734 -3276 437818
rect -3876 437498 -3694 437734
rect -3458 437498 -3276 437734
rect -3876 402054 -3276 437498
rect -3876 401818 -3694 402054
rect -3458 401818 -3276 402054
rect -3876 401734 -3276 401818
rect -3876 401498 -3694 401734
rect -3458 401498 -3276 401734
rect -3876 366054 -3276 401498
rect -3876 365818 -3694 366054
rect -3458 365818 -3276 366054
rect -3876 365734 -3276 365818
rect -3876 365498 -3694 365734
rect -3458 365498 -3276 365734
rect -3876 330054 -3276 365498
rect -3876 329818 -3694 330054
rect -3458 329818 -3276 330054
rect -3876 329734 -3276 329818
rect -3876 329498 -3694 329734
rect -3458 329498 -3276 329734
rect -3876 294054 -3276 329498
rect -3876 293818 -3694 294054
rect -3458 293818 -3276 294054
rect -3876 293734 -3276 293818
rect -3876 293498 -3694 293734
rect -3458 293498 -3276 293734
rect -3876 258054 -3276 293498
rect -3876 257818 -3694 258054
rect -3458 257818 -3276 258054
rect -3876 257734 -3276 257818
rect -3876 257498 -3694 257734
rect -3458 257498 -3276 257734
rect -3876 222054 -3276 257498
rect -3876 221818 -3694 222054
rect -3458 221818 -3276 222054
rect -3876 221734 -3276 221818
rect -3876 221498 -3694 221734
rect -3458 221498 -3276 221734
rect -3876 186054 -3276 221498
rect -3876 185818 -3694 186054
rect -3458 185818 -3276 186054
rect -3876 185734 -3276 185818
rect -3876 185498 -3694 185734
rect -3458 185498 -3276 185734
rect -3876 150054 -3276 185498
rect -3876 149818 -3694 150054
rect -3458 149818 -3276 150054
rect -3876 149734 -3276 149818
rect -3876 149498 -3694 149734
rect -3458 149498 -3276 149734
rect -3876 114054 -3276 149498
rect -3876 113818 -3694 114054
rect -3458 113818 -3276 114054
rect -3876 113734 -3276 113818
rect -3876 113498 -3694 113734
rect -3458 113498 -3276 113734
rect -3876 78054 -3276 113498
rect -3876 77818 -3694 78054
rect -3458 77818 -3276 78054
rect -3876 77734 -3276 77818
rect -3876 77498 -3694 77734
rect -3458 77498 -3276 77734
rect -3876 42054 -3276 77498
rect -3876 41818 -3694 42054
rect -3458 41818 -3276 42054
rect -3876 41734 -3276 41818
rect -3876 41498 -3694 41734
rect -3458 41498 -3276 41734
rect -3876 6054 -3276 41498
rect -3876 5818 -3694 6054
rect -3458 5818 -3276 6054
rect -3876 5734 -3276 5818
rect -3876 5498 -3694 5734
rect -3458 5498 -3276 5734
rect -3876 -2226 -3276 5498
rect -2936 705778 -2336 705800
rect -2936 705542 -2754 705778
rect -2518 705542 -2336 705778
rect -2936 705458 -2336 705542
rect -2936 705222 -2754 705458
rect -2518 705222 -2336 705458
rect -2936 668454 -2336 705222
rect -2936 668218 -2754 668454
rect -2518 668218 -2336 668454
rect -2936 668134 -2336 668218
rect -2936 667898 -2754 668134
rect -2518 667898 -2336 668134
rect -2936 632454 -2336 667898
rect -2936 632218 -2754 632454
rect -2518 632218 -2336 632454
rect -2936 632134 -2336 632218
rect -2936 631898 -2754 632134
rect -2518 631898 -2336 632134
rect -2936 596454 -2336 631898
rect -2936 596218 -2754 596454
rect -2518 596218 -2336 596454
rect -2936 596134 -2336 596218
rect -2936 595898 -2754 596134
rect -2518 595898 -2336 596134
rect -2936 560454 -2336 595898
rect -2936 560218 -2754 560454
rect -2518 560218 -2336 560454
rect -2936 560134 -2336 560218
rect -2936 559898 -2754 560134
rect -2518 559898 -2336 560134
rect -2936 524454 -2336 559898
rect -2936 524218 -2754 524454
rect -2518 524218 -2336 524454
rect -2936 524134 -2336 524218
rect -2936 523898 -2754 524134
rect -2518 523898 -2336 524134
rect -2936 488454 -2336 523898
rect -2936 488218 -2754 488454
rect -2518 488218 -2336 488454
rect -2936 488134 -2336 488218
rect -2936 487898 -2754 488134
rect -2518 487898 -2336 488134
rect -2936 452454 -2336 487898
rect -2936 452218 -2754 452454
rect -2518 452218 -2336 452454
rect -2936 452134 -2336 452218
rect -2936 451898 -2754 452134
rect -2518 451898 -2336 452134
rect -2936 416454 -2336 451898
rect -2936 416218 -2754 416454
rect -2518 416218 -2336 416454
rect -2936 416134 -2336 416218
rect -2936 415898 -2754 416134
rect -2518 415898 -2336 416134
rect -2936 380454 -2336 415898
rect -2936 380218 -2754 380454
rect -2518 380218 -2336 380454
rect -2936 380134 -2336 380218
rect -2936 379898 -2754 380134
rect -2518 379898 -2336 380134
rect -2936 344454 -2336 379898
rect -2936 344218 -2754 344454
rect -2518 344218 -2336 344454
rect -2936 344134 -2336 344218
rect -2936 343898 -2754 344134
rect -2518 343898 -2336 344134
rect -2936 308454 -2336 343898
rect -2936 308218 -2754 308454
rect -2518 308218 -2336 308454
rect -2936 308134 -2336 308218
rect -2936 307898 -2754 308134
rect -2518 307898 -2336 308134
rect -2936 272454 -2336 307898
rect -2936 272218 -2754 272454
rect -2518 272218 -2336 272454
rect -2936 272134 -2336 272218
rect -2936 271898 -2754 272134
rect -2518 271898 -2336 272134
rect -2936 236454 -2336 271898
rect -2936 236218 -2754 236454
rect -2518 236218 -2336 236454
rect -2936 236134 -2336 236218
rect -2936 235898 -2754 236134
rect -2518 235898 -2336 236134
rect -2936 200454 -2336 235898
rect -2936 200218 -2754 200454
rect -2518 200218 -2336 200454
rect -2936 200134 -2336 200218
rect -2936 199898 -2754 200134
rect -2518 199898 -2336 200134
rect -2936 164454 -2336 199898
rect -2936 164218 -2754 164454
rect -2518 164218 -2336 164454
rect -2936 164134 -2336 164218
rect -2936 163898 -2754 164134
rect -2518 163898 -2336 164134
rect -2936 128454 -2336 163898
rect -2936 128218 -2754 128454
rect -2518 128218 -2336 128454
rect -2936 128134 -2336 128218
rect -2936 127898 -2754 128134
rect -2518 127898 -2336 128134
rect -2936 92454 -2336 127898
rect -2936 92218 -2754 92454
rect -2518 92218 -2336 92454
rect -2936 92134 -2336 92218
rect -2936 91898 -2754 92134
rect -2518 91898 -2336 92134
rect -2936 56454 -2336 91898
rect -2936 56218 -2754 56454
rect -2518 56218 -2336 56454
rect -2936 56134 -2336 56218
rect -2936 55898 -2754 56134
rect -2518 55898 -2336 56134
rect -2936 20454 -2336 55898
rect -2936 20218 -2754 20454
rect -2518 20218 -2336 20454
rect -2936 20134 -2336 20218
rect -2936 19898 -2754 20134
rect -2518 19898 -2336 20134
rect -2936 -1286 -2336 19898
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 686454 -1396 704282
rect -1996 686218 -1814 686454
rect -1578 686218 -1396 686454
rect -1996 686134 -1396 686218
rect -1996 685898 -1814 686134
rect -1578 685898 -1396 686134
rect -1996 650454 -1396 685898
rect -1996 650218 -1814 650454
rect -1578 650218 -1396 650454
rect -1996 650134 -1396 650218
rect -1996 649898 -1814 650134
rect -1578 649898 -1396 650134
rect -1996 614454 -1396 649898
rect -1996 614218 -1814 614454
rect -1578 614218 -1396 614454
rect -1996 614134 -1396 614218
rect -1996 613898 -1814 614134
rect -1578 613898 -1396 614134
rect -1996 578454 -1396 613898
rect -1996 578218 -1814 578454
rect -1578 578218 -1396 578454
rect -1996 578134 -1396 578218
rect -1996 577898 -1814 578134
rect -1578 577898 -1396 578134
rect -1996 542454 -1396 577898
rect -1996 542218 -1814 542454
rect -1578 542218 -1396 542454
rect -1996 542134 -1396 542218
rect -1996 541898 -1814 542134
rect -1578 541898 -1396 542134
rect -1996 506454 -1396 541898
rect -1996 506218 -1814 506454
rect -1578 506218 -1396 506454
rect -1996 506134 -1396 506218
rect -1996 505898 -1814 506134
rect -1578 505898 -1396 506134
rect -1996 470454 -1396 505898
rect -1996 470218 -1814 470454
rect -1578 470218 -1396 470454
rect -1996 470134 -1396 470218
rect -1996 469898 -1814 470134
rect -1578 469898 -1396 470134
rect -1996 434454 -1396 469898
rect -1996 434218 -1814 434454
rect -1578 434218 -1396 434454
rect -1996 434134 -1396 434218
rect -1996 433898 -1814 434134
rect -1578 433898 -1396 434134
rect -1996 398454 -1396 433898
rect -1996 398218 -1814 398454
rect -1578 398218 -1396 398454
rect -1996 398134 -1396 398218
rect -1996 397898 -1814 398134
rect -1578 397898 -1396 398134
rect -1996 362454 -1396 397898
rect -1996 362218 -1814 362454
rect -1578 362218 -1396 362454
rect -1996 362134 -1396 362218
rect -1996 361898 -1814 362134
rect -1578 361898 -1396 362134
rect -1996 326454 -1396 361898
rect -1996 326218 -1814 326454
rect -1578 326218 -1396 326454
rect -1996 326134 -1396 326218
rect -1996 325898 -1814 326134
rect -1578 325898 -1396 326134
rect -1996 290454 -1396 325898
rect -1996 290218 -1814 290454
rect -1578 290218 -1396 290454
rect -1996 290134 -1396 290218
rect -1996 289898 -1814 290134
rect -1578 289898 -1396 290134
rect -1996 254454 -1396 289898
rect -1996 254218 -1814 254454
rect -1578 254218 -1396 254454
rect -1996 254134 -1396 254218
rect -1996 253898 -1814 254134
rect -1578 253898 -1396 254134
rect -1996 218454 -1396 253898
rect -1996 218218 -1814 218454
rect -1578 218218 -1396 218454
rect -1996 218134 -1396 218218
rect -1996 217898 -1814 218134
rect -1578 217898 -1396 218134
rect -1996 182454 -1396 217898
rect -1996 182218 -1814 182454
rect -1578 182218 -1396 182454
rect -1996 182134 -1396 182218
rect -1996 181898 -1814 182134
rect -1578 181898 -1396 182134
rect -1996 146454 -1396 181898
rect -1996 146218 -1814 146454
rect -1578 146218 -1396 146454
rect -1996 146134 -1396 146218
rect -1996 145898 -1814 146134
rect -1578 145898 -1396 146134
rect -1996 110454 -1396 145898
rect -1996 110218 -1814 110454
rect -1578 110218 -1396 110454
rect -1996 110134 -1396 110218
rect -1996 109898 -1814 110134
rect -1578 109898 -1396 110134
rect -1996 74454 -1396 109898
rect -1996 74218 -1814 74454
rect -1578 74218 -1396 74454
rect -1996 74134 -1396 74218
rect -1996 73898 -1814 74134
rect -1578 73898 -1396 74134
rect -1996 38454 -1396 73898
rect -1996 38218 -1814 38454
rect -1578 38218 -1396 38454
rect -1996 38134 -1396 38218
rect -1996 37898 -1814 38134
rect -1578 37898 -1396 38134
rect -1996 2454 -1396 37898
rect -1996 2218 -1814 2454
rect -1578 2218 -1396 2454
rect -1996 2134 -1396 2218
rect -1996 1898 -1814 2134
rect -1578 1898 -1396 2134
rect -1996 -346 -1396 1898
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 804 704838 1404 705800
rect 804 704602 986 704838
rect 1222 704602 1404 704838
rect 804 704518 1404 704602
rect 804 704282 986 704518
rect 1222 704282 1404 704518
rect 804 686454 1404 704282
rect 804 686218 986 686454
rect 1222 686218 1404 686454
rect 804 686134 1404 686218
rect 804 685898 986 686134
rect 1222 685898 1404 686134
rect 804 650454 1404 685898
rect 804 650218 986 650454
rect 1222 650218 1404 650454
rect 804 650134 1404 650218
rect 804 649898 986 650134
rect 1222 649898 1404 650134
rect 804 614454 1404 649898
rect 804 614218 986 614454
rect 1222 614218 1404 614454
rect 804 614134 1404 614218
rect 804 613898 986 614134
rect 1222 613898 1404 614134
rect 804 578454 1404 613898
rect 804 578218 986 578454
rect 1222 578218 1404 578454
rect 804 578134 1404 578218
rect 804 577898 986 578134
rect 1222 577898 1404 578134
rect 804 542454 1404 577898
rect 804 542218 986 542454
rect 1222 542218 1404 542454
rect 804 542134 1404 542218
rect 804 541898 986 542134
rect 1222 541898 1404 542134
rect 804 506454 1404 541898
rect 804 506218 986 506454
rect 1222 506218 1404 506454
rect 804 506134 1404 506218
rect 804 505898 986 506134
rect 1222 505898 1404 506134
rect 804 470454 1404 505898
rect 804 470218 986 470454
rect 1222 470218 1404 470454
rect 804 470134 1404 470218
rect 804 469898 986 470134
rect 1222 469898 1404 470134
rect 804 434454 1404 469898
rect 804 434218 986 434454
rect 1222 434218 1404 434454
rect 804 434134 1404 434218
rect 804 433898 986 434134
rect 1222 433898 1404 434134
rect 804 398454 1404 433898
rect 804 398218 986 398454
rect 1222 398218 1404 398454
rect 804 398134 1404 398218
rect 804 397898 986 398134
rect 1222 397898 1404 398134
rect 804 362454 1404 397898
rect 804 362218 986 362454
rect 1222 362218 1404 362454
rect 804 362134 1404 362218
rect 804 361898 986 362134
rect 1222 361898 1404 362134
rect 804 326454 1404 361898
rect 804 326218 986 326454
rect 1222 326218 1404 326454
rect 804 326134 1404 326218
rect 804 325898 986 326134
rect 1222 325898 1404 326134
rect 804 290454 1404 325898
rect 804 290218 986 290454
rect 1222 290218 1404 290454
rect 804 290134 1404 290218
rect 804 289898 986 290134
rect 1222 289898 1404 290134
rect 804 254454 1404 289898
rect 804 254218 986 254454
rect 1222 254218 1404 254454
rect 804 254134 1404 254218
rect 804 253898 986 254134
rect 1222 253898 1404 254134
rect 804 218454 1404 253898
rect 804 218218 986 218454
rect 1222 218218 1404 218454
rect 804 218134 1404 218218
rect 804 217898 986 218134
rect 1222 217898 1404 218134
rect 804 182454 1404 217898
rect 804 182218 986 182454
rect 1222 182218 1404 182454
rect 804 182134 1404 182218
rect 804 181898 986 182134
rect 1222 181898 1404 182134
rect 804 146454 1404 181898
rect 804 146218 986 146454
rect 1222 146218 1404 146454
rect 804 146134 1404 146218
rect 804 145898 986 146134
rect 1222 145898 1404 146134
rect 804 110454 1404 145898
rect 804 110218 986 110454
rect 1222 110218 1404 110454
rect 804 110134 1404 110218
rect 804 109898 986 110134
rect 1222 109898 1404 110134
rect 804 74454 1404 109898
rect 804 74218 986 74454
rect 1222 74218 1404 74454
rect 804 74134 1404 74218
rect 804 73898 986 74134
rect 1222 73898 1404 74134
rect 804 38454 1404 73898
rect 804 38218 986 38454
rect 1222 38218 1404 38454
rect 804 38134 1404 38218
rect 804 37898 986 38134
rect 1222 37898 1404 38134
rect 804 2454 1404 37898
rect 804 2218 986 2454
rect 1222 2218 1404 2454
rect 804 2134 1404 2218
rect 804 1898 986 2134
rect 1222 1898 1404 2134
rect 804 -346 1404 1898
rect 804 -582 986 -346
rect 1222 -582 1404 -346
rect 804 -666 1404 -582
rect 804 -902 986 -666
rect 1222 -902 1404 -666
rect -2936 -1522 -2754 -1286
rect -2518 -1522 -2336 -1286
rect -2936 -1606 -2336 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 -2336 -1606
rect -2936 -1864 -2336 -1842
rect 804 -1864 1404 -902
rect 4404 690054 5004 706162
rect 4404 689818 4586 690054
rect 4822 689818 5004 690054
rect 4404 689734 5004 689818
rect 4404 689498 4586 689734
rect 4822 689498 5004 689734
rect 4404 654054 5004 689498
rect 4404 653818 4586 654054
rect 4822 653818 5004 654054
rect 4404 653734 5004 653818
rect 4404 653498 4586 653734
rect 4822 653498 5004 653734
rect 4404 618054 5004 653498
rect 4404 617818 4586 618054
rect 4822 617818 5004 618054
rect 4404 617734 5004 617818
rect 4404 617498 4586 617734
rect 4822 617498 5004 617734
rect 4404 582054 5004 617498
rect 4404 581818 4586 582054
rect 4822 581818 5004 582054
rect 4404 581734 5004 581818
rect 4404 581498 4586 581734
rect 4822 581498 5004 581734
rect 4404 546054 5004 581498
rect 4404 545818 4586 546054
rect 4822 545818 5004 546054
rect 4404 545734 5004 545818
rect 4404 545498 4586 545734
rect 4822 545498 5004 545734
rect 4404 510054 5004 545498
rect 4404 509818 4586 510054
rect 4822 509818 5004 510054
rect 4404 509734 5004 509818
rect 4404 509498 4586 509734
rect 4822 509498 5004 509734
rect 4404 474054 5004 509498
rect 4404 473818 4586 474054
rect 4822 473818 5004 474054
rect 4404 473734 5004 473818
rect 4404 473498 4586 473734
rect 4822 473498 5004 473734
rect 4404 438054 5004 473498
rect 4404 437818 4586 438054
rect 4822 437818 5004 438054
rect 4404 437734 5004 437818
rect 4404 437498 4586 437734
rect 4822 437498 5004 437734
rect 4404 402054 5004 437498
rect 4404 401818 4586 402054
rect 4822 401818 5004 402054
rect 4404 401734 5004 401818
rect 4404 401498 4586 401734
rect 4822 401498 5004 401734
rect 4404 366054 5004 401498
rect 4404 365818 4586 366054
rect 4822 365818 5004 366054
rect 4404 365734 5004 365818
rect 4404 365498 4586 365734
rect 4822 365498 5004 365734
rect 4404 330054 5004 365498
rect 4404 329818 4586 330054
rect 4822 329818 5004 330054
rect 4404 329734 5004 329818
rect 4404 329498 4586 329734
rect 4822 329498 5004 329734
rect 4404 294054 5004 329498
rect 4404 293818 4586 294054
rect 4822 293818 5004 294054
rect 4404 293734 5004 293818
rect 4404 293498 4586 293734
rect 4822 293498 5004 293734
rect 4404 258054 5004 293498
rect 4404 257818 4586 258054
rect 4822 257818 5004 258054
rect 4404 257734 5004 257818
rect 4404 257498 4586 257734
rect 4822 257498 5004 257734
rect 4404 222054 5004 257498
rect 4404 221818 4586 222054
rect 4822 221818 5004 222054
rect 4404 221734 5004 221818
rect 4404 221498 4586 221734
rect 4822 221498 5004 221734
rect 4404 186054 5004 221498
rect 4404 185818 4586 186054
rect 4822 185818 5004 186054
rect 4404 185734 5004 185818
rect 4404 185498 4586 185734
rect 4822 185498 5004 185734
rect 4404 150054 5004 185498
rect 4404 149818 4586 150054
rect 4822 149818 5004 150054
rect 4404 149734 5004 149818
rect 4404 149498 4586 149734
rect 4822 149498 5004 149734
rect 4404 114054 5004 149498
rect 4404 113818 4586 114054
rect 4822 113818 5004 114054
rect 4404 113734 5004 113818
rect 4404 113498 4586 113734
rect 4822 113498 5004 113734
rect 4404 78054 5004 113498
rect 4404 77818 4586 78054
rect 4822 77818 5004 78054
rect 4404 77734 5004 77818
rect 4404 77498 4586 77734
rect 4822 77498 5004 77734
rect 4404 42054 5004 77498
rect 4404 41818 4586 42054
rect 4822 41818 5004 42054
rect 4404 41734 5004 41818
rect 4404 41498 4586 41734
rect 4822 41498 5004 41734
rect 4404 6054 5004 41498
rect 4404 5818 4586 6054
rect 4822 5818 5004 6054
rect 4404 5734 5004 5818
rect 4404 5498 4586 5734
rect 4822 5498 5004 5734
rect -3876 -2462 -3694 -2226
rect -3458 -2462 -3276 -2226
rect -3876 -2546 -3276 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 -3276 -2546
rect -3876 -2804 -3276 -2782
rect 4404 -2226 5004 5498
rect 4404 -2462 4586 -2226
rect 4822 -2462 5004 -2226
rect 4404 -2546 5004 -2462
rect 4404 -2782 4586 -2546
rect 4822 -2782 5004 -2546
rect -4816 -3402 -4634 -3166
rect -4398 -3402 -4216 -3166
rect -4816 -3486 -4216 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 -4216 -3486
rect -4816 -3744 -4216 -3722
rect 4404 -3744 5004 -2782
rect 8004 693654 8604 708042
rect 8004 693418 8186 693654
rect 8422 693418 8604 693654
rect 8004 693334 8604 693418
rect 8004 693098 8186 693334
rect 8422 693098 8604 693334
rect 8004 657654 8604 693098
rect 8004 657418 8186 657654
rect 8422 657418 8604 657654
rect 8004 657334 8604 657418
rect 8004 657098 8186 657334
rect 8422 657098 8604 657334
rect 8004 621654 8604 657098
rect 8004 621418 8186 621654
rect 8422 621418 8604 621654
rect 8004 621334 8604 621418
rect 8004 621098 8186 621334
rect 8422 621098 8604 621334
rect 8004 585654 8604 621098
rect 8004 585418 8186 585654
rect 8422 585418 8604 585654
rect 8004 585334 8604 585418
rect 8004 585098 8186 585334
rect 8422 585098 8604 585334
rect 8004 549654 8604 585098
rect 8004 549418 8186 549654
rect 8422 549418 8604 549654
rect 8004 549334 8604 549418
rect 8004 549098 8186 549334
rect 8422 549098 8604 549334
rect 8004 513654 8604 549098
rect 8004 513418 8186 513654
rect 8422 513418 8604 513654
rect 8004 513334 8604 513418
rect 8004 513098 8186 513334
rect 8422 513098 8604 513334
rect 8004 477654 8604 513098
rect 8004 477418 8186 477654
rect 8422 477418 8604 477654
rect 8004 477334 8604 477418
rect 8004 477098 8186 477334
rect 8422 477098 8604 477334
rect 8004 441654 8604 477098
rect 8004 441418 8186 441654
rect 8422 441418 8604 441654
rect 8004 441334 8604 441418
rect 8004 441098 8186 441334
rect 8422 441098 8604 441334
rect 8004 405654 8604 441098
rect 8004 405418 8186 405654
rect 8422 405418 8604 405654
rect 8004 405334 8604 405418
rect 8004 405098 8186 405334
rect 8422 405098 8604 405334
rect 8004 369654 8604 405098
rect 8004 369418 8186 369654
rect 8422 369418 8604 369654
rect 8004 369334 8604 369418
rect 8004 369098 8186 369334
rect 8422 369098 8604 369334
rect 8004 333654 8604 369098
rect 8004 333418 8186 333654
rect 8422 333418 8604 333654
rect 8004 333334 8604 333418
rect 8004 333098 8186 333334
rect 8422 333098 8604 333334
rect 8004 297654 8604 333098
rect 8004 297418 8186 297654
rect 8422 297418 8604 297654
rect 8004 297334 8604 297418
rect 8004 297098 8186 297334
rect 8422 297098 8604 297334
rect 8004 261654 8604 297098
rect 8004 261418 8186 261654
rect 8422 261418 8604 261654
rect 8004 261334 8604 261418
rect 8004 261098 8186 261334
rect 8422 261098 8604 261334
rect 8004 225654 8604 261098
rect 8004 225418 8186 225654
rect 8422 225418 8604 225654
rect 8004 225334 8604 225418
rect 8004 225098 8186 225334
rect 8422 225098 8604 225334
rect 8004 189654 8604 225098
rect 8004 189418 8186 189654
rect 8422 189418 8604 189654
rect 8004 189334 8604 189418
rect 8004 189098 8186 189334
rect 8422 189098 8604 189334
rect 8004 153654 8604 189098
rect 8004 153418 8186 153654
rect 8422 153418 8604 153654
rect 8004 153334 8604 153418
rect 8004 153098 8186 153334
rect 8422 153098 8604 153334
rect 8004 117654 8604 153098
rect 8004 117418 8186 117654
rect 8422 117418 8604 117654
rect 8004 117334 8604 117418
rect 8004 117098 8186 117334
rect 8422 117098 8604 117334
rect 8004 81654 8604 117098
rect 8004 81418 8186 81654
rect 8422 81418 8604 81654
rect 8004 81334 8604 81418
rect 8004 81098 8186 81334
rect 8422 81098 8604 81334
rect 8004 45654 8604 81098
rect 8004 45418 8186 45654
rect 8422 45418 8604 45654
rect 8004 45334 8604 45418
rect 8004 45098 8186 45334
rect 8422 45098 8604 45334
rect 8004 9654 8604 45098
rect 8004 9418 8186 9654
rect 8422 9418 8604 9654
rect 8004 9334 8604 9418
rect 8004 9098 8186 9334
rect 8422 9098 8604 9334
rect -5756 -4342 -5574 -4106
rect -5338 -4342 -5156 -4106
rect -5756 -4426 -5156 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 -5156 -4426
rect -5756 -4684 -5156 -4662
rect 8004 -4106 8604 9098
rect 8004 -4342 8186 -4106
rect 8422 -4342 8604 -4106
rect 8004 -4426 8604 -4342
rect 8004 -4662 8186 -4426
rect 8422 -4662 8604 -4426
rect -6696 -5282 -6514 -5046
rect -6278 -5282 -6096 -5046
rect -6696 -5366 -6096 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 -6096 -5366
rect -6696 -5624 -6096 -5602
rect 8004 -5624 8604 -4662
rect 11604 697254 12204 709922
rect 29604 711418 30204 711440
rect 29604 711182 29786 711418
rect 30022 711182 30204 711418
rect 29604 711098 30204 711182
rect 29604 710862 29786 711098
rect 30022 710862 30204 711098
rect 26004 709538 26604 709560
rect 26004 709302 26186 709538
rect 26422 709302 26604 709538
rect 26004 709218 26604 709302
rect 26004 708982 26186 709218
rect 26422 708982 26604 709218
rect 22404 707658 23004 707680
rect 22404 707422 22586 707658
rect 22822 707422 23004 707658
rect 22404 707338 23004 707422
rect 22404 707102 22586 707338
rect 22822 707102 23004 707338
rect 11604 697018 11786 697254
rect 12022 697018 12204 697254
rect 11604 696934 12204 697018
rect 11604 696698 11786 696934
rect 12022 696698 12204 696934
rect 11604 661254 12204 696698
rect 11604 661018 11786 661254
rect 12022 661018 12204 661254
rect 11604 660934 12204 661018
rect 11604 660698 11786 660934
rect 12022 660698 12204 660934
rect 11604 625254 12204 660698
rect 11604 625018 11786 625254
rect 12022 625018 12204 625254
rect 11604 624934 12204 625018
rect 11604 624698 11786 624934
rect 12022 624698 12204 624934
rect 11604 589254 12204 624698
rect 11604 589018 11786 589254
rect 12022 589018 12204 589254
rect 11604 588934 12204 589018
rect 11604 588698 11786 588934
rect 12022 588698 12204 588934
rect 11604 553254 12204 588698
rect 11604 553018 11786 553254
rect 12022 553018 12204 553254
rect 11604 552934 12204 553018
rect 11604 552698 11786 552934
rect 12022 552698 12204 552934
rect 11604 517254 12204 552698
rect 11604 517018 11786 517254
rect 12022 517018 12204 517254
rect 11604 516934 12204 517018
rect 11604 516698 11786 516934
rect 12022 516698 12204 516934
rect 11604 481254 12204 516698
rect 11604 481018 11786 481254
rect 12022 481018 12204 481254
rect 11604 480934 12204 481018
rect 11604 480698 11786 480934
rect 12022 480698 12204 480934
rect 11604 445254 12204 480698
rect 11604 445018 11786 445254
rect 12022 445018 12204 445254
rect 11604 444934 12204 445018
rect 11604 444698 11786 444934
rect 12022 444698 12204 444934
rect 11604 409254 12204 444698
rect 11604 409018 11786 409254
rect 12022 409018 12204 409254
rect 11604 408934 12204 409018
rect 11604 408698 11786 408934
rect 12022 408698 12204 408934
rect 11604 373254 12204 408698
rect 11604 373018 11786 373254
rect 12022 373018 12204 373254
rect 11604 372934 12204 373018
rect 11604 372698 11786 372934
rect 12022 372698 12204 372934
rect 11604 337254 12204 372698
rect 11604 337018 11786 337254
rect 12022 337018 12204 337254
rect 11604 336934 12204 337018
rect 11604 336698 11786 336934
rect 12022 336698 12204 336934
rect 11604 301254 12204 336698
rect 11604 301018 11786 301254
rect 12022 301018 12204 301254
rect 11604 300934 12204 301018
rect 11604 300698 11786 300934
rect 12022 300698 12204 300934
rect 11604 265254 12204 300698
rect 11604 265018 11786 265254
rect 12022 265018 12204 265254
rect 11604 264934 12204 265018
rect 11604 264698 11786 264934
rect 12022 264698 12204 264934
rect 11604 229254 12204 264698
rect 11604 229018 11786 229254
rect 12022 229018 12204 229254
rect 11604 228934 12204 229018
rect 11604 228698 11786 228934
rect 12022 228698 12204 228934
rect 11604 193254 12204 228698
rect 11604 193018 11786 193254
rect 12022 193018 12204 193254
rect 11604 192934 12204 193018
rect 11604 192698 11786 192934
rect 12022 192698 12204 192934
rect 11604 157254 12204 192698
rect 11604 157018 11786 157254
rect 12022 157018 12204 157254
rect 11604 156934 12204 157018
rect 11604 156698 11786 156934
rect 12022 156698 12204 156934
rect 11604 121254 12204 156698
rect 11604 121018 11786 121254
rect 12022 121018 12204 121254
rect 11604 120934 12204 121018
rect 11604 120698 11786 120934
rect 12022 120698 12204 120934
rect 11604 85254 12204 120698
rect 11604 85018 11786 85254
rect 12022 85018 12204 85254
rect 11604 84934 12204 85018
rect 11604 84698 11786 84934
rect 12022 84698 12204 84934
rect 11604 49254 12204 84698
rect 11604 49018 11786 49254
rect 12022 49018 12204 49254
rect 11604 48934 12204 49018
rect 11604 48698 11786 48934
rect 12022 48698 12204 48934
rect 11604 13254 12204 48698
rect 11604 13018 11786 13254
rect 12022 13018 12204 13254
rect 11604 12934 12204 13018
rect 11604 12698 11786 12934
rect 12022 12698 12204 12934
rect -7636 -6222 -7454 -5986
rect -7218 -6222 -7036 -5986
rect -7636 -6306 -7036 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 -7036 -6306
rect -7636 -6564 -7036 -6542
rect 11604 -5986 12204 12698
rect 18804 705778 19404 705800
rect 18804 705542 18986 705778
rect 19222 705542 19404 705778
rect 18804 705458 19404 705542
rect 18804 705222 18986 705458
rect 19222 705222 19404 705458
rect 18804 668454 19404 705222
rect 18804 668218 18986 668454
rect 19222 668218 19404 668454
rect 18804 668134 19404 668218
rect 18804 667898 18986 668134
rect 19222 667898 19404 668134
rect 18804 632454 19404 667898
rect 18804 632218 18986 632454
rect 19222 632218 19404 632454
rect 18804 632134 19404 632218
rect 18804 631898 18986 632134
rect 19222 631898 19404 632134
rect 18804 596454 19404 631898
rect 18804 596218 18986 596454
rect 19222 596218 19404 596454
rect 18804 596134 19404 596218
rect 18804 595898 18986 596134
rect 19222 595898 19404 596134
rect 18804 560454 19404 595898
rect 18804 560218 18986 560454
rect 19222 560218 19404 560454
rect 18804 560134 19404 560218
rect 18804 559898 18986 560134
rect 19222 559898 19404 560134
rect 18804 524454 19404 559898
rect 18804 524218 18986 524454
rect 19222 524218 19404 524454
rect 18804 524134 19404 524218
rect 18804 523898 18986 524134
rect 19222 523898 19404 524134
rect 18804 488454 19404 523898
rect 18804 488218 18986 488454
rect 19222 488218 19404 488454
rect 18804 488134 19404 488218
rect 18804 487898 18986 488134
rect 19222 487898 19404 488134
rect 18804 452454 19404 487898
rect 18804 452218 18986 452454
rect 19222 452218 19404 452454
rect 18804 452134 19404 452218
rect 18804 451898 18986 452134
rect 19222 451898 19404 452134
rect 18804 416454 19404 451898
rect 18804 416218 18986 416454
rect 19222 416218 19404 416454
rect 18804 416134 19404 416218
rect 18804 415898 18986 416134
rect 19222 415898 19404 416134
rect 18804 380454 19404 415898
rect 18804 380218 18986 380454
rect 19222 380218 19404 380454
rect 18804 380134 19404 380218
rect 18804 379898 18986 380134
rect 19222 379898 19404 380134
rect 18804 344454 19404 379898
rect 18804 344218 18986 344454
rect 19222 344218 19404 344454
rect 18804 344134 19404 344218
rect 18804 343898 18986 344134
rect 19222 343898 19404 344134
rect 18804 308454 19404 343898
rect 18804 308218 18986 308454
rect 19222 308218 19404 308454
rect 18804 308134 19404 308218
rect 18804 307898 18986 308134
rect 19222 307898 19404 308134
rect 18804 272454 19404 307898
rect 18804 272218 18986 272454
rect 19222 272218 19404 272454
rect 18804 272134 19404 272218
rect 18804 271898 18986 272134
rect 19222 271898 19404 272134
rect 18804 236454 19404 271898
rect 18804 236218 18986 236454
rect 19222 236218 19404 236454
rect 18804 236134 19404 236218
rect 18804 235898 18986 236134
rect 19222 235898 19404 236134
rect 18804 200454 19404 235898
rect 18804 200218 18986 200454
rect 19222 200218 19404 200454
rect 18804 200134 19404 200218
rect 18804 199898 18986 200134
rect 19222 199898 19404 200134
rect 18804 164454 19404 199898
rect 18804 164218 18986 164454
rect 19222 164218 19404 164454
rect 18804 164134 19404 164218
rect 18804 163898 18986 164134
rect 19222 163898 19404 164134
rect 18804 128454 19404 163898
rect 18804 128218 18986 128454
rect 19222 128218 19404 128454
rect 18804 128134 19404 128218
rect 18804 127898 18986 128134
rect 19222 127898 19404 128134
rect 18804 92454 19404 127898
rect 18804 92218 18986 92454
rect 19222 92218 19404 92454
rect 18804 92134 19404 92218
rect 18804 91898 18986 92134
rect 19222 91898 19404 92134
rect 18804 56454 19404 91898
rect 18804 56218 18986 56454
rect 19222 56218 19404 56454
rect 18804 56134 19404 56218
rect 18804 55898 18986 56134
rect 19222 55898 19404 56134
rect 18804 20454 19404 55898
rect 18804 20218 18986 20454
rect 19222 20218 19404 20454
rect 18804 20134 19404 20218
rect 18804 19898 18986 20134
rect 19222 19898 19404 20134
rect 18804 -1286 19404 19898
rect 18804 -1522 18986 -1286
rect 19222 -1522 19404 -1286
rect 18804 -1606 19404 -1522
rect 18804 -1842 18986 -1606
rect 19222 -1842 19404 -1606
rect 18804 -1864 19404 -1842
rect 22404 672054 23004 707102
rect 22404 671818 22586 672054
rect 22822 671818 23004 672054
rect 22404 671734 23004 671818
rect 22404 671498 22586 671734
rect 22822 671498 23004 671734
rect 22404 636054 23004 671498
rect 22404 635818 22586 636054
rect 22822 635818 23004 636054
rect 22404 635734 23004 635818
rect 22404 635498 22586 635734
rect 22822 635498 23004 635734
rect 22404 600054 23004 635498
rect 22404 599818 22586 600054
rect 22822 599818 23004 600054
rect 22404 599734 23004 599818
rect 22404 599498 22586 599734
rect 22822 599498 23004 599734
rect 22404 564054 23004 599498
rect 22404 563818 22586 564054
rect 22822 563818 23004 564054
rect 22404 563734 23004 563818
rect 22404 563498 22586 563734
rect 22822 563498 23004 563734
rect 22404 528054 23004 563498
rect 22404 527818 22586 528054
rect 22822 527818 23004 528054
rect 22404 527734 23004 527818
rect 22404 527498 22586 527734
rect 22822 527498 23004 527734
rect 22404 492054 23004 527498
rect 22404 491818 22586 492054
rect 22822 491818 23004 492054
rect 22404 491734 23004 491818
rect 22404 491498 22586 491734
rect 22822 491498 23004 491734
rect 22404 456054 23004 491498
rect 22404 455818 22586 456054
rect 22822 455818 23004 456054
rect 22404 455734 23004 455818
rect 22404 455498 22586 455734
rect 22822 455498 23004 455734
rect 22404 420054 23004 455498
rect 22404 419818 22586 420054
rect 22822 419818 23004 420054
rect 22404 419734 23004 419818
rect 22404 419498 22586 419734
rect 22822 419498 23004 419734
rect 22404 384054 23004 419498
rect 22404 383818 22586 384054
rect 22822 383818 23004 384054
rect 22404 383734 23004 383818
rect 22404 383498 22586 383734
rect 22822 383498 23004 383734
rect 22404 348054 23004 383498
rect 22404 347818 22586 348054
rect 22822 347818 23004 348054
rect 22404 347734 23004 347818
rect 22404 347498 22586 347734
rect 22822 347498 23004 347734
rect 22404 312054 23004 347498
rect 22404 311818 22586 312054
rect 22822 311818 23004 312054
rect 22404 311734 23004 311818
rect 22404 311498 22586 311734
rect 22822 311498 23004 311734
rect 22404 276054 23004 311498
rect 22404 275818 22586 276054
rect 22822 275818 23004 276054
rect 22404 275734 23004 275818
rect 22404 275498 22586 275734
rect 22822 275498 23004 275734
rect 22404 240054 23004 275498
rect 22404 239818 22586 240054
rect 22822 239818 23004 240054
rect 22404 239734 23004 239818
rect 22404 239498 22586 239734
rect 22822 239498 23004 239734
rect 22404 204054 23004 239498
rect 22404 203818 22586 204054
rect 22822 203818 23004 204054
rect 22404 203734 23004 203818
rect 22404 203498 22586 203734
rect 22822 203498 23004 203734
rect 22404 168054 23004 203498
rect 22404 167818 22586 168054
rect 22822 167818 23004 168054
rect 22404 167734 23004 167818
rect 22404 167498 22586 167734
rect 22822 167498 23004 167734
rect 22404 132054 23004 167498
rect 22404 131818 22586 132054
rect 22822 131818 23004 132054
rect 22404 131734 23004 131818
rect 22404 131498 22586 131734
rect 22822 131498 23004 131734
rect 22404 96054 23004 131498
rect 22404 95818 22586 96054
rect 22822 95818 23004 96054
rect 22404 95734 23004 95818
rect 22404 95498 22586 95734
rect 22822 95498 23004 95734
rect 22404 60054 23004 95498
rect 22404 59818 22586 60054
rect 22822 59818 23004 60054
rect 22404 59734 23004 59818
rect 22404 59498 22586 59734
rect 22822 59498 23004 59734
rect 22404 24054 23004 59498
rect 22404 23818 22586 24054
rect 22822 23818 23004 24054
rect 22404 23734 23004 23818
rect 22404 23498 22586 23734
rect 22822 23498 23004 23734
rect 22404 -3166 23004 23498
rect 22404 -3402 22586 -3166
rect 22822 -3402 23004 -3166
rect 22404 -3486 23004 -3402
rect 22404 -3722 22586 -3486
rect 22822 -3722 23004 -3486
rect 22404 -3744 23004 -3722
rect 26004 675654 26604 708982
rect 26004 675418 26186 675654
rect 26422 675418 26604 675654
rect 26004 675334 26604 675418
rect 26004 675098 26186 675334
rect 26422 675098 26604 675334
rect 26004 639654 26604 675098
rect 26004 639418 26186 639654
rect 26422 639418 26604 639654
rect 26004 639334 26604 639418
rect 26004 639098 26186 639334
rect 26422 639098 26604 639334
rect 26004 603654 26604 639098
rect 26004 603418 26186 603654
rect 26422 603418 26604 603654
rect 26004 603334 26604 603418
rect 26004 603098 26186 603334
rect 26422 603098 26604 603334
rect 26004 567654 26604 603098
rect 26004 567418 26186 567654
rect 26422 567418 26604 567654
rect 26004 567334 26604 567418
rect 26004 567098 26186 567334
rect 26422 567098 26604 567334
rect 26004 531654 26604 567098
rect 26004 531418 26186 531654
rect 26422 531418 26604 531654
rect 26004 531334 26604 531418
rect 26004 531098 26186 531334
rect 26422 531098 26604 531334
rect 26004 495654 26604 531098
rect 26004 495418 26186 495654
rect 26422 495418 26604 495654
rect 26004 495334 26604 495418
rect 26004 495098 26186 495334
rect 26422 495098 26604 495334
rect 26004 459654 26604 495098
rect 26004 459418 26186 459654
rect 26422 459418 26604 459654
rect 26004 459334 26604 459418
rect 26004 459098 26186 459334
rect 26422 459098 26604 459334
rect 26004 423654 26604 459098
rect 26004 423418 26186 423654
rect 26422 423418 26604 423654
rect 26004 423334 26604 423418
rect 26004 423098 26186 423334
rect 26422 423098 26604 423334
rect 26004 387654 26604 423098
rect 26004 387418 26186 387654
rect 26422 387418 26604 387654
rect 26004 387334 26604 387418
rect 26004 387098 26186 387334
rect 26422 387098 26604 387334
rect 26004 351654 26604 387098
rect 26004 351418 26186 351654
rect 26422 351418 26604 351654
rect 26004 351334 26604 351418
rect 26004 351098 26186 351334
rect 26422 351098 26604 351334
rect 26004 315654 26604 351098
rect 26004 315418 26186 315654
rect 26422 315418 26604 315654
rect 26004 315334 26604 315418
rect 26004 315098 26186 315334
rect 26422 315098 26604 315334
rect 26004 279654 26604 315098
rect 26004 279418 26186 279654
rect 26422 279418 26604 279654
rect 26004 279334 26604 279418
rect 26004 279098 26186 279334
rect 26422 279098 26604 279334
rect 26004 243654 26604 279098
rect 26004 243418 26186 243654
rect 26422 243418 26604 243654
rect 26004 243334 26604 243418
rect 26004 243098 26186 243334
rect 26422 243098 26604 243334
rect 26004 207654 26604 243098
rect 26004 207418 26186 207654
rect 26422 207418 26604 207654
rect 26004 207334 26604 207418
rect 26004 207098 26186 207334
rect 26422 207098 26604 207334
rect 26004 171654 26604 207098
rect 26004 171418 26186 171654
rect 26422 171418 26604 171654
rect 26004 171334 26604 171418
rect 26004 171098 26186 171334
rect 26422 171098 26604 171334
rect 26004 135654 26604 171098
rect 26004 135418 26186 135654
rect 26422 135418 26604 135654
rect 26004 135334 26604 135418
rect 26004 135098 26186 135334
rect 26422 135098 26604 135334
rect 26004 99654 26604 135098
rect 26004 99418 26186 99654
rect 26422 99418 26604 99654
rect 26004 99334 26604 99418
rect 26004 99098 26186 99334
rect 26422 99098 26604 99334
rect 26004 63654 26604 99098
rect 26004 63418 26186 63654
rect 26422 63418 26604 63654
rect 26004 63334 26604 63418
rect 26004 63098 26186 63334
rect 26422 63098 26604 63334
rect 26004 27654 26604 63098
rect 26004 27418 26186 27654
rect 26422 27418 26604 27654
rect 26004 27334 26604 27418
rect 26004 27098 26186 27334
rect 26422 27098 26604 27334
rect 26004 -5046 26604 27098
rect 26004 -5282 26186 -5046
rect 26422 -5282 26604 -5046
rect 26004 -5366 26604 -5282
rect 26004 -5602 26186 -5366
rect 26422 -5602 26604 -5366
rect 26004 -5624 26604 -5602
rect 29604 679254 30204 710862
rect 47604 710478 48204 711440
rect 47604 710242 47786 710478
rect 48022 710242 48204 710478
rect 47604 710158 48204 710242
rect 47604 709922 47786 710158
rect 48022 709922 48204 710158
rect 44004 708598 44604 709560
rect 44004 708362 44186 708598
rect 44422 708362 44604 708598
rect 44004 708278 44604 708362
rect 44004 708042 44186 708278
rect 44422 708042 44604 708278
rect 40404 706718 41004 707680
rect 40404 706482 40586 706718
rect 40822 706482 41004 706718
rect 40404 706398 41004 706482
rect 40404 706162 40586 706398
rect 40822 706162 41004 706398
rect 29604 679018 29786 679254
rect 30022 679018 30204 679254
rect 29604 678934 30204 679018
rect 29604 678698 29786 678934
rect 30022 678698 30204 678934
rect 29604 643254 30204 678698
rect 29604 643018 29786 643254
rect 30022 643018 30204 643254
rect 29604 642934 30204 643018
rect 29604 642698 29786 642934
rect 30022 642698 30204 642934
rect 29604 607254 30204 642698
rect 29604 607018 29786 607254
rect 30022 607018 30204 607254
rect 29604 606934 30204 607018
rect 29604 606698 29786 606934
rect 30022 606698 30204 606934
rect 29604 571254 30204 606698
rect 29604 571018 29786 571254
rect 30022 571018 30204 571254
rect 29604 570934 30204 571018
rect 29604 570698 29786 570934
rect 30022 570698 30204 570934
rect 29604 535254 30204 570698
rect 29604 535018 29786 535254
rect 30022 535018 30204 535254
rect 29604 534934 30204 535018
rect 29604 534698 29786 534934
rect 30022 534698 30204 534934
rect 29604 499254 30204 534698
rect 29604 499018 29786 499254
rect 30022 499018 30204 499254
rect 29604 498934 30204 499018
rect 29604 498698 29786 498934
rect 30022 498698 30204 498934
rect 29604 463254 30204 498698
rect 29604 463018 29786 463254
rect 30022 463018 30204 463254
rect 29604 462934 30204 463018
rect 29604 462698 29786 462934
rect 30022 462698 30204 462934
rect 29604 427254 30204 462698
rect 29604 427018 29786 427254
rect 30022 427018 30204 427254
rect 29604 426934 30204 427018
rect 29604 426698 29786 426934
rect 30022 426698 30204 426934
rect 29604 391254 30204 426698
rect 29604 391018 29786 391254
rect 30022 391018 30204 391254
rect 29604 390934 30204 391018
rect 29604 390698 29786 390934
rect 30022 390698 30204 390934
rect 29604 355254 30204 390698
rect 29604 355018 29786 355254
rect 30022 355018 30204 355254
rect 29604 354934 30204 355018
rect 29604 354698 29786 354934
rect 30022 354698 30204 354934
rect 29604 319254 30204 354698
rect 29604 319018 29786 319254
rect 30022 319018 30204 319254
rect 29604 318934 30204 319018
rect 29604 318698 29786 318934
rect 30022 318698 30204 318934
rect 29604 283254 30204 318698
rect 29604 283018 29786 283254
rect 30022 283018 30204 283254
rect 29604 282934 30204 283018
rect 29604 282698 29786 282934
rect 30022 282698 30204 282934
rect 29604 247254 30204 282698
rect 29604 247018 29786 247254
rect 30022 247018 30204 247254
rect 29604 246934 30204 247018
rect 29604 246698 29786 246934
rect 30022 246698 30204 246934
rect 29604 211254 30204 246698
rect 29604 211018 29786 211254
rect 30022 211018 30204 211254
rect 29604 210934 30204 211018
rect 29604 210698 29786 210934
rect 30022 210698 30204 210934
rect 29604 175254 30204 210698
rect 29604 175018 29786 175254
rect 30022 175018 30204 175254
rect 29604 174934 30204 175018
rect 29604 174698 29786 174934
rect 30022 174698 30204 174934
rect 29604 139254 30204 174698
rect 29604 139018 29786 139254
rect 30022 139018 30204 139254
rect 29604 138934 30204 139018
rect 29604 138698 29786 138934
rect 30022 138698 30204 138934
rect 29604 103254 30204 138698
rect 29604 103018 29786 103254
rect 30022 103018 30204 103254
rect 29604 102934 30204 103018
rect 29604 102698 29786 102934
rect 30022 102698 30204 102934
rect 29604 67254 30204 102698
rect 29604 67018 29786 67254
rect 30022 67018 30204 67254
rect 29604 66934 30204 67018
rect 29604 66698 29786 66934
rect 30022 66698 30204 66934
rect 29604 31254 30204 66698
rect 29604 31018 29786 31254
rect 30022 31018 30204 31254
rect 29604 30934 30204 31018
rect 29604 30698 29786 30934
rect 30022 30698 30204 30934
rect 11604 -6222 11786 -5986
rect 12022 -6222 12204 -5986
rect 11604 -6306 12204 -6222
rect 11604 -6542 11786 -6306
rect 12022 -6542 12204 -6306
rect -8576 -7162 -8394 -6926
rect -8158 -7162 -7976 -6926
rect -8576 -7246 -7976 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 -7976 -7246
rect -8576 -7504 -7976 -7482
rect 11604 -7504 12204 -6542
rect 29604 -6926 30204 30698
rect 36804 704838 37404 705800
rect 36804 704602 36986 704838
rect 37222 704602 37404 704838
rect 36804 704518 37404 704602
rect 36804 704282 36986 704518
rect 37222 704282 37404 704518
rect 36804 686454 37404 704282
rect 36804 686218 36986 686454
rect 37222 686218 37404 686454
rect 36804 686134 37404 686218
rect 36804 685898 36986 686134
rect 37222 685898 37404 686134
rect 36804 650454 37404 685898
rect 36804 650218 36986 650454
rect 37222 650218 37404 650454
rect 36804 650134 37404 650218
rect 36804 649898 36986 650134
rect 37222 649898 37404 650134
rect 36804 614454 37404 649898
rect 36804 614218 36986 614454
rect 37222 614218 37404 614454
rect 36804 614134 37404 614218
rect 36804 613898 36986 614134
rect 37222 613898 37404 614134
rect 36804 578454 37404 613898
rect 36804 578218 36986 578454
rect 37222 578218 37404 578454
rect 36804 578134 37404 578218
rect 36804 577898 36986 578134
rect 37222 577898 37404 578134
rect 36804 542454 37404 577898
rect 36804 542218 36986 542454
rect 37222 542218 37404 542454
rect 36804 542134 37404 542218
rect 36804 541898 36986 542134
rect 37222 541898 37404 542134
rect 36804 506454 37404 541898
rect 36804 506218 36986 506454
rect 37222 506218 37404 506454
rect 36804 506134 37404 506218
rect 36804 505898 36986 506134
rect 37222 505898 37404 506134
rect 36804 470454 37404 505898
rect 36804 470218 36986 470454
rect 37222 470218 37404 470454
rect 36804 470134 37404 470218
rect 36804 469898 36986 470134
rect 37222 469898 37404 470134
rect 36804 434454 37404 469898
rect 36804 434218 36986 434454
rect 37222 434218 37404 434454
rect 36804 434134 37404 434218
rect 36804 433898 36986 434134
rect 37222 433898 37404 434134
rect 36804 398454 37404 433898
rect 36804 398218 36986 398454
rect 37222 398218 37404 398454
rect 36804 398134 37404 398218
rect 36804 397898 36986 398134
rect 37222 397898 37404 398134
rect 36804 362454 37404 397898
rect 36804 362218 36986 362454
rect 37222 362218 37404 362454
rect 36804 362134 37404 362218
rect 36804 361898 36986 362134
rect 37222 361898 37404 362134
rect 36804 326454 37404 361898
rect 36804 326218 36986 326454
rect 37222 326218 37404 326454
rect 36804 326134 37404 326218
rect 36804 325898 36986 326134
rect 37222 325898 37404 326134
rect 36804 290454 37404 325898
rect 36804 290218 36986 290454
rect 37222 290218 37404 290454
rect 36804 290134 37404 290218
rect 36804 289898 36986 290134
rect 37222 289898 37404 290134
rect 36804 254454 37404 289898
rect 36804 254218 36986 254454
rect 37222 254218 37404 254454
rect 36804 254134 37404 254218
rect 36804 253898 36986 254134
rect 37222 253898 37404 254134
rect 36804 218454 37404 253898
rect 36804 218218 36986 218454
rect 37222 218218 37404 218454
rect 36804 218134 37404 218218
rect 36804 217898 36986 218134
rect 37222 217898 37404 218134
rect 36804 182454 37404 217898
rect 36804 182218 36986 182454
rect 37222 182218 37404 182454
rect 36804 182134 37404 182218
rect 36804 181898 36986 182134
rect 37222 181898 37404 182134
rect 36804 146454 37404 181898
rect 36804 146218 36986 146454
rect 37222 146218 37404 146454
rect 36804 146134 37404 146218
rect 36804 145898 36986 146134
rect 37222 145898 37404 146134
rect 36804 110454 37404 145898
rect 36804 110218 36986 110454
rect 37222 110218 37404 110454
rect 36804 110134 37404 110218
rect 36804 109898 36986 110134
rect 37222 109898 37404 110134
rect 36804 74454 37404 109898
rect 36804 74218 36986 74454
rect 37222 74218 37404 74454
rect 36804 74134 37404 74218
rect 36804 73898 36986 74134
rect 37222 73898 37404 74134
rect 36804 38454 37404 73898
rect 36804 38218 36986 38454
rect 37222 38218 37404 38454
rect 36804 38134 37404 38218
rect 36804 37898 36986 38134
rect 37222 37898 37404 38134
rect 36804 2454 37404 37898
rect 36804 2218 36986 2454
rect 37222 2218 37404 2454
rect 36804 2134 37404 2218
rect 36804 1898 36986 2134
rect 37222 1898 37404 2134
rect 36804 -346 37404 1898
rect 36804 -582 36986 -346
rect 37222 -582 37404 -346
rect 36804 -666 37404 -582
rect 36804 -902 36986 -666
rect 37222 -902 37404 -666
rect 36804 -1864 37404 -902
rect 40404 690054 41004 706162
rect 40404 689818 40586 690054
rect 40822 689818 41004 690054
rect 40404 689734 41004 689818
rect 40404 689498 40586 689734
rect 40822 689498 41004 689734
rect 40404 654054 41004 689498
rect 40404 653818 40586 654054
rect 40822 653818 41004 654054
rect 40404 653734 41004 653818
rect 40404 653498 40586 653734
rect 40822 653498 41004 653734
rect 40404 618054 41004 653498
rect 40404 617818 40586 618054
rect 40822 617818 41004 618054
rect 40404 617734 41004 617818
rect 40404 617498 40586 617734
rect 40822 617498 41004 617734
rect 40404 582054 41004 617498
rect 40404 581818 40586 582054
rect 40822 581818 41004 582054
rect 40404 581734 41004 581818
rect 40404 581498 40586 581734
rect 40822 581498 41004 581734
rect 40404 546054 41004 581498
rect 40404 545818 40586 546054
rect 40822 545818 41004 546054
rect 40404 545734 41004 545818
rect 40404 545498 40586 545734
rect 40822 545498 41004 545734
rect 40404 510054 41004 545498
rect 40404 509818 40586 510054
rect 40822 509818 41004 510054
rect 40404 509734 41004 509818
rect 40404 509498 40586 509734
rect 40822 509498 41004 509734
rect 40404 474054 41004 509498
rect 40404 473818 40586 474054
rect 40822 473818 41004 474054
rect 40404 473734 41004 473818
rect 40404 473498 40586 473734
rect 40822 473498 41004 473734
rect 40404 438054 41004 473498
rect 40404 437818 40586 438054
rect 40822 437818 41004 438054
rect 40404 437734 41004 437818
rect 40404 437498 40586 437734
rect 40822 437498 41004 437734
rect 40404 402054 41004 437498
rect 40404 401818 40586 402054
rect 40822 401818 41004 402054
rect 40404 401734 41004 401818
rect 40404 401498 40586 401734
rect 40822 401498 41004 401734
rect 40404 366054 41004 401498
rect 40404 365818 40586 366054
rect 40822 365818 41004 366054
rect 40404 365734 41004 365818
rect 40404 365498 40586 365734
rect 40822 365498 41004 365734
rect 40404 330054 41004 365498
rect 40404 329818 40586 330054
rect 40822 329818 41004 330054
rect 40404 329734 41004 329818
rect 40404 329498 40586 329734
rect 40822 329498 41004 329734
rect 40404 294054 41004 329498
rect 40404 293818 40586 294054
rect 40822 293818 41004 294054
rect 40404 293734 41004 293818
rect 40404 293498 40586 293734
rect 40822 293498 41004 293734
rect 40404 258054 41004 293498
rect 40404 257818 40586 258054
rect 40822 257818 41004 258054
rect 40404 257734 41004 257818
rect 40404 257498 40586 257734
rect 40822 257498 41004 257734
rect 40404 222054 41004 257498
rect 40404 221818 40586 222054
rect 40822 221818 41004 222054
rect 40404 221734 41004 221818
rect 40404 221498 40586 221734
rect 40822 221498 41004 221734
rect 40404 186054 41004 221498
rect 40404 185818 40586 186054
rect 40822 185818 41004 186054
rect 40404 185734 41004 185818
rect 40404 185498 40586 185734
rect 40822 185498 41004 185734
rect 40404 150054 41004 185498
rect 40404 149818 40586 150054
rect 40822 149818 41004 150054
rect 40404 149734 41004 149818
rect 40404 149498 40586 149734
rect 40822 149498 41004 149734
rect 40404 114054 41004 149498
rect 40404 113818 40586 114054
rect 40822 113818 41004 114054
rect 40404 113734 41004 113818
rect 40404 113498 40586 113734
rect 40822 113498 41004 113734
rect 40404 78054 41004 113498
rect 40404 77818 40586 78054
rect 40822 77818 41004 78054
rect 40404 77734 41004 77818
rect 40404 77498 40586 77734
rect 40822 77498 41004 77734
rect 40404 42054 41004 77498
rect 40404 41818 40586 42054
rect 40822 41818 41004 42054
rect 40404 41734 41004 41818
rect 40404 41498 40586 41734
rect 40822 41498 41004 41734
rect 40404 6054 41004 41498
rect 40404 5818 40586 6054
rect 40822 5818 41004 6054
rect 40404 5734 41004 5818
rect 40404 5498 40586 5734
rect 40822 5498 41004 5734
rect 40404 -2226 41004 5498
rect 40404 -2462 40586 -2226
rect 40822 -2462 41004 -2226
rect 40404 -2546 41004 -2462
rect 40404 -2782 40586 -2546
rect 40822 -2782 41004 -2546
rect 40404 -3744 41004 -2782
rect 44004 693654 44604 708042
rect 44004 693418 44186 693654
rect 44422 693418 44604 693654
rect 44004 693334 44604 693418
rect 44004 693098 44186 693334
rect 44422 693098 44604 693334
rect 44004 657654 44604 693098
rect 44004 657418 44186 657654
rect 44422 657418 44604 657654
rect 44004 657334 44604 657418
rect 44004 657098 44186 657334
rect 44422 657098 44604 657334
rect 44004 621654 44604 657098
rect 44004 621418 44186 621654
rect 44422 621418 44604 621654
rect 44004 621334 44604 621418
rect 44004 621098 44186 621334
rect 44422 621098 44604 621334
rect 44004 585654 44604 621098
rect 44004 585418 44186 585654
rect 44422 585418 44604 585654
rect 44004 585334 44604 585418
rect 44004 585098 44186 585334
rect 44422 585098 44604 585334
rect 44004 549654 44604 585098
rect 44004 549418 44186 549654
rect 44422 549418 44604 549654
rect 44004 549334 44604 549418
rect 44004 549098 44186 549334
rect 44422 549098 44604 549334
rect 44004 513654 44604 549098
rect 44004 513418 44186 513654
rect 44422 513418 44604 513654
rect 44004 513334 44604 513418
rect 44004 513098 44186 513334
rect 44422 513098 44604 513334
rect 44004 477654 44604 513098
rect 44004 477418 44186 477654
rect 44422 477418 44604 477654
rect 44004 477334 44604 477418
rect 44004 477098 44186 477334
rect 44422 477098 44604 477334
rect 44004 441654 44604 477098
rect 44004 441418 44186 441654
rect 44422 441418 44604 441654
rect 44004 441334 44604 441418
rect 44004 441098 44186 441334
rect 44422 441098 44604 441334
rect 44004 405654 44604 441098
rect 44004 405418 44186 405654
rect 44422 405418 44604 405654
rect 44004 405334 44604 405418
rect 44004 405098 44186 405334
rect 44422 405098 44604 405334
rect 44004 369654 44604 405098
rect 44004 369418 44186 369654
rect 44422 369418 44604 369654
rect 44004 369334 44604 369418
rect 44004 369098 44186 369334
rect 44422 369098 44604 369334
rect 44004 333654 44604 369098
rect 44004 333418 44186 333654
rect 44422 333418 44604 333654
rect 44004 333334 44604 333418
rect 44004 333098 44186 333334
rect 44422 333098 44604 333334
rect 44004 297654 44604 333098
rect 44004 297418 44186 297654
rect 44422 297418 44604 297654
rect 44004 297334 44604 297418
rect 44004 297098 44186 297334
rect 44422 297098 44604 297334
rect 44004 261654 44604 297098
rect 44004 261418 44186 261654
rect 44422 261418 44604 261654
rect 44004 261334 44604 261418
rect 44004 261098 44186 261334
rect 44422 261098 44604 261334
rect 44004 225654 44604 261098
rect 44004 225418 44186 225654
rect 44422 225418 44604 225654
rect 44004 225334 44604 225418
rect 44004 225098 44186 225334
rect 44422 225098 44604 225334
rect 44004 189654 44604 225098
rect 44004 189418 44186 189654
rect 44422 189418 44604 189654
rect 44004 189334 44604 189418
rect 44004 189098 44186 189334
rect 44422 189098 44604 189334
rect 44004 153654 44604 189098
rect 44004 153418 44186 153654
rect 44422 153418 44604 153654
rect 44004 153334 44604 153418
rect 44004 153098 44186 153334
rect 44422 153098 44604 153334
rect 44004 117654 44604 153098
rect 44004 117418 44186 117654
rect 44422 117418 44604 117654
rect 44004 117334 44604 117418
rect 44004 117098 44186 117334
rect 44422 117098 44604 117334
rect 44004 81654 44604 117098
rect 44004 81418 44186 81654
rect 44422 81418 44604 81654
rect 44004 81334 44604 81418
rect 44004 81098 44186 81334
rect 44422 81098 44604 81334
rect 44004 45654 44604 81098
rect 44004 45418 44186 45654
rect 44422 45418 44604 45654
rect 44004 45334 44604 45418
rect 44004 45098 44186 45334
rect 44422 45098 44604 45334
rect 44004 9654 44604 45098
rect 44004 9418 44186 9654
rect 44422 9418 44604 9654
rect 44004 9334 44604 9418
rect 44004 9098 44186 9334
rect 44422 9098 44604 9334
rect 44004 -4106 44604 9098
rect 44004 -4342 44186 -4106
rect 44422 -4342 44604 -4106
rect 44004 -4426 44604 -4342
rect 44004 -4662 44186 -4426
rect 44422 -4662 44604 -4426
rect 44004 -5624 44604 -4662
rect 47604 697254 48204 709922
rect 65604 711418 66204 711440
rect 65604 711182 65786 711418
rect 66022 711182 66204 711418
rect 65604 711098 66204 711182
rect 65604 710862 65786 711098
rect 66022 710862 66204 711098
rect 62004 709538 62604 709560
rect 62004 709302 62186 709538
rect 62422 709302 62604 709538
rect 62004 709218 62604 709302
rect 62004 708982 62186 709218
rect 62422 708982 62604 709218
rect 58404 707658 59004 707680
rect 58404 707422 58586 707658
rect 58822 707422 59004 707658
rect 58404 707338 59004 707422
rect 58404 707102 58586 707338
rect 58822 707102 59004 707338
rect 47604 697018 47786 697254
rect 48022 697018 48204 697254
rect 47604 696934 48204 697018
rect 47604 696698 47786 696934
rect 48022 696698 48204 696934
rect 47604 661254 48204 696698
rect 47604 661018 47786 661254
rect 48022 661018 48204 661254
rect 47604 660934 48204 661018
rect 47604 660698 47786 660934
rect 48022 660698 48204 660934
rect 47604 625254 48204 660698
rect 47604 625018 47786 625254
rect 48022 625018 48204 625254
rect 47604 624934 48204 625018
rect 47604 624698 47786 624934
rect 48022 624698 48204 624934
rect 47604 589254 48204 624698
rect 47604 589018 47786 589254
rect 48022 589018 48204 589254
rect 47604 588934 48204 589018
rect 47604 588698 47786 588934
rect 48022 588698 48204 588934
rect 47604 553254 48204 588698
rect 47604 553018 47786 553254
rect 48022 553018 48204 553254
rect 47604 552934 48204 553018
rect 47604 552698 47786 552934
rect 48022 552698 48204 552934
rect 47604 517254 48204 552698
rect 47604 517018 47786 517254
rect 48022 517018 48204 517254
rect 47604 516934 48204 517018
rect 47604 516698 47786 516934
rect 48022 516698 48204 516934
rect 47604 481254 48204 516698
rect 47604 481018 47786 481254
rect 48022 481018 48204 481254
rect 47604 480934 48204 481018
rect 47604 480698 47786 480934
rect 48022 480698 48204 480934
rect 47604 445254 48204 480698
rect 47604 445018 47786 445254
rect 48022 445018 48204 445254
rect 47604 444934 48204 445018
rect 47604 444698 47786 444934
rect 48022 444698 48204 444934
rect 47604 409254 48204 444698
rect 47604 409018 47786 409254
rect 48022 409018 48204 409254
rect 47604 408934 48204 409018
rect 47604 408698 47786 408934
rect 48022 408698 48204 408934
rect 47604 373254 48204 408698
rect 47604 373018 47786 373254
rect 48022 373018 48204 373254
rect 47604 372934 48204 373018
rect 47604 372698 47786 372934
rect 48022 372698 48204 372934
rect 47604 337254 48204 372698
rect 47604 337018 47786 337254
rect 48022 337018 48204 337254
rect 47604 336934 48204 337018
rect 47604 336698 47786 336934
rect 48022 336698 48204 336934
rect 47604 301254 48204 336698
rect 47604 301018 47786 301254
rect 48022 301018 48204 301254
rect 47604 300934 48204 301018
rect 47604 300698 47786 300934
rect 48022 300698 48204 300934
rect 47604 265254 48204 300698
rect 47604 265018 47786 265254
rect 48022 265018 48204 265254
rect 47604 264934 48204 265018
rect 47604 264698 47786 264934
rect 48022 264698 48204 264934
rect 47604 229254 48204 264698
rect 47604 229018 47786 229254
rect 48022 229018 48204 229254
rect 47604 228934 48204 229018
rect 47604 228698 47786 228934
rect 48022 228698 48204 228934
rect 47604 193254 48204 228698
rect 47604 193018 47786 193254
rect 48022 193018 48204 193254
rect 47604 192934 48204 193018
rect 47604 192698 47786 192934
rect 48022 192698 48204 192934
rect 47604 157254 48204 192698
rect 47604 157018 47786 157254
rect 48022 157018 48204 157254
rect 47604 156934 48204 157018
rect 47604 156698 47786 156934
rect 48022 156698 48204 156934
rect 47604 121254 48204 156698
rect 47604 121018 47786 121254
rect 48022 121018 48204 121254
rect 47604 120934 48204 121018
rect 47604 120698 47786 120934
rect 48022 120698 48204 120934
rect 47604 85254 48204 120698
rect 47604 85018 47786 85254
rect 48022 85018 48204 85254
rect 47604 84934 48204 85018
rect 47604 84698 47786 84934
rect 48022 84698 48204 84934
rect 47604 49254 48204 84698
rect 47604 49018 47786 49254
rect 48022 49018 48204 49254
rect 47604 48934 48204 49018
rect 47604 48698 47786 48934
rect 48022 48698 48204 48934
rect 47604 13254 48204 48698
rect 47604 13018 47786 13254
rect 48022 13018 48204 13254
rect 47604 12934 48204 13018
rect 47604 12698 47786 12934
rect 48022 12698 48204 12934
rect 29604 -7162 29786 -6926
rect 30022 -7162 30204 -6926
rect 29604 -7246 30204 -7162
rect 29604 -7482 29786 -7246
rect 30022 -7482 30204 -7246
rect 29604 -7504 30204 -7482
rect 47604 -5986 48204 12698
rect 54804 705778 55404 705800
rect 54804 705542 54986 705778
rect 55222 705542 55404 705778
rect 54804 705458 55404 705542
rect 54804 705222 54986 705458
rect 55222 705222 55404 705458
rect 54804 668454 55404 705222
rect 57835 700364 57901 700365
rect 57835 700300 57836 700364
rect 57900 700300 57901 700364
rect 57835 700299 57901 700300
rect 57651 686220 57717 686221
rect 57651 686156 57652 686220
rect 57716 686156 57717 686220
rect 57651 686155 57717 686156
rect 54804 668218 54986 668454
rect 55222 668218 55404 668454
rect 54804 668134 55404 668218
rect 54804 667898 54986 668134
rect 55222 667898 55404 668134
rect 54804 632454 55404 667898
rect 54804 632218 54986 632454
rect 55222 632218 55404 632454
rect 54804 632134 55404 632218
rect 54804 631898 54986 632134
rect 55222 631898 55404 632134
rect 54804 596454 55404 631898
rect 54804 596218 54986 596454
rect 55222 596218 55404 596454
rect 54804 596134 55404 596218
rect 54804 595898 54986 596134
rect 55222 595898 55404 596134
rect 54804 560454 55404 595898
rect 54804 560218 54986 560454
rect 55222 560218 55404 560454
rect 54804 560134 55404 560218
rect 54804 559898 54986 560134
rect 55222 559898 55404 560134
rect 54804 524454 55404 559898
rect 57467 545596 57533 545597
rect 57467 545532 57468 545596
rect 57532 545532 57533 545596
rect 57467 545531 57533 545532
rect 57283 540292 57349 540293
rect 57283 540228 57284 540292
rect 57348 540228 57349 540292
rect 57283 540227 57349 540228
rect 54804 524218 54986 524454
rect 55222 524218 55404 524454
rect 54804 524134 55404 524218
rect 54804 523898 54986 524134
rect 55222 523898 55404 524134
rect 54804 488454 55404 523898
rect 54804 488218 54986 488454
rect 55222 488218 55404 488454
rect 54804 488134 55404 488218
rect 54804 487898 54986 488134
rect 55222 487898 55404 488134
rect 54804 452454 55404 487898
rect 54804 452218 54986 452454
rect 55222 452218 55404 452454
rect 54804 452134 55404 452218
rect 54804 451898 54986 452134
rect 55222 451898 55404 452134
rect 54804 416454 55404 451898
rect 54804 416218 54986 416454
rect 55222 416218 55404 416454
rect 54804 416134 55404 416218
rect 54804 415898 54986 416134
rect 55222 415898 55404 416134
rect 54804 380454 55404 415898
rect 57286 394365 57346 540227
rect 57283 394364 57349 394365
rect 57283 394300 57284 394364
rect 57348 394300 57349 394364
rect 57283 394299 57349 394300
rect 57470 388517 57530 545531
rect 57654 405925 57714 686155
rect 57838 411773 57898 700299
rect 58404 672054 59004 707102
rect 59123 697236 59189 697237
rect 59123 697172 59124 697236
rect 59188 697172 59189 697236
rect 59123 697171 59189 697172
rect 58404 671818 58586 672054
rect 58822 671818 59004 672054
rect 58404 671734 59004 671818
rect 58404 671498 58586 671734
rect 58822 671498 59004 671734
rect 58404 654247 59004 671498
rect 58203 650860 58269 650861
rect 58203 650796 58204 650860
rect 58268 650796 58269 650860
rect 58203 650795 58269 650796
rect 57835 411772 57901 411773
rect 57835 411708 57836 411772
rect 57900 411708 57901 411772
rect 57835 411707 57901 411708
rect 57651 405924 57717 405925
rect 57651 405860 57652 405924
rect 57716 405860 57717 405924
rect 57651 405859 57717 405860
rect 58206 398173 58266 650795
rect 58404 543000 59004 557000
rect 59126 404021 59186 697171
rect 62004 675654 62604 708982
rect 62004 675418 62186 675654
rect 62422 675418 62604 675654
rect 62004 675334 62604 675418
rect 62004 675098 62186 675334
rect 62422 675098 62604 675334
rect 59307 673844 59373 673845
rect 59307 673780 59308 673844
rect 59372 673780 59373 673844
rect 59307 673779 59373 673780
rect 59123 404020 59189 404021
rect 59123 403956 59124 404020
rect 59188 403956 59189 404020
rect 59123 403955 59189 403956
rect 59310 402117 59370 673779
rect 62004 654247 62604 675098
rect 65604 679254 66204 710862
rect 83604 710478 84204 711440
rect 83604 710242 83786 710478
rect 84022 710242 84204 710478
rect 83604 710158 84204 710242
rect 83604 709922 83786 710158
rect 84022 709922 84204 710158
rect 80004 708598 80604 709560
rect 80004 708362 80186 708598
rect 80422 708362 80604 708598
rect 80004 708278 80604 708362
rect 80004 708042 80186 708278
rect 80422 708042 80604 708278
rect 76404 706718 77004 707680
rect 76404 706482 76586 706718
rect 76822 706482 77004 706718
rect 76404 706398 77004 706482
rect 76404 706162 76586 706398
rect 76822 706162 77004 706398
rect 65604 679018 65786 679254
rect 66022 679018 66204 679254
rect 65604 678934 66204 679018
rect 65604 678698 65786 678934
rect 66022 678698 66204 678934
rect 65604 654247 66204 678698
rect 72804 704838 73404 705800
rect 72804 704602 72986 704838
rect 73222 704602 73404 704838
rect 72804 704518 73404 704602
rect 72804 704282 72986 704518
rect 73222 704282 73404 704518
rect 72804 686454 73404 704282
rect 72804 686218 72986 686454
rect 73222 686218 73404 686454
rect 72804 686134 73404 686218
rect 72804 685898 72986 686134
rect 73222 685898 73404 686134
rect 72804 654247 73404 685898
rect 76404 690054 77004 706162
rect 76404 689818 76586 690054
rect 76822 689818 77004 690054
rect 76404 689734 77004 689818
rect 76404 689498 76586 689734
rect 76822 689498 77004 689734
rect 76404 654247 77004 689498
rect 80004 693654 80604 708042
rect 80004 693418 80186 693654
rect 80422 693418 80604 693654
rect 80004 693334 80604 693418
rect 80004 693098 80186 693334
rect 80422 693098 80604 693334
rect 80004 657654 80604 693098
rect 80004 657418 80186 657654
rect 80422 657418 80604 657654
rect 80004 657334 80604 657418
rect 80004 657098 80186 657334
rect 80422 657098 80604 657334
rect 80004 654247 80604 657098
rect 83604 697254 84204 709922
rect 101604 711418 102204 711440
rect 101604 711182 101786 711418
rect 102022 711182 102204 711418
rect 101604 711098 102204 711182
rect 101604 710862 101786 711098
rect 102022 710862 102204 711098
rect 98004 709538 98604 709560
rect 98004 709302 98186 709538
rect 98422 709302 98604 709538
rect 98004 709218 98604 709302
rect 98004 708982 98186 709218
rect 98422 708982 98604 709218
rect 94404 707658 95004 707680
rect 94404 707422 94586 707658
rect 94822 707422 95004 707658
rect 94404 707338 95004 707422
rect 94404 707102 94586 707338
rect 94822 707102 95004 707338
rect 83604 697018 83786 697254
rect 84022 697018 84204 697254
rect 83604 696934 84204 697018
rect 83604 696698 83786 696934
rect 84022 696698 84204 696934
rect 83604 661254 84204 696698
rect 83604 661018 83786 661254
rect 84022 661018 84204 661254
rect 83604 660934 84204 661018
rect 83604 660698 83786 660934
rect 84022 660698 84204 660934
rect 83604 654247 84204 660698
rect 90804 705778 91404 705800
rect 90804 705542 90986 705778
rect 91222 705542 91404 705778
rect 90804 705458 91404 705542
rect 90804 705222 90986 705458
rect 91222 705222 91404 705458
rect 90804 668454 91404 705222
rect 90804 668218 90986 668454
rect 91222 668218 91404 668454
rect 90804 668134 91404 668218
rect 90804 667898 90986 668134
rect 91222 667898 91404 668134
rect 90804 654247 91404 667898
rect 94404 672054 95004 707102
rect 94404 671818 94586 672054
rect 94822 671818 95004 672054
rect 94404 671734 95004 671818
rect 94404 671498 94586 671734
rect 94822 671498 95004 671734
rect 94404 654247 95004 671498
rect 98004 675654 98604 708982
rect 98004 675418 98186 675654
rect 98422 675418 98604 675654
rect 98004 675334 98604 675418
rect 98004 675098 98186 675334
rect 98422 675098 98604 675334
rect 98004 654247 98604 675098
rect 101604 679254 102204 710862
rect 119604 710478 120204 711440
rect 119604 710242 119786 710478
rect 120022 710242 120204 710478
rect 119604 710158 120204 710242
rect 119604 709922 119786 710158
rect 120022 709922 120204 710158
rect 116004 708598 116604 709560
rect 116004 708362 116186 708598
rect 116422 708362 116604 708598
rect 116004 708278 116604 708362
rect 116004 708042 116186 708278
rect 116422 708042 116604 708278
rect 112404 706718 113004 707680
rect 112404 706482 112586 706718
rect 112822 706482 113004 706718
rect 112404 706398 113004 706482
rect 112404 706162 112586 706398
rect 112822 706162 113004 706398
rect 101604 679018 101786 679254
rect 102022 679018 102204 679254
rect 101604 678934 102204 679018
rect 101604 678698 101786 678934
rect 102022 678698 102204 678934
rect 101604 654247 102204 678698
rect 108804 704838 109404 705800
rect 108804 704602 108986 704838
rect 109222 704602 109404 704838
rect 108804 704518 109404 704602
rect 108804 704282 108986 704518
rect 109222 704282 109404 704518
rect 108804 686454 109404 704282
rect 108804 686218 108986 686454
rect 109222 686218 109404 686454
rect 108804 686134 109404 686218
rect 108804 685898 108986 686134
rect 109222 685898 109404 686134
rect 108804 654247 109404 685898
rect 112404 690054 113004 706162
rect 112404 689818 112586 690054
rect 112822 689818 113004 690054
rect 112404 689734 113004 689818
rect 112404 689498 112586 689734
rect 112822 689498 113004 689734
rect 112404 654247 113004 689498
rect 116004 693654 116604 708042
rect 116004 693418 116186 693654
rect 116422 693418 116604 693654
rect 116004 693334 116604 693418
rect 116004 693098 116186 693334
rect 116422 693098 116604 693334
rect 116004 657654 116604 693098
rect 116004 657418 116186 657654
rect 116422 657418 116604 657654
rect 116004 657334 116604 657418
rect 116004 657098 116186 657334
rect 116422 657098 116604 657334
rect 116004 654247 116604 657098
rect 119604 697254 120204 709922
rect 137604 711418 138204 711440
rect 137604 711182 137786 711418
rect 138022 711182 138204 711418
rect 137604 711098 138204 711182
rect 137604 710862 137786 711098
rect 138022 710862 138204 711098
rect 134004 709538 134604 709560
rect 134004 709302 134186 709538
rect 134422 709302 134604 709538
rect 134004 709218 134604 709302
rect 134004 708982 134186 709218
rect 134422 708982 134604 709218
rect 130404 707658 131004 707680
rect 130404 707422 130586 707658
rect 130822 707422 131004 707658
rect 130404 707338 131004 707422
rect 130404 707102 130586 707338
rect 130822 707102 131004 707338
rect 119604 697018 119786 697254
rect 120022 697018 120204 697254
rect 119604 696934 120204 697018
rect 119604 696698 119786 696934
rect 120022 696698 120204 696934
rect 119604 661254 120204 696698
rect 119604 661018 119786 661254
rect 120022 661018 120204 661254
rect 119604 660934 120204 661018
rect 119604 660698 119786 660934
rect 120022 660698 120204 660934
rect 119604 654247 120204 660698
rect 126804 705778 127404 705800
rect 126804 705542 126986 705778
rect 127222 705542 127404 705778
rect 126804 705458 127404 705542
rect 126804 705222 126986 705458
rect 127222 705222 127404 705458
rect 126804 668454 127404 705222
rect 126804 668218 126986 668454
rect 127222 668218 127404 668454
rect 126804 668134 127404 668218
rect 126804 667898 126986 668134
rect 127222 667898 127404 668134
rect 126804 654247 127404 667898
rect 130404 672054 131004 707102
rect 130404 671818 130586 672054
rect 130822 671818 131004 672054
rect 130404 671734 131004 671818
rect 130404 671498 130586 671734
rect 130822 671498 131004 671734
rect 130404 654247 131004 671498
rect 134004 675654 134604 708982
rect 134004 675418 134186 675654
rect 134422 675418 134604 675654
rect 134004 675334 134604 675418
rect 134004 675098 134186 675334
rect 134422 675098 134604 675334
rect 134004 654247 134604 675098
rect 137604 679254 138204 710862
rect 155604 710478 156204 711440
rect 155604 710242 155786 710478
rect 156022 710242 156204 710478
rect 155604 710158 156204 710242
rect 155604 709922 155786 710158
rect 156022 709922 156204 710158
rect 152004 708598 152604 709560
rect 152004 708362 152186 708598
rect 152422 708362 152604 708598
rect 152004 708278 152604 708362
rect 152004 708042 152186 708278
rect 152422 708042 152604 708278
rect 148404 706718 149004 707680
rect 148404 706482 148586 706718
rect 148822 706482 149004 706718
rect 148404 706398 149004 706482
rect 148404 706162 148586 706398
rect 148822 706162 149004 706398
rect 137604 679018 137786 679254
rect 138022 679018 138204 679254
rect 137604 678934 138204 679018
rect 137604 678698 137786 678934
rect 138022 678698 138204 678934
rect 137604 654247 138204 678698
rect 144804 704838 145404 705800
rect 144804 704602 144986 704838
rect 145222 704602 145404 704838
rect 144804 704518 145404 704602
rect 144804 704282 144986 704518
rect 145222 704282 145404 704518
rect 144804 686454 145404 704282
rect 144804 686218 144986 686454
rect 145222 686218 145404 686454
rect 144804 686134 145404 686218
rect 144804 685898 144986 686134
rect 145222 685898 145404 686134
rect 129227 652900 129293 652901
rect 129227 652836 129228 652900
rect 129292 652836 129293 652900
rect 129227 652835 129293 652836
rect 133643 652900 133709 652901
rect 133643 652836 133644 652900
rect 133708 652836 133709 652900
rect 133643 652835 133709 652836
rect 129230 651130 129290 652835
rect 133646 651810 133706 652835
rect 128608 651070 129290 651130
rect 133573 651750 133706 651810
rect 133573 651100 133633 651750
rect 125547 650860 125613 650861
rect 125547 650796 125548 650860
rect 125612 650796 125613 650860
rect 125547 650795 125613 650796
rect 125550 650589 125610 650795
rect 125547 650588 125613 650589
rect 125547 650524 125548 650588
rect 125612 650524 125613 650588
rect 125547 650523 125613 650524
rect 144804 650454 145404 685898
rect 144804 650218 144986 650454
rect 145222 650218 145404 650454
rect 144804 650134 145404 650218
rect 144804 649898 144986 650134
rect 145222 649898 145404 650134
rect 136938 643254 137262 643276
rect 136938 643018 136982 643254
rect 137218 643018 137262 643254
rect 136938 642934 137262 643018
rect 136938 642698 136982 642934
rect 137218 642698 137262 642934
rect 136938 642676 137262 642698
rect 136938 639654 137262 639676
rect 136938 639418 136982 639654
rect 137218 639418 137262 639654
rect 136938 639334 137262 639418
rect 136938 639098 136982 639334
rect 137218 639098 137262 639334
rect 136938 639076 137262 639098
rect 136938 636054 137262 636076
rect 136938 635818 136982 636054
rect 137218 635818 137262 636054
rect 136938 635734 137262 635818
rect 136938 635498 136982 635734
rect 137218 635498 137262 635734
rect 136938 635476 137262 635498
rect 136938 632454 137262 632476
rect 136938 632218 136982 632454
rect 137218 632218 137262 632454
rect 136938 632134 137262 632218
rect 136938 631898 136982 632134
rect 137218 631898 137262 632134
rect 136938 631876 137262 631898
rect 136494 625254 136814 625276
rect 136494 625018 136536 625254
rect 136772 625018 136814 625254
rect 136494 624934 136814 625018
rect 136494 624698 136536 624934
rect 136772 624698 136814 624934
rect 136494 624676 136814 624698
rect 136494 621654 136814 621676
rect 136494 621418 136536 621654
rect 136772 621418 136814 621654
rect 136494 621334 136814 621418
rect 136494 621098 136536 621334
rect 136772 621098 136814 621334
rect 136494 621076 136814 621098
rect 136494 618054 136814 618076
rect 136494 617818 136536 618054
rect 136772 617818 136814 618054
rect 136494 617734 136814 617818
rect 136494 617498 136536 617734
rect 136772 617498 136814 617734
rect 136494 617476 136814 617498
rect 136494 614454 136814 614476
rect 136494 614218 136536 614454
rect 136772 614218 136814 614454
rect 136494 614134 136814 614218
rect 136494 613898 136536 614134
rect 136772 613898 136814 614134
rect 136494 613876 136814 613898
rect 144804 614454 145404 649898
rect 144804 614218 144986 614454
rect 145222 614218 145404 614454
rect 144804 614134 145404 614218
rect 144804 613898 144986 614134
rect 145222 613898 145404 614134
rect 136938 607254 137262 607276
rect 136938 607018 136982 607254
rect 137218 607018 137262 607254
rect 136938 606934 137262 607018
rect 136938 606698 136982 606934
rect 137218 606698 137262 606934
rect 136938 606676 137262 606698
rect 136938 603654 137262 603676
rect 136938 603418 136982 603654
rect 137218 603418 137262 603654
rect 136938 603334 137262 603418
rect 136938 603098 136982 603334
rect 137218 603098 137262 603334
rect 136938 603076 137262 603098
rect 136938 600054 137262 600076
rect 136938 599818 136982 600054
rect 137218 599818 137262 600054
rect 136938 599734 137262 599818
rect 136938 599498 136982 599734
rect 137218 599498 137262 599734
rect 136938 599476 137262 599498
rect 136938 596454 137262 596476
rect 136938 596218 136982 596454
rect 137218 596218 137262 596454
rect 136938 596134 137262 596218
rect 136938 595898 136982 596134
rect 137218 595898 137262 596134
rect 136938 595876 137262 595898
rect 136494 589254 136814 589276
rect 136494 589018 136536 589254
rect 136772 589018 136814 589254
rect 136494 588934 136814 589018
rect 136494 588698 136536 588934
rect 136772 588698 136814 588934
rect 136494 588676 136814 588698
rect 136494 585654 136814 585676
rect 136494 585418 136536 585654
rect 136772 585418 136814 585654
rect 136494 585334 136814 585418
rect 136494 585098 136536 585334
rect 136772 585098 136814 585334
rect 136494 585076 136814 585098
rect 136494 582054 136814 582076
rect 136494 581818 136536 582054
rect 136772 581818 136814 582054
rect 136494 581734 136814 581818
rect 136494 581498 136536 581734
rect 136772 581498 136814 581734
rect 136494 581476 136814 581498
rect 136494 578454 136814 578476
rect 136494 578218 136536 578454
rect 136772 578218 136814 578454
rect 136494 578134 136814 578218
rect 136494 577898 136536 578134
rect 136772 577898 136814 578134
rect 136494 577876 136814 577898
rect 144804 578454 145404 613898
rect 144804 578218 144986 578454
rect 145222 578218 145404 578454
rect 144804 578134 145404 578218
rect 144804 577898 144986 578134
rect 145222 577898 145404 578134
rect 136938 571254 137262 571276
rect 136938 571018 136982 571254
rect 137218 571018 137262 571254
rect 136938 570934 137262 571018
rect 136938 570698 136982 570934
rect 137218 570698 137262 570934
rect 136938 570676 137262 570698
rect 136938 567654 137262 567676
rect 136938 567418 136982 567654
rect 137218 567418 137262 567654
rect 136938 567334 137262 567418
rect 136938 567098 136982 567334
rect 137218 567098 137262 567334
rect 136938 567076 137262 567098
rect 136938 564054 137262 564076
rect 136938 563818 136982 564054
rect 137218 563818 137262 564054
rect 136938 563734 137262 563818
rect 136938 563498 136982 563734
rect 137218 563498 137262 563734
rect 136938 563476 137262 563498
rect 72374 560430 72672 560490
rect 79366 560430 79680 560490
rect 86358 560430 86688 560490
rect 95742 560430 96032 560490
rect 102734 560430 103040 560490
rect 106230 560430 106544 560490
rect 63833 560290 64338 560350
rect 66832 560290 67466 560350
rect 68000 560290 68570 560350
rect 69168 560290 69858 560350
rect 64278 558789 64338 560290
rect 67406 558925 67466 560290
rect 68510 558925 68570 560290
rect 67403 558924 67469 558925
rect 67403 558860 67404 558924
rect 67468 558860 67469 558924
rect 67403 558859 67469 558860
rect 68507 558924 68573 558925
rect 68507 558860 68508 558924
rect 68572 558860 68573 558924
rect 68507 558859 68573 558860
rect 64275 558788 64341 558789
rect 64275 558724 64276 558788
rect 64340 558724 64341 558788
rect 64275 558723 64341 558724
rect 69798 558653 69858 560290
rect 70166 560290 70336 560350
rect 71504 560290 71698 560350
rect 70166 558925 70226 560290
rect 71638 558925 71698 560290
rect 72374 558925 72434 560430
rect 72796 560290 72986 560350
rect 72926 558925 72986 560290
rect 73662 560290 73840 560350
rect 73964 560290 74274 560350
rect 73662 558925 73722 560290
rect 74214 558925 74274 560290
rect 74950 558925 75010 560350
rect 75132 560290 75746 560350
rect 70163 558924 70229 558925
rect 70163 558860 70164 558924
rect 70228 558860 70229 558924
rect 70163 558859 70229 558860
rect 71635 558924 71701 558925
rect 71635 558860 71636 558924
rect 71700 558860 71701 558924
rect 71635 558859 71701 558860
rect 72371 558924 72437 558925
rect 72371 558860 72372 558924
rect 72436 558860 72437 558924
rect 72371 558859 72437 558860
rect 72923 558924 72989 558925
rect 72923 558860 72924 558924
rect 72988 558860 72989 558924
rect 72923 558859 72989 558860
rect 73659 558924 73725 558925
rect 73659 558860 73660 558924
rect 73724 558860 73725 558924
rect 73659 558859 73725 558860
rect 74211 558924 74277 558925
rect 74211 558860 74212 558924
rect 74276 558860 74277 558924
rect 74211 558859 74277 558860
rect 74947 558924 75013 558925
rect 74947 558860 74948 558924
rect 75012 558860 75013 558924
rect 74947 558859 75013 558860
rect 69795 558652 69861 558653
rect 69795 558588 69796 558652
rect 69860 558588 69861 558652
rect 69795 558587 69861 558588
rect 75686 558245 75746 560290
rect 75870 560290 76176 560350
rect 76300 560290 76850 560350
rect 75870 558925 75930 560290
rect 76790 558925 76850 560290
rect 77314 559330 77374 560320
rect 77468 560290 78138 560350
rect 77314 559270 77402 559330
rect 77342 558925 77402 559270
rect 75867 558924 75933 558925
rect 75867 558860 75868 558924
rect 75932 558860 75933 558924
rect 75867 558859 75933 558860
rect 76787 558924 76853 558925
rect 76787 558860 76788 558924
rect 76852 558860 76853 558924
rect 76787 558859 76853 558860
rect 77339 558924 77405 558925
rect 77339 558860 77340 558924
rect 77404 558860 77405 558924
rect 77339 558859 77405 558860
rect 78078 558381 78138 560290
rect 78446 560290 78512 560350
rect 78636 560290 79242 560350
rect 78446 558925 78506 560290
rect 79182 558925 79242 560290
rect 78443 558924 78509 558925
rect 78443 558860 78444 558924
rect 78508 558860 78509 558924
rect 78443 558859 78509 558860
rect 79179 558924 79245 558925
rect 79179 558860 79180 558924
rect 79244 558860 79245 558924
rect 79179 558859 79245 558860
rect 79366 558653 79426 560430
rect 79804 560290 79978 560350
rect 79918 558925 79978 560290
rect 80654 560290 80848 560350
rect 80972 560290 81266 560350
rect 80654 558925 80714 560290
rect 81206 558925 81266 560290
rect 81942 560290 82016 560350
rect 82140 560290 82738 560350
rect 81942 558925 82002 560290
rect 82678 558925 82738 560290
rect 82862 560290 83184 560350
rect 83308 560290 83842 560350
rect 79915 558924 79981 558925
rect 79915 558860 79916 558924
rect 79980 558860 79981 558924
rect 79915 558859 79981 558860
rect 80651 558924 80717 558925
rect 80651 558860 80652 558924
rect 80716 558860 80717 558924
rect 80651 558859 80717 558860
rect 81203 558924 81269 558925
rect 81203 558860 81204 558924
rect 81268 558860 81269 558924
rect 81203 558859 81269 558860
rect 81939 558924 82005 558925
rect 81939 558860 81940 558924
rect 82004 558860 82005 558924
rect 81939 558859 82005 558860
rect 82675 558924 82741 558925
rect 82675 558860 82676 558924
rect 82740 558860 82741 558924
rect 82675 558859 82741 558860
rect 82862 558653 82922 560290
rect 83782 558925 83842 560290
rect 84150 560290 84352 560350
rect 84476 560290 85130 560350
rect 84150 558925 84210 560290
rect 85070 558925 85130 560290
rect 85438 560290 85520 560350
rect 85644 560290 86234 560350
rect 83779 558924 83845 558925
rect 83779 558860 83780 558924
rect 83844 558860 83845 558924
rect 83779 558859 83845 558860
rect 84147 558924 84213 558925
rect 84147 558860 84148 558924
rect 84212 558860 84213 558924
rect 84147 558859 84213 558860
rect 85067 558924 85133 558925
rect 85067 558860 85068 558924
rect 85132 558860 85133 558924
rect 85067 558859 85133 558860
rect 85438 558653 85498 560290
rect 86174 558653 86234 560290
rect 86358 558925 86418 560430
rect 86782 559330 86842 560320
rect 87826 560010 87886 560320
rect 87980 560290 88258 560350
rect 87826 559950 87890 560010
rect 86726 559270 86842 559330
rect 86726 558925 86786 559270
rect 87830 558925 87890 559950
rect 88198 558925 88258 560290
rect 88934 560290 89024 560350
rect 88934 558925 88994 560290
rect 89118 558925 89178 560320
rect 89854 560290 90192 560350
rect 90316 560290 91018 560350
rect 89854 558925 89914 560290
rect 90958 558925 91018 560290
rect 91142 560290 91360 560350
rect 91484 560290 92122 560350
rect 86355 558924 86421 558925
rect 86355 558860 86356 558924
rect 86420 558860 86421 558924
rect 86355 558859 86421 558860
rect 86723 558924 86789 558925
rect 86723 558860 86724 558924
rect 86788 558860 86789 558924
rect 86723 558859 86789 558860
rect 87827 558924 87893 558925
rect 87827 558860 87828 558924
rect 87892 558860 87893 558924
rect 87827 558859 87893 558860
rect 88195 558924 88261 558925
rect 88195 558860 88196 558924
rect 88260 558860 88261 558924
rect 88195 558859 88261 558860
rect 88931 558924 88997 558925
rect 88931 558860 88932 558924
rect 88996 558860 88997 558924
rect 88931 558859 88997 558860
rect 89115 558924 89181 558925
rect 89115 558860 89116 558924
rect 89180 558860 89181 558924
rect 89115 558859 89181 558860
rect 89851 558924 89917 558925
rect 89851 558860 89852 558924
rect 89916 558860 89917 558924
rect 89851 558859 89917 558860
rect 90955 558924 91021 558925
rect 90955 558860 90956 558924
rect 91020 558860 91021 558924
rect 90955 558859 91021 558860
rect 91142 558653 91202 560290
rect 79363 558652 79429 558653
rect 79363 558588 79364 558652
rect 79428 558588 79429 558652
rect 79363 558587 79429 558588
rect 82859 558652 82925 558653
rect 82859 558588 82860 558652
rect 82924 558588 82925 558652
rect 82859 558587 82925 558588
rect 85435 558652 85501 558653
rect 85435 558588 85436 558652
rect 85500 558588 85501 558652
rect 85435 558587 85501 558588
rect 86171 558652 86237 558653
rect 86171 558588 86172 558652
rect 86236 558588 86237 558652
rect 86171 558587 86237 558588
rect 91139 558652 91205 558653
rect 91139 558588 91140 558652
rect 91204 558588 91205 558652
rect 91139 558587 91205 558588
rect 92062 558381 92122 560290
rect 92498 560010 92558 560320
rect 92652 560290 93226 560350
rect 92430 559950 92558 560010
rect 92430 558925 92490 559950
rect 93166 558925 93226 560290
rect 93350 560290 93696 560350
rect 92427 558924 92493 558925
rect 92427 558860 92428 558924
rect 92492 558860 92493 558924
rect 92427 558859 92493 558860
rect 93163 558924 93229 558925
rect 93163 558860 93164 558924
rect 93228 558860 93229 558924
rect 93163 558859 93229 558860
rect 93350 558653 93410 560290
rect 93790 559330 93850 560320
rect 93718 559270 93850 559330
rect 93718 558653 93778 559270
rect 94822 558925 94882 560350
rect 94988 560290 95066 560350
rect 95006 558925 95066 560290
rect 95742 558925 95802 560430
rect 96156 560290 96538 560350
rect 96478 558925 96538 560290
rect 97030 560290 97200 560350
rect 97324 560290 97826 560350
rect 97030 558925 97090 560290
rect 97766 558925 97826 560290
rect 98134 560290 98368 560350
rect 98492 560290 99114 560350
rect 98134 558925 98194 560290
rect 99054 558925 99114 560290
rect 99506 559330 99566 560320
rect 99660 560290 100218 560350
rect 99506 559270 99666 559330
rect 99606 558925 99666 559270
rect 100158 558925 100218 560290
rect 100342 560290 100704 560350
rect 100828 560290 101506 560350
rect 94819 558924 94885 558925
rect 94819 558860 94820 558924
rect 94884 558860 94885 558924
rect 94819 558859 94885 558860
rect 95003 558924 95069 558925
rect 95003 558860 95004 558924
rect 95068 558860 95069 558924
rect 95003 558859 95069 558860
rect 95739 558924 95805 558925
rect 95739 558860 95740 558924
rect 95804 558860 95805 558924
rect 95739 558859 95805 558860
rect 96475 558924 96541 558925
rect 96475 558860 96476 558924
rect 96540 558860 96541 558924
rect 96475 558859 96541 558860
rect 97027 558924 97093 558925
rect 97027 558860 97028 558924
rect 97092 558860 97093 558924
rect 97027 558859 97093 558860
rect 97763 558924 97829 558925
rect 97763 558860 97764 558924
rect 97828 558860 97829 558924
rect 97763 558859 97829 558860
rect 98131 558924 98197 558925
rect 98131 558860 98132 558924
rect 98196 558860 98197 558924
rect 98131 558859 98197 558860
rect 99051 558924 99117 558925
rect 99051 558860 99052 558924
rect 99116 558860 99117 558924
rect 99051 558859 99117 558860
rect 99603 558924 99669 558925
rect 99603 558860 99604 558924
rect 99668 558860 99669 558924
rect 99603 558859 99669 558860
rect 100155 558924 100221 558925
rect 100155 558860 100156 558924
rect 100220 558860 100221 558924
rect 100155 558859 100221 558860
rect 100342 558653 100402 560290
rect 101446 558925 101506 560290
rect 101630 560290 101872 560350
rect 101996 560290 102058 560350
rect 101443 558924 101509 558925
rect 101443 558860 101444 558924
rect 101508 558860 101509 558924
rect 101443 558859 101509 558860
rect 93347 558652 93413 558653
rect 93347 558588 93348 558652
rect 93412 558588 93413 558652
rect 93347 558587 93413 558588
rect 93715 558652 93781 558653
rect 93715 558588 93716 558652
rect 93780 558588 93781 558652
rect 93715 558587 93781 558588
rect 100339 558652 100405 558653
rect 100339 558588 100340 558652
rect 100404 558588 100405 558652
rect 100339 558587 100405 558588
rect 101630 558381 101690 560290
rect 101998 558653 102058 560290
rect 102734 558653 102794 560430
rect 103164 560290 103346 560350
rect 103286 558925 103346 560290
rect 104022 560290 104208 560350
rect 104332 560290 104818 560350
rect 103283 558924 103349 558925
rect 103283 558860 103284 558924
rect 103348 558860 103349 558924
rect 103283 558859 103349 558860
rect 104022 558653 104082 560290
rect 104758 558925 104818 560290
rect 105310 560290 105376 560350
rect 105500 560290 106106 560350
rect 105310 558925 105370 560290
rect 106046 558925 106106 560290
rect 104755 558924 104821 558925
rect 104755 558860 104756 558924
rect 104820 558860 104821 558924
rect 104755 558859 104821 558860
rect 105307 558924 105373 558925
rect 105307 558860 105308 558924
rect 105372 558860 105373 558924
rect 105307 558859 105373 558860
rect 106043 558924 106109 558925
rect 106043 558860 106044 558924
rect 106108 558860 106109 558924
rect 106043 558859 106109 558860
rect 106230 558653 106290 560430
rect 106668 560290 107210 560350
rect 107150 558925 107210 560290
rect 107682 559330 107742 560320
rect 107836 560290 108498 560350
rect 107682 559270 107762 559330
rect 107147 558924 107213 558925
rect 107147 558860 107148 558924
rect 107212 558860 107213 558924
rect 107147 558859 107213 558860
rect 107702 558653 107762 559270
rect 108438 558925 108498 560290
rect 108622 560290 108880 560350
rect 109004 560290 109602 560350
rect 108435 558924 108501 558925
rect 108435 558860 108436 558924
rect 108500 558860 108501 558924
rect 108435 558859 108501 558860
rect 108622 558653 108682 560290
rect 109542 558925 109602 560290
rect 109539 558924 109605 558925
rect 109539 558860 109540 558924
rect 109604 558860 109605 558924
rect 109539 558859 109605 558860
rect 101995 558652 102061 558653
rect 101995 558588 101996 558652
rect 102060 558588 102061 558652
rect 101995 558587 102061 558588
rect 102731 558652 102797 558653
rect 102731 558588 102732 558652
rect 102796 558588 102797 558652
rect 102731 558587 102797 558588
rect 104019 558652 104085 558653
rect 104019 558588 104020 558652
rect 104084 558588 104085 558652
rect 104019 558587 104085 558588
rect 106227 558652 106293 558653
rect 106227 558588 106228 558652
rect 106292 558588 106293 558652
rect 106227 558587 106293 558588
rect 107699 558652 107765 558653
rect 107699 558588 107700 558652
rect 107764 558588 107765 558652
rect 107699 558587 107765 558588
rect 108619 558652 108685 558653
rect 108619 558588 108620 558652
rect 108684 558588 108685 558652
rect 108619 558587 108685 558588
rect 78075 558380 78141 558381
rect 78075 558316 78076 558380
rect 78140 558316 78141 558380
rect 78075 558315 78141 558316
rect 92059 558380 92125 558381
rect 92059 558316 92060 558380
rect 92124 558316 92125 558380
rect 92059 558315 92125 558316
rect 101627 558380 101693 558381
rect 101627 558316 101628 558380
rect 101692 558316 101693 558380
rect 101627 558315 101693 558316
rect 75683 558244 75749 558245
rect 75683 558180 75684 558244
rect 75748 558180 75749 558244
rect 75683 558179 75749 558180
rect 62004 543000 62604 557000
rect 65604 543000 66204 557000
rect 72804 543000 73404 557000
rect 76404 546054 77004 557000
rect 76404 545818 76586 546054
rect 76822 545818 77004 546054
rect 76404 545734 77004 545818
rect 76404 545498 76586 545734
rect 76822 545498 77004 545734
rect 75867 545188 75933 545189
rect 75867 545124 75868 545188
rect 75932 545124 75933 545188
rect 75867 545123 75933 545124
rect 75870 544917 75930 545123
rect 75867 544916 75933 544917
rect 75867 544852 75868 544916
rect 75932 544852 75933 544916
rect 75867 544851 75933 544852
rect 76404 543000 77004 545498
rect 80004 549654 80604 557000
rect 80004 549418 80186 549654
rect 80422 549418 80604 549654
rect 80004 549334 80604 549418
rect 80004 549098 80186 549334
rect 80422 549098 80604 549334
rect 80004 543000 80604 549098
rect 83604 553254 84204 557000
rect 83604 553018 83786 553254
rect 84022 553018 84204 553254
rect 83604 552934 84204 553018
rect 83604 552698 83786 552934
rect 84022 552698 84204 552934
rect 83604 543000 84204 552698
rect 90804 543000 91404 557000
rect 94404 543000 95004 557000
rect 98004 543000 98604 557000
rect 101604 543000 102204 557000
rect 108804 543000 109404 557000
rect 112404 546054 113004 557000
rect 112404 545818 112586 546054
rect 112822 545818 113004 546054
rect 112404 545734 113004 545818
rect 112404 545498 112586 545734
rect 112822 545498 113004 545734
rect 112404 543000 113004 545498
rect 116004 549654 116604 557000
rect 116004 549418 116186 549654
rect 116422 549418 116604 549654
rect 116004 549334 116604 549418
rect 116004 549098 116186 549334
rect 116422 549098 116604 549334
rect 116004 543000 116604 549098
rect 119604 553254 120204 557000
rect 119604 553018 119786 553254
rect 120022 553018 120204 553254
rect 119604 552934 120204 553018
rect 119604 552698 119786 552934
rect 120022 552698 120204 552934
rect 119604 543000 120204 552698
rect 126804 543000 127404 557000
rect 130404 543000 131004 557000
rect 134004 543000 134604 557000
rect 137604 543000 138204 557000
rect 144804 543000 145404 577898
rect 148404 690054 149004 706162
rect 148404 689818 148586 690054
rect 148822 689818 149004 690054
rect 148404 689734 149004 689818
rect 148404 689498 148586 689734
rect 148822 689498 149004 689734
rect 148404 654054 149004 689498
rect 148404 653818 148586 654054
rect 148822 653818 149004 654054
rect 148404 653734 149004 653818
rect 148404 653498 148586 653734
rect 148822 653498 149004 653734
rect 148404 618054 149004 653498
rect 148404 617818 148586 618054
rect 148822 617818 149004 618054
rect 148404 617734 149004 617818
rect 148404 617498 148586 617734
rect 148822 617498 149004 617734
rect 148404 582054 149004 617498
rect 148404 581818 148586 582054
rect 148822 581818 149004 582054
rect 148404 581734 149004 581818
rect 148404 581498 148586 581734
rect 148822 581498 149004 581734
rect 148404 546054 149004 581498
rect 148404 545818 148586 546054
rect 148822 545818 149004 546054
rect 148404 545734 149004 545818
rect 148404 545498 148586 545734
rect 148822 545498 149004 545734
rect 148404 543000 149004 545498
rect 152004 693654 152604 708042
rect 152004 693418 152186 693654
rect 152422 693418 152604 693654
rect 152004 693334 152604 693418
rect 152004 693098 152186 693334
rect 152422 693098 152604 693334
rect 152004 657654 152604 693098
rect 152004 657418 152186 657654
rect 152422 657418 152604 657654
rect 152004 657334 152604 657418
rect 152004 657098 152186 657334
rect 152422 657098 152604 657334
rect 152004 621654 152604 657098
rect 152004 621418 152186 621654
rect 152422 621418 152604 621654
rect 152004 621334 152604 621418
rect 152004 621098 152186 621334
rect 152422 621098 152604 621334
rect 152004 585654 152604 621098
rect 152004 585418 152186 585654
rect 152422 585418 152604 585654
rect 152004 585334 152604 585418
rect 152004 585098 152186 585334
rect 152422 585098 152604 585334
rect 152004 549654 152604 585098
rect 152004 549418 152186 549654
rect 152422 549418 152604 549654
rect 152004 549334 152604 549418
rect 152004 549098 152186 549334
rect 152422 549098 152604 549334
rect 152004 543000 152604 549098
rect 155604 697254 156204 709922
rect 173604 711418 174204 711440
rect 173604 711182 173786 711418
rect 174022 711182 174204 711418
rect 173604 711098 174204 711182
rect 173604 710862 173786 711098
rect 174022 710862 174204 711098
rect 170004 709538 170604 709560
rect 170004 709302 170186 709538
rect 170422 709302 170604 709538
rect 170004 709218 170604 709302
rect 170004 708982 170186 709218
rect 170422 708982 170604 709218
rect 166404 707658 167004 707680
rect 166404 707422 166586 707658
rect 166822 707422 167004 707658
rect 166404 707338 167004 707422
rect 166404 707102 166586 707338
rect 166822 707102 167004 707338
rect 155604 697018 155786 697254
rect 156022 697018 156204 697254
rect 155604 696934 156204 697018
rect 155604 696698 155786 696934
rect 156022 696698 156204 696934
rect 155604 661254 156204 696698
rect 155604 661018 155786 661254
rect 156022 661018 156204 661254
rect 155604 660934 156204 661018
rect 155604 660698 155786 660934
rect 156022 660698 156204 660934
rect 155604 625254 156204 660698
rect 155604 625018 155786 625254
rect 156022 625018 156204 625254
rect 155604 624934 156204 625018
rect 155604 624698 155786 624934
rect 156022 624698 156204 624934
rect 155604 589254 156204 624698
rect 155604 589018 155786 589254
rect 156022 589018 156204 589254
rect 155604 588934 156204 589018
rect 155604 588698 155786 588934
rect 156022 588698 156204 588934
rect 155604 553254 156204 588698
rect 155604 553018 155786 553254
rect 156022 553018 156204 553254
rect 155604 552934 156204 553018
rect 155604 552698 155786 552934
rect 156022 552698 156204 552934
rect 155604 543000 156204 552698
rect 162804 705778 163404 705800
rect 162804 705542 162986 705778
rect 163222 705542 163404 705778
rect 162804 705458 163404 705542
rect 162804 705222 162986 705458
rect 163222 705222 163404 705458
rect 162804 668454 163404 705222
rect 164187 686356 164253 686357
rect 164187 686292 164188 686356
rect 164252 686292 164253 686356
rect 164187 686291 164253 686292
rect 164190 685949 164250 686291
rect 164187 685948 164253 685949
rect 164187 685884 164188 685948
rect 164252 685884 164253 685948
rect 164187 685883 164253 685884
rect 162804 668218 162986 668454
rect 163222 668218 163404 668454
rect 162804 668134 163404 668218
rect 162804 667898 162986 668134
rect 163222 667898 163404 668134
rect 162804 632454 163404 667898
rect 162804 632218 162986 632454
rect 163222 632218 163404 632454
rect 162804 632134 163404 632218
rect 162804 631898 162986 632134
rect 163222 631898 163404 632134
rect 162804 596454 163404 631898
rect 162804 596218 162986 596454
rect 163222 596218 163404 596454
rect 162804 596134 163404 596218
rect 162804 595898 162986 596134
rect 163222 595898 163404 596134
rect 162804 560454 163404 595898
rect 162804 560218 162986 560454
rect 163222 560218 163404 560454
rect 162804 560134 163404 560218
rect 162804 559898 162986 560134
rect 163222 559898 163404 560134
rect 162804 543000 163404 559898
rect 166404 672054 167004 707102
rect 166404 671818 166586 672054
rect 166822 671818 167004 672054
rect 166404 671734 167004 671818
rect 166404 671498 166586 671734
rect 166822 671498 167004 671734
rect 166404 636054 167004 671498
rect 166404 635818 166586 636054
rect 166822 635818 167004 636054
rect 166404 635734 167004 635818
rect 166404 635498 166586 635734
rect 166822 635498 167004 635734
rect 166404 600054 167004 635498
rect 166404 599818 166586 600054
rect 166822 599818 167004 600054
rect 166404 599734 167004 599818
rect 166404 599498 166586 599734
rect 166822 599498 167004 599734
rect 166404 564054 167004 599498
rect 166404 563818 166586 564054
rect 166822 563818 167004 564054
rect 166404 563734 167004 563818
rect 166404 563498 166586 563734
rect 166822 563498 167004 563734
rect 166404 543000 167004 563498
rect 170004 675654 170604 708982
rect 170004 675418 170186 675654
rect 170422 675418 170604 675654
rect 170004 675334 170604 675418
rect 170004 675098 170186 675334
rect 170422 675098 170604 675334
rect 170004 639654 170604 675098
rect 170004 639418 170186 639654
rect 170422 639418 170604 639654
rect 170004 639334 170604 639418
rect 170004 639098 170186 639334
rect 170422 639098 170604 639334
rect 170004 603654 170604 639098
rect 170004 603418 170186 603654
rect 170422 603418 170604 603654
rect 170004 603334 170604 603418
rect 170004 603098 170186 603334
rect 170422 603098 170604 603334
rect 170004 567654 170604 603098
rect 170004 567418 170186 567654
rect 170422 567418 170604 567654
rect 170004 567334 170604 567418
rect 170004 567098 170186 567334
rect 170422 567098 170604 567334
rect 170004 543000 170604 567098
rect 173604 679254 174204 710862
rect 191604 710478 192204 711440
rect 191604 710242 191786 710478
rect 192022 710242 192204 710478
rect 191604 710158 192204 710242
rect 191604 709922 191786 710158
rect 192022 709922 192204 710158
rect 188004 708598 188604 709560
rect 188004 708362 188186 708598
rect 188422 708362 188604 708598
rect 188004 708278 188604 708362
rect 188004 708042 188186 708278
rect 188422 708042 188604 708278
rect 184404 706718 185004 707680
rect 184404 706482 184586 706718
rect 184822 706482 185004 706718
rect 184404 706398 185004 706482
rect 184404 706162 184586 706398
rect 184822 706162 185004 706398
rect 173604 679018 173786 679254
rect 174022 679018 174204 679254
rect 173604 678934 174204 679018
rect 173604 678698 173786 678934
rect 174022 678698 174204 678934
rect 173604 643254 174204 678698
rect 173604 643018 173786 643254
rect 174022 643018 174204 643254
rect 173604 642934 174204 643018
rect 173604 642698 173786 642934
rect 174022 642698 174204 642934
rect 173604 607254 174204 642698
rect 173604 607018 173786 607254
rect 174022 607018 174204 607254
rect 173604 606934 174204 607018
rect 173604 606698 173786 606934
rect 174022 606698 174204 606934
rect 173604 571254 174204 606698
rect 173604 571018 173786 571254
rect 174022 571018 174204 571254
rect 173604 570934 174204 571018
rect 173604 570698 173786 570934
rect 174022 570698 174204 570934
rect 173604 543000 174204 570698
rect 180804 704838 181404 705800
rect 180804 704602 180986 704838
rect 181222 704602 181404 704838
rect 180804 704518 181404 704602
rect 180804 704282 180986 704518
rect 181222 704282 181404 704518
rect 180804 686454 181404 704282
rect 184404 690054 185004 706162
rect 184404 689818 184586 690054
rect 184822 689818 185004 690054
rect 184404 689734 185004 689818
rect 184404 689498 184586 689734
rect 184822 689498 185004 689734
rect 180804 686218 180986 686454
rect 181222 686218 181404 686454
rect 183507 686492 183573 686493
rect 183507 686428 183508 686492
rect 183572 686428 183573 686492
rect 183507 686427 183573 686428
rect 183510 686221 183570 686427
rect 180804 686134 181404 686218
rect 183507 686220 183573 686221
rect 183507 686156 183508 686220
rect 183572 686156 183573 686220
rect 183507 686155 183573 686156
rect 180804 685898 180986 686134
rect 181222 685898 181404 686134
rect 180804 650454 181404 685898
rect 183507 674116 183573 674117
rect 183507 674052 183508 674116
rect 183572 674052 183573 674116
rect 183507 674051 183573 674052
rect 183510 673845 183570 674051
rect 183507 673844 183573 673845
rect 183507 673780 183508 673844
rect 183572 673780 183573 673844
rect 183507 673779 183573 673780
rect 180804 650218 180986 650454
rect 181222 650218 181404 650454
rect 180804 650134 181404 650218
rect 180804 649898 180986 650134
rect 181222 649898 181404 650134
rect 180804 614454 181404 649898
rect 180804 614218 180986 614454
rect 181222 614218 181404 614454
rect 180804 614134 181404 614218
rect 180804 613898 180986 614134
rect 181222 613898 181404 614134
rect 180804 578454 181404 613898
rect 180804 578218 180986 578454
rect 181222 578218 181404 578454
rect 180804 578134 181404 578218
rect 180804 577898 180986 578134
rect 181222 577898 181404 578134
rect 180804 543000 181404 577898
rect 184404 654054 185004 689498
rect 188004 693654 188604 708042
rect 188004 693418 188186 693654
rect 188422 693418 188604 693654
rect 188004 693334 188604 693418
rect 188004 693098 188186 693334
rect 188422 693098 188604 693334
rect 188004 657654 188604 693098
rect 188004 657418 188186 657654
rect 188422 657418 188604 657654
rect 188004 657334 188604 657418
rect 188004 657098 188186 657334
rect 188422 657098 188604 657334
rect 188004 654247 188604 657098
rect 191604 697254 192204 709922
rect 209604 711418 210204 711440
rect 209604 711182 209786 711418
rect 210022 711182 210204 711418
rect 209604 711098 210204 711182
rect 209604 710862 209786 711098
rect 210022 710862 210204 711098
rect 206004 709538 206604 709560
rect 206004 709302 206186 709538
rect 206422 709302 206604 709538
rect 206004 709218 206604 709302
rect 206004 708982 206186 709218
rect 206422 708982 206604 709218
rect 202404 707658 203004 707680
rect 202404 707422 202586 707658
rect 202822 707422 203004 707658
rect 202404 707338 203004 707422
rect 202404 707102 202586 707338
rect 202822 707102 203004 707338
rect 191604 697018 191786 697254
rect 192022 697018 192204 697254
rect 191604 696934 192204 697018
rect 191604 696698 191786 696934
rect 192022 696698 192204 696934
rect 191604 661254 192204 696698
rect 191604 661018 191786 661254
rect 192022 661018 192204 661254
rect 191604 660934 192204 661018
rect 191604 660698 191786 660934
rect 192022 660698 192204 660934
rect 191604 654247 192204 660698
rect 198804 705778 199404 705800
rect 198804 705542 198986 705778
rect 199222 705542 199404 705778
rect 198804 705458 199404 705542
rect 198804 705222 198986 705458
rect 199222 705222 199404 705458
rect 198804 668454 199404 705222
rect 198804 668218 198986 668454
rect 199222 668218 199404 668454
rect 198804 668134 199404 668218
rect 198804 667898 198986 668134
rect 199222 667898 199404 668134
rect 198804 654247 199404 667898
rect 202404 672054 203004 707102
rect 202404 671818 202586 672054
rect 202822 671818 203004 672054
rect 202404 671734 203004 671818
rect 202404 671498 202586 671734
rect 202822 671498 203004 671734
rect 202404 654247 203004 671498
rect 206004 675654 206604 708982
rect 206004 675418 206186 675654
rect 206422 675418 206604 675654
rect 206004 675334 206604 675418
rect 206004 675098 206186 675334
rect 206422 675098 206604 675334
rect 206004 654247 206604 675098
rect 209604 679254 210204 710862
rect 227604 710478 228204 711440
rect 227604 710242 227786 710478
rect 228022 710242 228204 710478
rect 227604 710158 228204 710242
rect 227604 709922 227786 710158
rect 228022 709922 228204 710158
rect 224004 708598 224604 709560
rect 224004 708362 224186 708598
rect 224422 708362 224604 708598
rect 224004 708278 224604 708362
rect 224004 708042 224186 708278
rect 224422 708042 224604 708278
rect 220404 706718 221004 707680
rect 220404 706482 220586 706718
rect 220822 706482 221004 706718
rect 220404 706398 221004 706482
rect 220404 706162 220586 706398
rect 220822 706162 221004 706398
rect 209604 679018 209786 679254
rect 210022 679018 210204 679254
rect 209604 678934 210204 679018
rect 209604 678698 209786 678934
rect 210022 678698 210204 678934
rect 209604 654247 210204 678698
rect 216804 704838 217404 705800
rect 216804 704602 216986 704838
rect 217222 704602 217404 704838
rect 216804 704518 217404 704602
rect 216804 704282 216986 704518
rect 217222 704282 217404 704518
rect 216804 686454 217404 704282
rect 216804 686218 216986 686454
rect 217222 686218 217404 686454
rect 216804 686134 217404 686218
rect 216804 685898 216986 686134
rect 217222 685898 217404 686134
rect 216804 654247 217404 685898
rect 220404 690054 221004 706162
rect 220404 689818 220586 690054
rect 220822 689818 221004 690054
rect 220404 689734 221004 689818
rect 220404 689498 220586 689734
rect 220822 689498 221004 689734
rect 220404 654247 221004 689498
rect 224004 693654 224604 708042
rect 224004 693418 224186 693654
rect 224422 693418 224604 693654
rect 224004 693334 224604 693418
rect 224004 693098 224186 693334
rect 224422 693098 224604 693334
rect 224004 657654 224604 693098
rect 224004 657418 224186 657654
rect 224422 657418 224604 657654
rect 224004 657334 224604 657418
rect 224004 657098 224186 657334
rect 224422 657098 224604 657334
rect 224004 654247 224604 657098
rect 227604 697254 228204 709922
rect 245604 711418 246204 711440
rect 245604 711182 245786 711418
rect 246022 711182 246204 711418
rect 245604 711098 246204 711182
rect 245604 710862 245786 711098
rect 246022 710862 246204 711098
rect 242004 709538 242604 709560
rect 242004 709302 242186 709538
rect 242422 709302 242604 709538
rect 242004 709218 242604 709302
rect 242004 708982 242186 709218
rect 242422 708982 242604 709218
rect 238404 707658 239004 707680
rect 238404 707422 238586 707658
rect 238822 707422 239004 707658
rect 238404 707338 239004 707422
rect 238404 707102 238586 707338
rect 238822 707102 239004 707338
rect 227604 697018 227786 697254
rect 228022 697018 228204 697254
rect 227604 696934 228204 697018
rect 227604 696698 227786 696934
rect 228022 696698 228204 696934
rect 227604 661254 228204 696698
rect 227604 661018 227786 661254
rect 228022 661018 228204 661254
rect 227604 660934 228204 661018
rect 227604 660698 227786 660934
rect 228022 660698 228204 660934
rect 227604 654247 228204 660698
rect 234804 705778 235404 705800
rect 234804 705542 234986 705778
rect 235222 705542 235404 705778
rect 234804 705458 235404 705542
rect 234804 705222 234986 705458
rect 235222 705222 235404 705458
rect 234804 668454 235404 705222
rect 234804 668218 234986 668454
rect 235222 668218 235404 668454
rect 234804 668134 235404 668218
rect 234804 667898 234986 668134
rect 235222 667898 235404 668134
rect 234804 654247 235404 667898
rect 238404 672054 239004 707102
rect 238404 671818 238586 672054
rect 238822 671818 239004 672054
rect 238404 671734 239004 671818
rect 238404 671498 238586 671734
rect 238822 671498 239004 671734
rect 238404 654247 239004 671498
rect 242004 675654 242604 708982
rect 242004 675418 242186 675654
rect 242422 675418 242604 675654
rect 242004 675334 242604 675418
rect 242004 675098 242186 675334
rect 242422 675098 242604 675334
rect 242004 654247 242604 675098
rect 245604 679254 246204 710862
rect 263604 710478 264204 711440
rect 263604 710242 263786 710478
rect 264022 710242 264204 710478
rect 263604 710158 264204 710242
rect 263604 709922 263786 710158
rect 264022 709922 264204 710158
rect 260004 708598 260604 709560
rect 260004 708362 260186 708598
rect 260422 708362 260604 708598
rect 260004 708278 260604 708362
rect 260004 708042 260186 708278
rect 260422 708042 260604 708278
rect 256404 706718 257004 707680
rect 256404 706482 256586 706718
rect 256822 706482 257004 706718
rect 256404 706398 257004 706482
rect 256404 706162 256586 706398
rect 256822 706162 257004 706398
rect 245604 679018 245786 679254
rect 246022 679018 246204 679254
rect 245604 678934 246204 679018
rect 245604 678698 245786 678934
rect 246022 678698 246204 678934
rect 245604 654247 246204 678698
rect 252804 704838 253404 705800
rect 252804 704602 252986 704838
rect 253222 704602 253404 704838
rect 252804 704518 253404 704602
rect 252804 704282 252986 704518
rect 253222 704282 253404 704518
rect 252804 686454 253404 704282
rect 252804 686218 252986 686454
rect 253222 686218 253404 686454
rect 252804 686134 253404 686218
rect 252804 685898 252986 686134
rect 253222 685898 253404 686134
rect 252804 654247 253404 685898
rect 256404 690054 257004 706162
rect 256404 689818 256586 690054
rect 256822 689818 257004 690054
rect 256404 689734 257004 689818
rect 256404 689498 256586 689734
rect 256822 689498 257004 689734
rect 256404 654247 257004 689498
rect 260004 693654 260604 708042
rect 260004 693418 260186 693654
rect 260422 693418 260604 693654
rect 260004 693334 260604 693418
rect 260004 693098 260186 693334
rect 260422 693098 260604 693334
rect 260004 657654 260604 693098
rect 260004 657418 260186 657654
rect 260422 657418 260604 657654
rect 260004 657334 260604 657418
rect 260004 657098 260186 657334
rect 260422 657098 260604 657334
rect 260004 654247 260604 657098
rect 263604 697254 264204 709922
rect 281604 711418 282204 711440
rect 281604 711182 281786 711418
rect 282022 711182 282204 711418
rect 281604 711098 282204 711182
rect 281604 710862 281786 711098
rect 282022 710862 282204 711098
rect 278004 709538 278604 709560
rect 278004 709302 278186 709538
rect 278422 709302 278604 709538
rect 278004 709218 278604 709302
rect 278004 708982 278186 709218
rect 278422 708982 278604 709218
rect 274404 707658 275004 707680
rect 274404 707422 274586 707658
rect 274822 707422 275004 707658
rect 274404 707338 275004 707422
rect 274404 707102 274586 707338
rect 274822 707102 275004 707338
rect 263604 697018 263786 697254
rect 264022 697018 264204 697254
rect 263604 696934 264204 697018
rect 263604 696698 263786 696934
rect 264022 696698 264204 696934
rect 263604 661254 264204 696698
rect 263604 661018 263786 661254
rect 264022 661018 264204 661254
rect 263604 660934 264204 661018
rect 263604 660698 263786 660934
rect 264022 660698 264204 660934
rect 263604 654247 264204 660698
rect 270804 705778 271404 705800
rect 270804 705542 270986 705778
rect 271222 705542 271404 705778
rect 270804 705458 271404 705542
rect 270804 705222 270986 705458
rect 271222 705222 271404 705458
rect 270804 668454 271404 705222
rect 270804 668218 270986 668454
rect 271222 668218 271404 668454
rect 270804 668134 271404 668218
rect 270804 667898 270986 668134
rect 271222 667898 271404 668134
rect 184404 653818 184586 654054
rect 184822 653818 185004 654054
rect 184404 653734 185004 653818
rect 184404 653498 184586 653734
rect 184822 653498 185004 653734
rect 184404 618054 185004 653498
rect 258579 652900 258645 652901
rect 258579 652836 258580 652900
rect 258644 652836 258645 652900
rect 258579 652835 258645 652836
rect 258582 651070 258642 652835
rect 263570 651676 263636 651677
rect 263570 651612 263571 651676
rect 263635 651612 263636 651676
rect 263570 651611 263636 651612
rect 263573 651100 263633 651611
rect 266938 643254 267262 643276
rect 266938 643018 266982 643254
rect 267218 643018 267262 643254
rect 266938 642934 267262 643018
rect 266938 642698 266982 642934
rect 267218 642698 267262 642934
rect 266938 642676 267262 642698
rect 266938 639654 267262 639676
rect 266938 639418 266982 639654
rect 267218 639418 267262 639654
rect 266938 639334 267262 639418
rect 266938 639098 266982 639334
rect 267218 639098 267262 639334
rect 266938 639076 267262 639098
rect 266938 636054 267262 636076
rect 266938 635818 266982 636054
rect 267218 635818 267262 636054
rect 266938 635734 267262 635818
rect 266938 635498 266982 635734
rect 267218 635498 267262 635734
rect 266938 635476 267262 635498
rect 266938 632454 267262 632476
rect 266938 632218 266982 632454
rect 267218 632218 267262 632454
rect 266938 632134 267262 632218
rect 266938 631898 266982 632134
rect 267218 631898 267262 632134
rect 266938 631876 267262 631898
rect 270804 632454 271404 667898
rect 270804 632218 270986 632454
rect 271222 632218 271404 632454
rect 270804 632134 271404 632218
rect 270804 631898 270986 632134
rect 271222 631898 271404 632134
rect 266494 625254 266814 625276
rect 266494 625018 266536 625254
rect 266772 625018 266814 625254
rect 266494 624934 266814 625018
rect 266494 624698 266536 624934
rect 266772 624698 266814 624934
rect 266494 624676 266814 624698
rect 266494 621654 266814 621676
rect 266494 621418 266536 621654
rect 266772 621418 266814 621654
rect 266494 621334 266814 621418
rect 266494 621098 266536 621334
rect 266772 621098 266814 621334
rect 266494 621076 266814 621098
rect 184404 617818 184586 618054
rect 184822 617818 185004 618054
rect 184404 617734 185004 617818
rect 184404 617498 184586 617734
rect 184822 617498 185004 617734
rect 184404 582054 185004 617498
rect 266494 618054 266814 618076
rect 266494 617818 266536 618054
rect 266772 617818 266814 618054
rect 266494 617734 266814 617818
rect 266494 617498 266536 617734
rect 266772 617498 266814 617734
rect 266494 617476 266814 617498
rect 266494 614454 266814 614476
rect 266494 614218 266536 614454
rect 266772 614218 266814 614454
rect 266494 614134 266814 614218
rect 266494 613898 266536 614134
rect 266772 613898 266814 614134
rect 266494 613876 266814 613898
rect 266938 607254 267262 607276
rect 266938 607018 266982 607254
rect 267218 607018 267262 607254
rect 266938 606934 267262 607018
rect 266938 606698 266982 606934
rect 267218 606698 267262 606934
rect 266938 606676 267262 606698
rect 266938 603654 267262 603676
rect 266938 603418 266982 603654
rect 267218 603418 267262 603654
rect 266938 603334 267262 603418
rect 266938 603098 266982 603334
rect 267218 603098 267262 603334
rect 266938 603076 267262 603098
rect 266938 600054 267262 600076
rect 266938 599818 266982 600054
rect 267218 599818 267262 600054
rect 266938 599734 267262 599818
rect 266938 599498 266982 599734
rect 267218 599498 267262 599734
rect 266938 599476 267262 599498
rect 266938 596454 267262 596476
rect 266938 596218 266982 596454
rect 267218 596218 267262 596454
rect 266938 596134 267262 596218
rect 266938 595898 266982 596134
rect 267218 595898 267262 596134
rect 266938 595876 267262 595898
rect 270804 596454 271404 631898
rect 270804 596218 270986 596454
rect 271222 596218 271404 596454
rect 270804 596134 271404 596218
rect 270804 595898 270986 596134
rect 271222 595898 271404 596134
rect 266494 589254 266814 589276
rect 266494 589018 266536 589254
rect 266772 589018 266814 589254
rect 266494 588934 266814 589018
rect 266494 588698 266536 588934
rect 266772 588698 266814 588934
rect 266494 588676 266814 588698
rect 266494 585654 266814 585676
rect 266494 585418 266536 585654
rect 266772 585418 266814 585654
rect 266494 585334 266814 585418
rect 266494 585098 266536 585334
rect 266772 585098 266814 585334
rect 266494 585076 266814 585098
rect 184404 581818 184586 582054
rect 184822 581818 185004 582054
rect 184404 581734 185004 581818
rect 184404 581498 184586 581734
rect 184822 581498 185004 581734
rect 184404 546054 185004 581498
rect 266494 582054 266814 582076
rect 266494 581818 266536 582054
rect 266772 581818 266814 582054
rect 266494 581734 266814 581818
rect 266494 581498 266536 581734
rect 266772 581498 266814 581734
rect 266494 581476 266814 581498
rect 266494 578454 266814 578476
rect 266494 578218 266536 578454
rect 266772 578218 266814 578454
rect 266494 578134 266814 578218
rect 266494 577898 266536 578134
rect 266772 577898 266814 578134
rect 266494 577876 266814 577898
rect 266938 571254 267262 571276
rect 266938 571018 266982 571254
rect 267218 571018 267262 571254
rect 266938 570934 267262 571018
rect 266938 570698 266982 570934
rect 267218 570698 267262 570934
rect 266938 570676 267262 570698
rect 266938 567654 267262 567676
rect 266938 567418 266982 567654
rect 267218 567418 267262 567654
rect 266938 567334 267262 567418
rect 266938 567098 266982 567334
rect 267218 567098 267262 567334
rect 266938 567076 267262 567098
rect 266938 564054 267262 564076
rect 266938 563818 266982 564054
rect 267218 563818 267262 564054
rect 266938 563734 267262 563818
rect 266938 563498 266982 563734
rect 267218 563498 267262 563734
rect 266938 563476 267262 563498
rect 201504 560430 201786 560490
rect 193833 560290 194426 560350
rect 194366 558789 194426 560290
rect 196206 560290 196832 560350
rect 197494 560290 198000 560350
rect 198782 560290 199168 560350
rect 200254 560290 200336 560350
rect 196206 558925 196266 560290
rect 197494 558925 197554 560290
rect 196203 558924 196269 558925
rect 196203 558860 196204 558924
rect 196268 558860 196269 558924
rect 196203 558859 196269 558860
rect 197491 558924 197557 558925
rect 197491 558860 197492 558924
rect 197556 558860 197557 558924
rect 197491 558859 197557 558860
rect 194363 558788 194429 558789
rect 194363 558724 194364 558788
rect 194428 558724 194429 558788
rect 194363 558723 194429 558724
rect 198782 557701 198842 560290
rect 200254 557837 200314 560290
rect 201726 558925 201786 560430
rect 207062 560430 207344 560490
rect 217550 560430 217856 560490
rect 221046 560430 221360 560490
rect 270804 560454 271404 595898
rect 202462 560290 202672 560350
rect 201723 558924 201789 558925
rect 201723 558860 201724 558924
rect 201788 558860 201789 558924
rect 201723 558859 201789 558860
rect 202462 558653 202522 560290
rect 202766 559330 202826 560320
rect 202646 559270 202826 559330
rect 203750 560290 203840 560350
rect 202646 558925 202706 559270
rect 202643 558924 202709 558925
rect 202643 558860 202644 558924
rect 202708 558860 202709 558924
rect 202643 558859 202709 558860
rect 203750 558789 203810 560290
rect 203934 558925 203994 560320
rect 204854 560290 205008 560350
rect 205132 560290 205466 560350
rect 203931 558924 203997 558925
rect 203931 558860 203932 558924
rect 203996 558860 203997 558924
rect 203931 558859 203997 558860
rect 203747 558788 203813 558789
rect 203747 558724 203748 558788
rect 203812 558724 203813 558788
rect 203747 558723 203813 558724
rect 204854 558653 204914 560290
rect 205406 558925 205466 560290
rect 206142 558925 206202 560350
rect 206300 560290 206938 560350
rect 205403 558924 205469 558925
rect 205403 558860 205404 558924
rect 205468 558860 205469 558924
rect 205403 558859 205469 558860
rect 206139 558924 206205 558925
rect 206139 558860 206140 558924
rect 206204 558860 206205 558924
rect 206139 558859 206205 558860
rect 202459 558652 202525 558653
rect 202459 558588 202460 558652
rect 202524 558588 202525 558652
rect 202459 558587 202525 558588
rect 204851 558652 204917 558653
rect 204851 558588 204852 558652
rect 204916 558588 204917 558652
rect 204851 558587 204917 558588
rect 200251 557836 200317 557837
rect 200251 557772 200252 557836
rect 200316 557772 200317 557836
rect 200251 557771 200317 557772
rect 198779 557700 198845 557701
rect 198779 557636 198780 557700
rect 198844 557636 198845 557700
rect 198779 557635 198845 557636
rect 206878 557565 206938 560290
rect 207062 557701 207122 560430
rect 207468 560290 208042 560350
rect 207059 557700 207125 557701
rect 207059 557636 207060 557700
rect 207124 557636 207125 557700
rect 207059 557635 207125 557636
rect 207982 557565 208042 560290
rect 208350 560290 208512 560350
rect 208636 560290 209330 560350
rect 208350 558925 208410 560290
rect 208347 558924 208413 558925
rect 208347 558860 208348 558924
rect 208412 558860 208413 558924
rect 208347 558859 208413 558860
rect 209270 557565 209330 560290
rect 209638 558653 209698 560350
rect 209804 560290 210434 560350
rect 209635 558652 209701 558653
rect 209635 558588 209636 558652
rect 209700 558588 209701 558652
rect 209635 558587 209701 558588
rect 210374 557701 210434 560290
rect 210558 560290 210848 560350
rect 210558 558925 210618 560290
rect 210942 560010 211002 560320
rect 211846 560290 212016 560350
rect 212140 560290 212458 560350
rect 211107 560012 211173 560013
rect 211107 560010 211108 560012
rect 210942 559950 211108 560010
rect 211107 559948 211108 559950
rect 211172 559948 211173 560012
rect 211107 559947 211173 559948
rect 211846 558925 211906 560290
rect 210555 558924 210621 558925
rect 210555 558860 210556 558924
rect 210620 558860 210621 558924
rect 210555 558859 210621 558860
rect 211843 558924 211909 558925
rect 211843 558860 211844 558924
rect 211908 558860 211909 558924
rect 211843 558859 211909 558860
rect 210371 557700 210437 557701
rect 210371 557636 210372 557700
rect 210436 557636 210437 557700
rect 210371 557635 210437 557636
rect 212398 557565 212458 560290
rect 213134 558925 213194 560350
rect 213308 560290 213562 560350
rect 213131 558924 213197 558925
rect 213131 558860 213132 558924
rect 213196 558860 213197 558924
rect 213131 558859 213197 558860
rect 213502 557565 213562 560290
rect 214054 560290 214352 560350
rect 214476 560290 214850 560350
rect 214054 558925 214114 560290
rect 214051 558924 214117 558925
rect 214051 558860 214052 558924
rect 214116 558860 214117 558924
rect 214051 558859 214117 558860
rect 214790 557565 214850 560290
rect 215342 560290 215520 560350
rect 215644 560290 216322 560350
rect 215342 558925 215402 560290
rect 215339 558924 215405 558925
rect 215339 558860 215340 558924
rect 215404 558860 215405 558924
rect 215339 558859 215405 558860
rect 216262 557565 216322 560290
rect 216630 558789 216690 560350
rect 216812 560290 217426 560350
rect 216627 558788 216693 558789
rect 216627 558724 216628 558788
rect 216692 558724 216693 558788
rect 216627 558723 216693 558724
rect 217366 557701 217426 560290
rect 217550 558925 217610 560430
rect 217950 559330 218010 560320
rect 217918 559270 218010 559330
rect 218838 560290 219024 560350
rect 217547 558924 217613 558925
rect 217547 558860 217548 558924
rect 217612 558860 217613 558924
rect 217547 558859 217613 558860
rect 217363 557700 217429 557701
rect 217363 557636 217364 557700
rect 217428 557636 217429 557700
rect 217363 557635 217429 557636
rect 217918 557565 217978 559270
rect 218838 558925 218898 560290
rect 219118 560010 219178 560320
rect 220126 560290 220192 560350
rect 220316 560290 220738 560350
rect 219118 559950 219266 560010
rect 218835 558924 218901 558925
rect 218835 558860 218836 558924
rect 218900 558860 218901 558924
rect 218835 558859 218901 558860
rect 219206 557565 219266 559950
rect 220126 559061 220186 560290
rect 220123 559060 220189 559061
rect 220123 558996 220124 559060
rect 220188 558996 220189 559060
rect 220123 558995 220189 558996
rect 220678 557565 220738 560290
rect 221046 558381 221106 560430
rect 221484 560290 222026 560350
rect 221043 558380 221109 558381
rect 221043 558316 221044 558380
rect 221108 558316 221109 558380
rect 221043 558315 221109 558316
rect 221966 557565 222026 560290
rect 222334 560290 222528 560350
rect 222652 560290 223314 560350
rect 222334 558925 222394 560290
rect 222331 558924 222397 558925
rect 222331 558860 222332 558924
rect 222396 558860 222397 558924
rect 222331 558859 222397 558860
rect 223254 557565 223314 560290
rect 223622 560290 223696 560350
rect 223820 560290 224418 560350
rect 223622 558925 223682 560290
rect 223619 558924 223685 558925
rect 223619 558860 223620 558924
rect 223684 558860 223685 558924
rect 223619 558859 223685 558860
rect 224358 557565 224418 560290
rect 224542 560290 224864 560350
rect 224988 560290 225706 560350
rect 224542 558925 224602 560290
rect 224539 558924 224605 558925
rect 224539 558860 224540 558924
rect 224604 558860 224605 558924
rect 224539 558859 224605 558860
rect 225646 557701 225706 560290
rect 225830 560290 226032 560350
rect 225830 558925 225890 560290
rect 226126 560010 226186 560320
rect 227118 560290 227200 560350
rect 227324 560290 227546 560350
rect 226126 559950 226258 560010
rect 225827 558924 225893 558925
rect 225827 558860 225828 558924
rect 225892 558860 225893 558924
rect 225827 558859 225893 558860
rect 225643 557700 225709 557701
rect 225643 557636 225644 557700
rect 225708 557636 225709 557700
rect 225643 557635 225709 557636
rect 226198 557565 226258 559950
rect 227118 558925 227178 560290
rect 227115 558924 227181 558925
rect 227115 558860 227116 558924
rect 227180 558860 227181 558924
rect 227115 558859 227181 558860
rect 227486 557565 227546 560290
rect 228338 559330 228398 560320
rect 228492 560290 228834 560350
rect 228222 559270 228398 559330
rect 228222 558925 228282 559270
rect 228219 558924 228285 558925
rect 228219 558860 228220 558924
rect 228284 558860 228285 558924
rect 228219 558859 228285 558860
rect 228774 557565 228834 560290
rect 229506 560010 229566 560320
rect 229660 560290 230306 560350
rect 229506 559950 229570 560010
rect 229510 558925 229570 559950
rect 229507 558924 229573 558925
rect 229507 558860 229508 558924
rect 229572 558860 229573 558924
rect 229507 558859 229573 558860
rect 230246 557565 230306 560290
rect 230614 560290 230704 560350
rect 230614 558381 230674 560290
rect 230611 558380 230677 558381
rect 230611 558316 230612 558380
rect 230676 558316 230677 558380
rect 230611 558315 230677 558316
rect 230798 557565 230858 560320
rect 231842 559330 231902 560320
rect 231996 560290 232698 560350
rect 231842 559270 231962 559330
rect 231902 558381 231962 559270
rect 231899 558380 231965 558381
rect 231899 558316 231900 558380
rect 231964 558316 231965 558380
rect 231899 558315 231965 558316
rect 232638 557701 232698 560290
rect 232822 560290 233040 560350
rect 232822 558789 232882 560290
rect 233134 559330 233194 560320
rect 233006 559270 233194 559330
rect 233558 560290 234208 560350
rect 234332 560290 234538 560350
rect 232819 558788 232885 558789
rect 232819 558724 232820 558788
rect 232884 558724 232885 558788
rect 232819 558723 232885 558724
rect 232635 557700 232701 557701
rect 232635 557636 232636 557700
rect 232700 557636 232701 557700
rect 232635 557635 232701 557636
rect 233006 557565 233066 559270
rect 233558 558789 233618 560290
rect 233555 558788 233621 558789
rect 233555 558724 233556 558788
rect 233620 558724 233621 558788
rect 233555 558723 233621 558724
rect 234478 557565 234538 560290
rect 235030 560290 235376 560350
rect 235500 560290 235826 560350
rect 235030 558653 235090 560290
rect 235027 558652 235093 558653
rect 235027 558588 235028 558652
rect 235092 558588 235093 558652
rect 235027 558587 235093 558588
rect 235766 557565 235826 560290
rect 236134 560290 236544 560350
rect 236668 560290 237298 560350
rect 236134 558517 236194 560290
rect 236131 558516 236197 558517
rect 236131 558452 236132 558516
rect 236196 558452 236197 558516
rect 236131 558451 236197 558452
rect 237238 557565 237298 560290
rect 237422 560290 237712 560350
rect 237836 560290 238402 560350
rect 237422 558653 237482 560290
rect 237419 558652 237485 558653
rect 237419 558588 237420 558652
rect 237484 558588 237485 558652
rect 237419 558587 237485 558588
rect 238342 557565 238402 560290
rect 238710 560290 238880 560350
rect 239004 560290 239690 560350
rect 238710 558517 238770 560290
rect 238707 558516 238773 558517
rect 238707 558452 238708 558516
rect 238772 558452 238773 558516
rect 238707 558451 238773 558452
rect 239630 557565 239690 560290
rect 270804 560218 270986 560454
rect 271222 560218 271404 560454
rect 270804 560134 271404 560218
rect 270804 559898 270986 560134
rect 271222 559898 271404 560134
rect 206875 557564 206941 557565
rect 206875 557500 206876 557564
rect 206940 557500 206941 557564
rect 206875 557499 206941 557500
rect 207979 557564 208045 557565
rect 207979 557500 207980 557564
rect 208044 557500 208045 557564
rect 207979 557499 208045 557500
rect 209267 557564 209333 557565
rect 209267 557500 209268 557564
rect 209332 557500 209333 557564
rect 209267 557499 209333 557500
rect 212395 557564 212461 557565
rect 212395 557500 212396 557564
rect 212460 557500 212461 557564
rect 212395 557499 212461 557500
rect 213499 557564 213565 557565
rect 213499 557500 213500 557564
rect 213564 557500 213565 557564
rect 213499 557499 213565 557500
rect 214787 557564 214853 557565
rect 214787 557500 214788 557564
rect 214852 557500 214853 557564
rect 214787 557499 214853 557500
rect 216259 557564 216325 557565
rect 216259 557500 216260 557564
rect 216324 557500 216325 557564
rect 216259 557499 216325 557500
rect 217915 557564 217981 557565
rect 217915 557500 217916 557564
rect 217980 557500 217981 557564
rect 217915 557499 217981 557500
rect 219203 557564 219269 557565
rect 219203 557500 219204 557564
rect 219268 557500 219269 557564
rect 219203 557499 219269 557500
rect 220675 557564 220741 557565
rect 220675 557500 220676 557564
rect 220740 557500 220741 557564
rect 220675 557499 220741 557500
rect 221963 557564 222029 557565
rect 221963 557500 221964 557564
rect 222028 557500 222029 557564
rect 221963 557499 222029 557500
rect 223251 557564 223317 557565
rect 223251 557500 223252 557564
rect 223316 557500 223317 557564
rect 223251 557499 223317 557500
rect 224355 557564 224421 557565
rect 224355 557500 224356 557564
rect 224420 557500 224421 557564
rect 224355 557499 224421 557500
rect 226195 557564 226261 557565
rect 226195 557500 226196 557564
rect 226260 557500 226261 557564
rect 226195 557499 226261 557500
rect 227483 557564 227549 557565
rect 227483 557500 227484 557564
rect 227548 557500 227549 557564
rect 227483 557499 227549 557500
rect 228771 557564 228837 557565
rect 228771 557500 228772 557564
rect 228836 557500 228837 557564
rect 228771 557499 228837 557500
rect 230243 557564 230309 557565
rect 230243 557500 230244 557564
rect 230308 557500 230309 557564
rect 230243 557499 230309 557500
rect 230795 557564 230861 557565
rect 230795 557500 230796 557564
rect 230860 557500 230861 557564
rect 230795 557499 230861 557500
rect 233003 557564 233069 557565
rect 233003 557500 233004 557564
rect 233068 557500 233069 557564
rect 233003 557499 233069 557500
rect 234475 557564 234541 557565
rect 234475 557500 234476 557564
rect 234540 557500 234541 557564
rect 234475 557499 234541 557500
rect 235763 557564 235829 557565
rect 235763 557500 235764 557564
rect 235828 557500 235829 557564
rect 235763 557499 235829 557500
rect 237235 557564 237301 557565
rect 237235 557500 237236 557564
rect 237300 557500 237301 557564
rect 237235 557499 237301 557500
rect 238339 557564 238405 557565
rect 238339 557500 238340 557564
rect 238404 557500 238405 557564
rect 238339 557499 238405 557500
rect 239627 557564 239693 557565
rect 239627 557500 239628 557564
rect 239692 557500 239693 557564
rect 239627 557499 239693 557500
rect 184404 545818 184586 546054
rect 184822 545818 185004 546054
rect 184404 545734 185004 545818
rect 184404 545498 184586 545734
rect 184822 545498 185004 545734
rect 184404 543000 185004 545498
rect 188004 549654 188604 557000
rect 188004 549418 188186 549654
rect 188422 549418 188604 549654
rect 188004 549334 188604 549418
rect 188004 549098 188186 549334
rect 188422 549098 188604 549334
rect 188004 543000 188604 549098
rect 191604 553254 192204 557000
rect 191604 553018 191786 553254
rect 192022 553018 192204 553254
rect 191604 552934 192204 553018
rect 191604 552698 191786 552934
rect 192022 552698 192204 552934
rect 191604 543000 192204 552698
rect 198804 543000 199404 557000
rect 202404 543000 203004 557000
rect 206004 543000 206604 557000
rect 209604 543000 210204 557000
rect 216804 543000 217404 557000
rect 220404 546054 221004 557000
rect 220404 545818 220586 546054
rect 220822 545818 221004 546054
rect 220404 545734 221004 545818
rect 220404 545498 220586 545734
rect 220822 545498 221004 545734
rect 220404 543000 221004 545498
rect 224004 549654 224604 557000
rect 224004 549418 224186 549654
rect 224422 549418 224604 549654
rect 224004 549334 224604 549418
rect 224004 549098 224186 549334
rect 224422 549098 224604 549334
rect 224004 543000 224604 549098
rect 227604 553254 228204 557000
rect 227604 553018 227786 553254
rect 228022 553018 228204 553254
rect 227604 552934 228204 553018
rect 227604 552698 227786 552934
rect 228022 552698 228204 552934
rect 227604 543000 228204 552698
rect 234804 543000 235404 557000
rect 238404 543000 239004 557000
rect 242004 543000 242604 557000
rect 245604 543000 246204 557000
rect 252804 543000 253404 557000
rect 256404 546054 257004 557000
rect 256404 545818 256586 546054
rect 256822 545818 257004 546054
rect 256404 545734 257004 545818
rect 256404 545498 256586 545734
rect 256822 545498 257004 545734
rect 256404 543000 257004 545498
rect 260004 549654 260604 557000
rect 260004 549418 260186 549654
rect 260422 549418 260604 549654
rect 260004 549334 260604 549418
rect 260004 549098 260186 549334
rect 260422 549098 260604 549334
rect 260004 543000 260604 549098
rect 263604 553254 264204 557000
rect 263604 553018 263786 553254
rect 264022 553018 264204 553254
rect 263604 552934 264204 553018
rect 263604 552698 263786 552934
rect 264022 552698 264204 552934
rect 263604 543000 264204 552698
rect 270804 543000 271404 559898
rect 274404 672054 275004 707102
rect 274404 671818 274586 672054
rect 274822 671818 275004 672054
rect 274404 671734 275004 671818
rect 274404 671498 274586 671734
rect 274822 671498 275004 671734
rect 274404 636054 275004 671498
rect 274404 635818 274586 636054
rect 274822 635818 275004 636054
rect 274404 635734 275004 635818
rect 274404 635498 274586 635734
rect 274822 635498 275004 635734
rect 274404 600054 275004 635498
rect 274404 599818 274586 600054
rect 274822 599818 275004 600054
rect 274404 599734 275004 599818
rect 274404 599498 274586 599734
rect 274822 599498 275004 599734
rect 274404 564054 275004 599498
rect 274404 563818 274586 564054
rect 274822 563818 275004 564054
rect 274404 563734 275004 563818
rect 274404 563498 274586 563734
rect 274822 563498 275004 563734
rect 274404 543000 275004 563498
rect 278004 675654 278604 708982
rect 278004 675418 278186 675654
rect 278422 675418 278604 675654
rect 278004 675334 278604 675418
rect 278004 675098 278186 675334
rect 278422 675098 278604 675334
rect 278004 639654 278604 675098
rect 278004 639418 278186 639654
rect 278422 639418 278604 639654
rect 278004 639334 278604 639418
rect 278004 639098 278186 639334
rect 278422 639098 278604 639334
rect 278004 603654 278604 639098
rect 278004 603418 278186 603654
rect 278422 603418 278604 603654
rect 278004 603334 278604 603418
rect 278004 603098 278186 603334
rect 278422 603098 278604 603334
rect 278004 567654 278604 603098
rect 278004 567418 278186 567654
rect 278422 567418 278604 567654
rect 278004 567334 278604 567418
rect 278004 567098 278186 567334
rect 278422 567098 278604 567334
rect 278004 543000 278604 567098
rect 281604 679254 282204 710862
rect 299604 710478 300204 711440
rect 299604 710242 299786 710478
rect 300022 710242 300204 710478
rect 299604 710158 300204 710242
rect 299604 709922 299786 710158
rect 300022 709922 300204 710158
rect 296004 708598 296604 709560
rect 296004 708362 296186 708598
rect 296422 708362 296604 708598
rect 296004 708278 296604 708362
rect 296004 708042 296186 708278
rect 296422 708042 296604 708278
rect 292404 706718 293004 707680
rect 292404 706482 292586 706718
rect 292822 706482 293004 706718
rect 292404 706398 293004 706482
rect 292404 706162 292586 706398
rect 292822 706162 293004 706398
rect 281604 679018 281786 679254
rect 282022 679018 282204 679254
rect 281604 678934 282204 679018
rect 281604 678698 281786 678934
rect 282022 678698 282204 678934
rect 281604 643254 282204 678698
rect 281604 643018 281786 643254
rect 282022 643018 282204 643254
rect 281604 642934 282204 643018
rect 281604 642698 281786 642934
rect 282022 642698 282204 642934
rect 281604 607254 282204 642698
rect 281604 607018 281786 607254
rect 282022 607018 282204 607254
rect 281604 606934 282204 607018
rect 281604 606698 281786 606934
rect 282022 606698 282204 606934
rect 281604 571254 282204 606698
rect 281604 571018 281786 571254
rect 282022 571018 282204 571254
rect 281604 570934 282204 571018
rect 281604 570698 281786 570934
rect 282022 570698 282204 570934
rect 281604 543000 282204 570698
rect 288804 704838 289404 705800
rect 288804 704602 288986 704838
rect 289222 704602 289404 704838
rect 288804 704518 289404 704602
rect 288804 704282 288986 704518
rect 289222 704282 289404 704518
rect 288804 686454 289404 704282
rect 288804 686218 288986 686454
rect 289222 686218 289404 686454
rect 288804 686134 289404 686218
rect 288804 685898 288986 686134
rect 289222 685898 289404 686134
rect 288804 650454 289404 685898
rect 288804 650218 288986 650454
rect 289222 650218 289404 650454
rect 288804 650134 289404 650218
rect 288804 649898 288986 650134
rect 289222 649898 289404 650134
rect 288804 614454 289404 649898
rect 288804 614218 288986 614454
rect 289222 614218 289404 614454
rect 288804 614134 289404 614218
rect 288804 613898 288986 614134
rect 289222 613898 289404 614134
rect 288804 578454 289404 613898
rect 288804 578218 288986 578454
rect 289222 578218 289404 578454
rect 288804 578134 289404 578218
rect 288804 577898 288986 578134
rect 289222 577898 289404 578134
rect 282315 558652 282381 558653
rect 282315 558588 282316 558652
rect 282380 558588 282381 558652
rect 282315 558587 282381 558588
rect 59491 540428 59557 540429
rect 59491 540364 59492 540428
rect 59556 540364 59557 540428
rect 59491 540363 59557 540364
rect 59494 407829 59554 540363
rect 79568 535254 79888 535276
rect 79568 535018 79610 535254
rect 79846 535018 79888 535254
rect 79568 534934 79888 535018
rect 79568 534698 79610 534934
rect 79846 534698 79888 534934
rect 79568 534676 79888 534698
rect 79568 531654 79888 531676
rect 79568 531418 79610 531654
rect 79846 531418 79888 531654
rect 79568 531334 79888 531418
rect 79568 531098 79610 531334
rect 79846 531098 79888 531334
rect 79568 531076 79888 531098
rect 79568 528054 79888 528076
rect 79568 527818 79610 528054
rect 79846 527818 79888 528054
rect 79568 527734 79888 527818
rect 79568 527498 79610 527734
rect 79846 527498 79888 527734
rect 79568 527476 79888 527498
rect 79568 524454 79888 524476
rect 79568 524218 79610 524454
rect 79846 524218 79888 524454
rect 79568 524134 79888 524218
rect 79568 523898 79610 524134
rect 79846 523898 79888 524134
rect 79568 523876 79888 523898
rect 64208 517254 64528 517276
rect 64208 517018 64250 517254
rect 64486 517018 64528 517254
rect 64208 516934 64528 517018
rect 64208 516698 64250 516934
rect 64486 516698 64528 516934
rect 64208 516676 64528 516698
rect 64208 513654 64528 513676
rect 64208 513418 64250 513654
rect 64486 513418 64528 513654
rect 64208 513334 64528 513418
rect 64208 513098 64250 513334
rect 64486 513098 64528 513334
rect 64208 513076 64528 513098
rect 64208 510054 64528 510076
rect 64208 509818 64250 510054
rect 64486 509818 64528 510054
rect 64208 509734 64528 509818
rect 64208 509498 64250 509734
rect 64486 509498 64528 509734
rect 64208 509476 64528 509498
rect 64208 506454 64528 506476
rect 64208 506218 64250 506454
rect 64486 506218 64528 506454
rect 64208 506134 64528 506218
rect 64208 505898 64250 506134
rect 64486 505898 64528 506134
rect 64208 505876 64528 505898
rect 79568 499254 79888 499276
rect 79568 499018 79610 499254
rect 79846 499018 79888 499254
rect 79568 498934 79888 499018
rect 79568 498698 79610 498934
rect 79846 498698 79888 498934
rect 79568 498676 79888 498698
rect 79568 495654 79888 495676
rect 79568 495418 79610 495654
rect 79846 495418 79888 495654
rect 79568 495334 79888 495418
rect 79568 495098 79610 495334
rect 79846 495098 79888 495334
rect 79568 495076 79888 495098
rect 79568 492054 79888 492076
rect 79568 491818 79610 492054
rect 79846 491818 79888 492054
rect 79568 491734 79888 491818
rect 79568 491498 79610 491734
rect 79846 491498 79888 491734
rect 79568 491476 79888 491498
rect 79568 488454 79888 488476
rect 79568 488218 79610 488454
rect 79846 488218 79888 488454
rect 79568 488134 79888 488218
rect 79568 487898 79610 488134
rect 79846 487898 79888 488134
rect 79568 487876 79888 487898
rect 64208 481254 64528 481276
rect 64208 481018 64250 481254
rect 64486 481018 64528 481254
rect 64208 480934 64528 481018
rect 64208 480698 64250 480934
rect 64486 480698 64528 480934
rect 64208 480676 64528 480698
rect 64208 477654 64528 477676
rect 64208 477418 64250 477654
rect 64486 477418 64528 477654
rect 64208 477334 64528 477418
rect 64208 477098 64250 477334
rect 64486 477098 64528 477334
rect 64208 477076 64528 477098
rect 64208 474054 64528 474076
rect 64208 473818 64250 474054
rect 64486 473818 64528 474054
rect 64208 473734 64528 473818
rect 64208 473498 64250 473734
rect 64486 473498 64528 473734
rect 64208 473476 64528 473498
rect 64208 470454 64528 470476
rect 64208 470218 64250 470454
rect 64486 470218 64528 470454
rect 64208 470134 64528 470218
rect 64208 469898 64250 470134
rect 64486 469898 64528 470134
rect 64208 469876 64528 469898
rect 79568 463254 79888 463276
rect 79568 463018 79610 463254
rect 79846 463018 79888 463254
rect 79568 462934 79888 463018
rect 79568 462698 79610 462934
rect 79846 462698 79888 462934
rect 79568 462676 79888 462698
rect 79568 459654 79888 459676
rect 79568 459418 79610 459654
rect 79846 459418 79888 459654
rect 79568 459334 79888 459418
rect 79568 459098 79610 459334
rect 79846 459098 79888 459334
rect 79568 459076 79888 459098
rect 79568 456054 79888 456076
rect 79568 455818 79610 456054
rect 79846 455818 79888 456054
rect 79568 455734 79888 455818
rect 79568 455498 79610 455734
rect 79846 455498 79888 455734
rect 79568 455476 79888 455498
rect 79568 452454 79888 452476
rect 79568 452218 79610 452454
rect 79846 452218 79888 452454
rect 79568 452134 79888 452218
rect 79568 451898 79610 452134
rect 79846 451898 79888 452134
rect 79568 451876 79888 451898
rect 64208 445254 64528 445276
rect 64208 445018 64250 445254
rect 64486 445018 64528 445254
rect 64208 444934 64528 445018
rect 64208 444698 64250 444934
rect 64486 444698 64528 444934
rect 64208 444676 64528 444698
rect 64208 441654 64528 441676
rect 64208 441418 64250 441654
rect 64486 441418 64528 441654
rect 64208 441334 64528 441418
rect 64208 441098 64250 441334
rect 64486 441098 64528 441334
rect 64208 441076 64528 441098
rect 64208 438054 64528 438076
rect 64208 437818 64250 438054
rect 64486 437818 64528 438054
rect 64208 437734 64528 437818
rect 64208 437498 64250 437734
rect 64486 437498 64528 437734
rect 64208 437476 64528 437498
rect 64208 434454 64528 434476
rect 64208 434218 64250 434454
rect 64486 434218 64528 434454
rect 64208 434134 64528 434218
rect 64208 433898 64250 434134
rect 64486 433898 64528 434134
rect 64208 433876 64528 433898
rect 79568 427254 79888 427276
rect 79568 427018 79610 427254
rect 79846 427018 79888 427254
rect 79568 426934 79888 427018
rect 79568 426698 79610 426934
rect 79846 426698 79888 426934
rect 79568 426676 79888 426698
rect 79568 423654 79888 423676
rect 79568 423418 79610 423654
rect 79846 423418 79888 423654
rect 79568 423334 79888 423418
rect 79568 423098 79610 423334
rect 79846 423098 79888 423334
rect 79568 423076 79888 423098
rect 79568 420054 79888 420076
rect 79568 419818 79610 420054
rect 79846 419818 79888 420054
rect 79568 419734 79888 419818
rect 79568 419498 79610 419734
rect 79846 419498 79888 419734
rect 79568 419476 79888 419498
rect 79568 416454 79888 416476
rect 79568 416218 79610 416454
rect 79846 416218 79888 416454
rect 79568 416134 79888 416218
rect 79568 415898 79610 416134
rect 79846 415898 79888 416134
rect 79568 415876 79888 415898
rect 281579 413948 281645 413949
rect 281579 413884 281580 413948
rect 281644 413884 281645 413948
rect 281579 413883 281645 413884
rect 64208 409254 64528 409276
rect 64208 409018 64250 409254
rect 64486 409018 64528 409254
rect 64208 408934 64528 409018
rect 64208 408698 64250 408934
rect 64486 408698 64528 408934
rect 64208 408676 64528 408698
rect 59491 407828 59557 407829
rect 59491 407764 59492 407828
rect 59556 407764 59557 407828
rect 59491 407763 59557 407764
rect 64208 405654 64528 405676
rect 64208 405418 64250 405654
rect 64486 405418 64528 405654
rect 64208 405334 64528 405418
rect 64208 405098 64250 405334
rect 64486 405098 64528 405334
rect 64208 405076 64528 405098
rect 59307 402116 59373 402117
rect 59307 402052 59308 402116
rect 59372 402052 59373 402116
rect 59307 402051 59373 402052
rect 64208 402054 64528 402076
rect 64208 401818 64250 402054
rect 64486 401818 64528 402054
rect 64208 401734 64528 401818
rect 64208 401498 64250 401734
rect 64486 401498 64528 401734
rect 64208 401476 64528 401498
rect 64208 398454 64528 398476
rect 64208 398218 64250 398454
rect 64486 398218 64528 398454
rect 58203 398172 58269 398173
rect 58203 398108 58204 398172
rect 58268 398108 58269 398172
rect 58203 398107 58269 398108
rect 64208 398134 64528 398218
rect 64208 397898 64250 398134
rect 64486 397898 64528 398134
rect 64208 397876 64528 397898
rect 79568 391254 79888 391276
rect 79568 391018 79610 391254
rect 79846 391018 79888 391254
rect 79568 390934 79888 391018
rect 79568 390698 79610 390934
rect 79846 390698 79888 390934
rect 79568 390676 79888 390698
rect 57467 388516 57533 388517
rect 57467 388452 57468 388516
rect 57532 388452 57533 388516
rect 57467 388451 57533 388452
rect 79568 387654 79888 387676
rect 79568 387418 79610 387654
rect 79846 387418 79888 387654
rect 79568 387334 79888 387418
rect 79568 387098 79610 387334
rect 79846 387098 79888 387334
rect 79568 387076 79888 387098
rect 79568 384054 79888 384076
rect 79568 383818 79610 384054
rect 79846 383818 79888 384054
rect 79568 383734 79888 383818
rect 79568 383498 79610 383734
rect 79846 383498 79888 383734
rect 79568 383476 79888 383498
rect 54804 380218 54986 380454
rect 55222 380218 55404 380454
rect 54804 380134 55404 380218
rect 54804 379898 54986 380134
rect 55222 379898 55404 380134
rect 54804 344454 55404 379898
rect 79568 380454 79888 380476
rect 79568 380218 79610 380454
rect 79846 380218 79888 380454
rect 79568 380134 79888 380218
rect 79568 379898 79610 380134
rect 79846 379898 79888 380134
rect 79568 379876 79888 379898
rect 57835 375052 57901 375053
rect 57835 374988 57836 375052
rect 57900 374988 57901 375052
rect 57835 374987 57901 374988
rect 56915 353836 56981 353837
rect 56915 353772 56916 353836
rect 56980 353772 56981 353836
rect 56915 353771 56981 353772
rect 54804 344218 54986 344454
rect 55222 344218 55404 344454
rect 54804 344134 55404 344218
rect 54804 343898 54986 344134
rect 55222 343898 55404 344134
rect 54804 308454 55404 343898
rect 54804 308218 54986 308454
rect 55222 308218 55404 308454
rect 54804 308134 55404 308218
rect 54804 307898 54986 308134
rect 55222 307898 55404 308134
rect 54804 272454 55404 307898
rect 54804 272218 54986 272454
rect 55222 272218 55404 272454
rect 54804 272134 55404 272218
rect 54804 271898 54986 272134
rect 55222 271898 55404 272134
rect 54804 236454 55404 271898
rect 56918 263941 56978 353771
rect 57283 347988 57349 347989
rect 57283 347924 57284 347988
rect 57348 347924 57349 347988
rect 57283 347923 57349 347924
rect 57099 346084 57165 346085
rect 57099 346020 57100 346084
rect 57164 346020 57165 346084
rect 57099 346019 57165 346020
rect 56915 263940 56981 263941
rect 56915 263876 56916 263940
rect 56980 263876 56981 263940
rect 56915 263875 56981 263876
rect 54804 236218 54986 236454
rect 55222 236218 55404 236454
rect 54804 236134 55404 236218
rect 54804 235898 54986 236134
rect 55222 235898 55404 236134
rect 54804 200454 55404 235898
rect 57102 228037 57162 346019
rect 57099 228036 57165 228037
rect 57099 227972 57100 228036
rect 57164 227972 57165 228036
rect 57099 227971 57165 227972
rect 57286 217021 57346 347923
rect 57651 342276 57717 342277
rect 57651 342212 57652 342276
rect 57716 342212 57717 342276
rect 57651 342211 57717 342212
rect 57467 340236 57533 340237
rect 57467 340172 57468 340236
rect 57532 340172 57533 340236
rect 57467 340171 57533 340172
rect 57283 217020 57349 217021
rect 57283 216956 57284 217020
rect 57348 216956 57349 217020
rect 57283 216955 57349 216956
rect 54804 200218 54986 200454
rect 55222 200218 55404 200454
rect 54804 200134 55404 200218
rect 54804 199898 54986 200134
rect 55222 199898 55404 200134
rect 54804 164454 55404 199898
rect 57470 181117 57530 340171
rect 57467 181116 57533 181117
rect 57467 181052 57468 181116
rect 57532 181052 57533 181116
rect 57467 181051 57533 181052
rect 57654 170101 57714 342211
rect 57838 330717 57898 374987
rect 64208 373254 64528 373276
rect 64208 373018 64250 373254
rect 64486 373018 64528 373254
rect 64208 372934 64528 373018
rect 64208 372698 64250 372934
rect 64486 372698 64528 372934
rect 64208 372676 64528 372698
rect 64208 369654 64528 369676
rect 64208 369418 64250 369654
rect 64486 369418 64528 369654
rect 64208 369334 64528 369418
rect 64208 369098 64250 369334
rect 64486 369098 64528 369334
rect 64208 369076 64528 369098
rect 64208 366054 64528 366076
rect 64208 365818 64250 366054
rect 64486 365818 64528 366054
rect 64208 365734 64528 365818
rect 64208 365498 64250 365734
rect 64486 365498 64528 365734
rect 64208 365476 64528 365498
rect 64208 362454 64528 362476
rect 64208 362218 64250 362454
rect 64486 362218 64528 362454
rect 64208 362134 64528 362218
rect 64208 361898 64250 362134
rect 64486 361898 64528 362134
rect 64208 361876 64528 361898
rect 79568 355254 79888 355276
rect 79568 355018 79610 355254
rect 79846 355018 79888 355254
rect 79568 354934 79888 355018
rect 79568 354698 79610 354934
rect 79846 354698 79888 354934
rect 79568 354676 79888 354698
rect 79568 351654 79888 351676
rect 79568 351418 79610 351654
rect 79846 351418 79888 351654
rect 79568 351334 79888 351418
rect 79568 351098 79610 351334
rect 79846 351098 79888 351334
rect 79568 351076 79888 351098
rect 79568 348054 79888 348076
rect 79568 347818 79610 348054
rect 79846 347818 79888 348054
rect 79568 347734 79888 347818
rect 79568 347498 79610 347734
rect 79846 347498 79888 347734
rect 79568 347476 79888 347498
rect 79568 344454 79888 344476
rect 79568 344218 79610 344454
rect 79846 344218 79888 344454
rect 79568 344134 79888 344218
rect 79568 343898 79610 344134
rect 79846 343898 79888 344134
rect 79568 343876 79888 343898
rect 64208 337254 64528 337276
rect 64208 337018 64250 337254
rect 64486 337018 64528 337254
rect 64208 336934 64528 337018
rect 64208 336698 64250 336934
rect 64486 336698 64528 336934
rect 64208 336676 64528 336698
rect 64208 333654 64528 333676
rect 64208 333418 64250 333654
rect 64486 333418 64528 333654
rect 64208 333334 64528 333418
rect 64208 333098 64250 333334
rect 64486 333098 64528 333334
rect 64208 333076 64528 333098
rect 57835 330716 57901 330717
rect 57835 330652 57836 330716
rect 57900 330652 57901 330716
rect 57835 330651 57901 330652
rect 57835 330580 57901 330581
rect 57835 330516 57836 330580
rect 57900 330516 57901 330580
rect 57835 330515 57901 330516
rect 57651 170100 57717 170101
rect 57651 170036 57652 170100
rect 57716 170036 57717 170100
rect 57651 170035 57717 170036
rect 54804 164218 54986 164454
rect 55222 164218 55404 164454
rect 54804 164134 55404 164218
rect 54804 163898 54986 164134
rect 55222 163898 55404 164134
rect 54804 128454 55404 163898
rect 54804 128218 54986 128454
rect 55222 128218 55404 128454
rect 54804 128134 55404 128218
rect 54804 127898 54986 128134
rect 55222 127898 55404 128134
rect 54804 92454 55404 127898
rect 54804 92218 54986 92454
rect 55222 92218 55404 92454
rect 54804 92134 55404 92218
rect 54804 91898 54986 92134
rect 55222 91898 55404 92134
rect 54804 56454 55404 91898
rect 57838 76261 57898 330515
rect 64208 330054 64528 330076
rect 64208 329818 64250 330054
rect 64486 329818 64528 330054
rect 64208 329734 64528 329818
rect 64208 329498 64250 329734
rect 64486 329498 64528 329734
rect 64208 329476 64528 329498
rect 64208 326454 64528 326476
rect 64208 326218 64250 326454
rect 64486 326218 64528 326454
rect 64208 326134 64528 326218
rect 64208 325898 64250 326134
rect 64486 325898 64528 326134
rect 64208 325876 64528 325898
rect 281582 317389 281642 413883
rect 282318 391101 282378 558587
rect 283419 558516 283485 558517
rect 283419 558452 283420 558516
rect 283484 558452 283485 558516
rect 283419 558451 283485 558452
rect 283422 395181 283482 558451
rect 283787 558380 283853 558381
rect 283787 558316 283788 558380
rect 283852 558316 283853 558380
rect 283787 558315 283853 558316
rect 283603 558244 283669 558245
rect 283603 558180 283604 558244
rect 283668 558180 283669 558244
rect 283603 558179 283669 558180
rect 283606 397221 283666 558179
rect 283603 397220 283669 397221
rect 283603 397156 283604 397220
rect 283668 397156 283669 397220
rect 283603 397155 283669 397156
rect 283790 396133 283850 558315
rect 288804 542454 289404 577898
rect 288804 542218 288986 542454
rect 289222 542218 289404 542454
rect 288804 542134 289404 542218
rect 288804 541898 288986 542134
rect 289222 541898 289404 542134
rect 288804 506454 289404 541898
rect 288804 506218 288986 506454
rect 289222 506218 289404 506454
rect 288804 506134 289404 506218
rect 288804 505898 288986 506134
rect 289222 505898 289404 506134
rect 288804 470454 289404 505898
rect 288804 470218 288986 470454
rect 289222 470218 289404 470454
rect 288804 470134 289404 470218
rect 288804 469898 288986 470134
rect 289222 469898 289404 470134
rect 288804 434454 289404 469898
rect 288804 434218 288986 434454
rect 289222 434218 289404 434454
rect 288804 434134 289404 434218
rect 288804 433898 288986 434134
rect 289222 433898 289404 434134
rect 288804 398454 289404 433898
rect 288804 398218 288986 398454
rect 289222 398218 289404 398454
rect 288804 398134 289404 398218
rect 288804 397898 288986 398134
rect 289222 397898 289404 398134
rect 283787 396132 283853 396133
rect 283787 396068 283788 396132
rect 283852 396068 283853 396132
rect 283787 396067 283853 396068
rect 283419 395180 283485 395181
rect 283419 395116 283420 395180
rect 283484 395116 283485 395180
rect 283419 395115 283485 395116
rect 282315 391100 282381 391101
rect 282315 391036 282316 391100
rect 282380 391036 282381 391100
rect 282315 391035 282381 391036
rect 288804 362454 289404 397898
rect 288804 362218 288986 362454
rect 289222 362218 289404 362454
rect 288804 362134 289404 362218
rect 288804 361898 288986 362134
rect 289222 361898 289404 362134
rect 288804 326454 289404 361898
rect 288804 326218 288986 326454
rect 289222 326218 289404 326454
rect 288804 326134 289404 326218
rect 288804 325898 288986 326134
rect 289222 325898 289404 326134
rect 281579 317388 281645 317389
rect 281579 317324 281580 317388
rect 281644 317324 281645 317388
rect 281579 317323 281645 317324
rect 58404 312054 59004 317000
rect 58404 311818 58586 312054
rect 58822 311818 59004 312054
rect 58404 311734 59004 311818
rect 58404 311498 58586 311734
rect 58822 311498 59004 311734
rect 58404 276054 59004 311498
rect 58404 275818 58586 276054
rect 58822 275818 59004 276054
rect 58404 275734 59004 275818
rect 58404 275498 58586 275734
rect 58822 275498 59004 275734
rect 58404 240054 59004 275498
rect 58404 239818 58586 240054
rect 58822 239818 59004 240054
rect 58404 239734 59004 239818
rect 58404 239498 58586 239734
rect 58822 239498 59004 239734
rect 58404 204054 59004 239498
rect 58404 203818 58586 204054
rect 58822 203818 59004 204054
rect 58404 203734 59004 203818
rect 58404 203498 58586 203734
rect 58822 203498 59004 203734
rect 58404 168054 59004 203498
rect 58404 167818 58586 168054
rect 58822 167818 59004 168054
rect 58404 167734 59004 167818
rect 58404 167498 58586 167734
rect 58822 167498 59004 167734
rect 58404 132054 59004 167498
rect 58404 131818 58586 132054
rect 58822 131818 59004 132054
rect 58404 131734 59004 131818
rect 58404 131498 58586 131734
rect 58822 131498 59004 131734
rect 58404 96054 59004 131498
rect 58404 95818 58586 96054
rect 58822 95818 59004 96054
rect 58404 95734 59004 95818
rect 58404 95498 58586 95734
rect 58822 95498 59004 95734
rect 57835 76260 57901 76261
rect 57835 76196 57836 76260
rect 57900 76196 57901 76260
rect 57835 76195 57901 76196
rect 54804 56218 54986 56454
rect 55222 56218 55404 56454
rect 54804 56134 55404 56218
rect 54804 55898 54986 56134
rect 55222 55898 55404 56134
rect 54804 20454 55404 55898
rect 54804 20218 54986 20454
rect 55222 20218 55404 20454
rect 54804 20134 55404 20218
rect 54804 19898 54986 20134
rect 55222 19898 55404 20134
rect 54804 -1286 55404 19898
rect 54804 -1522 54986 -1286
rect 55222 -1522 55404 -1286
rect 54804 -1606 55404 -1522
rect 54804 -1842 54986 -1606
rect 55222 -1842 55404 -1606
rect 54804 -1864 55404 -1842
rect 58404 60054 59004 95498
rect 58404 59818 58586 60054
rect 58822 59818 59004 60054
rect 58404 59734 59004 59818
rect 58404 59498 58586 59734
rect 58822 59498 59004 59734
rect 58404 24054 59004 59498
rect 58404 23818 58586 24054
rect 58822 23818 59004 24054
rect 58404 23734 59004 23818
rect 58404 23498 58586 23734
rect 58822 23498 59004 23734
rect 58404 -3166 59004 23498
rect 58404 -3402 58586 -3166
rect 58822 -3402 59004 -3166
rect 58404 -3486 59004 -3402
rect 58404 -3722 58586 -3486
rect 58822 -3722 59004 -3486
rect 58404 -3744 59004 -3722
rect 62004 315654 62604 317000
rect 62004 315418 62186 315654
rect 62422 315418 62604 315654
rect 62004 315334 62604 315418
rect 62004 315098 62186 315334
rect 62422 315098 62604 315334
rect 62004 279654 62604 315098
rect 62004 279418 62186 279654
rect 62422 279418 62604 279654
rect 62004 279334 62604 279418
rect 62004 279098 62186 279334
rect 62422 279098 62604 279334
rect 62004 243654 62604 279098
rect 62004 243418 62186 243654
rect 62422 243418 62604 243654
rect 62004 243334 62604 243418
rect 62004 243098 62186 243334
rect 62422 243098 62604 243334
rect 62004 207654 62604 243098
rect 62004 207418 62186 207654
rect 62422 207418 62604 207654
rect 62004 207334 62604 207418
rect 62004 207098 62186 207334
rect 62422 207098 62604 207334
rect 62004 171654 62604 207098
rect 62004 171418 62186 171654
rect 62422 171418 62604 171654
rect 62004 171334 62604 171418
rect 62004 171098 62186 171334
rect 62422 171098 62604 171334
rect 62004 135654 62604 171098
rect 62004 135418 62186 135654
rect 62422 135418 62604 135654
rect 62004 135334 62604 135418
rect 62004 135098 62186 135334
rect 62422 135098 62604 135334
rect 62004 99654 62604 135098
rect 62004 99418 62186 99654
rect 62422 99418 62604 99654
rect 62004 99334 62604 99418
rect 62004 99098 62186 99334
rect 62422 99098 62604 99334
rect 62004 63654 62604 99098
rect 62004 63418 62186 63654
rect 62422 63418 62604 63654
rect 62004 63334 62604 63418
rect 62004 63098 62186 63334
rect 62422 63098 62604 63334
rect 62004 27654 62604 63098
rect 62004 27418 62186 27654
rect 62422 27418 62604 27654
rect 62004 27334 62604 27418
rect 62004 27098 62186 27334
rect 62422 27098 62604 27334
rect 62004 -5046 62604 27098
rect 62004 -5282 62186 -5046
rect 62422 -5282 62604 -5046
rect 62004 -5366 62604 -5282
rect 62004 -5602 62186 -5366
rect 62422 -5602 62604 -5366
rect 62004 -5624 62604 -5602
rect 65604 283254 66204 317000
rect 65604 283018 65786 283254
rect 66022 283018 66204 283254
rect 65604 282934 66204 283018
rect 65604 282698 65786 282934
rect 66022 282698 66204 282934
rect 65604 247254 66204 282698
rect 65604 247018 65786 247254
rect 66022 247018 66204 247254
rect 65604 246934 66204 247018
rect 65604 246698 65786 246934
rect 66022 246698 66204 246934
rect 65604 211254 66204 246698
rect 65604 211018 65786 211254
rect 66022 211018 66204 211254
rect 65604 210934 66204 211018
rect 65604 210698 65786 210934
rect 66022 210698 66204 210934
rect 65604 175254 66204 210698
rect 65604 175018 65786 175254
rect 66022 175018 66204 175254
rect 65604 174934 66204 175018
rect 65604 174698 65786 174934
rect 66022 174698 66204 174934
rect 65604 139254 66204 174698
rect 65604 139018 65786 139254
rect 66022 139018 66204 139254
rect 65604 138934 66204 139018
rect 65604 138698 65786 138934
rect 66022 138698 66204 138934
rect 65604 103254 66204 138698
rect 65604 103018 65786 103254
rect 66022 103018 66204 103254
rect 65604 102934 66204 103018
rect 65604 102698 65786 102934
rect 66022 102698 66204 102934
rect 65604 67254 66204 102698
rect 65604 67018 65786 67254
rect 66022 67018 66204 67254
rect 65604 66934 66204 67018
rect 65604 66698 65786 66934
rect 66022 66698 66204 66934
rect 65604 31254 66204 66698
rect 65604 31018 65786 31254
rect 66022 31018 66204 31254
rect 65604 30934 66204 31018
rect 65604 30698 65786 30934
rect 66022 30698 66204 30934
rect 47604 -6222 47786 -5986
rect 48022 -6222 48204 -5986
rect 47604 -6306 48204 -6222
rect 47604 -6542 47786 -6306
rect 48022 -6542 48204 -6306
rect 47604 -7504 48204 -6542
rect 65604 -6926 66204 30698
rect 72804 290454 73404 317000
rect 72804 290218 72986 290454
rect 73222 290218 73404 290454
rect 72804 290134 73404 290218
rect 72804 289898 72986 290134
rect 73222 289898 73404 290134
rect 72804 254454 73404 289898
rect 72804 254218 72986 254454
rect 73222 254218 73404 254454
rect 72804 254134 73404 254218
rect 72804 253898 72986 254134
rect 73222 253898 73404 254134
rect 72804 218454 73404 253898
rect 72804 218218 72986 218454
rect 73222 218218 73404 218454
rect 72804 218134 73404 218218
rect 72804 217898 72986 218134
rect 73222 217898 73404 218134
rect 72804 182454 73404 217898
rect 72804 182218 72986 182454
rect 73222 182218 73404 182454
rect 72804 182134 73404 182218
rect 72804 181898 72986 182134
rect 73222 181898 73404 182134
rect 72804 146454 73404 181898
rect 72804 146218 72986 146454
rect 73222 146218 73404 146454
rect 72804 146134 73404 146218
rect 72804 145898 72986 146134
rect 73222 145898 73404 146134
rect 72804 110454 73404 145898
rect 72804 110218 72986 110454
rect 73222 110218 73404 110454
rect 72804 110134 73404 110218
rect 72804 109898 72986 110134
rect 73222 109898 73404 110134
rect 72804 74454 73404 109898
rect 72804 74218 72986 74454
rect 73222 74218 73404 74454
rect 72804 74134 73404 74218
rect 72804 73898 72986 74134
rect 73222 73898 73404 74134
rect 72804 38454 73404 73898
rect 72804 38218 72986 38454
rect 73222 38218 73404 38454
rect 72804 38134 73404 38218
rect 72804 37898 72986 38134
rect 73222 37898 73404 38134
rect 72804 2454 73404 37898
rect 72804 2218 72986 2454
rect 73222 2218 73404 2454
rect 72804 2134 73404 2218
rect 72804 1898 72986 2134
rect 73222 1898 73404 2134
rect 72804 -346 73404 1898
rect 72804 -582 72986 -346
rect 73222 -582 73404 -346
rect 72804 -666 73404 -582
rect 72804 -902 72986 -666
rect 73222 -902 73404 -666
rect 72804 -1864 73404 -902
rect 76404 294054 77004 317000
rect 76404 293818 76586 294054
rect 76822 293818 77004 294054
rect 76404 293734 77004 293818
rect 76404 293498 76586 293734
rect 76822 293498 77004 293734
rect 76404 258054 77004 293498
rect 76404 257818 76586 258054
rect 76822 257818 77004 258054
rect 76404 257734 77004 257818
rect 76404 257498 76586 257734
rect 76822 257498 77004 257734
rect 76404 222054 77004 257498
rect 76404 221818 76586 222054
rect 76822 221818 77004 222054
rect 76404 221734 77004 221818
rect 76404 221498 76586 221734
rect 76822 221498 77004 221734
rect 76404 186054 77004 221498
rect 76404 185818 76586 186054
rect 76822 185818 77004 186054
rect 76404 185734 77004 185818
rect 76404 185498 76586 185734
rect 76822 185498 77004 185734
rect 76404 150054 77004 185498
rect 76404 149818 76586 150054
rect 76822 149818 77004 150054
rect 76404 149734 77004 149818
rect 76404 149498 76586 149734
rect 76822 149498 77004 149734
rect 76404 114054 77004 149498
rect 76404 113818 76586 114054
rect 76822 113818 77004 114054
rect 76404 113734 77004 113818
rect 76404 113498 76586 113734
rect 76822 113498 77004 113734
rect 76404 78054 77004 113498
rect 76404 77818 76586 78054
rect 76822 77818 77004 78054
rect 76404 77734 77004 77818
rect 76404 77498 76586 77734
rect 76822 77498 77004 77734
rect 76404 42054 77004 77498
rect 76404 41818 76586 42054
rect 76822 41818 77004 42054
rect 76404 41734 77004 41818
rect 76404 41498 76586 41734
rect 76822 41498 77004 41734
rect 76404 6054 77004 41498
rect 76404 5818 76586 6054
rect 76822 5818 77004 6054
rect 76404 5734 77004 5818
rect 76404 5498 76586 5734
rect 76822 5498 77004 5734
rect 76404 -2226 77004 5498
rect 76404 -2462 76586 -2226
rect 76822 -2462 77004 -2226
rect 76404 -2546 77004 -2462
rect 76404 -2782 76586 -2546
rect 76822 -2782 77004 -2546
rect 76404 -3744 77004 -2782
rect 80004 297654 80604 317000
rect 80004 297418 80186 297654
rect 80422 297418 80604 297654
rect 80004 297334 80604 297418
rect 80004 297098 80186 297334
rect 80422 297098 80604 297334
rect 80004 261654 80604 297098
rect 80004 261418 80186 261654
rect 80422 261418 80604 261654
rect 80004 261334 80604 261418
rect 80004 261098 80186 261334
rect 80422 261098 80604 261334
rect 80004 225654 80604 261098
rect 80004 225418 80186 225654
rect 80422 225418 80604 225654
rect 80004 225334 80604 225418
rect 80004 225098 80186 225334
rect 80422 225098 80604 225334
rect 80004 189654 80604 225098
rect 80004 189418 80186 189654
rect 80422 189418 80604 189654
rect 80004 189334 80604 189418
rect 80004 189098 80186 189334
rect 80422 189098 80604 189334
rect 80004 153654 80604 189098
rect 80004 153418 80186 153654
rect 80422 153418 80604 153654
rect 80004 153334 80604 153418
rect 80004 153098 80186 153334
rect 80422 153098 80604 153334
rect 80004 117654 80604 153098
rect 80004 117418 80186 117654
rect 80422 117418 80604 117654
rect 80004 117334 80604 117418
rect 80004 117098 80186 117334
rect 80422 117098 80604 117334
rect 80004 81654 80604 117098
rect 80004 81418 80186 81654
rect 80422 81418 80604 81654
rect 80004 81334 80604 81418
rect 80004 81098 80186 81334
rect 80422 81098 80604 81334
rect 80004 45654 80604 81098
rect 80004 45418 80186 45654
rect 80422 45418 80604 45654
rect 80004 45334 80604 45418
rect 80004 45098 80186 45334
rect 80422 45098 80604 45334
rect 80004 9654 80604 45098
rect 80004 9418 80186 9654
rect 80422 9418 80604 9654
rect 80004 9334 80604 9418
rect 80004 9098 80186 9334
rect 80422 9098 80604 9334
rect 80004 -4106 80604 9098
rect 80004 -4342 80186 -4106
rect 80422 -4342 80604 -4106
rect 80004 -4426 80604 -4342
rect 80004 -4662 80186 -4426
rect 80422 -4662 80604 -4426
rect 80004 -5624 80604 -4662
rect 83604 301254 84204 317000
rect 83604 301018 83786 301254
rect 84022 301018 84204 301254
rect 83604 300934 84204 301018
rect 83604 300698 83786 300934
rect 84022 300698 84204 300934
rect 83604 265254 84204 300698
rect 83604 265018 83786 265254
rect 84022 265018 84204 265254
rect 83604 264934 84204 265018
rect 83604 264698 83786 264934
rect 84022 264698 84204 264934
rect 83604 229254 84204 264698
rect 90804 308454 91404 317000
rect 90804 308218 90986 308454
rect 91222 308218 91404 308454
rect 90804 308134 91404 308218
rect 90804 307898 90986 308134
rect 91222 307898 91404 308134
rect 90804 272454 91404 307898
rect 90804 272218 90986 272454
rect 91222 272218 91404 272454
rect 90804 272134 91404 272218
rect 90804 271898 90986 272134
rect 91222 271898 91404 272134
rect 86907 264076 86973 264077
rect 86907 264012 86908 264076
rect 86972 264012 86973 264076
rect 86907 264011 86973 264012
rect 86910 263669 86970 264011
rect 86907 263668 86973 263669
rect 86907 263604 86908 263668
rect 86972 263604 86973 263668
rect 86907 263603 86973 263604
rect 83604 229018 83786 229254
rect 84022 229018 84204 229254
rect 83604 228934 84204 229018
rect 83604 228698 83786 228934
rect 84022 228698 84204 228934
rect 83604 193254 84204 228698
rect 90804 236454 91404 271898
rect 90804 236218 90986 236454
rect 91222 236218 91404 236454
rect 90804 236134 91404 236218
rect 90804 235898 90986 236134
rect 91222 235898 91404 236134
rect 86907 227764 86973 227765
rect 86907 227700 86908 227764
rect 86972 227700 86973 227764
rect 86907 227699 86973 227700
rect 86910 227493 86970 227699
rect 86907 227492 86973 227493
rect 86907 227428 86908 227492
rect 86972 227428 86973 227492
rect 86907 227427 86973 227428
rect 83604 193018 83786 193254
rect 84022 193018 84204 193254
rect 83604 192934 84204 193018
rect 83604 192698 83786 192934
rect 84022 192698 84204 192934
rect 83604 157254 84204 192698
rect 83604 157018 83786 157254
rect 84022 157018 84204 157254
rect 83604 156934 84204 157018
rect 83604 156698 83786 156934
rect 84022 156698 84204 156934
rect 83604 121254 84204 156698
rect 83604 121018 83786 121254
rect 84022 121018 84204 121254
rect 83604 120934 84204 121018
rect 83604 120698 83786 120934
rect 84022 120698 84204 120934
rect 83604 85254 84204 120698
rect 83604 85018 83786 85254
rect 84022 85018 84204 85254
rect 83604 84934 84204 85018
rect 83604 84698 83786 84934
rect 84022 84698 84204 84934
rect 83604 49254 84204 84698
rect 83604 49018 83786 49254
rect 84022 49018 84204 49254
rect 83604 48934 84204 49018
rect 83604 48698 83786 48934
rect 84022 48698 84204 48934
rect 83604 13254 84204 48698
rect 90804 200454 91404 235898
rect 90804 200218 90986 200454
rect 91222 200218 91404 200454
rect 90804 200134 91404 200218
rect 90804 199898 90986 200134
rect 91222 199898 91404 200134
rect 90804 164454 91404 199898
rect 90804 164218 90986 164454
rect 91222 164218 91404 164454
rect 90804 164134 91404 164218
rect 90804 163898 90986 164134
rect 91222 163898 91404 164134
rect 90804 128454 91404 163898
rect 90804 128218 90986 128454
rect 91222 128218 91404 128454
rect 90804 128134 91404 128218
rect 90804 127898 90986 128134
rect 91222 127898 91404 128134
rect 90804 92454 91404 127898
rect 90804 92218 90986 92454
rect 91222 92218 91404 92454
rect 90804 92134 91404 92218
rect 90804 91898 90986 92134
rect 91222 91898 91404 92134
rect 90804 56454 91404 91898
rect 90804 56218 90986 56454
rect 91222 56218 91404 56454
rect 90804 56134 91404 56218
rect 90804 55898 90986 56134
rect 91222 55898 91404 56134
rect 89299 31788 89365 31789
rect 89299 31724 89300 31788
rect 89364 31724 89365 31788
rect 89299 31723 89365 31724
rect 89302 26349 89362 31723
rect 89299 26348 89365 26349
rect 89299 26284 89300 26348
rect 89364 26284 89365 26348
rect 89299 26283 89365 26284
rect 83604 13018 83786 13254
rect 84022 13018 84204 13254
rect 83604 12934 84204 13018
rect 83604 12698 83786 12934
rect 84022 12698 84204 12934
rect 65604 -7162 65786 -6926
rect 66022 -7162 66204 -6926
rect 65604 -7246 66204 -7162
rect 65604 -7482 65786 -7246
rect 66022 -7482 66204 -7246
rect 65604 -7504 66204 -7482
rect 83604 -5986 84204 12698
rect 90804 20454 91404 55898
rect 90804 20218 90986 20454
rect 91222 20218 91404 20454
rect 90804 20134 91404 20218
rect 90804 19898 90986 20134
rect 91222 19898 91404 20134
rect 90804 -1286 91404 19898
rect 90804 -1522 90986 -1286
rect 91222 -1522 91404 -1286
rect 90804 -1606 91404 -1522
rect 90804 -1842 90986 -1606
rect 91222 -1842 91404 -1606
rect 90804 -1864 91404 -1842
rect 94404 312054 95004 317000
rect 94404 311818 94586 312054
rect 94822 311818 95004 312054
rect 94404 311734 95004 311818
rect 94404 311498 94586 311734
rect 94822 311498 95004 311734
rect 94404 276054 95004 311498
rect 94404 275818 94586 276054
rect 94822 275818 95004 276054
rect 94404 275734 95004 275818
rect 94404 275498 94586 275734
rect 94822 275498 95004 275734
rect 94404 240054 95004 275498
rect 98004 315654 98604 317000
rect 98004 315418 98186 315654
rect 98422 315418 98604 315654
rect 98004 315334 98604 315418
rect 98004 315098 98186 315334
rect 98422 315098 98604 315334
rect 98004 279654 98604 315098
rect 98004 279418 98186 279654
rect 98422 279418 98604 279654
rect 98004 279334 98604 279418
rect 98004 279098 98186 279334
rect 98422 279098 98604 279334
rect 96475 264076 96541 264077
rect 96475 264012 96476 264076
rect 96540 264012 96541 264076
rect 96475 264011 96541 264012
rect 96478 263805 96538 264011
rect 96475 263804 96541 263805
rect 96475 263740 96476 263804
rect 96540 263740 96541 263804
rect 96475 263739 96541 263740
rect 94404 239818 94586 240054
rect 94822 239818 95004 240054
rect 94404 239734 95004 239818
rect 94404 239498 94586 239734
rect 94822 239498 95004 239734
rect 94404 204054 95004 239498
rect 98004 243654 98604 279098
rect 98004 243418 98186 243654
rect 98422 243418 98604 243654
rect 98004 243334 98604 243418
rect 98004 243098 98186 243334
rect 98422 243098 98604 243334
rect 96475 227900 96541 227901
rect 96475 227836 96476 227900
rect 96540 227836 96541 227900
rect 96475 227835 96541 227836
rect 96478 227493 96538 227835
rect 96475 227492 96541 227493
rect 96475 227428 96476 227492
rect 96540 227428 96541 227492
rect 96475 227427 96541 227428
rect 94404 203818 94586 204054
rect 94822 203818 95004 204054
rect 94404 203734 95004 203818
rect 94404 203498 94586 203734
rect 94822 203498 95004 203734
rect 94404 168054 95004 203498
rect 98004 207654 98604 243098
rect 98004 207418 98186 207654
rect 98422 207418 98604 207654
rect 98004 207334 98604 207418
rect 98004 207098 98186 207334
rect 98422 207098 98604 207334
rect 96475 180980 96541 180981
rect 96475 180916 96476 180980
rect 96540 180916 96541 180980
rect 96475 180915 96541 180916
rect 96478 180845 96538 180915
rect 96475 180844 96541 180845
rect 96475 180780 96476 180844
rect 96540 180780 96541 180844
rect 96475 180779 96541 180780
rect 94404 167818 94586 168054
rect 94822 167818 95004 168054
rect 94404 167734 95004 167818
rect 94404 167498 94586 167734
rect 94822 167498 95004 167734
rect 94404 132054 95004 167498
rect 94404 131818 94586 132054
rect 94822 131818 95004 132054
rect 94404 131734 95004 131818
rect 94404 131498 94586 131734
rect 94822 131498 95004 131734
rect 94404 96054 95004 131498
rect 94404 95818 94586 96054
rect 94822 95818 95004 96054
rect 94404 95734 95004 95818
rect 94404 95498 94586 95734
rect 94822 95498 95004 95734
rect 94404 60054 95004 95498
rect 94404 59818 94586 60054
rect 94822 59818 95004 60054
rect 94404 59734 95004 59818
rect 94404 59498 94586 59734
rect 94822 59498 95004 59734
rect 94404 24054 95004 59498
rect 94404 23818 94586 24054
rect 94822 23818 95004 24054
rect 94404 23734 95004 23818
rect 94404 23498 94586 23734
rect 94822 23498 95004 23734
rect 94404 -3166 95004 23498
rect 94404 -3402 94586 -3166
rect 94822 -3402 95004 -3166
rect 94404 -3486 95004 -3402
rect 94404 -3722 94586 -3486
rect 94822 -3722 95004 -3486
rect 94404 -3744 95004 -3722
rect 98004 171654 98604 207098
rect 98004 171418 98186 171654
rect 98422 171418 98604 171654
rect 98004 171334 98604 171418
rect 98004 171098 98186 171334
rect 98422 171098 98604 171334
rect 98004 135654 98604 171098
rect 98004 135418 98186 135654
rect 98422 135418 98604 135654
rect 98004 135334 98604 135418
rect 98004 135098 98186 135334
rect 98422 135098 98604 135334
rect 98004 99654 98604 135098
rect 98004 99418 98186 99654
rect 98422 99418 98604 99654
rect 98004 99334 98604 99418
rect 98004 99098 98186 99334
rect 98422 99098 98604 99334
rect 98004 63654 98604 99098
rect 98004 63418 98186 63654
rect 98422 63418 98604 63654
rect 98004 63334 98604 63418
rect 98004 63098 98186 63334
rect 98422 63098 98604 63334
rect 98004 27654 98604 63098
rect 98004 27418 98186 27654
rect 98422 27418 98604 27654
rect 98004 27334 98604 27418
rect 98004 27098 98186 27334
rect 98422 27098 98604 27334
rect 98004 -5046 98604 27098
rect 98004 -5282 98186 -5046
rect 98422 -5282 98604 -5046
rect 98004 -5366 98604 -5282
rect 98004 -5602 98186 -5366
rect 98422 -5602 98604 -5366
rect 98004 -5624 98604 -5602
rect 101604 283254 102204 317000
rect 101604 283018 101786 283254
rect 102022 283018 102204 283254
rect 101604 282934 102204 283018
rect 101604 282698 101786 282934
rect 102022 282698 102204 282934
rect 101604 247254 102204 282698
rect 108804 290454 109404 317000
rect 108804 290218 108986 290454
rect 109222 290218 109404 290454
rect 108804 290134 109404 290218
rect 108804 289898 108986 290134
rect 109222 289898 109404 290134
rect 106227 264348 106293 264349
rect 106227 264284 106228 264348
rect 106292 264284 106293 264348
rect 106227 264283 106293 264284
rect 106230 264077 106290 264283
rect 106227 264076 106293 264077
rect 106227 264012 106228 264076
rect 106292 264012 106293 264076
rect 106227 264011 106293 264012
rect 101604 247018 101786 247254
rect 102022 247018 102204 247254
rect 101604 246934 102204 247018
rect 101604 246698 101786 246934
rect 102022 246698 102204 246934
rect 101604 211254 102204 246698
rect 108804 254454 109404 289898
rect 108804 254218 108986 254454
rect 109222 254218 109404 254454
rect 108804 254134 109404 254218
rect 108804 253898 108986 254134
rect 109222 253898 109404 254134
rect 106227 228444 106293 228445
rect 106227 228380 106228 228444
rect 106292 228380 106293 228444
rect 106227 228379 106293 228380
rect 106230 228173 106290 228379
rect 106227 228172 106293 228173
rect 106227 228108 106228 228172
rect 106292 228108 106293 228172
rect 106227 228107 106293 228108
rect 101604 211018 101786 211254
rect 102022 211018 102204 211254
rect 101604 210934 102204 211018
rect 101604 210698 101786 210934
rect 102022 210698 102204 210934
rect 101604 175254 102204 210698
rect 108804 218454 109404 253898
rect 108804 218218 108986 218454
rect 109222 218218 109404 218454
rect 108804 218134 109404 218218
rect 108804 217898 108986 218134
rect 109222 217898 109404 218134
rect 108804 182454 109404 217898
rect 108804 182218 108986 182454
rect 109222 182218 109404 182454
rect 108804 182134 109404 182218
rect 108804 181898 108986 182134
rect 109222 181898 109404 182134
rect 106227 181524 106293 181525
rect 106227 181460 106228 181524
rect 106292 181460 106293 181524
rect 106227 181459 106293 181460
rect 106230 181253 106290 181459
rect 106227 181252 106293 181253
rect 106227 181188 106228 181252
rect 106292 181188 106293 181252
rect 106227 181187 106293 181188
rect 101604 175018 101786 175254
rect 102022 175018 102204 175254
rect 101604 174934 102204 175018
rect 101604 174698 101786 174934
rect 102022 174698 102204 174934
rect 101604 139254 102204 174698
rect 106227 170508 106293 170509
rect 106227 170444 106228 170508
rect 106292 170444 106293 170508
rect 106227 170443 106293 170444
rect 106230 170237 106290 170443
rect 106227 170236 106293 170237
rect 106227 170172 106228 170236
rect 106292 170172 106293 170236
rect 106227 170171 106293 170172
rect 101604 139018 101786 139254
rect 102022 139018 102204 139254
rect 101604 138934 102204 139018
rect 101604 138698 101786 138934
rect 102022 138698 102204 138934
rect 101604 103254 102204 138698
rect 101604 103018 101786 103254
rect 102022 103018 102204 103254
rect 101604 102934 102204 103018
rect 101604 102698 101786 102934
rect 102022 102698 102204 102934
rect 101604 67254 102204 102698
rect 101604 67018 101786 67254
rect 102022 67018 102204 67254
rect 101604 66934 102204 67018
rect 101604 66698 101786 66934
rect 102022 66698 102204 66934
rect 101604 31254 102204 66698
rect 101604 31018 101786 31254
rect 102022 31018 102204 31254
rect 101604 30934 102204 31018
rect 101604 30698 101786 30934
rect 102022 30698 102204 30934
rect 83604 -6222 83786 -5986
rect 84022 -6222 84204 -5986
rect 83604 -6306 84204 -6222
rect 83604 -6542 83786 -6306
rect 84022 -6542 84204 -6306
rect 83604 -7504 84204 -6542
rect 101604 -6926 102204 30698
rect 108804 146454 109404 181898
rect 108804 146218 108986 146454
rect 109222 146218 109404 146454
rect 108804 146134 109404 146218
rect 108804 145898 108986 146134
rect 109222 145898 109404 146134
rect 108804 110454 109404 145898
rect 108804 110218 108986 110454
rect 109222 110218 109404 110454
rect 108804 110134 109404 110218
rect 108804 109898 108986 110134
rect 109222 109898 109404 110134
rect 108804 74454 109404 109898
rect 108804 74218 108986 74454
rect 109222 74218 109404 74454
rect 108804 74134 109404 74218
rect 108804 73898 108986 74134
rect 109222 73898 109404 74134
rect 108804 38454 109404 73898
rect 108804 38218 108986 38454
rect 109222 38218 109404 38454
rect 108804 38134 109404 38218
rect 108804 37898 108986 38134
rect 109222 37898 109404 38134
rect 108804 2454 109404 37898
rect 108804 2218 108986 2454
rect 109222 2218 109404 2454
rect 108804 2134 109404 2218
rect 108804 1898 108986 2134
rect 109222 1898 109404 2134
rect 108804 -346 109404 1898
rect 108804 -582 108986 -346
rect 109222 -582 109404 -346
rect 108804 -666 109404 -582
rect 108804 -902 108986 -666
rect 109222 -902 109404 -666
rect 108804 -1864 109404 -902
rect 112404 294054 113004 317000
rect 112404 293818 112586 294054
rect 112822 293818 113004 294054
rect 112404 293734 113004 293818
rect 112404 293498 112586 293734
rect 112822 293498 113004 293734
rect 112404 258054 113004 293498
rect 112404 257818 112586 258054
rect 112822 257818 113004 258054
rect 112404 257734 113004 257818
rect 112404 257498 112586 257734
rect 112822 257498 113004 257734
rect 112404 222054 113004 257498
rect 112404 221818 112586 222054
rect 112822 221818 113004 222054
rect 112404 221734 113004 221818
rect 112404 221498 112586 221734
rect 112822 221498 113004 221734
rect 112404 186054 113004 221498
rect 112404 185818 112586 186054
rect 112822 185818 113004 186054
rect 112404 185734 113004 185818
rect 112404 185498 112586 185734
rect 112822 185498 113004 185734
rect 112404 150054 113004 185498
rect 112404 149818 112586 150054
rect 112822 149818 113004 150054
rect 112404 149734 113004 149818
rect 112404 149498 112586 149734
rect 112822 149498 113004 149734
rect 112404 114054 113004 149498
rect 112404 113818 112586 114054
rect 112822 113818 113004 114054
rect 112404 113734 113004 113818
rect 112404 113498 112586 113734
rect 112822 113498 113004 113734
rect 112404 78054 113004 113498
rect 112404 77818 112586 78054
rect 112822 77818 113004 78054
rect 112404 77734 113004 77818
rect 112404 77498 112586 77734
rect 112822 77498 113004 77734
rect 112404 42054 113004 77498
rect 112404 41818 112586 42054
rect 112822 41818 113004 42054
rect 112404 41734 113004 41818
rect 112404 41498 112586 41734
rect 112822 41498 113004 41734
rect 112404 6054 113004 41498
rect 112404 5818 112586 6054
rect 112822 5818 113004 6054
rect 112404 5734 113004 5818
rect 112404 5498 112586 5734
rect 112822 5498 113004 5734
rect 112404 -2226 113004 5498
rect 112404 -2462 112586 -2226
rect 112822 -2462 113004 -2226
rect 112404 -2546 113004 -2462
rect 112404 -2782 112586 -2546
rect 112822 -2782 113004 -2546
rect 112404 -3744 113004 -2782
rect 116004 297654 116604 317000
rect 116004 297418 116186 297654
rect 116422 297418 116604 297654
rect 116004 297334 116604 297418
rect 116004 297098 116186 297334
rect 116422 297098 116604 297334
rect 116004 261654 116604 297098
rect 116004 261418 116186 261654
rect 116422 261418 116604 261654
rect 116004 261334 116604 261418
rect 116004 261098 116186 261334
rect 116422 261098 116604 261334
rect 116004 225654 116604 261098
rect 116004 225418 116186 225654
rect 116422 225418 116604 225654
rect 116004 225334 116604 225418
rect 116004 225098 116186 225334
rect 116422 225098 116604 225334
rect 116004 189654 116604 225098
rect 116004 189418 116186 189654
rect 116422 189418 116604 189654
rect 116004 189334 116604 189418
rect 116004 189098 116186 189334
rect 116422 189098 116604 189334
rect 116004 153654 116604 189098
rect 116004 153418 116186 153654
rect 116422 153418 116604 153654
rect 116004 153334 116604 153418
rect 116004 153098 116186 153334
rect 116422 153098 116604 153334
rect 116004 117654 116604 153098
rect 116004 117418 116186 117654
rect 116422 117418 116604 117654
rect 116004 117334 116604 117418
rect 116004 117098 116186 117334
rect 116422 117098 116604 117334
rect 116004 81654 116604 117098
rect 116004 81418 116186 81654
rect 116422 81418 116604 81654
rect 116004 81334 116604 81418
rect 116004 81098 116186 81334
rect 116422 81098 116604 81334
rect 116004 45654 116604 81098
rect 116004 45418 116186 45654
rect 116422 45418 116604 45654
rect 116004 45334 116604 45418
rect 116004 45098 116186 45334
rect 116422 45098 116604 45334
rect 116004 9654 116604 45098
rect 116004 9418 116186 9654
rect 116422 9418 116604 9654
rect 116004 9334 116604 9418
rect 116004 9098 116186 9334
rect 116422 9098 116604 9334
rect 116004 -4106 116604 9098
rect 116004 -4342 116186 -4106
rect 116422 -4342 116604 -4106
rect 116004 -4426 116604 -4342
rect 116004 -4662 116186 -4426
rect 116422 -4662 116604 -4426
rect 116004 -5624 116604 -4662
rect 119604 301254 120204 317000
rect 119604 301018 119786 301254
rect 120022 301018 120204 301254
rect 119604 300934 120204 301018
rect 119604 300698 119786 300934
rect 120022 300698 120204 300934
rect 119604 265254 120204 300698
rect 119604 265018 119786 265254
rect 120022 265018 120204 265254
rect 119604 264934 120204 265018
rect 119604 264698 119786 264934
rect 120022 264698 120204 264934
rect 119604 229254 120204 264698
rect 126804 308454 127404 317000
rect 126804 308218 126986 308454
rect 127222 308218 127404 308454
rect 126804 308134 127404 308218
rect 126804 307898 126986 308134
rect 127222 307898 127404 308134
rect 126804 272454 127404 307898
rect 126804 272218 126986 272454
rect 127222 272218 127404 272454
rect 126804 272134 127404 272218
rect 126804 271898 126986 272134
rect 127222 271898 127404 272134
rect 125547 264212 125613 264213
rect 125547 264148 125548 264212
rect 125612 264148 125613 264212
rect 125547 264147 125613 264148
rect 125550 263941 125610 264147
rect 125547 263940 125613 263941
rect 125547 263876 125548 263940
rect 125612 263876 125613 263940
rect 125547 263875 125613 263876
rect 119604 229018 119786 229254
rect 120022 229018 120204 229254
rect 119604 228934 120204 229018
rect 119604 228698 119786 228934
rect 120022 228698 120204 228934
rect 119604 193254 120204 228698
rect 126804 236454 127404 271898
rect 126804 236218 126986 236454
rect 127222 236218 127404 236454
rect 126804 236134 127404 236218
rect 126804 235898 126986 236134
rect 127222 235898 127404 236134
rect 125547 228308 125613 228309
rect 125547 228244 125548 228308
rect 125612 228244 125613 228308
rect 125547 228243 125613 228244
rect 125550 228037 125610 228243
rect 125547 228036 125613 228037
rect 125547 227972 125548 228036
rect 125612 227972 125613 228036
rect 125547 227971 125613 227972
rect 125547 217292 125613 217293
rect 125547 217228 125548 217292
rect 125612 217228 125613 217292
rect 125547 217227 125613 217228
rect 125550 217021 125610 217227
rect 125547 217020 125613 217021
rect 125547 216956 125548 217020
rect 125612 216956 125613 217020
rect 125547 216955 125613 216956
rect 119604 193018 119786 193254
rect 120022 193018 120204 193254
rect 119604 192934 120204 193018
rect 119604 192698 119786 192934
rect 120022 192698 120204 192934
rect 119604 157254 120204 192698
rect 126804 200454 127404 235898
rect 126804 200218 126986 200454
rect 127222 200218 127404 200454
rect 126804 200134 127404 200218
rect 126804 199898 126986 200134
rect 127222 199898 127404 200134
rect 125547 170372 125613 170373
rect 125547 170308 125548 170372
rect 125612 170308 125613 170372
rect 125547 170307 125613 170308
rect 125550 170101 125610 170307
rect 125547 170100 125613 170101
rect 125547 170036 125548 170100
rect 125612 170036 125613 170100
rect 125547 170035 125613 170036
rect 119604 157018 119786 157254
rect 120022 157018 120204 157254
rect 119604 156934 120204 157018
rect 119604 156698 119786 156934
rect 120022 156698 120204 156934
rect 119604 121254 120204 156698
rect 119604 121018 119786 121254
rect 120022 121018 120204 121254
rect 119604 120934 120204 121018
rect 119604 120698 119786 120934
rect 120022 120698 120204 120934
rect 119604 85254 120204 120698
rect 119604 85018 119786 85254
rect 120022 85018 120204 85254
rect 119604 84934 120204 85018
rect 119604 84698 119786 84934
rect 120022 84698 120204 84934
rect 119604 49254 120204 84698
rect 126804 164454 127404 199898
rect 126804 164218 126986 164454
rect 127222 164218 127404 164454
rect 126804 164134 127404 164218
rect 126804 163898 126986 164134
rect 127222 163898 127404 164134
rect 126804 128454 127404 163898
rect 126804 128218 126986 128454
rect 127222 128218 127404 128454
rect 126804 128134 127404 128218
rect 126804 127898 126986 128134
rect 127222 127898 127404 128134
rect 126804 92454 127404 127898
rect 126804 92218 126986 92454
rect 127222 92218 127404 92454
rect 126804 92134 127404 92218
rect 126804 91898 126986 92134
rect 127222 91898 127404 92134
rect 125547 76532 125613 76533
rect 125547 76468 125548 76532
rect 125612 76468 125613 76532
rect 125547 76467 125613 76468
rect 125550 76261 125610 76467
rect 125547 76260 125613 76261
rect 125547 76196 125548 76260
rect 125612 76196 125613 76260
rect 125547 76195 125613 76196
rect 119604 49018 119786 49254
rect 120022 49018 120204 49254
rect 119604 48934 120204 49018
rect 119604 48698 119786 48934
rect 120022 48698 120204 48934
rect 119604 13254 120204 48698
rect 119604 13018 119786 13254
rect 120022 13018 120204 13254
rect 119604 12934 120204 13018
rect 119604 12698 119786 12934
rect 120022 12698 120204 12934
rect 101604 -7162 101786 -6926
rect 102022 -7162 102204 -6926
rect 101604 -7246 102204 -7162
rect 101604 -7482 101786 -7246
rect 102022 -7482 102204 -7246
rect 101604 -7504 102204 -7482
rect 119604 -5986 120204 12698
rect 126804 56454 127404 91898
rect 126804 56218 126986 56454
rect 127222 56218 127404 56454
rect 126804 56134 127404 56218
rect 126804 55898 126986 56134
rect 127222 55898 127404 56134
rect 126804 20454 127404 55898
rect 126804 20218 126986 20454
rect 127222 20218 127404 20454
rect 126804 20134 127404 20218
rect 126804 19898 126986 20134
rect 127222 19898 127404 20134
rect 126804 -1286 127404 19898
rect 126804 -1522 126986 -1286
rect 127222 -1522 127404 -1286
rect 126804 -1606 127404 -1522
rect 126804 -1842 126986 -1606
rect 127222 -1842 127404 -1606
rect 126804 -1864 127404 -1842
rect 130404 312054 131004 317000
rect 130404 311818 130586 312054
rect 130822 311818 131004 312054
rect 130404 311734 131004 311818
rect 130404 311498 130586 311734
rect 130822 311498 131004 311734
rect 130404 276054 131004 311498
rect 130404 275818 130586 276054
rect 130822 275818 131004 276054
rect 130404 275734 131004 275818
rect 130404 275498 130586 275734
rect 130822 275498 131004 275734
rect 130404 240054 131004 275498
rect 130404 239818 130586 240054
rect 130822 239818 131004 240054
rect 130404 239734 131004 239818
rect 130404 239498 130586 239734
rect 130822 239498 131004 239734
rect 130404 204054 131004 239498
rect 130404 203818 130586 204054
rect 130822 203818 131004 204054
rect 130404 203734 131004 203818
rect 130404 203498 130586 203734
rect 130822 203498 131004 203734
rect 130404 168054 131004 203498
rect 130404 167818 130586 168054
rect 130822 167818 131004 168054
rect 130404 167734 131004 167818
rect 130404 167498 130586 167734
rect 130822 167498 131004 167734
rect 130404 132054 131004 167498
rect 130404 131818 130586 132054
rect 130822 131818 131004 132054
rect 130404 131734 131004 131818
rect 130404 131498 130586 131734
rect 130822 131498 131004 131734
rect 130404 96054 131004 131498
rect 130404 95818 130586 96054
rect 130822 95818 131004 96054
rect 130404 95734 131004 95818
rect 130404 95498 130586 95734
rect 130822 95498 131004 95734
rect 130404 60054 131004 95498
rect 130404 59818 130586 60054
rect 130822 59818 131004 60054
rect 130404 59734 131004 59818
rect 130404 59498 130586 59734
rect 130822 59498 131004 59734
rect 130404 24054 131004 59498
rect 130404 23818 130586 24054
rect 130822 23818 131004 24054
rect 130404 23734 131004 23818
rect 130404 23498 130586 23734
rect 130822 23498 131004 23734
rect 130404 -3166 131004 23498
rect 130404 -3402 130586 -3166
rect 130822 -3402 131004 -3166
rect 130404 -3486 131004 -3402
rect 130404 -3722 130586 -3486
rect 130822 -3722 131004 -3486
rect 130404 -3744 131004 -3722
rect 134004 315654 134604 317000
rect 134004 315418 134186 315654
rect 134422 315418 134604 315654
rect 134004 315334 134604 315418
rect 134004 315098 134186 315334
rect 134422 315098 134604 315334
rect 134004 279654 134604 315098
rect 134004 279418 134186 279654
rect 134422 279418 134604 279654
rect 134004 279334 134604 279418
rect 134004 279098 134186 279334
rect 134422 279098 134604 279334
rect 134004 243654 134604 279098
rect 134004 243418 134186 243654
rect 134422 243418 134604 243654
rect 134004 243334 134604 243418
rect 134004 243098 134186 243334
rect 134422 243098 134604 243334
rect 134004 207654 134604 243098
rect 134004 207418 134186 207654
rect 134422 207418 134604 207654
rect 134004 207334 134604 207418
rect 134004 207098 134186 207334
rect 134422 207098 134604 207334
rect 134004 171654 134604 207098
rect 134004 171418 134186 171654
rect 134422 171418 134604 171654
rect 134004 171334 134604 171418
rect 134004 171098 134186 171334
rect 134422 171098 134604 171334
rect 134004 135654 134604 171098
rect 134004 135418 134186 135654
rect 134422 135418 134604 135654
rect 134004 135334 134604 135418
rect 134004 135098 134186 135334
rect 134422 135098 134604 135334
rect 134004 99654 134604 135098
rect 134004 99418 134186 99654
rect 134422 99418 134604 99654
rect 134004 99334 134604 99418
rect 134004 99098 134186 99334
rect 134422 99098 134604 99334
rect 134004 63654 134604 99098
rect 134004 63418 134186 63654
rect 134422 63418 134604 63654
rect 134004 63334 134604 63418
rect 134004 63098 134186 63334
rect 134422 63098 134604 63334
rect 134004 27654 134604 63098
rect 134004 27418 134186 27654
rect 134422 27418 134604 27654
rect 134004 27334 134604 27418
rect 134004 27098 134186 27334
rect 134422 27098 134604 27334
rect 134004 -5046 134604 27098
rect 134004 -5282 134186 -5046
rect 134422 -5282 134604 -5046
rect 134004 -5366 134604 -5282
rect 134004 -5602 134186 -5366
rect 134422 -5602 134604 -5366
rect 134004 -5624 134604 -5602
rect 137604 283254 138204 317000
rect 137604 283018 137786 283254
rect 138022 283018 138204 283254
rect 137604 282934 138204 283018
rect 137604 282698 137786 282934
rect 138022 282698 138204 282934
rect 137604 247254 138204 282698
rect 137604 247018 137786 247254
rect 138022 247018 138204 247254
rect 137604 246934 138204 247018
rect 137604 246698 137786 246934
rect 138022 246698 138204 246934
rect 137604 211254 138204 246698
rect 137604 211018 137786 211254
rect 138022 211018 138204 211254
rect 137604 210934 138204 211018
rect 137604 210698 137786 210934
rect 138022 210698 138204 210934
rect 137604 175254 138204 210698
rect 137604 175018 137786 175254
rect 138022 175018 138204 175254
rect 137604 174934 138204 175018
rect 137604 174698 137786 174934
rect 138022 174698 138204 174934
rect 137604 139254 138204 174698
rect 137604 139018 137786 139254
rect 138022 139018 138204 139254
rect 137604 138934 138204 139018
rect 137604 138698 137786 138934
rect 138022 138698 138204 138934
rect 137604 103254 138204 138698
rect 137604 103018 137786 103254
rect 138022 103018 138204 103254
rect 137604 102934 138204 103018
rect 137604 102698 137786 102934
rect 138022 102698 138204 102934
rect 137604 67254 138204 102698
rect 137604 67018 137786 67254
rect 138022 67018 138204 67254
rect 137604 66934 138204 67018
rect 137604 66698 137786 66934
rect 138022 66698 138204 66934
rect 137604 31254 138204 66698
rect 137604 31018 137786 31254
rect 138022 31018 138204 31254
rect 137604 30934 138204 31018
rect 137604 30698 137786 30934
rect 138022 30698 138204 30934
rect 119604 -6222 119786 -5986
rect 120022 -6222 120204 -5986
rect 119604 -6306 120204 -6222
rect 119604 -6542 119786 -6306
rect 120022 -6542 120204 -6306
rect 119604 -7504 120204 -6542
rect 137604 -6926 138204 30698
rect 144804 290454 145404 317000
rect 144804 290218 144986 290454
rect 145222 290218 145404 290454
rect 144804 290134 145404 290218
rect 144804 289898 144986 290134
rect 145222 289898 145404 290134
rect 144804 254454 145404 289898
rect 144804 254218 144986 254454
rect 145222 254218 145404 254454
rect 144804 254134 145404 254218
rect 144804 253898 144986 254134
rect 145222 253898 145404 254134
rect 144804 218454 145404 253898
rect 144804 218218 144986 218454
rect 145222 218218 145404 218454
rect 144804 218134 145404 218218
rect 144804 217898 144986 218134
rect 145222 217898 145404 218134
rect 144804 182454 145404 217898
rect 144804 182218 144986 182454
rect 145222 182218 145404 182454
rect 144804 182134 145404 182218
rect 144804 181898 144986 182134
rect 145222 181898 145404 182134
rect 144804 146454 145404 181898
rect 144804 146218 144986 146454
rect 145222 146218 145404 146454
rect 144804 146134 145404 146218
rect 144804 145898 144986 146134
rect 145222 145898 145404 146134
rect 144804 110454 145404 145898
rect 144804 110218 144986 110454
rect 145222 110218 145404 110454
rect 144804 110134 145404 110218
rect 144804 109898 144986 110134
rect 145222 109898 145404 110134
rect 144804 74454 145404 109898
rect 144804 74218 144986 74454
rect 145222 74218 145404 74454
rect 144804 74134 145404 74218
rect 144804 73898 144986 74134
rect 145222 73898 145404 74134
rect 144804 38454 145404 73898
rect 144804 38218 144986 38454
rect 145222 38218 145404 38454
rect 144804 38134 145404 38218
rect 144804 37898 144986 38134
rect 145222 37898 145404 38134
rect 144804 2454 145404 37898
rect 144804 2218 144986 2454
rect 145222 2218 145404 2454
rect 144804 2134 145404 2218
rect 144804 1898 144986 2134
rect 145222 1898 145404 2134
rect 144804 -346 145404 1898
rect 144804 -582 144986 -346
rect 145222 -582 145404 -346
rect 144804 -666 145404 -582
rect 144804 -902 144986 -666
rect 145222 -902 145404 -666
rect 144804 -1864 145404 -902
rect 148404 294054 149004 317000
rect 148404 293818 148586 294054
rect 148822 293818 149004 294054
rect 148404 293734 149004 293818
rect 148404 293498 148586 293734
rect 148822 293498 149004 293734
rect 148404 258054 149004 293498
rect 148404 257818 148586 258054
rect 148822 257818 149004 258054
rect 148404 257734 149004 257818
rect 148404 257498 148586 257734
rect 148822 257498 149004 257734
rect 148404 222054 149004 257498
rect 148404 221818 148586 222054
rect 148822 221818 149004 222054
rect 148404 221734 149004 221818
rect 148404 221498 148586 221734
rect 148822 221498 149004 221734
rect 148404 186054 149004 221498
rect 148404 185818 148586 186054
rect 148822 185818 149004 186054
rect 148404 185734 149004 185818
rect 148404 185498 148586 185734
rect 148822 185498 149004 185734
rect 148404 150054 149004 185498
rect 148404 149818 148586 150054
rect 148822 149818 149004 150054
rect 148404 149734 149004 149818
rect 148404 149498 148586 149734
rect 148822 149498 149004 149734
rect 148404 114054 149004 149498
rect 148404 113818 148586 114054
rect 148822 113818 149004 114054
rect 148404 113734 149004 113818
rect 148404 113498 148586 113734
rect 148822 113498 149004 113734
rect 148404 78054 149004 113498
rect 148404 77818 148586 78054
rect 148822 77818 149004 78054
rect 148404 77734 149004 77818
rect 148404 77498 148586 77734
rect 148822 77498 149004 77734
rect 148404 42054 149004 77498
rect 148404 41818 148586 42054
rect 148822 41818 149004 42054
rect 148404 41734 149004 41818
rect 148404 41498 148586 41734
rect 148822 41498 149004 41734
rect 148404 6054 149004 41498
rect 148404 5818 148586 6054
rect 148822 5818 149004 6054
rect 148404 5734 149004 5818
rect 148404 5498 148586 5734
rect 148822 5498 149004 5734
rect 148404 -2226 149004 5498
rect 148404 -2462 148586 -2226
rect 148822 -2462 149004 -2226
rect 148404 -2546 149004 -2462
rect 148404 -2782 148586 -2546
rect 148822 -2782 149004 -2546
rect 148404 -3744 149004 -2782
rect 152004 297654 152604 317000
rect 152004 297418 152186 297654
rect 152422 297418 152604 297654
rect 152004 297334 152604 297418
rect 152004 297098 152186 297334
rect 152422 297098 152604 297334
rect 152004 261654 152604 297098
rect 152004 261418 152186 261654
rect 152422 261418 152604 261654
rect 152004 261334 152604 261418
rect 152004 261098 152186 261334
rect 152422 261098 152604 261334
rect 152004 225654 152604 261098
rect 152004 225418 152186 225654
rect 152422 225418 152604 225654
rect 152004 225334 152604 225418
rect 152004 225098 152186 225334
rect 152422 225098 152604 225334
rect 152004 189654 152604 225098
rect 152004 189418 152186 189654
rect 152422 189418 152604 189654
rect 152004 189334 152604 189418
rect 152004 189098 152186 189334
rect 152422 189098 152604 189334
rect 152004 153654 152604 189098
rect 152004 153418 152186 153654
rect 152422 153418 152604 153654
rect 152004 153334 152604 153418
rect 152004 153098 152186 153334
rect 152422 153098 152604 153334
rect 152004 117654 152604 153098
rect 152004 117418 152186 117654
rect 152422 117418 152604 117654
rect 152004 117334 152604 117418
rect 152004 117098 152186 117334
rect 152422 117098 152604 117334
rect 152004 81654 152604 117098
rect 152004 81418 152186 81654
rect 152422 81418 152604 81654
rect 152004 81334 152604 81418
rect 152004 81098 152186 81334
rect 152422 81098 152604 81334
rect 152004 45654 152604 81098
rect 152004 45418 152186 45654
rect 152422 45418 152604 45654
rect 152004 45334 152604 45418
rect 152004 45098 152186 45334
rect 152422 45098 152604 45334
rect 152004 9654 152604 45098
rect 152004 9418 152186 9654
rect 152422 9418 152604 9654
rect 152004 9334 152604 9418
rect 152004 9098 152186 9334
rect 152422 9098 152604 9334
rect 152004 -4106 152604 9098
rect 152004 -4342 152186 -4106
rect 152422 -4342 152604 -4106
rect 152004 -4426 152604 -4342
rect 152004 -4662 152186 -4426
rect 152422 -4662 152604 -4426
rect 152004 -5624 152604 -4662
rect 155604 301254 156204 317000
rect 155604 301018 155786 301254
rect 156022 301018 156204 301254
rect 155604 300934 156204 301018
rect 155604 300698 155786 300934
rect 156022 300698 156204 300934
rect 155604 265254 156204 300698
rect 155604 265018 155786 265254
rect 156022 265018 156204 265254
rect 155604 264934 156204 265018
rect 155604 264698 155786 264934
rect 156022 264698 156204 264934
rect 155604 229254 156204 264698
rect 155604 229018 155786 229254
rect 156022 229018 156204 229254
rect 155604 228934 156204 229018
rect 155604 228698 155786 228934
rect 156022 228698 156204 228934
rect 155604 193254 156204 228698
rect 155604 193018 155786 193254
rect 156022 193018 156204 193254
rect 155604 192934 156204 193018
rect 155604 192698 155786 192934
rect 156022 192698 156204 192934
rect 155604 157254 156204 192698
rect 155604 157018 155786 157254
rect 156022 157018 156204 157254
rect 155604 156934 156204 157018
rect 155604 156698 155786 156934
rect 156022 156698 156204 156934
rect 155604 121254 156204 156698
rect 155604 121018 155786 121254
rect 156022 121018 156204 121254
rect 155604 120934 156204 121018
rect 155604 120698 155786 120934
rect 156022 120698 156204 120934
rect 155604 85254 156204 120698
rect 155604 85018 155786 85254
rect 156022 85018 156204 85254
rect 155604 84934 156204 85018
rect 155604 84698 155786 84934
rect 156022 84698 156204 84934
rect 155604 49254 156204 84698
rect 155604 49018 155786 49254
rect 156022 49018 156204 49254
rect 155604 48934 156204 49018
rect 155604 48698 155786 48934
rect 156022 48698 156204 48934
rect 155604 13254 156204 48698
rect 155604 13018 155786 13254
rect 156022 13018 156204 13254
rect 155604 12934 156204 13018
rect 155604 12698 155786 12934
rect 156022 12698 156204 12934
rect 137604 -7162 137786 -6926
rect 138022 -7162 138204 -6926
rect 137604 -7246 138204 -7162
rect 137604 -7482 137786 -7246
rect 138022 -7482 138204 -7246
rect 137604 -7504 138204 -7482
rect 155604 -5986 156204 12698
rect 162804 308454 163404 317000
rect 162804 308218 162986 308454
rect 163222 308218 163404 308454
rect 162804 308134 163404 308218
rect 162804 307898 162986 308134
rect 163222 307898 163404 308134
rect 162804 272454 163404 307898
rect 162804 272218 162986 272454
rect 163222 272218 163404 272454
rect 162804 272134 163404 272218
rect 162804 271898 162986 272134
rect 163222 271898 163404 272134
rect 162804 236454 163404 271898
rect 162804 236218 162986 236454
rect 163222 236218 163404 236454
rect 162804 236134 163404 236218
rect 162804 235898 162986 236134
rect 163222 235898 163404 236134
rect 162804 200454 163404 235898
rect 162804 200218 162986 200454
rect 163222 200218 163404 200454
rect 162804 200134 163404 200218
rect 162804 199898 162986 200134
rect 163222 199898 163404 200134
rect 162804 164454 163404 199898
rect 162804 164218 162986 164454
rect 163222 164218 163404 164454
rect 162804 164134 163404 164218
rect 162804 163898 162986 164134
rect 163222 163898 163404 164134
rect 162804 128454 163404 163898
rect 162804 128218 162986 128454
rect 163222 128218 163404 128454
rect 162804 128134 163404 128218
rect 162804 127898 162986 128134
rect 163222 127898 163404 128134
rect 162804 92454 163404 127898
rect 162804 92218 162986 92454
rect 163222 92218 163404 92454
rect 162804 92134 163404 92218
rect 162804 91898 162986 92134
rect 163222 91898 163404 92134
rect 162804 56454 163404 91898
rect 162804 56218 162986 56454
rect 163222 56218 163404 56454
rect 162804 56134 163404 56218
rect 162804 55898 162986 56134
rect 163222 55898 163404 56134
rect 162804 20454 163404 55898
rect 162804 20218 162986 20454
rect 163222 20218 163404 20454
rect 162804 20134 163404 20218
rect 162804 19898 162986 20134
rect 163222 19898 163404 20134
rect 162804 -1286 163404 19898
rect 162804 -1522 162986 -1286
rect 163222 -1522 163404 -1286
rect 162804 -1606 163404 -1522
rect 162804 -1842 162986 -1606
rect 163222 -1842 163404 -1606
rect 162804 -1864 163404 -1842
rect 166404 312054 167004 317000
rect 166404 311818 166586 312054
rect 166822 311818 167004 312054
rect 166404 311734 167004 311818
rect 166404 311498 166586 311734
rect 166822 311498 167004 311734
rect 166404 276054 167004 311498
rect 166404 275818 166586 276054
rect 166822 275818 167004 276054
rect 166404 275734 167004 275818
rect 166404 275498 166586 275734
rect 166822 275498 167004 275734
rect 166404 240054 167004 275498
rect 166404 239818 166586 240054
rect 166822 239818 167004 240054
rect 166404 239734 167004 239818
rect 166404 239498 166586 239734
rect 166822 239498 167004 239734
rect 166404 204054 167004 239498
rect 166404 203818 166586 204054
rect 166822 203818 167004 204054
rect 166404 203734 167004 203818
rect 166404 203498 166586 203734
rect 166822 203498 167004 203734
rect 166404 168054 167004 203498
rect 166404 167818 166586 168054
rect 166822 167818 167004 168054
rect 166404 167734 167004 167818
rect 166404 167498 166586 167734
rect 166822 167498 167004 167734
rect 166404 132054 167004 167498
rect 166404 131818 166586 132054
rect 166822 131818 167004 132054
rect 166404 131734 167004 131818
rect 166404 131498 166586 131734
rect 166822 131498 167004 131734
rect 166404 96054 167004 131498
rect 166404 95818 166586 96054
rect 166822 95818 167004 96054
rect 166404 95734 167004 95818
rect 166404 95498 166586 95734
rect 166822 95498 167004 95734
rect 166404 60054 167004 95498
rect 166404 59818 166586 60054
rect 166822 59818 167004 60054
rect 166404 59734 167004 59818
rect 166404 59498 166586 59734
rect 166822 59498 167004 59734
rect 166404 24054 167004 59498
rect 166404 23818 166586 24054
rect 166822 23818 167004 24054
rect 166404 23734 167004 23818
rect 166404 23498 166586 23734
rect 166822 23498 167004 23734
rect 166404 -3166 167004 23498
rect 166404 -3402 166586 -3166
rect 166822 -3402 167004 -3166
rect 166404 -3486 167004 -3402
rect 166404 -3722 166586 -3486
rect 166822 -3722 167004 -3486
rect 166404 -3744 167004 -3722
rect 170004 315654 170604 317000
rect 170004 315418 170186 315654
rect 170422 315418 170604 315654
rect 170004 315334 170604 315418
rect 170004 315098 170186 315334
rect 170422 315098 170604 315334
rect 170004 279654 170604 315098
rect 170004 279418 170186 279654
rect 170422 279418 170604 279654
rect 170004 279334 170604 279418
rect 170004 279098 170186 279334
rect 170422 279098 170604 279334
rect 170004 243654 170604 279098
rect 170004 243418 170186 243654
rect 170422 243418 170604 243654
rect 170004 243334 170604 243418
rect 170004 243098 170186 243334
rect 170422 243098 170604 243334
rect 170004 207654 170604 243098
rect 170004 207418 170186 207654
rect 170422 207418 170604 207654
rect 170004 207334 170604 207418
rect 170004 207098 170186 207334
rect 170422 207098 170604 207334
rect 170004 171654 170604 207098
rect 170004 171418 170186 171654
rect 170422 171418 170604 171654
rect 170004 171334 170604 171418
rect 170004 171098 170186 171334
rect 170422 171098 170604 171334
rect 170004 135654 170604 171098
rect 170004 135418 170186 135654
rect 170422 135418 170604 135654
rect 170004 135334 170604 135418
rect 170004 135098 170186 135334
rect 170422 135098 170604 135334
rect 170004 99654 170604 135098
rect 170004 99418 170186 99654
rect 170422 99418 170604 99654
rect 170004 99334 170604 99418
rect 170004 99098 170186 99334
rect 170422 99098 170604 99334
rect 170004 63654 170604 99098
rect 170004 63418 170186 63654
rect 170422 63418 170604 63654
rect 170004 63334 170604 63418
rect 170004 63098 170186 63334
rect 170422 63098 170604 63334
rect 170004 27654 170604 63098
rect 170004 27418 170186 27654
rect 170422 27418 170604 27654
rect 170004 27334 170604 27418
rect 170004 27098 170186 27334
rect 170422 27098 170604 27334
rect 170004 -5046 170604 27098
rect 170004 -5282 170186 -5046
rect 170422 -5282 170604 -5046
rect 170004 -5366 170604 -5282
rect 170004 -5602 170186 -5366
rect 170422 -5602 170604 -5366
rect 170004 -5624 170604 -5602
rect 173604 283254 174204 317000
rect 173604 283018 173786 283254
rect 174022 283018 174204 283254
rect 173604 282934 174204 283018
rect 173604 282698 173786 282934
rect 174022 282698 174204 282934
rect 173604 247254 174204 282698
rect 173604 247018 173786 247254
rect 174022 247018 174204 247254
rect 173604 246934 174204 247018
rect 173604 246698 173786 246934
rect 174022 246698 174204 246934
rect 173604 211254 174204 246698
rect 173604 211018 173786 211254
rect 174022 211018 174204 211254
rect 173604 210934 174204 211018
rect 173604 210698 173786 210934
rect 174022 210698 174204 210934
rect 173604 175254 174204 210698
rect 173604 175018 173786 175254
rect 174022 175018 174204 175254
rect 173604 174934 174204 175018
rect 173604 174698 173786 174934
rect 174022 174698 174204 174934
rect 173604 139254 174204 174698
rect 173604 139018 173786 139254
rect 174022 139018 174204 139254
rect 173604 138934 174204 139018
rect 173604 138698 173786 138934
rect 174022 138698 174204 138934
rect 173604 103254 174204 138698
rect 173604 103018 173786 103254
rect 174022 103018 174204 103254
rect 173604 102934 174204 103018
rect 173604 102698 173786 102934
rect 174022 102698 174204 102934
rect 173604 67254 174204 102698
rect 173604 67018 173786 67254
rect 174022 67018 174204 67254
rect 173604 66934 174204 67018
rect 173604 66698 173786 66934
rect 174022 66698 174204 66934
rect 173604 31254 174204 66698
rect 173604 31018 173786 31254
rect 174022 31018 174204 31254
rect 173604 30934 174204 31018
rect 173604 30698 173786 30934
rect 174022 30698 174204 30934
rect 155604 -6222 155786 -5986
rect 156022 -6222 156204 -5986
rect 155604 -6306 156204 -6222
rect 155604 -6542 155786 -6306
rect 156022 -6542 156204 -6306
rect 155604 -7504 156204 -6542
rect 173604 -6926 174204 30698
rect 180804 290454 181404 317000
rect 180804 290218 180986 290454
rect 181222 290218 181404 290454
rect 180804 290134 181404 290218
rect 180804 289898 180986 290134
rect 181222 289898 181404 290134
rect 180804 254454 181404 289898
rect 180804 254218 180986 254454
rect 181222 254218 181404 254454
rect 180804 254134 181404 254218
rect 180804 253898 180986 254134
rect 181222 253898 181404 254134
rect 180804 218454 181404 253898
rect 180804 218218 180986 218454
rect 181222 218218 181404 218454
rect 180804 218134 181404 218218
rect 180804 217898 180986 218134
rect 181222 217898 181404 218134
rect 180804 182454 181404 217898
rect 180804 182218 180986 182454
rect 181222 182218 181404 182454
rect 180804 182134 181404 182218
rect 180804 181898 180986 182134
rect 181222 181898 181404 182134
rect 180804 146454 181404 181898
rect 180804 146218 180986 146454
rect 181222 146218 181404 146454
rect 180804 146134 181404 146218
rect 180804 145898 180986 146134
rect 181222 145898 181404 146134
rect 180804 110454 181404 145898
rect 180804 110218 180986 110454
rect 181222 110218 181404 110454
rect 180804 110134 181404 110218
rect 180804 109898 180986 110134
rect 181222 109898 181404 110134
rect 180804 74454 181404 109898
rect 180804 74218 180986 74454
rect 181222 74218 181404 74454
rect 180804 74134 181404 74218
rect 180804 73898 180986 74134
rect 181222 73898 181404 74134
rect 180804 38454 181404 73898
rect 180804 38218 180986 38454
rect 181222 38218 181404 38454
rect 180804 38134 181404 38218
rect 180804 37898 180986 38134
rect 181222 37898 181404 38134
rect 180804 2454 181404 37898
rect 180804 2218 180986 2454
rect 181222 2218 181404 2454
rect 180804 2134 181404 2218
rect 180804 1898 180986 2134
rect 181222 1898 181404 2134
rect 180804 -346 181404 1898
rect 180804 -582 180986 -346
rect 181222 -582 181404 -346
rect 180804 -666 181404 -582
rect 180804 -902 180986 -666
rect 181222 -902 181404 -666
rect 180804 -1864 181404 -902
rect 184404 294054 185004 317000
rect 184404 293818 184586 294054
rect 184822 293818 185004 294054
rect 184404 293734 185004 293818
rect 184404 293498 184586 293734
rect 184822 293498 185004 293734
rect 184404 258054 185004 293498
rect 184404 257818 184586 258054
rect 184822 257818 185004 258054
rect 184404 257734 185004 257818
rect 184404 257498 184586 257734
rect 184822 257498 185004 257734
rect 184404 222054 185004 257498
rect 184404 221818 184586 222054
rect 184822 221818 185004 222054
rect 184404 221734 185004 221818
rect 184404 221498 184586 221734
rect 184822 221498 185004 221734
rect 184404 186054 185004 221498
rect 184404 185818 184586 186054
rect 184822 185818 185004 186054
rect 184404 185734 185004 185818
rect 184404 185498 184586 185734
rect 184822 185498 185004 185734
rect 184404 150054 185004 185498
rect 184404 149818 184586 150054
rect 184822 149818 185004 150054
rect 184404 149734 185004 149818
rect 184404 149498 184586 149734
rect 184822 149498 185004 149734
rect 184404 114054 185004 149498
rect 184404 113818 184586 114054
rect 184822 113818 185004 114054
rect 184404 113734 185004 113818
rect 184404 113498 184586 113734
rect 184822 113498 185004 113734
rect 184404 78054 185004 113498
rect 184404 77818 184586 78054
rect 184822 77818 185004 78054
rect 184404 77734 185004 77818
rect 184404 77498 184586 77734
rect 184822 77498 185004 77734
rect 184404 42054 185004 77498
rect 184404 41818 184586 42054
rect 184822 41818 185004 42054
rect 184404 41734 185004 41818
rect 184404 41498 184586 41734
rect 184822 41498 185004 41734
rect 184404 6054 185004 41498
rect 184404 5818 184586 6054
rect 184822 5818 185004 6054
rect 184404 5734 185004 5818
rect 184404 5498 184586 5734
rect 184822 5498 185004 5734
rect 184404 -2226 185004 5498
rect 184404 -2462 184586 -2226
rect 184822 -2462 185004 -2226
rect 184404 -2546 185004 -2462
rect 184404 -2782 184586 -2546
rect 184822 -2782 185004 -2546
rect 184404 -3744 185004 -2782
rect 188004 297654 188604 317000
rect 188004 297418 188186 297654
rect 188422 297418 188604 297654
rect 188004 297334 188604 297418
rect 188004 297098 188186 297334
rect 188422 297098 188604 297334
rect 188004 261654 188604 297098
rect 188004 261418 188186 261654
rect 188422 261418 188604 261654
rect 188004 261334 188604 261418
rect 188004 261098 188186 261334
rect 188422 261098 188604 261334
rect 188004 225654 188604 261098
rect 188004 225418 188186 225654
rect 188422 225418 188604 225654
rect 188004 225334 188604 225418
rect 188004 225098 188186 225334
rect 188422 225098 188604 225334
rect 188004 189654 188604 225098
rect 188004 189418 188186 189654
rect 188422 189418 188604 189654
rect 188004 189334 188604 189418
rect 188004 189098 188186 189334
rect 188422 189098 188604 189334
rect 188004 153654 188604 189098
rect 188004 153418 188186 153654
rect 188422 153418 188604 153654
rect 188004 153334 188604 153418
rect 188004 153098 188186 153334
rect 188422 153098 188604 153334
rect 188004 117654 188604 153098
rect 188004 117418 188186 117654
rect 188422 117418 188604 117654
rect 188004 117334 188604 117418
rect 188004 117098 188186 117334
rect 188422 117098 188604 117334
rect 188004 81654 188604 117098
rect 188004 81418 188186 81654
rect 188422 81418 188604 81654
rect 188004 81334 188604 81418
rect 188004 81098 188186 81334
rect 188422 81098 188604 81334
rect 188004 45654 188604 81098
rect 188004 45418 188186 45654
rect 188422 45418 188604 45654
rect 188004 45334 188604 45418
rect 188004 45098 188186 45334
rect 188422 45098 188604 45334
rect 188004 9654 188604 45098
rect 188004 9418 188186 9654
rect 188422 9418 188604 9654
rect 188004 9334 188604 9418
rect 188004 9098 188186 9334
rect 188422 9098 188604 9334
rect 188004 -4106 188604 9098
rect 188004 -4342 188186 -4106
rect 188422 -4342 188604 -4106
rect 188004 -4426 188604 -4342
rect 188004 -4662 188186 -4426
rect 188422 -4662 188604 -4426
rect 188004 -5624 188604 -4662
rect 191604 301254 192204 317000
rect 191604 301018 191786 301254
rect 192022 301018 192204 301254
rect 191604 300934 192204 301018
rect 191604 300698 191786 300934
rect 192022 300698 192204 300934
rect 191604 265254 192204 300698
rect 191604 265018 191786 265254
rect 192022 265018 192204 265254
rect 191604 264934 192204 265018
rect 191604 264698 191786 264934
rect 192022 264698 192204 264934
rect 191604 229254 192204 264698
rect 191604 229018 191786 229254
rect 192022 229018 192204 229254
rect 191604 228934 192204 229018
rect 191604 228698 191786 228934
rect 192022 228698 192204 228934
rect 191604 193254 192204 228698
rect 191604 193018 191786 193254
rect 192022 193018 192204 193254
rect 191604 192934 192204 193018
rect 191604 192698 191786 192934
rect 192022 192698 192204 192934
rect 191604 157254 192204 192698
rect 191604 157018 191786 157254
rect 192022 157018 192204 157254
rect 191604 156934 192204 157018
rect 191604 156698 191786 156934
rect 192022 156698 192204 156934
rect 191604 121254 192204 156698
rect 191604 121018 191786 121254
rect 192022 121018 192204 121254
rect 191604 120934 192204 121018
rect 191604 120698 191786 120934
rect 192022 120698 192204 120934
rect 191604 85254 192204 120698
rect 191604 85018 191786 85254
rect 192022 85018 192204 85254
rect 191604 84934 192204 85018
rect 191604 84698 191786 84934
rect 192022 84698 192204 84934
rect 191604 49254 192204 84698
rect 191604 49018 191786 49254
rect 192022 49018 192204 49254
rect 191604 48934 192204 49018
rect 191604 48698 191786 48934
rect 192022 48698 192204 48934
rect 191604 13254 192204 48698
rect 191604 13018 191786 13254
rect 192022 13018 192204 13254
rect 191604 12934 192204 13018
rect 191604 12698 191786 12934
rect 192022 12698 192204 12934
rect 173604 -7162 173786 -6926
rect 174022 -7162 174204 -6926
rect 173604 -7246 174204 -7162
rect 173604 -7482 173786 -7246
rect 174022 -7482 174204 -7246
rect 173604 -7504 174204 -7482
rect 191604 -5986 192204 12698
rect 198804 308454 199404 317000
rect 198804 308218 198986 308454
rect 199222 308218 199404 308454
rect 198804 308134 199404 308218
rect 198804 307898 198986 308134
rect 199222 307898 199404 308134
rect 198804 272454 199404 307898
rect 198804 272218 198986 272454
rect 199222 272218 199404 272454
rect 198804 272134 199404 272218
rect 198804 271898 198986 272134
rect 199222 271898 199404 272134
rect 198804 236454 199404 271898
rect 198804 236218 198986 236454
rect 199222 236218 199404 236454
rect 198804 236134 199404 236218
rect 198804 235898 198986 236134
rect 199222 235898 199404 236134
rect 198804 200454 199404 235898
rect 198804 200218 198986 200454
rect 199222 200218 199404 200454
rect 198804 200134 199404 200218
rect 198804 199898 198986 200134
rect 199222 199898 199404 200134
rect 198804 164454 199404 199898
rect 198804 164218 198986 164454
rect 199222 164218 199404 164454
rect 198804 164134 199404 164218
rect 198804 163898 198986 164134
rect 199222 163898 199404 164134
rect 198804 128454 199404 163898
rect 198804 128218 198986 128454
rect 199222 128218 199404 128454
rect 198804 128134 199404 128218
rect 198804 127898 198986 128134
rect 199222 127898 199404 128134
rect 198804 92454 199404 127898
rect 198804 92218 198986 92454
rect 199222 92218 199404 92454
rect 198804 92134 199404 92218
rect 198804 91898 198986 92134
rect 199222 91898 199404 92134
rect 198804 56454 199404 91898
rect 198804 56218 198986 56454
rect 199222 56218 199404 56454
rect 198804 56134 199404 56218
rect 198804 55898 198986 56134
rect 199222 55898 199404 56134
rect 198804 20454 199404 55898
rect 198804 20218 198986 20454
rect 199222 20218 199404 20454
rect 198804 20134 199404 20218
rect 198804 19898 198986 20134
rect 199222 19898 199404 20134
rect 198804 -1286 199404 19898
rect 198804 -1522 198986 -1286
rect 199222 -1522 199404 -1286
rect 198804 -1606 199404 -1522
rect 198804 -1842 198986 -1606
rect 199222 -1842 199404 -1606
rect 198804 -1864 199404 -1842
rect 202404 312054 203004 317000
rect 202404 311818 202586 312054
rect 202822 311818 203004 312054
rect 202404 311734 203004 311818
rect 202404 311498 202586 311734
rect 202822 311498 203004 311734
rect 202404 276054 203004 311498
rect 202404 275818 202586 276054
rect 202822 275818 203004 276054
rect 202404 275734 203004 275818
rect 202404 275498 202586 275734
rect 202822 275498 203004 275734
rect 202404 240054 203004 275498
rect 202404 239818 202586 240054
rect 202822 239818 203004 240054
rect 202404 239734 203004 239818
rect 202404 239498 202586 239734
rect 202822 239498 203004 239734
rect 202404 204054 203004 239498
rect 202404 203818 202586 204054
rect 202822 203818 203004 204054
rect 202404 203734 203004 203818
rect 202404 203498 202586 203734
rect 202822 203498 203004 203734
rect 202404 168054 203004 203498
rect 202404 167818 202586 168054
rect 202822 167818 203004 168054
rect 202404 167734 203004 167818
rect 202404 167498 202586 167734
rect 202822 167498 203004 167734
rect 202404 132054 203004 167498
rect 202404 131818 202586 132054
rect 202822 131818 203004 132054
rect 202404 131734 203004 131818
rect 202404 131498 202586 131734
rect 202822 131498 203004 131734
rect 202404 96054 203004 131498
rect 202404 95818 202586 96054
rect 202822 95818 203004 96054
rect 202404 95734 203004 95818
rect 202404 95498 202586 95734
rect 202822 95498 203004 95734
rect 202404 60054 203004 95498
rect 202404 59818 202586 60054
rect 202822 59818 203004 60054
rect 202404 59734 203004 59818
rect 202404 59498 202586 59734
rect 202822 59498 203004 59734
rect 202404 24054 203004 59498
rect 202404 23818 202586 24054
rect 202822 23818 203004 24054
rect 202404 23734 203004 23818
rect 202404 23498 202586 23734
rect 202822 23498 203004 23734
rect 202404 -3166 203004 23498
rect 202404 -3402 202586 -3166
rect 202822 -3402 203004 -3166
rect 202404 -3486 203004 -3402
rect 202404 -3722 202586 -3486
rect 202822 -3722 203004 -3486
rect 202404 -3744 203004 -3722
rect 206004 315654 206604 317000
rect 206004 315418 206186 315654
rect 206422 315418 206604 315654
rect 206004 315334 206604 315418
rect 206004 315098 206186 315334
rect 206422 315098 206604 315334
rect 206004 279654 206604 315098
rect 206004 279418 206186 279654
rect 206422 279418 206604 279654
rect 206004 279334 206604 279418
rect 206004 279098 206186 279334
rect 206422 279098 206604 279334
rect 206004 243654 206604 279098
rect 206004 243418 206186 243654
rect 206422 243418 206604 243654
rect 206004 243334 206604 243418
rect 206004 243098 206186 243334
rect 206422 243098 206604 243334
rect 206004 207654 206604 243098
rect 206004 207418 206186 207654
rect 206422 207418 206604 207654
rect 206004 207334 206604 207418
rect 206004 207098 206186 207334
rect 206422 207098 206604 207334
rect 206004 171654 206604 207098
rect 206004 171418 206186 171654
rect 206422 171418 206604 171654
rect 206004 171334 206604 171418
rect 206004 171098 206186 171334
rect 206422 171098 206604 171334
rect 206004 135654 206604 171098
rect 206004 135418 206186 135654
rect 206422 135418 206604 135654
rect 206004 135334 206604 135418
rect 206004 135098 206186 135334
rect 206422 135098 206604 135334
rect 206004 99654 206604 135098
rect 206004 99418 206186 99654
rect 206422 99418 206604 99654
rect 206004 99334 206604 99418
rect 206004 99098 206186 99334
rect 206422 99098 206604 99334
rect 206004 63654 206604 99098
rect 206004 63418 206186 63654
rect 206422 63418 206604 63654
rect 206004 63334 206604 63418
rect 206004 63098 206186 63334
rect 206422 63098 206604 63334
rect 206004 27654 206604 63098
rect 206004 27418 206186 27654
rect 206422 27418 206604 27654
rect 206004 27334 206604 27418
rect 206004 27098 206186 27334
rect 206422 27098 206604 27334
rect 206004 -5046 206604 27098
rect 206004 -5282 206186 -5046
rect 206422 -5282 206604 -5046
rect 206004 -5366 206604 -5282
rect 206004 -5602 206186 -5366
rect 206422 -5602 206604 -5366
rect 206004 -5624 206604 -5602
rect 209604 283254 210204 317000
rect 209604 283018 209786 283254
rect 210022 283018 210204 283254
rect 209604 282934 210204 283018
rect 209604 282698 209786 282934
rect 210022 282698 210204 282934
rect 209604 247254 210204 282698
rect 209604 247018 209786 247254
rect 210022 247018 210204 247254
rect 209604 246934 210204 247018
rect 209604 246698 209786 246934
rect 210022 246698 210204 246934
rect 209604 211254 210204 246698
rect 209604 211018 209786 211254
rect 210022 211018 210204 211254
rect 209604 210934 210204 211018
rect 209604 210698 209786 210934
rect 210022 210698 210204 210934
rect 209604 175254 210204 210698
rect 209604 175018 209786 175254
rect 210022 175018 210204 175254
rect 209604 174934 210204 175018
rect 209604 174698 209786 174934
rect 210022 174698 210204 174934
rect 209604 139254 210204 174698
rect 209604 139018 209786 139254
rect 210022 139018 210204 139254
rect 209604 138934 210204 139018
rect 209604 138698 209786 138934
rect 210022 138698 210204 138934
rect 209604 103254 210204 138698
rect 209604 103018 209786 103254
rect 210022 103018 210204 103254
rect 209604 102934 210204 103018
rect 209604 102698 209786 102934
rect 210022 102698 210204 102934
rect 209604 67254 210204 102698
rect 209604 67018 209786 67254
rect 210022 67018 210204 67254
rect 209604 66934 210204 67018
rect 209604 66698 209786 66934
rect 210022 66698 210204 66934
rect 209604 31254 210204 66698
rect 209604 31018 209786 31254
rect 210022 31018 210204 31254
rect 209604 30934 210204 31018
rect 209604 30698 209786 30934
rect 210022 30698 210204 30934
rect 191604 -6222 191786 -5986
rect 192022 -6222 192204 -5986
rect 191604 -6306 192204 -6222
rect 191604 -6542 191786 -6306
rect 192022 -6542 192204 -6306
rect 191604 -7504 192204 -6542
rect 209604 -6926 210204 30698
rect 216804 290454 217404 317000
rect 216804 290218 216986 290454
rect 217222 290218 217404 290454
rect 216804 290134 217404 290218
rect 216804 289898 216986 290134
rect 217222 289898 217404 290134
rect 216804 254454 217404 289898
rect 216804 254218 216986 254454
rect 217222 254218 217404 254454
rect 216804 254134 217404 254218
rect 216804 253898 216986 254134
rect 217222 253898 217404 254134
rect 216804 218454 217404 253898
rect 216804 218218 216986 218454
rect 217222 218218 217404 218454
rect 216804 218134 217404 218218
rect 216804 217898 216986 218134
rect 217222 217898 217404 218134
rect 216804 182454 217404 217898
rect 216804 182218 216986 182454
rect 217222 182218 217404 182454
rect 216804 182134 217404 182218
rect 216804 181898 216986 182134
rect 217222 181898 217404 182134
rect 216804 146454 217404 181898
rect 216804 146218 216986 146454
rect 217222 146218 217404 146454
rect 216804 146134 217404 146218
rect 216804 145898 216986 146134
rect 217222 145898 217404 146134
rect 216804 110454 217404 145898
rect 216804 110218 216986 110454
rect 217222 110218 217404 110454
rect 216804 110134 217404 110218
rect 216804 109898 216986 110134
rect 217222 109898 217404 110134
rect 216804 74454 217404 109898
rect 216804 74218 216986 74454
rect 217222 74218 217404 74454
rect 216804 74134 217404 74218
rect 216804 73898 216986 74134
rect 217222 73898 217404 74134
rect 216804 38454 217404 73898
rect 216804 38218 216986 38454
rect 217222 38218 217404 38454
rect 216804 38134 217404 38218
rect 216804 37898 216986 38134
rect 217222 37898 217404 38134
rect 216804 2454 217404 37898
rect 216804 2218 216986 2454
rect 217222 2218 217404 2454
rect 216804 2134 217404 2218
rect 216804 1898 216986 2134
rect 217222 1898 217404 2134
rect 216804 -346 217404 1898
rect 216804 -582 216986 -346
rect 217222 -582 217404 -346
rect 216804 -666 217404 -582
rect 216804 -902 216986 -666
rect 217222 -902 217404 -666
rect 216804 -1864 217404 -902
rect 220404 294054 221004 317000
rect 220404 293818 220586 294054
rect 220822 293818 221004 294054
rect 220404 293734 221004 293818
rect 220404 293498 220586 293734
rect 220822 293498 221004 293734
rect 220404 258054 221004 293498
rect 220404 257818 220586 258054
rect 220822 257818 221004 258054
rect 220404 257734 221004 257818
rect 220404 257498 220586 257734
rect 220822 257498 221004 257734
rect 220404 222054 221004 257498
rect 220404 221818 220586 222054
rect 220822 221818 221004 222054
rect 220404 221734 221004 221818
rect 220404 221498 220586 221734
rect 220822 221498 221004 221734
rect 220404 186054 221004 221498
rect 220404 185818 220586 186054
rect 220822 185818 221004 186054
rect 220404 185734 221004 185818
rect 220404 185498 220586 185734
rect 220822 185498 221004 185734
rect 220404 150054 221004 185498
rect 220404 149818 220586 150054
rect 220822 149818 221004 150054
rect 220404 149734 221004 149818
rect 220404 149498 220586 149734
rect 220822 149498 221004 149734
rect 220404 114054 221004 149498
rect 220404 113818 220586 114054
rect 220822 113818 221004 114054
rect 220404 113734 221004 113818
rect 220404 113498 220586 113734
rect 220822 113498 221004 113734
rect 220404 78054 221004 113498
rect 220404 77818 220586 78054
rect 220822 77818 221004 78054
rect 220404 77734 221004 77818
rect 220404 77498 220586 77734
rect 220822 77498 221004 77734
rect 220404 42054 221004 77498
rect 220404 41818 220586 42054
rect 220822 41818 221004 42054
rect 220404 41734 221004 41818
rect 220404 41498 220586 41734
rect 220822 41498 221004 41734
rect 220404 6054 221004 41498
rect 220404 5818 220586 6054
rect 220822 5818 221004 6054
rect 220404 5734 221004 5818
rect 220404 5498 220586 5734
rect 220822 5498 221004 5734
rect 220404 -2226 221004 5498
rect 220404 -2462 220586 -2226
rect 220822 -2462 221004 -2226
rect 220404 -2546 221004 -2462
rect 220404 -2782 220586 -2546
rect 220822 -2782 221004 -2546
rect 220404 -3744 221004 -2782
rect 224004 297654 224604 317000
rect 224004 297418 224186 297654
rect 224422 297418 224604 297654
rect 224004 297334 224604 297418
rect 224004 297098 224186 297334
rect 224422 297098 224604 297334
rect 224004 261654 224604 297098
rect 224004 261418 224186 261654
rect 224422 261418 224604 261654
rect 224004 261334 224604 261418
rect 224004 261098 224186 261334
rect 224422 261098 224604 261334
rect 224004 225654 224604 261098
rect 224004 225418 224186 225654
rect 224422 225418 224604 225654
rect 224004 225334 224604 225418
rect 224004 225098 224186 225334
rect 224422 225098 224604 225334
rect 224004 189654 224604 225098
rect 224004 189418 224186 189654
rect 224422 189418 224604 189654
rect 224004 189334 224604 189418
rect 224004 189098 224186 189334
rect 224422 189098 224604 189334
rect 224004 153654 224604 189098
rect 224004 153418 224186 153654
rect 224422 153418 224604 153654
rect 224004 153334 224604 153418
rect 224004 153098 224186 153334
rect 224422 153098 224604 153334
rect 224004 117654 224604 153098
rect 224004 117418 224186 117654
rect 224422 117418 224604 117654
rect 224004 117334 224604 117418
rect 224004 117098 224186 117334
rect 224422 117098 224604 117334
rect 224004 81654 224604 117098
rect 224004 81418 224186 81654
rect 224422 81418 224604 81654
rect 224004 81334 224604 81418
rect 224004 81098 224186 81334
rect 224422 81098 224604 81334
rect 224004 45654 224604 81098
rect 224004 45418 224186 45654
rect 224422 45418 224604 45654
rect 224004 45334 224604 45418
rect 224004 45098 224186 45334
rect 224422 45098 224604 45334
rect 224004 9654 224604 45098
rect 224004 9418 224186 9654
rect 224422 9418 224604 9654
rect 224004 9334 224604 9418
rect 224004 9098 224186 9334
rect 224422 9098 224604 9334
rect 224004 -4106 224604 9098
rect 224004 -4342 224186 -4106
rect 224422 -4342 224604 -4106
rect 224004 -4426 224604 -4342
rect 224004 -4662 224186 -4426
rect 224422 -4662 224604 -4426
rect 224004 -5624 224604 -4662
rect 227604 301254 228204 317000
rect 227604 301018 227786 301254
rect 228022 301018 228204 301254
rect 227604 300934 228204 301018
rect 227604 300698 227786 300934
rect 228022 300698 228204 300934
rect 227604 265254 228204 300698
rect 227604 265018 227786 265254
rect 228022 265018 228204 265254
rect 227604 264934 228204 265018
rect 227604 264698 227786 264934
rect 228022 264698 228204 264934
rect 227604 229254 228204 264698
rect 227604 229018 227786 229254
rect 228022 229018 228204 229254
rect 227604 228934 228204 229018
rect 227604 228698 227786 228934
rect 228022 228698 228204 228934
rect 227604 193254 228204 228698
rect 227604 193018 227786 193254
rect 228022 193018 228204 193254
rect 227604 192934 228204 193018
rect 227604 192698 227786 192934
rect 228022 192698 228204 192934
rect 227604 157254 228204 192698
rect 227604 157018 227786 157254
rect 228022 157018 228204 157254
rect 227604 156934 228204 157018
rect 227604 156698 227786 156934
rect 228022 156698 228204 156934
rect 227604 121254 228204 156698
rect 227604 121018 227786 121254
rect 228022 121018 228204 121254
rect 227604 120934 228204 121018
rect 227604 120698 227786 120934
rect 228022 120698 228204 120934
rect 227604 85254 228204 120698
rect 227604 85018 227786 85254
rect 228022 85018 228204 85254
rect 227604 84934 228204 85018
rect 227604 84698 227786 84934
rect 228022 84698 228204 84934
rect 227604 49254 228204 84698
rect 227604 49018 227786 49254
rect 228022 49018 228204 49254
rect 227604 48934 228204 49018
rect 227604 48698 227786 48934
rect 228022 48698 228204 48934
rect 227604 13254 228204 48698
rect 227604 13018 227786 13254
rect 228022 13018 228204 13254
rect 227604 12934 228204 13018
rect 227604 12698 227786 12934
rect 228022 12698 228204 12934
rect 209604 -7162 209786 -6926
rect 210022 -7162 210204 -6926
rect 209604 -7246 210204 -7162
rect 209604 -7482 209786 -7246
rect 210022 -7482 210204 -7246
rect 209604 -7504 210204 -7482
rect 227604 -5986 228204 12698
rect 234804 308454 235404 317000
rect 234804 308218 234986 308454
rect 235222 308218 235404 308454
rect 234804 308134 235404 308218
rect 234804 307898 234986 308134
rect 235222 307898 235404 308134
rect 234804 272454 235404 307898
rect 234804 272218 234986 272454
rect 235222 272218 235404 272454
rect 234804 272134 235404 272218
rect 234804 271898 234986 272134
rect 235222 271898 235404 272134
rect 234804 236454 235404 271898
rect 234804 236218 234986 236454
rect 235222 236218 235404 236454
rect 234804 236134 235404 236218
rect 234804 235898 234986 236134
rect 235222 235898 235404 236134
rect 234804 200454 235404 235898
rect 234804 200218 234986 200454
rect 235222 200218 235404 200454
rect 234804 200134 235404 200218
rect 234804 199898 234986 200134
rect 235222 199898 235404 200134
rect 234804 164454 235404 199898
rect 234804 164218 234986 164454
rect 235222 164218 235404 164454
rect 234804 164134 235404 164218
rect 234804 163898 234986 164134
rect 235222 163898 235404 164134
rect 234804 128454 235404 163898
rect 234804 128218 234986 128454
rect 235222 128218 235404 128454
rect 234804 128134 235404 128218
rect 234804 127898 234986 128134
rect 235222 127898 235404 128134
rect 234804 92454 235404 127898
rect 234804 92218 234986 92454
rect 235222 92218 235404 92454
rect 234804 92134 235404 92218
rect 234804 91898 234986 92134
rect 235222 91898 235404 92134
rect 234804 56454 235404 91898
rect 234804 56218 234986 56454
rect 235222 56218 235404 56454
rect 234804 56134 235404 56218
rect 234804 55898 234986 56134
rect 235222 55898 235404 56134
rect 234804 20454 235404 55898
rect 234804 20218 234986 20454
rect 235222 20218 235404 20454
rect 234804 20134 235404 20218
rect 234804 19898 234986 20134
rect 235222 19898 235404 20134
rect 234804 -1286 235404 19898
rect 234804 -1522 234986 -1286
rect 235222 -1522 235404 -1286
rect 234804 -1606 235404 -1522
rect 234804 -1842 234986 -1606
rect 235222 -1842 235404 -1606
rect 234804 -1864 235404 -1842
rect 238404 312054 239004 317000
rect 238404 311818 238586 312054
rect 238822 311818 239004 312054
rect 238404 311734 239004 311818
rect 238404 311498 238586 311734
rect 238822 311498 239004 311734
rect 238404 276054 239004 311498
rect 238404 275818 238586 276054
rect 238822 275818 239004 276054
rect 238404 275734 239004 275818
rect 238404 275498 238586 275734
rect 238822 275498 239004 275734
rect 238404 240054 239004 275498
rect 238404 239818 238586 240054
rect 238822 239818 239004 240054
rect 238404 239734 239004 239818
rect 238404 239498 238586 239734
rect 238822 239498 239004 239734
rect 238404 204054 239004 239498
rect 238404 203818 238586 204054
rect 238822 203818 239004 204054
rect 238404 203734 239004 203818
rect 238404 203498 238586 203734
rect 238822 203498 239004 203734
rect 238404 168054 239004 203498
rect 238404 167818 238586 168054
rect 238822 167818 239004 168054
rect 238404 167734 239004 167818
rect 238404 167498 238586 167734
rect 238822 167498 239004 167734
rect 238404 132054 239004 167498
rect 238404 131818 238586 132054
rect 238822 131818 239004 132054
rect 238404 131734 239004 131818
rect 238404 131498 238586 131734
rect 238822 131498 239004 131734
rect 238404 96054 239004 131498
rect 238404 95818 238586 96054
rect 238822 95818 239004 96054
rect 238404 95734 239004 95818
rect 238404 95498 238586 95734
rect 238822 95498 239004 95734
rect 238404 60054 239004 95498
rect 238404 59818 238586 60054
rect 238822 59818 239004 60054
rect 238404 59734 239004 59818
rect 238404 59498 238586 59734
rect 238822 59498 239004 59734
rect 238404 24054 239004 59498
rect 238404 23818 238586 24054
rect 238822 23818 239004 24054
rect 238404 23734 239004 23818
rect 238404 23498 238586 23734
rect 238822 23498 239004 23734
rect 238404 -3166 239004 23498
rect 238404 -3402 238586 -3166
rect 238822 -3402 239004 -3166
rect 238404 -3486 239004 -3402
rect 238404 -3722 238586 -3486
rect 238822 -3722 239004 -3486
rect 238404 -3744 239004 -3722
rect 242004 315654 242604 317000
rect 242004 315418 242186 315654
rect 242422 315418 242604 315654
rect 242004 315334 242604 315418
rect 242004 315098 242186 315334
rect 242422 315098 242604 315334
rect 242004 279654 242604 315098
rect 242004 279418 242186 279654
rect 242422 279418 242604 279654
rect 242004 279334 242604 279418
rect 242004 279098 242186 279334
rect 242422 279098 242604 279334
rect 242004 243654 242604 279098
rect 242004 243418 242186 243654
rect 242422 243418 242604 243654
rect 242004 243334 242604 243418
rect 242004 243098 242186 243334
rect 242422 243098 242604 243334
rect 242004 207654 242604 243098
rect 242004 207418 242186 207654
rect 242422 207418 242604 207654
rect 242004 207334 242604 207418
rect 242004 207098 242186 207334
rect 242422 207098 242604 207334
rect 242004 171654 242604 207098
rect 242004 171418 242186 171654
rect 242422 171418 242604 171654
rect 242004 171334 242604 171418
rect 242004 171098 242186 171334
rect 242422 171098 242604 171334
rect 242004 135654 242604 171098
rect 242004 135418 242186 135654
rect 242422 135418 242604 135654
rect 242004 135334 242604 135418
rect 242004 135098 242186 135334
rect 242422 135098 242604 135334
rect 242004 99654 242604 135098
rect 242004 99418 242186 99654
rect 242422 99418 242604 99654
rect 242004 99334 242604 99418
rect 242004 99098 242186 99334
rect 242422 99098 242604 99334
rect 242004 63654 242604 99098
rect 242004 63418 242186 63654
rect 242422 63418 242604 63654
rect 242004 63334 242604 63418
rect 242004 63098 242186 63334
rect 242422 63098 242604 63334
rect 242004 27654 242604 63098
rect 242004 27418 242186 27654
rect 242422 27418 242604 27654
rect 242004 27334 242604 27418
rect 242004 27098 242186 27334
rect 242422 27098 242604 27334
rect 242004 -5046 242604 27098
rect 242004 -5282 242186 -5046
rect 242422 -5282 242604 -5046
rect 242004 -5366 242604 -5282
rect 242004 -5602 242186 -5366
rect 242422 -5602 242604 -5366
rect 242004 -5624 242604 -5602
rect 245604 283254 246204 317000
rect 245604 283018 245786 283254
rect 246022 283018 246204 283254
rect 245604 282934 246204 283018
rect 245604 282698 245786 282934
rect 246022 282698 246204 282934
rect 245604 247254 246204 282698
rect 245604 247018 245786 247254
rect 246022 247018 246204 247254
rect 245604 246934 246204 247018
rect 245604 246698 245786 246934
rect 246022 246698 246204 246934
rect 245604 211254 246204 246698
rect 245604 211018 245786 211254
rect 246022 211018 246204 211254
rect 245604 210934 246204 211018
rect 245604 210698 245786 210934
rect 246022 210698 246204 210934
rect 245604 175254 246204 210698
rect 245604 175018 245786 175254
rect 246022 175018 246204 175254
rect 245604 174934 246204 175018
rect 245604 174698 245786 174934
rect 246022 174698 246204 174934
rect 245604 139254 246204 174698
rect 245604 139018 245786 139254
rect 246022 139018 246204 139254
rect 245604 138934 246204 139018
rect 245604 138698 245786 138934
rect 246022 138698 246204 138934
rect 245604 103254 246204 138698
rect 245604 103018 245786 103254
rect 246022 103018 246204 103254
rect 245604 102934 246204 103018
rect 245604 102698 245786 102934
rect 246022 102698 246204 102934
rect 245604 67254 246204 102698
rect 245604 67018 245786 67254
rect 246022 67018 246204 67254
rect 245604 66934 246204 67018
rect 245604 66698 245786 66934
rect 246022 66698 246204 66934
rect 245604 31254 246204 66698
rect 245604 31018 245786 31254
rect 246022 31018 246204 31254
rect 245604 30934 246204 31018
rect 245604 30698 245786 30934
rect 246022 30698 246204 30934
rect 227604 -6222 227786 -5986
rect 228022 -6222 228204 -5986
rect 227604 -6306 228204 -6222
rect 227604 -6542 227786 -6306
rect 228022 -6542 228204 -6306
rect 227604 -7504 228204 -6542
rect 245604 -6926 246204 30698
rect 252804 290454 253404 317000
rect 252804 290218 252986 290454
rect 253222 290218 253404 290454
rect 252804 290134 253404 290218
rect 252804 289898 252986 290134
rect 253222 289898 253404 290134
rect 252804 254454 253404 289898
rect 252804 254218 252986 254454
rect 253222 254218 253404 254454
rect 252804 254134 253404 254218
rect 252804 253898 252986 254134
rect 253222 253898 253404 254134
rect 252804 218454 253404 253898
rect 252804 218218 252986 218454
rect 253222 218218 253404 218454
rect 252804 218134 253404 218218
rect 252804 217898 252986 218134
rect 253222 217898 253404 218134
rect 252804 182454 253404 217898
rect 252804 182218 252986 182454
rect 253222 182218 253404 182454
rect 252804 182134 253404 182218
rect 252804 181898 252986 182134
rect 253222 181898 253404 182134
rect 252804 146454 253404 181898
rect 252804 146218 252986 146454
rect 253222 146218 253404 146454
rect 252804 146134 253404 146218
rect 252804 145898 252986 146134
rect 253222 145898 253404 146134
rect 252804 110454 253404 145898
rect 252804 110218 252986 110454
rect 253222 110218 253404 110454
rect 252804 110134 253404 110218
rect 252804 109898 252986 110134
rect 253222 109898 253404 110134
rect 252804 74454 253404 109898
rect 252804 74218 252986 74454
rect 253222 74218 253404 74454
rect 252804 74134 253404 74218
rect 252804 73898 252986 74134
rect 253222 73898 253404 74134
rect 252804 38454 253404 73898
rect 252804 38218 252986 38454
rect 253222 38218 253404 38454
rect 252804 38134 253404 38218
rect 252804 37898 252986 38134
rect 253222 37898 253404 38134
rect 252804 2454 253404 37898
rect 252804 2218 252986 2454
rect 253222 2218 253404 2454
rect 252804 2134 253404 2218
rect 252804 1898 252986 2134
rect 253222 1898 253404 2134
rect 252804 -346 253404 1898
rect 252804 -582 252986 -346
rect 253222 -582 253404 -346
rect 252804 -666 253404 -582
rect 252804 -902 252986 -666
rect 253222 -902 253404 -666
rect 252804 -1864 253404 -902
rect 256404 294054 257004 317000
rect 256404 293818 256586 294054
rect 256822 293818 257004 294054
rect 256404 293734 257004 293818
rect 256404 293498 256586 293734
rect 256822 293498 257004 293734
rect 256404 258054 257004 293498
rect 256404 257818 256586 258054
rect 256822 257818 257004 258054
rect 256404 257734 257004 257818
rect 256404 257498 256586 257734
rect 256822 257498 257004 257734
rect 256404 222054 257004 257498
rect 256404 221818 256586 222054
rect 256822 221818 257004 222054
rect 256404 221734 257004 221818
rect 256404 221498 256586 221734
rect 256822 221498 257004 221734
rect 256404 186054 257004 221498
rect 256404 185818 256586 186054
rect 256822 185818 257004 186054
rect 256404 185734 257004 185818
rect 256404 185498 256586 185734
rect 256822 185498 257004 185734
rect 256404 150054 257004 185498
rect 256404 149818 256586 150054
rect 256822 149818 257004 150054
rect 256404 149734 257004 149818
rect 256404 149498 256586 149734
rect 256822 149498 257004 149734
rect 256404 114054 257004 149498
rect 256404 113818 256586 114054
rect 256822 113818 257004 114054
rect 256404 113734 257004 113818
rect 256404 113498 256586 113734
rect 256822 113498 257004 113734
rect 256404 78054 257004 113498
rect 256404 77818 256586 78054
rect 256822 77818 257004 78054
rect 256404 77734 257004 77818
rect 256404 77498 256586 77734
rect 256822 77498 257004 77734
rect 256404 42054 257004 77498
rect 256404 41818 256586 42054
rect 256822 41818 257004 42054
rect 256404 41734 257004 41818
rect 256404 41498 256586 41734
rect 256822 41498 257004 41734
rect 256404 6054 257004 41498
rect 256404 5818 256586 6054
rect 256822 5818 257004 6054
rect 256404 5734 257004 5818
rect 256404 5498 256586 5734
rect 256822 5498 257004 5734
rect 256404 -2226 257004 5498
rect 256404 -2462 256586 -2226
rect 256822 -2462 257004 -2226
rect 256404 -2546 257004 -2462
rect 256404 -2782 256586 -2546
rect 256822 -2782 257004 -2546
rect 256404 -3744 257004 -2782
rect 260004 297654 260604 317000
rect 260004 297418 260186 297654
rect 260422 297418 260604 297654
rect 260004 297334 260604 297418
rect 260004 297098 260186 297334
rect 260422 297098 260604 297334
rect 260004 261654 260604 297098
rect 260004 261418 260186 261654
rect 260422 261418 260604 261654
rect 260004 261334 260604 261418
rect 260004 261098 260186 261334
rect 260422 261098 260604 261334
rect 260004 225654 260604 261098
rect 260004 225418 260186 225654
rect 260422 225418 260604 225654
rect 260004 225334 260604 225418
rect 260004 225098 260186 225334
rect 260422 225098 260604 225334
rect 260004 189654 260604 225098
rect 260004 189418 260186 189654
rect 260422 189418 260604 189654
rect 260004 189334 260604 189418
rect 260004 189098 260186 189334
rect 260422 189098 260604 189334
rect 260004 153654 260604 189098
rect 260004 153418 260186 153654
rect 260422 153418 260604 153654
rect 260004 153334 260604 153418
rect 260004 153098 260186 153334
rect 260422 153098 260604 153334
rect 260004 117654 260604 153098
rect 260004 117418 260186 117654
rect 260422 117418 260604 117654
rect 260004 117334 260604 117418
rect 260004 117098 260186 117334
rect 260422 117098 260604 117334
rect 260004 81654 260604 117098
rect 260004 81418 260186 81654
rect 260422 81418 260604 81654
rect 260004 81334 260604 81418
rect 260004 81098 260186 81334
rect 260422 81098 260604 81334
rect 260004 45654 260604 81098
rect 260004 45418 260186 45654
rect 260422 45418 260604 45654
rect 260004 45334 260604 45418
rect 260004 45098 260186 45334
rect 260422 45098 260604 45334
rect 260004 9654 260604 45098
rect 260004 9418 260186 9654
rect 260422 9418 260604 9654
rect 260004 9334 260604 9418
rect 260004 9098 260186 9334
rect 260422 9098 260604 9334
rect 260004 -4106 260604 9098
rect 260004 -4342 260186 -4106
rect 260422 -4342 260604 -4106
rect 260004 -4426 260604 -4342
rect 260004 -4662 260186 -4426
rect 260422 -4662 260604 -4426
rect 260004 -5624 260604 -4662
rect 263604 301254 264204 317000
rect 263604 301018 263786 301254
rect 264022 301018 264204 301254
rect 263604 300934 264204 301018
rect 263604 300698 263786 300934
rect 264022 300698 264204 300934
rect 263604 265254 264204 300698
rect 263604 265018 263786 265254
rect 264022 265018 264204 265254
rect 263604 264934 264204 265018
rect 263604 264698 263786 264934
rect 264022 264698 264204 264934
rect 263604 229254 264204 264698
rect 263604 229018 263786 229254
rect 264022 229018 264204 229254
rect 263604 228934 264204 229018
rect 263604 228698 263786 228934
rect 264022 228698 264204 228934
rect 263604 193254 264204 228698
rect 263604 193018 263786 193254
rect 264022 193018 264204 193254
rect 263604 192934 264204 193018
rect 263604 192698 263786 192934
rect 264022 192698 264204 192934
rect 263604 157254 264204 192698
rect 263604 157018 263786 157254
rect 264022 157018 264204 157254
rect 263604 156934 264204 157018
rect 263604 156698 263786 156934
rect 264022 156698 264204 156934
rect 263604 121254 264204 156698
rect 263604 121018 263786 121254
rect 264022 121018 264204 121254
rect 263604 120934 264204 121018
rect 263604 120698 263786 120934
rect 264022 120698 264204 120934
rect 263604 85254 264204 120698
rect 263604 85018 263786 85254
rect 264022 85018 264204 85254
rect 263604 84934 264204 85018
rect 263604 84698 263786 84934
rect 264022 84698 264204 84934
rect 263604 49254 264204 84698
rect 263604 49018 263786 49254
rect 264022 49018 264204 49254
rect 263604 48934 264204 49018
rect 263604 48698 263786 48934
rect 264022 48698 264204 48934
rect 263604 13254 264204 48698
rect 263604 13018 263786 13254
rect 264022 13018 264204 13254
rect 263604 12934 264204 13018
rect 263604 12698 263786 12934
rect 264022 12698 264204 12934
rect 245604 -7162 245786 -6926
rect 246022 -7162 246204 -6926
rect 245604 -7246 246204 -7162
rect 245604 -7482 245786 -7246
rect 246022 -7482 246204 -7246
rect 245604 -7504 246204 -7482
rect 263604 -5986 264204 12698
rect 270804 308454 271404 317000
rect 270804 308218 270986 308454
rect 271222 308218 271404 308454
rect 270804 308134 271404 308218
rect 270804 307898 270986 308134
rect 271222 307898 271404 308134
rect 270804 272454 271404 307898
rect 270804 272218 270986 272454
rect 271222 272218 271404 272454
rect 270804 272134 271404 272218
rect 270804 271898 270986 272134
rect 271222 271898 271404 272134
rect 270804 236454 271404 271898
rect 270804 236218 270986 236454
rect 271222 236218 271404 236454
rect 270804 236134 271404 236218
rect 270804 235898 270986 236134
rect 271222 235898 271404 236134
rect 270804 200454 271404 235898
rect 270804 200218 270986 200454
rect 271222 200218 271404 200454
rect 270804 200134 271404 200218
rect 270804 199898 270986 200134
rect 271222 199898 271404 200134
rect 270804 164454 271404 199898
rect 270804 164218 270986 164454
rect 271222 164218 271404 164454
rect 270804 164134 271404 164218
rect 270804 163898 270986 164134
rect 271222 163898 271404 164134
rect 270804 128454 271404 163898
rect 270804 128218 270986 128454
rect 271222 128218 271404 128454
rect 270804 128134 271404 128218
rect 270804 127898 270986 128134
rect 271222 127898 271404 128134
rect 270804 92454 271404 127898
rect 270804 92218 270986 92454
rect 271222 92218 271404 92454
rect 270804 92134 271404 92218
rect 270804 91898 270986 92134
rect 271222 91898 271404 92134
rect 270804 56454 271404 91898
rect 270804 56218 270986 56454
rect 271222 56218 271404 56454
rect 270804 56134 271404 56218
rect 270804 55898 270986 56134
rect 271222 55898 271404 56134
rect 270804 20454 271404 55898
rect 270804 20218 270986 20454
rect 271222 20218 271404 20454
rect 270804 20134 271404 20218
rect 270804 19898 270986 20134
rect 271222 19898 271404 20134
rect 270804 -1286 271404 19898
rect 270804 -1522 270986 -1286
rect 271222 -1522 271404 -1286
rect 270804 -1606 271404 -1522
rect 270804 -1842 270986 -1606
rect 271222 -1842 271404 -1606
rect 270804 -1864 271404 -1842
rect 274404 312054 275004 317000
rect 274404 311818 274586 312054
rect 274822 311818 275004 312054
rect 274404 311734 275004 311818
rect 274404 311498 274586 311734
rect 274822 311498 275004 311734
rect 274404 276054 275004 311498
rect 274404 275818 274586 276054
rect 274822 275818 275004 276054
rect 274404 275734 275004 275818
rect 274404 275498 274586 275734
rect 274822 275498 275004 275734
rect 274404 240054 275004 275498
rect 274404 239818 274586 240054
rect 274822 239818 275004 240054
rect 274404 239734 275004 239818
rect 274404 239498 274586 239734
rect 274822 239498 275004 239734
rect 274404 204054 275004 239498
rect 274404 203818 274586 204054
rect 274822 203818 275004 204054
rect 274404 203734 275004 203818
rect 274404 203498 274586 203734
rect 274822 203498 275004 203734
rect 274404 168054 275004 203498
rect 274404 167818 274586 168054
rect 274822 167818 275004 168054
rect 274404 167734 275004 167818
rect 274404 167498 274586 167734
rect 274822 167498 275004 167734
rect 274404 132054 275004 167498
rect 274404 131818 274586 132054
rect 274822 131818 275004 132054
rect 274404 131734 275004 131818
rect 274404 131498 274586 131734
rect 274822 131498 275004 131734
rect 274404 96054 275004 131498
rect 274404 95818 274586 96054
rect 274822 95818 275004 96054
rect 274404 95734 275004 95818
rect 274404 95498 274586 95734
rect 274822 95498 275004 95734
rect 274404 60054 275004 95498
rect 274404 59818 274586 60054
rect 274822 59818 275004 60054
rect 274404 59734 275004 59818
rect 274404 59498 274586 59734
rect 274822 59498 275004 59734
rect 274404 24054 275004 59498
rect 274404 23818 274586 24054
rect 274822 23818 275004 24054
rect 274404 23734 275004 23818
rect 274404 23498 274586 23734
rect 274822 23498 275004 23734
rect 274404 -3166 275004 23498
rect 274404 -3402 274586 -3166
rect 274822 -3402 275004 -3166
rect 274404 -3486 275004 -3402
rect 274404 -3722 274586 -3486
rect 274822 -3722 275004 -3486
rect 274404 -3744 275004 -3722
rect 278004 315654 278604 317000
rect 278004 315418 278186 315654
rect 278422 315418 278604 315654
rect 278004 315334 278604 315418
rect 278004 315098 278186 315334
rect 278422 315098 278604 315334
rect 278004 279654 278604 315098
rect 278004 279418 278186 279654
rect 278422 279418 278604 279654
rect 278004 279334 278604 279418
rect 278004 279098 278186 279334
rect 278422 279098 278604 279334
rect 278004 243654 278604 279098
rect 278004 243418 278186 243654
rect 278422 243418 278604 243654
rect 278004 243334 278604 243418
rect 278004 243098 278186 243334
rect 278422 243098 278604 243334
rect 278004 207654 278604 243098
rect 278004 207418 278186 207654
rect 278422 207418 278604 207654
rect 278004 207334 278604 207418
rect 278004 207098 278186 207334
rect 278422 207098 278604 207334
rect 278004 171654 278604 207098
rect 278004 171418 278186 171654
rect 278422 171418 278604 171654
rect 278004 171334 278604 171418
rect 278004 171098 278186 171334
rect 278422 171098 278604 171334
rect 278004 135654 278604 171098
rect 278004 135418 278186 135654
rect 278422 135418 278604 135654
rect 278004 135334 278604 135418
rect 278004 135098 278186 135334
rect 278422 135098 278604 135334
rect 278004 99654 278604 135098
rect 278004 99418 278186 99654
rect 278422 99418 278604 99654
rect 278004 99334 278604 99418
rect 278004 99098 278186 99334
rect 278422 99098 278604 99334
rect 278004 63654 278604 99098
rect 278004 63418 278186 63654
rect 278422 63418 278604 63654
rect 278004 63334 278604 63418
rect 278004 63098 278186 63334
rect 278422 63098 278604 63334
rect 278004 27654 278604 63098
rect 278004 27418 278186 27654
rect 278422 27418 278604 27654
rect 278004 27334 278604 27418
rect 278004 27098 278186 27334
rect 278422 27098 278604 27334
rect 278004 -5046 278604 27098
rect 278004 -5282 278186 -5046
rect 278422 -5282 278604 -5046
rect 278004 -5366 278604 -5282
rect 278004 -5602 278186 -5366
rect 278422 -5602 278604 -5366
rect 278004 -5624 278604 -5602
rect 281604 283254 282204 317000
rect 281604 283018 281786 283254
rect 282022 283018 282204 283254
rect 281604 282934 282204 283018
rect 281604 282698 281786 282934
rect 282022 282698 282204 282934
rect 281604 247254 282204 282698
rect 281604 247018 281786 247254
rect 282022 247018 282204 247254
rect 281604 246934 282204 247018
rect 281604 246698 281786 246934
rect 282022 246698 282204 246934
rect 281604 211254 282204 246698
rect 281604 211018 281786 211254
rect 282022 211018 282204 211254
rect 281604 210934 282204 211018
rect 281604 210698 281786 210934
rect 282022 210698 282204 210934
rect 281604 175254 282204 210698
rect 281604 175018 281786 175254
rect 282022 175018 282204 175254
rect 281604 174934 282204 175018
rect 281604 174698 281786 174934
rect 282022 174698 282204 174934
rect 281604 139254 282204 174698
rect 281604 139018 281786 139254
rect 282022 139018 282204 139254
rect 281604 138934 282204 139018
rect 281604 138698 281786 138934
rect 282022 138698 282204 138934
rect 281604 103254 282204 138698
rect 281604 103018 281786 103254
rect 282022 103018 282204 103254
rect 281604 102934 282204 103018
rect 281604 102698 281786 102934
rect 282022 102698 282204 102934
rect 281604 67254 282204 102698
rect 281604 67018 281786 67254
rect 282022 67018 282204 67254
rect 281604 66934 282204 67018
rect 281604 66698 281786 66934
rect 282022 66698 282204 66934
rect 281604 31254 282204 66698
rect 281604 31018 281786 31254
rect 282022 31018 282204 31254
rect 281604 30934 282204 31018
rect 281604 30698 281786 30934
rect 282022 30698 282204 30934
rect 263604 -6222 263786 -5986
rect 264022 -6222 264204 -5986
rect 263604 -6306 264204 -6222
rect 263604 -6542 263786 -6306
rect 264022 -6542 264204 -6306
rect 263604 -7504 264204 -6542
rect 281604 -6926 282204 30698
rect 288804 290454 289404 325898
rect 288804 290218 288986 290454
rect 289222 290218 289404 290454
rect 288804 290134 289404 290218
rect 288804 289898 288986 290134
rect 289222 289898 289404 290134
rect 288804 254454 289404 289898
rect 288804 254218 288986 254454
rect 289222 254218 289404 254454
rect 288804 254134 289404 254218
rect 288804 253898 288986 254134
rect 289222 253898 289404 254134
rect 288804 218454 289404 253898
rect 288804 218218 288986 218454
rect 289222 218218 289404 218454
rect 288804 218134 289404 218218
rect 288804 217898 288986 218134
rect 289222 217898 289404 218134
rect 288804 182454 289404 217898
rect 288804 182218 288986 182454
rect 289222 182218 289404 182454
rect 288804 182134 289404 182218
rect 288804 181898 288986 182134
rect 289222 181898 289404 182134
rect 288804 146454 289404 181898
rect 288804 146218 288986 146454
rect 289222 146218 289404 146454
rect 288804 146134 289404 146218
rect 288804 145898 288986 146134
rect 289222 145898 289404 146134
rect 288804 110454 289404 145898
rect 288804 110218 288986 110454
rect 289222 110218 289404 110454
rect 288804 110134 289404 110218
rect 288804 109898 288986 110134
rect 289222 109898 289404 110134
rect 288804 74454 289404 109898
rect 288804 74218 288986 74454
rect 289222 74218 289404 74454
rect 288804 74134 289404 74218
rect 288804 73898 288986 74134
rect 289222 73898 289404 74134
rect 288804 38454 289404 73898
rect 288804 38218 288986 38454
rect 289222 38218 289404 38454
rect 288804 38134 289404 38218
rect 288804 37898 288986 38134
rect 289222 37898 289404 38134
rect 288804 2454 289404 37898
rect 288804 2218 288986 2454
rect 289222 2218 289404 2454
rect 288804 2134 289404 2218
rect 288804 1898 288986 2134
rect 289222 1898 289404 2134
rect 288804 -346 289404 1898
rect 288804 -582 288986 -346
rect 289222 -582 289404 -346
rect 288804 -666 289404 -582
rect 288804 -902 288986 -666
rect 289222 -902 289404 -666
rect 288804 -1864 289404 -902
rect 292404 690054 293004 706162
rect 292404 689818 292586 690054
rect 292822 689818 293004 690054
rect 292404 689734 293004 689818
rect 292404 689498 292586 689734
rect 292822 689498 293004 689734
rect 292404 654054 293004 689498
rect 292404 653818 292586 654054
rect 292822 653818 293004 654054
rect 292404 653734 293004 653818
rect 292404 653498 292586 653734
rect 292822 653498 293004 653734
rect 292404 618054 293004 653498
rect 292404 617818 292586 618054
rect 292822 617818 293004 618054
rect 292404 617734 293004 617818
rect 292404 617498 292586 617734
rect 292822 617498 293004 617734
rect 292404 582054 293004 617498
rect 292404 581818 292586 582054
rect 292822 581818 293004 582054
rect 292404 581734 293004 581818
rect 292404 581498 292586 581734
rect 292822 581498 293004 581734
rect 292404 546054 293004 581498
rect 292404 545818 292586 546054
rect 292822 545818 293004 546054
rect 292404 545734 293004 545818
rect 292404 545498 292586 545734
rect 292822 545498 293004 545734
rect 292404 510054 293004 545498
rect 292404 509818 292586 510054
rect 292822 509818 293004 510054
rect 292404 509734 293004 509818
rect 292404 509498 292586 509734
rect 292822 509498 293004 509734
rect 292404 474054 293004 509498
rect 292404 473818 292586 474054
rect 292822 473818 293004 474054
rect 292404 473734 293004 473818
rect 292404 473498 292586 473734
rect 292822 473498 293004 473734
rect 292404 438054 293004 473498
rect 292404 437818 292586 438054
rect 292822 437818 293004 438054
rect 292404 437734 293004 437818
rect 292404 437498 292586 437734
rect 292822 437498 293004 437734
rect 292404 402054 293004 437498
rect 292404 401818 292586 402054
rect 292822 401818 293004 402054
rect 292404 401734 293004 401818
rect 292404 401498 292586 401734
rect 292822 401498 293004 401734
rect 292404 366054 293004 401498
rect 292404 365818 292586 366054
rect 292822 365818 293004 366054
rect 292404 365734 293004 365818
rect 292404 365498 292586 365734
rect 292822 365498 293004 365734
rect 292404 330054 293004 365498
rect 292404 329818 292586 330054
rect 292822 329818 293004 330054
rect 292404 329734 293004 329818
rect 292404 329498 292586 329734
rect 292822 329498 293004 329734
rect 292404 294054 293004 329498
rect 292404 293818 292586 294054
rect 292822 293818 293004 294054
rect 292404 293734 293004 293818
rect 292404 293498 292586 293734
rect 292822 293498 293004 293734
rect 292404 258054 293004 293498
rect 292404 257818 292586 258054
rect 292822 257818 293004 258054
rect 292404 257734 293004 257818
rect 292404 257498 292586 257734
rect 292822 257498 293004 257734
rect 292404 222054 293004 257498
rect 292404 221818 292586 222054
rect 292822 221818 293004 222054
rect 292404 221734 293004 221818
rect 292404 221498 292586 221734
rect 292822 221498 293004 221734
rect 292404 186054 293004 221498
rect 292404 185818 292586 186054
rect 292822 185818 293004 186054
rect 292404 185734 293004 185818
rect 292404 185498 292586 185734
rect 292822 185498 293004 185734
rect 292404 150054 293004 185498
rect 292404 149818 292586 150054
rect 292822 149818 293004 150054
rect 292404 149734 293004 149818
rect 292404 149498 292586 149734
rect 292822 149498 293004 149734
rect 292404 114054 293004 149498
rect 292404 113818 292586 114054
rect 292822 113818 293004 114054
rect 292404 113734 293004 113818
rect 292404 113498 292586 113734
rect 292822 113498 293004 113734
rect 292404 78054 293004 113498
rect 292404 77818 292586 78054
rect 292822 77818 293004 78054
rect 292404 77734 293004 77818
rect 292404 77498 292586 77734
rect 292822 77498 293004 77734
rect 292404 42054 293004 77498
rect 292404 41818 292586 42054
rect 292822 41818 293004 42054
rect 292404 41734 293004 41818
rect 292404 41498 292586 41734
rect 292822 41498 293004 41734
rect 292404 6054 293004 41498
rect 292404 5818 292586 6054
rect 292822 5818 293004 6054
rect 292404 5734 293004 5818
rect 292404 5498 292586 5734
rect 292822 5498 293004 5734
rect 292404 -2226 293004 5498
rect 292404 -2462 292586 -2226
rect 292822 -2462 293004 -2226
rect 292404 -2546 293004 -2462
rect 292404 -2782 292586 -2546
rect 292822 -2782 293004 -2546
rect 292404 -3744 293004 -2782
rect 296004 693654 296604 708042
rect 296004 693418 296186 693654
rect 296422 693418 296604 693654
rect 296004 693334 296604 693418
rect 296004 693098 296186 693334
rect 296422 693098 296604 693334
rect 296004 657654 296604 693098
rect 299604 697254 300204 709922
rect 317604 711418 318204 711440
rect 317604 711182 317786 711418
rect 318022 711182 318204 711418
rect 317604 711098 318204 711182
rect 317604 710862 317786 711098
rect 318022 710862 318204 711098
rect 314004 709538 314604 709560
rect 314004 709302 314186 709538
rect 314422 709302 314604 709538
rect 314004 709218 314604 709302
rect 314004 708982 314186 709218
rect 314422 708982 314604 709218
rect 310404 707658 311004 707680
rect 310404 707422 310586 707658
rect 310822 707422 311004 707658
rect 310404 707338 311004 707422
rect 310404 707102 310586 707338
rect 310822 707102 311004 707338
rect 299604 697018 299786 697254
rect 300022 697018 300204 697254
rect 299604 696934 300204 697018
rect 299604 696698 299786 696934
rect 300022 696698 300204 696934
rect 299427 686220 299493 686221
rect 299427 686156 299428 686220
rect 299492 686156 299493 686220
rect 299427 686155 299493 686156
rect 299430 685949 299490 686155
rect 299427 685948 299493 685949
rect 299427 685884 299428 685948
rect 299492 685884 299493 685948
rect 299427 685883 299493 685884
rect 299427 673844 299493 673845
rect 299427 673780 299428 673844
rect 299492 673780 299493 673844
rect 299427 673779 299493 673780
rect 299430 673573 299490 673779
rect 299427 673572 299493 673573
rect 299427 673508 299428 673572
rect 299492 673508 299493 673572
rect 299427 673507 299493 673508
rect 296004 657418 296186 657654
rect 296422 657418 296604 657654
rect 296004 657334 296604 657418
rect 296004 657098 296186 657334
rect 296422 657098 296604 657334
rect 296004 621654 296604 657098
rect 299604 661254 300204 696698
rect 299604 661018 299786 661254
rect 300022 661018 300204 661254
rect 299604 660934 300204 661018
rect 299604 660698 299786 660934
rect 300022 660698 300204 660934
rect 299427 650724 299493 650725
rect 299427 650660 299428 650724
rect 299492 650660 299493 650724
rect 299427 650659 299493 650660
rect 299430 650453 299490 650659
rect 299427 650452 299493 650453
rect 299427 650388 299428 650452
rect 299492 650388 299493 650452
rect 299427 650387 299493 650388
rect 296004 621418 296186 621654
rect 296422 621418 296604 621654
rect 296004 621334 296604 621418
rect 296004 621098 296186 621334
rect 296422 621098 296604 621334
rect 296004 585654 296604 621098
rect 296004 585418 296186 585654
rect 296422 585418 296604 585654
rect 296004 585334 296604 585418
rect 296004 585098 296186 585334
rect 296422 585098 296604 585334
rect 296004 549654 296604 585098
rect 296004 549418 296186 549654
rect 296422 549418 296604 549654
rect 296004 549334 296604 549418
rect 296004 549098 296186 549334
rect 296422 549098 296604 549334
rect 296004 513654 296604 549098
rect 296004 513418 296186 513654
rect 296422 513418 296604 513654
rect 296004 513334 296604 513418
rect 296004 513098 296186 513334
rect 296422 513098 296604 513334
rect 296004 477654 296604 513098
rect 296004 477418 296186 477654
rect 296422 477418 296604 477654
rect 296004 477334 296604 477418
rect 296004 477098 296186 477334
rect 296422 477098 296604 477334
rect 296004 441654 296604 477098
rect 296004 441418 296186 441654
rect 296422 441418 296604 441654
rect 296004 441334 296604 441418
rect 296004 441098 296186 441334
rect 296422 441098 296604 441334
rect 296004 405654 296604 441098
rect 296004 405418 296186 405654
rect 296422 405418 296604 405654
rect 296004 405334 296604 405418
rect 296004 405098 296186 405334
rect 296422 405098 296604 405334
rect 296004 369654 296604 405098
rect 296004 369418 296186 369654
rect 296422 369418 296604 369654
rect 296004 369334 296604 369418
rect 296004 369098 296186 369334
rect 296422 369098 296604 369334
rect 296004 333654 296604 369098
rect 296004 333418 296186 333654
rect 296422 333418 296604 333654
rect 296004 333334 296604 333418
rect 296004 333098 296186 333334
rect 296422 333098 296604 333334
rect 296004 297654 296604 333098
rect 296004 297418 296186 297654
rect 296422 297418 296604 297654
rect 296004 297334 296604 297418
rect 296004 297098 296186 297334
rect 296422 297098 296604 297334
rect 296004 261654 296604 297098
rect 296004 261418 296186 261654
rect 296422 261418 296604 261654
rect 296004 261334 296604 261418
rect 296004 261098 296186 261334
rect 296422 261098 296604 261334
rect 296004 225654 296604 261098
rect 296004 225418 296186 225654
rect 296422 225418 296604 225654
rect 296004 225334 296604 225418
rect 296004 225098 296186 225334
rect 296422 225098 296604 225334
rect 296004 189654 296604 225098
rect 296004 189418 296186 189654
rect 296422 189418 296604 189654
rect 296004 189334 296604 189418
rect 296004 189098 296186 189334
rect 296422 189098 296604 189334
rect 296004 153654 296604 189098
rect 296004 153418 296186 153654
rect 296422 153418 296604 153654
rect 296004 153334 296604 153418
rect 296004 153098 296186 153334
rect 296422 153098 296604 153334
rect 296004 117654 296604 153098
rect 296004 117418 296186 117654
rect 296422 117418 296604 117654
rect 296004 117334 296604 117418
rect 296004 117098 296186 117334
rect 296422 117098 296604 117334
rect 296004 81654 296604 117098
rect 296004 81418 296186 81654
rect 296422 81418 296604 81654
rect 296004 81334 296604 81418
rect 296004 81098 296186 81334
rect 296422 81098 296604 81334
rect 296004 45654 296604 81098
rect 296004 45418 296186 45654
rect 296422 45418 296604 45654
rect 296004 45334 296604 45418
rect 296004 45098 296186 45334
rect 296422 45098 296604 45334
rect 296004 9654 296604 45098
rect 296004 9418 296186 9654
rect 296422 9418 296604 9654
rect 296004 9334 296604 9418
rect 296004 9098 296186 9334
rect 296422 9098 296604 9334
rect 296004 -4106 296604 9098
rect 296004 -4342 296186 -4106
rect 296422 -4342 296604 -4106
rect 296004 -4426 296604 -4342
rect 296004 -4662 296186 -4426
rect 296422 -4662 296604 -4426
rect 296004 -5624 296604 -4662
rect 299604 625254 300204 660698
rect 306804 705778 307404 705800
rect 306804 705542 306986 705778
rect 307222 705542 307404 705778
rect 306804 705458 307404 705542
rect 306804 705222 306986 705458
rect 307222 705222 307404 705458
rect 306804 668454 307404 705222
rect 306804 668218 306986 668454
rect 307222 668218 307404 668454
rect 306804 668134 307404 668218
rect 306804 667898 306986 668134
rect 307222 667898 307404 668134
rect 306804 654247 307404 667898
rect 310404 672054 311004 707102
rect 310404 671818 310586 672054
rect 310822 671818 311004 672054
rect 310404 671734 311004 671818
rect 310404 671498 310586 671734
rect 310822 671498 311004 671734
rect 310404 654247 311004 671498
rect 314004 675654 314604 708982
rect 314004 675418 314186 675654
rect 314422 675418 314604 675654
rect 314004 675334 314604 675418
rect 314004 675098 314186 675334
rect 314422 675098 314604 675334
rect 314004 654247 314604 675098
rect 317604 679254 318204 710862
rect 335604 710478 336204 711440
rect 335604 710242 335786 710478
rect 336022 710242 336204 710478
rect 335604 710158 336204 710242
rect 335604 709922 335786 710158
rect 336022 709922 336204 710158
rect 332004 708598 332604 709560
rect 332004 708362 332186 708598
rect 332422 708362 332604 708598
rect 332004 708278 332604 708362
rect 332004 708042 332186 708278
rect 332422 708042 332604 708278
rect 328404 706718 329004 707680
rect 328404 706482 328586 706718
rect 328822 706482 329004 706718
rect 328404 706398 329004 706482
rect 328404 706162 328586 706398
rect 328822 706162 329004 706398
rect 317604 679018 317786 679254
rect 318022 679018 318204 679254
rect 317604 678934 318204 679018
rect 317604 678698 317786 678934
rect 318022 678698 318204 678934
rect 317604 654247 318204 678698
rect 324804 704838 325404 705800
rect 324804 704602 324986 704838
rect 325222 704602 325404 704838
rect 324804 704518 325404 704602
rect 324804 704282 324986 704518
rect 325222 704282 325404 704518
rect 324804 686454 325404 704282
rect 324804 686218 324986 686454
rect 325222 686218 325404 686454
rect 324804 686134 325404 686218
rect 324804 685898 324986 686134
rect 325222 685898 325404 686134
rect 324804 654247 325404 685898
rect 328404 690054 329004 706162
rect 328404 689818 328586 690054
rect 328822 689818 329004 690054
rect 328404 689734 329004 689818
rect 328404 689498 328586 689734
rect 328822 689498 329004 689734
rect 328404 654247 329004 689498
rect 332004 693654 332604 708042
rect 332004 693418 332186 693654
rect 332422 693418 332604 693654
rect 332004 693334 332604 693418
rect 332004 693098 332186 693334
rect 332422 693098 332604 693334
rect 332004 657654 332604 693098
rect 332004 657418 332186 657654
rect 332422 657418 332604 657654
rect 332004 657334 332604 657418
rect 332004 657098 332186 657334
rect 332422 657098 332604 657334
rect 332004 654247 332604 657098
rect 335604 697254 336204 709922
rect 353604 711418 354204 711440
rect 353604 711182 353786 711418
rect 354022 711182 354204 711418
rect 353604 711098 354204 711182
rect 353604 710862 353786 711098
rect 354022 710862 354204 711098
rect 350004 709538 350604 709560
rect 350004 709302 350186 709538
rect 350422 709302 350604 709538
rect 350004 709218 350604 709302
rect 350004 708982 350186 709218
rect 350422 708982 350604 709218
rect 346404 707658 347004 707680
rect 346404 707422 346586 707658
rect 346822 707422 347004 707658
rect 346404 707338 347004 707422
rect 346404 707102 346586 707338
rect 346822 707102 347004 707338
rect 335604 697018 335786 697254
rect 336022 697018 336204 697254
rect 335604 696934 336204 697018
rect 335604 696698 335786 696934
rect 336022 696698 336204 696934
rect 335604 661254 336204 696698
rect 335604 661018 335786 661254
rect 336022 661018 336204 661254
rect 335604 660934 336204 661018
rect 335604 660698 335786 660934
rect 336022 660698 336204 660934
rect 335604 654247 336204 660698
rect 342804 705778 343404 705800
rect 342804 705542 342986 705778
rect 343222 705542 343404 705778
rect 342804 705458 343404 705542
rect 342804 705222 342986 705458
rect 343222 705222 343404 705458
rect 342804 668454 343404 705222
rect 342804 668218 342986 668454
rect 343222 668218 343404 668454
rect 342804 668134 343404 668218
rect 342804 667898 342986 668134
rect 343222 667898 343404 668134
rect 342804 654247 343404 667898
rect 346404 672054 347004 707102
rect 346404 671818 346586 672054
rect 346822 671818 347004 672054
rect 346404 671734 347004 671818
rect 346404 671498 346586 671734
rect 346822 671498 347004 671734
rect 346404 654247 347004 671498
rect 350004 675654 350604 708982
rect 350004 675418 350186 675654
rect 350422 675418 350604 675654
rect 350004 675334 350604 675418
rect 350004 675098 350186 675334
rect 350422 675098 350604 675334
rect 350004 654247 350604 675098
rect 353604 679254 354204 710862
rect 371604 710478 372204 711440
rect 371604 710242 371786 710478
rect 372022 710242 372204 710478
rect 371604 710158 372204 710242
rect 371604 709922 371786 710158
rect 372022 709922 372204 710158
rect 368004 708598 368604 709560
rect 368004 708362 368186 708598
rect 368422 708362 368604 708598
rect 368004 708278 368604 708362
rect 368004 708042 368186 708278
rect 368422 708042 368604 708278
rect 364404 706718 365004 707680
rect 364404 706482 364586 706718
rect 364822 706482 365004 706718
rect 364404 706398 365004 706482
rect 364404 706162 364586 706398
rect 364822 706162 365004 706398
rect 360804 704838 361404 705800
rect 360804 704602 360986 704838
rect 361222 704602 361404 704838
rect 360804 704518 361404 704602
rect 360804 704282 360986 704518
rect 361222 704282 361404 704518
rect 360804 686454 361404 704282
rect 357387 686356 357453 686357
rect 357387 686292 357388 686356
rect 357452 686292 357453 686356
rect 357387 686291 357453 686292
rect 357390 685949 357450 686291
rect 360804 686218 360986 686454
rect 361222 686218 361404 686454
rect 360804 686134 361404 686218
rect 357387 685948 357453 685949
rect 357387 685884 357388 685948
rect 357452 685884 357453 685948
rect 357387 685883 357453 685884
rect 360804 685898 360986 686134
rect 361222 685898 361404 686134
rect 353604 679018 353786 679254
rect 354022 679018 354204 679254
rect 353604 678934 354204 679018
rect 353604 678698 353786 678934
rect 354022 678698 354204 678934
rect 353604 654247 354204 678698
rect 357387 673980 357453 673981
rect 357387 673916 357388 673980
rect 357452 673916 357453 673980
rect 357387 673915 357453 673916
rect 357390 673573 357450 673915
rect 357387 673572 357453 673573
rect 357387 673508 357388 673572
rect 357452 673508 357453 673572
rect 357387 673507 357453 673508
rect 360804 654247 361404 685898
rect 364404 690054 365004 706162
rect 364404 689818 364586 690054
rect 364822 689818 365004 690054
rect 364404 689734 365004 689818
rect 364404 689498 364586 689734
rect 364822 689498 365004 689734
rect 364404 654247 365004 689498
rect 368004 693654 368604 708042
rect 368004 693418 368186 693654
rect 368422 693418 368604 693654
rect 368004 693334 368604 693418
rect 368004 693098 368186 693334
rect 368422 693098 368604 693334
rect 368004 657654 368604 693098
rect 368004 657418 368186 657654
rect 368422 657418 368604 657654
rect 368004 657334 368604 657418
rect 368004 657098 368186 657334
rect 368422 657098 368604 657334
rect 368004 654247 368604 657098
rect 371604 697254 372204 709922
rect 389604 711418 390204 711440
rect 389604 711182 389786 711418
rect 390022 711182 390204 711418
rect 389604 711098 390204 711182
rect 389604 710862 389786 711098
rect 390022 710862 390204 711098
rect 386004 709538 386604 709560
rect 386004 709302 386186 709538
rect 386422 709302 386604 709538
rect 386004 709218 386604 709302
rect 386004 708982 386186 709218
rect 386422 708982 386604 709218
rect 382404 707658 383004 707680
rect 382404 707422 382586 707658
rect 382822 707422 383004 707658
rect 382404 707338 383004 707422
rect 382404 707102 382586 707338
rect 382822 707102 383004 707338
rect 371604 697018 371786 697254
rect 372022 697018 372204 697254
rect 371604 696934 372204 697018
rect 371604 696698 371786 696934
rect 372022 696698 372204 696934
rect 371604 661254 372204 696698
rect 378804 705778 379404 705800
rect 378804 705542 378986 705778
rect 379222 705542 379404 705778
rect 378804 705458 379404 705542
rect 378804 705222 378986 705458
rect 379222 705222 379404 705458
rect 376707 686492 376773 686493
rect 376707 686428 376708 686492
rect 376772 686428 376773 686492
rect 376707 686427 376773 686428
rect 376710 686221 376770 686427
rect 376707 686220 376773 686221
rect 376707 686156 376708 686220
rect 376772 686156 376773 686220
rect 376707 686155 376773 686156
rect 376707 674116 376773 674117
rect 376707 674052 376708 674116
rect 376772 674052 376773 674116
rect 376707 674051 376773 674052
rect 376710 673845 376770 674051
rect 376707 673844 376773 673845
rect 376707 673780 376708 673844
rect 376772 673780 376773 673844
rect 376707 673779 376773 673780
rect 371604 661018 371786 661254
rect 372022 661018 372204 661254
rect 371604 660934 372204 661018
rect 371604 660698 371786 660934
rect 372022 660698 372204 660934
rect 371604 654247 372204 660698
rect 378804 668454 379404 705222
rect 378804 668218 378986 668454
rect 379222 668218 379404 668454
rect 378804 668134 379404 668218
rect 378804 667898 378986 668134
rect 379222 667898 379404 668134
rect 378804 654247 379404 667898
rect 382404 672054 383004 707102
rect 382404 671818 382586 672054
rect 382822 671818 383004 672054
rect 382404 671734 383004 671818
rect 382404 671498 382586 671734
rect 382822 671498 383004 671734
rect 382404 654247 383004 671498
rect 386004 675654 386604 708982
rect 386004 675418 386186 675654
rect 386422 675418 386604 675654
rect 386004 675334 386604 675418
rect 386004 675098 386186 675334
rect 386422 675098 386604 675334
rect 386004 654247 386604 675098
rect 389604 679254 390204 710862
rect 407604 710478 408204 711440
rect 407604 710242 407786 710478
rect 408022 710242 408204 710478
rect 407604 710158 408204 710242
rect 407604 709922 407786 710158
rect 408022 709922 408204 710158
rect 404004 708598 404604 709560
rect 404004 708362 404186 708598
rect 404422 708362 404604 708598
rect 404004 708278 404604 708362
rect 404004 708042 404186 708278
rect 404422 708042 404604 708278
rect 400404 706718 401004 707680
rect 400404 706482 400586 706718
rect 400822 706482 401004 706718
rect 400404 706398 401004 706482
rect 400404 706162 400586 706398
rect 400822 706162 401004 706398
rect 389604 679018 389786 679254
rect 390022 679018 390204 679254
rect 389604 678934 390204 679018
rect 389604 678698 389786 678934
rect 390022 678698 390204 678934
rect 389604 654247 390204 678698
rect 396804 704838 397404 705800
rect 396804 704602 396986 704838
rect 397222 704602 397404 704838
rect 396804 704518 397404 704602
rect 396804 704282 396986 704518
rect 397222 704282 397404 704518
rect 396804 686454 397404 704282
rect 396804 686218 396986 686454
rect 397222 686218 397404 686454
rect 396804 686134 397404 686218
rect 396804 685898 396986 686134
rect 397222 685898 397404 686134
rect 378179 652900 378245 652901
rect 378179 652836 378180 652900
rect 378244 652836 378245 652900
rect 378179 652835 378245 652836
rect 383515 652900 383581 652901
rect 383515 652836 383516 652900
rect 383580 652836 383581 652900
rect 383515 652835 383581 652836
rect 376707 651404 376773 651405
rect 376707 651340 376708 651404
rect 376772 651340 376773 651404
rect 376707 651339 376773 651340
rect 376710 651133 376770 651339
rect 376707 651132 376773 651133
rect 376707 651068 376708 651132
rect 376772 651068 376773 651132
rect 378182 651130 378242 652835
rect 383518 651130 383578 652835
rect 396027 651132 396093 651133
rect 378182 651070 378608 651130
rect 383518 651070 383603 651130
rect 376707 651067 376773 651068
rect 396027 651068 396028 651132
rect 396092 651068 396093 651132
rect 396027 651067 396093 651068
rect 318747 650996 318813 650997
rect 318747 650932 318748 650996
rect 318812 650932 318813 650996
rect 318747 650931 318813 650932
rect 318750 650589 318810 650931
rect 396030 650861 396090 651067
rect 396027 650860 396093 650861
rect 396027 650796 396028 650860
rect 396092 650796 396093 650860
rect 396027 650795 396093 650796
rect 318747 650588 318813 650589
rect 318747 650524 318748 650588
rect 318812 650524 318813 650588
rect 318747 650523 318813 650524
rect 396804 650454 397404 685898
rect 396804 650218 396986 650454
rect 397222 650218 397404 650454
rect 396804 650134 397404 650218
rect 396804 649898 396986 650134
rect 397222 649898 397404 650134
rect 386938 643254 387262 643276
rect 386938 643018 386982 643254
rect 387218 643018 387262 643254
rect 386938 642934 387262 643018
rect 386938 642698 386982 642934
rect 387218 642698 387262 642934
rect 386938 642676 387262 642698
rect 386938 639654 387262 639676
rect 386938 639418 386982 639654
rect 387218 639418 387262 639654
rect 386938 639334 387262 639418
rect 386938 639098 386982 639334
rect 387218 639098 387262 639334
rect 386938 639076 387262 639098
rect 386938 636054 387262 636076
rect 386938 635818 386982 636054
rect 387218 635818 387262 636054
rect 386938 635734 387262 635818
rect 386938 635498 386982 635734
rect 387218 635498 387262 635734
rect 386938 635476 387262 635498
rect 386938 632454 387262 632476
rect 386938 632218 386982 632454
rect 387218 632218 387262 632454
rect 386938 632134 387262 632218
rect 386938 631898 386982 632134
rect 387218 631898 387262 632134
rect 386938 631876 387262 631898
rect 299604 625018 299786 625254
rect 300022 625018 300204 625254
rect 299604 624934 300204 625018
rect 299604 624698 299786 624934
rect 300022 624698 300204 624934
rect 299604 589254 300204 624698
rect 386494 625254 386814 625276
rect 386494 625018 386536 625254
rect 386772 625018 386814 625254
rect 386494 624934 386814 625018
rect 386494 624698 386536 624934
rect 386772 624698 386814 624934
rect 386494 624676 386814 624698
rect 386494 621654 386814 621676
rect 386494 621418 386536 621654
rect 386772 621418 386814 621654
rect 386494 621334 386814 621418
rect 386494 621098 386536 621334
rect 386772 621098 386814 621334
rect 386494 621076 386814 621098
rect 386494 618054 386814 618076
rect 386494 617818 386536 618054
rect 386772 617818 386814 618054
rect 386494 617734 386814 617818
rect 386494 617498 386536 617734
rect 386772 617498 386814 617734
rect 386494 617476 386814 617498
rect 386494 614454 386814 614476
rect 386494 614218 386536 614454
rect 386772 614218 386814 614454
rect 386494 614134 386814 614218
rect 386494 613898 386536 614134
rect 386772 613898 386814 614134
rect 386494 613876 386814 613898
rect 396804 614454 397404 649898
rect 396804 614218 396986 614454
rect 397222 614218 397404 614454
rect 396804 614134 397404 614218
rect 396804 613898 396986 614134
rect 397222 613898 397404 614134
rect 386938 607254 387262 607276
rect 386938 607018 386982 607254
rect 387218 607018 387262 607254
rect 386938 606934 387262 607018
rect 386938 606698 386982 606934
rect 387218 606698 387262 606934
rect 386938 606676 387262 606698
rect 386938 603654 387262 603676
rect 386938 603418 386982 603654
rect 387218 603418 387262 603654
rect 386938 603334 387262 603418
rect 386938 603098 386982 603334
rect 387218 603098 387262 603334
rect 386938 603076 387262 603098
rect 386938 600054 387262 600076
rect 386938 599818 386982 600054
rect 387218 599818 387262 600054
rect 386938 599734 387262 599818
rect 386938 599498 386982 599734
rect 387218 599498 387262 599734
rect 386938 599476 387262 599498
rect 386938 596454 387262 596476
rect 386938 596218 386982 596454
rect 387218 596218 387262 596454
rect 386938 596134 387262 596218
rect 386938 595898 386982 596134
rect 387218 595898 387262 596134
rect 386938 595876 387262 595898
rect 299604 589018 299786 589254
rect 300022 589018 300204 589254
rect 299604 588934 300204 589018
rect 299604 588698 299786 588934
rect 300022 588698 300204 588934
rect 299604 553254 300204 588698
rect 386494 589254 386814 589276
rect 386494 589018 386536 589254
rect 386772 589018 386814 589254
rect 386494 588934 386814 589018
rect 386494 588698 386536 588934
rect 386772 588698 386814 588934
rect 386494 588676 386814 588698
rect 386494 585654 386814 585676
rect 386494 585418 386536 585654
rect 386772 585418 386814 585654
rect 386494 585334 386814 585418
rect 386494 585098 386536 585334
rect 386772 585098 386814 585334
rect 386494 585076 386814 585098
rect 386494 582054 386814 582076
rect 386494 581818 386536 582054
rect 386772 581818 386814 582054
rect 386494 581734 386814 581818
rect 386494 581498 386536 581734
rect 386772 581498 386814 581734
rect 386494 581476 386814 581498
rect 386494 578454 386814 578476
rect 386494 578218 386536 578454
rect 386772 578218 386814 578454
rect 386494 578134 386814 578218
rect 386494 577898 386536 578134
rect 386772 577898 386814 578134
rect 386494 577876 386814 577898
rect 396804 578454 397404 613898
rect 396804 578218 396986 578454
rect 397222 578218 397404 578454
rect 396804 578134 397404 578218
rect 396804 577898 396986 578134
rect 397222 577898 397404 578134
rect 386938 571254 387262 571276
rect 386938 571018 386982 571254
rect 387218 571018 387262 571254
rect 386938 570934 387262 571018
rect 386938 570698 386982 570934
rect 387218 570698 387262 570934
rect 386938 570676 387262 570698
rect 386938 567654 387262 567676
rect 386938 567418 386982 567654
rect 387218 567418 387262 567654
rect 386938 567334 387262 567418
rect 386938 567098 386982 567334
rect 387218 567098 387262 567334
rect 386938 567076 387262 567098
rect 386938 564054 387262 564076
rect 386938 563818 386982 564054
rect 387218 563818 387262 564054
rect 386938 563734 387262 563818
rect 386938 563498 386982 563734
rect 387218 563498 387262 563734
rect 386938 563476 387262 563498
rect 359004 560630 359474 560690
rect 320336 560430 320650 560490
rect 313414 560290 313833 560350
rect 316358 560290 316832 560350
rect 317462 560290 318000 560350
rect 318934 560290 319168 560350
rect 313414 558925 313474 560290
rect 313411 558924 313477 558925
rect 313411 558860 313412 558924
rect 313476 558860 313477 558924
rect 313411 558859 313477 558860
rect 316358 557565 316418 560290
rect 317462 557973 317522 560290
rect 317459 557972 317525 557973
rect 317459 557908 317460 557972
rect 317524 557908 317525 557972
rect 317459 557907 317525 557908
rect 318934 557565 318994 560290
rect 320590 557973 320650 560430
rect 323534 560430 323840 560490
rect 327030 560430 327344 560490
rect 328636 560430 328930 560490
rect 320958 560290 321504 560350
rect 322246 560290 322672 560350
rect 322796 560290 322858 560350
rect 320587 557972 320653 557973
rect 320587 557908 320588 557972
rect 320652 557908 320653 557972
rect 320587 557907 320653 557908
rect 320958 557565 321018 560290
rect 322246 558789 322306 560290
rect 322798 558925 322858 560290
rect 322795 558924 322861 558925
rect 322795 558860 322796 558924
rect 322860 558860 322861 558924
rect 322795 558859 322861 558860
rect 323534 558789 323594 560430
rect 323964 560290 324146 560350
rect 324086 558925 324146 560290
rect 324822 560290 325008 560350
rect 324083 558924 324149 558925
rect 324083 558860 324084 558924
rect 324148 558860 324149 558924
rect 324083 558859 324149 558860
rect 324822 558789 324882 560290
rect 325102 560010 325162 560320
rect 326110 560290 326176 560350
rect 325102 559950 325250 560010
rect 325190 558925 325250 559950
rect 325187 558924 325253 558925
rect 325187 558860 325188 558924
rect 325252 558860 325253 558924
rect 325187 558859 325253 558860
rect 326110 558789 326170 560290
rect 326294 558925 326354 560350
rect 326291 558924 326357 558925
rect 326291 558860 326292 558924
rect 326356 558860 326357 558924
rect 326291 558859 326357 558860
rect 327030 558789 327090 560430
rect 327468 560290 327642 560350
rect 327582 558925 327642 560290
rect 328482 559877 328542 560320
rect 328479 559876 328545 559877
rect 328479 559812 328480 559876
rect 328544 559812 328545 559876
rect 328479 559811 328545 559812
rect 327579 558924 327645 558925
rect 327579 558860 327580 558924
rect 327644 558860 327645 558924
rect 327579 558859 327645 558860
rect 322243 558788 322309 558789
rect 322243 558724 322244 558788
rect 322308 558724 322309 558788
rect 322243 558723 322309 558724
rect 323531 558788 323597 558789
rect 323531 558724 323532 558788
rect 323596 558724 323597 558788
rect 323531 558723 323597 558724
rect 324819 558788 324885 558789
rect 324819 558724 324820 558788
rect 324884 558724 324885 558788
rect 324819 558723 324885 558724
rect 326107 558788 326173 558789
rect 326107 558724 326108 558788
rect 326172 558724 326173 558788
rect 326107 558723 326173 558724
rect 327027 558788 327093 558789
rect 327027 558724 327028 558788
rect 327092 558724 327093 558788
rect 327027 558723 327093 558724
rect 316355 557564 316421 557565
rect 316355 557500 316356 557564
rect 316420 557500 316421 557564
rect 316355 557499 316421 557500
rect 318931 557564 318997 557565
rect 318931 557500 318932 557564
rect 318996 557500 318997 557564
rect 318931 557499 318997 557500
rect 320955 557564 321021 557565
rect 320955 557500 320956 557564
rect 321020 557500 321021 557564
rect 320955 557499 321021 557500
rect 328870 557157 328930 560430
rect 330526 560430 330848 560490
rect 332140 560430 332426 560490
rect 329606 560290 329680 560350
rect 329606 558925 329666 560290
rect 329790 558925 329850 560350
rect 330526 558925 330586 560430
rect 330972 560290 331138 560350
rect 329603 558924 329669 558925
rect 329603 558860 329604 558924
rect 329668 558860 329669 558924
rect 329603 558859 329669 558860
rect 329787 558924 329853 558925
rect 329787 558860 329788 558924
rect 329852 558860 329853 558924
rect 329787 558859 329853 558860
rect 330523 558924 330589 558925
rect 330523 558860 330524 558924
rect 330588 558860 330589 558924
rect 330523 558859 330589 558860
rect 331078 558789 331138 560290
rect 331814 560290 332016 560350
rect 331814 558789 331874 560290
rect 332366 558925 332426 560430
rect 334022 560430 334352 560490
rect 335644 560430 335922 560490
rect 332734 560290 333184 560350
rect 332363 558924 332429 558925
rect 332363 558860 332364 558924
rect 332428 558860 332429 558924
rect 332363 558859 332429 558860
rect 332734 558789 332794 560290
rect 333286 558925 333346 560350
rect 333283 558924 333349 558925
rect 333283 558860 333284 558924
rect 333348 558860 333349 558924
rect 333283 558859 333349 558860
rect 334022 558789 334082 560430
rect 334476 560290 334634 560350
rect 334574 558925 334634 560290
rect 335490 560010 335550 560320
rect 335490 559950 335554 560010
rect 334571 558924 334637 558925
rect 334571 558860 334572 558924
rect 334636 558860 334637 558924
rect 334571 558859 334637 558860
rect 335494 558789 335554 559950
rect 335862 558925 335922 560430
rect 339910 560430 340192 560490
rect 341484 560430 341810 560490
rect 336598 560290 336688 560350
rect 335859 558924 335925 558925
rect 335859 558860 335860 558924
rect 335924 558860 335925 558924
rect 335859 558859 335925 558860
rect 336598 558789 336658 560290
rect 336782 558925 336842 560320
rect 337702 560290 337856 560350
rect 337702 559877 337762 560290
rect 337699 559876 337765 559877
rect 337699 559812 337700 559876
rect 337764 559812 337765 559876
rect 337699 559811 337765 559812
rect 337950 559330 338010 560320
rect 337886 559270 338010 559330
rect 336779 558924 336845 558925
rect 336779 558860 336780 558924
rect 336844 558860 336845 558924
rect 336779 558859 336845 558860
rect 331075 558788 331141 558789
rect 331075 558724 331076 558788
rect 331140 558724 331141 558788
rect 331075 558723 331141 558724
rect 331811 558788 331877 558789
rect 331811 558724 331812 558788
rect 331876 558724 331877 558788
rect 331811 558723 331877 558724
rect 332731 558788 332797 558789
rect 332731 558724 332732 558788
rect 332796 558724 332797 558788
rect 332731 558723 332797 558724
rect 334019 558788 334085 558789
rect 334019 558724 334020 558788
rect 334084 558724 334085 558788
rect 334019 558723 334085 558724
rect 335491 558788 335557 558789
rect 335491 558724 335492 558788
rect 335556 558724 335557 558788
rect 335491 558723 335557 558724
rect 336595 558788 336661 558789
rect 336595 558724 336596 558788
rect 336660 558724 336661 558788
rect 336595 558723 336661 558724
rect 337886 557973 337946 559270
rect 338990 558789 339050 560350
rect 339148 560290 339234 560350
rect 339174 558925 339234 560290
rect 339171 558924 339237 558925
rect 339171 558860 339172 558924
rect 339236 558860 339237 558924
rect 339171 558859 339237 558860
rect 339910 558789 339970 560430
rect 340316 560290 340522 560350
rect 340462 558925 340522 560290
rect 341198 560290 341360 560350
rect 341198 558925 341258 560290
rect 340459 558924 340525 558925
rect 340459 558860 340460 558924
rect 340524 558860 340525 558924
rect 340459 558859 340525 558860
rect 341195 558924 341261 558925
rect 341195 558860 341196 558924
rect 341260 558860 341261 558924
rect 341195 558859 341261 558860
rect 338987 558788 339053 558789
rect 338987 558724 338988 558788
rect 339052 558724 339053 558788
rect 338987 558723 339053 558724
rect 339907 558788 339973 558789
rect 339907 558724 339908 558788
rect 339972 558724 339973 558788
rect 339907 558723 339973 558724
rect 337883 557972 337949 557973
rect 337883 557908 337884 557972
rect 337948 557908 337949 557972
rect 337883 557907 337949 557908
rect 341750 557565 341810 560430
rect 346902 560430 347200 560490
rect 348492 560430 348802 560490
rect 351996 560430 352298 560490
rect 355500 560430 355794 560490
rect 342486 558925 342546 560350
rect 342652 560290 342730 560350
rect 342483 558924 342549 558925
rect 342483 558860 342484 558924
rect 342548 558860 342549 558924
rect 342483 558859 342549 558860
rect 342670 557565 342730 560290
rect 343666 560010 343726 560320
rect 343820 560290 344018 560350
rect 343590 559950 343726 560010
rect 343590 558925 343650 559950
rect 343587 558924 343653 558925
rect 343587 558860 343588 558924
rect 343652 558860 343653 558924
rect 343587 558859 343653 558860
rect 343958 557565 344018 560290
rect 344694 560290 344864 560350
rect 344694 558925 344754 560290
rect 344958 559330 345018 560320
rect 344878 559270 345018 559330
rect 345798 560290 346032 560350
rect 346156 560290 346226 560350
rect 344691 558924 344757 558925
rect 344691 558860 344692 558924
rect 344756 558860 344757 558924
rect 344691 558859 344757 558860
rect 344878 557701 344938 559270
rect 345798 558925 345858 560290
rect 345795 558924 345861 558925
rect 345795 558860 345796 558924
rect 345860 558860 345861 558924
rect 345795 558859 345861 558860
rect 344875 557700 344941 557701
rect 344875 557636 344876 557700
rect 344940 557636 344941 557700
rect 344875 557635 344941 557636
rect 346166 557565 346226 560290
rect 346902 558925 346962 560430
rect 347324 560290 347514 560350
rect 346899 558924 346965 558925
rect 346899 558860 346900 558924
rect 346964 558860 346965 558924
rect 346899 558859 346965 558860
rect 347454 557565 347514 560290
rect 348190 560290 348368 560350
rect 348190 558925 348250 560290
rect 348187 558924 348253 558925
rect 348187 558860 348188 558924
rect 348252 558860 348253 558924
rect 348187 558859 348253 558860
rect 348742 557565 348802 560430
rect 349478 558925 349538 560350
rect 349660 560290 349722 560350
rect 349475 558924 349541 558925
rect 349475 558860 349476 558924
rect 349540 558860 349541 558924
rect 349475 558859 349541 558860
rect 349662 557565 349722 560290
rect 350674 560010 350734 560320
rect 350828 560290 351010 560350
rect 350582 559950 350734 560010
rect 350582 558517 350642 559950
rect 350579 558516 350645 558517
rect 350579 558452 350580 558516
rect 350644 558452 350645 558516
rect 350579 558451 350645 558452
rect 350950 557565 351010 560290
rect 351842 559333 351902 560320
rect 351842 559332 351933 559333
rect 351842 559270 351868 559332
rect 351867 559268 351868 559270
rect 351932 559268 351933 559332
rect 351867 559267 351933 559268
rect 352238 559197 352298 560430
rect 352422 560290 353040 560350
rect 352235 559196 352301 559197
rect 352235 559132 352236 559196
rect 352300 559132 352301 559196
rect 352235 559131 352301 559132
rect 352422 558245 352482 560290
rect 352419 558244 352485 558245
rect 352419 558180 352420 558244
rect 352484 558180 352485 558244
rect 352419 558179 352485 558180
rect 353158 558109 353218 560350
rect 353526 560290 354208 560350
rect 354332 560290 354506 560350
rect 353526 558789 353586 560290
rect 353523 558788 353589 558789
rect 353523 558724 353524 558788
rect 353588 558724 353589 558788
rect 353523 558723 353589 558724
rect 353155 558108 353221 558109
rect 353155 558044 353156 558108
rect 353220 558044 353221 558108
rect 353155 558043 353221 558044
rect 354446 557973 354506 560290
rect 354814 560290 355376 560350
rect 354814 558789 354874 560290
rect 354811 558788 354877 558789
rect 354811 558724 354812 558788
rect 354876 558724 354877 558788
rect 354811 558723 354877 558724
rect 355734 558245 355794 560430
rect 356102 560290 356544 560350
rect 356102 558789 356162 560290
rect 356099 558788 356165 558789
rect 356099 558724 356100 558788
rect 356164 558724 356165 558788
rect 356099 558723 356165 558724
rect 355731 558244 355797 558245
rect 355731 558180 355732 558244
rect 355796 558180 355797 558244
rect 355731 558179 355797 558180
rect 354443 557972 354509 557973
rect 354443 557908 354444 557972
rect 354508 557908 354509 557972
rect 354443 557907 354509 557908
rect 356654 557701 356714 560350
rect 357682 560010 357742 560320
rect 357836 560290 358002 560350
rect 357574 559950 357742 560010
rect 357574 558517 357634 559950
rect 357942 558653 358002 560290
rect 358850 559877 358910 560320
rect 358847 559876 358913 559877
rect 358847 559812 358848 559876
rect 358912 559812 358913 559876
rect 358847 559811 358913 559812
rect 359414 559741 359474 560630
rect 358859 559740 358925 559741
rect 358859 559676 358860 559740
rect 358924 559676 358925 559740
rect 358859 559675 358925 559676
rect 359411 559740 359477 559741
rect 359411 559676 359412 559740
rect 359476 559676 359477 559740
rect 359411 559675 359477 559676
rect 358862 558925 358922 559675
rect 358859 558924 358925 558925
rect 358859 558860 358860 558924
rect 358924 558860 358925 558924
rect 358859 558859 358925 558860
rect 357939 558652 358005 558653
rect 357939 558588 357940 558652
rect 358004 558588 358005 558652
rect 357939 558587 358005 558588
rect 357571 558516 357637 558517
rect 357571 558452 357572 558516
rect 357636 558452 357637 558516
rect 357571 558451 357637 558452
rect 356651 557700 356717 557701
rect 356651 557636 356652 557700
rect 356716 557636 356717 557700
rect 356651 557635 356717 557636
rect 341747 557564 341813 557565
rect 341747 557500 341748 557564
rect 341812 557500 341813 557564
rect 341747 557499 341813 557500
rect 342667 557564 342733 557565
rect 342667 557500 342668 557564
rect 342732 557500 342733 557564
rect 342667 557499 342733 557500
rect 343955 557564 344021 557565
rect 343955 557500 343956 557564
rect 344020 557500 344021 557564
rect 343955 557499 344021 557500
rect 346163 557564 346229 557565
rect 346163 557500 346164 557564
rect 346228 557500 346229 557564
rect 346163 557499 346229 557500
rect 347451 557564 347517 557565
rect 347451 557500 347452 557564
rect 347516 557500 347517 557564
rect 347451 557499 347517 557500
rect 348739 557564 348805 557565
rect 348739 557500 348740 557564
rect 348804 557500 348805 557564
rect 348739 557499 348805 557500
rect 349659 557564 349725 557565
rect 349659 557500 349660 557564
rect 349724 557500 349725 557564
rect 349659 557499 349725 557500
rect 350947 557564 351013 557565
rect 350947 557500 350948 557564
rect 351012 557500 351013 557564
rect 350947 557499 351013 557500
rect 328867 557156 328933 557157
rect 328867 557092 328868 557156
rect 328932 557092 328933 557156
rect 328867 557091 328933 557092
rect 299604 553018 299786 553254
rect 300022 553018 300204 553254
rect 299604 552934 300204 553018
rect 299604 552698 299786 552934
rect 300022 552698 300204 552934
rect 299604 517254 300204 552698
rect 299604 517018 299786 517254
rect 300022 517018 300204 517254
rect 299604 516934 300204 517018
rect 299604 516698 299786 516934
rect 300022 516698 300204 516934
rect 299604 481254 300204 516698
rect 299604 481018 299786 481254
rect 300022 481018 300204 481254
rect 299604 480934 300204 481018
rect 299604 480698 299786 480934
rect 300022 480698 300204 480934
rect 299604 445254 300204 480698
rect 299604 445018 299786 445254
rect 300022 445018 300204 445254
rect 299604 444934 300204 445018
rect 299604 444698 299786 444934
rect 300022 444698 300204 444934
rect 299604 409254 300204 444698
rect 299604 409018 299786 409254
rect 300022 409018 300204 409254
rect 299604 408934 300204 409018
rect 299604 408698 299786 408934
rect 300022 408698 300204 408934
rect 299604 373254 300204 408698
rect 299604 373018 299786 373254
rect 300022 373018 300204 373254
rect 299604 372934 300204 373018
rect 299604 372698 299786 372934
rect 300022 372698 300204 372934
rect 299604 337254 300204 372698
rect 299604 337018 299786 337254
rect 300022 337018 300204 337254
rect 299604 336934 300204 337018
rect 299604 336698 299786 336934
rect 300022 336698 300204 336934
rect 299604 301254 300204 336698
rect 299604 301018 299786 301254
rect 300022 301018 300204 301254
rect 299604 300934 300204 301018
rect 299604 300698 299786 300934
rect 300022 300698 300204 300934
rect 299604 265254 300204 300698
rect 299604 265018 299786 265254
rect 300022 265018 300204 265254
rect 299604 264934 300204 265018
rect 299604 264698 299786 264934
rect 300022 264698 300204 264934
rect 299604 229254 300204 264698
rect 299604 229018 299786 229254
rect 300022 229018 300204 229254
rect 299604 228934 300204 229018
rect 299604 228698 299786 228934
rect 300022 228698 300204 228934
rect 299604 193254 300204 228698
rect 299604 193018 299786 193254
rect 300022 193018 300204 193254
rect 299604 192934 300204 193018
rect 299604 192698 299786 192934
rect 300022 192698 300204 192934
rect 299604 157254 300204 192698
rect 299604 157018 299786 157254
rect 300022 157018 300204 157254
rect 299604 156934 300204 157018
rect 299604 156698 299786 156934
rect 300022 156698 300204 156934
rect 299604 121254 300204 156698
rect 299604 121018 299786 121254
rect 300022 121018 300204 121254
rect 299604 120934 300204 121018
rect 299604 120698 299786 120934
rect 300022 120698 300204 120934
rect 299604 85254 300204 120698
rect 299604 85018 299786 85254
rect 300022 85018 300204 85254
rect 299604 84934 300204 85018
rect 299604 84698 299786 84934
rect 300022 84698 300204 84934
rect 299604 49254 300204 84698
rect 299604 49018 299786 49254
rect 300022 49018 300204 49254
rect 299604 48934 300204 49018
rect 299604 48698 299786 48934
rect 300022 48698 300204 48934
rect 299604 13254 300204 48698
rect 299604 13018 299786 13254
rect 300022 13018 300204 13254
rect 299604 12934 300204 13018
rect 299604 12698 299786 12934
rect 300022 12698 300204 12934
rect 281604 -7162 281786 -6926
rect 282022 -7162 282204 -6926
rect 281604 -7246 282204 -7162
rect 281604 -7482 281786 -7246
rect 282022 -7482 282204 -7246
rect 281604 -7504 282204 -7482
rect 299604 -5986 300204 12698
rect 306804 524454 307404 557000
rect 306804 524218 306986 524454
rect 307222 524218 307404 524454
rect 306804 524134 307404 524218
rect 306804 523898 306986 524134
rect 307222 523898 307404 524134
rect 306804 488454 307404 523898
rect 306804 488218 306986 488454
rect 307222 488218 307404 488454
rect 306804 488134 307404 488218
rect 306804 487898 306986 488134
rect 307222 487898 307404 488134
rect 306804 452454 307404 487898
rect 306804 452218 306986 452454
rect 307222 452218 307404 452454
rect 306804 452134 307404 452218
rect 306804 451898 306986 452134
rect 307222 451898 307404 452134
rect 306804 416454 307404 451898
rect 306804 416218 306986 416454
rect 307222 416218 307404 416454
rect 306804 416134 307404 416218
rect 306804 415898 306986 416134
rect 307222 415898 307404 416134
rect 306804 380454 307404 415898
rect 306804 380218 306986 380454
rect 307222 380218 307404 380454
rect 306804 380134 307404 380218
rect 306804 379898 306986 380134
rect 307222 379898 307404 380134
rect 306804 344454 307404 379898
rect 306804 344218 306986 344454
rect 307222 344218 307404 344454
rect 306804 344134 307404 344218
rect 306804 343898 306986 344134
rect 307222 343898 307404 344134
rect 306804 308454 307404 343898
rect 306804 308218 306986 308454
rect 307222 308218 307404 308454
rect 306804 308134 307404 308218
rect 306804 307898 306986 308134
rect 307222 307898 307404 308134
rect 306804 272454 307404 307898
rect 306804 272218 306986 272454
rect 307222 272218 307404 272454
rect 306804 272134 307404 272218
rect 306804 271898 306986 272134
rect 307222 271898 307404 272134
rect 306804 236454 307404 271898
rect 306804 236218 306986 236454
rect 307222 236218 307404 236454
rect 306804 236134 307404 236218
rect 306804 235898 306986 236134
rect 307222 235898 307404 236134
rect 306804 200454 307404 235898
rect 306804 200218 306986 200454
rect 307222 200218 307404 200454
rect 306804 200134 307404 200218
rect 306804 199898 306986 200134
rect 307222 199898 307404 200134
rect 306804 164454 307404 199898
rect 306804 164218 306986 164454
rect 307222 164218 307404 164454
rect 306804 164134 307404 164218
rect 306804 163898 306986 164134
rect 307222 163898 307404 164134
rect 306804 128454 307404 163898
rect 306804 128218 306986 128454
rect 307222 128218 307404 128454
rect 306804 128134 307404 128218
rect 306804 127898 306986 128134
rect 307222 127898 307404 128134
rect 306804 92454 307404 127898
rect 306804 92218 306986 92454
rect 307222 92218 307404 92454
rect 306804 92134 307404 92218
rect 306804 91898 306986 92134
rect 307222 91898 307404 92134
rect 306804 56454 307404 91898
rect 306804 56218 306986 56454
rect 307222 56218 307404 56454
rect 306804 56134 307404 56218
rect 306804 55898 306986 56134
rect 307222 55898 307404 56134
rect 306804 20454 307404 55898
rect 306804 20218 306986 20454
rect 307222 20218 307404 20454
rect 306804 20134 307404 20218
rect 306804 19898 306986 20134
rect 307222 19898 307404 20134
rect 306804 -1286 307404 19898
rect 306804 -1522 306986 -1286
rect 307222 -1522 307404 -1286
rect 306804 -1606 307404 -1522
rect 306804 -1842 306986 -1606
rect 307222 -1842 307404 -1606
rect 306804 -1864 307404 -1842
rect 310404 528054 311004 557000
rect 310404 527818 310586 528054
rect 310822 527818 311004 528054
rect 310404 527734 311004 527818
rect 310404 527498 310586 527734
rect 310822 527498 311004 527734
rect 310404 492054 311004 527498
rect 310404 491818 310586 492054
rect 310822 491818 311004 492054
rect 310404 491734 311004 491818
rect 310404 491498 310586 491734
rect 310822 491498 311004 491734
rect 310404 456054 311004 491498
rect 310404 455818 310586 456054
rect 310822 455818 311004 456054
rect 310404 455734 311004 455818
rect 310404 455498 310586 455734
rect 310822 455498 311004 455734
rect 310404 420054 311004 455498
rect 310404 419818 310586 420054
rect 310822 419818 311004 420054
rect 310404 419734 311004 419818
rect 310404 419498 310586 419734
rect 310822 419498 311004 419734
rect 310404 384054 311004 419498
rect 310404 383818 310586 384054
rect 310822 383818 311004 384054
rect 310404 383734 311004 383818
rect 310404 383498 310586 383734
rect 310822 383498 311004 383734
rect 310404 348054 311004 383498
rect 310404 347818 310586 348054
rect 310822 347818 311004 348054
rect 310404 347734 311004 347818
rect 310404 347498 310586 347734
rect 310822 347498 311004 347734
rect 310404 312054 311004 347498
rect 310404 311818 310586 312054
rect 310822 311818 311004 312054
rect 310404 311734 311004 311818
rect 310404 311498 310586 311734
rect 310822 311498 311004 311734
rect 310404 276054 311004 311498
rect 310404 275818 310586 276054
rect 310822 275818 311004 276054
rect 310404 275734 311004 275818
rect 310404 275498 310586 275734
rect 310822 275498 311004 275734
rect 310404 240054 311004 275498
rect 310404 239818 310586 240054
rect 310822 239818 311004 240054
rect 310404 239734 311004 239818
rect 310404 239498 310586 239734
rect 310822 239498 311004 239734
rect 310404 204054 311004 239498
rect 310404 203818 310586 204054
rect 310822 203818 311004 204054
rect 310404 203734 311004 203818
rect 310404 203498 310586 203734
rect 310822 203498 311004 203734
rect 310404 168054 311004 203498
rect 310404 167818 310586 168054
rect 310822 167818 311004 168054
rect 310404 167734 311004 167818
rect 310404 167498 310586 167734
rect 310822 167498 311004 167734
rect 310404 132054 311004 167498
rect 310404 131818 310586 132054
rect 310822 131818 311004 132054
rect 310404 131734 311004 131818
rect 310404 131498 310586 131734
rect 310822 131498 311004 131734
rect 310404 96054 311004 131498
rect 310404 95818 310586 96054
rect 310822 95818 311004 96054
rect 310404 95734 311004 95818
rect 310404 95498 310586 95734
rect 310822 95498 311004 95734
rect 310404 60054 311004 95498
rect 310404 59818 310586 60054
rect 310822 59818 311004 60054
rect 310404 59734 311004 59818
rect 310404 59498 310586 59734
rect 310822 59498 311004 59734
rect 310404 24054 311004 59498
rect 310404 23818 310586 24054
rect 310822 23818 311004 24054
rect 310404 23734 311004 23818
rect 310404 23498 310586 23734
rect 310822 23498 311004 23734
rect 310404 -3166 311004 23498
rect 310404 -3402 310586 -3166
rect 310822 -3402 311004 -3166
rect 310404 -3486 311004 -3402
rect 310404 -3722 310586 -3486
rect 310822 -3722 311004 -3486
rect 310404 -3744 311004 -3722
rect 314004 531654 314604 557000
rect 314004 531418 314186 531654
rect 314422 531418 314604 531654
rect 314004 531334 314604 531418
rect 314004 531098 314186 531334
rect 314422 531098 314604 531334
rect 314004 495654 314604 531098
rect 314004 495418 314186 495654
rect 314422 495418 314604 495654
rect 314004 495334 314604 495418
rect 314004 495098 314186 495334
rect 314422 495098 314604 495334
rect 314004 459654 314604 495098
rect 314004 459418 314186 459654
rect 314422 459418 314604 459654
rect 314004 459334 314604 459418
rect 314004 459098 314186 459334
rect 314422 459098 314604 459334
rect 314004 423654 314604 459098
rect 314004 423418 314186 423654
rect 314422 423418 314604 423654
rect 314004 423334 314604 423418
rect 314004 423098 314186 423334
rect 314422 423098 314604 423334
rect 314004 387654 314604 423098
rect 314004 387418 314186 387654
rect 314422 387418 314604 387654
rect 314004 387334 314604 387418
rect 314004 387098 314186 387334
rect 314422 387098 314604 387334
rect 314004 351654 314604 387098
rect 314004 351418 314186 351654
rect 314422 351418 314604 351654
rect 314004 351334 314604 351418
rect 314004 351098 314186 351334
rect 314422 351098 314604 351334
rect 314004 315654 314604 351098
rect 314004 315418 314186 315654
rect 314422 315418 314604 315654
rect 314004 315334 314604 315418
rect 314004 315098 314186 315334
rect 314422 315098 314604 315334
rect 314004 279654 314604 315098
rect 314004 279418 314186 279654
rect 314422 279418 314604 279654
rect 314004 279334 314604 279418
rect 314004 279098 314186 279334
rect 314422 279098 314604 279334
rect 314004 243654 314604 279098
rect 314004 243418 314186 243654
rect 314422 243418 314604 243654
rect 314004 243334 314604 243418
rect 314004 243098 314186 243334
rect 314422 243098 314604 243334
rect 314004 207654 314604 243098
rect 314004 207418 314186 207654
rect 314422 207418 314604 207654
rect 314004 207334 314604 207418
rect 314004 207098 314186 207334
rect 314422 207098 314604 207334
rect 314004 171654 314604 207098
rect 314004 171418 314186 171654
rect 314422 171418 314604 171654
rect 314004 171334 314604 171418
rect 314004 171098 314186 171334
rect 314422 171098 314604 171334
rect 314004 135654 314604 171098
rect 314004 135418 314186 135654
rect 314422 135418 314604 135654
rect 314004 135334 314604 135418
rect 314004 135098 314186 135334
rect 314422 135098 314604 135334
rect 314004 99654 314604 135098
rect 314004 99418 314186 99654
rect 314422 99418 314604 99654
rect 314004 99334 314604 99418
rect 314004 99098 314186 99334
rect 314422 99098 314604 99334
rect 314004 63654 314604 99098
rect 314004 63418 314186 63654
rect 314422 63418 314604 63654
rect 314004 63334 314604 63418
rect 314004 63098 314186 63334
rect 314422 63098 314604 63334
rect 314004 27654 314604 63098
rect 314004 27418 314186 27654
rect 314422 27418 314604 27654
rect 314004 27334 314604 27418
rect 314004 27098 314186 27334
rect 314422 27098 314604 27334
rect 314004 -5046 314604 27098
rect 314004 -5282 314186 -5046
rect 314422 -5282 314604 -5046
rect 314004 -5366 314604 -5282
rect 314004 -5602 314186 -5366
rect 314422 -5602 314604 -5366
rect 314004 -5624 314604 -5602
rect 317604 535254 318204 557000
rect 317604 535018 317786 535254
rect 318022 535018 318204 535254
rect 317604 534934 318204 535018
rect 317604 534698 317786 534934
rect 318022 534698 318204 534934
rect 317604 499254 318204 534698
rect 317604 499018 317786 499254
rect 318022 499018 318204 499254
rect 317604 498934 318204 499018
rect 317604 498698 317786 498934
rect 318022 498698 318204 498934
rect 317604 463254 318204 498698
rect 317604 463018 317786 463254
rect 318022 463018 318204 463254
rect 317604 462934 318204 463018
rect 317604 462698 317786 462934
rect 318022 462698 318204 462934
rect 317604 427254 318204 462698
rect 317604 427018 317786 427254
rect 318022 427018 318204 427254
rect 317604 426934 318204 427018
rect 317604 426698 317786 426934
rect 318022 426698 318204 426934
rect 317604 391254 318204 426698
rect 317604 391018 317786 391254
rect 318022 391018 318204 391254
rect 317604 390934 318204 391018
rect 317604 390698 317786 390934
rect 318022 390698 318204 390934
rect 317604 355254 318204 390698
rect 317604 355018 317786 355254
rect 318022 355018 318204 355254
rect 317604 354934 318204 355018
rect 317604 354698 317786 354934
rect 318022 354698 318204 354934
rect 317604 319254 318204 354698
rect 317604 319018 317786 319254
rect 318022 319018 318204 319254
rect 317604 318934 318204 319018
rect 317604 318698 317786 318934
rect 318022 318698 318204 318934
rect 317604 283254 318204 318698
rect 317604 283018 317786 283254
rect 318022 283018 318204 283254
rect 317604 282934 318204 283018
rect 317604 282698 317786 282934
rect 318022 282698 318204 282934
rect 317604 247254 318204 282698
rect 317604 247018 317786 247254
rect 318022 247018 318204 247254
rect 317604 246934 318204 247018
rect 317604 246698 317786 246934
rect 318022 246698 318204 246934
rect 317604 211254 318204 246698
rect 317604 211018 317786 211254
rect 318022 211018 318204 211254
rect 317604 210934 318204 211018
rect 317604 210698 317786 210934
rect 318022 210698 318204 210934
rect 317604 175254 318204 210698
rect 317604 175018 317786 175254
rect 318022 175018 318204 175254
rect 317604 174934 318204 175018
rect 317604 174698 317786 174934
rect 318022 174698 318204 174934
rect 317604 139254 318204 174698
rect 317604 139018 317786 139254
rect 318022 139018 318204 139254
rect 317604 138934 318204 139018
rect 317604 138698 317786 138934
rect 318022 138698 318204 138934
rect 317604 103254 318204 138698
rect 317604 103018 317786 103254
rect 318022 103018 318204 103254
rect 317604 102934 318204 103018
rect 317604 102698 317786 102934
rect 318022 102698 318204 102934
rect 317604 67254 318204 102698
rect 317604 67018 317786 67254
rect 318022 67018 318204 67254
rect 317604 66934 318204 67018
rect 317604 66698 317786 66934
rect 318022 66698 318204 66934
rect 317604 31254 318204 66698
rect 317604 31018 317786 31254
rect 318022 31018 318204 31254
rect 317604 30934 318204 31018
rect 317604 30698 317786 30934
rect 318022 30698 318204 30934
rect 299604 -6222 299786 -5986
rect 300022 -6222 300204 -5986
rect 299604 -6306 300204 -6222
rect 299604 -6542 299786 -6306
rect 300022 -6542 300204 -6306
rect 299604 -7504 300204 -6542
rect 317604 -6926 318204 30698
rect 324804 542454 325404 557000
rect 324804 542218 324986 542454
rect 325222 542218 325404 542454
rect 324804 542134 325404 542218
rect 324804 541898 324986 542134
rect 325222 541898 325404 542134
rect 324804 506454 325404 541898
rect 324804 506218 324986 506454
rect 325222 506218 325404 506454
rect 324804 506134 325404 506218
rect 324804 505898 324986 506134
rect 325222 505898 325404 506134
rect 324804 470454 325404 505898
rect 324804 470218 324986 470454
rect 325222 470218 325404 470454
rect 324804 470134 325404 470218
rect 324804 469898 324986 470134
rect 325222 469898 325404 470134
rect 324804 434454 325404 469898
rect 324804 434218 324986 434454
rect 325222 434218 325404 434454
rect 324804 434134 325404 434218
rect 324804 433898 324986 434134
rect 325222 433898 325404 434134
rect 324804 398454 325404 433898
rect 324804 398218 324986 398454
rect 325222 398218 325404 398454
rect 324804 398134 325404 398218
rect 324804 397898 324986 398134
rect 325222 397898 325404 398134
rect 324804 362454 325404 397898
rect 324804 362218 324986 362454
rect 325222 362218 325404 362454
rect 324804 362134 325404 362218
rect 324804 361898 324986 362134
rect 325222 361898 325404 362134
rect 324804 326454 325404 361898
rect 324804 326218 324986 326454
rect 325222 326218 325404 326454
rect 324804 326134 325404 326218
rect 324804 325898 324986 326134
rect 325222 325898 325404 326134
rect 324804 290454 325404 325898
rect 324804 290218 324986 290454
rect 325222 290218 325404 290454
rect 324804 290134 325404 290218
rect 324804 289898 324986 290134
rect 325222 289898 325404 290134
rect 324804 254454 325404 289898
rect 324804 254218 324986 254454
rect 325222 254218 325404 254454
rect 324804 254134 325404 254218
rect 324804 253898 324986 254134
rect 325222 253898 325404 254134
rect 324804 218454 325404 253898
rect 324804 218218 324986 218454
rect 325222 218218 325404 218454
rect 324804 218134 325404 218218
rect 324804 217898 324986 218134
rect 325222 217898 325404 218134
rect 324804 182454 325404 217898
rect 324804 182218 324986 182454
rect 325222 182218 325404 182454
rect 324804 182134 325404 182218
rect 324804 181898 324986 182134
rect 325222 181898 325404 182134
rect 324804 146454 325404 181898
rect 324804 146218 324986 146454
rect 325222 146218 325404 146454
rect 324804 146134 325404 146218
rect 324804 145898 324986 146134
rect 325222 145898 325404 146134
rect 324804 110454 325404 145898
rect 324804 110218 324986 110454
rect 325222 110218 325404 110454
rect 324804 110134 325404 110218
rect 324804 109898 324986 110134
rect 325222 109898 325404 110134
rect 324804 74454 325404 109898
rect 324804 74218 324986 74454
rect 325222 74218 325404 74454
rect 324804 74134 325404 74218
rect 324804 73898 324986 74134
rect 325222 73898 325404 74134
rect 324804 38454 325404 73898
rect 324804 38218 324986 38454
rect 325222 38218 325404 38454
rect 324804 38134 325404 38218
rect 324804 37898 324986 38134
rect 325222 37898 325404 38134
rect 324804 2454 325404 37898
rect 324804 2218 324986 2454
rect 325222 2218 325404 2454
rect 324804 2134 325404 2218
rect 324804 1898 324986 2134
rect 325222 1898 325404 2134
rect 324804 -346 325404 1898
rect 324804 -582 324986 -346
rect 325222 -582 325404 -346
rect 324804 -666 325404 -582
rect 324804 -902 324986 -666
rect 325222 -902 325404 -666
rect 324804 -1864 325404 -902
rect 328404 546054 329004 557000
rect 328404 545818 328586 546054
rect 328822 545818 329004 546054
rect 328404 545734 329004 545818
rect 328404 545498 328586 545734
rect 328822 545498 329004 545734
rect 328404 510054 329004 545498
rect 328404 509818 328586 510054
rect 328822 509818 329004 510054
rect 328404 509734 329004 509818
rect 328404 509498 328586 509734
rect 328822 509498 329004 509734
rect 328404 474054 329004 509498
rect 328404 473818 328586 474054
rect 328822 473818 329004 474054
rect 328404 473734 329004 473818
rect 328404 473498 328586 473734
rect 328822 473498 329004 473734
rect 328404 438054 329004 473498
rect 328404 437818 328586 438054
rect 328822 437818 329004 438054
rect 328404 437734 329004 437818
rect 328404 437498 328586 437734
rect 328822 437498 329004 437734
rect 328404 402054 329004 437498
rect 328404 401818 328586 402054
rect 328822 401818 329004 402054
rect 328404 401734 329004 401818
rect 328404 401498 328586 401734
rect 328822 401498 329004 401734
rect 328404 366054 329004 401498
rect 328404 365818 328586 366054
rect 328822 365818 329004 366054
rect 328404 365734 329004 365818
rect 328404 365498 328586 365734
rect 328822 365498 329004 365734
rect 328404 330054 329004 365498
rect 328404 329818 328586 330054
rect 328822 329818 329004 330054
rect 328404 329734 329004 329818
rect 328404 329498 328586 329734
rect 328822 329498 329004 329734
rect 328404 294054 329004 329498
rect 328404 293818 328586 294054
rect 328822 293818 329004 294054
rect 328404 293734 329004 293818
rect 328404 293498 328586 293734
rect 328822 293498 329004 293734
rect 328404 258054 329004 293498
rect 328404 257818 328586 258054
rect 328822 257818 329004 258054
rect 328404 257734 329004 257818
rect 328404 257498 328586 257734
rect 328822 257498 329004 257734
rect 328404 222054 329004 257498
rect 328404 221818 328586 222054
rect 328822 221818 329004 222054
rect 328404 221734 329004 221818
rect 328404 221498 328586 221734
rect 328822 221498 329004 221734
rect 328404 186054 329004 221498
rect 328404 185818 328586 186054
rect 328822 185818 329004 186054
rect 328404 185734 329004 185818
rect 328404 185498 328586 185734
rect 328822 185498 329004 185734
rect 328404 150054 329004 185498
rect 328404 149818 328586 150054
rect 328822 149818 329004 150054
rect 328404 149734 329004 149818
rect 328404 149498 328586 149734
rect 328822 149498 329004 149734
rect 328404 114054 329004 149498
rect 328404 113818 328586 114054
rect 328822 113818 329004 114054
rect 328404 113734 329004 113818
rect 328404 113498 328586 113734
rect 328822 113498 329004 113734
rect 328404 78054 329004 113498
rect 328404 77818 328586 78054
rect 328822 77818 329004 78054
rect 328404 77734 329004 77818
rect 328404 77498 328586 77734
rect 328822 77498 329004 77734
rect 328404 42054 329004 77498
rect 328404 41818 328586 42054
rect 328822 41818 329004 42054
rect 328404 41734 329004 41818
rect 328404 41498 328586 41734
rect 328822 41498 329004 41734
rect 328404 6054 329004 41498
rect 328404 5818 328586 6054
rect 328822 5818 329004 6054
rect 328404 5734 329004 5818
rect 328404 5498 328586 5734
rect 328822 5498 329004 5734
rect 328404 -2226 329004 5498
rect 328404 -2462 328586 -2226
rect 328822 -2462 329004 -2226
rect 328404 -2546 329004 -2462
rect 328404 -2782 328586 -2546
rect 328822 -2782 329004 -2546
rect 328404 -3744 329004 -2782
rect 332004 549654 332604 557000
rect 332004 549418 332186 549654
rect 332422 549418 332604 549654
rect 332004 549334 332604 549418
rect 332004 549098 332186 549334
rect 332422 549098 332604 549334
rect 332004 513654 332604 549098
rect 332004 513418 332186 513654
rect 332422 513418 332604 513654
rect 332004 513334 332604 513418
rect 332004 513098 332186 513334
rect 332422 513098 332604 513334
rect 332004 477654 332604 513098
rect 332004 477418 332186 477654
rect 332422 477418 332604 477654
rect 332004 477334 332604 477418
rect 332004 477098 332186 477334
rect 332422 477098 332604 477334
rect 332004 441654 332604 477098
rect 332004 441418 332186 441654
rect 332422 441418 332604 441654
rect 332004 441334 332604 441418
rect 332004 441098 332186 441334
rect 332422 441098 332604 441334
rect 332004 405654 332604 441098
rect 332004 405418 332186 405654
rect 332422 405418 332604 405654
rect 332004 405334 332604 405418
rect 332004 405098 332186 405334
rect 332422 405098 332604 405334
rect 332004 369654 332604 405098
rect 332004 369418 332186 369654
rect 332422 369418 332604 369654
rect 332004 369334 332604 369418
rect 332004 369098 332186 369334
rect 332422 369098 332604 369334
rect 332004 333654 332604 369098
rect 332004 333418 332186 333654
rect 332422 333418 332604 333654
rect 332004 333334 332604 333418
rect 332004 333098 332186 333334
rect 332422 333098 332604 333334
rect 332004 297654 332604 333098
rect 332004 297418 332186 297654
rect 332422 297418 332604 297654
rect 332004 297334 332604 297418
rect 332004 297098 332186 297334
rect 332422 297098 332604 297334
rect 332004 261654 332604 297098
rect 332004 261418 332186 261654
rect 332422 261418 332604 261654
rect 332004 261334 332604 261418
rect 332004 261098 332186 261334
rect 332422 261098 332604 261334
rect 332004 225654 332604 261098
rect 332004 225418 332186 225654
rect 332422 225418 332604 225654
rect 332004 225334 332604 225418
rect 332004 225098 332186 225334
rect 332422 225098 332604 225334
rect 332004 189654 332604 225098
rect 332004 189418 332186 189654
rect 332422 189418 332604 189654
rect 332004 189334 332604 189418
rect 332004 189098 332186 189334
rect 332422 189098 332604 189334
rect 332004 153654 332604 189098
rect 332004 153418 332186 153654
rect 332422 153418 332604 153654
rect 332004 153334 332604 153418
rect 332004 153098 332186 153334
rect 332422 153098 332604 153334
rect 332004 117654 332604 153098
rect 332004 117418 332186 117654
rect 332422 117418 332604 117654
rect 332004 117334 332604 117418
rect 332004 117098 332186 117334
rect 332422 117098 332604 117334
rect 332004 81654 332604 117098
rect 332004 81418 332186 81654
rect 332422 81418 332604 81654
rect 332004 81334 332604 81418
rect 332004 81098 332186 81334
rect 332422 81098 332604 81334
rect 332004 45654 332604 81098
rect 332004 45418 332186 45654
rect 332422 45418 332604 45654
rect 332004 45334 332604 45418
rect 332004 45098 332186 45334
rect 332422 45098 332604 45334
rect 332004 9654 332604 45098
rect 332004 9418 332186 9654
rect 332422 9418 332604 9654
rect 332004 9334 332604 9418
rect 332004 9098 332186 9334
rect 332422 9098 332604 9334
rect 332004 -4106 332604 9098
rect 332004 -4342 332186 -4106
rect 332422 -4342 332604 -4106
rect 332004 -4426 332604 -4342
rect 332004 -4662 332186 -4426
rect 332422 -4662 332604 -4426
rect 332004 -5624 332604 -4662
rect 335604 553254 336204 557000
rect 335604 553018 335786 553254
rect 336022 553018 336204 553254
rect 335604 552934 336204 553018
rect 335604 552698 335786 552934
rect 336022 552698 336204 552934
rect 335604 517254 336204 552698
rect 335604 517018 335786 517254
rect 336022 517018 336204 517254
rect 335604 516934 336204 517018
rect 335604 516698 335786 516934
rect 336022 516698 336204 516934
rect 335604 481254 336204 516698
rect 335604 481018 335786 481254
rect 336022 481018 336204 481254
rect 335604 480934 336204 481018
rect 335604 480698 335786 480934
rect 336022 480698 336204 480934
rect 335604 445254 336204 480698
rect 335604 445018 335786 445254
rect 336022 445018 336204 445254
rect 335604 444934 336204 445018
rect 335604 444698 335786 444934
rect 336022 444698 336204 444934
rect 335604 409254 336204 444698
rect 342804 524454 343404 557000
rect 342804 524218 342986 524454
rect 343222 524218 343404 524454
rect 342804 524134 343404 524218
rect 342804 523898 342986 524134
rect 343222 523898 343404 524134
rect 342804 488454 343404 523898
rect 342804 488218 342986 488454
rect 343222 488218 343404 488454
rect 342804 488134 343404 488218
rect 342804 487898 342986 488134
rect 343222 487898 343404 488134
rect 342804 452454 343404 487898
rect 342804 452218 342986 452454
rect 343222 452218 343404 452454
rect 342804 452134 343404 452218
rect 342804 451898 342986 452134
rect 343222 451898 343404 452134
rect 342804 416454 343404 451898
rect 342804 416218 342986 416454
rect 343222 416218 343404 416454
rect 342804 416134 343404 416218
rect 342804 415898 342986 416134
rect 343222 415898 343404 416134
rect 342804 414247 343404 415898
rect 346404 528054 347004 557000
rect 347819 545460 347885 545461
rect 347819 545396 347820 545460
rect 347884 545396 347885 545460
rect 347819 545395 347885 545396
rect 347822 545189 347882 545395
rect 347819 545188 347885 545189
rect 347819 545124 347820 545188
rect 347884 545124 347885 545188
rect 347819 545123 347885 545124
rect 346404 527818 346586 528054
rect 346822 527818 347004 528054
rect 346404 527734 347004 527818
rect 346404 527498 346586 527734
rect 346822 527498 347004 527734
rect 346404 492054 347004 527498
rect 346404 491818 346586 492054
rect 346822 491818 347004 492054
rect 346404 491734 347004 491818
rect 346404 491498 346586 491734
rect 346822 491498 347004 491734
rect 346404 456054 347004 491498
rect 346404 455818 346586 456054
rect 346822 455818 347004 456054
rect 346404 455734 347004 455818
rect 346404 455498 346586 455734
rect 346822 455498 347004 455734
rect 346404 420054 347004 455498
rect 346404 419818 346586 420054
rect 346822 419818 347004 420054
rect 346404 419734 347004 419818
rect 346404 419498 346586 419734
rect 346822 419498 347004 419734
rect 346404 414247 347004 419498
rect 350004 531654 350604 557000
rect 350004 531418 350186 531654
rect 350422 531418 350604 531654
rect 350004 531334 350604 531418
rect 350004 531098 350186 531334
rect 350422 531098 350604 531334
rect 350004 495654 350604 531098
rect 350004 495418 350186 495654
rect 350422 495418 350604 495654
rect 350004 495334 350604 495418
rect 350004 495098 350186 495334
rect 350422 495098 350604 495334
rect 350004 459654 350604 495098
rect 350004 459418 350186 459654
rect 350422 459418 350604 459654
rect 350004 459334 350604 459418
rect 350004 459098 350186 459334
rect 350422 459098 350604 459334
rect 350004 423654 350604 459098
rect 350004 423418 350186 423654
rect 350422 423418 350604 423654
rect 350004 423334 350604 423418
rect 350004 423098 350186 423334
rect 350422 423098 350604 423334
rect 350004 414247 350604 423098
rect 353604 535254 354204 557000
rect 357387 545188 357453 545189
rect 357387 545124 357388 545188
rect 357452 545124 357453 545188
rect 357387 545123 357453 545124
rect 357390 544917 357450 545123
rect 357387 544916 357453 544917
rect 357387 544852 357388 544916
rect 357452 544852 357453 544916
rect 357387 544851 357453 544852
rect 353604 535018 353786 535254
rect 354022 535018 354204 535254
rect 353604 534934 354204 535018
rect 353604 534698 353786 534934
rect 354022 534698 354204 534934
rect 353604 499254 354204 534698
rect 353604 499018 353786 499254
rect 354022 499018 354204 499254
rect 353604 498934 354204 499018
rect 353604 498698 353786 498934
rect 354022 498698 354204 498934
rect 353604 463254 354204 498698
rect 353604 463018 353786 463254
rect 354022 463018 354204 463254
rect 353604 462934 354204 463018
rect 353604 462698 353786 462934
rect 354022 462698 354204 462934
rect 353604 427254 354204 462698
rect 353604 427018 353786 427254
rect 354022 427018 354204 427254
rect 353604 426934 354204 427018
rect 353604 426698 353786 426934
rect 354022 426698 354204 426934
rect 353604 414247 354204 426698
rect 360804 542454 361404 557000
rect 360804 542218 360986 542454
rect 361222 542218 361404 542454
rect 360804 542134 361404 542218
rect 360804 541898 360986 542134
rect 361222 541898 361404 542134
rect 360804 506454 361404 541898
rect 360804 506218 360986 506454
rect 361222 506218 361404 506454
rect 360804 506134 361404 506218
rect 360804 505898 360986 506134
rect 361222 505898 361404 506134
rect 360804 470454 361404 505898
rect 360804 470218 360986 470454
rect 361222 470218 361404 470454
rect 360804 470134 361404 470218
rect 360804 469898 360986 470134
rect 361222 469898 361404 470134
rect 360804 434454 361404 469898
rect 360804 434218 360986 434454
rect 361222 434218 361404 434454
rect 360804 434134 361404 434218
rect 360804 433898 360986 434134
rect 361222 433898 361404 434134
rect 360804 414247 361404 433898
rect 364404 546054 365004 557000
rect 364404 545818 364586 546054
rect 364822 545818 365004 546054
rect 364404 545734 365004 545818
rect 364404 545498 364586 545734
rect 364822 545498 365004 545734
rect 364404 510054 365004 545498
rect 364404 509818 364586 510054
rect 364822 509818 365004 510054
rect 364404 509734 365004 509818
rect 364404 509498 364586 509734
rect 364822 509498 365004 509734
rect 364404 474054 365004 509498
rect 364404 473818 364586 474054
rect 364822 473818 365004 474054
rect 364404 473734 365004 473818
rect 364404 473498 364586 473734
rect 364822 473498 365004 473734
rect 364404 438054 365004 473498
rect 364404 437818 364586 438054
rect 364822 437818 365004 438054
rect 364404 437734 365004 437818
rect 364404 437498 364586 437734
rect 364822 437498 365004 437734
rect 364404 414247 365004 437498
rect 368004 549654 368604 557000
rect 368004 549418 368186 549654
rect 368422 549418 368604 549654
rect 368004 549334 368604 549418
rect 368004 549098 368186 549334
rect 368422 549098 368604 549334
rect 368004 513654 368604 549098
rect 368004 513418 368186 513654
rect 368422 513418 368604 513654
rect 368004 513334 368604 513418
rect 368004 513098 368186 513334
rect 368422 513098 368604 513334
rect 368004 477654 368604 513098
rect 368004 477418 368186 477654
rect 368422 477418 368604 477654
rect 368004 477334 368604 477418
rect 368004 477098 368186 477334
rect 368422 477098 368604 477334
rect 368004 441654 368604 477098
rect 368004 441418 368186 441654
rect 368422 441418 368604 441654
rect 368004 441334 368604 441418
rect 368004 441098 368186 441334
rect 368422 441098 368604 441334
rect 368004 414247 368604 441098
rect 371604 553254 372204 557000
rect 371604 553018 371786 553254
rect 372022 553018 372204 553254
rect 371604 552934 372204 553018
rect 371604 552698 371786 552934
rect 372022 552698 372204 552934
rect 371604 517254 372204 552698
rect 376707 545460 376773 545461
rect 376707 545396 376708 545460
rect 376772 545396 376773 545460
rect 376707 545395 376773 545396
rect 376710 545189 376770 545395
rect 376707 545188 376773 545189
rect 376707 545124 376708 545188
rect 376772 545124 376773 545188
rect 376707 545123 376773 545124
rect 371604 517018 371786 517254
rect 372022 517018 372204 517254
rect 371604 516934 372204 517018
rect 371604 516698 371786 516934
rect 372022 516698 372204 516934
rect 371604 481254 372204 516698
rect 371604 481018 371786 481254
rect 372022 481018 372204 481254
rect 371604 480934 372204 481018
rect 371604 480698 371786 480934
rect 372022 480698 372204 480934
rect 371604 445254 372204 480698
rect 371604 445018 371786 445254
rect 372022 445018 372204 445254
rect 371604 444934 372204 445018
rect 371604 444698 371786 444934
rect 372022 444698 372204 444934
rect 371604 414247 372204 444698
rect 378804 524454 379404 557000
rect 378804 524218 378986 524454
rect 379222 524218 379404 524454
rect 378804 524134 379404 524218
rect 378804 523898 378986 524134
rect 379222 523898 379404 524134
rect 378804 488454 379404 523898
rect 378804 488218 378986 488454
rect 379222 488218 379404 488454
rect 378804 488134 379404 488218
rect 378804 487898 378986 488134
rect 379222 487898 379404 488134
rect 378804 452454 379404 487898
rect 378804 452218 378986 452454
rect 379222 452218 379404 452454
rect 378804 452134 379404 452218
rect 378804 451898 378986 452134
rect 379222 451898 379404 452134
rect 378804 416454 379404 451898
rect 378804 416218 378986 416454
rect 379222 416218 379404 416454
rect 378804 416134 379404 416218
rect 378804 415898 378986 416134
rect 379222 415898 379404 416134
rect 378804 414247 379404 415898
rect 382404 528054 383004 557000
rect 382404 527818 382586 528054
rect 382822 527818 383004 528054
rect 382404 527734 383004 527818
rect 382404 527498 382586 527734
rect 382822 527498 383004 527734
rect 382404 492054 383004 527498
rect 382404 491818 382586 492054
rect 382822 491818 383004 492054
rect 382404 491734 383004 491818
rect 382404 491498 382586 491734
rect 382822 491498 383004 491734
rect 382404 456054 383004 491498
rect 382404 455818 382586 456054
rect 382822 455818 383004 456054
rect 382404 455734 383004 455818
rect 382404 455498 382586 455734
rect 382822 455498 383004 455734
rect 382404 420054 383004 455498
rect 382404 419818 382586 420054
rect 382822 419818 383004 420054
rect 382404 419734 383004 419818
rect 382404 419498 382586 419734
rect 382822 419498 383004 419734
rect 382404 414247 383004 419498
rect 386004 531654 386604 557000
rect 386004 531418 386186 531654
rect 386422 531418 386604 531654
rect 386004 531334 386604 531418
rect 386004 531098 386186 531334
rect 386422 531098 386604 531334
rect 386004 495654 386604 531098
rect 386004 495418 386186 495654
rect 386422 495418 386604 495654
rect 386004 495334 386604 495418
rect 386004 495098 386186 495334
rect 386422 495098 386604 495334
rect 386004 459654 386604 495098
rect 386004 459418 386186 459654
rect 386422 459418 386604 459654
rect 386004 459334 386604 459418
rect 386004 459098 386186 459334
rect 386422 459098 386604 459334
rect 386004 423654 386604 459098
rect 386004 423418 386186 423654
rect 386422 423418 386604 423654
rect 386004 423334 386604 423418
rect 386004 423098 386186 423334
rect 386422 423098 386604 423334
rect 386004 414247 386604 423098
rect 389604 535254 390204 557000
rect 389604 535018 389786 535254
rect 390022 535018 390204 535254
rect 389604 534934 390204 535018
rect 389604 534698 389786 534934
rect 390022 534698 390204 534934
rect 389604 499254 390204 534698
rect 389604 499018 389786 499254
rect 390022 499018 390204 499254
rect 389604 498934 390204 499018
rect 389604 498698 389786 498934
rect 390022 498698 390204 498934
rect 389604 463254 390204 498698
rect 389604 463018 389786 463254
rect 390022 463018 390204 463254
rect 389604 462934 390204 463018
rect 389604 462698 389786 462934
rect 390022 462698 390204 462934
rect 389604 427254 390204 462698
rect 389604 427018 389786 427254
rect 390022 427018 390204 427254
rect 389604 426934 390204 427018
rect 389604 426698 389786 426934
rect 390022 426698 390204 426934
rect 389604 414247 390204 426698
rect 396804 542454 397404 577898
rect 396804 542218 396986 542454
rect 397222 542218 397404 542454
rect 396804 542134 397404 542218
rect 396804 541898 396986 542134
rect 397222 541898 397404 542134
rect 396804 506454 397404 541898
rect 396804 506218 396986 506454
rect 397222 506218 397404 506454
rect 396804 506134 397404 506218
rect 396804 505898 396986 506134
rect 397222 505898 397404 506134
rect 396804 470454 397404 505898
rect 396804 470218 396986 470454
rect 397222 470218 397404 470454
rect 396804 470134 397404 470218
rect 396804 469898 396986 470134
rect 397222 469898 397404 470134
rect 396804 434454 397404 469898
rect 396804 434218 396986 434454
rect 397222 434218 397404 434454
rect 396804 434134 397404 434218
rect 396804 433898 396986 434134
rect 397222 433898 397404 434134
rect 396804 414247 397404 433898
rect 400404 690054 401004 706162
rect 400404 689818 400586 690054
rect 400822 689818 401004 690054
rect 400404 689734 401004 689818
rect 400404 689498 400586 689734
rect 400822 689498 401004 689734
rect 400404 654054 401004 689498
rect 400404 653818 400586 654054
rect 400822 653818 401004 654054
rect 400404 653734 401004 653818
rect 400404 653498 400586 653734
rect 400822 653498 401004 653734
rect 400404 618054 401004 653498
rect 400404 617818 400586 618054
rect 400822 617818 401004 618054
rect 400404 617734 401004 617818
rect 400404 617498 400586 617734
rect 400822 617498 401004 617734
rect 400404 582054 401004 617498
rect 400404 581818 400586 582054
rect 400822 581818 401004 582054
rect 400404 581734 401004 581818
rect 400404 581498 400586 581734
rect 400822 581498 401004 581734
rect 400404 546054 401004 581498
rect 400404 545818 400586 546054
rect 400822 545818 401004 546054
rect 400404 545734 401004 545818
rect 400404 545498 400586 545734
rect 400822 545498 401004 545734
rect 400404 510054 401004 545498
rect 400404 509818 400586 510054
rect 400822 509818 401004 510054
rect 400404 509734 401004 509818
rect 400404 509498 400586 509734
rect 400822 509498 401004 509734
rect 400404 474054 401004 509498
rect 400404 473818 400586 474054
rect 400822 473818 401004 474054
rect 400404 473734 401004 473818
rect 400404 473498 400586 473734
rect 400822 473498 401004 473734
rect 400404 438054 401004 473498
rect 400404 437818 400586 438054
rect 400822 437818 401004 438054
rect 400404 437734 401004 437818
rect 400404 437498 400586 437734
rect 400822 437498 401004 437734
rect 400404 414247 401004 437498
rect 404004 693654 404604 708042
rect 404004 693418 404186 693654
rect 404422 693418 404604 693654
rect 404004 693334 404604 693418
rect 404004 693098 404186 693334
rect 404422 693098 404604 693334
rect 404004 657654 404604 693098
rect 404004 657418 404186 657654
rect 404422 657418 404604 657654
rect 404004 657334 404604 657418
rect 404004 657098 404186 657334
rect 404422 657098 404604 657334
rect 404004 621654 404604 657098
rect 404004 621418 404186 621654
rect 404422 621418 404604 621654
rect 404004 621334 404604 621418
rect 404004 621098 404186 621334
rect 404422 621098 404604 621334
rect 404004 585654 404604 621098
rect 404004 585418 404186 585654
rect 404422 585418 404604 585654
rect 404004 585334 404604 585418
rect 404004 585098 404186 585334
rect 404422 585098 404604 585334
rect 404004 549654 404604 585098
rect 404004 549418 404186 549654
rect 404422 549418 404604 549654
rect 404004 549334 404604 549418
rect 404004 549098 404186 549334
rect 404422 549098 404604 549334
rect 404004 513654 404604 549098
rect 404004 513418 404186 513654
rect 404422 513418 404604 513654
rect 404004 513334 404604 513418
rect 404004 513098 404186 513334
rect 404422 513098 404604 513334
rect 404004 477654 404604 513098
rect 404004 477418 404186 477654
rect 404422 477418 404604 477654
rect 404004 477334 404604 477418
rect 404004 477098 404186 477334
rect 404422 477098 404604 477334
rect 404004 441654 404604 477098
rect 404004 441418 404186 441654
rect 404422 441418 404604 441654
rect 404004 441334 404604 441418
rect 404004 441098 404186 441334
rect 404422 441098 404604 441334
rect 404004 414247 404604 441098
rect 407604 697254 408204 709922
rect 425604 711418 426204 711440
rect 425604 711182 425786 711418
rect 426022 711182 426204 711418
rect 425604 711098 426204 711182
rect 425604 710862 425786 711098
rect 426022 710862 426204 711098
rect 422004 709538 422604 709560
rect 422004 709302 422186 709538
rect 422422 709302 422604 709538
rect 422004 709218 422604 709302
rect 422004 708982 422186 709218
rect 422422 708982 422604 709218
rect 418404 707658 419004 707680
rect 418404 707422 418586 707658
rect 418822 707422 419004 707658
rect 418404 707338 419004 707422
rect 418404 707102 418586 707338
rect 418822 707102 419004 707338
rect 407604 697018 407786 697254
rect 408022 697018 408204 697254
rect 407604 696934 408204 697018
rect 407604 696698 407786 696934
rect 408022 696698 408204 696934
rect 407604 661254 408204 696698
rect 407604 661018 407786 661254
rect 408022 661018 408204 661254
rect 407604 660934 408204 661018
rect 407604 660698 407786 660934
rect 408022 660698 408204 660934
rect 407604 625254 408204 660698
rect 407604 625018 407786 625254
rect 408022 625018 408204 625254
rect 407604 624934 408204 625018
rect 407604 624698 407786 624934
rect 408022 624698 408204 624934
rect 407604 589254 408204 624698
rect 407604 589018 407786 589254
rect 408022 589018 408204 589254
rect 407604 588934 408204 589018
rect 407604 588698 407786 588934
rect 408022 588698 408204 588934
rect 407604 553254 408204 588698
rect 407604 553018 407786 553254
rect 408022 553018 408204 553254
rect 407604 552934 408204 553018
rect 407604 552698 407786 552934
rect 408022 552698 408204 552934
rect 407604 517254 408204 552698
rect 407604 517018 407786 517254
rect 408022 517018 408204 517254
rect 407604 516934 408204 517018
rect 407604 516698 407786 516934
rect 408022 516698 408204 516934
rect 407604 481254 408204 516698
rect 407604 481018 407786 481254
rect 408022 481018 408204 481254
rect 407604 480934 408204 481018
rect 407604 480698 407786 480934
rect 408022 480698 408204 480934
rect 407604 445254 408204 480698
rect 407604 445018 407786 445254
rect 408022 445018 408204 445254
rect 407604 444934 408204 445018
rect 407604 444698 407786 444934
rect 408022 444698 408204 444934
rect 407604 414247 408204 444698
rect 414804 705778 415404 705800
rect 414804 705542 414986 705778
rect 415222 705542 415404 705778
rect 414804 705458 415404 705542
rect 414804 705222 414986 705458
rect 415222 705222 415404 705458
rect 414804 668454 415404 705222
rect 414804 668218 414986 668454
rect 415222 668218 415404 668454
rect 414804 668134 415404 668218
rect 414804 667898 414986 668134
rect 415222 667898 415404 668134
rect 414804 632454 415404 667898
rect 414804 632218 414986 632454
rect 415222 632218 415404 632454
rect 414804 632134 415404 632218
rect 414804 631898 414986 632134
rect 415222 631898 415404 632134
rect 414804 596454 415404 631898
rect 414804 596218 414986 596454
rect 415222 596218 415404 596454
rect 414804 596134 415404 596218
rect 414804 595898 414986 596134
rect 415222 595898 415404 596134
rect 414804 560454 415404 595898
rect 414804 560218 414986 560454
rect 415222 560218 415404 560454
rect 414804 560134 415404 560218
rect 414804 559898 414986 560134
rect 415222 559898 415404 560134
rect 414804 524454 415404 559898
rect 414804 524218 414986 524454
rect 415222 524218 415404 524454
rect 414804 524134 415404 524218
rect 414804 523898 414986 524134
rect 415222 523898 415404 524134
rect 414804 488454 415404 523898
rect 414804 488218 414986 488454
rect 415222 488218 415404 488454
rect 414804 488134 415404 488218
rect 414804 487898 414986 488134
rect 415222 487898 415404 488134
rect 414804 452454 415404 487898
rect 414804 452218 414986 452454
rect 415222 452218 415404 452454
rect 414804 452134 415404 452218
rect 414804 451898 414986 452134
rect 415222 451898 415404 452134
rect 414804 416454 415404 451898
rect 414804 416218 414986 416454
rect 415222 416218 415404 416454
rect 414804 416134 415404 416218
rect 414804 415898 414986 416134
rect 415222 415898 415404 416134
rect 414804 414247 415404 415898
rect 418404 672054 419004 707102
rect 418404 671818 418586 672054
rect 418822 671818 419004 672054
rect 418404 671734 419004 671818
rect 418404 671498 418586 671734
rect 418822 671498 419004 671734
rect 418404 636054 419004 671498
rect 418404 635818 418586 636054
rect 418822 635818 419004 636054
rect 418404 635734 419004 635818
rect 418404 635498 418586 635734
rect 418822 635498 419004 635734
rect 418404 600054 419004 635498
rect 418404 599818 418586 600054
rect 418822 599818 419004 600054
rect 418404 599734 419004 599818
rect 418404 599498 418586 599734
rect 418822 599498 419004 599734
rect 418404 564054 419004 599498
rect 418404 563818 418586 564054
rect 418822 563818 419004 564054
rect 418404 563734 419004 563818
rect 418404 563498 418586 563734
rect 418822 563498 419004 563734
rect 418404 528054 419004 563498
rect 418404 527818 418586 528054
rect 418822 527818 419004 528054
rect 418404 527734 419004 527818
rect 418404 527498 418586 527734
rect 418822 527498 419004 527734
rect 418404 492054 419004 527498
rect 418404 491818 418586 492054
rect 418822 491818 419004 492054
rect 418404 491734 419004 491818
rect 418404 491498 418586 491734
rect 418822 491498 419004 491734
rect 418404 456054 419004 491498
rect 418404 455818 418586 456054
rect 418822 455818 419004 456054
rect 418404 455734 419004 455818
rect 418404 455498 418586 455734
rect 418822 455498 419004 455734
rect 418404 420054 419004 455498
rect 418404 419818 418586 420054
rect 418822 419818 419004 420054
rect 418404 419734 419004 419818
rect 418404 419498 418586 419734
rect 418822 419498 419004 419734
rect 418404 414247 419004 419498
rect 422004 675654 422604 708982
rect 422004 675418 422186 675654
rect 422422 675418 422604 675654
rect 422004 675334 422604 675418
rect 422004 675098 422186 675334
rect 422422 675098 422604 675334
rect 422004 639654 422604 675098
rect 422004 639418 422186 639654
rect 422422 639418 422604 639654
rect 422004 639334 422604 639418
rect 422004 639098 422186 639334
rect 422422 639098 422604 639334
rect 422004 603654 422604 639098
rect 422004 603418 422186 603654
rect 422422 603418 422604 603654
rect 422004 603334 422604 603418
rect 422004 603098 422186 603334
rect 422422 603098 422604 603334
rect 422004 567654 422604 603098
rect 422004 567418 422186 567654
rect 422422 567418 422604 567654
rect 422004 567334 422604 567418
rect 422004 567098 422186 567334
rect 422422 567098 422604 567334
rect 422004 531654 422604 567098
rect 422004 531418 422186 531654
rect 422422 531418 422604 531654
rect 422004 531334 422604 531418
rect 422004 531098 422186 531334
rect 422422 531098 422604 531334
rect 422004 495654 422604 531098
rect 422004 495418 422186 495654
rect 422422 495418 422604 495654
rect 422004 495334 422604 495418
rect 422004 495098 422186 495334
rect 422422 495098 422604 495334
rect 422004 459654 422604 495098
rect 422004 459418 422186 459654
rect 422422 459418 422604 459654
rect 422004 459334 422604 459418
rect 422004 459098 422186 459334
rect 422422 459098 422604 459334
rect 422004 423654 422604 459098
rect 422004 423418 422186 423654
rect 422422 423418 422604 423654
rect 422004 423334 422604 423418
rect 422004 423098 422186 423334
rect 422422 423098 422604 423334
rect 367691 413948 367757 413949
rect 367691 413884 367692 413948
rect 367756 413884 367757 413948
rect 367691 413883 367757 413884
rect 368979 413948 369045 413949
rect 368979 413884 368980 413948
rect 369044 413884 369045 413948
rect 368979 413883 369045 413884
rect 370267 413948 370333 413949
rect 370267 413884 370268 413948
rect 370332 413884 370333 413948
rect 370267 413883 370333 413884
rect 371555 413948 371621 413949
rect 371555 413884 371556 413948
rect 371620 413884 371621 413948
rect 371555 413883 371621 413884
rect 372659 413948 372725 413949
rect 372659 413884 372660 413948
rect 372724 413884 372725 413948
rect 372659 413883 372725 413884
rect 373947 413948 374013 413949
rect 373947 413884 373948 413948
rect 374012 413884 374013 413948
rect 373947 413883 374013 413884
rect 375971 413948 376037 413949
rect 375971 413884 375972 413948
rect 376036 413884 376037 413948
rect 375971 413883 376037 413884
rect 377259 413948 377325 413949
rect 377259 413884 377260 413948
rect 377324 413884 377325 413948
rect 377259 413883 377325 413884
rect 378363 413948 378429 413949
rect 378363 413884 378364 413948
rect 378428 413884 378429 413948
rect 378363 413883 378429 413884
rect 379651 413948 379717 413949
rect 379651 413884 379652 413948
rect 379716 413884 379717 413948
rect 379651 413883 379717 413884
rect 380939 413948 381005 413949
rect 380939 413884 380940 413948
rect 381004 413884 381005 413948
rect 380939 413883 381005 413884
rect 382227 413948 382293 413949
rect 382227 413884 382228 413948
rect 382292 413884 382293 413948
rect 382227 413883 382293 413884
rect 385171 413948 385237 413949
rect 385171 413884 385172 413948
rect 385236 413884 385237 413948
rect 385171 413883 385237 413884
rect 367694 411090 367754 413883
rect 368243 413404 368309 413405
rect 368243 413340 368244 413404
rect 368308 413340 368309 413404
rect 368243 413339 368309 413340
rect 368246 411770 368306 413339
rect 368246 411710 368446 411770
rect 367694 411030 368292 411090
rect 368386 411060 368446 411710
rect 368982 411090 369042 413883
rect 369715 413404 369781 413405
rect 369715 413340 369716 413404
rect 369780 413340 369781 413404
rect 369715 413339 369781 413340
rect 369718 411090 369778 413339
rect 368982 411030 369460 411090
rect 369584 411030 369778 411090
rect 370270 411090 370330 413883
rect 371003 413268 371069 413269
rect 371003 413204 371004 413268
rect 371068 413204 371069 413268
rect 371003 413203 371069 413204
rect 371006 411090 371066 413203
rect 370270 411030 370628 411090
rect 370752 411030 371066 411090
rect 371558 411090 371618 413883
rect 371923 413132 371989 413133
rect 371923 413068 371924 413132
rect 371988 413068 371989 413132
rect 371923 413067 371989 413068
rect 371926 411090 371986 413067
rect 371558 411030 371796 411090
rect 371920 411030 371986 411090
rect 372662 410750 372722 413883
rect 373027 413132 373093 413133
rect 373027 413068 373028 413132
rect 373092 413068 373093 413132
rect 373027 413067 373093 413068
rect 373030 411770 373090 413067
rect 373030 411710 373118 411770
rect 373058 411060 373118 411710
rect 373950 411090 374010 413883
rect 374683 413812 374749 413813
rect 374683 413748 374684 413812
rect 374748 413748 374749 413812
rect 374683 413747 374749 413748
rect 374315 412996 374381 412997
rect 374315 412932 374316 412996
rect 374380 412932 374381 412996
rect 374315 412931 374381 412932
rect 374318 411770 374378 412931
rect 374226 411710 374378 411770
rect 373950 411030 374132 411090
rect 374226 411060 374286 411710
rect 374686 411090 374746 413747
rect 375419 412860 375485 412861
rect 375419 412796 375420 412860
rect 375484 412796 375485 412860
rect 375419 412795 375485 412796
rect 374686 411030 375300 411090
rect 375422 411030 375482 412795
rect 375974 411090 376034 413883
rect 376523 412860 376589 412861
rect 376523 412796 376524 412860
rect 376588 412796 376589 412860
rect 376523 412795 376589 412796
rect 376526 411770 376586 412795
rect 376526 411710 376622 411770
rect 375974 411030 376468 411090
rect 376562 411060 376622 411710
rect 377262 411090 377322 413883
rect 377995 413404 378061 413405
rect 377995 413340 377996 413404
rect 378060 413340 378061 413404
rect 377995 413339 378061 413340
rect 377998 411090 378058 413339
rect 377262 411030 377636 411090
rect 377760 411030 378058 411090
rect 378366 411090 378426 413883
rect 378915 413132 378981 413133
rect 378915 413068 378916 413132
rect 378980 413068 378981 413132
rect 378915 413067 378981 413068
rect 378366 411030 378804 411090
rect 378918 411030 378978 413067
rect 379654 411090 379714 413883
rect 380203 413268 380269 413269
rect 380203 413204 380204 413268
rect 380268 413204 380269 413268
rect 380203 413203 380269 413204
rect 380206 411090 380266 413203
rect 379654 411030 379972 411090
rect 380096 411030 380266 411090
rect 380942 411090 381002 413883
rect 381491 413132 381557 413133
rect 381491 413068 381492 413132
rect 381556 413068 381557 413132
rect 381491 413067 381557 413068
rect 381494 411090 381554 413067
rect 380942 411030 381140 411090
rect 381264 411030 381554 411090
rect 382230 411090 382290 413883
rect 382963 413812 383029 413813
rect 382963 413748 382964 413812
rect 383028 413748 383029 413812
rect 382963 413747 383029 413748
rect 384067 413812 384133 413813
rect 384067 413748 384068 413812
rect 384132 413748 384133 413812
rect 384067 413747 384133 413748
rect 382411 413132 382477 413133
rect 382411 413068 382412 413132
rect 382476 413068 382477 413132
rect 382411 413067 382477 413068
rect 382230 411030 382308 411090
rect 382414 411030 382474 413067
rect 382966 411090 383026 413747
rect 383515 412996 383581 412997
rect 383515 412932 383516 412996
rect 383580 412932 383581 412996
rect 383515 412931 383581 412932
rect 383518 411770 383578 412931
rect 383518 411710 383630 411770
rect 382966 411030 383476 411090
rect 383570 411060 383630 411710
rect 384070 411090 384130 413747
rect 384803 412996 384869 412997
rect 384803 412932 384804 412996
rect 384868 412932 384869 412996
rect 384803 412931 384869 412932
rect 384806 411770 384866 412931
rect 384738 411710 384866 411770
rect 384070 411030 384644 411090
rect 384738 411060 384798 411710
rect 385174 411090 385234 413883
rect 412771 413812 412837 413813
rect 412771 413748 412772 413812
rect 412836 413748 412837 413812
rect 412771 413747 412837 413748
rect 396395 413676 396461 413677
rect 396395 413612 396396 413676
rect 396460 413612 396461 413676
rect 396395 413611 396461 413612
rect 397499 413676 397565 413677
rect 397499 413612 397500 413676
rect 397564 413612 397565 413676
rect 397499 413611 397565 413612
rect 388299 413404 388365 413405
rect 388299 413340 388300 413404
rect 388364 413340 388365 413404
rect 388299 413339 388365 413340
rect 386827 413268 386893 413269
rect 386827 413204 386828 413268
rect 386892 413204 386893 413268
rect 386827 413203 386893 413204
rect 385907 412996 385973 412997
rect 385907 412932 385908 412996
rect 385972 412932 385973 412996
rect 385907 412931 385973 412932
rect 385174 411030 385812 411090
rect 385910 411030 385970 412931
rect 386830 411090 386890 413203
rect 387195 413132 387261 413133
rect 387195 413068 387196 413132
rect 387260 413068 387261 413132
rect 387195 413067 387261 413068
rect 387198 411090 387258 413067
rect 388115 411772 388181 411773
rect 388115 411708 388116 411772
rect 388180 411708 388181 411772
rect 388115 411707 388181 411708
rect 386830 411030 386980 411090
rect 387104 411030 387258 411090
rect 388118 411060 388178 411707
rect 388302 411090 388362 413339
rect 393451 412860 393517 412861
rect 393451 412796 393452 412860
rect 393516 412796 393517 412860
rect 393451 412795 393517 412796
rect 389587 412724 389653 412725
rect 389587 412660 389588 412724
rect 389652 412660 389653 412724
rect 389587 412659 389653 412660
rect 390875 412724 390941 412725
rect 390875 412660 390876 412724
rect 390940 412660 390941 412724
rect 390875 412659 390941 412660
rect 391795 412724 391861 412725
rect 391795 412660 391796 412724
rect 391860 412660 391861 412724
rect 391795 412659 391861 412660
rect 393083 412724 393149 412725
rect 393083 412660 393084 412724
rect 393148 412660 393149 412724
rect 393083 412659 393149 412660
rect 389283 411500 389349 411501
rect 389283 411436 389284 411500
rect 389348 411436 389349 411500
rect 389283 411435 389349 411436
rect 388272 411030 388362 411090
rect 389286 411060 389346 411435
rect 389590 411090 389650 412659
rect 389440 411030 389650 411090
rect 389771 411092 389837 411093
rect 389771 411028 389772 411092
rect 389836 411090 389837 411092
rect 389836 411030 390484 411090
rect 389836 411028 389837 411030
rect 389771 411027 389837 411028
rect 390878 410750 390938 412659
rect 391059 411636 391125 411637
rect 391059 411572 391060 411636
rect 391124 411572 391125 411636
rect 391059 411571 391125 411572
rect 391062 411090 391122 411571
rect 391798 411090 391858 412659
rect 393086 411090 393146 412659
rect 391062 411030 391652 411090
rect 391776 411030 391858 411090
rect 392944 411030 393146 411090
rect 393454 411090 393514 412795
rect 394003 412724 394069 412725
rect 394003 412660 394004 412724
rect 394068 412660 394069 412724
rect 394003 412659 394069 412660
rect 394739 412724 394805 412725
rect 394739 412660 394740 412724
rect 394804 412660 394805 412724
rect 394739 412659 394805 412660
rect 395291 412724 395357 412725
rect 395291 412660 395292 412724
rect 395356 412660 395357 412724
rect 395291 412659 395357 412660
rect 396027 412724 396093 412725
rect 396027 412660 396028 412724
rect 396092 412660 396093 412724
rect 396027 412659 396093 412660
rect 394006 411634 394066 412659
rect 394006 411574 394142 411634
rect 393454 411030 393988 411090
rect 394082 411060 394142 411574
rect 394742 411090 394802 412659
rect 395294 411090 395354 412659
rect 394742 411030 395156 411090
rect 395280 411030 395354 411090
rect 372662 410690 372964 410750
rect 390608 410690 390938 410750
rect 396030 410750 396090 412659
rect 396398 411634 396458 413611
rect 397502 411770 397562 413611
rect 405779 413540 405845 413541
rect 405779 413476 405780 413540
rect 405844 413476 405845 413540
rect 405779 413475 405845 413476
rect 404675 413404 404741 413405
rect 404675 413340 404676 413404
rect 404740 413340 404741 413404
rect 404675 413339 404741 413340
rect 402283 413268 402349 413269
rect 402283 413204 402284 413268
rect 402348 413204 402349 413268
rect 402283 413203 402349 413204
rect 403387 413268 403453 413269
rect 403387 413204 403388 413268
rect 403452 413204 403453 413268
rect 403387 413203 403453 413204
rect 399891 413132 399957 413133
rect 399891 413068 399892 413132
rect 399956 413068 399957 413132
rect 399891 413067 399957 413068
rect 398603 412860 398669 412861
rect 398603 412796 398604 412860
rect 398668 412796 398669 412860
rect 398603 412795 398669 412796
rect 397502 411710 397646 411770
rect 397459 411636 397525 411637
rect 396398 411574 396478 411634
rect 396418 411060 396478 411574
rect 397459 411572 397460 411636
rect 397524 411572 397525 411636
rect 397459 411571 397525 411572
rect 397462 411060 397522 411571
rect 397586 411060 397646 411710
rect 398606 411634 398666 412795
rect 399155 411636 399221 411637
rect 398606 411574 398814 411634
rect 398051 411500 398117 411501
rect 398051 411436 398052 411500
rect 398116 411436 398117 411500
rect 398051 411435 398117 411436
rect 398054 411090 398114 411435
rect 398054 411030 398660 411090
rect 398754 411060 398814 411574
rect 399155 411572 399156 411636
rect 399220 411572 399221 411636
rect 399155 411571 399221 411572
rect 399158 411090 399218 411571
rect 399894 411498 399954 413067
rect 401179 412996 401245 412997
rect 401179 412932 401180 412996
rect 401244 412932 401245 412996
rect 401179 412931 401245 412932
rect 400963 411500 401029 411501
rect 399894 411438 399982 411498
rect 399158 411030 399828 411090
rect 399922 411060 399982 411438
rect 400963 411436 400964 411500
rect 401028 411436 401029 411500
rect 401182 411498 401242 412931
rect 400963 411435 401029 411436
rect 401090 411438 401242 411498
rect 400966 411060 401026 411435
rect 401090 411060 401150 411438
rect 401731 411364 401797 411365
rect 401731 411300 401732 411364
rect 401796 411300 401797 411364
rect 401731 411299 401797 411300
rect 401734 411090 401794 411299
rect 401734 411030 402164 411090
rect 402286 411030 402346 413203
rect 403390 411770 403450 413203
rect 404678 411770 404738 413339
rect 403390 411710 403486 411770
rect 403299 411500 403365 411501
rect 403299 411436 403300 411500
rect 403364 411436 403365 411500
rect 403299 411435 403365 411436
rect 403302 411060 403362 411435
rect 403426 411060 403486 411710
rect 404594 411710 404738 411770
rect 404307 411364 404373 411365
rect 404307 411300 404308 411364
rect 404372 411300 404373 411364
rect 404307 411299 404373 411300
rect 404310 411090 404370 411299
rect 404310 411030 404500 411090
rect 404594 411060 404654 411710
rect 405782 411030 405842 413475
rect 407435 413268 407501 413269
rect 407435 413204 407436 413268
rect 407500 413204 407501 413268
rect 407435 413203 407501 413204
rect 406331 412724 406397 412725
rect 406331 412660 406332 412724
rect 406396 412660 406397 412724
rect 406331 412659 406397 412660
rect 406334 411090 406394 412659
rect 407438 411090 407498 413203
rect 408723 413132 408789 413133
rect 408723 413068 408724 413132
rect 408788 413068 408789 413132
rect 408723 413067 408789 413068
rect 408726 411090 408786 413067
rect 412774 411090 412834 413747
rect 406334 411030 406960 411090
rect 407438 411030 408128 411090
rect 408726 411030 409296 411090
rect 412774 411030 413463 411090
rect 396030 410690 396324 410750
rect 392301 410412 392367 410413
rect 392301 410348 392302 410412
rect 392366 410410 392367 410412
rect 410011 410412 410077 410413
rect 392366 410350 392820 410410
rect 392366 410348 392367 410350
rect 392301 410347 392367 410348
rect 410011 410348 410012 410412
rect 410076 410410 410077 410412
rect 410076 410350 410464 410410
rect 410076 410348 410077 410350
rect 410011 410347 410077 410348
rect 335604 409018 335786 409254
rect 336022 409018 336204 409254
rect 335604 408934 336204 409018
rect 335604 408698 335786 408934
rect 336022 408698 336204 408934
rect 335604 373254 336204 408698
rect 340482 409254 340802 409276
rect 340482 409018 340524 409254
rect 340760 409018 340802 409254
rect 340482 408934 340802 409018
rect 340482 408698 340524 408934
rect 340760 408698 340802 408934
rect 340482 408676 340802 408698
rect 340482 405654 340802 405676
rect 340482 405418 340524 405654
rect 340760 405418 340802 405654
rect 340482 405334 340802 405418
rect 340482 405098 340524 405334
rect 340760 405098 340802 405334
rect 340482 405076 340802 405098
rect 340482 402054 340802 402076
rect 340482 401818 340524 402054
rect 340760 401818 340802 402054
rect 340482 401734 340802 401818
rect 340482 401498 340524 401734
rect 340760 401498 340802 401734
rect 340482 401476 340802 401498
rect 340482 398454 340802 398476
rect 340482 398218 340524 398454
rect 340760 398218 340802 398454
rect 340482 398134 340802 398218
rect 340482 397898 340524 398134
rect 340760 397898 340802 398134
rect 340482 397876 340802 397898
rect 340034 391254 340358 391276
rect 340034 391018 340078 391254
rect 340314 391018 340358 391254
rect 340034 390934 340358 391018
rect 340034 390698 340078 390934
rect 340314 390698 340358 390934
rect 340034 390676 340358 390698
rect 340034 387654 340358 387676
rect 340034 387418 340078 387654
rect 340314 387418 340358 387654
rect 340034 387334 340358 387418
rect 340034 387098 340078 387334
rect 340314 387098 340358 387334
rect 340034 387076 340358 387098
rect 422004 387654 422604 423098
rect 422004 387418 422186 387654
rect 422422 387418 422604 387654
rect 422004 387334 422604 387418
rect 422004 387098 422186 387334
rect 422422 387098 422604 387334
rect 340034 384054 340358 384076
rect 340034 383818 340078 384054
rect 340314 383818 340358 384054
rect 340034 383734 340358 383818
rect 340034 383498 340078 383734
rect 340314 383498 340358 383734
rect 340034 383476 340358 383498
rect 340034 380454 340358 380476
rect 340034 380218 340078 380454
rect 340314 380218 340358 380454
rect 340034 380134 340358 380218
rect 340034 379898 340078 380134
rect 340314 379898 340358 380134
rect 340034 379876 340358 379898
rect 335604 373018 335786 373254
rect 336022 373018 336204 373254
rect 335604 372934 336204 373018
rect 335604 372698 335786 372934
rect 336022 372698 336204 372934
rect 335604 337254 336204 372698
rect 340482 373254 340802 373276
rect 340482 373018 340524 373254
rect 340760 373018 340802 373254
rect 340482 372934 340802 373018
rect 340482 372698 340524 372934
rect 340760 372698 340802 372934
rect 340482 372676 340802 372698
rect 340482 369654 340802 369676
rect 340482 369418 340524 369654
rect 340760 369418 340802 369654
rect 340482 369334 340802 369418
rect 340482 369098 340524 369334
rect 340760 369098 340802 369334
rect 340482 369076 340802 369098
rect 340482 366054 340802 366076
rect 340482 365818 340524 366054
rect 340760 365818 340802 366054
rect 340482 365734 340802 365818
rect 340482 365498 340524 365734
rect 340760 365498 340802 365734
rect 340482 365476 340802 365498
rect 340482 362454 340802 362476
rect 340482 362218 340524 362454
rect 340760 362218 340802 362454
rect 340482 362134 340802 362218
rect 340482 361898 340524 362134
rect 340760 361898 340802 362134
rect 340482 361876 340802 361898
rect 340034 355254 340358 355276
rect 340034 355018 340078 355254
rect 340314 355018 340358 355254
rect 340034 354934 340358 355018
rect 340034 354698 340078 354934
rect 340314 354698 340358 354934
rect 340034 354676 340358 354698
rect 340034 351654 340358 351676
rect 340034 351418 340078 351654
rect 340314 351418 340358 351654
rect 340034 351334 340358 351418
rect 340034 351098 340078 351334
rect 340314 351098 340358 351334
rect 340034 351076 340358 351098
rect 422004 351654 422604 387098
rect 422004 351418 422186 351654
rect 422422 351418 422604 351654
rect 422004 351334 422604 351418
rect 422004 351098 422186 351334
rect 422422 351098 422604 351334
rect 340034 348054 340358 348076
rect 340034 347818 340078 348054
rect 340314 347818 340358 348054
rect 340034 347734 340358 347818
rect 340034 347498 340078 347734
rect 340314 347498 340358 347734
rect 340034 347476 340358 347498
rect 340034 344454 340358 344476
rect 340034 344218 340078 344454
rect 340314 344218 340358 344454
rect 340034 344134 340358 344218
rect 340034 343898 340078 344134
rect 340314 343898 340358 344134
rect 340034 343876 340358 343898
rect 335604 337018 335786 337254
rect 336022 337018 336204 337254
rect 335604 336934 336204 337018
rect 335604 336698 335786 336934
rect 336022 336698 336204 336934
rect 335604 301254 336204 336698
rect 340482 337254 340802 337276
rect 340482 337018 340524 337254
rect 340760 337018 340802 337254
rect 340482 336934 340802 337018
rect 340482 336698 340524 336934
rect 340760 336698 340802 336934
rect 340482 336676 340802 336698
rect 340482 333654 340802 333676
rect 340482 333418 340524 333654
rect 340760 333418 340802 333654
rect 340482 333334 340802 333418
rect 340482 333098 340524 333334
rect 340760 333098 340802 333334
rect 340482 333076 340802 333098
rect 340482 330054 340802 330076
rect 340482 329818 340524 330054
rect 340760 329818 340802 330054
rect 340482 329734 340802 329818
rect 340482 329498 340524 329734
rect 340760 329498 340802 329734
rect 340482 329476 340802 329498
rect 340482 326454 340802 326476
rect 340482 326218 340524 326454
rect 340760 326218 340802 326454
rect 340482 326134 340802 326218
rect 340482 325898 340524 326134
rect 340760 325898 340802 326134
rect 340482 325876 340802 325898
rect 343693 320430 344018 320490
rect 343958 318749 344018 320430
rect 348006 320250 348688 320310
rect 343955 318748 344021 318749
rect 343955 318684 343956 318748
rect 344020 318684 344021 318748
rect 343955 318683 344021 318684
rect 348006 318477 348066 320250
rect 348003 318476 348069 318477
rect 348003 318412 348004 318476
rect 348068 318412 348069 318476
rect 348003 318411 348069 318412
rect 335604 301018 335786 301254
rect 336022 301018 336204 301254
rect 335604 300934 336204 301018
rect 335604 300698 335786 300934
rect 336022 300698 336204 300934
rect 335604 265254 336204 300698
rect 335604 265018 335786 265254
rect 336022 265018 336204 265254
rect 335604 264934 336204 265018
rect 335604 264698 335786 264934
rect 336022 264698 336204 264934
rect 335604 229254 336204 264698
rect 335604 229018 335786 229254
rect 336022 229018 336204 229254
rect 335604 228934 336204 229018
rect 335604 228698 335786 228934
rect 336022 228698 336204 228934
rect 335604 193254 336204 228698
rect 335604 193018 335786 193254
rect 336022 193018 336204 193254
rect 335604 192934 336204 193018
rect 335604 192698 335786 192934
rect 336022 192698 336204 192934
rect 335604 157254 336204 192698
rect 335604 157018 335786 157254
rect 336022 157018 336204 157254
rect 335604 156934 336204 157018
rect 335604 156698 335786 156934
rect 336022 156698 336204 156934
rect 335604 121254 336204 156698
rect 335604 121018 335786 121254
rect 336022 121018 336204 121254
rect 335604 120934 336204 121018
rect 335604 120698 335786 120934
rect 336022 120698 336204 120934
rect 335604 85254 336204 120698
rect 335604 85018 335786 85254
rect 336022 85018 336204 85254
rect 335604 84934 336204 85018
rect 335604 84698 335786 84934
rect 336022 84698 336204 84934
rect 335604 49254 336204 84698
rect 335604 49018 335786 49254
rect 336022 49018 336204 49254
rect 335604 48934 336204 49018
rect 335604 48698 335786 48934
rect 336022 48698 336204 48934
rect 335604 13254 336204 48698
rect 335604 13018 335786 13254
rect 336022 13018 336204 13254
rect 335604 12934 336204 13018
rect 335604 12698 335786 12934
rect 336022 12698 336204 12934
rect 317604 -7162 317786 -6926
rect 318022 -7162 318204 -6926
rect 317604 -7246 318204 -7162
rect 317604 -7482 317786 -7246
rect 318022 -7482 318204 -7246
rect 317604 -7504 318204 -7482
rect 335604 -5986 336204 12698
rect 342804 308454 343404 317000
rect 342804 308218 342986 308454
rect 343222 308218 343404 308454
rect 342804 308134 343404 308218
rect 342804 307898 342986 308134
rect 343222 307898 343404 308134
rect 342804 272454 343404 307898
rect 342804 272218 342986 272454
rect 343222 272218 343404 272454
rect 342804 272134 343404 272218
rect 342804 271898 342986 272134
rect 343222 271898 343404 272134
rect 342804 236454 343404 271898
rect 342804 236218 342986 236454
rect 343222 236218 343404 236454
rect 342804 236134 343404 236218
rect 342804 235898 342986 236134
rect 343222 235898 343404 236134
rect 342804 200454 343404 235898
rect 342804 200218 342986 200454
rect 343222 200218 343404 200454
rect 342804 200134 343404 200218
rect 342804 199898 342986 200134
rect 343222 199898 343404 200134
rect 342804 164454 343404 199898
rect 342804 164218 342986 164454
rect 343222 164218 343404 164454
rect 342804 164134 343404 164218
rect 342804 163898 342986 164134
rect 343222 163898 343404 164134
rect 342804 128454 343404 163898
rect 342804 128218 342986 128454
rect 343222 128218 343404 128454
rect 342804 128134 343404 128218
rect 342804 127898 342986 128134
rect 343222 127898 343404 128134
rect 342804 92454 343404 127898
rect 342804 92218 342986 92454
rect 343222 92218 343404 92454
rect 342804 92134 343404 92218
rect 342804 91898 342986 92134
rect 343222 91898 343404 92134
rect 342804 56454 343404 91898
rect 342804 56218 342986 56454
rect 343222 56218 343404 56454
rect 342804 56134 343404 56218
rect 342804 55898 342986 56134
rect 343222 55898 343404 56134
rect 342804 20454 343404 55898
rect 342804 20218 342986 20454
rect 343222 20218 343404 20454
rect 342804 20134 343404 20218
rect 342804 19898 342986 20134
rect 343222 19898 343404 20134
rect 342804 -1286 343404 19898
rect 342804 -1522 342986 -1286
rect 343222 -1522 343404 -1286
rect 342804 -1606 343404 -1522
rect 342804 -1842 342986 -1606
rect 343222 -1842 343404 -1606
rect 342804 -1864 343404 -1842
rect 346404 312054 347004 317000
rect 346404 311818 346586 312054
rect 346822 311818 347004 312054
rect 346404 311734 347004 311818
rect 346404 311498 346586 311734
rect 346822 311498 347004 311734
rect 346404 276054 347004 311498
rect 346404 275818 346586 276054
rect 346822 275818 347004 276054
rect 346404 275734 347004 275818
rect 346404 275498 346586 275734
rect 346822 275498 347004 275734
rect 346404 240054 347004 275498
rect 346404 239818 346586 240054
rect 346822 239818 347004 240054
rect 346404 239734 347004 239818
rect 346404 239498 346586 239734
rect 346822 239498 347004 239734
rect 346404 204054 347004 239498
rect 346404 203818 346586 204054
rect 346822 203818 347004 204054
rect 346404 203734 347004 203818
rect 346404 203498 346586 203734
rect 346822 203498 347004 203734
rect 346404 168054 347004 203498
rect 346404 167818 346586 168054
rect 346822 167818 347004 168054
rect 346404 167734 347004 167818
rect 346404 167498 346586 167734
rect 346822 167498 347004 167734
rect 346404 132054 347004 167498
rect 346404 131818 346586 132054
rect 346822 131818 347004 132054
rect 346404 131734 347004 131818
rect 346404 131498 346586 131734
rect 346822 131498 347004 131734
rect 346404 96054 347004 131498
rect 346404 95818 346586 96054
rect 346822 95818 347004 96054
rect 346404 95734 347004 95818
rect 346404 95498 346586 95734
rect 346822 95498 347004 95734
rect 346404 60054 347004 95498
rect 346404 59818 346586 60054
rect 346822 59818 347004 60054
rect 346404 59734 347004 59818
rect 346404 59498 346586 59734
rect 346822 59498 347004 59734
rect 346404 24054 347004 59498
rect 346404 23818 346586 24054
rect 346822 23818 347004 24054
rect 346404 23734 347004 23818
rect 346404 23498 346586 23734
rect 346822 23498 347004 23734
rect 346404 -3166 347004 23498
rect 346404 -3402 346586 -3166
rect 346822 -3402 347004 -3166
rect 346404 -3486 347004 -3402
rect 346404 -3722 346586 -3486
rect 346822 -3722 347004 -3486
rect 346404 -3744 347004 -3722
rect 350004 315654 350604 317000
rect 350004 315418 350186 315654
rect 350422 315418 350604 315654
rect 350004 315334 350604 315418
rect 350004 315098 350186 315334
rect 350422 315098 350604 315334
rect 350004 279654 350604 315098
rect 350004 279418 350186 279654
rect 350422 279418 350604 279654
rect 350004 279334 350604 279418
rect 350004 279098 350186 279334
rect 350422 279098 350604 279334
rect 350004 243654 350604 279098
rect 350004 243418 350186 243654
rect 350422 243418 350604 243654
rect 350004 243334 350604 243418
rect 350004 243098 350186 243334
rect 350422 243098 350604 243334
rect 350004 207654 350604 243098
rect 350004 207418 350186 207654
rect 350422 207418 350604 207654
rect 350004 207334 350604 207418
rect 350004 207098 350186 207334
rect 350422 207098 350604 207334
rect 350004 171654 350604 207098
rect 350004 171418 350186 171654
rect 350422 171418 350604 171654
rect 350004 171334 350604 171418
rect 350004 171098 350186 171334
rect 350422 171098 350604 171334
rect 350004 135654 350604 171098
rect 350004 135418 350186 135654
rect 350422 135418 350604 135654
rect 350004 135334 350604 135418
rect 350004 135098 350186 135334
rect 350422 135098 350604 135334
rect 350004 99654 350604 135098
rect 350004 99418 350186 99654
rect 350422 99418 350604 99654
rect 350004 99334 350604 99418
rect 350004 99098 350186 99334
rect 350422 99098 350604 99334
rect 350004 63654 350604 99098
rect 350004 63418 350186 63654
rect 350422 63418 350604 63654
rect 350004 63334 350604 63418
rect 350004 63098 350186 63334
rect 350422 63098 350604 63334
rect 350004 27654 350604 63098
rect 350004 27418 350186 27654
rect 350422 27418 350604 27654
rect 350004 27334 350604 27418
rect 350004 27098 350186 27334
rect 350422 27098 350604 27334
rect 350004 -5046 350604 27098
rect 350004 -5282 350186 -5046
rect 350422 -5282 350604 -5046
rect 350004 -5366 350604 -5282
rect 350004 -5602 350186 -5366
rect 350422 -5602 350604 -5366
rect 350004 -5624 350604 -5602
rect 353604 283254 354204 317000
rect 353604 283018 353786 283254
rect 354022 283018 354204 283254
rect 353604 282934 354204 283018
rect 353604 282698 353786 282934
rect 354022 282698 354204 282934
rect 353604 247254 354204 282698
rect 353604 247018 353786 247254
rect 354022 247018 354204 247254
rect 353604 246934 354204 247018
rect 353604 246698 353786 246934
rect 354022 246698 354204 246934
rect 353604 211254 354204 246698
rect 353604 211018 353786 211254
rect 354022 211018 354204 211254
rect 353604 210934 354204 211018
rect 353604 210698 353786 210934
rect 354022 210698 354204 210934
rect 353604 175254 354204 210698
rect 353604 175018 353786 175254
rect 354022 175018 354204 175254
rect 353604 174934 354204 175018
rect 353604 174698 353786 174934
rect 354022 174698 354204 174934
rect 353604 139254 354204 174698
rect 353604 139018 353786 139254
rect 354022 139018 354204 139254
rect 353604 138934 354204 139018
rect 353604 138698 353786 138934
rect 354022 138698 354204 138934
rect 353604 103254 354204 138698
rect 353604 103018 353786 103254
rect 354022 103018 354204 103254
rect 353604 102934 354204 103018
rect 353604 102698 353786 102934
rect 354022 102698 354204 102934
rect 353604 67254 354204 102698
rect 353604 67018 353786 67254
rect 354022 67018 354204 67254
rect 353604 66934 354204 67018
rect 353604 66698 353786 66934
rect 354022 66698 354204 66934
rect 353604 31254 354204 66698
rect 353604 31018 353786 31254
rect 354022 31018 354204 31254
rect 353604 30934 354204 31018
rect 353604 30698 353786 30934
rect 354022 30698 354204 30934
rect 335604 -6222 335786 -5986
rect 336022 -6222 336204 -5986
rect 335604 -6306 336204 -6222
rect 335604 -6542 335786 -6306
rect 336022 -6542 336204 -6306
rect 335604 -7504 336204 -6542
rect 353604 -6926 354204 30698
rect 360804 290454 361404 317000
rect 360804 290218 360986 290454
rect 361222 290218 361404 290454
rect 360804 290134 361404 290218
rect 360804 289898 360986 290134
rect 361222 289898 361404 290134
rect 360804 254454 361404 289898
rect 360804 254218 360986 254454
rect 361222 254218 361404 254454
rect 360804 254134 361404 254218
rect 360804 253898 360986 254134
rect 361222 253898 361404 254134
rect 360804 218454 361404 253898
rect 360804 218218 360986 218454
rect 361222 218218 361404 218454
rect 360804 218134 361404 218218
rect 360804 217898 360986 218134
rect 361222 217898 361404 218134
rect 360804 182454 361404 217898
rect 360804 182218 360986 182454
rect 361222 182218 361404 182454
rect 360804 182134 361404 182218
rect 360804 181898 360986 182134
rect 361222 181898 361404 182134
rect 360804 146454 361404 181898
rect 360804 146218 360986 146454
rect 361222 146218 361404 146454
rect 360804 146134 361404 146218
rect 360804 145898 360986 146134
rect 361222 145898 361404 146134
rect 360804 110454 361404 145898
rect 360804 110218 360986 110454
rect 361222 110218 361404 110454
rect 360804 110134 361404 110218
rect 360804 109898 360986 110134
rect 361222 109898 361404 110134
rect 360804 74454 361404 109898
rect 360804 74218 360986 74454
rect 361222 74218 361404 74454
rect 360804 74134 361404 74218
rect 360804 73898 360986 74134
rect 361222 73898 361404 74134
rect 360804 38454 361404 73898
rect 360804 38218 360986 38454
rect 361222 38218 361404 38454
rect 360804 38134 361404 38218
rect 360804 37898 360986 38134
rect 361222 37898 361404 38134
rect 360804 2454 361404 37898
rect 360804 2218 360986 2454
rect 361222 2218 361404 2454
rect 360804 2134 361404 2218
rect 360804 1898 360986 2134
rect 361222 1898 361404 2134
rect 360804 -346 361404 1898
rect 360804 -582 360986 -346
rect 361222 -582 361404 -346
rect 360804 -666 361404 -582
rect 360804 -902 360986 -666
rect 361222 -902 361404 -666
rect 360804 -1864 361404 -902
rect 364404 294054 365004 317000
rect 364404 293818 364586 294054
rect 364822 293818 365004 294054
rect 364404 293734 365004 293818
rect 364404 293498 364586 293734
rect 364822 293498 365004 293734
rect 364404 258054 365004 293498
rect 364404 257818 364586 258054
rect 364822 257818 365004 258054
rect 364404 257734 365004 257818
rect 364404 257498 364586 257734
rect 364822 257498 365004 257734
rect 364404 222054 365004 257498
rect 364404 221818 364586 222054
rect 364822 221818 365004 222054
rect 364404 221734 365004 221818
rect 364404 221498 364586 221734
rect 364822 221498 365004 221734
rect 364404 186054 365004 221498
rect 364404 185818 364586 186054
rect 364822 185818 365004 186054
rect 364404 185734 365004 185818
rect 364404 185498 364586 185734
rect 364822 185498 365004 185734
rect 364404 150054 365004 185498
rect 364404 149818 364586 150054
rect 364822 149818 365004 150054
rect 364404 149734 365004 149818
rect 364404 149498 364586 149734
rect 364822 149498 365004 149734
rect 364404 114054 365004 149498
rect 364404 113818 364586 114054
rect 364822 113818 365004 114054
rect 364404 113734 365004 113818
rect 364404 113498 364586 113734
rect 364822 113498 365004 113734
rect 364404 78054 365004 113498
rect 364404 77818 364586 78054
rect 364822 77818 365004 78054
rect 364404 77734 365004 77818
rect 364404 77498 364586 77734
rect 364822 77498 365004 77734
rect 364404 42054 365004 77498
rect 364404 41818 364586 42054
rect 364822 41818 365004 42054
rect 364404 41734 365004 41818
rect 364404 41498 364586 41734
rect 364822 41498 365004 41734
rect 364404 6054 365004 41498
rect 364404 5818 364586 6054
rect 364822 5818 365004 6054
rect 364404 5734 365004 5818
rect 364404 5498 364586 5734
rect 364822 5498 365004 5734
rect 364404 -2226 365004 5498
rect 364404 -2462 364586 -2226
rect 364822 -2462 365004 -2226
rect 364404 -2546 365004 -2462
rect 364404 -2782 364586 -2546
rect 364822 -2782 365004 -2546
rect 364404 -3744 365004 -2782
rect 368004 297654 368604 317000
rect 368004 297418 368186 297654
rect 368422 297418 368604 297654
rect 368004 297334 368604 297418
rect 368004 297098 368186 297334
rect 368422 297098 368604 297334
rect 368004 261654 368604 297098
rect 368004 261418 368186 261654
rect 368422 261418 368604 261654
rect 368004 261334 368604 261418
rect 368004 261098 368186 261334
rect 368422 261098 368604 261334
rect 368004 225654 368604 261098
rect 368004 225418 368186 225654
rect 368422 225418 368604 225654
rect 368004 225334 368604 225418
rect 368004 225098 368186 225334
rect 368422 225098 368604 225334
rect 368004 189654 368604 225098
rect 368004 189418 368186 189654
rect 368422 189418 368604 189654
rect 368004 189334 368604 189418
rect 368004 189098 368186 189334
rect 368422 189098 368604 189334
rect 368004 153654 368604 189098
rect 368004 153418 368186 153654
rect 368422 153418 368604 153654
rect 368004 153334 368604 153418
rect 368004 153098 368186 153334
rect 368422 153098 368604 153334
rect 368004 117654 368604 153098
rect 368004 117418 368186 117654
rect 368422 117418 368604 117654
rect 368004 117334 368604 117418
rect 368004 117098 368186 117334
rect 368422 117098 368604 117334
rect 368004 81654 368604 117098
rect 368004 81418 368186 81654
rect 368422 81418 368604 81654
rect 368004 81334 368604 81418
rect 368004 81098 368186 81334
rect 368422 81098 368604 81334
rect 368004 45654 368604 81098
rect 368004 45418 368186 45654
rect 368422 45418 368604 45654
rect 368004 45334 368604 45418
rect 368004 45098 368186 45334
rect 368422 45098 368604 45334
rect 368004 9654 368604 45098
rect 368004 9418 368186 9654
rect 368422 9418 368604 9654
rect 368004 9334 368604 9418
rect 368004 9098 368186 9334
rect 368422 9098 368604 9334
rect 368004 -4106 368604 9098
rect 368004 -4342 368186 -4106
rect 368422 -4342 368604 -4106
rect 368004 -4426 368604 -4342
rect 368004 -4662 368186 -4426
rect 368422 -4662 368604 -4426
rect 368004 -5624 368604 -4662
rect 371604 301254 372204 317000
rect 371604 301018 371786 301254
rect 372022 301018 372204 301254
rect 371604 300934 372204 301018
rect 371604 300698 371786 300934
rect 372022 300698 372204 300934
rect 371604 265254 372204 300698
rect 371604 265018 371786 265254
rect 372022 265018 372204 265254
rect 371604 264934 372204 265018
rect 371604 264698 371786 264934
rect 372022 264698 372204 264934
rect 371604 229254 372204 264698
rect 371604 229018 371786 229254
rect 372022 229018 372204 229254
rect 371604 228934 372204 229018
rect 371604 228698 371786 228934
rect 372022 228698 372204 228934
rect 371604 193254 372204 228698
rect 371604 193018 371786 193254
rect 372022 193018 372204 193254
rect 371604 192934 372204 193018
rect 371604 192698 371786 192934
rect 372022 192698 372204 192934
rect 371604 157254 372204 192698
rect 371604 157018 371786 157254
rect 372022 157018 372204 157254
rect 371604 156934 372204 157018
rect 371604 156698 371786 156934
rect 372022 156698 372204 156934
rect 371604 121254 372204 156698
rect 371604 121018 371786 121254
rect 372022 121018 372204 121254
rect 371604 120934 372204 121018
rect 371604 120698 371786 120934
rect 372022 120698 372204 120934
rect 371604 85254 372204 120698
rect 371604 85018 371786 85254
rect 372022 85018 372204 85254
rect 371604 84934 372204 85018
rect 371604 84698 371786 84934
rect 372022 84698 372204 84934
rect 371604 49254 372204 84698
rect 371604 49018 371786 49254
rect 372022 49018 372204 49254
rect 371604 48934 372204 49018
rect 371604 48698 371786 48934
rect 372022 48698 372204 48934
rect 371604 13254 372204 48698
rect 371604 13018 371786 13254
rect 372022 13018 372204 13254
rect 371604 12934 372204 13018
rect 371604 12698 371786 12934
rect 372022 12698 372204 12934
rect 353604 -7162 353786 -6926
rect 354022 -7162 354204 -6926
rect 353604 -7246 354204 -7162
rect 353604 -7482 353786 -7246
rect 354022 -7482 354204 -7246
rect 353604 -7504 354204 -7482
rect 371604 -5986 372204 12698
rect 378804 308454 379404 317000
rect 378804 308218 378986 308454
rect 379222 308218 379404 308454
rect 378804 308134 379404 308218
rect 378804 307898 378986 308134
rect 379222 307898 379404 308134
rect 378804 272454 379404 307898
rect 378804 272218 378986 272454
rect 379222 272218 379404 272454
rect 378804 272134 379404 272218
rect 378804 271898 378986 272134
rect 379222 271898 379404 272134
rect 378804 236454 379404 271898
rect 378804 236218 378986 236454
rect 379222 236218 379404 236454
rect 378804 236134 379404 236218
rect 378804 235898 378986 236134
rect 379222 235898 379404 236134
rect 378804 200454 379404 235898
rect 378804 200218 378986 200454
rect 379222 200218 379404 200454
rect 378804 200134 379404 200218
rect 378804 199898 378986 200134
rect 379222 199898 379404 200134
rect 378804 164454 379404 199898
rect 378804 164218 378986 164454
rect 379222 164218 379404 164454
rect 378804 164134 379404 164218
rect 378804 163898 378986 164134
rect 379222 163898 379404 164134
rect 378804 128454 379404 163898
rect 378804 128218 378986 128454
rect 379222 128218 379404 128454
rect 378804 128134 379404 128218
rect 378804 127898 378986 128134
rect 379222 127898 379404 128134
rect 378804 92454 379404 127898
rect 378804 92218 378986 92454
rect 379222 92218 379404 92454
rect 378804 92134 379404 92218
rect 378804 91898 378986 92134
rect 379222 91898 379404 92134
rect 378804 56454 379404 91898
rect 378804 56218 378986 56454
rect 379222 56218 379404 56454
rect 378804 56134 379404 56218
rect 378804 55898 378986 56134
rect 379222 55898 379404 56134
rect 378804 20454 379404 55898
rect 378804 20218 378986 20454
rect 379222 20218 379404 20454
rect 378804 20134 379404 20218
rect 378804 19898 378986 20134
rect 379222 19898 379404 20134
rect 378804 -1286 379404 19898
rect 378804 -1522 378986 -1286
rect 379222 -1522 379404 -1286
rect 378804 -1606 379404 -1522
rect 378804 -1842 378986 -1606
rect 379222 -1842 379404 -1606
rect 378804 -1864 379404 -1842
rect 382404 312054 383004 317000
rect 382404 311818 382586 312054
rect 382822 311818 383004 312054
rect 382404 311734 383004 311818
rect 382404 311498 382586 311734
rect 382822 311498 383004 311734
rect 382404 276054 383004 311498
rect 382404 275818 382586 276054
rect 382822 275818 383004 276054
rect 382404 275734 383004 275818
rect 382404 275498 382586 275734
rect 382822 275498 383004 275734
rect 382404 240054 383004 275498
rect 382404 239818 382586 240054
rect 382822 239818 383004 240054
rect 382404 239734 383004 239818
rect 382404 239498 382586 239734
rect 382822 239498 383004 239734
rect 382404 204054 383004 239498
rect 382404 203818 382586 204054
rect 382822 203818 383004 204054
rect 382404 203734 383004 203818
rect 382404 203498 382586 203734
rect 382822 203498 383004 203734
rect 382404 168054 383004 203498
rect 382404 167818 382586 168054
rect 382822 167818 383004 168054
rect 382404 167734 383004 167818
rect 382404 167498 382586 167734
rect 382822 167498 383004 167734
rect 382404 132054 383004 167498
rect 382404 131818 382586 132054
rect 382822 131818 383004 132054
rect 382404 131734 383004 131818
rect 382404 131498 382586 131734
rect 382822 131498 383004 131734
rect 382404 96054 383004 131498
rect 382404 95818 382586 96054
rect 382822 95818 383004 96054
rect 382404 95734 383004 95818
rect 382404 95498 382586 95734
rect 382822 95498 383004 95734
rect 382404 60054 383004 95498
rect 382404 59818 382586 60054
rect 382822 59818 383004 60054
rect 382404 59734 383004 59818
rect 382404 59498 382586 59734
rect 382822 59498 383004 59734
rect 382404 24054 383004 59498
rect 382404 23818 382586 24054
rect 382822 23818 383004 24054
rect 382404 23734 383004 23818
rect 382404 23498 382586 23734
rect 382822 23498 383004 23734
rect 382404 -3166 383004 23498
rect 382404 -3402 382586 -3166
rect 382822 -3402 383004 -3166
rect 382404 -3486 383004 -3402
rect 382404 -3722 382586 -3486
rect 382822 -3722 383004 -3486
rect 382404 -3744 383004 -3722
rect 386004 315654 386604 317000
rect 386004 315418 386186 315654
rect 386422 315418 386604 315654
rect 386004 315334 386604 315418
rect 386004 315098 386186 315334
rect 386422 315098 386604 315334
rect 386004 279654 386604 315098
rect 386004 279418 386186 279654
rect 386422 279418 386604 279654
rect 386004 279334 386604 279418
rect 386004 279098 386186 279334
rect 386422 279098 386604 279334
rect 386004 243654 386604 279098
rect 386004 243418 386186 243654
rect 386422 243418 386604 243654
rect 386004 243334 386604 243418
rect 386004 243098 386186 243334
rect 386422 243098 386604 243334
rect 386004 207654 386604 243098
rect 386004 207418 386186 207654
rect 386422 207418 386604 207654
rect 386004 207334 386604 207418
rect 386004 207098 386186 207334
rect 386422 207098 386604 207334
rect 386004 171654 386604 207098
rect 386004 171418 386186 171654
rect 386422 171418 386604 171654
rect 386004 171334 386604 171418
rect 386004 171098 386186 171334
rect 386422 171098 386604 171334
rect 386004 135654 386604 171098
rect 386004 135418 386186 135654
rect 386422 135418 386604 135654
rect 386004 135334 386604 135418
rect 386004 135098 386186 135334
rect 386422 135098 386604 135334
rect 386004 99654 386604 135098
rect 386004 99418 386186 99654
rect 386422 99418 386604 99654
rect 386004 99334 386604 99418
rect 386004 99098 386186 99334
rect 386422 99098 386604 99334
rect 386004 63654 386604 99098
rect 386004 63418 386186 63654
rect 386422 63418 386604 63654
rect 386004 63334 386604 63418
rect 386004 63098 386186 63334
rect 386422 63098 386604 63334
rect 386004 27654 386604 63098
rect 386004 27418 386186 27654
rect 386422 27418 386604 27654
rect 386004 27334 386604 27418
rect 386004 27098 386186 27334
rect 386422 27098 386604 27334
rect 386004 -5046 386604 27098
rect 386004 -5282 386186 -5046
rect 386422 -5282 386604 -5046
rect 386004 -5366 386604 -5282
rect 386004 -5602 386186 -5366
rect 386422 -5602 386604 -5366
rect 386004 -5624 386604 -5602
rect 389604 283254 390204 317000
rect 389604 283018 389786 283254
rect 390022 283018 390204 283254
rect 389604 282934 390204 283018
rect 389604 282698 389786 282934
rect 390022 282698 390204 282934
rect 389604 247254 390204 282698
rect 389604 247018 389786 247254
rect 390022 247018 390204 247254
rect 389604 246934 390204 247018
rect 389604 246698 389786 246934
rect 390022 246698 390204 246934
rect 389604 211254 390204 246698
rect 389604 211018 389786 211254
rect 390022 211018 390204 211254
rect 389604 210934 390204 211018
rect 389604 210698 389786 210934
rect 390022 210698 390204 210934
rect 389604 175254 390204 210698
rect 389604 175018 389786 175254
rect 390022 175018 390204 175254
rect 389604 174934 390204 175018
rect 389604 174698 389786 174934
rect 390022 174698 390204 174934
rect 389604 139254 390204 174698
rect 389604 139018 389786 139254
rect 390022 139018 390204 139254
rect 389604 138934 390204 139018
rect 389604 138698 389786 138934
rect 390022 138698 390204 138934
rect 389604 103254 390204 138698
rect 389604 103018 389786 103254
rect 390022 103018 390204 103254
rect 389604 102934 390204 103018
rect 389604 102698 389786 102934
rect 390022 102698 390204 102934
rect 389604 67254 390204 102698
rect 389604 67018 389786 67254
rect 390022 67018 390204 67254
rect 389604 66934 390204 67018
rect 389604 66698 389786 66934
rect 390022 66698 390204 66934
rect 389604 31254 390204 66698
rect 389604 31018 389786 31254
rect 390022 31018 390204 31254
rect 389604 30934 390204 31018
rect 389604 30698 389786 30934
rect 390022 30698 390204 30934
rect 371604 -6222 371786 -5986
rect 372022 -6222 372204 -5986
rect 371604 -6306 372204 -6222
rect 371604 -6542 371786 -6306
rect 372022 -6542 372204 -6306
rect 371604 -7504 372204 -6542
rect 389604 -6926 390204 30698
rect 396804 290454 397404 317000
rect 396804 290218 396986 290454
rect 397222 290218 397404 290454
rect 396804 290134 397404 290218
rect 396804 289898 396986 290134
rect 397222 289898 397404 290134
rect 396804 254454 397404 289898
rect 396804 254218 396986 254454
rect 397222 254218 397404 254454
rect 396804 254134 397404 254218
rect 396804 253898 396986 254134
rect 397222 253898 397404 254134
rect 396804 218454 397404 253898
rect 396804 218218 396986 218454
rect 397222 218218 397404 218454
rect 396804 218134 397404 218218
rect 396804 217898 396986 218134
rect 397222 217898 397404 218134
rect 396804 182454 397404 217898
rect 396804 182218 396986 182454
rect 397222 182218 397404 182454
rect 396804 182134 397404 182218
rect 396804 181898 396986 182134
rect 397222 181898 397404 182134
rect 396804 146454 397404 181898
rect 396804 146218 396986 146454
rect 397222 146218 397404 146454
rect 396804 146134 397404 146218
rect 396804 145898 396986 146134
rect 397222 145898 397404 146134
rect 396804 110454 397404 145898
rect 396804 110218 396986 110454
rect 397222 110218 397404 110454
rect 396804 110134 397404 110218
rect 396804 109898 396986 110134
rect 397222 109898 397404 110134
rect 396804 74454 397404 109898
rect 396804 74218 396986 74454
rect 397222 74218 397404 74454
rect 396804 74134 397404 74218
rect 396804 73898 396986 74134
rect 397222 73898 397404 74134
rect 396804 38454 397404 73898
rect 396804 38218 396986 38454
rect 397222 38218 397404 38454
rect 396804 38134 397404 38218
rect 396804 37898 396986 38134
rect 397222 37898 397404 38134
rect 396804 2454 397404 37898
rect 396804 2218 396986 2454
rect 397222 2218 397404 2454
rect 396804 2134 397404 2218
rect 396804 1898 396986 2134
rect 397222 1898 397404 2134
rect 396804 -346 397404 1898
rect 396804 -582 396986 -346
rect 397222 -582 397404 -346
rect 396804 -666 397404 -582
rect 396804 -902 396986 -666
rect 397222 -902 397404 -666
rect 396804 -1864 397404 -902
rect 400404 294054 401004 317000
rect 400404 293818 400586 294054
rect 400822 293818 401004 294054
rect 400404 293734 401004 293818
rect 400404 293498 400586 293734
rect 400822 293498 401004 293734
rect 400404 258054 401004 293498
rect 400404 257818 400586 258054
rect 400822 257818 401004 258054
rect 400404 257734 401004 257818
rect 400404 257498 400586 257734
rect 400822 257498 401004 257734
rect 400404 222054 401004 257498
rect 400404 221818 400586 222054
rect 400822 221818 401004 222054
rect 400404 221734 401004 221818
rect 400404 221498 400586 221734
rect 400822 221498 401004 221734
rect 400404 186054 401004 221498
rect 400404 185818 400586 186054
rect 400822 185818 401004 186054
rect 400404 185734 401004 185818
rect 400404 185498 400586 185734
rect 400822 185498 401004 185734
rect 400404 150054 401004 185498
rect 400404 149818 400586 150054
rect 400822 149818 401004 150054
rect 400404 149734 401004 149818
rect 400404 149498 400586 149734
rect 400822 149498 401004 149734
rect 400404 114054 401004 149498
rect 400404 113818 400586 114054
rect 400822 113818 401004 114054
rect 400404 113734 401004 113818
rect 400404 113498 400586 113734
rect 400822 113498 401004 113734
rect 400404 78054 401004 113498
rect 400404 77818 400586 78054
rect 400822 77818 401004 78054
rect 400404 77734 401004 77818
rect 400404 77498 400586 77734
rect 400822 77498 401004 77734
rect 400404 42054 401004 77498
rect 400404 41818 400586 42054
rect 400822 41818 401004 42054
rect 400404 41734 401004 41818
rect 400404 41498 400586 41734
rect 400822 41498 401004 41734
rect 400404 6054 401004 41498
rect 400404 5818 400586 6054
rect 400822 5818 401004 6054
rect 400404 5734 401004 5818
rect 400404 5498 400586 5734
rect 400822 5498 401004 5734
rect 400404 -2226 401004 5498
rect 400404 -2462 400586 -2226
rect 400822 -2462 401004 -2226
rect 400404 -2546 401004 -2462
rect 400404 -2782 400586 -2546
rect 400822 -2782 401004 -2546
rect 400404 -3744 401004 -2782
rect 404004 297654 404604 317000
rect 404004 297418 404186 297654
rect 404422 297418 404604 297654
rect 404004 297334 404604 297418
rect 404004 297098 404186 297334
rect 404422 297098 404604 297334
rect 404004 261654 404604 297098
rect 404004 261418 404186 261654
rect 404422 261418 404604 261654
rect 404004 261334 404604 261418
rect 404004 261098 404186 261334
rect 404422 261098 404604 261334
rect 404004 225654 404604 261098
rect 404004 225418 404186 225654
rect 404422 225418 404604 225654
rect 404004 225334 404604 225418
rect 404004 225098 404186 225334
rect 404422 225098 404604 225334
rect 404004 189654 404604 225098
rect 404004 189418 404186 189654
rect 404422 189418 404604 189654
rect 404004 189334 404604 189418
rect 404004 189098 404186 189334
rect 404422 189098 404604 189334
rect 404004 153654 404604 189098
rect 404004 153418 404186 153654
rect 404422 153418 404604 153654
rect 404004 153334 404604 153418
rect 404004 153098 404186 153334
rect 404422 153098 404604 153334
rect 404004 117654 404604 153098
rect 404004 117418 404186 117654
rect 404422 117418 404604 117654
rect 404004 117334 404604 117418
rect 404004 117098 404186 117334
rect 404422 117098 404604 117334
rect 404004 81654 404604 117098
rect 404004 81418 404186 81654
rect 404422 81418 404604 81654
rect 404004 81334 404604 81418
rect 404004 81098 404186 81334
rect 404422 81098 404604 81334
rect 404004 45654 404604 81098
rect 404004 45418 404186 45654
rect 404422 45418 404604 45654
rect 404004 45334 404604 45418
rect 404004 45098 404186 45334
rect 404422 45098 404604 45334
rect 404004 9654 404604 45098
rect 404004 9418 404186 9654
rect 404422 9418 404604 9654
rect 404004 9334 404604 9418
rect 404004 9098 404186 9334
rect 404422 9098 404604 9334
rect 404004 -4106 404604 9098
rect 404004 -4342 404186 -4106
rect 404422 -4342 404604 -4106
rect 404004 -4426 404604 -4342
rect 404004 -4662 404186 -4426
rect 404422 -4662 404604 -4426
rect 404004 -5624 404604 -4662
rect 407604 301254 408204 317000
rect 407604 301018 407786 301254
rect 408022 301018 408204 301254
rect 407604 300934 408204 301018
rect 407604 300698 407786 300934
rect 408022 300698 408204 300934
rect 407604 265254 408204 300698
rect 407604 265018 407786 265254
rect 408022 265018 408204 265254
rect 407604 264934 408204 265018
rect 407604 264698 407786 264934
rect 408022 264698 408204 264934
rect 407604 229254 408204 264698
rect 407604 229018 407786 229254
rect 408022 229018 408204 229254
rect 407604 228934 408204 229018
rect 407604 228698 407786 228934
rect 408022 228698 408204 228934
rect 407604 193254 408204 228698
rect 407604 193018 407786 193254
rect 408022 193018 408204 193254
rect 407604 192934 408204 193018
rect 407604 192698 407786 192934
rect 408022 192698 408204 192934
rect 407604 157254 408204 192698
rect 407604 157018 407786 157254
rect 408022 157018 408204 157254
rect 407604 156934 408204 157018
rect 407604 156698 407786 156934
rect 408022 156698 408204 156934
rect 407604 121254 408204 156698
rect 407604 121018 407786 121254
rect 408022 121018 408204 121254
rect 407604 120934 408204 121018
rect 407604 120698 407786 120934
rect 408022 120698 408204 120934
rect 407604 85254 408204 120698
rect 407604 85018 407786 85254
rect 408022 85018 408204 85254
rect 407604 84934 408204 85018
rect 407604 84698 407786 84934
rect 408022 84698 408204 84934
rect 407604 49254 408204 84698
rect 407604 49018 407786 49254
rect 408022 49018 408204 49254
rect 407604 48934 408204 49018
rect 407604 48698 407786 48934
rect 408022 48698 408204 48934
rect 407604 13254 408204 48698
rect 407604 13018 407786 13254
rect 408022 13018 408204 13254
rect 407604 12934 408204 13018
rect 407604 12698 407786 12934
rect 408022 12698 408204 12934
rect 389604 -7162 389786 -6926
rect 390022 -7162 390204 -6926
rect 389604 -7246 390204 -7162
rect 389604 -7482 389786 -7246
rect 390022 -7482 390204 -7246
rect 389604 -7504 390204 -7482
rect 407604 -5986 408204 12698
rect 414804 308454 415404 317000
rect 414804 308218 414986 308454
rect 415222 308218 415404 308454
rect 414804 308134 415404 308218
rect 414804 307898 414986 308134
rect 415222 307898 415404 308134
rect 414804 272454 415404 307898
rect 414804 272218 414986 272454
rect 415222 272218 415404 272454
rect 414804 272134 415404 272218
rect 414804 271898 414986 272134
rect 415222 271898 415404 272134
rect 414804 236454 415404 271898
rect 414804 236218 414986 236454
rect 415222 236218 415404 236454
rect 414804 236134 415404 236218
rect 414804 235898 414986 236134
rect 415222 235898 415404 236134
rect 414804 200454 415404 235898
rect 414804 200218 414986 200454
rect 415222 200218 415404 200454
rect 414804 200134 415404 200218
rect 414804 199898 414986 200134
rect 415222 199898 415404 200134
rect 414804 164454 415404 199898
rect 414804 164218 414986 164454
rect 415222 164218 415404 164454
rect 414804 164134 415404 164218
rect 414804 163898 414986 164134
rect 415222 163898 415404 164134
rect 414804 128454 415404 163898
rect 414804 128218 414986 128454
rect 415222 128218 415404 128454
rect 414804 128134 415404 128218
rect 414804 127898 414986 128134
rect 415222 127898 415404 128134
rect 414804 92454 415404 127898
rect 414804 92218 414986 92454
rect 415222 92218 415404 92454
rect 414804 92134 415404 92218
rect 414804 91898 414986 92134
rect 415222 91898 415404 92134
rect 414804 56454 415404 91898
rect 414804 56218 414986 56454
rect 415222 56218 415404 56454
rect 414804 56134 415404 56218
rect 414804 55898 414986 56134
rect 415222 55898 415404 56134
rect 414804 20454 415404 55898
rect 414804 20218 414986 20454
rect 415222 20218 415404 20454
rect 414804 20134 415404 20218
rect 414804 19898 414986 20134
rect 415222 19898 415404 20134
rect 414804 -1286 415404 19898
rect 414804 -1522 414986 -1286
rect 415222 -1522 415404 -1286
rect 414804 -1606 415404 -1522
rect 414804 -1842 414986 -1606
rect 415222 -1842 415404 -1606
rect 414804 -1864 415404 -1842
rect 418404 312054 419004 317000
rect 418404 311818 418586 312054
rect 418822 311818 419004 312054
rect 418404 311734 419004 311818
rect 418404 311498 418586 311734
rect 418822 311498 419004 311734
rect 418404 276054 419004 311498
rect 418404 275818 418586 276054
rect 418822 275818 419004 276054
rect 418404 275734 419004 275818
rect 418404 275498 418586 275734
rect 418822 275498 419004 275734
rect 418404 240054 419004 275498
rect 418404 239818 418586 240054
rect 418822 239818 419004 240054
rect 418404 239734 419004 239818
rect 418404 239498 418586 239734
rect 418822 239498 419004 239734
rect 418404 204054 419004 239498
rect 418404 203818 418586 204054
rect 418822 203818 419004 204054
rect 418404 203734 419004 203818
rect 418404 203498 418586 203734
rect 418822 203498 419004 203734
rect 418404 168054 419004 203498
rect 418404 167818 418586 168054
rect 418822 167818 419004 168054
rect 418404 167734 419004 167818
rect 418404 167498 418586 167734
rect 418822 167498 419004 167734
rect 418404 132054 419004 167498
rect 418404 131818 418586 132054
rect 418822 131818 419004 132054
rect 418404 131734 419004 131818
rect 418404 131498 418586 131734
rect 418822 131498 419004 131734
rect 418404 96054 419004 131498
rect 418404 95818 418586 96054
rect 418822 95818 419004 96054
rect 418404 95734 419004 95818
rect 418404 95498 418586 95734
rect 418822 95498 419004 95734
rect 418404 60054 419004 95498
rect 418404 59818 418586 60054
rect 418822 59818 419004 60054
rect 418404 59734 419004 59818
rect 418404 59498 418586 59734
rect 418822 59498 419004 59734
rect 418404 24054 419004 59498
rect 418404 23818 418586 24054
rect 418822 23818 419004 24054
rect 418404 23734 419004 23818
rect 418404 23498 418586 23734
rect 418822 23498 419004 23734
rect 418404 -3166 419004 23498
rect 418404 -3402 418586 -3166
rect 418822 -3402 419004 -3166
rect 418404 -3486 419004 -3402
rect 418404 -3722 418586 -3486
rect 418822 -3722 419004 -3486
rect 418404 -3744 419004 -3722
rect 422004 315654 422604 351098
rect 422004 315418 422186 315654
rect 422422 315418 422604 315654
rect 422004 315334 422604 315418
rect 422004 315098 422186 315334
rect 422422 315098 422604 315334
rect 422004 279654 422604 315098
rect 422004 279418 422186 279654
rect 422422 279418 422604 279654
rect 422004 279334 422604 279418
rect 422004 279098 422186 279334
rect 422422 279098 422604 279334
rect 422004 243654 422604 279098
rect 422004 243418 422186 243654
rect 422422 243418 422604 243654
rect 422004 243334 422604 243418
rect 422004 243098 422186 243334
rect 422422 243098 422604 243334
rect 422004 207654 422604 243098
rect 422004 207418 422186 207654
rect 422422 207418 422604 207654
rect 422004 207334 422604 207418
rect 422004 207098 422186 207334
rect 422422 207098 422604 207334
rect 422004 171654 422604 207098
rect 422004 171418 422186 171654
rect 422422 171418 422604 171654
rect 422004 171334 422604 171418
rect 422004 171098 422186 171334
rect 422422 171098 422604 171334
rect 422004 135654 422604 171098
rect 422004 135418 422186 135654
rect 422422 135418 422604 135654
rect 422004 135334 422604 135418
rect 422004 135098 422186 135334
rect 422422 135098 422604 135334
rect 422004 99654 422604 135098
rect 422004 99418 422186 99654
rect 422422 99418 422604 99654
rect 422004 99334 422604 99418
rect 422004 99098 422186 99334
rect 422422 99098 422604 99334
rect 422004 63654 422604 99098
rect 422004 63418 422186 63654
rect 422422 63418 422604 63654
rect 422004 63334 422604 63418
rect 422004 63098 422186 63334
rect 422422 63098 422604 63334
rect 422004 27654 422604 63098
rect 422004 27418 422186 27654
rect 422422 27418 422604 27654
rect 422004 27334 422604 27418
rect 422004 27098 422186 27334
rect 422422 27098 422604 27334
rect 422004 -5046 422604 27098
rect 422004 -5282 422186 -5046
rect 422422 -5282 422604 -5046
rect 422004 -5366 422604 -5282
rect 422004 -5602 422186 -5366
rect 422422 -5602 422604 -5366
rect 422004 -5624 422604 -5602
rect 425604 679254 426204 710862
rect 443604 710478 444204 711440
rect 443604 710242 443786 710478
rect 444022 710242 444204 710478
rect 443604 710158 444204 710242
rect 443604 709922 443786 710158
rect 444022 709922 444204 710158
rect 440004 708598 440604 709560
rect 440004 708362 440186 708598
rect 440422 708362 440604 708598
rect 440004 708278 440604 708362
rect 440004 708042 440186 708278
rect 440422 708042 440604 708278
rect 436404 706718 437004 707680
rect 436404 706482 436586 706718
rect 436822 706482 437004 706718
rect 436404 706398 437004 706482
rect 436404 706162 436586 706398
rect 436822 706162 437004 706398
rect 425604 679018 425786 679254
rect 426022 679018 426204 679254
rect 425604 678934 426204 679018
rect 425604 678698 425786 678934
rect 426022 678698 426204 678934
rect 425604 643254 426204 678698
rect 425604 643018 425786 643254
rect 426022 643018 426204 643254
rect 425604 642934 426204 643018
rect 425604 642698 425786 642934
rect 426022 642698 426204 642934
rect 425604 607254 426204 642698
rect 425604 607018 425786 607254
rect 426022 607018 426204 607254
rect 425604 606934 426204 607018
rect 425604 606698 425786 606934
rect 426022 606698 426204 606934
rect 425604 571254 426204 606698
rect 425604 571018 425786 571254
rect 426022 571018 426204 571254
rect 425604 570934 426204 571018
rect 425604 570698 425786 570934
rect 426022 570698 426204 570934
rect 425604 535254 426204 570698
rect 425604 535018 425786 535254
rect 426022 535018 426204 535254
rect 425604 534934 426204 535018
rect 425604 534698 425786 534934
rect 426022 534698 426204 534934
rect 425604 499254 426204 534698
rect 425604 499018 425786 499254
rect 426022 499018 426204 499254
rect 425604 498934 426204 499018
rect 425604 498698 425786 498934
rect 426022 498698 426204 498934
rect 425604 463254 426204 498698
rect 425604 463018 425786 463254
rect 426022 463018 426204 463254
rect 425604 462934 426204 463018
rect 425604 462698 425786 462934
rect 426022 462698 426204 462934
rect 425604 427254 426204 462698
rect 425604 427018 425786 427254
rect 426022 427018 426204 427254
rect 425604 426934 426204 427018
rect 425604 426698 425786 426934
rect 426022 426698 426204 426934
rect 425604 391254 426204 426698
rect 425604 391018 425786 391254
rect 426022 391018 426204 391254
rect 425604 390934 426204 391018
rect 425604 390698 425786 390934
rect 426022 390698 426204 390934
rect 425604 355254 426204 390698
rect 425604 355018 425786 355254
rect 426022 355018 426204 355254
rect 425604 354934 426204 355018
rect 425604 354698 425786 354934
rect 426022 354698 426204 354934
rect 425604 319254 426204 354698
rect 425604 319018 425786 319254
rect 426022 319018 426204 319254
rect 425604 318934 426204 319018
rect 425604 318698 425786 318934
rect 426022 318698 426204 318934
rect 425604 283254 426204 318698
rect 425604 283018 425786 283254
rect 426022 283018 426204 283254
rect 425604 282934 426204 283018
rect 425604 282698 425786 282934
rect 426022 282698 426204 282934
rect 425604 247254 426204 282698
rect 425604 247018 425786 247254
rect 426022 247018 426204 247254
rect 425604 246934 426204 247018
rect 425604 246698 425786 246934
rect 426022 246698 426204 246934
rect 425604 211254 426204 246698
rect 425604 211018 425786 211254
rect 426022 211018 426204 211254
rect 425604 210934 426204 211018
rect 425604 210698 425786 210934
rect 426022 210698 426204 210934
rect 425604 175254 426204 210698
rect 425604 175018 425786 175254
rect 426022 175018 426204 175254
rect 425604 174934 426204 175018
rect 425604 174698 425786 174934
rect 426022 174698 426204 174934
rect 425604 139254 426204 174698
rect 425604 139018 425786 139254
rect 426022 139018 426204 139254
rect 425604 138934 426204 139018
rect 425604 138698 425786 138934
rect 426022 138698 426204 138934
rect 425604 103254 426204 138698
rect 425604 103018 425786 103254
rect 426022 103018 426204 103254
rect 425604 102934 426204 103018
rect 425604 102698 425786 102934
rect 426022 102698 426204 102934
rect 425604 67254 426204 102698
rect 425604 67018 425786 67254
rect 426022 67018 426204 67254
rect 425604 66934 426204 67018
rect 425604 66698 425786 66934
rect 426022 66698 426204 66934
rect 425604 31254 426204 66698
rect 425604 31018 425786 31254
rect 426022 31018 426204 31254
rect 425604 30934 426204 31018
rect 425604 30698 425786 30934
rect 426022 30698 426204 30934
rect 407604 -6222 407786 -5986
rect 408022 -6222 408204 -5986
rect 407604 -6306 408204 -6222
rect 407604 -6542 407786 -6306
rect 408022 -6542 408204 -6306
rect 407604 -7504 408204 -6542
rect 425604 -6926 426204 30698
rect 432804 704838 433404 705800
rect 432804 704602 432986 704838
rect 433222 704602 433404 704838
rect 432804 704518 433404 704602
rect 432804 704282 432986 704518
rect 433222 704282 433404 704518
rect 432804 686454 433404 704282
rect 436404 690054 437004 706162
rect 436404 689818 436586 690054
rect 436822 689818 437004 690054
rect 436404 689734 437004 689818
rect 436404 689498 436586 689734
rect 436822 689498 437004 689734
rect 432804 686218 432986 686454
rect 433222 686218 433404 686454
rect 434667 686492 434733 686493
rect 434667 686428 434668 686492
rect 434732 686428 434733 686492
rect 434667 686427 434733 686428
rect 432804 686134 433404 686218
rect 432804 685898 432986 686134
rect 433222 685898 433404 686134
rect 434670 686085 434730 686427
rect 434667 686084 434733 686085
rect 434667 686020 434668 686084
rect 434732 686020 434733 686084
rect 434667 686019 434733 686020
rect 432804 650454 433404 685898
rect 436404 654054 437004 689498
rect 436404 653818 436586 654054
rect 436822 653818 437004 654054
rect 436404 653734 437004 653818
rect 436404 653498 436586 653734
rect 436822 653498 437004 653734
rect 434667 650860 434733 650861
rect 434667 650796 434668 650860
rect 434732 650796 434733 650860
rect 434667 650795 434733 650796
rect 432804 650218 432986 650454
rect 433222 650218 433404 650454
rect 434670 650453 434730 650795
rect 434667 650452 434733 650453
rect 434667 650388 434668 650452
rect 434732 650388 434733 650452
rect 434667 650387 434733 650388
rect 432804 650134 433404 650218
rect 432804 649898 432986 650134
rect 433222 649898 433404 650134
rect 432804 614454 433404 649898
rect 432804 614218 432986 614454
rect 433222 614218 433404 614454
rect 432804 614134 433404 614218
rect 432804 613898 432986 614134
rect 433222 613898 433404 614134
rect 432804 578454 433404 613898
rect 432804 578218 432986 578454
rect 433222 578218 433404 578454
rect 432804 578134 433404 578218
rect 432804 577898 432986 578134
rect 433222 577898 433404 578134
rect 432804 542454 433404 577898
rect 432804 542218 432986 542454
rect 433222 542218 433404 542454
rect 432804 542134 433404 542218
rect 432804 541898 432986 542134
rect 433222 541898 433404 542134
rect 432804 506454 433404 541898
rect 432804 506218 432986 506454
rect 433222 506218 433404 506454
rect 432804 506134 433404 506218
rect 432804 505898 432986 506134
rect 433222 505898 433404 506134
rect 432804 470454 433404 505898
rect 432804 470218 432986 470454
rect 433222 470218 433404 470454
rect 432804 470134 433404 470218
rect 432804 469898 432986 470134
rect 433222 469898 433404 470134
rect 432804 434454 433404 469898
rect 432804 434218 432986 434454
rect 433222 434218 433404 434454
rect 432804 434134 433404 434218
rect 432804 433898 432986 434134
rect 433222 433898 433404 434134
rect 432804 398454 433404 433898
rect 432804 398218 432986 398454
rect 433222 398218 433404 398454
rect 432804 398134 433404 398218
rect 432804 397898 432986 398134
rect 433222 397898 433404 398134
rect 432804 362454 433404 397898
rect 432804 362218 432986 362454
rect 433222 362218 433404 362454
rect 432804 362134 433404 362218
rect 432804 361898 432986 362134
rect 433222 361898 433404 362134
rect 432804 326454 433404 361898
rect 432804 326218 432986 326454
rect 433222 326218 433404 326454
rect 432804 326134 433404 326218
rect 432804 325898 432986 326134
rect 433222 325898 433404 326134
rect 432804 290454 433404 325898
rect 432804 290218 432986 290454
rect 433222 290218 433404 290454
rect 432804 290134 433404 290218
rect 432804 289898 432986 290134
rect 433222 289898 433404 290134
rect 432804 254454 433404 289898
rect 432804 254218 432986 254454
rect 433222 254218 433404 254454
rect 432804 254134 433404 254218
rect 432804 253898 432986 254134
rect 433222 253898 433404 254134
rect 432804 218454 433404 253898
rect 432804 218218 432986 218454
rect 433222 218218 433404 218454
rect 432804 218134 433404 218218
rect 432804 217898 432986 218134
rect 433222 217898 433404 218134
rect 432804 182454 433404 217898
rect 432804 182218 432986 182454
rect 433222 182218 433404 182454
rect 432804 182134 433404 182218
rect 432804 181898 432986 182134
rect 433222 181898 433404 182134
rect 432804 146454 433404 181898
rect 432804 146218 432986 146454
rect 433222 146218 433404 146454
rect 432804 146134 433404 146218
rect 432804 145898 432986 146134
rect 433222 145898 433404 146134
rect 432804 110454 433404 145898
rect 432804 110218 432986 110454
rect 433222 110218 433404 110454
rect 432804 110134 433404 110218
rect 432804 109898 432986 110134
rect 433222 109898 433404 110134
rect 432804 74454 433404 109898
rect 432804 74218 432986 74454
rect 433222 74218 433404 74454
rect 432804 74134 433404 74218
rect 432804 73898 432986 74134
rect 433222 73898 433404 74134
rect 432804 38454 433404 73898
rect 432804 38218 432986 38454
rect 433222 38218 433404 38454
rect 432804 38134 433404 38218
rect 432804 37898 432986 38134
rect 433222 37898 433404 38134
rect 432804 2454 433404 37898
rect 432804 2218 432986 2454
rect 433222 2218 433404 2454
rect 432804 2134 433404 2218
rect 432804 1898 432986 2134
rect 433222 1898 433404 2134
rect 432804 -346 433404 1898
rect 432804 -582 432986 -346
rect 433222 -582 433404 -346
rect 432804 -666 433404 -582
rect 432804 -902 432986 -666
rect 433222 -902 433404 -666
rect 432804 -1864 433404 -902
rect 436404 618054 437004 653498
rect 436404 617818 436586 618054
rect 436822 617818 437004 618054
rect 436404 617734 437004 617818
rect 436404 617498 436586 617734
rect 436822 617498 437004 617734
rect 436404 582054 437004 617498
rect 436404 581818 436586 582054
rect 436822 581818 437004 582054
rect 436404 581734 437004 581818
rect 436404 581498 436586 581734
rect 436822 581498 437004 581734
rect 436404 546054 437004 581498
rect 436404 545818 436586 546054
rect 436822 545818 437004 546054
rect 436404 545734 437004 545818
rect 436404 545498 436586 545734
rect 436822 545498 437004 545734
rect 436404 510054 437004 545498
rect 436404 509818 436586 510054
rect 436822 509818 437004 510054
rect 436404 509734 437004 509818
rect 436404 509498 436586 509734
rect 436822 509498 437004 509734
rect 436404 474054 437004 509498
rect 436404 473818 436586 474054
rect 436822 473818 437004 474054
rect 436404 473734 437004 473818
rect 436404 473498 436586 473734
rect 436822 473498 437004 473734
rect 436404 438054 437004 473498
rect 436404 437818 436586 438054
rect 436822 437818 437004 438054
rect 436404 437734 437004 437818
rect 436404 437498 436586 437734
rect 436822 437498 437004 437734
rect 436404 402054 437004 437498
rect 436404 401818 436586 402054
rect 436822 401818 437004 402054
rect 436404 401734 437004 401818
rect 436404 401498 436586 401734
rect 436822 401498 437004 401734
rect 436404 366054 437004 401498
rect 436404 365818 436586 366054
rect 436822 365818 437004 366054
rect 436404 365734 437004 365818
rect 436404 365498 436586 365734
rect 436822 365498 437004 365734
rect 436404 330054 437004 365498
rect 436404 329818 436586 330054
rect 436822 329818 437004 330054
rect 436404 329734 437004 329818
rect 436404 329498 436586 329734
rect 436822 329498 437004 329734
rect 436404 294054 437004 329498
rect 436404 293818 436586 294054
rect 436822 293818 437004 294054
rect 436404 293734 437004 293818
rect 436404 293498 436586 293734
rect 436822 293498 437004 293734
rect 436404 258054 437004 293498
rect 436404 257818 436586 258054
rect 436822 257818 437004 258054
rect 436404 257734 437004 257818
rect 436404 257498 436586 257734
rect 436822 257498 437004 257734
rect 436404 222054 437004 257498
rect 436404 221818 436586 222054
rect 436822 221818 437004 222054
rect 436404 221734 437004 221818
rect 436404 221498 436586 221734
rect 436822 221498 437004 221734
rect 436404 186054 437004 221498
rect 436404 185818 436586 186054
rect 436822 185818 437004 186054
rect 436404 185734 437004 185818
rect 436404 185498 436586 185734
rect 436822 185498 437004 185734
rect 436404 150054 437004 185498
rect 436404 149818 436586 150054
rect 436822 149818 437004 150054
rect 436404 149734 437004 149818
rect 436404 149498 436586 149734
rect 436822 149498 437004 149734
rect 436404 114054 437004 149498
rect 436404 113818 436586 114054
rect 436822 113818 437004 114054
rect 436404 113734 437004 113818
rect 436404 113498 436586 113734
rect 436822 113498 437004 113734
rect 436404 78054 437004 113498
rect 436404 77818 436586 78054
rect 436822 77818 437004 78054
rect 436404 77734 437004 77818
rect 436404 77498 436586 77734
rect 436822 77498 437004 77734
rect 436404 42054 437004 77498
rect 436404 41818 436586 42054
rect 436822 41818 437004 42054
rect 436404 41734 437004 41818
rect 436404 41498 436586 41734
rect 436822 41498 437004 41734
rect 436404 6054 437004 41498
rect 436404 5818 436586 6054
rect 436822 5818 437004 6054
rect 436404 5734 437004 5818
rect 436404 5498 436586 5734
rect 436822 5498 437004 5734
rect 436404 -2226 437004 5498
rect 436404 -2462 436586 -2226
rect 436822 -2462 437004 -2226
rect 436404 -2546 437004 -2462
rect 436404 -2782 436586 -2546
rect 436822 -2782 437004 -2546
rect 436404 -3744 437004 -2782
rect 440004 693654 440604 708042
rect 440004 693418 440186 693654
rect 440422 693418 440604 693654
rect 440004 693334 440604 693418
rect 440004 693098 440186 693334
rect 440422 693098 440604 693334
rect 440004 657654 440604 693098
rect 440004 657418 440186 657654
rect 440422 657418 440604 657654
rect 440004 657334 440604 657418
rect 440004 657098 440186 657334
rect 440422 657098 440604 657334
rect 440004 621654 440604 657098
rect 440004 621418 440186 621654
rect 440422 621418 440604 621654
rect 440004 621334 440604 621418
rect 440004 621098 440186 621334
rect 440422 621098 440604 621334
rect 440004 585654 440604 621098
rect 440004 585418 440186 585654
rect 440422 585418 440604 585654
rect 440004 585334 440604 585418
rect 440004 585098 440186 585334
rect 440422 585098 440604 585334
rect 440004 549654 440604 585098
rect 440004 549418 440186 549654
rect 440422 549418 440604 549654
rect 440004 549334 440604 549418
rect 440004 549098 440186 549334
rect 440422 549098 440604 549334
rect 440004 513654 440604 549098
rect 440004 513418 440186 513654
rect 440422 513418 440604 513654
rect 440004 513334 440604 513418
rect 440004 513098 440186 513334
rect 440422 513098 440604 513334
rect 440004 477654 440604 513098
rect 440004 477418 440186 477654
rect 440422 477418 440604 477654
rect 440004 477334 440604 477418
rect 440004 477098 440186 477334
rect 440422 477098 440604 477334
rect 440004 441654 440604 477098
rect 440004 441418 440186 441654
rect 440422 441418 440604 441654
rect 440004 441334 440604 441418
rect 440004 441098 440186 441334
rect 440422 441098 440604 441334
rect 440004 405654 440604 441098
rect 440004 405418 440186 405654
rect 440422 405418 440604 405654
rect 440004 405334 440604 405418
rect 440004 405098 440186 405334
rect 440422 405098 440604 405334
rect 440004 369654 440604 405098
rect 440004 369418 440186 369654
rect 440422 369418 440604 369654
rect 440004 369334 440604 369418
rect 440004 369098 440186 369334
rect 440422 369098 440604 369334
rect 440004 333654 440604 369098
rect 440004 333418 440186 333654
rect 440422 333418 440604 333654
rect 440004 333334 440604 333418
rect 440004 333098 440186 333334
rect 440422 333098 440604 333334
rect 440004 297654 440604 333098
rect 440004 297418 440186 297654
rect 440422 297418 440604 297654
rect 440004 297334 440604 297418
rect 440004 297098 440186 297334
rect 440422 297098 440604 297334
rect 440004 261654 440604 297098
rect 440004 261418 440186 261654
rect 440422 261418 440604 261654
rect 440004 261334 440604 261418
rect 440004 261098 440186 261334
rect 440422 261098 440604 261334
rect 440004 225654 440604 261098
rect 440004 225418 440186 225654
rect 440422 225418 440604 225654
rect 440004 225334 440604 225418
rect 440004 225098 440186 225334
rect 440422 225098 440604 225334
rect 440004 189654 440604 225098
rect 440004 189418 440186 189654
rect 440422 189418 440604 189654
rect 440004 189334 440604 189418
rect 440004 189098 440186 189334
rect 440422 189098 440604 189334
rect 440004 153654 440604 189098
rect 440004 153418 440186 153654
rect 440422 153418 440604 153654
rect 440004 153334 440604 153418
rect 440004 153098 440186 153334
rect 440422 153098 440604 153334
rect 440004 117654 440604 153098
rect 440004 117418 440186 117654
rect 440422 117418 440604 117654
rect 440004 117334 440604 117418
rect 440004 117098 440186 117334
rect 440422 117098 440604 117334
rect 440004 81654 440604 117098
rect 440004 81418 440186 81654
rect 440422 81418 440604 81654
rect 440004 81334 440604 81418
rect 440004 81098 440186 81334
rect 440422 81098 440604 81334
rect 440004 45654 440604 81098
rect 440004 45418 440186 45654
rect 440422 45418 440604 45654
rect 440004 45334 440604 45418
rect 440004 45098 440186 45334
rect 440422 45098 440604 45334
rect 440004 9654 440604 45098
rect 440004 9418 440186 9654
rect 440422 9418 440604 9654
rect 440004 9334 440604 9418
rect 440004 9098 440186 9334
rect 440422 9098 440604 9334
rect 440004 -4106 440604 9098
rect 440004 -4342 440186 -4106
rect 440422 -4342 440604 -4106
rect 440004 -4426 440604 -4342
rect 440004 -4662 440186 -4426
rect 440422 -4662 440604 -4426
rect 440004 -5624 440604 -4662
rect 443604 697254 444204 709922
rect 461604 711418 462204 711440
rect 461604 711182 461786 711418
rect 462022 711182 462204 711418
rect 461604 711098 462204 711182
rect 461604 710862 461786 711098
rect 462022 710862 462204 711098
rect 458004 709538 458604 709560
rect 458004 709302 458186 709538
rect 458422 709302 458604 709538
rect 458004 709218 458604 709302
rect 458004 708982 458186 709218
rect 458422 708982 458604 709218
rect 454404 707658 455004 707680
rect 454404 707422 454586 707658
rect 454822 707422 455004 707658
rect 454404 707338 455004 707422
rect 454404 707102 454586 707338
rect 454822 707102 455004 707338
rect 443604 697018 443786 697254
rect 444022 697018 444204 697254
rect 443604 696934 444204 697018
rect 443604 696698 443786 696934
rect 444022 696698 444204 696934
rect 443604 661254 444204 696698
rect 443604 661018 443786 661254
rect 444022 661018 444204 661254
rect 443604 660934 444204 661018
rect 443604 660698 443786 660934
rect 444022 660698 444204 660934
rect 443604 625254 444204 660698
rect 443604 625018 443786 625254
rect 444022 625018 444204 625254
rect 443604 624934 444204 625018
rect 443604 624698 443786 624934
rect 444022 624698 444204 624934
rect 443604 589254 444204 624698
rect 443604 589018 443786 589254
rect 444022 589018 444204 589254
rect 443604 588934 444204 589018
rect 443604 588698 443786 588934
rect 444022 588698 444204 588934
rect 443604 553254 444204 588698
rect 443604 553018 443786 553254
rect 444022 553018 444204 553254
rect 443604 552934 444204 553018
rect 443604 552698 443786 552934
rect 444022 552698 444204 552934
rect 443604 517254 444204 552698
rect 443604 517018 443786 517254
rect 444022 517018 444204 517254
rect 443604 516934 444204 517018
rect 443604 516698 443786 516934
rect 444022 516698 444204 516934
rect 443604 481254 444204 516698
rect 443604 481018 443786 481254
rect 444022 481018 444204 481254
rect 443604 480934 444204 481018
rect 443604 480698 443786 480934
rect 444022 480698 444204 480934
rect 443604 445254 444204 480698
rect 443604 445018 443786 445254
rect 444022 445018 444204 445254
rect 443604 444934 444204 445018
rect 443604 444698 443786 444934
rect 444022 444698 444204 444934
rect 443604 409254 444204 444698
rect 443604 409018 443786 409254
rect 444022 409018 444204 409254
rect 443604 408934 444204 409018
rect 443604 408698 443786 408934
rect 444022 408698 444204 408934
rect 443604 373254 444204 408698
rect 443604 373018 443786 373254
rect 444022 373018 444204 373254
rect 443604 372934 444204 373018
rect 443604 372698 443786 372934
rect 444022 372698 444204 372934
rect 443604 337254 444204 372698
rect 443604 337018 443786 337254
rect 444022 337018 444204 337254
rect 443604 336934 444204 337018
rect 443604 336698 443786 336934
rect 444022 336698 444204 336934
rect 443604 301254 444204 336698
rect 443604 301018 443786 301254
rect 444022 301018 444204 301254
rect 443604 300934 444204 301018
rect 443604 300698 443786 300934
rect 444022 300698 444204 300934
rect 443604 265254 444204 300698
rect 443604 265018 443786 265254
rect 444022 265018 444204 265254
rect 443604 264934 444204 265018
rect 443604 264698 443786 264934
rect 444022 264698 444204 264934
rect 443604 229254 444204 264698
rect 443604 229018 443786 229254
rect 444022 229018 444204 229254
rect 443604 228934 444204 229018
rect 443604 228698 443786 228934
rect 444022 228698 444204 228934
rect 443604 193254 444204 228698
rect 443604 193018 443786 193254
rect 444022 193018 444204 193254
rect 443604 192934 444204 193018
rect 443604 192698 443786 192934
rect 444022 192698 444204 192934
rect 443604 157254 444204 192698
rect 443604 157018 443786 157254
rect 444022 157018 444204 157254
rect 443604 156934 444204 157018
rect 443604 156698 443786 156934
rect 444022 156698 444204 156934
rect 443604 121254 444204 156698
rect 443604 121018 443786 121254
rect 444022 121018 444204 121254
rect 443604 120934 444204 121018
rect 443604 120698 443786 120934
rect 444022 120698 444204 120934
rect 443604 85254 444204 120698
rect 443604 85018 443786 85254
rect 444022 85018 444204 85254
rect 443604 84934 444204 85018
rect 443604 84698 443786 84934
rect 444022 84698 444204 84934
rect 443604 49254 444204 84698
rect 443604 49018 443786 49254
rect 444022 49018 444204 49254
rect 443604 48934 444204 49018
rect 443604 48698 443786 48934
rect 444022 48698 444204 48934
rect 443604 13254 444204 48698
rect 443604 13018 443786 13254
rect 444022 13018 444204 13254
rect 443604 12934 444204 13018
rect 443604 12698 443786 12934
rect 444022 12698 444204 12934
rect 425604 -7162 425786 -6926
rect 426022 -7162 426204 -6926
rect 425604 -7246 426204 -7162
rect 425604 -7482 425786 -7246
rect 426022 -7482 426204 -7246
rect 425604 -7504 426204 -7482
rect 443604 -5986 444204 12698
rect 450804 705778 451404 705800
rect 450804 705542 450986 705778
rect 451222 705542 451404 705778
rect 450804 705458 451404 705542
rect 450804 705222 450986 705458
rect 451222 705222 451404 705458
rect 450804 668454 451404 705222
rect 450804 668218 450986 668454
rect 451222 668218 451404 668454
rect 450804 668134 451404 668218
rect 450804 667898 450986 668134
rect 451222 667898 451404 668134
rect 450804 632454 451404 667898
rect 450804 632218 450986 632454
rect 451222 632218 451404 632454
rect 450804 632134 451404 632218
rect 450804 631898 450986 632134
rect 451222 631898 451404 632134
rect 450804 596454 451404 631898
rect 450804 596218 450986 596454
rect 451222 596218 451404 596454
rect 450804 596134 451404 596218
rect 450804 595898 450986 596134
rect 451222 595898 451404 596134
rect 450804 560454 451404 595898
rect 450804 560218 450986 560454
rect 451222 560218 451404 560454
rect 450804 560134 451404 560218
rect 450804 559898 450986 560134
rect 451222 559898 451404 560134
rect 450804 524454 451404 559898
rect 450804 524218 450986 524454
rect 451222 524218 451404 524454
rect 450804 524134 451404 524218
rect 450804 523898 450986 524134
rect 451222 523898 451404 524134
rect 450804 488454 451404 523898
rect 450804 488218 450986 488454
rect 451222 488218 451404 488454
rect 450804 488134 451404 488218
rect 450804 487898 450986 488134
rect 451222 487898 451404 488134
rect 450804 452454 451404 487898
rect 450804 452218 450986 452454
rect 451222 452218 451404 452454
rect 450804 452134 451404 452218
rect 450804 451898 450986 452134
rect 451222 451898 451404 452134
rect 450804 416454 451404 451898
rect 450804 416218 450986 416454
rect 451222 416218 451404 416454
rect 450804 416134 451404 416218
rect 450804 415898 450986 416134
rect 451222 415898 451404 416134
rect 450804 380454 451404 415898
rect 450804 380218 450986 380454
rect 451222 380218 451404 380454
rect 450804 380134 451404 380218
rect 450804 379898 450986 380134
rect 451222 379898 451404 380134
rect 450804 344454 451404 379898
rect 450804 344218 450986 344454
rect 451222 344218 451404 344454
rect 450804 344134 451404 344218
rect 450804 343898 450986 344134
rect 451222 343898 451404 344134
rect 450804 308454 451404 343898
rect 450804 308218 450986 308454
rect 451222 308218 451404 308454
rect 450804 308134 451404 308218
rect 450804 307898 450986 308134
rect 451222 307898 451404 308134
rect 450804 272454 451404 307898
rect 450804 272218 450986 272454
rect 451222 272218 451404 272454
rect 450804 272134 451404 272218
rect 450804 271898 450986 272134
rect 451222 271898 451404 272134
rect 450804 236454 451404 271898
rect 450804 236218 450986 236454
rect 451222 236218 451404 236454
rect 450804 236134 451404 236218
rect 450804 235898 450986 236134
rect 451222 235898 451404 236134
rect 450804 200454 451404 235898
rect 450804 200218 450986 200454
rect 451222 200218 451404 200454
rect 450804 200134 451404 200218
rect 450804 199898 450986 200134
rect 451222 199898 451404 200134
rect 450804 164454 451404 199898
rect 450804 164218 450986 164454
rect 451222 164218 451404 164454
rect 450804 164134 451404 164218
rect 450804 163898 450986 164134
rect 451222 163898 451404 164134
rect 450804 128454 451404 163898
rect 450804 128218 450986 128454
rect 451222 128218 451404 128454
rect 450804 128134 451404 128218
rect 450804 127898 450986 128134
rect 451222 127898 451404 128134
rect 450804 92454 451404 127898
rect 450804 92218 450986 92454
rect 451222 92218 451404 92454
rect 450804 92134 451404 92218
rect 450804 91898 450986 92134
rect 451222 91898 451404 92134
rect 450804 56454 451404 91898
rect 450804 56218 450986 56454
rect 451222 56218 451404 56454
rect 450804 56134 451404 56218
rect 450804 55898 450986 56134
rect 451222 55898 451404 56134
rect 450804 20454 451404 55898
rect 450804 20218 450986 20454
rect 451222 20218 451404 20454
rect 450804 20134 451404 20218
rect 450804 19898 450986 20134
rect 451222 19898 451404 20134
rect 450804 -1286 451404 19898
rect 450804 -1522 450986 -1286
rect 451222 -1522 451404 -1286
rect 450804 -1606 451404 -1522
rect 450804 -1842 450986 -1606
rect 451222 -1842 451404 -1606
rect 450804 -1864 451404 -1842
rect 454404 672054 455004 707102
rect 454404 671818 454586 672054
rect 454822 671818 455004 672054
rect 454404 671734 455004 671818
rect 454404 671498 454586 671734
rect 454822 671498 455004 671734
rect 454404 636054 455004 671498
rect 454404 635818 454586 636054
rect 454822 635818 455004 636054
rect 454404 635734 455004 635818
rect 454404 635498 454586 635734
rect 454822 635498 455004 635734
rect 454404 600054 455004 635498
rect 454404 599818 454586 600054
rect 454822 599818 455004 600054
rect 454404 599734 455004 599818
rect 454404 599498 454586 599734
rect 454822 599498 455004 599734
rect 454404 564054 455004 599498
rect 454404 563818 454586 564054
rect 454822 563818 455004 564054
rect 454404 563734 455004 563818
rect 454404 563498 454586 563734
rect 454822 563498 455004 563734
rect 454404 528054 455004 563498
rect 454404 527818 454586 528054
rect 454822 527818 455004 528054
rect 454404 527734 455004 527818
rect 454404 527498 454586 527734
rect 454822 527498 455004 527734
rect 454404 492054 455004 527498
rect 454404 491818 454586 492054
rect 454822 491818 455004 492054
rect 454404 491734 455004 491818
rect 454404 491498 454586 491734
rect 454822 491498 455004 491734
rect 454404 456054 455004 491498
rect 454404 455818 454586 456054
rect 454822 455818 455004 456054
rect 454404 455734 455004 455818
rect 454404 455498 454586 455734
rect 454822 455498 455004 455734
rect 454404 420054 455004 455498
rect 454404 419818 454586 420054
rect 454822 419818 455004 420054
rect 454404 419734 455004 419818
rect 454404 419498 454586 419734
rect 454822 419498 455004 419734
rect 454404 384054 455004 419498
rect 454404 383818 454586 384054
rect 454822 383818 455004 384054
rect 454404 383734 455004 383818
rect 454404 383498 454586 383734
rect 454822 383498 455004 383734
rect 454404 348054 455004 383498
rect 454404 347818 454586 348054
rect 454822 347818 455004 348054
rect 454404 347734 455004 347818
rect 454404 347498 454586 347734
rect 454822 347498 455004 347734
rect 454404 312054 455004 347498
rect 454404 311818 454586 312054
rect 454822 311818 455004 312054
rect 454404 311734 455004 311818
rect 454404 311498 454586 311734
rect 454822 311498 455004 311734
rect 454404 276054 455004 311498
rect 454404 275818 454586 276054
rect 454822 275818 455004 276054
rect 454404 275734 455004 275818
rect 454404 275498 454586 275734
rect 454822 275498 455004 275734
rect 454404 240054 455004 275498
rect 454404 239818 454586 240054
rect 454822 239818 455004 240054
rect 454404 239734 455004 239818
rect 454404 239498 454586 239734
rect 454822 239498 455004 239734
rect 454404 204054 455004 239498
rect 454404 203818 454586 204054
rect 454822 203818 455004 204054
rect 454404 203734 455004 203818
rect 454404 203498 454586 203734
rect 454822 203498 455004 203734
rect 454404 168054 455004 203498
rect 454404 167818 454586 168054
rect 454822 167818 455004 168054
rect 454404 167734 455004 167818
rect 454404 167498 454586 167734
rect 454822 167498 455004 167734
rect 454404 132054 455004 167498
rect 454404 131818 454586 132054
rect 454822 131818 455004 132054
rect 454404 131734 455004 131818
rect 454404 131498 454586 131734
rect 454822 131498 455004 131734
rect 454404 96054 455004 131498
rect 454404 95818 454586 96054
rect 454822 95818 455004 96054
rect 454404 95734 455004 95818
rect 454404 95498 454586 95734
rect 454822 95498 455004 95734
rect 454404 60054 455004 95498
rect 454404 59818 454586 60054
rect 454822 59818 455004 60054
rect 454404 59734 455004 59818
rect 454404 59498 454586 59734
rect 454822 59498 455004 59734
rect 454404 24054 455004 59498
rect 454404 23818 454586 24054
rect 454822 23818 455004 24054
rect 454404 23734 455004 23818
rect 454404 23498 454586 23734
rect 454822 23498 455004 23734
rect 454404 -3166 455004 23498
rect 454404 -3402 454586 -3166
rect 454822 -3402 455004 -3166
rect 454404 -3486 455004 -3402
rect 454404 -3722 454586 -3486
rect 454822 -3722 455004 -3486
rect 454404 -3744 455004 -3722
rect 458004 675654 458604 708982
rect 458004 675418 458186 675654
rect 458422 675418 458604 675654
rect 458004 675334 458604 675418
rect 458004 675098 458186 675334
rect 458422 675098 458604 675334
rect 458004 639654 458604 675098
rect 458004 639418 458186 639654
rect 458422 639418 458604 639654
rect 458004 639334 458604 639418
rect 458004 639098 458186 639334
rect 458422 639098 458604 639334
rect 458004 603654 458604 639098
rect 458004 603418 458186 603654
rect 458422 603418 458604 603654
rect 458004 603334 458604 603418
rect 458004 603098 458186 603334
rect 458422 603098 458604 603334
rect 458004 567654 458604 603098
rect 458004 567418 458186 567654
rect 458422 567418 458604 567654
rect 458004 567334 458604 567418
rect 458004 567098 458186 567334
rect 458422 567098 458604 567334
rect 458004 531654 458604 567098
rect 458004 531418 458186 531654
rect 458422 531418 458604 531654
rect 458004 531334 458604 531418
rect 458004 531098 458186 531334
rect 458422 531098 458604 531334
rect 458004 495654 458604 531098
rect 458004 495418 458186 495654
rect 458422 495418 458604 495654
rect 458004 495334 458604 495418
rect 458004 495098 458186 495334
rect 458422 495098 458604 495334
rect 458004 459654 458604 495098
rect 458004 459418 458186 459654
rect 458422 459418 458604 459654
rect 458004 459334 458604 459418
rect 458004 459098 458186 459334
rect 458422 459098 458604 459334
rect 458004 423654 458604 459098
rect 458004 423418 458186 423654
rect 458422 423418 458604 423654
rect 458004 423334 458604 423418
rect 458004 423098 458186 423334
rect 458422 423098 458604 423334
rect 458004 387654 458604 423098
rect 458004 387418 458186 387654
rect 458422 387418 458604 387654
rect 458004 387334 458604 387418
rect 458004 387098 458186 387334
rect 458422 387098 458604 387334
rect 458004 351654 458604 387098
rect 458004 351418 458186 351654
rect 458422 351418 458604 351654
rect 458004 351334 458604 351418
rect 458004 351098 458186 351334
rect 458422 351098 458604 351334
rect 458004 315654 458604 351098
rect 458004 315418 458186 315654
rect 458422 315418 458604 315654
rect 458004 315334 458604 315418
rect 458004 315098 458186 315334
rect 458422 315098 458604 315334
rect 458004 279654 458604 315098
rect 458004 279418 458186 279654
rect 458422 279418 458604 279654
rect 458004 279334 458604 279418
rect 458004 279098 458186 279334
rect 458422 279098 458604 279334
rect 458004 243654 458604 279098
rect 458004 243418 458186 243654
rect 458422 243418 458604 243654
rect 458004 243334 458604 243418
rect 458004 243098 458186 243334
rect 458422 243098 458604 243334
rect 458004 207654 458604 243098
rect 458004 207418 458186 207654
rect 458422 207418 458604 207654
rect 458004 207334 458604 207418
rect 458004 207098 458186 207334
rect 458422 207098 458604 207334
rect 458004 171654 458604 207098
rect 458004 171418 458186 171654
rect 458422 171418 458604 171654
rect 458004 171334 458604 171418
rect 458004 171098 458186 171334
rect 458422 171098 458604 171334
rect 458004 135654 458604 171098
rect 458004 135418 458186 135654
rect 458422 135418 458604 135654
rect 458004 135334 458604 135418
rect 458004 135098 458186 135334
rect 458422 135098 458604 135334
rect 458004 99654 458604 135098
rect 458004 99418 458186 99654
rect 458422 99418 458604 99654
rect 458004 99334 458604 99418
rect 458004 99098 458186 99334
rect 458422 99098 458604 99334
rect 458004 63654 458604 99098
rect 458004 63418 458186 63654
rect 458422 63418 458604 63654
rect 458004 63334 458604 63418
rect 458004 63098 458186 63334
rect 458422 63098 458604 63334
rect 458004 27654 458604 63098
rect 458004 27418 458186 27654
rect 458422 27418 458604 27654
rect 458004 27334 458604 27418
rect 458004 27098 458186 27334
rect 458422 27098 458604 27334
rect 458004 -5046 458604 27098
rect 458004 -5282 458186 -5046
rect 458422 -5282 458604 -5046
rect 458004 -5366 458604 -5282
rect 458004 -5602 458186 -5366
rect 458422 -5602 458604 -5366
rect 458004 -5624 458604 -5602
rect 461604 679254 462204 710862
rect 479604 710478 480204 711440
rect 479604 710242 479786 710478
rect 480022 710242 480204 710478
rect 479604 710158 480204 710242
rect 479604 709922 479786 710158
rect 480022 709922 480204 710158
rect 476004 708598 476604 709560
rect 476004 708362 476186 708598
rect 476422 708362 476604 708598
rect 476004 708278 476604 708362
rect 476004 708042 476186 708278
rect 476422 708042 476604 708278
rect 472404 706718 473004 707680
rect 472404 706482 472586 706718
rect 472822 706482 473004 706718
rect 472404 706398 473004 706482
rect 472404 706162 472586 706398
rect 472822 706162 473004 706398
rect 461604 679018 461786 679254
rect 462022 679018 462204 679254
rect 461604 678934 462204 679018
rect 461604 678698 461786 678934
rect 462022 678698 462204 678934
rect 461604 643254 462204 678698
rect 461604 643018 461786 643254
rect 462022 643018 462204 643254
rect 461604 642934 462204 643018
rect 461604 642698 461786 642934
rect 462022 642698 462204 642934
rect 461604 607254 462204 642698
rect 461604 607018 461786 607254
rect 462022 607018 462204 607254
rect 461604 606934 462204 607018
rect 461604 606698 461786 606934
rect 462022 606698 462204 606934
rect 461604 571254 462204 606698
rect 461604 571018 461786 571254
rect 462022 571018 462204 571254
rect 461604 570934 462204 571018
rect 461604 570698 461786 570934
rect 462022 570698 462204 570934
rect 461604 535254 462204 570698
rect 461604 535018 461786 535254
rect 462022 535018 462204 535254
rect 461604 534934 462204 535018
rect 461604 534698 461786 534934
rect 462022 534698 462204 534934
rect 461604 499254 462204 534698
rect 461604 499018 461786 499254
rect 462022 499018 462204 499254
rect 461604 498934 462204 499018
rect 461604 498698 461786 498934
rect 462022 498698 462204 498934
rect 461604 463254 462204 498698
rect 461604 463018 461786 463254
rect 462022 463018 462204 463254
rect 461604 462934 462204 463018
rect 461604 462698 461786 462934
rect 462022 462698 462204 462934
rect 461604 427254 462204 462698
rect 461604 427018 461786 427254
rect 462022 427018 462204 427254
rect 461604 426934 462204 427018
rect 461604 426698 461786 426934
rect 462022 426698 462204 426934
rect 461604 391254 462204 426698
rect 461604 391018 461786 391254
rect 462022 391018 462204 391254
rect 461604 390934 462204 391018
rect 461604 390698 461786 390934
rect 462022 390698 462204 390934
rect 461604 355254 462204 390698
rect 461604 355018 461786 355254
rect 462022 355018 462204 355254
rect 461604 354934 462204 355018
rect 461604 354698 461786 354934
rect 462022 354698 462204 354934
rect 461604 319254 462204 354698
rect 461604 319018 461786 319254
rect 462022 319018 462204 319254
rect 461604 318934 462204 319018
rect 461604 318698 461786 318934
rect 462022 318698 462204 318934
rect 461604 283254 462204 318698
rect 461604 283018 461786 283254
rect 462022 283018 462204 283254
rect 461604 282934 462204 283018
rect 461604 282698 461786 282934
rect 462022 282698 462204 282934
rect 461604 247254 462204 282698
rect 461604 247018 461786 247254
rect 462022 247018 462204 247254
rect 461604 246934 462204 247018
rect 461604 246698 461786 246934
rect 462022 246698 462204 246934
rect 461604 211254 462204 246698
rect 461604 211018 461786 211254
rect 462022 211018 462204 211254
rect 461604 210934 462204 211018
rect 461604 210698 461786 210934
rect 462022 210698 462204 210934
rect 461604 175254 462204 210698
rect 461604 175018 461786 175254
rect 462022 175018 462204 175254
rect 461604 174934 462204 175018
rect 461604 174698 461786 174934
rect 462022 174698 462204 174934
rect 461604 139254 462204 174698
rect 461604 139018 461786 139254
rect 462022 139018 462204 139254
rect 461604 138934 462204 139018
rect 461604 138698 461786 138934
rect 462022 138698 462204 138934
rect 461604 103254 462204 138698
rect 461604 103018 461786 103254
rect 462022 103018 462204 103254
rect 461604 102934 462204 103018
rect 461604 102698 461786 102934
rect 462022 102698 462204 102934
rect 461604 67254 462204 102698
rect 461604 67018 461786 67254
rect 462022 67018 462204 67254
rect 461604 66934 462204 67018
rect 461604 66698 461786 66934
rect 462022 66698 462204 66934
rect 461604 31254 462204 66698
rect 461604 31018 461786 31254
rect 462022 31018 462204 31254
rect 461604 30934 462204 31018
rect 461604 30698 461786 30934
rect 462022 30698 462204 30934
rect 443604 -6222 443786 -5986
rect 444022 -6222 444204 -5986
rect 443604 -6306 444204 -6222
rect 443604 -6542 443786 -6306
rect 444022 -6542 444204 -6306
rect 443604 -7504 444204 -6542
rect 461604 -6926 462204 30698
rect 468804 704838 469404 705800
rect 468804 704602 468986 704838
rect 469222 704602 469404 704838
rect 468804 704518 469404 704602
rect 468804 704282 468986 704518
rect 469222 704282 469404 704518
rect 468804 686454 469404 704282
rect 468804 686218 468986 686454
rect 469222 686218 469404 686454
rect 468804 686134 469404 686218
rect 468804 685898 468986 686134
rect 469222 685898 469404 686134
rect 468804 650454 469404 685898
rect 468804 650218 468986 650454
rect 469222 650218 469404 650454
rect 468804 650134 469404 650218
rect 468804 649898 468986 650134
rect 469222 649898 469404 650134
rect 468804 614454 469404 649898
rect 468804 614218 468986 614454
rect 469222 614218 469404 614454
rect 468804 614134 469404 614218
rect 468804 613898 468986 614134
rect 469222 613898 469404 614134
rect 468804 578454 469404 613898
rect 468804 578218 468986 578454
rect 469222 578218 469404 578454
rect 468804 578134 469404 578218
rect 468804 577898 468986 578134
rect 469222 577898 469404 578134
rect 468804 542454 469404 577898
rect 468804 542218 468986 542454
rect 469222 542218 469404 542454
rect 468804 542134 469404 542218
rect 468804 541898 468986 542134
rect 469222 541898 469404 542134
rect 468804 506454 469404 541898
rect 468804 506218 468986 506454
rect 469222 506218 469404 506454
rect 468804 506134 469404 506218
rect 468804 505898 468986 506134
rect 469222 505898 469404 506134
rect 468804 470454 469404 505898
rect 468804 470218 468986 470454
rect 469222 470218 469404 470454
rect 468804 470134 469404 470218
rect 468804 469898 468986 470134
rect 469222 469898 469404 470134
rect 468804 434454 469404 469898
rect 468804 434218 468986 434454
rect 469222 434218 469404 434454
rect 468804 434134 469404 434218
rect 468804 433898 468986 434134
rect 469222 433898 469404 434134
rect 468804 398454 469404 433898
rect 468804 398218 468986 398454
rect 469222 398218 469404 398454
rect 468804 398134 469404 398218
rect 468804 397898 468986 398134
rect 469222 397898 469404 398134
rect 468804 362454 469404 397898
rect 468804 362218 468986 362454
rect 469222 362218 469404 362454
rect 468804 362134 469404 362218
rect 468804 361898 468986 362134
rect 469222 361898 469404 362134
rect 468804 326454 469404 361898
rect 468804 326218 468986 326454
rect 469222 326218 469404 326454
rect 468804 326134 469404 326218
rect 468804 325898 468986 326134
rect 469222 325898 469404 326134
rect 468804 290454 469404 325898
rect 468804 290218 468986 290454
rect 469222 290218 469404 290454
rect 468804 290134 469404 290218
rect 468804 289898 468986 290134
rect 469222 289898 469404 290134
rect 468804 254454 469404 289898
rect 468804 254218 468986 254454
rect 469222 254218 469404 254454
rect 468804 254134 469404 254218
rect 468804 253898 468986 254134
rect 469222 253898 469404 254134
rect 468804 218454 469404 253898
rect 468804 218218 468986 218454
rect 469222 218218 469404 218454
rect 468804 218134 469404 218218
rect 468804 217898 468986 218134
rect 469222 217898 469404 218134
rect 468804 182454 469404 217898
rect 468804 182218 468986 182454
rect 469222 182218 469404 182454
rect 468804 182134 469404 182218
rect 468804 181898 468986 182134
rect 469222 181898 469404 182134
rect 468804 146454 469404 181898
rect 468804 146218 468986 146454
rect 469222 146218 469404 146454
rect 468804 146134 469404 146218
rect 468804 145898 468986 146134
rect 469222 145898 469404 146134
rect 468804 110454 469404 145898
rect 468804 110218 468986 110454
rect 469222 110218 469404 110454
rect 468804 110134 469404 110218
rect 468804 109898 468986 110134
rect 469222 109898 469404 110134
rect 468804 74454 469404 109898
rect 468804 74218 468986 74454
rect 469222 74218 469404 74454
rect 468804 74134 469404 74218
rect 468804 73898 468986 74134
rect 469222 73898 469404 74134
rect 468804 38454 469404 73898
rect 468804 38218 468986 38454
rect 469222 38218 469404 38454
rect 468804 38134 469404 38218
rect 468804 37898 468986 38134
rect 469222 37898 469404 38134
rect 468804 2454 469404 37898
rect 468804 2218 468986 2454
rect 469222 2218 469404 2454
rect 468804 2134 469404 2218
rect 468804 1898 468986 2134
rect 469222 1898 469404 2134
rect 468804 -346 469404 1898
rect 468804 -582 468986 -346
rect 469222 -582 469404 -346
rect 468804 -666 469404 -582
rect 468804 -902 468986 -666
rect 469222 -902 469404 -666
rect 468804 -1864 469404 -902
rect 472404 690054 473004 706162
rect 472404 689818 472586 690054
rect 472822 689818 473004 690054
rect 472404 689734 473004 689818
rect 472404 689498 472586 689734
rect 472822 689498 473004 689734
rect 472404 654054 473004 689498
rect 472404 653818 472586 654054
rect 472822 653818 473004 654054
rect 472404 653734 473004 653818
rect 472404 653498 472586 653734
rect 472822 653498 473004 653734
rect 472404 618054 473004 653498
rect 472404 617818 472586 618054
rect 472822 617818 473004 618054
rect 472404 617734 473004 617818
rect 472404 617498 472586 617734
rect 472822 617498 473004 617734
rect 472404 582054 473004 617498
rect 472404 581818 472586 582054
rect 472822 581818 473004 582054
rect 472404 581734 473004 581818
rect 472404 581498 472586 581734
rect 472822 581498 473004 581734
rect 472404 546054 473004 581498
rect 472404 545818 472586 546054
rect 472822 545818 473004 546054
rect 472404 545734 473004 545818
rect 472404 545498 472586 545734
rect 472822 545498 473004 545734
rect 472404 510054 473004 545498
rect 472404 509818 472586 510054
rect 472822 509818 473004 510054
rect 472404 509734 473004 509818
rect 472404 509498 472586 509734
rect 472822 509498 473004 509734
rect 472404 474054 473004 509498
rect 472404 473818 472586 474054
rect 472822 473818 473004 474054
rect 472404 473734 473004 473818
rect 472404 473498 472586 473734
rect 472822 473498 473004 473734
rect 472404 438054 473004 473498
rect 472404 437818 472586 438054
rect 472822 437818 473004 438054
rect 472404 437734 473004 437818
rect 472404 437498 472586 437734
rect 472822 437498 473004 437734
rect 472404 402054 473004 437498
rect 472404 401818 472586 402054
rect 472822 401818 473004 402054
rect 472404 401734 473004 401818
rect 472404 401498 472586 401734
rect 472822 401498 473004 401734
rect 472404 366054 473004 401498
rect 472404 365818 472586 366054
rect 472822 365818 473004 366054
rect 472404 365734 473004 365818
rect 472404 365498 472586 365734
rect 472822 365498 473004 365734
rect 472404 330054 473004 365498
rect 472404 329818 472586 330054
rect 472822 329818 473004 330054
rect 472404 329734 473004 329818
rect 472404 329498 472586 329734
rect 472822 329498 473004 329734
rect 472404 294054 473004 329498
rect 472404 293818 472586 294054
rect 472822 293818 473004 294054
rect 472404 293734 473004 293818
rect 472404 293498 472586 293734
rect 472822 293498 473004 293734
rect 472404 258054 473004 293498
rect 472404 257818 472586 258054
rect 472822 257818 473004 258054
rect 472404 257734 473004 257818
rect 472404 257498 472586 257734
rect 472822 257498 473004 257734
rect 472404 222054 473004 257498
rect 472404 221818 472586 222054
rect 472822 221818 473004 222054
rect 472404 221734 473004 221818
rect 472404 221498 472586 221734
rect 472822 221498 473004 221734
rect 472404 186054 473004 221498
rect 472404 185818 472586 186054
rect 472822 185818 473004 186054
rect 472404 185734 473004 185818
rect 472404 185498 472586 185734
rect 472822 185498 473004 185734
rect 472404 150054 473004 185498
rect 472404 149818 472586 150054
rect 472822 149818 473004 150054
rect 472404 149734 473004 149818
rect 472404 149498 472586 149734
rect 472822 149498 473004 149734
rect 472404 114054 473004 149498
rect 472404 113818 472586 114054
rect 472822 113818 473004 114054
rect 472404 113734 473004 113818
rect 472404 113498 472586 113734
rect 472822 113498 473004 113734
rect 472404 78054 473004 113498
rect 472404 77818 472586 78054
rect 472822 77818 473004 78054
rect 472404 77734 473004 77818
rect 472404 77498 472586 77734
rect 472822 77498 473004 77734
rect 472404 42054 473004 77498
rect 472404 41818 472586 42054
rect 472822 41818 473004 42054
rect 472404 41734 473004 41818
rect 472404 41498 472586 41734
rect 472822 41498 473004 41734
rect 472404 6054 473004 41498
rect 472404 5818 472586 6054
rect 472822 5818 473004 6054
rect 472404 5734 473004 5818
rect 472404 5498 472586 5734
rect 472822 5498 473004 5734
rect 472404 -2226 473004 5498
rect 472404 -2462 472586 -2226
rect 472822 -2462 473004 -2226
rect 472404 -2546 473004 -2462
rect 472404 -2782 472586 -2546
rect 472822 -2782 473004 -2546
rect 472404 -3744 473004 -2782
rect 476004 693654 476604 708042
rect 476004 693418 476186 693654
rect 476422 693418 476604 693654
rect 476004 693334 476604 693418
rect 476004 693098 476186 693334
rect 476422 693098 476604 693334
rect 476004 657654 476604 693098
rect 476004 657418 476186 657654
rect 476422 657418 476604 657654
rect 476004 657334 476604 657418
rect 476004 657098 476186 657334
rect 476422 657098 476604 657334
rect 476004 621654 476604 657098
rect 476004 621418 476186 621654
rect 476422 621418 476604 621654
rect 476004 621334 476604 621418
rect 476004 621098 476186 621334
rect 476422 621098 476604 621334
rect 476004 585654 476604 621098
rect 476004 585418 476186 585654
rect 476422 585418 476604 585654
rect 476004 585334 476604 585418
rect 476004 585098 476186 585334
rect 476422 585098 476604 585334
rect 476004 549654 476604 585098
rect 476004 549418 476186 549654
rect 476422 549418 476604 549654
rect 476004 549334 476604 549418
rect 476004 549098 476186 549334
rect 476422 549098 476604 549334
rect 476004 513654 476604 549098
rect 476004 513418 476186 513654
rect 476422 513418 476604 513654
rect 476004 513334 476604 513418
rect 476004 513098 476186 513334
rect 476422 513098 476604 513334
rect 476004 477654 476604 513098
rect 476004 477418 476186 477654
rect 476422 477418 476604 477654
rect 476004 477334 476604 477418
rect 476004 477098 476186 477334
rect 476422 477098 476604 477334
rect 476004 441654 476604 477098
rect 476004 441418 476186 441654
rect 476422 441418 476604 441654
rect 476004 441334 476604 441418
rect 476004 441098 476186 441334
rect 476422 441098 476604 441334
rect 476004 405654 476604 441098
rect 476004 405418 476186 405654
rect 476422 405418 476604 405654
rect 476004 405334 476604 405418
rect 476004 405098 476186 405334
rect 476422 405098 476604 405334
rect 476004 369654 476604 405098
rect 476004 369418 476186 369654
rect 476422 369418 476604 369654
rect 476004 369334 476604 369418
rect 476004 369098 476186 369334
rect 476422 369098 476604 369334
rect 476004 333654 476604 369098
rect 476004 333418 476186 333654
rect 476422 333418 476604 333654
rect 476004 333334 476604 333418
rect 476004 333098 476186 333334
rect 476422 333098 476604 333334
rect 476004 297654 476604 333098
rect 476004 297418 476186 297654
rect 476422 297418 476604 297654
rect 476004 297334 476604 297418
rect 476004 297098 476186 297334
rect 476422 297098 476604 297334
rect 476004 261654 476604 297098
rect 476004 261418 476186 261654
rect 476422 261418 476604 261654
rect 476004 261334 476604 261418
rect 476004 261098 476186 261334
rect 476422 261098 476604 261334
rect 476004 225654 476604 261098
rect 476004 225418 476186 225654
rect 476422 225418 476604 225654
rect 476004 225334 476604 225418
rect 476004 225098 476186 225334
rect 476422 225098 476604 225334
rect 476004 189654 476604 225098
rect 476004 189418 476186 189654
rect 476422 189418 476604 189654
rect 476004 189334 476604 189418
rect 476004 189098 476186 189334
rect 476422 189098 476604 189334
rect 476004 153654 476604 189098
rect 476004 153418 476186 153654
rect 476422 153418 476604 153654
rect 476004 153334 476604 153418
rect 476004 153098 476186 153334
rect 476422 153098 476604 153334
rect 476004 117654 476604 153098
rect 476004 117418 476186 117654
rect 476422 117418 476604 117654
rect 476004 117334 476604 117418
rect 476004 117098 476186 117334
rect 476422 117098 476604 117334
rect 476004 81654 476604 117098
rect 476004 81418 476186 81654
rect 476422 81418 476604 81654
rect 476004 81334 476604 81418
rect 476004 81098 476186 81334
rect 476422 81098 476604 81334
rect 476004 45654 476604 81098
rect 476004 45418 476186 45654
rect 476422 45418 476604 45654
rect 476004 45334 476604 45418
rect 476004 45098 476186 45334
rect 476422 45098 476604 45334
rect 476004 9654 476604 45098
rect 476004 9418 476186 9654
rect 476422 9418 476604 9654
rect 476004 9334 476604 9418
rect 476004 9098 476186 9334
rect 476422 9098 476604 9334
rect 476004 -4106 476604 9098
rect 476004 -4342 476186 -4106
rect 476422 -4342 476604 -4106
rect 476004 -4426 476604 -4342
rect 476004 -4662 476186 -4426
rect 476422 -4662 476604 -4426
rect 476004 -5624 476604 -4662
rect 479604 697254 480204 709922
rect 497604 711418 498204 711440
rect 497604 711182 497786 711418
rect 498022 711182 498204 711418
rect 497604 711098 498204 711182
rect 497604 710862 497786 711098
rect 498022 710862 498204 711098
rect 494004 709538 494604 709560
rect 494004 709302 494186 709538
rect 494422 709302 494604 709538
rect 494004 709218 494604 709302
rect 494004 708982 494186 709218
rect 494422 708982 494604 709218
rect 490404 707658 491004 707680
rect 490404 707422 490586 707658
rect 490822 707422 491004 707658
rect 490404 707338 491004 707422
rect 490404 707102 490586 707338
rect 490822 707102 491004 707338
rect 479604 697018 479786 697254
rect 480022 697018 480204 697254
rect 479604 696934 480204 697018
rect 479604 696698 479786 696934
rect 480022 696698 480204 696934
rect 479604 661254 480204 696698
rect 479604 661018 479786 661254
rect 480022 661018 480204 661254
rect 479604 660934 480204 661018
rect 479604 660698 479786 660934
rect 480022 660698 480204 660934
rect 479604 625254 480204 660698
rect 479604 625018 479786 625254
rect 480022 625018 480204 625254
rect 479604 624934 480204 625018
rect 479604 624698 479786 624934
rect 480022 624698 480204 624934
rect 479604 589254 480204 624698
rect 479604 589018 479786 589254
rect 480022 589018 480204 589254
rect 479604 588934 480204 589018
rect 479604 588698 479786 588934
rect 480022 588698 480204 588934
rect 479604 553254 480204 588698
rect 479604 553018 479786 553254
rect 480022 553018 480204 553254
rect 479604 552934 480204 553018
rect 479604 552698 479786 552934
rect 480022 552698 480204 552934
rect 479604 517254 480204 552698
rect 479604 517018 479786 517254
rect 480022 517018 480204 517254
rect 479604 516934 480204 517018
rect 479604 516698 479786 516934
rect 480022 516698 480204 516934
rect 479604 481254 480204 516698
rect 479604 481018 479786 481254
rect 480022 481018 480204 481254
rect 479604 480934 480204 481018
rect 479604 480698 479786 480934
rect 480022 480698 480204 480934
rect 479604 445254 480204 480698
rect 479604 445018 479786 445254
rect 480022 445018 480204 445254
rect 479604 444934 480204 445018
rect 479604 444698 479786 444934
rect 480022 444698 480204 444934
rect 479604 409254 480204 444698
rect 479604 409018 479786 409254
rect 480022 409018 480204 409254
rect 479604 408934 480204 409018
rect 479604 408698 479786 408934
rect 480022 408698 480204 408934
rect 479604 373254 480204 408698
rect 479604 373018 479786 373254
rect 480022 373018 480204 373254
rect 479604 372934 480204 373018
rect 479604 372698 479786 372934
rect 480022 372698 480204 372934
rect 479604 337254 480204 372698
rect 479604 337018 479786 337254
rect 480022 337018 480204 337254
rect 479604 336934 480204 337018
rect 479604 336698 479786 336934
rect 480022 336698 480204 336934
rect 479604 301254 480204 336698
rect 479604 301018 479786 301254
rect 480022 301018 480204 301254
rect 479604 300934 480204 301018
rect 479604 300698 479786 300934
rect 480022 300698 480204 300934
rect 479604 265254 480204 300698
rect 479604 265018 479786 265254
rect 480022 265018 480204 265254
rect 479604 264934 480204 265018
rect 479604 264698 479786 264934
rect 480022 264698 480204 264934
rect 479604 229254 480204 264698
rect 479604 229018 479786 229254
rect 480022 229018 480204 229254
rect 479604 228934 480204 229018
rect 479604 228698 479786 228934
rect 480022 228698 480204 228934
rect 479604 193254 480204 228698
rect 479604 193018 479786 193254
rect 480022 193018 480204 193254
rect 479604 192934 480204 193018
rect 479604 192698 479786 192934
rect 480022 192698 480204 192934
rect 479604 157254 480204 192698
rect 479604 157018 479786 157254
rect 480022 157018 480204 157254
rect 479604 156934 480204 157018
rect 479604 156698 479786 156934
rect 480022 156698 480204 156934
rect 479604 121254 480204 156698
rect 479604 121018 479786 121254
rect 480022 121018 480204 121254
rect 479604 120934 480204 121018
rect 479604 120698 479786 120934
rect 480022 120698 480204 120934
rect 479604 85254 480204 120698
rect 479604 85018 479786 85254
rect 480022 85018 480204 85254
rect 479604 84934 480204 85018
rect 479604 84698 479786 84934
rect 480022 84698 480204 84934
rect 479604 49254 480204 84698
rect 479604 49018 479786 49254
rect 480022 49018 480204 49254
rect 479604 48934 480204 49018
rect 479604 48698 479786 48934
rect 480022 48698 480204 48934
rect 479604 13254 480204 48698
rect 479604 13018 479786 13254
rect 480022 13018 480204 13254
rect 479604 12934 480204 13018
rect 479604 12698 479786 12934
rect 480022 12698 480204 12934
rect 461604 -7162 461786 -6926
rect 462022 -7162 462204 -6926
rect 461604 -7246 462204 -7162
rect 461604 -7482 461786 -7246
rect 462022 -7482 462204 -7246
rect 461604 -7504 462204 -7482
rect 479604 -5986 480204 12698
rect 486804 705778 487404 705800
rect 486804 705542 486986 705778
rect 487222 705542 487404 705778
rect 486804 705458 487404 705542
rect 486804 705222 486986 705458
rect 487222 705222 487404 705458
rect 486804 668454 487404 705222
rect 486804 668218 486986 668454
rect 487222 668218 487404 668454
rect 486804 668134 487404 668218
rect 486804 667898 486986 668134
rect 487222 667898 487404 668134
rect 486804 632454 487404 667898
rect 486804 632218 486986 632454
rect 487222 632218 487404 632454
rect 486804 632134 487404 632218
rect 486804 631898 486986 632134
rect 487222 631898 487404 632134
rect 486804 596454 487404 631898
rect 486804 596218 486986 596454
rect 487222 596218 487404 596454
rect 486804 596134 487404 596218
rect 486804 595898 486986 596134
rect 487222 595898 487404 596134
rect 486804 560454 487404 595898
rect 486804 560218 486986 560454
rect 487222 560218 487404 560454
rect 486804 560134 487404 560218
rect 486804 559898 486986 560134
rect 487222 559898 487404 560134
rect 486804 524454 487404 559898
rect 486804 524218 486986 524454
rect 487222 524218 487404 524454
rect 486804 524134 487404 524218
rect 486804 523898 486986 524134
rect 487222 523898 487404 524134
rect 486804 488454 487404 523898
rect 486804 488218 486986 488454
rect 487222 488218 487404 488454
rect 486804 488134 487404 488218
rect 486804 487898 486986 488134
rect 487222 487898 487404 488134
rect 486804 452454 487404 487898
rect 486804 452218 486986 452454
rect 487222 452218 487404 452454
rect 486804 452134 487404 452218
rect 486804 451898 486986 452134
rect 487222 451898 487404 452134
rect 486804 416454 487404 451898
rect 486804 416218 486986 416454
rect 487222 416218 487404 416454
rect 486804 416134 487404 416218
rect 486804 415898 486986 416134
rect 487222 415898 487404 416134
rect 486804 380454 487404 415898
rect 486804 380218 486986 380454
rect 487222 380218 487404 380454
rect 486804 380134 487404 380218
rect 486804 379898 486986 380134
rect 487222 379898 487404 380134
rect 486804 344454 487404 379898
rect 486804 344218 486986 344454
rect 487222 344218 487404 344454
rect 486804 344134 487404 344218
rect 486804 343898 486986 344134
rect 487222 343898 487404 344134
rect 486804 308454 487404 343898
rect 486804 308218 486986 308454
rect 487222 308218 487404 308454
rect 486804 308134 487404 308218
rect 486804 307898 486986 308134
rect 487222 307898 487404 308134
rect 486804 272454 487404 307898
rect 486804 272218 486986 272454
rect 487222 272218 487404 272454
rect 486804 272134 487404 272218
rect 486804 271898 486986 272134
rect 487222 271898 487404 272134
rect 486804 236454 487404 271898
rect 486804 236218 486986 236454
rect 487222 236218 487404 236454
rect 486804 236134 487404 236218
rect 486804 235898 486986 236134
rect 487222 235898 487404 236134
rect 486804 200454 487404 235898
rect 486804 200218 486986 200454
rect 487222 200218 487404 200454
rect 486804 200134 487404 200218
rect 486804 199898 486986 200134
rect 487222 199898 487404 200134
rect 486804 164454 487404 199898
rect 486804 164218 486986 164454
rect 487222 164218 487404 164454
rect 486804 164134 487404 164218
rect 486804 163898 486986 164134
rect 487222 163898 487404 164134
rect 486804 128454 487404 163898
rect 486804 128218 486986 128454
rect 487222 128218 487404 128454
rect 486804 128134 487404 128218
rect 486804 127898 486986 128134
rect 487222 127898 487404 128134
rect 486804 92454 487404 127898
rect 486804 92218 486986 92454
rect 487222 92218 487404 92454
rect 486804 92134 487404 92218
rect 486804 91898 486986 92134
rect 487222 91898 487404 92134
rect 486804 56454 487404 91898
rect 486804 56218 486986 56454
rect 487222 56218 487404 56454
rect 486804 56134 487404 56218
rect 486804 55898 486986 56134
rect 487222 55898 487404 56134
rect 486804 20454 487404 55898
rect 486804 20218 486986 20454
rect 487222 20218 487404 20454
rect 486804 20134 487404 20218
rect 486804 19898 486986 20134
rect 487222 19898 487404 20134
rect 486804 -1286 487404 19898
rect 486804 -1522 486986 -1286
rect 487222 -1522 487404 -1286
rect 486804 -1606 487404 -1522
rect 486804 -1842 486986 -1606
rect 487222 -1842 487404 -1606
rect 486804 -1864 487404 -1842
rect 490404 672054 491004 707102
rect 490404 671818 490586 672054
rect 490822 671818 491004 672054
rect 490404 671734 491004 671818
rect 490404 671498 490586 671734
rect 490822 671498 491004 671734
rect 490404 636054 491004 671498
rect 490404 635818 490586 636054
rect 490822 635818 491004 636054
rect 490404 635734 491004 635818
rect 490404 635498 490586 635734
rect 490822 635498 491004 635734
rect 490404 600054 491004 635498
rect 490404 599818 490586 600054
rect 490822 599818 491004 600054
rect 490404 599734 491004 599818
rect 490404 599498 490586 599734
rect 490822 599498 491004 599734
rect 490404 564054 491004 599498
rect 490404 563818 490586 564054
rect 490822 563818 491004 564054
rect 490404 563734 491004 563818
rect 490404 563498 490586 563734
rect 490822 563498 491004 563734
rect 490404 528054 491004 563498
rect 494004 675654 494604 708982
rect 494004 675418 494186 675654
rect 494422 675418 494604 675654
rect 494004 675334 494604 675418
rect 494004 675098 494186 675334
rect 494422 675098 494604 675334
rect 494004 639654 494604 675098
rect 494004 639418 494186 639654
rect 494422 639418 494604 639654
rect 494004 639334 494604 639418
rect 494004 639098 494186 639334
rect 494422 639098 494604 639334
rect 494004 603654 494604 639098
rect 494004 603418 494186 603654
rect 494422 603418 494604 603654
rect 494004 603334 494604 603418
rect 494004 603098 494186 603334
rect 494422 603098 494604 603334
rect 494004 567654 494604 603098
rect 494004 567418 494186 567654
rect 494422 567418 494604 567654
rect 494004 567334 494604 567418
rect 494004 567098 494186 567334
rect 494422 567098 494604 567334
rect 492627 545460 492693 545461
rect 492627 545396 492628 545460
rect 492692 545396 492693 545460
rect 492627 545395 492693 545396
rect 492630 545189 492690 545395
rect 492627 545188 492693 545189
rect 492627 545124 492628 545188
rect 492692 545124 492693 545188
rect 492627 545123 492693 545124
rect 490404 527818 490586 528054
rect 490822 527818 491004 528054
rect 490404 527734 491004 527818
rect 490404 527498 490586 527734
rect 490822 527498 491004 527734
rect 490404 492054 491004 527498
rect 490404 491818 490586 492054
rect 490822 491818 491004 492054
rect 490404 491734 491004 491818
rect 490404 491498 490586 491734
rect 490822 491498 491004 491734
rect 490404 456054 491004 491498
rect 490404 455818 490586 456054
rect 490822 455818 491004 456054
rect 490404 455734 491004 455818
rect 490404 455498 490586 455734
rect 490822 455498 491004 455734
rect 490404 420054 491004 455498
rect 490404 419818 490586 420054
rect 490822 419818 491004 420054
rect 490404 419734 491004 419818
rect 490404 419498 490586 419734
rect 490822 419498 491004 419734
rect 490404 384054 491004 419498
rect 490404 383818 490586 384054
rect 490822 383818 491004 384054
rect 490404 383734 491004 383818
rect 490404 383498 490586 383734
rect 490822 383498 491004 383734
rect 490404 348054 491004 383498
rect 490404 347818 490586 348054
rect 490822 347818 491004 348054
rect 490404 347734 491004 347818
rect 490404 347498 490586 347734
rect 490822 347498 491004 347734
rect 490404 312054 491004 347498
rect 490404 311818 490586 312054
rect 490822 311818 491004 312054
rect 490404 311734 491004 311818
rect 490404 311498 490586 311734
rect 490822 311498 491004 311734
rect 490404 276054 491004 311498
rect 490404 275818 490586 276054
rect 490822 275818 491004 276054
rect 490404 275734 491004 275818
rect 490404 275498 490586 275734
rect 490822 275498 491004 275734
rect 490404 240054 491004 275498
rect 490404 239818 490586 240054
rect 490822 239818 491004 240054
rect 490404 239734 491004 239818
rect 490404 239498 490586 239734
rect 490822 239498 491004 239734
rect 490404 204054 491004 239498
rect 490404 203818 490586 204054
rect 490822 203818 491004 204054
rect 490404 203734 491004 203818
rect 490404 203498 490586 203734
rect 490822 203498 491004 203734
rect 490404 168054 491004 203498
rect 490404 167818 490586 168054
rect 490822 167818 491004 168054
rect 490404 167734 491004 167818
rect 490404 167498 490586 167734
rect 490822 167498 491004 167734
rect 490404 132054 491004 167498
rect 490404 131818 490586 132054
rect 490822 131818 491004 132054
rect 490404 131734 491004 131818
rect 490404 131498 490586 131734
rect 490822 131498 491004 131734
rect 490404 96054 491004 131498
rect 490404 95818 490586 96054
rect 490822 95818 491004 96054
rect 490404 95734 491004 95818
rect 490404 95498 490586 95734
rect 490822 95498 491004 95734
rect 490404 60054 491004 95498
rect 490404 59818 490586 60054
rect 490822 59818 491004 60054
rect 490404 59734 491004 59818
rect 490404 59498 490586 59734
rect 490822 59498 491004 59734
rect 490404 24054 491004 59498
rect 490404 23818 490586 24054
rect 490822 23818 491004 24054
rect 490404 23734 491004 23818
rect 490404 23498 490586 23734
rect 490822 23498 491004 23734
rect 490404 -3166 491004 23498
rect 490404 -3402 490586 -3166
rect 490822 -3402 491004 -3166
rect 490404 -3486 491004 -3402
rect 490404 -3722 490586 -3486
rect 490822 -3722 491004 -3486
rect 490404 -3744 491004 -3722
rect 494004 531654 494604 567098
rect 494004 531418 494186 531654
rect 494422 531418 494604 531654
rect 494004 531334 494604 531418
rect 494004 531098 494186 531334
rect 494422 531098 494604 531334
rect 494004 495654 494604 531098
rect 494004 495418 494186 495654
rect 494422 495418 494604 495654
rect 494004 495334 494604 495418
rect 494004 495098 494186 495334
rect 494422 495098 494604 495334
rect 494004 459654 494604 495098
rect 494004 459418 494186 459654
rect 494422 459418 494604 459654
rect 494004 459334 494604 459418
rect 494004 459098 494186 459334
rect 494422 459098 494604 459334
rect 494004 423654 494604 459098
rect 494004 423418 494186 423654
rect 494422 423418 494604 423654
rect 494004 423334 494604 423418
rect 494004 423098 494186 423334
rect 494422 423098 494604 423334
rect 494004 387654 494604 423098
rect 494004 387418 494186 387654
rect 494422 387418 494604 387654
rect 494004 387334 494604 387418
rect 494004 387098 494186 387334
rect 494422 387098 494604 387334
rect 494004 351654 494604 387098
rect 494004 351418 494186 351654
rect 494422 351418 494604 351654
rect 494004 351334 494604 351418
rect 494004 351098 494186 351334
rect 494422 351098 494604 351334
rect 494004 315654 494604 351098
rect 494004 315418 494186 315654
rect 494422 315418 494604 315654
rect 494004 315334 494604 315418
rect 494004 315098 494186 315334
rect 494422 315098 494604 315334
rect 494004 279654 494604 315098
rect 494004 279418 494186 279654
rect 494422 279418 494604 279654
rect 494004 279334 494604 279418
rect 494004 279098 494186 279334
rect 494422 279098 494604 279334
rect 494004 243654 494604 279098
rect 494004 243418 494186 243654
rect 494422 243418 494604 243654
rect 494004 243334 494604 243418
rect 494004 243098 494186 243334
rect 494422 243098 494604 243334
rect 494004 207654 494604 243098
rect 494004 207418 494186 207654
rect 494422 207418 494604 207654
rect 494004 207334 494604 207418
rect 494004 207098 494186 207334
rect 494422 207098 494604 207334
rect 494004 171654 494604 207098
rect 494004 171418 494186 171654
rect 494422 171418 494604 171654
rect 494004 171334 494604 171418
rect 494004 171098 494186 171334
rect 494422 171098 494604 171334
rect 494004 135654 494604 171098
rect 494004 135418 494186 135654
rect 494422 135418 494604 135654
rect 494004 135334 494604 135418
rect 494004 135098 494186 135334
rect 494422 135098 494604 135334
rect 494004 99654 494604 135098
rect 494004 99418 494186 99654
rect 494422 99418 494604 99654
rect 494004 99334 494604 99418
rect 494004 99098 494186 99334
rect 494422 99098 494604 99334
rect 494004 63654 494604 99098
rect 494004 63418 494186 63654
rect 494422 63418 494604 63654
rect 494004 63334 494604 63418
rect 494004 63098 494186 63334
rect 494422 63098 494604 63334
rect 494004 27654 494604 63098
rect 494004 27418 494186 27654
rect 494422 27418 494604 27654
rect 494004 27334 494604 27418
rect 494004 27098 494186 27334
rect 494422 27098 494604 27334
rect 494004 -5046 494604 27098
rect 494004 -5282 494186 -5046
rect 494422 -5282 494604 -5046
rect 494004 -5366 494604 -5282
rect 494004 -5602 494186 -5366
rect 494422 -5602 494604 -5366
rect 494004 -5624 494604 -5602
rect 497604 679254 498204 710862
rect 515604 710478 516204 711440
rect 515604 710242 515786 710478
rect 516022 710242 516204 710478
rect 515604 710158 516204 710242
rect 515604 709922 515786 710158
rect 516022 709922 516204 710158
rect 512004 708598 512604 709560
rect 512004 708362 512186 708598
rect 512422 708362 512604 708598
rect 512004 708278 512604 708362
rect 512004 708042 512186 708278
rect 512422 708042 512604 708278
rect 508404 706718 509004 707680
rect 508404 706482 508586 706718
rect 508822 706482 509004 706718
rect 508404 706398 509004 706482
rect 508404 706162 508586 706398
rect 508822 706162 509004 706398
rect 497604 679018 497786 679254
rect 498022 679018 498204 679254
rect 497604 678934 498204 679018
rect 497604 678698 497786 678934
rect 498022 678698 498204 678934
rect 497604 643254 498204 678698
rect 497604 643018 497786 643254
rect 498022 643018 498204 643254
rect 497604 642934 498204 643018
rect 497604 642698 497786 642934
rect 498022 642698 498204 642934
rect 497604 607254 498204 642698
rect 497604 607018 497786 607254
rect 498022 607018 498204 607254
rect 497604 606934 498204 607018
rect 497604 606698 497786 606934
rect 498022 606698 498204 606934
rect 497604 571254 498204 606698
rect 497604 571018 497786 571254
rect 498022 571018 498204 571254
rect 497604 570934 498204 571018
rect 497604 570698 497786 570934
rect 498022 570698 498204 570934
rect 497604 535254 498204 570698
rect 497604 535018 497786 535254
rect 498022 535018 498204 535254
rect 497604 534934 498204 535018
rect 497604 534698 497786 534934
rect 498022 534698 498204 534934
rect 497604 499254 498204 534698
rect 497604 499018 497786 499254
rect 498022 499018 498204 499254
rect 497604 498934 498204 499018
rect 497604 498698 497786 498934
rect 498022 498698 498204 498934
rect 497604 463254 498204 498698
rect 497604 463018 497786 463254
rect 498022 463018 498204 463254
rect 497604 462934 498204 463018
rect 497604 462698 497786 462934
rect 498022 462698 498204 462934
rect 497604 427254 498204 462698
rect 497604 427018 497786 427254
rect 498022 427018 498204 427254
rect 497604 426934 498204 427018
rect 497604 426698 497786 426934
rect 498022 426698 498204 426934
rect 497604 391254 498204 426698
rect 497604 391018 497786 391254
rect 498022 391018 498204 391254
rect 497604 390934 498204 391018
rect 497604 390698 497786 390934
rect 498022 390698 498204 390934
rect 497604 355254 498204 390698
rect 497604 355018 497786 355254
rect 498022 355018 498204 355254
rect 497604 354934 498204 355018
rect 497604 354698 497786 354934
rect 498022 354698 498204 354934
rect 497604 319254 498204 354698
rect 497604 319018 497786 319254
rect 498022 319018 498204 319254
rect 497604 318934 498204 319018
rect 497604 318698 497786 318934
rect 498022 318698 498204 318934
rect 497604 283254 498204 318698
rect 497604 283018 497786 283254
rect 498022 283018 498204 283254
rect 497604 282934 498204 283018
rect 497604 282698 497786 282934
rect 498022 282698 498204 282934
rect 497604 247254 498204 282698
rect 497604 247018 497786 247254
rect 498022 247018 498204 247254
rect 497604 246934 498204 247018
rect 497604 246698 497786 246934
rect 498022 246698 498204 246934
rect 497604 211254 498204 246698
rect 497604 211018 497786 211254
rect 498022 211018 498204 211254
rect 497604 210934 498204 211018
rect 497604 210698 497786 210934
rect 498022 210698 498204 210934
rect 497604 175254 498204 210698
rect 497604 175018 497786 175254
rect 498022 175018 498204 175254
rect 497604 174934 498204 175018
rect 497604 174698 497786 174934
rect 498022 174698 498204 174934
rect 497604 139254 498204 174698
rect 497604 139018 497786 139254
rect 498022 139018 498204 139254
rect 497604 138934 498204 139018
rect 497604 138698 497786 138934
rect 498022 138698 498204 138934
rect 497604 103254 498204 138698
rect 497604 103018 497786 103254
rect 498022 103018 498204 103254
rect 497604 102934 498204 103018
rect 497604 102698 497786 102934
rect 498022 102698 498204 102934
rect 497604 67254 498204 102698
rect 497604 67018 497786 67254
rect 498022 67018 498204 67254
rect 497604 66934 498204 67018
rect 497604 66698 497786 66934
rect 498022 66698 498204 66934
rect 497604 31254 498204 66698
rect 497604 31018 497786 31254
rect 498022 31018 498204 31254
rect 497604 30934 498204 31018
rect 497604 30698 497786 30934
rect 498022 30698 498204 30934
rect 479604 -6222 479786 -5986
rect 480022 -6222 480204 -5986
rect 479604 -6306 480204 -6222
rect 479604 -6542 479786 -6306
rect 480022 -6542 480204 -6306
rect 479604 -7504 480204 -6542
rect 497604 -6926 498204 30698
rect 504804 704838 505404 705800
rect 504804 704602 504986 704838
rect 505222 704602 505404 704838
rect 504804 704518 505404 704602
rect 504804 704282 504986 704518
rect 505222 704282 505404 704518
rect 504804 686454 505404 704282
rect 504804 686218 504986 686454
rect 505222 686218 505404 686454
rect 504804 686134 505404 686218
rect 504804 685898 504986 686134
rect 505222 685898 505404 686134
rect 504804 650454 505404 685898
rect 504804 650218 504986 650454
rect 505222 650218 505404 650454
rect 504804 650134 505404 650218
rect 504804 649898 504986 650134
rect 505222 649898 505404 650134
rect 504804 614454 505404 649898
rect 504804 614218 504986 614454
rect 505222 614218 505404 614454
rect 504804 614134 505404 614218
rect 504804 613898 504986 614134
rect 505222 613898 505404 614134
rect 504804 578454 505404 613898
rect 504804 578218 504986 578454
rect 505222 578218 505404 578454
rect 504804 578134 505404 578218
rect 504804 577898 504986 578134
rect 505222 577898 505404 578134
rect 504804 542454 505404 577898
rect 504804 542218 504986 542454
rect 505222 542218 505404 542454
rect 504804 542134 505404 542218
rect 504804 541898 504986 542134
rect 505222 541898 505404 542134
rect 504804 506454 505404 541898
rect 504804 506218 504986 506454
rect 505222 506218 505404 506454
rect 504804 506134 505404 506218
rect 504804 505898 504986 506134
rect 505222 505898 505404 506134
rect 504804 470454 505404 505898
rect 504804 470218 504986 470454
rect 505222 470218 505404 470454
rect 504804 470134 505404 470218
rect 504804 469898 504986 470134
rect 505222 469898 505404 470134
rect 504804 434454 505404 469898
rect 504804 434218 504986 434454
rect 505222 434218 505404 434454
rect 504804 434134 505404 434218
rect 504804 433898 504986 434134
rect 505222 433898 505404 434134
rect 504804 398454 505404 433898
rect 504804 398218 504986 398454
rect 505222 398218 505404 398454
rect 504804 398134 505404 398218
rect 504804 397898 504986 398134
rect 505222 397898 505404 398134
rect 504804 362454 505404 397898
rect 504804 362218 504986 362454
rect 505222 362218 505404 362454
rect 504804 362134 505404 362218
rect 504804 361898 504986 362134
rect 505222 361898 505404 362134
rect 504804 326454 505404 361898
rect 504804 326218 504986 326454
rect 505222 326218 505404 326454
rect 504804 326134 505404 326218
rect 504804 325898 504986 326134
rect 505222 325898 505404 326134
rect 504804 290454 505404 325898
rect 504804 290218 504986 290454
rect 505222 290218 505404 290454
rect 504804 290134 505404 290218
rect 504804 289898 504986 290134
rect 505222 289898 505404 290134
rect 504804 254454 505404 289898
rect 504804 254218 504986 254454
rect 505222 254218 505404 254454
rect 504804 254134 505404 254218
rect 504804 253898 504986 254134
rect 505222 253898 505404 254134
rect 504804 218454 505404 253898
rect 504804 218218 504986 218454
rect 505222 218218 505404 218454
rect 504804 218134 505404 218218
rect 504804 217898 504986 218134
rect 505222 217898 505404 218134
rect 504804 182454 505404 217898
rect 504804 182218 504986 182454
rect 505222 182218 505404 182454
rect 504804 182134 505404 182218
rect 504804 181898 504986 182134
rect 505222 181898 505404 182134
rect 504804 146454 505404 181898
rect 504804 146218 504986 146454
rect 505222 146218 505404 146454
rect 504804 146134 505404 146218
rect 504804 145898 504986 146134
rect 505222 145898 505404 146134
rect 504804 110454 505404 145898
rect 504804 110218 504986 110454
rect 505222 110218 505404 110454
rect 504804 110134 505404 110218
rect 504804 109898 504986 110134
rect 505222 109898 505404 110134
rect 504804 74454 505404 109898
rect 504804 74218 504986 74454
rect 505222 74218 505404 74454
rect 504804 74134 505404 74218
rect 504804 73898 504986 74134
rect 505222 73898 505404 74134
rect 504804 38454 505404 73898
rect 504804 38218 504986 38454
rect 505222 38218 505404 38454
rect 504804 38134 505404 38218
rect 504804 37898 504986 38134
rect 505222 37898 505404 38134
rect 504804 2454 505404 37898
rect 504804 2218 504986 2454
rect 505222 2218 505404 2454
rect 504804 2134 505404 2218
rect 504804 1898 504986 2134
rect 505222 1898 505404 2134
rect 504804 -346 505404 1898
rect 504804 -582 504986 -346
rect 505222 -582 505404 -346
rect 504804 -666 505404 -582
rect 504804 -902 504986 -666
rect 505222 -902 505404 -666
rect 504804 -1864 505404 -902
rect 508404 690054 509004 706162
rect 508404 689818 508586 690054
rect 508822 689818 509004 690054
rect 508404 689734 509004 689818
rect 508404 689498 508586 689734
rect 508822 689498 509004 689734
rect 508404 654054 509004 689498
rect 508404 653818 508586 654054
rect 508822 653818 509004 654054
rect 508404 653734 509004 653818
rect 508404 653498 508586 653734
rect 508822 653498 509004 653734
rect 508404 618054 509004 653498
rect 508404 617818 508586 618054
rect 508822 617818 509004 618054
rect 508404 617734 509004 617818
rect 508404 617498 508586 617734
rect 508822 617498 509004 617734
rect 508404 582054 509004 617498
rect 508404 581818 508586 582054
rect 508822 581818 509004 582054
rect 508404 581734 509004 581818
rect 508404 581498 508586 581734
rect 508822 581498 509004 581734
rect 508404 546054 509004 581498
rect 508404 545818 508586 546054
rect 508822 545818 509004 546054
rect 508404 545734 509004 545818
rect 508404 545498 508586 545734
rect 508822 545498 509004 545734
rect 508404 510054 509004 545498
rect 508404 509818 508586 510054
rect 508822 509818 509004 510054
rect 508404 509734 509004 509818
rect 508404 509498 508586 509734
rect 508822 509498 509004 509734
rect 508404 474054 509004 509498
rect 508404 473818 508586 474054
rect 508822 473818 509004 474054
rect 508404 473734 509004 473818
rect 508404 473498 508586 473734
rect 508822 473498 509004 473734
rect 508404 438054 509004 473498
rect 508404 437818 508586 438054
rect 508822 437818 509004 438054
rect 508404 437734 509004 437818
rect 508404 437498 508586 437734
rect 508822 437498 509004 437734
rect 508404 402054 509004 437498
rect 508404 401818 508586 402054
rect 508822 401818 509004 402054
rect 508404 401734 509004 401818
rect 508404 401498 508586 401734
rect 508822 401498 509004 401734
rect 508404 366054 509004 401498
rect 508404 365818 508586 366054
rect 508822 365818 509004 366054
rect 508404 365734 509004 365818
rect 508404 365498 508586 365734
rect 508822 365498 509004 365734
rect 508404 330054 509004 365498
rect 508404 329818 508586 330054
rect 508822 329818 509004 330054
rect 508404 329734 509004 329818
rect 508404 329498 508586 329734
rect 508822 329498 509004 329734
rect 508404 294054 509004 329498
rect 508404 293818 508586 294054
rect 508822 293818 509004 294054
rect 508404 293734 509004 293818
rect 508404 293498 508586 293734
rect 508822 293498 509004 293734
rect 508404 258054 509004 293498
rect 508404 257818 508586 258054
rect 508822 257818 509004 258054
rect 508404 257734 509004 257818
rect 508404 257498 508586 257734
rect 508822 257498 509004 257734
rect 508404 222054 509004 257498
rect 508404 221818 508586 222054
rect 508822 221818 509004 222054
rect 508404 221734 509004 221818
rect 508404 221498 508586 221734
rect 508822 221498 509004 221734
rect 508404 186054 509004 221498
rect 508404 185818 508586 186054
rect 508822 185818 509004 186054
rect 508404 185734 509004 185818
rect 508404 185498 508586 185734
rect 508822 185498 509004 185734
rect 508404 150054 509004 185498
rect 508404 149818 508586 150054
rect 508822 149818 509004 150054
rect 508404 149734 509004 149818
rect 508404 149498 508586 149734
rect 508822 149498 509004 149734
rect 508404 114054 509004 149498
rect 508404 113818 508586 114054
rect 508822 113818 509004 114054
rect 508404 113734 509004 113818
rect 508404 113498 508586 113734
rect 508822 113498 509004 113734
rect 508404 78054 509004 113498
rect 508404 77818 508586 78054
rect 508822 77818 509004 78054
rect 508404 77734 509004 77818
rect 508404 77498 508586 77734
rect 508822 77498 509004 77734
rect 508404 42054 509004 77498
rect 508404 41818 508586 42054
rect 508822 41818 509004 42054
rect 508404 41734 509004 41818
rect 508404 41498 508586 41734
rect 508822 41498 509004 41734
rect 508404 6054 509004 41498
rect 508404 5818 508586 6054
rect 508822 5818 509004 6054
rect 508404 5734 509004 5818
rect 508404 5498 508586 5734
rect 508822 5498 509004 5734
rect 508404 -2226 509004 5498
rect 508404 -2462 508586 -2226
rect 508822 -2462 509004 -2226
rect 508404 -2546 509004 -2462
rect 508404 -2782 508586 -2546
rect 508822 -2782 509004 -2546
rect 508404 -3744 509004 -2782
rect 512004 693654 512604 708042
rect 512004 693418 512186 693654
rect 512422 693418 512604 693654
rect 512004 693334 512604 693418
rect 512004 693098 512186 693334
rect 512422 693098 512604 693334
rect 512004 657654 512604 693098
rect 512004 657418 512186 657654
rect 512422 657418 512604 657654
rect 512004 657334 512604 657418
rect 512004 657098 512186 657334
rect 512422 657098 512604 657334
rect 512004 621654 512604 657098
rect 512004 621418 512186 621654
rect 512422 621418 512604 621654
rect 512004 621334 512604 621418
rect 512004 621098 512186 621334
rect 512422 621098 512604 621334
rect 512004 585654 512604 621098
rect 512004 585418 512186 585654
rect 512422 585418 512604 585654
rect 512004 585334 512604 585418
rect 512004 585098 512186 585334
rect 512422 585098 512604 585334
rect 512004 549654 512604 585098
rect 512004 549418 512186 549654
rect 512422 549418 512604 549654
rect 512004 549334 512604 549418
rect 512004 549098 512186 549334
rect 512422 549098 512604 549334
rect 512004 513654 512604 549098
rect 512004 513418 512186 513654
rect 512422 513418 512604 513654
rect 512004 513334 512604 513418
rect 512004 513098 512186 513334
rect 512422 513098 512604 513334
rect 512004 477654 512604 513098
rect 512004 477418 512186 477654
rect 512422 477418 512604 477654
rect 512004 477334 512604 477418
rect 512004 477098 512186 477334
rect 512422 477098 512604 477334
rect 512004 441654 512604 477098
rect 512004 441418 512186 441654
rect 512422 441418 512604 441654
rect 512004 441334 512604 441418
rect 512004 441098 512186 441334
rect 512422 441098 512604 441334
rect 512004 405654 512604 441098
rect 512004 405418 512186 405654
rect 512422 405418 512604 405654
rect 512004 405334 512604 405418
rect 512004 405098 512186 405334
rect 512422 405098 512604 405334
rect 512004 369654 512604 405098
rect 512004 369418 512186 369654
rect 512422 369418 512604 369654
rect 512004 369334 512604 369418
rect 512004 369098 512186 369334
rect 512422 369098 512604 369334
rect 512004 333654 512604 369098
rect 512004 333418 512186 333654
rect 512422 333418 512604 333654
rect 512004 333334 512604 333418
rect 512004 333098 512186 333334
rect 512422 333098 512604 333334
rect 512004 297654 512604 333098
rect 512004 297418 512186 297654
rect 512422 297418 512604 297654
rect 512004 297334 512604 297418
rect 512004 297098 512186 297334
rect 512422 297098 512604 297334
rect 512004 261654 512604 297098
rect 512004 261418 512186 261654
rect 512422 261418 512604 261654
rect 512004 261334 512604 261418
rect 512004 261098 512186 261334
rect 512422 261098 512604 261334
rect 512004 225654 512604 261098
rect 512004 225418 512186 225654
rect 512422 225418 512604 225654
rect 512004 225334 512604 225418
rect 512004 225098 512186 225334
rect 512422 225098 512604 225334
rect 512004 189654 512604 225098
rect 512004 189418 512186 189654
rect 512422 189418 512604 189654
rect 512004 189334 512604 189418
rect 512004 189098 512186 189334
rect 512422 189098 512604 189334
rect 512004 153654 512604 189098
rect 512004 153418 512186 153654
rect 512422 153418 512604 153654
rect 512004 153334 512604 153418
rect 512004 153098 512186 153334
rect 512422 153098 512604 153334
rect 512004 117654 512604 153098
rect 512004 117418 512186 117654
rect 512422 117418 512604 117654
rect 512004 117334 512604 117418
rect 512004 117098 512186 117334
rect 512422 117098 512604 117334
rect 512004 81654 512604 117098
rect 512004 81418 512186 81654
rect 512422 81418 512604 81654
rect 512004 81334 512604 81418
rect 512004 81098 512186 81334
rect 512422 81098 512604 81334
rect 512004 45654 512604 81098
rect 512004 45418 512186 45654
rect 512422 45418 512604 45654
rect 512004 45334 512604 45418
rect 512004 45098 512186 45334
rect 512422 45098 512604 45334
rect 512004 9654 512604 45098
rect 512004 9418 512186 9654
rect 512422 9418 512604 9654
rect 512004 9334 512604 9418
rect 512004 9098 512186 9334
rect 512422 9098 512604 9334
rect 512004 -4106 512604 9098
rect 512004 -4342 512186 -4106
rect 512422 -4342 512604 -4106
rect 512004 -4426 512604 -4342
rect 512004 -4662 512186 -4426
rect 512422 -4662 512604 -4426
rect 512004 -5624 512604 -4662
rect 515604 697254 516204 709922
rect 533604 711418 534204 711440
rect 533604 711182 533786 711418
rect 534022 711182 534204 711418
rect 533604 711098 534204 711182
rect 533604 710862 533786 711098
rect 534022 710862 534204 711098
rect 530004 709538 530604 709560
rect 530004 709302 530186 709538
rect 530422 709302 530604 709538
rect 530004 709218 530604 709302
rect 530004 708982 530186 709218
rect 530422 708982 530604 709218
rect 526404 707658 527004 707680
rect 526404 707422 526586 707658
rect 526822 707422 527004 707658
rect 526404 707338 527004 707422
rect 526404 707102 526586 707338
rect 526822 707102 527004 707338
rect 515604 697018 515786 697254
rect 516022 697018 516204 697254
rect 515604 696934 516204 697018
rect 515604 696698 515786 696934
rect 516022 696698 516204 696934
rect 515604 661254 516204 696698
rect 515604 661018 515786 661254
rect 516022 661018 516204 661254
rect 515604 660934 516204 661018
rect 515604 660698 515786 660934
rect 516022 660698 516204 660934
rect 515604 625254 516204 660698
rect 515604 625018 515786 625254
rect 516022 625018 516204 625254
rect 515604 624934 516204 625018
rect 515604 624698 515786 624934
rect 516022 624698 516204 624934
rect 515604 589254 516204 624698
rect 515604 589018 515786 589254
rect 516022 589018 516204 589254
rect 515604 588934 516204 589018
rect 515604 588698 515786 588934
rect 516022 588698 516204 588934
rect 515604 553254 516204 588698
rect 515604 553018 515786 553254
rect 516022 553018 516204 553254
rect 515604 552934 516204 553018
rect 515604 552698 515786 552934
rect 516022 552698 516204 552934
rect 515604 517254 516204 552698
rect 515604 517018 515786 517254
rect 516022 517018 516204 517254
rect 515604 516934 516204 517018
rect 515604 516698 515786 516934
rect 516022 516698 516204 516934
rect 515604 481254 516204 516698
rect 515604 481018 515786 481254
rect 516022 481018 516204 481254
rect 515604 480934 516204 481018
rect 515604 480698 515786 480934
rect 516022 480698 516204 480934
rect 515604 445254 516204 480698
rect 515604 445018 515786 445254
rect 516022 445018 516204 445254
rect 515604 444934 516204 445018
rect 515604 444698 515786 444934
rect 516022 444698 516204 444934
rect 515604 409254 516204 444698
rect 515604 409018 515786 409254
rect 516022 409018 516204 409254
rect 515604 408934 516204 409018
rect 515604 408698 515786 408934
rect 516022 408698 516204 408934
rect 515604 373254 516204 408698
rect 515604 373018 515786 373254
rect 516022 373018 516204 373254
rect 515604 372934 516204 373018
rect 515604 372698 515786 372934
rect 516022 372698 516204 372934
rect 515604 337254 516204 372698
rect 515604 337018 515786 337254
rect 516022 337018 516204 337254
rect 515604 336934 516204 337018
rect 515604 336698 515786 336934
rect 516022 336698 516204 336934
rect 515604 301254 516204 336698
rect 515604 301018 515786 301254
rect 516022 301018 516204 301254
rect 515604 300934 516204 301018
rect 515604 300698 515786 300934
rect 516022 300698 516204 300934
rect 515604 265254 516204 300698
rect 515604 265018 515786 265254
rect 516022 265018 516204 265254
rect 515604 264934 516204 265018
rect 515604 264698 515786 264934
rect 516022 264698 516204 264934
rect 515604 229254 516204 264698
rect 515604 229018 515786 229254
rect 516022 229018 516204 229254
rect 515604 228934 516204 229018
rect 515604 228698 515786 228934
rect 516022 228698 516204 228934
rect 515604 193254 516204 228698
rect 515604 193018 515786 193254
rect 516022 193018 516204 193254
rect 515604 192934 516204 193018
rect 515604 192698 515786 192934
rect 516022 192698 516204 192934
rect 515604 157254 516204 192698
rect 515604 157018 515786 157254
rect 516022 157018 516204 157254
rect 515604 156934 516204 157018
rect 515604 156698 515786 156934
rect 516022 156698 516204 156934
rect 515604 121254 516204 156698
rect 515604 121018 515786 121254
rect 516022 121018 516204 121254
rect 515604 120934 516204 121018
rect 515604 120698 515786 120934
rect 516022 120698 516204 120934
rect 515604 85254 516204 120698
rect 515604 85018 515786 85254
rect 516022 85018 516204 85254
rect 515604 84934 516204 85018
rect 515604 84698 515786 84934
rect 516022 84698 516204 84934
rect 515604 49254 516204 84698
rect 515604 49018 515786 49254
rect 516022 49018 516204 49254
rect 515604 48934 516204 49018
rect 515604 48698 515786 48934
rect 516022 48698 516204 48934
rect 515604 13254 516204 48698
rect 515604 13018 515786 13254
rect 516022 13018 516204 13254
rect 515604 12934 516204 13018
rect 515604 12698 515786 12934
rect 516022 12698 516204 12934
rect 497604 -7162 497786 -6926
rect 498022 -7162 498204 -6926
rect 497604 -7246 498204 -7162
rect 497604 -7482 497786 -7246
rect 498022 -7482 498204 -7246
rect 497604 -7504 498204 -7482
rect 515604 -5986 516204 12698
rect 522804 705778 523404 705800
rect 522804 705542 522986 705778
rect 523222 705542 523404 705778
rect 522804 705458 523404 705542
rect 522804 705222 522986 705458
rect 523222 705222 523404 705458
rect 522804 668454 523404 705222
rect 522804 668218 522986 668454
rect 523222 668218 523404 668454
rect 522804 668134 523404 668218
rect 522804 667898 522986 668134
rect 523222 667898 523404 668134
rect 522804 632454 523404 667898
rect 522804 632218 522986 632454
rect 523222 632218 523404 632454
rect 522804 632134 523404 632218
rect 522804 631898 522986 632134
rect 523222 631898 523404 632134
rect 522804 596454 523404 631898
rect 522804 596218 522986 596454
rect 523222 596218 523404 596454
rect 522804 596134 523404 596218
rect 522804 595898 522986 596134
rect 523222 595898 523404 596134
rect 522804 560454 523404 595898
rect 522804 560218 522986 560454
rect 523222 560218 523404 560454
rect 522804 560134 523404 560218
rect 522804 559898 522986 560134
rect 523222 559898 523404 560134
rect 522804 524454 523404 559898
rect 522804 524218 522986 524454
rect 523222 524218 523404 524454
rect 522804 524134 523404 524218
rect 522804 523898 522986 524134
rect 523222 523898 523404 524134
rect 522804 488454 523404 523898
rect 522804 488218 522986 488454
rect 523222 488218 523404 488454
rect 522804 488134 523404 488218
rect 522804 487898 522986 488134
rect 523222 487898 523404 488134
rect 522804 452454 523404 487898
rect 522804 452218 522986 452454
rect 523222 452218 523404 452454
rect 522804 452134 523404 452218
rect 522804 451898 522986 452134
rect 523222 451898 523404 452134
rect 522804 416454 523404 451898
rect 522804 416218 522986 416454
rect 523222 416218 523404 416454
rect 522804 416134 523404 416218
rect 522804 415898 522986 416134
rect 523222 415898 523404 416134
rect 522804 380454 523404 415898
rect 522804 380218 522986 380454
rect 523222 380218 523404 380454
rect 522804 380134 523404 380218
rect 522804 379898 522986 380134
rect 523222 379898 523404 380134
rect 522804 344454 523404 379898
rect 522804 344218 522986 344454
rect 523222 344218 523404 344454
rect 522804 344134 523404 344218
rect 522804 343898 522986 344134
rect 523222 343898 523404 344134
rect 522804 308454 523404 343898
rect 522804 308218 522986 308454
rect 523222 308218 523404 308454
rect 522804 308134 523404 308218
rect 522804 307898 522986 308134
rect 523222 307898 523404 308134
rect 522804 272454 523404 307898
rect 522804 272218 522986 272454
rect 523222 272218 523404 272454
rect 522804 272134 523404 272218
rect 522804 271898 522986 272134
rect 523222 271898 523404 272134
rect 522804 236454 523404 271898
rect 522804 236218 522986 236454
rect 523222 236218 523404 236454
rect 522804 236134 523404 236218
rect 522804 235898 522986 236134
rect 523222 235898 523404 236134
rect 522804 200454 523404 235898
rect 522804 200218 522986 200454
rect 523222 200218 523404 200454
rect 522804 200134 523404 200218
rect 522804 199898 522986 200134
rect 523222 199898 523404 200134
rect 522804 164454 523404 199898
rect 522804 164218 522986 164454
rect 523222 164218 523404 164454
rect 522804 164134 523404 164218
rect 522804 163898 522986 164134
rect 523222 163898 523404 164134
rect 522804 128454 523404 163898
rect 522804 128218 522986 128454
rect 523222 128218 523404 128454
rect 522804 128134 523404 128218
rect 522804 127898 522986 128134
rect 523222 127898 523404 128134
rect 522804 92454 523404 127898
rect 522804 92218 522986 92454
rect 523222 92218 523404 92454
rect 522804 92134 523404 92218
rect 522804 91898 522986 92134
rect 523222 91898 523404 92134
rect 522804 56454 523404 91898
rect 522804 56218 522986 56454
rect 523222 56218 523404 56454
rect 522804 56134 523404 56218
rect 522804 55898 522986 56134
rect 523222 55898 523404 56134
rect 522804 20454 523404 55898
rect 522804 20218 522986 20454
rect 523222 20218 523404 20454
rect 522804 20134 523404 20218
rect 522804 19898 522986 20134
rect 523222 19898 523404 20134
rect 522804 -1286 523404 19898
rect 522804 -1522 522986 -1286
rect 523222 -1522 523404 -1286
rect 522804 -1606 523404 -1522
rect 522804 -1842 522986 -1606
rect 523222 -1842 523404 -1606
rect 522804 -1864 523404 -1842
rect 526404 672054 527004 707102
rect 526404 671818 526586 672054
rect 526822 671818 527004 672054
rect 526404 671734 527004 671818
rect 526404 671498 526586 671734
rect 526822 671498 527004 671734
rect 526404 636054 527004 671498
rect 526404 635818 526586 636054
rect 526822 635818 527004 636054
rect 526404 635734 527004 635818
rect 526404 635498 526586 635734
rect 526822 635498 527004 635734
rect 526404 600054 527004 635498
rect 526404 599818 526586 600054
rect 526822 599818 527004 600054
rect 526404 599734 527004 599818
rect 526404 599498 526586 599734
rect 526822 599498 527004 599734
rect 526404 564054 527004 599498
rect 526404 563818 526586 564054
rect 526822 563818 527004 564054
rect 526404 563734 527004 563818
rect 526404 563498 526586 563734
rect 526822 563498 527004 563734
rect 526404 528054 527004 563498
rect 526404 527818 526586 528054
rect 526822 527818 527004 528054
rect 526404 527734 527004 527818
rect 526404 527498 526586 527734
rect 526822 527498 527004 527734
rect 526404 492054 527004 527498
rect 526404 491818 526586 492054
rect 526822 491818 527004 492054
rect 526404 491734 527004 491818
rect 526404 491498 526586 491734
rect 526822 491498 527004 491734
rect 526404 456054 527004 491498
rect 526404 455818 526586 456054
rect 526822 455818 527004 456054
rect 526404 455734 527004 455818
rect 526404 455498 526586 455734
rect 526822 455498 527004 455734
rect 526404 420054 527004 455498
rect 526404 419818 526586 420054
rect 526822 419818 527004 420054
rect 526404 419734 527004 419818
rect 526404 419498 526586 419734
rect 526822 419498 527004 419734
rect 526404 384054 527004 419498
rect 526404 383818 526586 384054
rect 526822 383818 527004 384054
rect 526404 383734 527004 383818
rect 526404 383498 526586 383734
rect 526822 383498 527004 383734
rect 526404 348054 527004 383498
rect 526404 347818 526586 348054
rect 526822 347818 527004 348054
rect 526404 347734 527004 347818
rect 526404 347498 526586 347734
rect 526822 347498 527004 347734
rect 526404 312054 527004 347498
rect 526404 311818 526586 312054
rect 526822 311818 527004 312054
rect 526404 311734 527004 311818
rect 526404 311498 526586 311734
rect 526822 311498 527004 311734
rect 526404 276054 527004 311498
rect 526404 275818 526586 276054
rect 526822 275818 527004 276054
rect 526404 275734 527004 275818
rect 526404 275498 526586 275734
rect 526822 275498 527004 275734
rect 526404 240054 527004 275498
rect 526404 239818 526586 240054
rect 526822 239818 527004 240054
rect 526404 239734 527004 239818
rect 526404 239498 526586 239734
rect 526822 239498 527004 239734
rect 526404 204054 527004 239498
rect 526404 203818 526586 204054
rect 526822 203818 527004 204054
rect 526404 203734 527004 203818
rect 526404 203498 526586 203734
rect 526822 203498 527004 203734
rect 526404 168054 527004 203498
rect 526404 167818 526586 168054
rect 526822 167818 527004 168054
rect 526404 167734 527004 167818
rect 526404 167498 526586 167734
rect 526822 167498 527004 167734
rect 526404 132054 527004 167498
rect 526404 131818 526586 132054
rect 526822 131818 527004 132054
rect 526404 131734 527004 131818
rect 526404 131498 526586 131734
rect 526822 131498 527004 131734
rect 526404 96054 527004 131498
rect 526404 95818 526586 96054
rect 526822 95818 527004 96054
rect 526404 95734 527004 95818
rect 526404 95498 526586 95734
rect 526822 95498 527004 95734
rect 526404 60054 527004 95498
rect 526404 59818 526586 60054
rect 526822 59818 527004 60054
rect 526404 59734 527004 59818
rect 526404 59498 526586 59734
rect 526822 59498 527004 59734
rect 526404 24054 527004 59498
rect 526404 23818 526586 24054
rect 526822 23818 527004 24054
rect 526404 23734 527004 23818
rect 526404 23498 526586 23734
rect 526822 23498 527004 23734
rect 526404 -3166 527004 23498
rect 526404 -3402 526586 -3166
rect 526822 -3402 527004 -3166
rect 526404 -3486 527004 -3402
rect 526404 -3722 526586 -3486
rect 526822 -3722 527004 -3486
rect 526404 -3744 527004 -3722
rect 530004 675654 530604 708982
rect 530004 675418 530186 675654
rect 530422 675418 530604 675654
rect 530004 675334 530604 675418
rect 530004 675098 530186 675334
rect 530422 675098 530604 675334
rect 530004 639654 530604 675098
rect 530004 639418 530186 639654
rect 530422 639418 530604 639654
rect 530004 639334 530604 639418
rect 530004 639098 530186 639334
rect 530422 639098 530604 639334
rect 530004 603654 530604 639098
rect 530004 603418 530186 603654
rect 530422 603418 530604 603654
rect 530004 603334 530604 603418
rect 530004 603098 530186 603334
rect 530422 603098 530604 603334
rect 530004 567654 530604 603098
rect 530004 567418 530186 567654
rect 530422 567418 530604 567654
rect 530004 567334 530604 567418
rect 530004 567098 530186 567334
rect 530422 567098 530604 567334
rect 530004 531654 530604 567098
rect 530004 531418 530186 531654
rect 530422 531418 530604 531654
rect 530004 531334 530604 531418
rect 530004 531098 530186 531334
rect 530422 531098 530604 531334
rect 530004 495654 530604 531098
rect 530004 495418 530186 495654
rect 530422 495418 530604 495654
rect 530004 495334 530604 495418
rect 530004 495098 530186 495334
rect 530422 495098 530604 495334
rect 530004 459654 530604 495098
rect 530004 459418 530186 459654
rect 530422 459418 530604 459654
rect 530004 459334 530604 459418
rect 530004 459098 530186 459334
rect 530422 459098 530604 459334
rect 530004 423654 530604 459098
rect 530004 423418 530186 423654
rect 530422 423418 530604 423654
rect 530004 423334 530604 423418
rect 530004 423098 530186 423334
rect 530422 423098 530604 423334
rect 530004 387654 530604 423098
rect 530004 387418 530186 387654
rect 530422 387418 530604 387654
rect 530004 387334 530604 387418
rect 530004 387098 530186 387334
rect 530422 387098 530604 387334
rect 530004 351654 530604 387098
rect 530004 351418 530186 351654
rect 530422 351418 530604 351654
rect 530004 351334 530604 351418
rect 530004 351098 530186 351334
rect 530422 351098 530604 351334
rect 530004 315654 530604 351098
rect 530004 315418 530186 315654
rect 530422 315418 530604 315654
rect 530004 315334 530604 315418
rect 530004 315098 530186 315334
rect 530422 315098 530604 315334
rect 530004 279654 530604 315098
rect 530004 279418 530186 279654
rect 530422 279418 530604 279654
rect 530004 279334 530604 279418
rect 530004 279098 530186 279334
rect 530422 279098 530604 279334
rect 530004 243654 530604 279098
rect 530004 243418 530186 243654
rect 530422 243418 530604 243654
rect 530004 243334 530604 243418
rect 530004 243098 530186 243334
rect 530422 243098 530604 243334
rect 530004 207654 530604 243098
rect 530004 207418 530186 207654
rect 530422 207418 530604 207654
rect 530004 207334 530604 207418
rect 530004 207098 530186 207334
rect 530422 207098 530604 207334
rect 530004 171654 530604 207098
rect 530004 171418 530186 171654
rect 530422 171418 530604 171654
rect 530004 171334 530604 171418
rect 530004 171098 530186 171334
rect 530422 171098 530604 171334
rect 530004 135654 530604 171098
rect 530004 135418 530186 135654
rect 530422 135418 530604 135654
rect 530004 135334 530604 135418
rect 530004 135098 530186 135334
rect 530422 135098 530604 135334
rect 530004 99654 530604 135098
rect 530004 99418 530186 99654
rect 530422 99418 530604 99654
rect 530004 99334 530604 99418
rect 530004 99098 530186 99334
rect 530422 99098 530604 99334
rect 530004 63654 530604 99098
rect 530004 63418 530186 63654
rect 530422 63418 530604 63654
rect 530004 63334 530604 63418
rect 530004 63098 530186 63334
rect 530422 63098 530604 63334
rect 530004 27654 530604 63098
rect 530004 27418 530186 27654
rect 530422 27418 530604 27654
rect 530004 27334 530604 27418
rect 530004 27098 530186 27334
rect 530422 27098 530604 27334
rect 530004 -5046 530604 27098
rect 530004 -5282 530186 -5046
rect 530422 -5282 530604 -5046
rect 530004 -5366 530604 -5282
rect 530004 -5602 530186 -5366
rect 530422 -5602 530604 -5366
rect 530004 -5624 530604 -5602
rect 533604 679254 534204 710862
rect 551604 710478 552204 711440
rect 551604 710242 551786 710478
rect 552022 710242 552204 710478
rect 551604 710158 552204 710242
rect 551604 709922 551786 710158
rect 552022 709922 552204 710158
rect 548004 708598 548604 709560
rect 548004 708362 548186 708598
rect 548422 708362 548604 708598
rect 548004 708278 548604 708362
rect 548004 708042 548186 708278
rect 548422 708042 548604 708278
rect 544404 706718 545004 707680
rect 544404 706482 544586 706718
rect 544822 706482 545004 706718
rect 544404 706398 545004 706482
rect 544404 706162 544586 706398
rect 544822 706162 545004 706398
rect 533604 679018 533786 679254
rect 534022 679018 534204 679254
rect 533604 678934 534204 679018
rect 533604 678698 533786 678934
rect 534022 678698 534204 678934
rect 533604 643254 534204 678698
rect 533604 643018 533786 643254
rect 534022 643018 534204 643254
rect 533604 642934 534204 643018
rect 533604 642698 533786 642934
rect 534022 642698 534204 642934
rect 533604 607254 534204 642698
rect 533604 607018 533786 607254
rect 534022 607018 534204 607254
rect 533604 606934 534204 607018
rect 533604 606698 533786 606934
rect 534022 606698 534204 606934
rect 533604 571254 534204 606698
rect 533604 571018 533786 571254
rect 534022 571018 534204 571254
rect 533604 570934 534204 571018
rect 533604 570698 533786 570934
rect 534022 570698 534204 570934
rect 533604 535254 534204 570698
rect 533604 535018 533786 535254
rect 534022 535018 534204 535254
rect 533604 534934 534204 535018
rect 533604 534698 533786 534934
rect 534022 534698 534204 534934
rect 533604 499254 534204 534698
rect 533604 499018 533786 499254
rect 534022 499018 534204 499254
rect 533604 498934 534204 499018
rect 533604 498698 533786 498934
rect 534022 498698 534204 498934
rect 533604 463254 534204 498698
rect 533604 463018 533786 463254
rect 534022 463018 534204 463254
rect 533604 462934 534204 463018
rect 533604 462698 533786 462934
rect 534022 462698 534204 462934
rect 533604 427254 534204 462698
rect 533604 427018 533786 427254
rect 534022 427018 534204 427254
rect 533604 426934 534204 427018
rect 533604 426698 533786 426934
rect 534022 426698 534204 426934
rect 533604 391254 534204 426698
rect 533604 391018 533786 391254
rect 534022 391018 534204 391254
rect 533604 390934 534204 391018
rect 533604 390698 533786 390934
rect 534022 390698 534204 390934
rect 533604 355254 534204 390698
rect 533604 355018 533786 355254
rect 534022 355018 534204 355254
rect 533604 354934 534204 355018
rect 533604 354698 533786 354934
rect 534022 354698 534204 354934
rect 533604 319254 534204 354698
rect 533604 319018 533786 319254
rect 534022 319018 534204 319254
rect 533604 318934 534204 319018
rect 533604 318698 533786 318934
rect 534022 318698 534204 318934
rect 533604 283254 534204 318698
rect 533604 283018 533786 283254
rect 534022 283018 534204 283254
rect 533604 282934 534204 283018
rect 533604 282698 533786 282934
rect 534022 282698 534204 282934
rect 533604 247254 534204 282698
rect 533604 247018 533786 247254
rect 534022 247018 534204 247254
rect 533604 246934 534204 247018
rect 533604 246698 533786 246934
rect 534022 246698 534204 246934
rect 533604 211254 534204 246698
rect 533604 211018 533786 211254
rect 534022 211018 534204 211254
rect 533604 210934 534204 211018
rect 533604 210698 533786 210934
rect 534022 210698 534204 210934
rect 533604 175254 534204 210698
rect 533604 175018 533786 175254
rect 534022 175018 534204 175254
rect 533604 174934 534204 175018
rect 533604 174698 533786 174934
rect 534022 174698 534204 174934
rect 533604 139254 534204 174698
rect 533604 139018 533786 139254
rect 534022 139018 534204 139254
rect 533604 138934 534204 139018
rect 533604 138698 533786 138934
rect 534022 138698 534204 138934
rect 533604 103254 534204 138698
rect 533604 103018 533786 103254
rect 534022 103018 534204 103254
rect 533604 102934 534204 103018
rect 533604 102698 533786 102934
rect 534022 102698 534204 102934
rect 533604 67254 534204 102698
rect 533604 67018 533786 67254
rect 534022 67018 534204 67254
rect 533604 66934 534204 67018
rect 533604 66698 533786 66934
rect 534022 66698 534204 66934
rect 533604 31254 534204 66698
rect 533604 31018 533786 31254
rect 534022 31018 534204 31254
rect 533604 30934 534204 31018
rect 533604 30698 533786 30934
rect 534022 30698 534204 30934
rect 515604 -6222 515786 -5986
rect 516022 -6222 516204 -5986
rect 515604 -6306 516204 -6222
rect 515604 -6542 515786 -6306
rect 516022 -6542 516204 -6306
rect 515604 -7504 516204 -6542
rect 533604 -6926 534204 30698
rect 540804 704838 541404 705800
rect 540804 704602 540986 704838
rect 541222 704602 541404 704838
rect 540804 704518 541404 704602
rect 540804 704282 540986 704518
rect 541222 704282 541404 704518
rect 540804 686454 541404 704282
rect 540804 686218 540986 686454
rect 541222 686218 541404 686454
rect 540804 686134 541404 686218
rect 540804 685898 540986 686134
rect 541222 685898 541404 686134
rect 540804 650454 541404 685898
rect 540804 650218 540986 650454
rect 541222 650218 541404 650454
rect 540804 650134 541404 650218
rect 540804 649898 540986 650134
rect 541222 649898 541404 650134
rect 540804 614454 541404 649898
rect 540804 614218 540986 614454
rect 541222 614218 541404 614454
rect 540804 614134 541404 614218
rect 540804 613898 540986 614134
rect 541222 613898 541404 614134
rect 540804 578454 541404 613898
rect 540804 578218 540986 578454
rect 541222 578218 541404 578454
rect 540804 578134 541404 578218
rect 540804 577898 540986 578134
rect 541222 577898 541404 578134
rect 540804 542454 541404 577898
rect 540804 542218 540986 542454
rect 541222 542218 541404 542454
rect 540804 542134 541404 542218
rect 540804 541898 540986 542134
rect 541222 541898 541404 542134
rect 540804 506454 541404 541898
rect 540804 506218 540986 506454
rect 541222 506218 541404 506454
rect 540804 506134 541404 506218
rect 540804 505898 540986 506134
rect 541222 505898 541404 506134
rect 540804 470454 541404 505898
rect 540804 470218 540986 470454
rect 541222 470218 541404 470454
rect 540804 470134 541404 470218
rect 540804 469898 540986 470134
rect 541222 469898 541404 470134
rect 540804 434454 541404 469898
rect 540804 434218 540986 434454
rect 541222 434218 541404 434454
rect 540804 434134 541404 434218
rect 540804 433898 540986 434134
rect 541222 433898 541404 434134
rect 540804 398454 541404 433898
rect 540804 398218 540986 398454
rect 541222 398218 541404 398454
rect 540804 398134 541404 398218
rect 540804 397898 540986 398134
rect 541222 397898 541404 398134
rect 540804 362454 541404 397898
rect 540804 362218 540986 362454
rect 541222 362218 541404 362454
rect 540804 362134 541404 362218
rect 540804 361898 540986 362134
rect 541222 361898 541404 362134
rect 540804 326454 541404 361898
rect 540804 326218 540986 326454
rect 541222 326218 541404 326454
rect 540804 326134 541404 326218
rect 540804 325898 540986 326134
rect 541222 325898 541404 326134
rect 540804 290454 541404 325898
rect 540804 290218 540986 290454
rect 541222 290218 541404 290454
rect 540804 290134 541404 290218
rect 540804 289898 540986 290134
rect 541222 289898 541404 290134
rect 540804 254454 541404 289898
rect 540804 254218 540986 254454
rect 541222 254218 541404 254454
rect 540804 254134 541404 254218
rect 540804 253898 540986 254134
rect 541222 253898 541404 254134
rect 540804 218454 541404 253898
rect 540804 218218 540986 218454
rect 541222 218218 541404 218454
rect 540804 218134 541404 218218
rect 540804 217898 540986 218134
rect 541222 217898 541404 218134
rect 540804 182454 541404 217898
rect 540804 182218 540986 182454
rect 541222 182218 541404 182454
rect 540804 182134 541404 182218
rect 540804 181898 540986 182134
rect 541222 181898 541404 182134
rect 540804 146454 541404 181898
rect 540804 146218 540986 146454
rect 541222 146218 541404 146454
rect 540804 146134 541404 146218
rect 540804 145898 540986 146134
rect 541222 145898 541404 146134
rect 540804 110454 541404 145898
rect 540804 110218 540986 110454
rect 541222 110218 541404 110454
rect 540804 110134 541404 110218
rect 540804 109898 540986 110134
rect 541222 109898 541404 110134
rect 540804 74454 541404 109898
rect 540804 74218 540986 74454
rect 541222 74218 541404 74454
rect 540804 74134 541404 74218
rect 540804 73898 540986 74134
rect 541222 73898 541404 74134
rect 540804 38454 541404 73898
rect 540804 38218 540986 38454
rect 541222 38218 541404 38454
rect 540804 38134 541404 38218
rect 540804 37898 540986 38134
rect 541222 37898 541404 38134
rect 540804 2454 541404 37898
rect 540804 2218 540986 2454
rect 541222 2218 541404 2454
rect 540804 2134 541404 2218
rect 540804 1898 540986 2134
rect 541222 1898 541404 2134
rect 540804 -346 541404 1898
rect 540804 -582 540986 -346
rect 541222 -582 541404 -346
rect 540804 -666 541404 -582
rect 540804 -902 540986 -666
rect 541222 -902 541404 -666
rect 540804 -1864 541404 -902
rect 544404 690054 545004 706162
rect 544404 689818 544586 690054
rect 544822 689818 545004 690054
rect 544404 689734 545004 689818
rect 544404 689498 544586 689734
rect 544822 689498 545004 689734
rect 544404 654054 545004 689498
rect 544404 653818 544586 654054
rect 544822 653818 545004 654054
rect 544404 653734 545004 653818
rect 544404 653498 544586 653734
rect 544822 653498 545004 653734
rect 544404 618054 545004 653498
rect 544404 617818 544586 618054
rect 544822 617818 545004 618054
rect 544404 617734 545004 617818
rect 544404 617498 544586 617734
rect 544822 617498 545004 617734
rect 544404 582054 545004 617498
rect 544404 581818 544586 582054
rect 544822 581818 545004 582054
rect 544404 581734 545004 581818
rect 544404 581498 544586 581734
rect 544822 581498 545004 581734
rect 544404 546054 545004 581498
rect 544404 545818 544586 546054
rect 544822 545818 545004 546054
rect 544404 545734 545004 545818
rect 544404 545498 544586 545734
rect 544822 545498 545004 545734
rect 544404 510054 545004 545498
rect 544404 509818 544586 510054
rect 544822 509818 545004 510054
rect 544404 509734 545004 509818
rect 544404 509498 544586 509734
rect 544822 509498 545004 509734
rect 544404 474054 545004 509498
rect 544404 473818 544586 474054
rect 544822 473818 545004 474054
rect 544404 473734 545004 473818
rect 544404 473498 544586 473734
rect 544822 473498 545004 473734
rect 544404 438054 545004 473498
rect 544404 437818 544586 438054
rect 544822 437818 545004 438054
rect 544404 437734 545004 437818
rect 544404 437498 544586 437734
rect 544822 437498 545004 437734
rect 544404 402054 545004 437498
rect 544404 401818 544586 402054
rect 544822 401818 545004 402054
rect 544404 401734 545004 401818
rect 544404 401498 544586 401734
rect 544822 401498 545004 401734
rect 544404 366054 545004 401498
rect 544404 365818 544586 366054
rect 544822 365818 545004 366054
rect 544404 365734 545004 365818
rect 544404 365498 544586 365734
rect 544822 365498 545004 365734
rect 544404 330054 545004 365498
rect 544404 329818 544586 330054
rect 544822 329818 545004 330054
rect 544404 329734 545004 329818
rect 544404 329498 544586 329734
rect 544822 329498 545004 329734
rect 544404 294054 545004 329498
rect 544404 293818 544586 294054
rect 544822 293818 545004 294054
rect 544404 293734 545004 293818
rect 544404 293498 544586 293734
rect 544822 293498 545004 293734
rect 544404 258054 545004 293498
rect 544404 257818 544586 258054
rect 544822 257818 545004 258054
rect 544404 257734 545004 257818
rect 544404 257498 544586 257734
rect 544822 257498 545004 257734
rect 544404 222054 545004 257498
rect 544404 221818 544586 222054
rect 544822 221818 545004 222054
rect 544404 221734 545004 221818
rect 544404 221498 544586 221734
rect 544822 221498 545004 221734
rect 544404 186054 545004 221498
rect 544404 185818 544586 186054
rect 544822 185818 545004 186054
rect 544404 185734 545004 185818
rect 544404 185498 544586 185734
rect 544822 185498 545004 185734
rect 544404 150054 545004 185498
rect 544404 149818 544586 150054
rect 544822 149818 545004 150054
rect 544404 149734 545004 149818
rect 544404 149498 544586 149734
rect 544822 149498 545004 149734
rect 544404 114054 545004 149498
rect 544404 113818 544586 114054
rect 544822 113818 545004 114054
rect 544404 113734 545004 113818
rect 544404 113498 544586 113734
rect 544822 113498 545004 113734
rect 544404 78054 545004 113498
rect 544404 77818 544586 78054
rect 544822 77818 545004 78054
rect 544404 77734 545004 77818
rect 544404 77498 544586 77734
rect 544822 77498 545004 77734
rect 544404 42054 545004 77498
rect 544404 41818 544586 42054
rect 544822 41818 545004 42054
rect 544404 41734 545004 41818
rect 544404 41498 544586 41734
rect 544822 41498 545004 41734
rect 544404 6054 545004 41498
rect 544404 5818 544586 6054
rect 544822 5818 545004 6054
rect 544404 5734 545004 5818
rect 544404 5498 544586 5734
rect 544822 5498 545004 5734
rect 544404 -2226 545004 5498
rect 544404 -2462 544586 -2226
rect 544822 -2462 545004 -2226
rect 544404 -2546 545004 -2462
rect 544404 -2782 544586 -2546
rect 544822 -2782 545004 -2546
rect 544404 -3744 545004 -2782
rect 548004 693654 548604 708042
rect 550587 697372 550653 697373
rect 550587 697308 550588 697372
rect 550652 697308 550653 697372
rect 550587 697307 550653 697308
rect 550590 696965 550650 697307
rect 551604 697254 552204 709922
rect 569604 711418 570204 711440
rect 569604 711182 569786 711418
rect 570022 711182 570204 711418
rect 569604 711098 570204 711182
rect 569604 710862 569786 711098
rect 570022 710862 570204 711098
rect 566004 709538 566604 709560
rect 566004 709302 566186 709538
rect 566422 709302 566604 709538
rect 566004 709218 566604 709302
rect 566004 708982 566186 709218
rect 566422 708982 566604 709218
rect 562404 707658 563004 707680
rect 562404 707422 562586 707658
rect 562822 707422 563004 707658
rect 562404 707338 563004 707422
rect 562404 707102 562586 707338
rect 562822 707102 563004 707338
rect 551604 697018 551786 697254
rect 552022 697018 552204 697254
rect 550587 696964 550653 696965
rect 550587 696900 550588 696964
rect 550652 696900 550653 696964
rect 550587 696899 550653 696900
rect 551604 696934 552204 697018
rect 548004 693418 548186 693654
rect 548422 693418 548604 693654
rect 548004 693334 548604 693418
rect 548004 693098 548186 693334
rect 548422 693098 548604 693334
rect 548004 657654 548604 693098
rect 551604 696698 551786 696934
rect 552022 696698 552204 696934
rect 550587 686356 550653 686357
rect 550587 686292 550588 686356
rect 550652 686292 550653 686356
rect 550587 686291 550653 686292
rect 550590 685949 550650 686291
rect 550587 685948 550653 685949
rect 550587 685884 550588 685948
rect 550652 685884 550653 685948
rect 550587 685883 550653 685884
rect 548004 657418 548186 657654
rect 548422 657418 548604 657654
rect 548004 657334 548604 657418
rect 548004 657098 548186 657334
rect 548422 657098 548604 657334
rect 548004 621654 548604 657098
rect 548004 621418 548186 621654
rect 548422 621418 548604 621654
rect 548004 621334 548604 621418
rect 548004 621098 548186 621334
rect 548422 621098 548604 621334
rect 548004 585654 548604 621098
rect 548004 585418 548186 585654
rect 548422 585418 548604 585654
rect 548004 585334 548604 585418
rect 548004 585098 548186 585334
rect 548422 585098 548604 585334
rect 548004 549654 548604 585098
rect 548004 549418 548186 549654
rect 548422 549418 548604 549654
rect 548004 549334 548604 549418
rect 548004 549098 548186 549334
rect 548422 549098 548604 549334
rect 548004 513654 548604 549098
rect 551604 661254 552204 696698
rect 551604 661018 551786 661254
rect 552022 661018 552204 661254
rect 551604 660934 552204 661018
rect 551604 660698 551786 660934
rect 552022 660698 552204 660934
rect 551604 625254 552204 660698
rect 551604 625018 551786 625254
rect 552022 625018 552204 625254
rect 551604 624934 552204 625018
rect 551604 624698 551786 624934
rect 552022 624698 552204 624934
rect 551604 589254 552204 624698
rect 551604 589018 551786 589254
rect 552022 589018 552204 589254
rect 551604 588934 552204 589018
rect 551604 588698 551786 588934
rect 552022 588698 552204 588934
rect 551604 553254 552204 588698
rect 551604 553018 551786 553254
rect 552022 553018 552204 553254
rect 551604 552934 552204 553018
rect 551604 552698 551786 552934
rect 552022 552698 552204 552934
rect 550587 545596 550653 545597
rect 550587 545532 550588 545596
rect 550652 545532 550653 545596
rect 550587 545531 550653 545532
rect 550590 545189 550650 545531
rect 550587 545188 550653 545189
rect 550587 545124 550588 545188
rect 550652 545124 550653 545188
rect 550587 545123 550653 545124
rect 548004 513418 548186 513654
rect 548422 513418 548604 513654
rect 548004 513334 548604 513418
rect 548004 513098 548186 513334
rect 548422 513098 548604 513334
rect 548004 477654 548604 513098
rect 548004 477418 548186 477654
rect 548422 477418 548604 477654
rect 548004 477334 548604 477418
rect 548004 477098 548186 477334
rect 548422 477098 548604 477334
rect 548004 441654 548604 477098
rect 548004 441418 548186 441654
rect 548422 441418 548604 441654
rect 548004 441334 548604 441418
rect 548004 441098 548186 441334
rect 548422 441098 548604 441334
rect 548004 405654 548604 441098
rect 548004 405418 548186 405654
rect 548422 405418 548604 405654
rect 548004 405334 548604 405418
rect 548004 405098 548186 405334
rect 548422 405098 548604 405334
rect 548004 369654 548604 405098
rect 548004 369418 548186 369654
rect 548422 369418 548604 369654
rect 548004 369334 548604 369418
rect 548004 369098 548186 369334
rect 548422 369098 548604 369334
rect 548004 333654 548604 369098
rect 548004 333418 548186 333654
rect 548422 333418 548604 333654
rect 548004 333334 548604 333418
rect 548004 333098 548186 333334
rect 548422 333098 548604 333334
rect 548004 297654 548604 333098
rect 548004 297418 548186 297654
rect 548422 297418 548604 297654
rect 548004 297334 548604 297418
rect 548004 297098 548186 297334
rect 548422 297098 548604 297334
rect 548004 261654 548604 297098
rect 548004 261418 548186 261654
rect 548422 261418 548604 261654
rect 548004 261334 548604 261418
rect 548004 261098 548186 261334
rect 548422 261098 548604 261334
rect 548004 225654 548604 261098
rect 548004 225418 548186 225654
rect 548422 225418 548604 225654
rect 548004 225334 548604 225418
rect 548004 225098 548186 225334
rect 548422 225098 548604 225334
rect 548004 189654 548604 225098
rect 548004 189418 548186 189654
rect 548422 189418 548604 189654
rect 548004 189334 548604 189418
rect 548004 189098 548186 189334
rect 548422 189098 548604 189334
rect 548004 153654 548604 189098
rect 548004 153418 548186 153654
rect 548422 153418 548604 153654
rect 548004 153334 548604 153418
rect 548004 153098 548186 153334
rect 548422 153098 548604 153334
rect 548004 117654 548604 153098
rect 548004 117418 548186 117654
rect 548422 117418 548604 117654
rect 548004 117334 548604 117418
rect 548004 117098 548186 117334
rect 548422 117098 548604 117334
rect 548004 81654 548604 117098
rect 548004 81418 548186 81654
rect 548422 81418 548604 81654
rect 548004 81334 548604 81418
rect 548004 81098 548186 81334
rect 548422 81098 548604 81334
rect 548004 45654 548604 81098
rect 548004 45418 548186 45654
rect 548422 45418 548604 45654
rect 548004 45334 548604 45418
rect 548004 45098 548186 45334
rect 548422 45098 548604 45334
rect 548004 9654 548604 45098
rect 548004 9418 548186 9654
rect 548422 9418 548604 9654
rect 548004 9334 548604 9418
rect 548004 9098 548186 9334
rect 548422 9098 548604 9334
rect 548004 -4106 548604 9098
rect 548004 -4342 548186 -4106
rect 548422 -4342 548604 -4106
rect 548004 -4426 548604 -4342
rect 548004 -4662 548186 -4426
rect 548422 -4662 548604 -4426
rect 548004 -5624 548604 -4662
rect 551604 517254 552204 552698
rect 551604 517018 551786 517254
rect 552022 517018 552204 517254
rect 551604 516934 552204 517018
rect 551604 516698 551786 516934
rect 552022 516698 552204 516934
rect 551604 481254 552204 516698
rect 551604 481018 551786 481254
rect 552022 481018 552204 481254
rect 551604 480934 552204 481018
rect 551604 480698 551786 480934
rect 552022 480698 552204 480934
rect 551604 445254 552204 480698
rect 551604 445018 551786 445254
rect 552022 445018 552204 445254
rect 551604 444934 552204 445018
rect 551604 444698 551786 444934
rect 552022 444698 552204 444934
rect 551604 409254 552204 444698
rect 551604 409018 551786 409254
rect 552022 409018 552204 409254
rect 551604 408934 552204 409018
rect 551604 408698 551786 408934
rect 552022 408698 552204 408934
rect 551604 373254 552204 408698
rect 551604 373018 551786 373254
rect 552022 373018 552204 373254
rect 551604 372934 552204 373018
rect 551604 372698 551786 372934
rect 552022 372698 552204 372934
rect 551604 337254 552204 372698
rect 551604 337018 551786 337254
rect 552022 337018 552204 337254
rect 551604 336934 552204 337018
rect 551604 336698 551786 336934
rect 552022 336698 552204 336934
rect 551604 301254 552204 336698
rect 551604 301018 551786 301254
rect 552022 301018 552204 301254
rect 551604 300934 552204 301018
rect 551604 300698 551786 300934
rect 552022 300698 552204 300934
rect 551604 265254 552204 300698
rect 551604 265018 551786 265254
rect 552022 265018 552204 265254
rect 551604 264934 552204 265018
rect 551604 264698 551786 264934
rect 552022 264698 552204 264934
rect 551604 229254 552204 264698
rect 551604 229018 551786 229254
rect 552022 229018 552204 229254
rect 551604 228934 552204 229018
rect 551604 228698 551786 228934
rect 552022 228698 552204 228934
rect 551604 193254 552204 228698
rect 551604 193018 551786 193254
rect 552022 193018 552204 193254
rect 551604 192934 552204 193018
rect 551604 192698 551786 192934
rect 552022 192698 552204 192934
rect 551604 157254 552204 192698
rect 551604 157018 551786 157254
rect 552022 157018 552204 157254
rect 551604 156934 552204 157018
rect 551604 156698 551786 156934
rect 552022 156698 552204 156934
rect 551604 121254 552204 156698
rect 551604 121018 551786 121254
rect 552022 121018 552204 121254
rect 551604 120934 552204 121018
rect 551604 120698 551786 120934
rect 552022 120698 552204 120934
rect 551604 85254 552204 120698
rect 551604 85018 551786 85254
rect 552022 85018 552204 85254
rect 551604 84934 552204 85018
rect 551604 84698 551786 84934
rect 552022 84698 552204 84934
rect 551604 49254 552204 84698
rect 551604 49018 551786 49254
rect 552022 49018 552204 49254
rect 551604 48934 552204 49018
rect 551604 48698 551786 48934
rect 552022 48698 552204 48934
rect 551604 13254 552204 48698
rect 551604 13018 551786 13254
rect 552022 13018 552204 13254
rect 551604 12934 552204 13018
rect 551604 12698 551786 12934
rect 552022 12698 552204 12934
rect 533604 -7162 533786 -6926
rect 534022 -7162 534204 -6926
rect 533604 -7246 534204 -7162
rect 533604 -7482 533786 -7246
rect 534022 -7482 534204 -7246
rect 533604 -7504 534204 -7482
rect 551604 -5986 552204 12698
rect 558804 705778 559404 705800
rect 558804 705542 558986 705778
rect 559222 705542 559404 705778
rect 558804 705458 559404 705542
rect 558804 705222 558986 705458
rect 559222 705222 559404 705458
rect 558804 668454 559404 705222
rect 558804 668218 558986 668454
rect 559222 668218 559404 668454
rect 558804 668134 559404 668218
rect 558804 667898 558986 668134
rect 559222 667898 559404 668134
rect 558804 632454 559404 667898
rect 558804 632218 558986 632454
rect 559222 632218 559404 632454
rect 558804 632134 559404 632218
rect 558804 631898 558986 632134
rect 559222 631898 559404 632134
rect 558804 596454 559404 631898
rect 558804 596218 558986 596454
rect 559222 596218 559404 596454
rect 558804 596134 559404 596218
rect 558804 595898 558986 596134
rect 559222 595898 559404 596134
rect 558804 560454 559404 595898
rect 558804 560218 558986 560454
rect 559222 560218 559404 560454
rect 558804 560134 559404 560218
rect 558804 559898 558986 560134
rect 559222 559898 559404 560134
rect 558804 524454 559404 559898
rect 558804 524218 558986 524454
rect 559222 524218 559404 524454
rect 558804 524134 559404 524218
rect 558804 523898 558986 524134
rect 559222 523898 559404 524134
rect 558804 488454 559404 523898
rect 558804 488218 558986 488454
rect 559222 488218 559404 488454
rect 558804 488134 559404 488218
rect 558804 487898 558986 488134
rect 559222 487898 559404 488134
rect 558804 452454 559404 487898
rect 558804 452218 558986 452454
rect 559222 452218 559404 452454
rect 558804 452134 559404 452218
rect 558804 451898 558986 452134
rect 559222 451898 559404 452134
rect 558804 416454 559404 451898
rect 558804 416218 558986 416454
rect 559222 416218 559404 416454
rect 558804 416134 559404 416218
rect 558804 415898 558986 416134
rect 559222 415898 559404 416134
rect 558804 380454 559404 415898
rect 558804 380218 558986 380454
rect 559222 380218 559404 380454
rect 558804 380134 559404 380218
rect 558804 379898 558986 380134
rect 559222 379898 559404 380134
rect 558804 344454 559404 379898
rect 558804 344218 558986 344454
rect 559222 344218 559404 344454
rect 558804 344134 559404 344218
rect 558804 343898 558986 344134
rect 559222 343898 559404 344134
rect 558804 308454 559404 343898
rect 558804 308218 558986 308454
rect 559222 308218 559404 308454
rect 558804 308134 559404 308218
rect 558804 307898 558986 308134
rect 559222 307898 559404 308134
rect 558804 272454 559404 307898
rect 558804 272218 558986 272454
rect 559222 272218 559404 272454
rect 558804 272134 559404 272218
rect 558804 271898 558986 272134
rect 559222 271898 559404 272134
rect 558804 236454 559404 271898
rect 558804 236218 558986 236454
rect 559222 236218 559404 236454
rect 558804 236134 559404 236218
rect 558804 235898 558986 236134
rect 559222 235898 559404 236134
rect 558804 200454 559404 235898
rect 558804 200218 558986 200454
rect 559222 200218 559404 200454
rect 558804 200134 559404 200218
rect 558804 199898 558986 200134
rect 559222 199898 559404 200134
rect 558804 164454 559404 199898
rect 558804 164218 558986 164454
rect 559222 164218 559404 164454
rect 558804 164134 559404 164218
rect 558804 163898 558986 164134
rect 559222 163898 559404 164134
rect 558804 128454 559404 163898
rect 558804 128218 558986 128454
rect 559222 128218 559404 128454
rect 558804 128134 559404 128218
rect 558804 127898 558986 128134
rect 559222 127898 559404 128134
rect 558804 92454 559404 127898
rect 558804 92218 558986 92454
rect 559222 92218 559404 92454
rect 558804 92134 559404 92218
rect 558804 91898 558986 92134
rect 559222 91898 559404 92134
rect 558804 56454 559404 91898
rect 558804 56218 558986 56454
rect 559222 56218 559404 56454
rect 558804 56134 559404 56218
rect 558804 55898 558986 56134
rect 559222 55898 559404 56134
rect 558804 20454 559404 55898
rect 558804 20218 558986 20454
rect 559222 20218 559404 20454
rect 558804 20134 559404 20218
rect 558804 19898 558986 20134
rect 559222 19898 559404 20134
rect 558804 -1286 559404 19898
rect 558804 -1522 558986 -1286
rect 559222 -1522 559404 -1286
rect 558804 -1606 559404 -1522
rect 558804 -1842 558986 -1606
rect 559222 -1842 559404 -1606
rect 558804 -1864 559404 -1842
rect 562404 672054 563004 707102
rect 562404 671818 562586 672054
rect 562822 671818 563004 672054
rect 562404 671734 563004 671818
rect 562404 671498 562586 671734
rect 562822 671498 563004 671734
rect 562404 636054 563004 671498
rect 562404 635818 562586 636054
rect 562822 635818 563004 636054
rect 562404 635734 563004 635818
rect 562404 635498 562586 635734
rect 562822 635498 563004 635734
rect 562404 600054 563004 635498
rect 562404 599818 562586 600054
rect 562822 599818 563004 600054
rect 562404 599734 563004 599818
rect 562404 599498 562586 599734
rect 562822 599498 563004 599734
rect 562404 564054 563004 599498
rect 562404 563818 562586 564054
rect 562822 563818 563004 564054
rect 562404 563734 563004 563818
rect 562404 563498 562586 563734
rect 562822 563498 563004 563734
rect 562404 528054 563004 563498
rect 562404 527818 562586 528054
rect 562822 527818 563004 528054
rect 562404 527734 563004 527818
rect 562404 527498 562586 527734
rect 562822 527498 563004 527734
rect 562404 492054 563004 527498
rect 562404 491818 562586 492054
rect 562822 491818 563004 492054
rect 562404 491734 563004 491818
rect 562404 491498 562586 491734
rect 562822 491498 563004 491734
rect 562404 456054 563004 491498
rect 562404 455818 562586 456054
rect 562822 455818 563004 456054
rect 562404 455734 563004 455818
rect 562404 455498 562586 455734
rect 562822 455498 563004 455734
rect 562404 420054 563004 455498
rect 562404 419818 562586 420054
rect 562822 419818 563004 420054
rect 562404 419734 563004 419818
rect 562404 419498 562586 419734
rect 562822 419498 563004 419734
rect 562404 384054 563004 419498
rect 562404 383818 562586 384054
rect 562822 383818 563004 384054
rect 562404 383734 563004 383818
rect 562404 383498 562586 383734
rect 562822 383498 563004 383734
rect 562404 348054 563004 383498
rect 562404 347818 562586 348054
rect 562822 347818 563004 348054
rect 562404 347734 563004 347818
rect 562404 347498 562586 347734
rect 562822 347498 563004 347734
rect 562404 312054 563004 347498
rect 562404 311818 562586 312054
rect 562822 311818 563004 312054
rect 562404 311734 563004 311818
rect 562404 311498 562586 311734
rect 562822 311498 563004 311734
rect 562404 276054 563004 311498
rect 562404 275818 562586 276054
rect 562822 275818 563004 276054
rect 562404 275734 563004 275818
rect 562404 275498 562586 275734
rect 562822 275498 563004 275734
rect 562404 240054 563004 275498
rect 562404 239818 562586 240054
rect 562822 239818 563004 240054
rect 562404 239734 563004 239818
rect 562404 239498 562586 239734
rect 562822 239498 563004 239734
rect 562404 204054 563004 239498
rect 562404 203818 562586 204054
rect 562822 203818 563004 204054
rect 562404 203734 563004 203818
rect 562404 203498 562586 203734
rect 562822 203498 563004 203734
rect 562404 168054 563004 203498
rect 562404 167818 562586 168054
rect 562822 167818 563004 168054
rect 562404 167734 563004 167818
rect 562404 167498 562586 167734
rect 562822 167498 563004 167734
rect 562404 132054 563004 167498
rect 562404 131818 562586 132054
rect 562822 131818 563004 132054
rect 562404 131734 563004 131818
rect 562404 131498 562586 131734
rect 562822 131498 563004 131734
rect 562404 96054 563004 131498
rect 562404 95818 562586 96054
rect 562822 95818 563004 96054
rect 562404 95734 563004 95818
rect 562404 95498 562586 95734
rect 562822 95498 563004 95734
rect 562404 60054 563004 95498
rect 562404 59818 562586 60054
rect 562822 59818 563004 60054
rect 562404 59734 563004 59818
rect 562404 59498 562586 59734
rect 562822 59498 563004 59734
rect 562404 24054 563004 59498
rect 562404 23818 562586 24054
rect 562822 23818 563004 24054
rect 562404 23734 563004 23818
rect 562404 23498 562586 23734
rect 562822 23498 563004 23734
rect 562404 -3166 563004 23498
rect 562404 -3402 562586 -3166
rect 562822 -3402 563004 -3166
rect 562404 -3486 563004 -3402
rect 562404 -3722 562586 -3486
rect 562822 -3722 563004 -3486
rect 562404 -3744 563004 -3722
rect 566004 675654 566604 708982
rect 566004 675418 566186 675654
rect 566422 675418 566604 675654
rect 566004 675334 566604 675418
rect 566004 675098 566186 675334
rect 566422 675098 566604 675334
rect 566004 639654 566604 675098
rect 566004 639418 566186 639654
rect 566422 639418 566604 639654
rect 566004 639334 566604 639418
rect 566004 639098 566186 639334
rect 566422 639098 566604 639334
rect 566004 603654 566604 639098
rect 566004 603418 566186 603654
rect 566422 603418 566604 603654
rect 566004 603334 566604 603418
rect 566004 603098 566186 603334
rect 566422 603098 566604 603334
rect 566004 567654 566604 603098
rect 566004 567418 566186 567654
rect 566422 567418 566604 567654
rect 566004 567334 566604 567418
rect 566004 567098 566186 567334
rect 566422 567098 566604 567334
rect 566004 531654 566604 567098
rect 566004 531418 566186 531654
rect 566422 531418 566604 531654
rect 566004 531334 566604 531418
rect 566004 531098 566186 531334
rect 566422 531098 566604 531334
rect 566004 495654 566604 531098
rect 566004 495418 566186 495654
rect 566422 495418 566604 495654
rect 566004 495334 566604 495418
rect 566004 495098 566186 495334
rect 566422 495098 566604 495334
rect 566004 459654 566604 495098
rect 566004 459418 566186 459654
rect 566422 459418 566604 459654
rect 566004 459334 566604 459418
rect 566004 459098 566186 459334
rect 566422 459098 566604 459334
rect 566004 423654 566604 459098
rect 566004 423418 566186 423654
rect 566422 423418 566604 423654
rect 566004 423334 566604 423418
rect 566004 423098 566186 423334
rect 566422 423098 566604 423334
rect 566004 387654 566604 423098
rect 566004 387418 566186 387654
rect 566422 387418 566604 387654
rect 566004 387334 566604 387418
rect 566004 387098 566186 387334
rect 566422 387098 566604 387334
rect 566004 351654 566604 387098
rect 566004 351418 566186 351654
rect 566422 351418 566604 351654
rect 566004 351334 566604 351418
rect 566004 351098 566186 351334
rect 566422 351098 566604 351334
rect 566004 315654 566604 351098
rect 566004 315418 566186 315654
rect 566422 315418 566604 315654
rect 566004 315334 566604 315418
rect 566004 315098 566186 315334
rect 566422 315098 566604 315334
rect 566004 279654 566604 315098
rect 566004 279418 566186 279654
rect 566422 279418 566604 279654
rect 566004 279334 566604 279418
rect 566004 279098 566186 279334
rect 566422 279098 566604 279334
rect 566004 243654 566604 279098
rect 566004 243418 566186 243654
rect 566422 243418 566604 243654
rect 566004 243334 566604 243418
rect 566004 243098 566186 243334
rect 566422 243098 566604 243334
rect 566004 207654 566604 243098
rect 566004 207418 566186 207654
rect 566422 207418 566604 207654
rect 566004 207334 566604 207418
rect 566004 207098 566186 207334
rect 566422 207098 566604 207334
rect 566004 171654 566604 207098
rect 566004 171418 566186 171654
rect 566422 171418 566604 171654
rect 566004 171334 566604 171418
rect 566004 171098 566186 171334
rect 566422 171098 566604 171334
rect 566004 135654 566604 171098
rect 566004 135418 566186 135654
rect 566422 135418 566604 135654
rect 566004 135334 566604 135418
rect 566004 135098 566186 135334
rect 566422 135098 566604 135334
rect 566004 99654 566604 135098
rect 566004 99418 566186 99654
rect 566422 99418 566604 99654
rect 566004 99334 566604 99418
rect 566004 99098 566186 99334
rect 566422 99098 566604 99334
rect 566004 63654 566604 99098
rect 566004 63418 566186 63654
rect 566422 63418 566604 63654
rect 566004 63334 566604 63418
rect 566004 63098 566186 63334
rect 566422 63098 566604 63334
rect 566004 27654 566604 63098
rect 566004 27418 566186 27654
rect 566422 27418 566604 27654
rect 566004 27334 566604 27418
rect 566004 27098 566186 27334
rect 566422 27098 566604 27334
rect 566004 -5046 566604 27098
rect 566004 -5282 566186 -5046
rect 566422 -5282 566604 -5046
rect 566004 -5366 566604 -5282
rect 566004 -5602 566186 -5366
rect 566422 -5602 566604 -5366
rect 566004 -5624 566604 -5602
rect 569604 679254 570204 710862
rect 591900 711418 592500 711440
rect 591900 711182 592082 711418
rect 592318 711182 592500 711418
rect 591900 711098 592500 711182
rect 591900 710862 592082 711098
rect 592318 710862 592500 711098
rect 590960 710478 591560 710500
rect 590960 710242 591142 710478
rect 591378 710242 591560 710478
rect 590960 710158 591560 710242
rect 590960 709922 591142 710158
rect 591378 709922 591560 710158
rect 590020 709538 590620 709560
rect 590020 709302 590202 709538
rect 590438 709302 590620 709538
rect 590020 709218 590620 709302
rect 590020 708982 590202 709218
rect 590438 708982 590620 709218
rect 589080 708598 589680 708620
rect 589080 708362 589262 708598
rect 589498 708362 589680 708598
rect 589080 708278 589680 708362
rect 589080 708042 589262 708278
rect 589498 708042 589680 708278
rect 580404 706718 581004 707680
rect 588140 707658 588740 707680
rect 588140 707422 588322 707658
rect 588558 707422 588740 707658
rect 588140 707338 588740 707422
rect 588140 707102 588322 707338
rect 588558 707102 588740 707338
rect 580404 706482 580586 706718
rect 580822 706482 581004 706718
rect 580404 706398 581004 706482
rect 580404 706162 580586 706398
rect 580822 706162 581004 706398
rect 569604 679018 569786 679254
rect 570022 679018 570204 679254
rect 569604 678934 570204 679018
rect 569604 678698 569786 678934
rect 570022 678698 570204 678934
rect 569604 643254 570204 678698
rect 569604 643018 569786 643254
rect 570022 643018 570204 643254
rect 569604 642934 570204 643018
rect 569604 642698 569786 642934
rect 570022 642698 570204 642934
rect 569604 607254 570204 642698
rect 569604 607018 569786 607254
rect 570022 607018 570204 607254
rect 569604 606934 570204 607018
rect 569604 606698 569786 606934
rect 570022 606698 570204 606934
rect 569604 571254 570204 606698
rect 569604 571018 569786 571254
rect 570022 571018 570204 571254
rect 569604 570934 570204 571018
rect 569604 570698 569786 570934
rect 570022 570698 570204 570934
rect 569604 535254 570204 570698
rect 569604 535018 569786 535254
rect 570022 535018 570204 535254
rect 569604 534934 570204 535018
rect 569604 534698 569786 534934
rect 570022 534698 570204 534934
rect 569604 499254 570204 534698
rect 569604 499018 569786 499254
rect 570022 499018 570204 499254
rect 569604 498934 570204 499018
rect 569604 498698 569786 498934
rect 570022 498698 570204 498934
rect 569604 463254 570204 498698
rect 569604 463018 569786 463254
rect 570022 463018 570204 463254
rect 569604 462934 570204 463018
rect 569604 462698 569786 462934
rect 570022 462698 570204 462934
rect 569604 427254 570204 462698
rect 569604 427018 569786 427254
rect 570022 427018 570204 427254
rect 569604 426934 570204 427018
rect 569604 426698 569786 426934
rect 570022 426698 570204 426934
rect 569604 391254 570204 426698
rect 569604 391018 569786 391254
rect 570022 391018 570204 391254
rect 569604 390934 570204 391018
rect 569604 390698 569786 390934
rect 570022 390698 570204 390934
rect 569604 355254 570204 390698
rect 569604 355018 569786 355254
rect 570022 355018 570204 355254
rect 569604 354934 570204 355018
rect 569604 354698 569786 354934
rect 570022 354698 570204 354934
rect 569604 319254 570204 354698
rect 569604 319018 569786 319254
rect 570022 319018 570204 319254
rect 569604 318934 570204 319018
rect 569604 318698 569786 318934
rect 570022 318698 570204 318934
rect 569604 283254 570204 318698
rect 569604 283018 569786 283254
rect 570022 283018 570204 283254
rect 569604 282934 570204 283018
rect 569604 282698 569786 282934
rect 570022 282698 570204 282934
rect 569604 247254 570204 282698
rect 569604 247018 569786 247254
rect 570022 247018 570204 247254
rect 569604 246934 570204 247018
rect 569604 246698 569786 246934
rect 570022 246698 570204 246934
rect 569604 211254 570204 246698
rect 569604 211018 569786 211254
rect 570022 211018 570204 211254
rect 569604 210934 570204 211018
rect 569604 210698 569786 210934
rect 570022 210698 570204 210934
rect 569604 175254 570204 210698
rect 569604 175018 569786 175254
rect 570022 175018 570204 175254
rect 569604 174934 570204 175018
rect 569604 174698 569786 174934
rect 570022 174698 570204 174934
rect 569604 139254 570204 174698
rect 569604 139018 569786 139254
rect 570022 139018 570204 139254
rect 569604 138934 570204 139018
rect 569604 138698 569786 138934
rect 570022 138698 570204 138934
rect 569604 103254 570204 138698
rect 569604 103018 569786 103254
rect 570022 103018 570204 103254
rect 569604 102934 570204 103018
rect 569604 102698 569786 102934
rect 570022 102698 570204 102934
rect 569604 67254 570204 102698
rect 569604 67018 569786 67254
rect 570022 67018 570204 67254
rect 569604 66934 570204 67018
rect 569604 66698 569786 66934
rect 570022 66698 570204 66934
rect 569604 31254 570204 66698
rect 569604 31018 569786 31254
rect 570022 31018 570204 31254
rect 569604 30934 570204 31018
rect 569604 30698 569786 30934
rect 570022 30698 570204 30934
rect 551604 -6222 551786 -5986
rect 552022 -6222 552204 -5986
rect 551604 -6306 552204 -6222
rect 551604 -6542 551786 -6306
rect 552022 -6542 552204 -6306
rect 551604 -7504 552204 -6542
rect 569604 -6926 570204 30698
rect 576804 704838 577404 705800
rect 576804 704602 576986 704838
rect 577222 704602 577404 704838
rect 576804 704518 577404 704602
rect 576804 704282 576986 704518
rect 577222 704282 577404 704518
rect 576804 686454 577404 704282
rect 576804 686218 576986 686454
rect 577222 686218 577404 686454
rect 576804 686134 577404 686218
rect 576804 685898 576986 686134
rect 577222 685898 577404 686134
rect 576804 650454 577404 685898
rect 580404 690054 581004 706162
rect 587200 706718 587800 706740
rect 587200 706482 587382 706718
rect 587618 706482 587800 706718
rect 587200 706398 587800 706482
rect 587200 706162 587382 706398
rect 587618 706162 587800 706398
rect 586260 705778 586860 705800
rect 586260 705542 586442 705778
rect 586678 705542 586860 705778
rect 586260 705458 586860 705542
rect 586260 705222 586442 705458
rect 586678 705222 586860 705458
rect 580404 689818 580586 690054
rect 580822 689818 581004 690054
rect 580404 689734 581004 689818
rect 580404 689498 580586 689734
rect 580822 689498 581004 689734
rect 580404 654054 581004 689498
rect 580404 653818 580586 654054
rect 580822 653818 581004 654054
rect 580404 653734 581004 653818
rect 580404 653498 580586 653734
rect 580822 653498 581004 653734
rect 579659 650860 579725 650861
rect 579659 650796 579660 650860
rect 579724 650796 579725 650860
rect 579659 650795 579725 650796
rect 579662 650589 579722 650795
rect 579659 650588 579725 650589
rect 579659 650524 579660 650588
rect 579724 650524 579725 650588
rect 579659 650523 579725 650524
rect 576804 650218 576986 650454
rect 577222 650218 577404 650454
rect 576804 650134 577404 650218
rect 576804 649898 576986 650134
rect 577222 649898 577404 650134
rect 576804 614454 577404 649898
rect 576804 614218 576986 614454
rect 577222 614218 577404 614454
rect 576804 614134 577404 614218
rect 576804 613898 576986 614134
rect 577222 613898 577404 614134
rect 576804 578454 577404 613898
rect 576804 578218 576986 578454
rect 577222 578218 577404 578454
rect 576804 578134 577404 578218
rect 576804 577898 576986 578134
rect 577222 577898 577404 578134
rect 576804 542454 577404 577898
rect 576804 542218 576986 542454
rect 577222 542218 577404 542454
rect 576804 542134 577404 542218
rect 576804 541898 576986 542134
rect 577222 541898 577404 542134
rect 576804 506454 577404 541898
rect 576804 506218 576986 506454
rect 577222 506218 577404 506454
rect 576804 506134 577404 506218
rect 576804 505898 576986 506134
rect 577222 505898 577404 506134
rect 576804 470454 577404 505898
rect 576804 470218 576986 470454
rect 577222 470218 577404 470454
rect 576804 470134 577404 470218
rect 576804 469898 576986 470134
rect 577222 469898 577404 470134
rect 576804 434454 577404 469898
rect 576804 434218 576986 434454
rect 577222 434218 577404 434454
rect 576804 434134 577404 434218
rect 576804 433898 576986 434134
rect 577222 433898 577404 434134
rect 576804 398454 577404 433898
rect 576804 398218 576986 398454
rect 577222 398218 577404 398454
rect 576804 398134 577404 398218
rect 576804 397898 576986 398134
rect 577222 397898 577404 398134
rect 576804 362454 577404 397898
rect 576804 362218 576986 362454
rect 577222 362218 577404 362454
rect 576804 362134 577404 362218
rect 576804 361898 576986 362134
rect 577222 361898 577404 362134
rect 576804 326454 577404 361898
rect 576804 326218 576986 326454
rect 577222 326218 577404 326454
rect 576804 326134 577404 326218
rect 576804 325898 576986 326134
rect 577222 325898 577404 326134
rect 576804 290454 577404 325898
rect 576804 290218 576986 290454
rect 577222 290218 577404 290454
rect 576804 290134 577404 290218
rect 576804 289898 576986 290134
rect 577222 289898 577404 290134
rect 576804 254454 577404 289898
rect 576804 254218 576986 254454
rect 577222 254218 577404 254454
rect 576804 254134 577404 254218
rect 576804 253898 576986 254134
rect 577222 253898 577404 254134
rect 576804 218454 577404 253898
rect 576804 218218 576986 218454
rect 577222 218218 577404 218454
rect 576804 218134 577404 218218
rect 576804 217898 576986 218134
rect 577222 217898 577404 218134
rect 576804 182454 577404 217898
rect 576804 182218 576986 182454
rect 577222 182218 577404 182454
rect 576804 182134 577404 182218
rect 576804 181898 576986 182134
rect 577222 181898 577404 182134
rect 576804 146454 577404 181898
rect 576804 146218 576986 146454
rect 577222 146218 577404 146454
rect 576804 146134 577404 146218
rect 576804 145898 576986 146134
rect 577222 145898 577404 146134
rect 576804 110454 577404 145898
rect 576804 110218 576986 110454
rect 577222 110218 577404 110454
rect 576804 110134 577404 110218
rect 576804 109898 576986 110134
rect 577222 109898 577404 110134
rect 576804 74454 577404 109898
rect 576804 74218 576986 74454
rect 577222 74218 577404 74454
rect 576804 74134 577404 74218
rect 576804 73898 576986 74134
rect 577222 73898 577404 74134
rect 576804 38454 577404 73898
rect 576804 38218 576986 38454
rect 577222 38218 577404 38454
rect 576804 38134 577404 38218
rect 576804 37898 576986 38134
rect 577222 37898 577404 38134
rect 576804 2454 577404 37898
rect 576804 2218 576986 2454
rect 577222 2218 577404 2454
rect 576804 2134 577404 2218
rect 576804 1898 576986 2134
rect 577222 1898 577404 2134
rect 576804 -346 577404 1898
rect 576804 -582 576986 -346
rect 577222 -582 577404 -346
rect 576804 -666 577404 -582
rect 576804 -902 576986 -666
rect 577222 -902 577404 -666
rect 576804 -1864 577404 -902
rect 580404 618054 581004 653498
rect 580404 617818 580586 618054
rect 580822 617818 581004 618054
rect 580404 617734 581004 617818
rect 580404 617498 580586 617734
rect 580822 617498 581004 617734
rect 580404 582054 581004 617498
rect 580404 581818 580586 582054
rect 580822 581818 581004 582054
rect 580404 581734 581004 581818
rect 580404 581498 580586 581734
rect 580822 581498 581004 581734
rect 580404 546054 581004 581498
rect 580404 545818 580586 546054
rect 580822 545818 581004 546054
rect 580404 545734 581004 545818
rect 580404 545498 580586 545734
rect 580822 545498 581004 545734
rect 580404 510054 581004 545498
rect 580404 509818 580586 510054
rect 580822 509818 581004 510054
rect 580404 509734 581004 509818
rect 580404 509498 580586 509734
rect 580822 509498 581004 509734
rect 580404 474054 581004 509498
rect 580404 473818 580586 474054
rect 580822 473818 581004 474054
rect 580404 473734 581004 473818
rect 580404 473498 580586 473734
rect 580822 473498 581004 473734
rect 580404 438054 581004 473498
rect 580404 437818 580586 438054
rect 580822 437818 581004 438054
rect 580404 437734 581004 437818
rect 580404 437498 580586 437734
rect 580822 437498 581004 437734
rect 580404 402054 581004 437498
rect 580404 401818 580586 402054
rect 580822 401818 581004 402054
rect 580404 401734 581004 401818
rect 580404 401498 580586 401734
rect 580822 401498 581004 401734
rect 580404 366054 581004 401498
rect 580404 365818 580586 366054
rect 580822 365818 581004 366054
rect 580404 365734 581004 365818
rect 580404 365498 580586 365734
rect 580822 365498 581004 365734
rect 580404 330054 581004 365498
rect 580404 329818 580586 330054
rect 580822 329818 581004 330054
rect 580404 329734 581004 329818
rect 580404 329498 580586 329734
rect 580822 329498 581004 329734
rect 580404 294054 581004 329498
rect 580404 293818 580586 294054
rect 580822 293818 581004 294054
rect 580404 293734 581004 293818
rect 580404 293498 580586 293734
rect 580822 293498 581004 293734
rect 580404 258054 581004 293498
rect 580404 257818 580586 258054
rect 580822 257818 581004 258054
rect 580404 257734 581004 257818
rect 580404 257498 580586 257734
rect 580822 257498 581004 257734
rect 580404 222054 581004 257498
rect 580404 221818 580586 222054
rect 580822 221818 581004 222054
rect 580404 221734 581004 221818
rect 580404 221498 580586 221734
rect 580822 221498 581004 221734
rect 580404 186054 581004 221498
rect 580404 185818 580586 186054
rect 580822 185818 581004 186054
rect 580404 185734 581004 185818
rect 580404 185498 580586 185734
rect 580822 185498 581004 185734
rect 580404 150054 581004 185498
rect 580404 149818 580586 150054
rect 580822 149818 581004 150054
rect 580404 149734 581004 149818
rect 580404 149498 580586 149734
rect 580822 149498 581004 149734
rect 580404 114054 581004 149498
rect 580404 113818 580586 114054
rect 580822 113818 581004 114054
rect 580404 113734 581004 113818
rect 580404 113498 580586 113734
rect 580822 113498 581004 113734
rect 580404 78054 581004 113498
rect 580404 77818 580586 78054
rect 580822 77818 581004 78054
rect 580404 77734 581004 77818
rect 580404 77498 580586 77734
rect 580822 77498 581004 77734
rect 580404 42054 581004 77498
rect 580404 41818 580586 42054
rect 580822 41818 581004 42054
rect 580404 41734 581004 41818
rect 580404 41498 580586 41734
rect 580822 41498 581004 41734
rect 580404 6054 581004 41498
rect 580404 5818 580586 6054
rect 580822 5818 581004 6054
rect 580404 5734 581004 5818
rect 580404 5498 580586 5734
rect 580822 5498 581004 5734
rect 580404 -2226 581004 5498
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 585320 686454 585920 704282
rect 585320 686218 585502 686454
rect 585738 686218 585920 686454
rect 585320 686134 585920 686218
rect 585320 685898 585502 686134
rect 585738 685898 585920 686134
rect 585320 650454 585920 685898
rect 585320 650218 585502 650454
rect 585738 650218 585920 650454
rect 585320 650134 585920 650218
rect 585320 649898 585502 650134
rect 585738 649898 585920 650134
rect 585320 614454 585920 649898
rect 585320 614218 585502 614454
rect 585738 614218 585920 614454
rect 585320 614134 585920 614218
rect 585320 613898 585502 614134
rect 585738 613898 585920 614134
rect 585320 578454 585920 613898
rect 585320 578218 585502 578454
rect 585738 578218 585920 578454
rect 585320 578134 585920 578218
rect 585320 577898 585502 578134
rect 585738 577898 585920 578134
rect 585320 542454 585920 577898
rect 585320 542218 585502 542454
rect 585738 542218 585920 542454
rect 585320 542134 585920 542218
rect 585320 541898 585502 542134
rect 585738 541898 585920 542134
rect 585320 506454 585920 541898
rect 585320 506218 585502 506454
rect 585738 506218 585920 506454
rect 585320 506134 585920 506218
rect 585320 505898 585502 506134
rect 585738 505898 585920 506134
rect 585320 470454 585920 505898
rect 585320 470218 585502 470454
rect 585738 470218 585920 470454
rect 585320 470134 585920 470218
rect 585320 469898 585502 470134
rect 585738 469898 585920 470134
rect 585320 434454 585920 469898
rect 585320 434218 585502 434454
rect 585738 434218 585920 434454
rect 585320 434134 585920 434218
rect 585320 433898 585502 434134
rect 585738 433898 585920 434134
rect 585320 398454 585920 433898
rect 585320 398218 585502 398454
rect 585738 398218 585920 398454
rect 585320 398134 585920 398218
rect 585320 397898 585502 398134
rect 585738 397898 585920 398134
rect 585320 362454 585920 397898
rect 585320 362218 585502 362454
rect 585738 362218 585920 362454
rect 585320 362134 585920 362218
rect 585320 361898 585502 362134
rect 585738 361898 585920 362134
rect 585320 326454 585920 361898
rect 585320 326218 585502 326454
rect 585738 326218 585920 326454
rect 585320 326134 585920 326218
rect 585320 325898 585502 326134
rect 585738 325898 585920 326134
rect 585320 290454 585920 325898
rect 585320 290218 585502 290454
rect 585738 290218 585920 290454
rect 585320 290134 585920 290218
rect 585320 289898 585502 290134
rect 585738 289898 585920 290134
rect 585320 254454 585920 289898
rect 585320 254218 585502 254454
rect 585738 254218 585920 254454
rect 585320 254134 585920 254218
rect 585320 253898 585502 254134
rect 585738 253898 585920 254134
rect 585320 218454 585920 253898
rect 585320 218218 585502 218454
rect 585738 218218 585920 218454
rect 585320 218134 585920 218218
rect 585320 217898 585502 218134
rect 585738 217898 585920 218134
rect 585320 182454 585920 217898
rect 585320 182218 585502 182454
rect 585738 182218 585920 182454
rect 585320 182134 585920 182218
rect 585320 181898 585502 182134
rect 585738 181898 585920 182134
rect 585320 146454 585920 181898
rect 585320 146218 585502 146454
rect 585738 146218 585920 146454
rect 585320 146134 585920 146218
rect 585320 145898 585502 146134
rect 585738 145898 585920 146134
rect 585320 110454 585920 145898
rect 585320 110218 585502 110454
rect 585738 110218 585920 110454
rect 585320 110134 585920 110218
rect 585320 109898 585502 110134
rect 585738 109898 585920 110134
rect 585320 74454 585920 109898
rect 585320 74218 585502 74454
rect 585738 74218 585920 74454
rect 585320 74134 585920 74218
rect 585320 73898 585502 74134
rect 585738 73898 585920 74134
rect 585320 38454 585920 73898
rect 585320 38218 585502 38454
rect 585738 38218 585920 38454
rect 585320 38134 585920 38218
rect 585320 37898 585502 38134
rect 585738 37898 585920 38134
rect 585320 2454 585920 37898
rect 585320 2218 585502 2454
rect 585738 2218 585920 2454
rect 585320 2134 585920 2218
rect 585320 1898 585502 2134
rect 585738 1898 585920 2134
rect 585320 -346 585920 1898
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586260 668454 586860 705222
rect 586260 668218 586442 668454
rect 586678 668218 586860 668454
rect 586260 668134 586860 668218
rect 586260 667898 586442 668134
rect 586678 667898 586860 668134
rect 586260 632454 586860 667898
rect 586260 632218 586442 632454
rect 586678 632218 586860 632454
rect 586260 632134 586860 632218
rect 586260 631898 586442 632134
rect 586678 631898 586860 632134
rect 586260 596454 586860 631898
rect 586260 596218 586442 596454
rect 586678 596218 586860 596454
rect 586260 596134 586860 596218
rect 586260 595898 586442 596134
rect 586678 595898 586860 596134
rect 586260 560454 586860 595898
rect 586260 560218 586442 560454
rect 586678 560218 586860 560454
rect 586260 560134 586860 560218
rect 586260 559898 586442 560134
rect 586678 559898 586860 560134
rect 586260 524454 586860 559898
rect 586260 524218 586442 524454
rect 586678 524218 586860 524454
rect 586260 524134 586860 524218
rect 586260 523898 586442 524134
rect 586678 523898 586860 524134
rect 586260 488454 586860 523898
rect 586260 488218 586442 488454
rect 586678 488218 586860 488454
rect 586260 488134 586860 488218
rect 586260 487898 586442 488134
rect 586678 487898 586860 488134
rect 586260 452454 586860 487898
rect 586260 452218 586442 452454
rect 586678 452218 586860 452454
rect 586260 452134 586860 452218
rect 586260 451898 586442 452134
rect 586678 451898 586860 452134
rect 586260 416454 586860 451898
rect 586260 416218 586442 416454
rect 586678 416218 586860 416454
rect 586260 416134 586860 416218
rect 586260 415898 586442 416134
rect 586678 415898 586860 416134
rect 586260 380454 586860 415898
rect 586260 380218 586442 380454
rect 586678 380218 586860 380454
rect 586260 380134 586860 380218
rect 586260 379898 586442 380134
rect 586678 379898 586860 380134
rect 586260 344454 586860 379898
rect 586260 344218 586442 344454
rect 586678 344218 586860 344454
rect 586260 344134 586860 344218
rect 586260 343898 586442 344134
rect 586678 343898 586860 344134
rect 586260 308454 586860 343898
rect 586260 308218 586442 308454
rect 586678 308218 586860 308454
rect 586260 308134 586860 308218
rect 586260 307898 586442 308134
rect 586678 307898 586860 308134
rect 586260 272454 586860 307898
rect 586260 272218 586442 272454
rect 586678 272218 586860 272454
rect 586260 272134 586860 272218
rect 586260 271898 586442 272134
rect 586678 271898 586860 272134
rect 586260 236454 586860 271898
rect 586260 236218 586442 236454
rect 586678 236218 586860 236454
rect 586260 236134 586860 236218
rect 586260 235898 586442 236134
rect 586678 235898 586860 236134
rect 586260 200454 586860 235898
rect 586260 200218 586442 200454
rect 586678 200218 586860 200454
rect 586260 200134 586860 200218
rect 586260 199898 586442 200134
rect 586678 199898 586860 200134
rect 586260 164454 586860 199898
rect 586260 164218 586442 164454
rect 586678 164218 586860 164454
rect 586260 164134 586860 164218
rect 586260 163898 586442 164134
rect 586678 163898 586860 164134
rect 586260 128454 586860 163898
rect 586260 128218 586442 128454
rect 586678 128218 586860 128454
rect 586260 128134 586860 128218
rect 586260 127898 586442 128134
rect 586678 127898 586860 128134
rect 586260 92454 586860 127898
rect 586260 92218 586442 92454
rect 586678 92218 586860 92454
rect 586260 92134 586860 92218
rect 586260 91898 586442 92134
rect 586678 91898 586860 92134
rect 586260 56454 586860 91898
rect 586260 56218 586442 56454
rect 586678 56218 586860 56454
rect 586260 56134 586860 56218
rect 586260 55898 586442 56134
rect 586678 55898 586860 56134
rect 586260 20454 586860 55898
rect 586260 20218 586442 20454
rect 586678 20218 586860 20454
rect 586260 20134 586860 20218
rect 586260 19898 586442 20134
rect 586678 19898 586860 20134
rect 586260 -1286 586860 19898
rect 586260 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect 586260 -1606 586860 -1522
rect 586260 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect 586260 -1864 586860 -1842
rect 587200 690054 587800 706162
rect 587200 689818 587382 690054
rect 587618 689818 587800 690054
rect 587200 689734 587800 689818
rect 587200 689498 587382 689734
rect 587618 689498 587800 689734
rect 587200 654054 587800 689498
rect 587200 653818 587382 654054
rect 587618 653818 587800 654054
rect 587200 653734 587800 653818
rect 587200 653498 587382 653734
rect 587618 653498 587800 653734
rect 587200 618054 587800 653498
rect 587200 617818 587382 618054
rect 587618 617818 587800 618054
rect 587200 617734 587800 617818
rect 587200 617498 587382 617734
rect 587618 617498 587800 617734
rect 587200 582054 587800 617498
rect 587200 581818 587382 582054
rect 587618 581818 587800 582054
rect 587200 581734 587800 581818
rect 587200 581498 587382 581734
rect 587618 581498 587800 581734
rect 587200 546054 587800 581498
rect 587200 545818 587382 546054
rect 587618 545818 587800 546054
rect 587200 545734 587800 545818
rect 587200 545498 587382 545734
rect 587618 545498 587800 545734
rect 587200 510054 587800 545498
rect 587200 509818 587382 510054
rect 587618 509818 587800 510054
rect 587200 509734 587800 509818
rect 587200 509498 587382 509734
rect 587618 509498 587800 509734
rect 587200 474054 587800 509498
rect 587200 473818 587382 474054
rect 587618 473818 587800 474054
rect 587200 473734 587800 473818
rect 587200 473498 587382 473734
rect 587618 473498 587800 473734
rect 587200 438054 587800 473498
rect 587200 437818 587382 438054
rect 587618 437818 587800 438054
rect 587200 437734 587800 437818
rect 587200 437498 587382 437734
rect 587618 437498 587800 437734
rect 587200 402054 587800 437498
rect 587200 401818 587382 402054
rect 587618 401818 587800 402054
rect 587200 401734 587800 401818
rect 587200 401498 587382 401734
rect 587618 401498 587800 401734
rect 587200 366054 587800 401498
rect 587200 365818 587382 366054
rect 587618 365818 587800 366054
rect 587200 365734 587800 365818
rect 587200 365498 587382 365734
rect 587618 365498 587800 365734
rect 587200 330054 587800 365498
rect 587200 329818 587382 330054
rect 587618 329818 587800 330054
rect 587200 329734 587800 329818
rect 587200 329498 587382 329734
rect 587618 329498 587800 329734
rect 587200 294054 587800 329498
rect 587200 293818 587382 294054
rect 587618 293818 587800 294054
rect 587200 293734 587800 293818
rect 587200 293498 587382 293734
rect 587618 293498 587800 293734
rect 587200 258054 587800 293498
rect 587200 257818 587382 258054
rect 587618 257818 587800 258054
rect 587200 257734 587800 257818
rect 587200 257498 587382 257734
rect 587618 257498 587800 257734
rect 587200 222054 587800 257498
rect 587200 221818 587382 222054
rect 587618 221818 587800 222054
rect 587200 221734 587800 221818
rect 587200 221498 587382 221734
rect 587618 221498 587800 221734
rect 587200 186054 587800 221498
rect 587200 185818 587382 186054
rect 587618 185818 587800 186054
rect 587200 185734 587800 185818
rect 587200 185498 587382 185734
rect 587618 185498 587800 185734
rect 587200 150054 587800 185498
rect 587200 149818 587382 150054
rect 587618 149818 587800 150054
rect 587200 149734 587800 149818
rect 587200 149498 587382 149734
rect 587618 149498 587800 149734
rect 587200 114054 587800 149498
rect 587200 113818 587382 114054
rect 587618 113818 587800 114054
rect 587200 113734 587800 113818
rect 587200 113498 587382 113734
rect 587618 113498 587800 113734
rect 587200 78054 587800 113498
rect 587200 77818 587382 78054
rect 587618 77818 587800 78054
rect 587200 77734 587800 77818
rect 587200 77498 587382 77734
rect 587618 77498 587800 77734
rect 587200 42054 587800 77498
rect 587200 41818 587382 42054
rect 587618 41818 587800 42054
rect 587200 41734 587800 41818
rect 587200 41498 587382 41734
rect 587618 41498 587800 41734
rect 587200 6054 587800 41498
rect 587200 5818 587382 6054
rect 587618 5818 587800 6054
rect 587200 5734 587800 5818
rect 587200 5498 587382 5734
rect 587618 5498 587800 5734
rect 580404 -2462 580586 -2226
rect 580822 -2462 581004 -2226
rect 580404 -2546 581004 -2462
rect 580404 -2782 580586 -2546
rect 580822 -2782 581004 -2546
rect 580404 -3744 581004 -2782
rect 587200 -2226 587800 5498
rect 587200 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect 587200 -2546 587800 -2462
rect 587200 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect 587200 -2804 587800 -2782
rect 588140 672054 588740 707102
rect 588140 671818 588322 672054
rect 588558 671818 588740 672054
rect 588140 671734 588740 671818
rect 588140 671498 588322 671734
rect 588558 671498 588740 671734
rect 588140 636054 588740 671498
rect 588140 635818 588322 636054
rect 588558 635818 588740 636054
rect 588140 635734 588740 635818
rect 588140 635498 588322 635734
rect 588558 635498 588740 635734
rect 588140 600054 588740 635498
rect 588140 599818 588322 600054
rect 588558 599818 588740 600054
rect 588140 599734 588740 599818
rect 588140 599498 588322 599734
rect 588558 599498 588740 599734
rect 588140 564054 588740 599498
rect 588140 563818 588322 564054
rect 588558 563818 588740 564054
rect 588140 563734 588740 563818
rect 588140 563498 588322 563734
rect 588558 563498 588740 563734
rect 588140 528054 588740 563498
rect 588140 527818 588322 528054
rect 588558 527818 588740 528054
rect 588140 527734 588740 527818
rect 588140 527498 588322 527734
rect 588558 527498 588740 527734
rect 588140 492054 588740 527498
rect 588140 491818 588322 492054
rect 588558 491818 588740 492054
rect 588140 491734 588740 491818
rect 588140 491498 588322 491734
rect 588558 491498 588740 491734
rect 588140 456054 588740 491498
rect 588140 455818 588322 456054
rect 588558 455818 588740 456054
rect 588140 455734 588740 455818
rect 588140 455498 588322 455734
rect 588558 455498 588740 455734
rect 588140 420054 588740 455498
rect 588140 419818 588322 420054
rect 588558 419818 588740 420054
rect 588140 419734 588740 419818
rect 588140 419498 588322 419734
rect 588558 419498 588740 419734
rect 588140 384054 588740 419498
rect 588140 383818 588322 384054
rect 588558 383818 588740 384054
rect 588140 383734 588740 383818
rect 588140 383498 588322 383734
rect 588558 383498 588740 383734
rect 588140 348054 588740 383498
rect 588140 347818 588322 348054
rect 588558 347818 588740 348054
rect 588140 347734 588740 347818
rect 588140 347498 588322 347734
rect 588558 347498 588740 347734
rect 588140 312054 588740 347498
rect 588140 311818 588322 312054
rect 588558 311818 588740 312054
rect 588140 311734 588740 311818
rect 588140 311498 588322 311734
rect 588558 311498 588740 311734
rect 588140 276054 588740 311498
rect 588140 275818 588322 276054
rect 588558 275818 588740 276054
rect 588140 275734 588740 275818
rect 588140 275498 588322 275734
rect 588558 275498 588740 275734
rect 588140 240054 588740 275498
rect 588140 239818 588322 240054
rect 588558 239818 588740 240054
rect 588140 239734 588740 239818
rect 588140 239498 588322 239734
rect 588558 239498 588740 239734
rect 588140 204054 588740 239498
rect 588140 203818 588322 204054
rect 588558 203818 588740 204054
rect 588140 203734 588740 203818
rect 588140 203498 588322 203734
rect 588558 203498 588740 203734
rect 588140 168054 588740 203498
rect 588140 167818 588322 168054
rect 588558 167818 588740 168054
rect 588140 167734 588740 167818
rect 588140 167498 588322 167734
rect 588558 167498 588740 167734
rect 588140 132054 588740 167498
rect 588140 131818 588322 132054
rect 588558 131818 588740 132054
rect 588140 131734 588740 131818
rect 588140 131498 588322 131734
rect 588558 131498 588740 131734
rect 588140 96054 588740 131498
rect 588140 95818 588322 96054
rect 588558 95818 588740 96054
rect 588140 95734 588740 95818
rect 588140 95498 588322 95734
rect 588558 95498 588740 95734
rect 588140 60054 588740 95498
rect 588140 59818 588322 60054
rect 588558 59818 588740 60054
rect 588140 59734 588740 59818
rect 588140 59498 588322 59734
rect 588558 59498 588740 59734
rect 588140 24054 588740 59498
rect 588140 23818 588322 24054
rect 588558 23818 588740 24054
rect 588140 23734 588740 23818
rect 588140 23498 588322 23734
rect 588558 23498 588740 23734
rect 588140 -3166 588740 23498
rect 588140 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect 588140 -3486 588740 -3402
rect 588140 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect 588140 -3744 588740 -3722
rect 589080 693654 589680 708042
rect 589080 693418 589262 693654
rect 589498 693418 589680 693654
rect 589080 693334 589680 693418
rect 589080 693098 589262 693334
rect 589498 693098 589680 693334
rect 589080 657654 589680 693098
rect 589080 657418 589262 657654
rect 589498 657418 589680 657654
rect 589080 657334 589680 657418
rect 589080 657098 589262 657334
rect 589498 657098 589680 657334
rect 589080 621654 589680 657098
rect 589080 621418 589262 621654
rect 589498 621418 589680 621654
rect 589080 621334 589680 621418
rect 589080 621098 589262 621334
rect 589498 621098 589680 621334
rect 589080 585654 589680 621098
rect 589080 585418 589262 585654
rect 589498 585418 589680 585654
rect 589080 585334 589680 585418
rect 589080 585098 589262 585334
rect 589498 585098 589680 585334
rect 589080 549654 589680 585098
rect 589080 549418 589262 549654
rect 589498 549418 589680 549654
rect 589080 549334 589680 549418
rect 589080 549098 589262 549334
rect 589498 549098 589680 549334
rect 589080 513654 589680 549098
rect 589080 513418 589262 513654
rect 589498 513418 589680 513654
rect 589080 513334 589680 513418
rect 589080 513098 589262 513334
rect 589498 513098 589680 513334
rect 589080 477654 589680 513098
rect 589080 477418 589262 477654
rect 589498 477418 589680 477654
rect 589080 477334 589680 477418
rect 589080 477098 589262 477334
rect 589498 477098 589680 477334
rect 589080 441654 589680 477098
rect 589080 441418 589262 441654
rect 589498 441418 589680 441654
rect 589080 441334 589680 441418
rect 589080 441098 589262 441334
rect 589498 441098 589680 441334
rect 589080 405654 589680 441098
rect 589080 405418 589262 405654
rect 589498 405418 589680 405654
rect 589080 405334 589680 405418
rect 589080 405098 589262 405334
rect 589498 405098 589680 405334
rect 589080 369654 589680 405098
rect 589080 369418 589262 369654
rect 589498 369418 589680 369654
rect 589080 369334 589680 369418
rect 589080 369098 589262 369334
rect 589498 369098 589680 369334
rect 589080 333654 589680 369098
rect 589080 333418 589262 333654
rect 589498 333418 589680 333654
rect 589080 333334 589680 333418
rect 589080 333098 589262 333334
rect 589498 333098 589680 333334
rect 589080 297654 589680 333098
rect 589080 297418 589262 297654
rect 589498 297418 589680 297654
rect 589080 297334 589680 297418
rect 589080 297098 589262 297334
rect 589498 297098 589680 297334
rect 589080 261654 589680 297098
rect 589080 261418 589262 261654
rect 589498 261418 589680 261654
rect 589080 261334 589680 261418
rect 589080 261098 589262 261334
rect 589498 261098 589680 261334
rect 589080 225654 589680 261098
rect 589080 225418 589262 225654
rect 589498 225418 589680 225654
rect 589080 225334 589680 225418
rect 589080 225098 589262 225334
rect 589498 225098 589680 225334
rect 589080 189654 589680 225098
rect 589080 189418 589262 189654
rect 589498 189418 589680 189654
rect 589080 189334 589680 189418
rect 589080 189098 589262 189334
rect 589498 189098 589680 189334
rect 589080 153654 589680 189098
rect 589080 153418 589262 153654
rect 589498 153418 589680 153654
rect 589080 153334 589680 153418
rect 589080 153098 589262 153334
rect 589498 153098 589680 153334
rect 589080 117654 589680 153098
rect 589080 117418 589262 117654
rect 589498 117418 589680 117654
rect 589080 117334 589680 117418
rect 589080 117098 589262 117334
rect 589498 117098 589680 117334
rect 589080 81654 589680 117098
rect 589080 81418 589262 81654
rect 589498 81418 589680 81654
rect 589080 81334 589680 81418
rect 589080 81098 589262 81334
rect 589498 81098 589680 81334
rect 589080 45654 589680 81098
rect 589080 45418 589262 45654
rect 589498 45418 589680 45654
rect 589080 45334 589680 45418
rect 589080 45098 589262 45334
rect 589498 45098 589680 45334
rect 589080 9654 589680 45098
rect 589080 9418 589262 9654
rect 589498 9418 589680 9654
rect 589080 9334 589680 9418
rect 589080 9098 589262 9334
rect 589498 9098 589680 9334
rect 589080 -4106 589680 9098
rect 589080 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect 589080 -4426 589680 -4342
rect 589080 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect 589080 -4684 589680 -4662
rect 590020 675654 590620 708982
rect 590020 675418 590202 675654
rect 590438 675418 590620 675654
rect 590020 675334 590620 675418
rect 590020 675098 590202 675334
rect 590438 675098 590620 675334
rect 590020 639654 590620 675098
rect 590020 639418 590202 639654
rect 590438 639418 590620 639654
rect 590020 639334 590620 639418
rect 590020 639098 590202 639334
rect 590438 639098 590620 639334
rect 590020 603654 590620 639098
rect 590020 603418 590202 603654
rect 590438 603418 590620 603654
rect 590020 603334 590620 603418
rect 590020 603098 590202 603334
rect 590438 603098 590620 603334
rect 590020 567654 590620 603098
rect 590020 567418 590202 567654
rect 590438 567418 590620 567654
rect 590020 567334 590620 567418
rect 590020 567098 590202 567334
rect 590438 567098 590620 567334
rect 590020 531654 590620 567098
rect 590020 531418 590202 531654
rect 590438 531418 590620 531654
rect 590020 531334 590620 531418
rect 590020 531098 590202 531334
rect 590438 531098 590620 531334
rect 590020 495654 590620 531098
rect 590020 495418 590202 495654
rect 590438 495418 590620 495654
rect 590020 495334 590620 495418
rect 590020 495098 590202 495334
rect 590438 495098 590620 495334
rect 590020 459654 590620 495098
rect 590020 459418 590202 459654
rect 590438 459418 590620 459654
rect 590020 459334 590620 459418
rect 590020 459098 590202 459334
rect 590438 459098 590620 459334
rect 590020 423654 590620 459098
rect 590020 423418 590202 423654
rect 590438 423418 590620 423654
rect 590020 423334 590620 423418
rect 590020 423098 590202 423334
rect 590438 423098 590620 423334
rect 590020 387654 590620 423098
rect 590020 387418 590202 387654
rect 590438 387418 590620 387654
rect 590020 387334 590620 387418
rect 590020 387098 590202 387334
rect 590438 387098 590620 387334
rect 590020 351654 590620 387098
rect 590020 351418 590202 351654
rect 590438 351418 590620 351654
rect 590020 351334 590620 351418
rect 590020 351098 590202 351334
rect 590438 351098 590620 351334
rect 590020 315654 590620 351098
rect 590020 315418 590202 315654
rect 590438 315418 590620 315654
rect 590020 315334 590620 315418
rect 590020 315098 590202 315334
rect 590438 315098 590620 315334
rect 590020 279654 590620 315098
rect 590020 279418 590202 279654
rect 590438 279418 590620 279654
rect 590020 279334 590620 279418
rect 590020 279098 590202 279334
rect 590438 279098 590620 279334
rect 590020 243654 590620 279098
rect 590020 243418 590202 243654
rect 590438 243418 590620 243654
rect 590020 243334 590620 243418
rect 590020 243098 590202 243334
rect 590438 243098 590620 243334
rect 590020 207654 590620 243098
rect 590020 207418 590202 207654
rect 590438 207418 590620 207654
rect 590020 207334 590620 207418
rect 590020 207098 590202 207334
rect 590438 207098 590620 207334
rect 590020 171654 590620 207098
rect 590020 171418 590202 171654
rect 590438 171418 590620 171654
rect 590020 171334 590620 171418
rect 590020 171098 590202 171334
rect 590438 171098 590620 171334
rect 590020 135654 590620 171098
rect 590020 135418 590202 135654
rect 590438 135418 590620 135654
rect 590020 135334 590620 135418
rect 590020 135098 590202 135334
rect 590438 135098 590620 135334
rect 590020 99654 590620 135098
rect 590020 99418 590202 99654
rect 590438 99418 590620 99654
rect 590020 99334 590620 99418
rect 590020 99098 590202 99334
rect 590438 99098 590620 99334
rect 590020 63654 590620 99098
rect 590020 63418 590202 63654
rect 590438 63418 590620 63654
rect 590020 63334 590620 63418
rect 590020 63098 590202 63334
rect 590438 63098 590620 63334
rect 590020 27654 590620 63098
rect 590020 27418 590202 27654
rect 590438 27418 590620 27654
rect 590020 27334 590620 27418
rect 590020 27098 590202 27334
rect 590438 27098 590620 27334
rect 590020 -5046 590620 27098
rect 590020 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect 590020 -5366 590620 -5282
rect 590020 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect 590020 -5624 590620 -5602
rect 590960 697254 591560 709922
rect 590960 697018 591142 697254
rect 591378 697018 591560 697254
rect 590960 696934 591560 697018
rect 590960 696698 591142 696934
rect 591378 696698 591560 696934
rect 590960 661254 591560 696698
rect 590960 661018 591142 661254
rect 591378 661018 591560 661254
rect 590960 660934 591560 661018
rect 590960 660698 591142 660934
rect 591378 660698 591560 660934
rect 590960 625254 591560 660698
rect 590960 625018 591142 625254
rect 591378 625018 591560 625254
rect 590960 624934 591560 625018
rect 590960 624698 591142 624934
rect 591378 624698 591560 624934
rect 590960 589254 591560 624698
rect 590960 589018 591142 589254
rect 591378 589018 591560 589254
rect 590960 588934 591560 589018
rect 590960 588698 591142 588934
rect 591378 588698 591560 588934
rect 590960 553254 591560 588698
rect 590960 553018 591142 553254
rect 591378 553018 591560 553254
rect 590960 552934 591560 553018
rect 590960 552698 591142 552934
rect 591378 552698 591560 552934
rect 590960 517254 591560 552698
rect 590960 517018 591142 517254
rect 591378 517018 591560 517254
rect 590960 516934 591560 517018
rect 590960 516698 591142 516934
rect 591378 516698 591560 516934
rect 590960 481254 591560 516698
rect 590960 481018 591142 481254
rect 591378 481018 591560 481254
rect 590960 480934 591560 481018
rect 590960 480698 591142 480934
rect 591378 480698 591560 480934
rect 590960 445254 591560 480698
rect 590960 445018 591142 445254
rect 591378 445018 591560 445254
rect 590960 444934 591560 445018
rect 590960 444698 591142 444934
rect 591378 444698 591560 444934
rect 590960 409254 591560 444698
rect 590960 409018 591142 409254
rect 591378 409018 591560 409254
rect 590960 408934 591560 409018
rect 590960 408698 591142 408934
rect 591378 408698 591560 408934
rect 590960 373254 591560 408698
rect 590960 373018 591142 373254
rect 591378 373018 591560 373254
rect 590960 372934 591560 373018
rect 590960 372698 591142 372934
rect 591378 372698 591560 372934
rect 590960 337254 591560 372698
rect 590960 337018 591142 337254
rect 591378 337018 591560 337254
rect 590960 336934 591560 337018
rect 590960 336698 591142 336934
rect 591378 336698 591560 336934
rect 590960 301254 591560 336698
rect 590960 301018 591142 301254
rect 591378 301018 591560 301254
rect 590960 300934 591560 301018
rect 590960 300698 591142 300934
rect 591378 300698 591560 300934
rect 590960 265254 591560 300698
rect 590960 265018 591142 265254
rect 591378 265018 591560 265254
rect 590960 264934 591560 265018
rect 590960 264698 591142 264934
rect 591378 264698 591560 264934
rect 590960 229254 591560 264698
rect 590960 229018 591142 229254
rect 591378 229018 591560 229254
rect 590960 228934 591560 229018
rect 590960 228698 591142 228934
rect 591378 228698 591560 228934
rect 590960 193254 591560 228698
rect 590960 193018 591142 193254
rect 591378 193018 591560 193254
rect 590960 192934 591560 193018
rect 590960 192698 591142 192934
rect 591378 192698 591560 192934
rect 590960 157254 591560 192698
rect 590960 157018 591142 157254
rect 591378 157018 591560 157254
rect 590960 156934 591560 157018
rect 590960 156698 591142 156934
rect 591378 156698 591560 156934
rect 590960 121254 591560 156698
rect 590960 121018 591142 121254
rect 591378 121018 591560 121254
rect 590960 120934 591560 121018
rect 590960 120698 591142 120934
rect 591378 120698 591560 120934
rect 590960 85254 591560 120698
rect 590960 85018 591142 85254
rect 591378 85018 591560 85254
rect 590960 84934 591560 85018
rect 590960 84698 591142 84934
rect 591378 84698 591560 84934
rect 590960 49254 591560 84698
rect 590960 49018 591142 49254
rect 591378 49018 591560 49254
rect 590960 48934 591560 49018
rect 590960 48698 591142 48934
rect 591378 48698 591560 48934
rect 590960 13254 591560 48698
rect 590960 13018 591142 13254
rect 591378 13018 591560 13254
rect 590960 12934 591560 13018
rect 590960 12698 591142 12934
rect 591378 12698 591560 12934
rect 590960 -5986 591560 12698
rect 590960 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect 590960 -6306 591560 -6222
rect 590960 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect 590960 -6564 591560 -6542
rect 591900 679254 592500 710862
rect 591900 679018 592082 679254
rect 592318 679018 592500 679254
rect 591900 678934 592500 679018
rect 591900 678698 592082 678934
rect 592318 678698 592500 678934
rect 591900 643254 592500 678698
rect 591900 643018 592082 643254
rect 592318 643018 592500 643254
rect 591900 642934 592500 643018
rect 591900 642698 592082 642934
rect 592318 642698 592500 642934
rect 591900 607254 592500 642698
rect 591900 607018 592082 607254
rect 592318 607018 592500 607254
rect 591900 606934 592500 607018
rect 591900 606698 592082 606934
rect 592318 606698 592500 606934
rect 591900 571254 592500 606698
rect 591900 571018 592082 571254
rect 592318 571018 592500 571254
rect 591900 570934 592500 571018
rect 591900 570698 592082 570934
rect 592318 570698 592500 570934
rect 591900 535254 592500 570698
rect 591900 535018 592082 535254
rect 592318 535018 592500 535254
rect 591900 534934 592500 535018
rect 591900 534698 592082 534934
rect 592318 534698 592500 534934
rect 591900 499254 592500 534698
rect 591900 499018 592082 499254
rect 592318 499018 592500 499254
rect 591900 498934 592500 499018
rect 591900 498698 592082 498934
rect 592318 498698 592500 498934
rect 591900 463254 592500 498698
rect 591900 463018 592082 463254
rect 592318 463018 592500 463254
rect 591900 462934 592500 463018
rect 591900 462698 592082 462934
rect 592318 462698 592500 462934
rect 591900 427254 592500 462698
rect 591900 427018 592082 427254
rect 592318 427018 592500 427254
rect 591900 426934 592500 427018
rect 591900 426698 592082 426934
rect 592318 426698 592500 426934
rect 591900 391254 592500 426698
rect 591900 391018 592082 391254
rect 592318 391018 592500 391254
rect 591900 390934 592500 391018
rect 591900 390698 592082 390934
rect 592318 390698 592500 390934
rect 591900 355254 592500 390698
rect 591900 355018 592082 355254
rect 592318 355018 592500 355254
rect 591900 354934 592500 355018
rect 591900 354698 592082 354934
rect 592318 354698 592500 354934
rect 591900 319254 592500 354698
rect 591900 319018 592082 319254
rect 592318 319018 592500 319254
rect 591900 318934 592500 319018
rect 591900 318698 592082 318934
rect 592318 318698 592500 318934
rect 591900 283254 592500 318698
rect 591900 283018 592082 283254
rect 592318 283018 592500 283254
rect 591900 282934 592500 283018
rect 591900 282698 592082 282934
rect 592318 282698 592500 282934
rect 591900 247254 592500 282698
rect 591900 247018 592082 247254
rect 592318 247018 592500 247254
rect 591900 246934 592500 247018
rect 591900 246698 592082 246934
rect 592318 246698 592500 246934
rect 591900 211254 592500 246698
rect 591900 211018 592082 211254
rect 592318 211018 592500 211254
rect 591900 210934 592500 211018
rect 591900 210698 592082 210934
rect 592318 210698 592500 210934
rect 591900 175254 592500 210698
rect 591900 175018 592082 175254
rect 592318 175018 592500 175254
rect 591900 174934 592500 175018
rect 591900 174698 592082 174934
rect 592318 174698 592500 174934
rect 591900 139254 592500 174698
rect 591900 139018 592082 139254
rect 592318 139018 592500 139254
rect 591900 138934 592500 139018
rect 591900 138698 592082 138934
rect 592318 138698 592500 138934
rect 591900 103254 592500 138698
rect 591900 103018 592082 103254
rect 592318 103018 592500 103254
rect 591900 102934 592500 103018
rect 591900 102698 592082 102934
rect 592318 102698 592500 102934
rect 591900 67254 592500 102698
rect 591900 67018 592082 67254
rect 592318 67018 592500 67254
rect 591900 66934 592500 67018
rect 591900 66698 592082 66934
rect 592318 66698 592500 66934
rect 591900 31254 592500 66698
rect 591900 31018 592082 31254
rect 592318 31018 592500 31254
rect 591900 30934 592500 31018
rect 591900 30698 592082 30934
rect 592318 30698 592500 30934
rect 569604 -7162 569786 -6926
rect 570022 -7162 570204 -6926
rect 569604 -7246 570204 -7162
rect 569604 -7482 569786 -7246
rect 570022 -7482 570204 -7246
rect 569604 -7504 570204 -7482
rect 591900 -6926 592500 30698
rect 591900 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect 591900 -7246 592500 -7162
rect 591900 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect 591900 -7504 592500 -7482
<< via4 >>
rect -8394 711182 -8158 711418
rect -8394 710862 -8158 711098
rect -8394 679018 -8158 679254
rect -8394 678698 -8158 678934
rect -8394 643018 -8158 643254
rect -8394 642698 -8158 642934
rect -8394 607018 -8158 607254
rect -8394 606698 -8158 606934
rect -8394 571018 -8158 571254
rect -8394 570698 -8158 570934
rect -8394 535018 -8158 535254
rect -8394 534698 -8158 534934
rect -8394 499018 -8158 499254
rect -8394 498698 -8158 498934
rect -8394 463018 -8158 463254
rect -8394 462698 -8158 462934
rect -8394 427018 -8158 427254
rect -8394 426698 -8158 426934
rect -8394 391018 -8158 391254
rect -8394 390698 -8158 390934
rect -8394 355018 -8158 355254
rect -8394 354698 -8158 354934
rect -8394 319018 -8158 319254
rect -8394 318698 -8158 318934
rect -8394 283018 -8158 283254
rect -8394 282698 -8158 282934
rect -8394 247018 -8158 247254
rect -8394 246698 -8158 246934
rect -8394 211018 -8158 211254
rect -8394 210698 -8158 210934
rect -8394 175018 -8158 175254
rect -8394 174698 -8158 174934
rect -8394 139018 -8158 139254
rect -8394 138698 -8158 138934
rect -8394 103018 -8158 103254
rect -8394 102698 -8158 102934
rect -8394 67018 -8158 67254
rect -8394 66698 -8158 66934
rect -8394 31018 -8158 31254
rect -8394 30698 -8158 30934
rect -7454 710242 -7218 710478
rect -7454 709922 -7218 710158
rect 11786 710242 12022 710478
rect 11786 709922 12022 710158
rect -7454 697018 -7218 697254
rect -7454 696698 -7218 696934
rect -7454 661018 -7218 661254
rect -7454 660698 -7218 660934
rect -7454 625018 -7218 625254
rect -7454 624698 -7218 624934
rect -7454 589018 -7218 589254
rect -7454 588698 -7218 588934
rect -7454 553018 -7218 553254
rect -7454 552698 -7218 552934
rect -7454 517018 -7218 517254
rect -7454 516698 -7218 516934
rect -7454 481018 -7218 481254
rect -7454 480698 -7218 480934
rect -7454 445018 -7218 445254
rect -7454 444698 -7218 444934
rect -7454 409018 -7218 409254
rect -7454 408698 -7218 408934
rect -7454 373018 -7218 373254
rect -7454 372698 -7218 372934
rect -7454 337018 -7218 337254
rect -7454 336698 -7218 336934
rect -7454 301018 -7218 301254
rect -7454 300698 -7218 300934
rect -7454 265018 -7218 265254
rect -7454 264698 -7218 264934
rect -7454 229018 -7218 229254
rect -7454 228698 -7218 228934
rect -7454 193018 -7218 193254
rect -7454 192698 -7218 192934
rect -7454 157018 -7218 157254
rect -7454 156698 -7218 156934
rect -7454 121018 -7218 121254
rect -7454 120698 -7218 120934
rect -7454 85018 -7218 85254
rect -7454 84698 -7218 84934
rect -7454 49018 -7218 49254
rect -7454 48698 -7218 48934
rect -7454 13018 -7218 13254
rect -7454 12698 -7218 12934
rect -6514 709302 -6278 709538
rect -6514 708982 -6278 709218
rect -6514 675418 -6278 675654
rect -6514 675098 -6278 675334
rect -6514 639418 -6278 639654
rect -6514 639098 -6278 639334
rect -6514 603418 -6278 603654
rect -6514 603098 -6278 603334
rect -6514 567418 -6278 567654
rect -6514 567098 -6278 567334
rect -6514 531418 -6278 531654
rect -6514 531098 -6278 531334
rect -6514 495418 -6278 495654
rect -6514 495098 -6278 495334
rect -6514 459418 -6278 459654
rect -6514 459098 -6278 459334
rect -6514 423418 -6278 423654
rect -6514 423098 -6278 423334
rect -6514 387418 -6278 387654
rect -6514 387098 -6278 387334
rect -6514 351418 -6278 351654
rect -6514 351098 -6278 351334
rect -6514 315418 -6278 315654
rect -6514 315098 -6278 315334
rect -6514 279418 -6278 279654
rect -6514 279098 -6278 279334
rect -6514 243418 -6278 243654
rect -6514 243098 -6278 243334
rect -6514 207418 -6278 207654
rect -6514 207098 -6278 207334
rect -6514 171418 -6278 171654
rect -6514 171098 -6278 171334
rect -6514 135418 -6278 135654
rect -6514 135098 -6278 135334
rect -6514 99418 -6278 99654
rect -6514 99098 -6278 99334
rect -6514 63418 -6278 63654
rect -6514 63098 -6278 63334
rect -6514 27418 -6278 27654
rect -6514 27098 -6278 27334
rect -5574 708362 -5338 708598
rect -5574 708042 -5338 708278
rect 8186 708362 8422 708598
rect 8186 708042 8422 708278
rect -5574 693418 -5338 693654
rect -5574 693098 -5338 693334
rect -5574 657418 -5338 657654
rect -5574 657098 -5338 657334
rect -5574 621418 -5338 621654
rect -5574 621098 -5338 621334
rect -5574 585418 -5338 585654
rect -5574 585098 -5338 585334
rect -5574 549418 -5338 549654
rect -5574 549098 -5338 549334
rect -5574 513418 -5338 513654
rect -5574 513098 -5338 513334
rect -5574 477418 -5338 477654
rect -5574 477098 -5338 477334
rect -5574 441418 -5338 441654
rect -5574 441098 -5338 441334
rect -5574 405418 -5338 405654
rect -5574 405098 -5338 405334
rect -5574 369418 -5338 369654
rect -5574 369098 -5338 369334
rect -5574 333418 -5338 333654
rect -5574 333098 -5338 333334
rect -5574 297418 -5338 297654
rect -5574 297098 -5338 297334
rect -5574 261418 -5338 261654
rect -5574 261098 -5338 261334
rect -5574 225418 -5338 225654
rect -5574 225098 -5338 225334
rect -5574 189418 -5338 189654
rect -5574 189098 -5338 189334
rect -5574 153418 -5338 153654
rect -5574 153098 -5338 153334
rect -5574 117418 -5338 117654
rect -5574 117098 -5338 117334
rect -5574 81418 -5338 81654
rect -5574 81098 -5338 81334
rect -5574 45418 -5338 45654
rect -5574 45098 -5338 45334
rect -5574 9418 -5338 9654
rect -5574 9098 -5338 9334
rect -4634 707422 -4398 707658
rect -4634 707102 -4398 707338
rect -4634 671818 -4398 672054
rect -4634 671498 -4398 671734
rect -4634 635818 -4398 636054
rect -4634 635498 -4398 635734
rect -4634 599818 -4398 600054
rect -4634 599498 -4398 599734
rect -4634 563818 -4398 564054
rect -4634 563498 -4398 563734
rect -4634 527818 -4398 528054
rect -4634 527498 -4398 527734
rect -4634 491818 -4398 492054
rect -4634 491498 -4398 491734
rect -4634 455818 -4398 456054
rect -4634 455498 -4398 455734
rect -4634 419818 -4398 420054
rect -4634 419498 -4398 419734
rect -4634 383818 -4398 384054
rect -4634 383498 -4398 383734
rect -4634 347818 -4398 348054
rect -4634 347498 -4398 347734
rect -4634 311818 -4398 312054
rect -4634 311498 -4398 311734
rect -4634 275818 -4398 276054
rect -4634 275498 -4398 275734
rect -4634 239818 -4398 240054
rect -4634 239498 -4398 239734
rect -4634 203818 -4398 204054
rect -4634 203498 -4398 203734
rect -4634 167818 -4398 168054
rect -4634 167498 -4398 167734
rect -4634 131818 -4398 132054
rect -4634 131498 -4398 131734
rect -4634 95818 -4398 96054
rect -4634 95498 -4398 95734
rect -4634 59818 -4398 60054
rect -4634 59498 -4398 59734
rect -4634 23818 -4398 24054
rect -4634 23498 -4398 23734
rect -3694 706482 -3458 706718
rect -3694 706162 -3458 706398
rect 4586 706482 4822 706718
rect 4586 706162 4822 706398
rect -3694 689818 -3458 690054
rect -3694 689498 -3458 689734
rect -3694 653818 -3458 654054
rect -3694 653498 -3458 653734
rect -3694 617818 -3458 618054
rect -3694 617498 -3458 617734
rect -3694 581818 -3458 582054
rect -3694 581498 -3458 581734
rect -3694 545818 -3458 546054
rect -3694 545498 -3458 545734
rect -3694 509818 -3458 510054
rect -3694 509498 -3458 509734
rect -3694 473818 -3458 474054
rect -3694 473498 -3458 473734
rect -3694 437818 -3458 438054
rect -3694 437498 -3458 437734
rect -3694 401818 -3458 402054
rect -3694 401498 -3458 401734
rect -3694 365818 -3458 366054
rect -3694 365498 -3458 365734
rect -3694 329818 -3458 330054
rect -3694 329498 -3458 329734
rect -3694 293818 -3458 294054
rect -3694 293498 -3458 293734
rect -3694 257818 -3458 258054
rect -3694 257498 -3458 257734
rect -3694 221818 -3458 222054
rect -3694 221498 -3458 221734
rect -3694 185818 -3458 186054
rect -3694 185498 -3458 185734
rect -3694 149818 -3458 150054
rect -3694 149498 -3458 149734
rect -3694 113818 -3458 114054
rect -3694 113498 -3458 113734
rect -3694 77818 -3458 78054
rect -3694 77498 -3458 77734
rect -3694 41818 -3458 42054
rect -3694 41498 -3458 41734
rect -3694 5818 -3458 6054
rect -3694 5498 -3458 5734
rect -2754 705542 -2518 705778
rect -2754 705222 -2518 705458
rect -2754 668218 -2518 668454
rect -2754 667898 -2518 668134
rect -2754 632218 -2518 632454
rect -2754 631898 -2518 632134
rect -2754 596218 -2518 596454
rect -2754 595898 -2518 596134
rect -2754 560218 -2518 560454
rect -2754 559898 -2518 560134
rect -2754 524218 -2518 524454
rect -2754 523898 -2518 524134
rect -2754 488218 -2518 488454
rect -2754 487898 -2518 488134
rect -2754 452218 -2518 452454
rect -2754 451898 -2518 452134
rect -2754 416218 -2518 416454
rect -2754 415898 -2518 416134
rect -2754 380218 -2518 380454
rect -2754 379898 -2518 380134
rect -2754 344218 -2518 344454
rect -2754 343898 -2518 344134
rect -2754 308218 -2518 308454
rect -2754 307898 -2518 308134
rect -2754 272218 -2518 272454
rect -2754 271898 -2518 272134
rect -2754 236218 -2518 236454
rect -2754 235898 -2518 236134
rect -2754 200218 -2518 200454
rect -2754 199898 -2518 200134
rect -2754 164218 -2518 164454
rect -2754 163898 -2518 164134
rect -2754 128218 -2518 128454
rect -2754 127898 -2518 128134
rect -2754 92218 -2518 92454
rect -2754 91898 -2518 92134
rect -2754 56218 -2518 56454
rect -2754 55898 -2518 56134
rect -2754 20218 -2518 20454
rect -2754 19898 -2518 20134
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect -1814 686218 -1578 686454
rect -1814 685898 -1578 686134
rect -1814 650218 -1578 650454
rect -1814 649898 -1578 650134
rect -1814 614218 -1578 614454
rect -1814 613898 -1578 614134
rect -1814 578218 -1578 578454
rect -1814 577898 -1578 578134
rect -1814 542218 -1578 542454
rect -1814 541898 -1578 542134
rect -1814 506218 -1578 506454
rect -1814 505898 -1578 506134
rect -1814 470218 -1578 470454
rect -1814 469898 -1578 470134
rect -1814 434218 -1578 434454
rect -1814 433898 -1578 434134
rect -1814 398218 -1578 398454
rect -1814 397898 -1578 398134
rect -1814 362218 -1578 362454
rect -1814 361898 -1578 362134
rect -1814 326218 -1578 326454
rect -1814 325898 -1578 326134
rect -1814 290218 -1578 290454
rect -1814 289898 -1578 290134
rect -1814 254218 -1578 254454
rect -1814 253898 -1578 254134
rect -1814 218218 -1578 218454
rect -1814 217898 -1578 218134
rect -1814 182218 -1578 182454
rect -1814 181898 -1578 182134
rect -1814 146218 -1578 146454
rect -1814 145898 -1578 146134
rect -1814 110218 -1578 110454
rect -1814 109898 -1578 110134
rect -1814 74218 -1578 74454
rect -1814 73898 -1578 74134
rect -1814 38218 -1578 38454
rect -1814 37898 -1578 38134
rect -1814 2218 -1578 2454
rect -1814 1898 -1578 2134
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 986 704602 1222 704838
rect 986 704282 1222 704518
rect 986 686218 1222 686454
rect 986 685898 1222 686134
rect 986 650218 1222 650454
rect 986 649898 1222 650134
rect 986 614218 1222 614454
rect 986 613898 1222 614134
rect 986 578218 1222 578454
rect 986 577898 1222 578134
rect 986 542218 1222 542454
rect 986 541898 1222 542134
rect 986 506218 1222 506454
rect 986 505898 1222 506134
rect 986 470218 1222 470454
rect 986 469898 1222 470134
rect 986 434218 1222 434454
rect 986 433898 1222 434134
rect 986 398218 1222 398454
rect 986 397898 1222 398134
rect 986 362218 1222 362454
rect 986 361898 1222 362134
rect 986 326218 1222 326454
rect 986 325898 1222 326134
rect 986 290218 1222 290454
rect 986 289898 1222 290134
rect 986 254218 1222 254454
rect 986 253898 1222 254134
rect 986 218218 1222 218454
rect 986 217898 1222 218134
rect 986 182218 1222 182454
rect 986 181898 1222 182134
rect 986 146218 1222 146454
rect 986 145898 1222 146134
rect 986 110218 1222 110454
rect 986 109898 1222 110134
rect 986 74218 1222 74454
rect 986 73898 1222 74134
rect 986 38218 1222 38454
rect 986 37898 1222 38134
rect 986 2218 1222 2454
rect 986 1898 1222 2134
rect 986 -582 1222 -346
rect 986 -902 1222 -666
rect -2754 -1522 -2518 -1286
rect -2754 -1842 -2518 -1606
rect 4586 689818 4822 690054
rect 4586 689498 4822 689734
rect 4586 653818 4822 654054
rect 4586 653498 4822 653734
rect 4586 617818 4822 618054
rect 4586 617498 4822 617734
rect 4586 581818 4822 582054
rect 4586 581498 4822 581734
rect 4586 545818 4822 546054
rect 4586 545498 4822 545734
rect 4586 509818 4822 510054
rect 4586 509498 4822 509734
rect 4586 473818 4822 474054
rect 4586 473498 4822 473734
rect 4586 437818 4822 438054
rect 4586 437498 4822 437734
rect 4586 401818 4822 402054
rect 4586 401498 4822 401734
rect 4586 365818 4822 366054
rect 4586 365498 4822 365734
rect 4586 329818 4822 330054
rect 4586 329498 4822 329734
rect 4586 293818 4822 294054
rect 4586 293498 4822 293734
rect 4586 257818 4822 258054
rect 4586 257498 4822 257734
rect 4586 221818 4822 222054
rect 4586 221498 4822 221734
rect 4586 185818 4822 186054
rect 4586 185498 4822 185734
rect 4586 149818 4822 150054
rect 4586 149498 4822 149734
rect 4586 113818 4822 114054
rect 4586 113498 4822 113734
rect 4586 77818 4822 78054
rect 4586 77498 4822 77734
rect 4586 41818 4822 42054
rect 4586 41498 4822 41734
rect 4586 5818 4822 6054
rect 4586 5498 4822 5734
rect -3694 -2462 -3458 -2226
rect -3694 -2782 -3458 -2546
rect 4586 -2462 4822 -2226
rect 4586 -2782 4822 -2546
rect -4634 -3402 -4398 -3166
rect -4634 -3722 -4398 -3486
rect 8186 693418 8422 693654
rect 8186 693098 8422 693334
rect 8186 657418 8422 657654
rect 8186 657098 8422 657334
rect 8186 621418 8422 621654
rect 8186 621098 8422 621334
rect 8186 585418 8422 585654
rect 8186 585098 8422 585334
rect 8186 549418 8422 549654
rect 8186 549098 8422 549334
rect 8186 513418 8422 513654
rect 8186 513098 8422 513334
rect 8186 477418 8422 477654
rect 8186 477098 8422 477334
rect 8186 441418 8422 441654
rect 8186 441098 8422 441334
rect 8186 405418 8422 405654
rect 8186 405098 8422 405334
rect 8186 369418 8422 369654
rect 8186 369098 8422 369334
rect 8186 333418 8422 333654
rect 8186 333098 8422 333334
rect 8186 297418 8422 297654
rect 8186 297098 8422 297334
rect 8186 261418 8422 261654
rect 8186 261098 8422 261334
rect 8186 225418 8422 225654
rect 8186 225098 8422 225334
rect 8186 189418 8422 189654
rect 8186 189098 8422 189334
rect 8186 153418 8422 153654
rect 8186 153098 8422 153334
rect 8186 117418 8422 117654
rect 8186 117098 8422 117334
rect 8186 81418 8422 81654
rect 8186 81098 8422 81334
rect 8186 45418 8422 45654
rect 8186 45098 8422 45334
rect 8186 9418 8422 9654
rect 8186 9098 8422 9334
rect -5574 -4342 -5338 -4106
rect -5574 -4662 -5338 -4426
rect 8186 -4342 8422 -4106
rect 8186 -4662 8422 -4426
rect -6514 -5282 -6278 -5046
rect -6514 -5602 -6278 -5366
rect 29786 711182 30022 711418
rect 29786 710862 30022 711098
rect 26186 709302 26422 709538
rect 26186 708982 26422 709218
rect 22586 707422 22822 707658
rect 22586 707102 22822 707338
rect 11786 697018 12022 697254
rect 11786 696698 12022 696934
rect 11786 661018 12022 661254
rect 11786 660698 12022 660934
rect 11786 625018 12022 625254
rect 11786 624698 12022 624934
rect 11786 589018 12022 589254
rect 11786 588698 12022 588934
rect 11786 553018 12022 553254
rect 11786 552698 12022 552934
rect 11786 517018 12022 517254
rect 11786 516698 12022 516934
rect 11786 481018 12022 481254
rect 11786 480698 12022 480934
rect 11786 445018 12022 445254
rect 11786 444698 12022 444934
rect 11786 409018 12022 409254
rect 11786 408698 12022 408934
rect 11786 373018 12022 373254
rect 11786 372698 12022 372934
rect 11786 337018 12022 337254
rect 11786 336698 12022 336934
rect 11786 301018 12022 301254
rect 11786 300698 12022 300934
rect 11786 265018 12022 265254
rect 11786 264698 12022 264934
rect 11786 229018 12022 229254
rect 11786 228698 12022 228934
rect 11786 193018 12022 193254
rect 11786 192698 12022 192934
rect 11786 157018 12022 157254
rect 11786 156698 12022 156934
rect 11786 121018 12022 121254
rect 11786 120698 12022 120934
rect 11786 85018 12022 85254
rect 11786 84698 12022 84934
rect 11786 49018 12022 49254
rect 11786 48698 12022 48934
rect 11786 13018 12022 13254
rect 11786 12698 12022 12934
rect -7454 -6222 -7218 -5986
rect -7454 -6542 -7218 -6306
rect 18986 705542 19222 705778
rect 18986 705222 19222 705458
rect 18986 668218 19222 668454
rect 18986 667898 19222 668134
rect 18986 632218 19222 632454
rect 18986 631898 19222 632134
rect 18986 596218 19222 596454
rect 18986 595898 19222 596134
rect 18986 560218 19222 560454
rect 18986 559898 19222 560134
rect 18986 524218 19222 524454
rect 18986 523898 19222 524134
rect 18986 488218 19222 488454
rect 18986 487898 19222 488134
rect 18986 452218 19222 452454
rect 18986 451898 19222 452134
rect 18986 416218 19222 416454
rect 18986 415898 19222 416134
rect 18986 380218 19222 380454
rect 18986 379898 19222 380134
rect 18986 344218 19222 344454
rect 18986 343898 19222 344134
rect 18986 308218 19222 308454
rect 18986 307898 19222 308134
rect 18986 272218 19222 272454
rect 18986 271898 19222 272134
rect 18986 236218 19222 236454
rect 18986 235898 19222 236134
rect 18986 200218 19222 200454
rect 18986 199898 19222 200134
rect 18986 164218 19222 164454
rect 18986 163898 19222 164134
rect 18986 128218 19222 128454
rect 18986 127898 19222 128134
rect 18986 92218 19222 92454
rect 18986 91898 19222 92134
rect 18986 56218 19222 56454
rect 18986 55898 19222 56134
rect 18986 20218 19222 20454
rect 18986 19898 19222 20134
rect 18986 -1522 19222 -1286
rect 18986 -1842 19222 -1606
rect 22586 671818 22822 672054
rect 22586 671498 22822 671734
rect 22586 635818 22822 636054
rect 22586 635498 22822 635734
rect 22586 599818 22822 600054
rect 22586 599498 22822 599734
rect 22586 563818 22822 564054
rect 22586 563498 22822 563734
rect 22586 527818 22822 528054
rect 22586 527498 22822 527734
rect 22586 491818 22822 492054
rect 22586 491498 22822 491734
rect 22586 455818 22822 456054
rect 22586 455498 22822 455734
rect 22586 419818 22822 420054
rect 22586 419498 22822 419734
rect 22586 383818 22822 384054
rect 22586 383498 22822 383734
rect 22586 347818 22822 348054
rect 22586 347498 22822 347734
rect 22586 311818 22822 312054
rect 22586 311498 22822 311734
rect 22586 275818 22822 276054
rect 22586 275498 22822 275734
rect 22586 239818 22822 240054
rect 22586 239498 22822 239734
rect 22586 203818 22822 204054
rect 22586 203498 22822 203734
rect 22586 167818 22822 168054
rect 22586 167498 22822 167734
rect 22586 131818 22822 132054
rect 22586 131498 22822 131734
rect 22586 95818 22822 96054
rect 22586 95498 22822 95734
rect 22586 59818 22822 60054
rect 22586 59498 22822 59734
rect 22586 23818 22822 24054
rect 22586 23498 22822 23734
rect 22586 -3402 22822 -3166
rect 22586 -3722 22822 -3486
rect 26186 675418 26422 675654
rect 26186 675098 26422 675334
rect 26186 639418 26422 639654
rect 26186 639098 26422 639334
rect 26186 603418 26422 603654
rect 26186 603098 26422 603334
rect 26186 567418 26422 567654
rect 26186 567098 26422 567334
rect 26186 531418 26422 531654
rect 26186 531098 26422 531334
rect 26186 495418 26422 495654
rect 26186 495098 26422 495334
rect 26186 459418 26422 459654
rect 26186 459098 26422 459334
rect 26186 423418 26422 423654
rect 26186 423098 26422 423334
rect 26186 387418 26422 387654
rect 26186 387098 26422 387334
rect 26186 351418 26422 351654
rect 26186 351098 26422 351334
rect 26186 315418 26422 315654
rect 26186 315098 26422 315334
rect 26186 279418 26422 279654
rect 26186 279098 26422 279334
rect 26186 243418 26422 243654
rect 26186 243098 26422 243334
rect 26186 207418 26422 207654
rect 26186 207098 26422 207334
rect 26186 171418 26422 171654
rect 26186 171098 26422 171334
rect 26186 135418 26422 135654
rect 26186 135098 26422 135334
rect 26186 99418 26422 99654
rect 26186 99098 26422 99334
rect 26186 63418 26422 63654
rect 26186 63098 26422 63334
rect 26186 27418 26422 27654
rect 26186 27098 26422 27334
rect 26186 -5282 26422 -5046
rect 26186 -5602 26422 -5366
rect 47786 710242 48022 710478
rect 47786 709922 48022 710158
rect 44186 708362 44422 708598
rect 44186 708042 44422 708278
rect 40586 706482 40822 706718
rect 40586 706162 40822 706398
rect 29786 679018 30022 679254
rect 29786 678698 30022 678934
rect 29786 643018 30022 643254
rect 29786 642698 30022 642934
rect 29786 607018 30022 607254
rect 29786 606698 30022 606934
rect 29786 571018 30022 571254
rect 29786 570698 30022 570934
rect 29786 535018 30022 535254
rect 29786 534698 30022 534934
rect 29786 499018 30022 499254
rect 29786 498698 30022 498934
rect 29786 463018 30022 463254
rect 29786 462698 30022 462934
rect 29786 427018 30022 427254
rect 29786 426698 30022 426934
rect 29786 391018 30022 391254
rect 29786 390698 30022 390934
rect 29786 355018 30022 355254
rect 29786 354698 30022 354934
rect 29786 319018 30022 319254
rect 29786 318698 30022 318934
rect 29786 283018 30022 283254
rect 29786 282698 30022 282934
rect 29786 247018 30022 247254
rect 29786 246698 30022 246934
rect 29786 211018 30022 211254
rect 29786 210698 30022 210934
rect 29786 175018 30022 175254
rect 29786 174698 30022 174934
rect 29786 139018 30022 139254
rect 29786 138698 30022 138934
rect 29786 103018 30022 103254
rect 29786 102698 30022 102934
rect 29786 67018 30022 67254
rect 29786 66698 30022 66934
rect 29786 31018 30022 31254
rect 29786 30698 30022 30934
rect 11786 -6222 12022 -5986
rect 11786 -6542 12022 -6306
rect -8394 -7162 -8158 -6926
rect -8394 -7482 -8158 -7246
rect 36986 704602 37222 704838
rect 36986 704282 37222 704518
rect 36986 686218 37222 686454
rect 36986 685898 37222 686134
rect 36986 650218 37222 650454
rect 36986 649898 37222 650134
rect 36986 614218 37222 614454
rect 36986 613898 37222 614134
rect 36986 578218 37222 578454
rect 36986 577898 37222 578134
rect 36986 542218 37222 542454
rect 36986 541898 37222 542134
rect 36986 506218 37222 506454
rect 36986 505898 37222 506134
rect 36986 470218 37222 470454
rect 36986 469898 37222 470134
rect 36986 434218 37222 434454
rect 36986 433898 37222 434134
rect 36986 398218 37222 398454
rect 36986 397898 37222 398134
rect 36986 362218 37222 362454
rect 36986 361898 37222 362134
rect 36986 326218 37222 326454
rect 36986 325898 37222 326134
rect 36986 290218 37222 290454
rect 36986 289898 37222 290134
rect 36986 254218 37222 254454
rect 36986 253898 37222 254134
rect 36986 218218 37222 218454
rect 36986 217898 37222 218134
rect 36986 182218 37222 182454
rect 36986 181898 37222 182134
rect 36986 146218 37222 146454
rect 36986 145898 37222 146134
rect 36986 110218 37222 110454
rect 36986 109898 37222 110134
rect 36986 74218 37222 74454
rect 36986 73898 37222 74134
rect 36986 38218 37222 38454
rect 36986 37898 37222 38134
rect 36986 2218 37222 2454
rect 36986 1898 37222 2134
rect 36986 -582 37222 -346
rect 36986 -902 37222 -666
rect 40586 689818 40822 690054
rect 40586 689498 40822 689734
rect 40586 653818 40822 654054
rect 40586 653498 40822 653734
rect 40586 617818 40822 618054
rect 40586 617498 40822 617734
rect 40586 581818 40822 582054
rect 40586 581498 40822 581734
rect 40586 545818 40822 546054
rect 40586 545498 40822 545734
rect 40586 509818 40822 510054
rect 40586 509498 40822 509734
rect 40586 473818 40822 474054
rect 40586 473498 40822 473734
rect 40586 437818 40822 438054
rect 40586 437498 40822 437734
rect 40586 401818 40822 402054
rect 40586 401498 40822 401734
rect 40586 365818 40822 366054
rect 40586 365498 40822 365734
rect 40586 329818 40822 330054
rect 40586 329498 40822 329734
rect 40586 293818 40822 294054
rect 40586 293498 40822 293734
rect 40586 257818 40822 258054
rect 40586 257498 40822 257734
rect 40586 221818 40822 222054
rect 40586 221498 40822 221734
rect 40586 185818 40822 186054
rect 40586 185498 40822 185734
rect 40586 149818 40822 150054
rect 40586 149498 40822 149734
rect 40586 113818 40822 114054
rect 40586 113498 40822 113734
rect 40586 77818 40822 78054
rect 40586 77498 40822 77734
rect 40586 41818 40822 42054
rect 40586 41498 40822 41734
rect 40586 5818 40822 6054
rect 40586 5498 40822 5734
rect 40586 -2462 40822 -2226
rect 40586 -2782 40822 -2546
rect 44186 693418 44422 693654
rect 44186 693098 44422 693334
rect 44186 657418 44422 657654
rect 44186 657098 44422 657334
rect 44186 621418 44422 621654
rect 44186 621098 44422 621334
rect 44186 585418 44422 585654
rect 44186 585098 44422 585334
rect 44186 549418 44422 549654
rect 44186 549098 44422 549334
rect 44186 513418 44422 513654
rect 44186 513098 44422 513334
rect 44186 477418 44422 477654
rect 44186 477098 44422 477334
rect 44186 441418 44422 441654
rect 44186 441098 44422 441334
rect 44186 405418 44422 405654
rect 44186 405098 44422 405334
rect 44186 369418 44422 369654
rect 44186 369098 44422 369334
rect 44186 333418 44422 333654
rect 44186 333098 44422 333334
rect 44186 297418 44422 297654
rect 44186 297098 44422 297334
rect 44186 261418 44422 261654
rect 44186 261098 44422 261334
rect 44186 225418 44422 225654
rect 44186 225098 44422 225334
rect 44186 189418 44422 189654
rect 44186 189098 44422 189334
rect 44186 153418 44422 153654
rect 44186 153098 44422 153334
rect 44186 117418 44422 117654
rect 44186 117098 44422 117334
rect 44186 81418 44422 81654
rect 44186 81098 44422 81334
rect 44186 45418 44422 45654
rect 44186 45098 44422 45334
rect 44186 9418 44422 9654
rect 44186 9098 44422 9334
rect 44186 -4342 44422 -4106
rect 44186 -4662 44422 -4426
rect 65786 711182 66022 711418
rect 65786 710862 66022 711098
rect 62186 709302 62422 709538
rect 62186 708982 62422 709218
rect 58586 707422 58822 707658
rect 58586 707102 58822 707338
rect 47786 697018 48022 697254
rect 47786 696698 48022 696934
rect 47786 661018 48022 661254
rect 47786 660698 48022 660934
rect 47786 625018 48022 625254
rect 47786 624698 48022 624934
rect 47786 589018 48022 589254
rect 47786 588698 48022 588934
rect 47786 553018 48022 553254
rect 47786 552698 48022 552934
rect 47786 517018 48022 517254
rect 47786 516698 48022 516934
rect 47786 481018 48022 481254
rect 47786 480698 48022 480934
rect 47786 445018 48022 445254
rect 47786 444698 48022 444934
rect 47786 409018 48022 409254
rect 47786 408698 48022 408934
rect 47786 373018 48022 373254
rect 47786 372698 48022 372934
rect 47786 337018 48022 337254
rect 47786 336698 48022 336934
rect 47786 301018 48022 301254
rect 47786 300698 48022 300934
rect 47786 265018 48022 265254
rect 47786 264698 48022 264934
rect 47786 229018 48022 229254
rect 47786 228698 48022 228934
rect 47786 193018 48022 193254
rect 47786 192698 48022 192934
rect 47786 157018 48022 157254
rect 47786 156698 48022 156934
rect 47786 121018 48022 121254
rect 47786 120698 48022 120934
rect 47786 85018 48022 85254
rect 47786 84698 48022 84934
rect 47786 49018 48022 49254
rect 47786 48698 48022 48934
rect 47786 13018 48022 13254
rect 47786 12698 48022 12934
rect 29786 -7162 30022 -6926
rect 29786 -7482 30022 -7246
rect 54986 705542 55222 705778
rect 54986 705222 55222 705458
rect 54986 668218 55222 668454
rect 54986 667898 55222 668134
rect 54986 632218 55222 632454
rect 54986 631898 55222 632134
rect 54986 596218 55222 596454
rect 54986 595898 55222 596134
rect 54986 560218 55222 560454
rect 54986 559898 55222 560134
rect 54986 524218 55222 524454
rect 54986 523898 55222 524134
rect 54986 488218 55222 488454
rect 54986 487898 55222 488134
rect 54986 452218 55222 452454
rect 54986 451898 55222 452134
rect 54986 416218 55222 416454
rect 54986 415898 55222 416134
rect 58586 671818 58822 672054
rect 58586 671498 58822 671734
rect 62186 675418 62422 675654
rect 62186 675098 62422 675334
rect 83786 710242 84022 710478
rect 83786 709922 84022 710158
rect 80186 708362 80422 708598
rect 80186 708042 80422 708278
rect 76586 706482 76822 706718
rect 76586 706162 76822 706398
rect 65786 679018 66022 679254
rect 65786 678698 66022 678934
rect 72986 704602 73222 704838
rect 72986 704282 73222 704518
rect 72986 686218 73222 686454
rect 72986 685898 73222 686134
rect 76586 689818 76822 690054
rect 76586 689498 76822 689734
rect 80186 693418 80422 693654
rect 80186 693098 80422 693334
rect 80186 657418 80422 657654
rect 80186 657098 80422 657334
rect 101786 711182 102022 711418
rect 101786 710862 102022 711098
rect 98186 709302 98422 709538
rect 98186 708982 98422 709218
rect 94586 707422 94822 707658
rect 94586 707102 94822 707338
rect 83786 697018 84022 697254
rect 83786 696698 84022 696934
rect 83786 661018 84022 661254
rect 83786 660698 84022 660934
rect 90986 705542 91222 705778
rect 90986 705222 91222 705458
rect 90986 668218 91222 668454
rect 90986 667898 91222 668134
rect 94586 671818 94822 672054
rect 94586 671498 94822 671734
rect 98186 675418 98422 675654
rect 98186 675098 98422 675334
rect 119786 710242 120022 710478
rect 119786 709922 120022 710158
rect 116186 708362 116422 708598
rect 116186 708042 116422 708278
rect 112586 706482 112822 706718
rect 112586 706162 112822 706398
rect 101786 679018 102022 679254
rect 101786 678698 102022 678934
rect 108986 704602 109222 704838
rect 108986 704282 109222 704518
rect 108986 686218 109222 686454
rect 108986 685898 109222 686134
rect 112586 689818 112822 690054
rect 112586 689498 112822 689734
rect 116186 693418 116422 693654
rect 116186 693098 116422 693334
rect 116186 657418 116422 657654
rect 116186 657098 116422 657334
rect 137786 711182 138022 711418
rect 137786 710862 138022 711098
rect 134186 709302 134422 709538
rect 134186 708982 134422 709218
rect 130586 707422 130822 707658
rect 130586 707102 130822 707338
rect 119786 697018 120022 697254
rect 119786 696698 120022 696934
rect 119786 661018 120022 661254
rect 119786 660698 120022 660934
rect 126986 705542 127222 705778
rect 126986 705222 127222 705458
rect 126986 668218 127222 668454
rect 126986 667898 127222 668134
rect 130586 671818 130822 672054
rect 130586 671498 130822 671734
rect 134186 675418 134422 675654
rect 134186 675098 134422 675334
rect 155786 710242 156022 710478
rect 155786 709922 156022 710158
rect 152186 708362 152422 708598
rect 152186 708042 152422 708278
rect 148586 706482 148822 706718
rect 148586 706162 148822 706398
rect 137786 679018 138022 679254
rect 137786 678698 138022 678934
rect 144986 704602 145222 704838
rect 144986 704282 145222 704518
rect 144986 686218 145222 686454
rect 144986 685898 145222 686134
rect 144986 650218 145222 650454
rect 144986 649898 145222 650134
rect 136982 643018 137218 643254
rect 136982 642698 137218 642934
rect 136982 639418 137218 639654
rect 136982 639098 137218 639334
rect 136982 635818 137218 636054
rect 136982 635498 137218 635734
rect 136982 632218 137218 632454
rect 136982 631898 137218 632134
rect 136536 625018 136772 625254
rect 136536 624698 136772 624934
rect 136536 621418 136772 621654
rect 136536 621098 136772 621334
rect 136536 617818 136772 618054
rect 136536 617498 136772 617734
rect 136536 614218 136772 614454
rect 136536 613898 136772 614134
rect 144986 614218 145222 614454
rect 144986 613898 145222 614134
rect 136982 607018 137218 607254
rect 136982 606698 137218 606934
rect 136982 603418 137218 603654
rect 136982 603098 137218 603334
rect 136982 599818 137218 600054
rect 136982 599498 137218 599734
rect 136982 596218 137218 596454
rect 136982 595898 137218 596134
rect 136536 589018 136772 589254
rect 136536 588698 136772 588934
rect 136536 585418 136772 585654
rect 136536 585098 136772 585334
rect 136536 581818 136772 582054
rect 136536 581498 136772 581734
rect 136536 578218 136772 578454
rect 136536 577898 136772 578134
rect 144986 578218 145222 578454
rect 144986 577898 145222 578134
rect 136982 571018 137218 571254
rect 136982 570698 137218 570934
rect 136982 567418 137218 567654
rect 136982 567098 137218 567334
rect 136982 563818 137218 564054
rect 136982 563498 137218 563734
rect 76586 545818 76822 546054
rect 76586 545498 76822 545734
rect 80186 549418 80422 549654
rect 80186 549098 80422 549334
rect 83786 553018 84022 553254
rect 83786 552698 84022 552934
rect 112586 545818 112822 546054
rect 112586 545498 112822 545734
rect 116186 549418 116422 549654
rect 116186 549098 116422 549334
rect 119786 553018 120022 553254
rect 119786 552698 120022 552934
rect 148586 689818 148822 690054
rect 148586 689498 148822 689734
rect 148586 653818 148822 654054
rect 148586 653498 148822 653734
rect 148586 617818 148822 618054
rect 148586 617498 148822 617734
rect 148586 581818 148822 582054
rect 148586 581498 148822 581734
rect 148586 545818 148822 546054
rect 148586 545498 148822 545734
rect 152186 693418 152422 693654
rect 152186 693098 152422 693334
rect 152186 657418 152422 657654
rect 152186 657098 152422 657334
rect 152186 621418 152422 621654
rect 152186 621098 152422 621334
rect 152186 585418 152422 585654
rect 152186 585098 152422 585334
rect 152186 549418 152422 549654
rect 152186 549098 152422 549334
rect 173786 711182 174022 711418
rect 173786 710862 174022 711098
rect 170186 709302 170422 709538
rect 170186 708982 170422 709218
rect 166586 707422 166822 707658
rect 166586 707102 166822 707338
rect 155786 697018 156022 697254
rect 155786 696698 156022 696934
rect 155786 661018 156022 661254
rect 155786 660698 156022 660934
rect 155786 625018 156022 625254
rect 155786 624698 156022 624934
rect 155786 589018 156022 589254
rect 155786 588698 156022 588934
rect 155786 553018 156022 553254
rect 155786 552698 156022 552934
rect 162986 705542 163222 705778
rect 162986 705222 163222 705458
rect 162986 668218 163222 668454
rect 162986 667898 163222 668134
rect 162986 632218 163222 632454
rect 162986 631898 163222 632134
rect 162986 596218 163222 596454
rect 162986 595898 163222 596134
rect 162986 560218 163222 560454
rect 162986 559898 163222 560134
rect 166586 671818 166822 672054
rect 166586 671498 166822 671734
rect 166586 635818 166822 636054
rect 166586 635498 166822 635734
rect 166586 599818 166822 600054
rect 166586 599498 166822 599734
rect 166586 563818 166822 564054
rect 166586 563498 166822 563734
rect 170186 675418 170422 675654
rect 170186 675098 170422 675334
rect 170186 639418 170422 639654
rect 170186 639098 170422 639334
rect 170186 603418 170422 603654
rect 170186 603098 170422 603334
rect 170186 567418 170422 567654
rect 170186 567098 170422 567334
rect 191786 710242 192022 710478
rect 191786 709922 192022 710158
rect 188186 708362 188422 708598
rect 188186 708042 188422 708278
rect 184586 706482 184822 706718
rect 184586 706162 184822 706398
rect 173786 679018 174022 679254
rect 173786 678698 174022 678934
rect 173786 643018 174022 643254
rect 173786 642698 174022 642934
rect 173786 607018 174022 607254
rect 173786 606698 174022 606934
rect 173786 571018 174022 571254
rect 173786 570698 174022 570934
rect 180986 704602 181222 704838
rect 180986 704282 181222 704518
rect 184586 689818 184822 690054
rect 184586 689498 184822 689734
rect 180986 686218 181222 686454
rect 180986 685898 181222 686134
rect 180986 650218 181222 650454
rect 180986 649898 181222 650134
rect 180986 614218 181222 614454
rect 180986 613898 181222 614134
rect 180986 578218 181222 578454
rect 180986 577898 181222 578134
rect 188186 693418 188422 693654
rect 188186 693098 188422 693334
rect 188186 657418 188422 657654
rect 188186 657098 188422 657334
rect 209786 711182 210022 711418
rect 209786 710862 210022 711098
rect 206186 709302 206422 709538
rect 206186 708982 206422 709218
rect 202586 707422 202822 707658
rect 202586 707102 202822 707338
rect 191786 697018 192022 697254
rect 191786 696698 192022 696934
rect 191786 661018 192022 661254
rect 191786 660698 192022 660934
rect 198986 705542 199222 705778
rect 198986 705222 199222 705458
rect 198986 668218 199222 668454
rect 198986 667898 199222 668134
rect 202586 671818 202822 672054
rect 202586 671498 202822 671734
rect 206186 675418 206422 675654
rect 206186 675098 206422 675334
rect 227786 710242 228022 710478
rect 227786 709922 228022 710158
rect 224186 708362 224422 708598
rect 224186 708042 224422 708278
rect 220586 706482 220822 706718
rect 220586 706162 220822 706398
rect 209786 679018 210022 679254
rect 209786 678698 210022 678934
rect 216986 704602 217222 704838
rect 216986 704282 217222 704518
rect 216986 686218 217222 686454
rect 216986 685898 217222 686134
rect 220586 689818 220822 690054
rect 220586 689498 220822 689734
rect 224186 693418 224422 693654
rect 224186 693098 224422 693334
rect 224186 657418 224422 657654
rect 224186 657098 224422 657334
rect 245786 711182 246022 711418
rect 245786 710862 246022 711098
rect 242186 709302 242422 709538
rect 242186 708982 242422 709218
rect 238586 707422 238822 707658
rect 238586 707102 238822 707338
rect 227786 697018 228022 697254
rect 227786 696698 228022 696934
rect 227786 661018 228022 661254
rect 227786 660698 228022 660934
rect 234986 705542 235222 705778
rect 234986 705222 235222 705458
rect 234986 668218 235222 668454
rect 234986 667898 235222 668134
rect 238586 671818 238822 672054
rect 238586 671498 238822 671734
rect 242186 675418 242422 675654
rect 242186 675098 242422 675334
rect 263786 710242 264022 710478
rect 263786 709922 264022 710158
rect 260186 708362 260422 708598
rect 260186 708042 260422 708278
rect 256586 706482 256822 706718
rect 256586 706162 256822 706398
rect 245786 679018 246022 679254
rect 245786 678698 246022 678934
rect 252986 704602 253222 704838
rect 252986 704282 253222 704518
rect 252986 686218 253222 686454
rect 252986 685898 253222 686134
rect 256586 689818 256822 690054
rect 256586 689498 256822 689734
rect 260186 693418 260422 693654
rect 260186 693098 260422 693334
rect 260186 657418 260422 657654
rect 260186 657098 260422 657334
rect 281786 711182 282022 711418
rect 281786 710862 282022 711098
rect 278186 709302 278422 709538
rect 278186 708982 278422 709218
rect 274586 707422 274822 707658
rect 274586 707102 274822 707338
rect 263786 697018 264022 697254
rect 263786 696698 264022 696934
rect 263786 661018 264022 661254
rect 263786 660698 264022 660934
rect 270986 705542 271222 705778
rect 270986 705222 271222 705458
rect 270986 668218 271222 668454
rect 270986 667898 271222 668134
rect 184586 653818 184822 654054
rect 184586 653498 184822 653734
rect 266982 643018 267218 643254
rect 266982 642698 267218 642934
rect 266982 639418 267218 639654
rect 266982 639098 267218 639334
rect 266982 635818 267218 636054
rect 266982 635498 267218 635734
rect 266982 632218 267218 632454
rect 266982 631898 267218 632134
rect 270986 632218 271222 632454
rect 270986 631898 271222 632134
rect 266536 625018 266772 625254
rect 266536 624698 266772 624934
rect 266536 621418 266772 621654
rect 266536 621098 266772 621334
rect 184586 617818 184822 618054
rect 184586 617498 184822 617734
rect 266536 617818 266772 618054
rect 266536 617498 266772 617734
rect 266536 614218 266772 614454
rect 266536 613898 266772 614134
rect 266982 607018 267218 607254
rect 266982 606698 267218 606934
rect 266982 603418 267218 603654
rect 266982 603098 267218 603334
rect 266982 599818 267218 600054
rect 266982 599498 267218 599734
rect 266982 596218 267218 596454
rect 266982 595898 267218 596134
rect 270986 596218 271222 596454
rect 270986 595898 271222 596134
rect 266536 589018 266772 589254
rect 266536 588698 266772 588934
rect 266536 585418 266772 585654
rect 266536 585098 266772 585334
rect 184586 581818 184822 582054
rect 184586 581498 184822 581734
rect 266536 581818 266772 582054
rect 266536 581498 266772 581734
rect 266536 578218 266772 578454
rect 266536 577898 266772 578134
rect 266982 571018 267218 571254
rect 266982 570698 267218 570934
rect 266982 567418 267218 567654
rect 266982 567098 267218 567334
rect 266982 563818 267218 564054
rect 266982 563498 267218 563734
rect 270986 560218 271222 560454
rect 270986 559898 271222 560134
rect 184586 545818 184822 546054
rect 184586 545498 184822 545734
rect 188186 549418 188422 549654
rect 188186 549098 188422 549334
rect 191786 553018 192022 553254
rect 191786 552698 192022 552934
rect 220586 545818 220822 546054
rect 220586 545498 220822 545734
rect 224186 549418 224422 549654
rect 224186 549098 224422 549334
rect 227786 553018 228022 553254
rect 227786 552698 228022 552934
rect 256586 545818 256822 546054
rect 256586 545498 256822 545734
rect 260186 549418 260422 549654
rect 260186 549098 260422 549334
rect 263786 553018 264022 553254
rect 263786 552698 264022 552934
rect 274586 671818 274822 672054
rect 274586 671498 274822 671734
rect 274586 635818 274822 636054
rect 274586 635498 274822 635734
rect 274586 599818 274822 600054
rect 274586 599498 274822 599734
rect 274586 563818 274822 564054
rect 274586 563498 274822 563734
rect 278186 675418 278422 675654
rect 278186 675098 278422 675334
rect 278186 639418 278422 639654
rect 278186 639098 278422 639334
rect 278186 603418 278422 603654
rect 278186 603098 278422 603334
rect 278186 567418 278422 567654
rect 278186 567098 278422 567334
rect 299786 710242 300022 710478
rect 299786 709922 300022 710158
rect 296186 708362 296422 708598
rect 296186 708042 296422 708278
rect 292586 706482 292822 706718
rect 292586 706162 292822 706398
rect 281786 679018 282022 679254
rect 281786 678698 282022 678934
rect 281786 643018 282022 643254
rect 281786 642698 282022 642934
rect 281786 607018 282022 607254
rect 281786 606698 282022 606934
rect 281786 571018 282022 571254
rect 281786 570698 282022 570934
rect 288986 704602 289222 704838
rect 288986 704282 289222 704518
rect 288986 686218 289222 686454
rect 288986 685898 289222 686134
rect 288986 650218 289222 650454
rect 288986 649898 289222 650134
rect 288986 614218 289222 614454
rect 288986 613898 289222 614134
rect 288986 578218 289222 578454
rect 288986 577898 289222 578134
rect 79610 535018 79846 535254
rect 79610 534698 79846 534934
rect 79610 531418 79846 531654
rect 79610 531098 79846 531334
rect 79610 527818 79846 528054
rect 79610 527498 79846 527734
rect 79610 524218 79846 524454
rect 79610 523898 79846 524134
rect 64250 517018 64486 517254
rect 64250 516698 64486 516934
rect 64250 513418 64486 513654
rect 64250 513098 64486 513334
rect 64250 509818 64486 510054
rect 64250 509498 64486 509734
rect 64250 506218 64486 506454
rect 64250 505898 64486 506134
rect 79610 499018 79846 499254
rect 79610 498698 79846 498934
rect 79610 495418 79846 495654
rect 79610 495098 79846 495334
rect 79610 491818 79846 492054
rect 79610 491498 79846 491734
rect 79610 488218 79846 488454
rect 79610 487898 79846 488134
rect 64250 481018 64486 481254
rect 64250 480698 64486 480934
rect 64250 477418 64486 477654
rect 64250 477098 64486 477334
rect 64250 473818 64486 474054
rect 64250 473498 64486 473734
rect 64250 470218 64486 470454
rect 64250 469898 64486 470134
rect 79610 463018 79846 463254
rect 79610 462698 79846 462934
rect 79610 459418 79846 459654
rect 79610 459098 79846 459334
rect 79610 455818 79846 456054
rect 79610 455498 79846 455734
rect 79610 452218 79846 452454
rect 79610 451898 79846 452134
rect 64250 445018 64486 445254
rect 64250 444698 64486 444934
rect 64250 441418 64486 441654
rect 64250 441098 64486 441334
rect 64250 437818 64486 438054
rect 64250 437498 64486 437734
rect 64250 434218 64486 434454
rect 64250 433898 64486 434134
rect 79610 427018 79846 427254
rect 79610 426698 79846 426934
rect 79610 423418 79846 423654
rect 79610 423098 79846 423334
rect 79610 419818 79846 420054
rect 79610 419498 79846 419734
rect 79610 416218 79846 416454
rect 79610 415898 79846 416134
rect 64250 409018 64486 409254
rect 64250 408698 64486 408934
rect 64250 405418 64486 405654
rect 64250 405098 64486 405334
rect 64250 401818 64486 402054
rect 64250 401498 64486 401734
rect 64250 398218 64486 398454
rect 64250 397898 64486 398134
rect 79610 391018 79846 391254
rect 79610 390698 79846 390934
rect 79610 387418 79846 387654
rect 79610 387098 79846 387334
rect 79610 383818 79846 384054
rect 79610 383498 79846 383734
rect 54986 380218 55222 380454
rect 54986 379898 55222 380134
rect 79610 380218 79846 380454
rect 79610 379898 79846 380134
rect 54986 344218 55222 344454
rect 54986 343898 55222 344134
rect 54986 308218 55222 308454
rect 54986 307898 55222 308134
rect 54986 272218 55222 272454
rect 54986 271898 55222 272134
rect 54986 236218 55222 236454
rect 54986 235898 55222 236134
rect 54986 200218 55222 200454
rect 54986 199898 55222 200134
rect 64250 373018 64486 373254
rect 64250 372698 64486 372934
rect 64250 369418 64486 369654
rect 64250 369098 64486 369334
rect 64250 365818 64486 366054
rect 64250 365498 64486 365734
rect 64250 362218 64486 362454
rect 64250 361898 64486 362134
rect 79610 355018 79846 355254
rect 79610 354698 79846 354934
rect 79610 351418 79846 351654
rect 79610 351098 79846 351334
rect 79610 347818 79846 348054
rect 79610 347498 79846 347734
rect 79610 344218 79846 344454
rect 79610 343898 79846 344134
rect 64250 337018 64486 337254
rect 64250 336698 64486 336934
rect 64250 333418 64486 333654
rect 64250 333098 64486 333334
rect 54986 164218 55222 164454
rect 54986 163898 55222 164134
rect 54986 128218 55222 128454
rect 54986 127898 55222 128134
rect 54986 92218 55222 92454
rect 54986 91898 55222 92134
rect 64250 329818 64486 330054
rect 64250 329498 64486 329734
rect 64250 326218 64486 326454
rect 64250 325898 64486 326134
rect 288986 542218 289222 542454
rect 288986 541898 289222 542134
rect 288986 506218 289222 506454
rect 288986 505898 289222 506134
rect 288986 470218 289222 470454
rect 288986 469898 289222 470134
rect 288986 434218 289222 434454
rect 288986 433898 289222 434134
rect 288986 398218 289222 398454
rect 288986 397898 289222 398134
rect 288986 362218 289222 362454
rect 288986 361898 289222 362134
rect 288986 326218 289222 326454
rect 288986 325898 289222 326134
rect 58586 311818 58822 312054
rect 58586 311498 58822 311734
rect 58586 275818 58822 276054
rect 58586 275498 58822 275734
rect 58586 239818 58822 240054
rect 58586 239498 58822 239734
rect 58586 203818 58822 204054
rect 58586 203498 58822 203734
rect 58586 167818 58822 168054
rect 58586 167498 58822 167734
rect 58586 131818 58822 132054
rect 58586 131498 58822 131734
rect 58586 95818 58822 96054
rect 58586 95498 58822 95734
rect 54986 56218 55222 56454
rect 54986 55898 55222 56134
rect 54986 20218 55222 20454
rect 54986 19898 55222 20134
rect 54986 -1522 55222 -1286
rect 54986 -1842 55222 -1606
rect 58586 59818 58822 60054
rect 58586 59498 58822 59734
rect 58586 23818 58822 24054
rect 58586 23498 58822 23734
rect 58586 -3402 58822 -3166
rect 58586 -3722 58822 -3486
rect 62186 315418 62422 315654
rect 62186 315098 62422 315334
rect 62186 279418 62422 279654
rect 62186 279098 62422 279334
rect 62186 243418 62422 243654
rect 62186 243098 62422 243334
rect 62186 207418 62422 207654
rect 62186 207098 62422 207334
rect 62186 171418 62422 171654
rect 62186 171098 62422 171334
rect 62186 135418 62422 135654
rect 62186 135098 62422 135334
rect 62186 99418 62422 99654
rect 62186 99098 62422 99334
rect 62186 63418 62422 63654
rect 62186 63098 62422 63334
rect 62186 27418 62422 27654
rect 62186 27098 62422 27334
rect 62186 -5282 62422 -5046
rect 62186 -5602 62422 -5366
rect 65786 283018 66022 283254
rect 65786 282698 66022 282934
rect 65786 247018 66022 247254
rect 65786 246698 66022 246934
rect 65786 211018 66022 211254
rect 65786 210698 66022 210934
rect 65786 175018 66022 175254
rect 65786 174698 66022 174934
rect 65786 139018 66022 139254
rect 65786 138698 66022 138934
rect 65786 103018 66022 103254
rect 65786 102698 66022 102934
rect 65786 67018 66022 67254
rect 65786 66698 66022 66934
rect 65786 31018 66022 31254
rect 65786 30698 66022 30934
rect 47786 -6222 48022 -5986
rect 47786 -6542 48022 -6306
rect 72986 290218 73222 290454
rect 72986 289898 73222 290134
rect 72986 254218 73222 254454
rect 72986 253898 73222 254134
rect 72986 218218 73222 218454
rect 72986 217898 73222 218134
rect 72986 182218 73222 182454
rect 72986 181898 73222 182134
rect 72986 146218 73222 146454
rect 72986 145898 73222 146134
rect 72986 110218 73222 110454
rect 72986 109898 73222 110134
rect 72986 74218 73222 74454
rect 72986 73898 73222 74134
rect 72986 38218 73222 38454
rect 72986 37898 73222 38134
rect 72986 2218 73222 2454
rect 72986 1898 73222 2134
rect 72986 -582 73222 -346
rect 72986 -902 73222 -666
rect 76586 293818 76822 294054
rect 76586 293498 76822 293734
rect 76586 257818 76822 258054
rect 76586 257498 76822 257734
rect 76586 221818 76822 222054
rect 76586 221498 76822 221734
rect 76586 185818 76822 186054
rect 76586 185498 76822 185734
rect 76586 149818 76822 150054
rect 76586 149498 76822 149734
rect 76586 113818 76822 114054
rect 76586 113498 76822 113734
rect 76586 77818 76822 78054
rect 76586 77498 76822 77734
rect 76586 41818 76822 42054
rect 76586 41498 76822 41734
rect 76586 5818 76822 6054
rect 76586 5498 76822 5734
rect 76586 -2462 76822 -2226
rect 76586 -2782 76822 -2546
rect 80186 297418 80422 297654
rect 80186 297098 80422 297334
rect 80186 261418 80422 261654
rect 80186 261098 80422 261334
rect 80186 225418 80422 225654
rect 80186 225098 80422 225334
rect 80186 189418 80422 189654
rect 80186 189098 80422 189334
rect 80186 153418 80422 153654
rect 80186 153098 80422 153334
rect 80186 117418 80422 117654
rect 80186 117098 80422 117334
rect 80186 81418 80422 81654
rect 80186 81098 80422 81334
rect 80186 45418 80422 45654
rect 80186 45098 80422 45334
rect 80186 9418 80422 9654
rect 80186 9098 80422 9334
rect 80186 -4342 80422 -4106
rect 80186 -4662 80422 -4426
rect 83786 301018 84022 301254
rect 83786 300698 84022 300934
rect 83786 265018 84022 265254
rect 83786 264698 84022 264934
rect 90986 308218 91222 308454
rect 90986 307898 91222 308134
rect 90986 272218 91222 272454
rect 90986 271898 91222 272134
rect 83786 229018 84022 229254
rect 83786 228698 84022 228934
rect 90986 236218 91222 236454
rect 90986 235898 91222 236134
rect 83786 193018 84022 193254
rect 83786 192698 84022 192934
rect 83786 157018 84022 157254
rect 83786 156698 84022 156934
rect 83786 121018 84022 121254
rect 83786 120698 84022 120934
rect 83786 85018 84022 85254
rect 83786 84698 84022 84934
rect 83786 49018 84022 49254
rect 83786 48698 84022 48934
rect 90986 200218 91222 200454
rect 90986 199898 91222 200134
rect 90986 164218 91222 164454
rect 90986 163898 91222 164134
rect 90986 128218 91222 128454
rect 90986 127898 91222 128134
rect 90986 92218 91222 92454
rect 90986 91898 91222 92134
rect 90986 56218 91222 56454
rect 90986 55898 91222 56134
rect 83786 13018 84022 13254
rect 83786 12698 84022 12934
rect 65786 -7162 66022 -6926
rect 65786 -7482 66022 -7246
rect 90986 20218 91222 20454
rect 90986 19898 91222 20134
rect 90986 -1522 91222 -1286
rect 90986 -1842 91222 -1606
rect 94586 311818 94822 312054
rect 94586 311498 94822 311734
rect 94586 275818 94822 276054
rect 94586 275498 94822 275734
rect 98186 315418 98422 315654
rect 98186 315098 98422 315334
rect 98186 279418 98422 279654
rect 98186 279098 98422 279334
rect 94586 239818 94822 240054
rect 94586 239498 94822 239734
rect 98186 243418 98422 243654
rect 98186 243098 98422 243334
rect 94586 203818 94822 204054
rect 94586 203498 94822 203734
rect 98186 207418 98422 207654
rect 98186 207098 98422 207334
rect 94586 167818 94822 168054
rect 94586 167498 94822 167734
rect 94586 131818 94822 132054
rect 94586 131498 94822 131734
rect 94586 95818 94822 96054
rect 94586 95498 94822 95734
rect 94586 59818 94822 60054
rect 94586 59498 94822 59734
rect 94586 23818 94822 24054
rect 94586 23498 94822 23734
rect 94586 -3402 94822 -3166
rect 94586 -3722 94822 -3486
rect 98186 171418 98422 171654
rect 98186 171098 98422 171334
rect 98186 135418 98422 135654
rect 98186 135098 98422 135334
rect 98186 99418 98422 99654
rect 98186 99098 98422 99334
rect 98186 63418 98422 63654
rect 98186 63098 98422 63334
rect 98186 27418 98422 27654
rect 98186 27098 98422 27334
rect 98186 -5282 98422 -5046
rect 98186 -5602 98422 -5366
rect 101786 283018 102022 283254
rect 101786 282698 102022 282934
rect 108986 290218 109222 290454
rect 108986 289898 109222 290134
rect 101786 247018 102022 247254
rect 101786 246698 102022 246934
rect 108986 254218 109222 254454
rect 108986 253898 109222 254134
rect 101786 211018 102022 211254
rect 101786 210698 102022 210934
rect 108986 218218 109222 218454
rect 108986 217898 109222 218134
rect 108986 182218 109222 182454
rect 108986 181898 109222 182134
rect 101786 175018 102022 175254
rect 101786 174698 102022 174934
rect 101786 139018 102022 139254
rect 101786 138698 102022 138934
rect 101786 103018 102022 103254
rect 101786 102698 102022 102934
rect 101786 67018 102022 67254
rect 101786 66698 102022 66934
rect 101786 31018 102022 31254
rect 101786 30698 102022 30934
rect 83786 -6222 84022 -5986
rect 83786 -6542 84022 -6306
rect 108986 146218 109222 146454
rect 108986 145898 109222 146134
rect 108986 110218 109222 110454
rect 108986 109898 109222 110134
rect 108986 74218 109222 74454
rect 108986 73898 109222 74134
rect 108986 38218 109222 38454
rect 108986 37898 109222 38134
rect 108986 2218 109222 2454
rect 108986 1898 109222 2134
rect 108986 -582 109222 -346
rect 108986 -902 109222 -666
rect 112586 293818 112822 294054
rect 112586 293498 112822 293734
rect 112586 257818 112822 258054
rect 112586 257498 112822 257734
rect 112586 221818 112822 222054
rect 112586 221498 112822 221734
rect 112586 185818 112822 186054
rect 112586 185498 112822 185734
rect 112586 149818 112822 150054
rect 112586 149498 112822 149734
rect 112586 113818 112822 114054
rect 112586 113498 112822 113734
rect 112586 77818 112822 78054
rect 112586 77498 112822 77734
rect 112586 41818 112822 42054
rect 112586 41498 112822 41734
rect 112586 5818 112822 6054
rect 112586 5498 112822 5734
rect 112586 -2462 112822 -2226
rect 112586 -2782 112822 -2546
rect 116186 297418 116422 297654
rect 116186 297098 116422 297334
rect 116186 261418 116422 261654
rect 116186 261098 116422 261334
rect 116186 225418 116422 225654
rect 116186 225098 116422 225334
rect 116186 189418 116422 189654
rect 116186 189098 116422 189334
rect 116186 153418 116422 153654
rect 116186 153098 116422 153334
rect 116186 117418 116422 117654
rect 116186 117098 116422 117334
rect 116186 81418 116422 81654
rect 116186 81098 116422 81334
rect 116186 45418 116422 45654
rect 116186 45098 116422 45334
rect 116186 9418 116422 9654
rect 116186 9098 116422 9334
rect 116186 -4342 116422 -4106
rect 116186 -4662 116422 -4426
rect 119786 301018 120022 301254
rect 119786 300698 120022 300934
rect 119786 265018 120022 265254
rect 119786 264698 120022 264934
rect 126986 308218 127222 308454
rect 126986 307898 127222 308134
rect 126986 272218 127222 272454
rect 126986 271898 127222 272134
rect 119786 229018 120022 229254
rect 119786 228698 120022 228934
rect 126986 236218 127222 236454
rect 126986 235898 127222 236134
rect 119786 193018 120022 193254
rect 119786 192698 120022 192934
rect 126986 200218 127222 200454
rect 126986 199898 127222 200134
rect 119786 157018 120022 157254
rect 119786 156698 120022 156934
rect 119786 121018 120022 121254
rect 119786 120698 120022 120934
rect 119786 85018 120022 85254
rect 119786 84698 120022 84934
rect 126986 164218 127222 164454
rect 126986 163898 127222 164134
rect 126986 128218 127222 128454
rect 126986 127898 127222 128134
rect 126986 92218 127222 92454
rect 126986 91898 127222 92134
rect 119786 49018 120022 49254
rect 119786 48698 120022 48934
rect 119786 13018 120022 13254
rect 119786 12698 120022 12934
rect 101786 -7162 102022 -6926
rect 101786 -7482 102022 -7246
rect 126986 56218 127222 56454
rect 126986 55898 127222 56134
rect 126986 20218 127222 20454
rect 126986 19898 127222 20134
rect 126986 -1522 127222 -1286
rect 126986 -1842 127222 -1606
rect 130586 311818 130822 312054
rect 130586 311498 130822 311734
rect 130586 275818 130822 276054
rect 130586 275498 130822 275734
rect 130586 239818 130822 240054
rect 130586 239498 130822 239734
rect 130586 203818 130822 204054
rect 130586 203498 130822 203734
rect 130586 167818 130822 168054
rect 130586 167498 130822 167734
rect 130586 131818 130822 132054
rect 130586 131498 130822 131734
rect 130586 95818 130822 96054
rect 130586 95498 130822 95734
rect 130586 59818 130822 60054
rect 130586 59498 130822 59734
rect 130586 23818 130822 24054
rect 130586 23498 130822 23734
rect 130586 -3402 130822 -3166
rect 130586 -3722 130822 -3486
rect 134186 315418 134422 315654
rect 134186 315098 134422 315334
rect 134186 279418 134422 279654
rect 134186 279098 134422 279334
rect 134186 243418 134422 243654
rect 134186 243098 134422 243334
rect 134186 207418 134422 207654
rect 134186 207098 134422 207334
rect 134186 171418 134422 171654
rect 134186 171098 134422 171334
rect 134186 135418 134422 135654
rect 134186 135098 134422 135334
rect 134186 99418 134422 99654
rect 134186 99098 134422 99334
rect 134186 63418 134422 63654
rect 134186 63098 134422 63334
rect 134186 27418 134422 27654
rect 134186 27098 134422 27334
rect 134186 -5282 134422 -5046
rect 134186 -5602 134422 -5366
rect 137786 283018 138022 283254
rect 137786 282698 138022 282934
rect 137786 247018 138022 247254
rect 137786 246698 138022 246934
rect 137786 211018 138022 211254
rect 137786 210698 138022 210934
rect 137786 175018 138022 175254
rect 137786 174698 138022 174934
rect 137786 139018 138022 139254
rect 137786 138698 138022 138934
rect 137786 103018 138022 103254
rect 137786 102698 138022 102934
rect 137786 67018 138022 67254
rect 137786 66698 138022 66934
rect 137786 31018 138022 31254
rect 137786 30698 138022 30934
rect 119786 -6222 120022 -5986
rect 119786 -6542 120022 -6306
rect 144986 290218 145222 290454
rect 144986 289898 145222 290134
rect 144986 254218 145222 254454
rect 144986 253898 145222 254134
rect 144986 218218 145222 218454
rect 144986 217898 145222 218134
rect 144986 182218 145222 182454
rect 144986 181898 145222 182134
rect 144986 146218 145222 146454
rect 144986 145898 145222 146134
rect 144986 110218 145222 110454
rect 144986 109898 145222 110134
rect 144986 74218 145222 74454
rect 144986 73898 145222 74134
rect 144986 38218 145222 38454
rect 144986 37898 145222 38134
rect 144986 2218 145222 2454
rect 144986 1898 145222 2134
rect 144986 -582 145222 -346
rect 144986 -902 145222 -666
rect 148586 293818 148822 294054
rect 148586 293498 148822 293734
rect 148586 257818 148822 258054
rect 148586 257498 148822 257734
rect 148586 221818 148822 222054
rect 148586 221498 148822 221734
rect 148586 185818 148822 186054
rect 148586 185498 148822 185734
rect 148586 149818 148822 150054
rect 148586 149498 148822 149734
rect 148586 113818 148822 114054
rect 148586 113498 148822 113734
rect 148586 77818 148822 78054
rect 148586 77498 148822 77734
rect 148586 41818 148822 42054
rect 148586 41498 148822 41734
rect 148586 5818 148822 6054
rect 148586 5498 148822 5734
rect 148586 -2462 148822 -2226
rect 148586 -2782 148822 -2546
rect 152186 297418 152422 297654
rect 152186 297098 152422 297334
rect 152186 261418 152422 261654
rect 152186 261098 152422 261334
rect 152186 225418 152422 225654
rect 152186 225098 152422 225334
rect 152186 189418 152422 189654
rect 152186 189098 152422 189334
rect 152186 153418 152422 153654
rect 152186 153098 152422 153334
rect 152186 117418 152422 117654
rect 152186 117098 152422 117334
rect 152186 81418 152422 81654
rect 152186 81098 152422 81334
rect 152186 45418 152422 45654
rect 152186 45098 152422 45334
rect 152186 9418 152422 9654
rect 152186 9098 152422 9334
rect 152186 -4342 152422 -4106
rect 152186 -4662 152422 -4426
rect 155786 301018 156022 301254
rect 155786 300698 156022 300934
rect 155786 265018 156022 265254
rect 155786 264698 156022 264934
rect 155786 229018 156022 229254
rect 155786 228698 156022 228934
rect 155786 193018 156022 193254
rect 155786 192698 156022 192934
rect 155786 157018 156022 157254
rect 155786 156698 156022 156934
rect 155786 121018 156022 121254
rect 155786 120698 156022 120934
rect 155786 85018 156022 85254
rect 155786 84698 156022 84934
rect 155786 49018 156022 49254
rect 155786 48698 156022 48934
rect 155786 13018 156022 13254
rect 155786 12698 156022 12934
rect 137786 -7162 138022 -6926
rect 137786 -7482 138022 -7246
rect 162986 308218 163222 308454
rect 162986 307898 163222 308134
rect 162986 272218 163222 272454
rect 162986 271898 163222 272134
rect 162986 236218 163222 236454
rect 162986 235898 163222 236134
rect 162986 200218 163222 200454
rect 162986 199898 163222 200134
rect 162986 164218 163222 164454
rect 162986 163898 163222 164134
rect 162986 128218 163222 128454
rect 162986 127898 163222 128134
rect 162986 92218 163222 92454
rect 162986 91898 163222 92134
rect 162986 56218 163222 56454
rect 162986 55898 163222 56134
rect 162986 20218 163222 20454
rect 162986 19898 163222 20134
rect 162986 -1522 163222 -1286
rect 162986 -1842 163222 -1606
rect 166586 311818 166822 312054
rect 166586 311498 166822 311734
rect 166586 275818 166822 276054
rect 166586 275498 166822 275734
rect 166586 239818 166822 240054
rect 166586 239498 166822 239734
rect 166586 203818 166822 204054
rect 166586 203498 166822 203734
rect 166586 167818 166822 168054
rect 166586 167498 166822 167734
rect 166586 131818 166822 132054
rect 166586 131498 166822 131734
rect 166586 95818 166822 96054
rect 166586 95498 166822 95734
rect 166586 59818 166822 60054
rect 166586 59498 166822 59734
rect 166586 23818 166822 24054
rect 166586 23498 166822 23734
rect 166586 -3402 166822 -3166
rect 166586 -3722 166822 -3486
rect 170186 315418 170422 315654
rect 170186 315098 170422 315334
rect 170186 279418 170422 279654
rect 170186 279098 170422 279334
rect 170186 243418 170422 243654
rect 170186 243098 170422 243334
rect 170186 207418 170422 207654
rect 170186 207098 170422 207334
rect 170186 171418 170422 171654
rect 170186 171098 170422 171334
rect 170186 135418 170422 135654
rect 170186 135098 170422 135334
rect 170186 99418 170422 99654
rect 170186 99098 170422 99334
rect 170186 63418 170422 63654
rect 170186 63098 170422 63334
rect 170186 27418 170422 27654
rect 170186 27098 170422 27334
rect 170186 -5282 170422 -5046
rect 170186 -5602 170422 -5366
rect 173786 283018 174022 283254
rect 173786 282698 174022 282934
rect 173786 247018 174022 247254
rect 173786 246698 174022 246934
rect 173786 211018 174022 211254
rect 173786 210698 174022 210934
rect 173786 175018 174022 175254
rect 173786 174698 174022 174934
rect 173786 139018 174022 139254
rect 173786 138698 174022 138934
rect 173786 103018 174022 103254
rect 173786 102698 174022 102934
rect 173786 67018 174022 67254
rect 173786 66698 174022 66934
rect 173786 31018 174022 31254
rect 173786 30698 174022 30934
rect 155786 -6222 156022 -5986
rect 155786 -6542 156022 -6306
rect 180986 290218 181222 290454
rect 180986 289898 181222 290134
rect 180986 254218 181222 254454
rect 180986 253898 181222 254134
rect 180986 218218 181222 218454
rect 180986 217898 181222 218134
rect 180986 182218 181222 182454
rect 180986 181898 181222 182134
rect 180986 146218 181222 146454
rect 180986 145898 181222 146134
rect 180986 110218 181222 110454
rect 180986 109898 181222 110134
rect 180986 74218 181222 74454
rect 180986 73898 181222 74134
rect 180986 38218 181222 38454
rect 180986 37898 181222 38134
rect 180986 2218 181222 2454
rect 180986 1898 181222 2134
rect 180986 -582 181222 -346
rect 180986 -902 181222 -666
rect 184586 293818 184822 294054
rect 184586 293498 184822 293734
rect 184586 257818 184822 258054
rect 184586 257498 184822 257734
rect 184586 221818 184822 222054
rect 184586 221498 184822 221734
rect 184586 185818 184822 186054
rect 184586 185498 184822 185734
rect 184586 149818 184822 150054
rect 184586 149498 184822 149734
rect 184586 113818 184822 114054
rect 184586 113498 184822 113734
rect 184586 77818 184822 78054
rect 184586 77498 184822 77734
rect 184586 41818 184822 42054
rect 184586 41498 184822 41734
rect 184586 5818 184822 6054
rect 184586 5498 184822 5734
rect 184586 -2462 184822 -2226
rect 184586 -2782 184822 -2546
rect 188186 297418 188422 297654
rect 188186 297098 188422 297334
rect 188186 261418 188422 261654
rect 188186 261098 188422 261334
rect 188186 225418 188422 225654
rect 188186 225098 188422 225334
rect 188186 189418 188422 189654
rect 188186 189098 188422 189334
rect 188186 153418 188422 153654
rect 188186 153098 188422 153334
rect 188186 117418 188422 117654
rect 188186 117098 188422 117334
rect 188186 81418 188422 81654
rect 188186 81098 188422 81334
rect 188186 45418 188422 45654
rect 188186 45098 188422 45334
rect 188186 9418 188422 9654
rect 188186 9098 188422 9334
rect 188186 -4342 188422 -4106
rect 188186 -4662 188422 -4426
rect 191786 301018 192022 301254
rect 191786 300698 192022 300934
rect 191786 265018 192022 265254
rect 191786 264698 192022 264934
rect 191786 229018 192022 229254
rect 191786 228698 192022 228934
rect 191786 193018 192022 193254
rect 191786 192698 192022 192934
rect 191786 157018 192022 157254
rect 191786 156698 192022 156934
rect 191786 121018 192022 121254
rect 191786 120698 192022 120934
rect 191786 85018 192022 85254
rect 191786 84698 192022 84934
rect 191786 49018 192022 49254
rect 191786 48698 192022 48934
rect 191786 13018 192022 13254
rect 191786 12698 192022 12934
rect 173786 -7162 174022 -6926
rect 173786 -7482 174022 -7246
rect 198986 308218 199222 308454
rect 198986 307898 199222 308134
rect 198986 272218 199222 272454
rect 198986 271898 199222 272134
rect 198986 236218 199222 236454
rect 198986 235898 199222 236134
rect 198986 200218 199222 200454
rect 198986 199898 199222 200134
rect 198986 164218 199222 164454
rect 198986 163898 199222 164134
rect 198986 128218 199222 128454
rect 198986 127898 199222 128134
rect 198986 92218 199222 92454
rect 198986 91898 199222 92134
rect 198986 56218 199222 56454
rect 198986 55898 199222 56134
rect 198986 20218 199222 20454
rect 198986 19898 199222 20134
rect 198986 -1522 199222 -1286
rect 198986 -1842 199222 -1606
rect 202586 311818 202822 312054
rect 202586 311498 202822 311734
rect 202586 275818 202822 276054
rect 202586 275498 202822 275734
rect 202586 239818 202822 240054
rect 202586 239498 202822 239734
rect 202586 203818 202822 204054
rect 202586 203498 202822 203734
rect 202586 167818 202822 168054
rect 202586 167498 202822 167734
rect 202586 131818 202822 132054
rect 202586 131498 202822 131734
rect 202586 95818 202822 96054
rect 202586 95498 202822 95734
rect 202586 59818 202822 60054
rect 202586 59498 202822 59734
rect 202586 23818 202822 24054
rect 202586 23498 202822 23734
rect 202586 -3402 202822 -3166
rect 202586 -3722 202822 -3486
rect 206186 315418 206422 315654
rect 206186 315098 206422 315334
rect 206186 279418 206422 279654
rect 206186 279098 206422 279334
rect 206186 243418 206422 243654
rect 206186 243098 206422 243334
rect 206186 207418 206422 207654
rect 206186 207098 206422 207334
rect 206186 171418 206422 171654
rect 206186 171098 206422 171334
rect 206186 135418 206422 135654
rect 206186 135098 206422 135334
rect 206186 99418 206422 99654
rect 206186 99098 206422 99334
rect 206186 63418 206422 63654
rect 206186 63098 206422 63334
rect 206186 27418 206422 27654
rect 206186 27098 206422 27334
rect 206186 -5282 206422 -5046
rect 206186 -5602 206422 -5366
rect 209786 283018 210022 283254
rect 209786 282698 210022 282934
rect 209786 247018 210022 247254
rect 209786 246698 210022 246934
rect 209786 211018 210022 211254
rect 209786 210698 210022 210934
rect 209786 175018 210022 175254
rect 209786 174698 210022 174934
rect 209786 139018 210022 139254
rect 209786 138698 210022 138934
rect 209786 103018 210022 103254
rect 209786 102698 210022 102934
rect 209786 67018 210022 67254
rect 209786 66698 210022 66934
rect 209786 31018 210022 31254
rect 209786 30698 210022 30934
rect 191786 -6222 192022 -5986
rect 191786 -6542 192022 -6306
rect 216986 290218 217222 290454
rect 216986 289898 217222 290134
rect 216986 254218 217222 254454
rect 216986 253898 217222 254134
rect 216986 218218 217222 218454
rect 216986 217898 217222 218134
rect 216986 182218 217222 182454
rect 216986 181898 217222 182134
rect 216986 146218 217222 146454
rect 216986 145898 217222 146134
rect 216986 110218 217222 110454
rect 216986 109898 217222 110134
rect 216986 74218 217222 74454
rect 216986 73898 217222 74134
rect 216986 38218 217222 38454
rect 216986 37898 217222 38134
rect 216986 2218 217222 2454
rect 216986 1898 217222 2134
rect 216986 -582 217222 -346
rect 216986 -902 217222 -666
rect 220586 293818 220822 294054
rect 220586 293498 220822 293734
rect 220586 257818 220822 258054
rect 220586 257498 220822 257734
rect 220586 221818 220822 222054
rect 220586 221498 220822 221734
rect 220586 185818 220822 186054
rect 220586 185498 220822 185734
rect 220586 149818 220822 150054
rect 220586 149498 220822 149734
rect 220586 113818 220822 114054
rect 220586 113498 220822 113734
rect 220586 77818 220822 78054
rect 220586 77498 220822 77734
rect 220586 41818 220822 42054
rect 220586 41498 220822 41734
rect 220586 5818 220822 6054
rect 220586 5498 220822 5734
rect 220586 -2462 220822 -2226
rect 220586 -2782 220822 -2546
rect 224186 297418 224422 297654
rect 224186 297098 224422 297334
rect 224186 261418 224422 261654
rect 224186 261098 224422 261334
rect 224186 225418 224422 225654
rect 224186 225098 224422 225334
rect 224186 189418 224422 189654
rect 224186 189098 224422 189334
rect 224186 153418 224422 153654
rect 224186 153098 224422 153334
rect 224186 117418 224422 117654
rect 224186 117098 224422 117334
rect 224186 81418 224422 81654
rect 224186 81098 224422 81334
rect 224186 45418 224422 45654
rect 224186 45098 224422 45334
rect 224186 9418 224422 9654
rect 224186 9098 224422 9334
rect 224186 -4342 224422 -4106
rect 224186 -4662 224422 -4426
rect 227786 301018 228022 301254
rect 227786 300698 228022 300934
rect 227786 265018 228022 265254
rect 227786 264698 228022 264934
rect 227786 229018 228022 229254
rect 227786 228698 228022 228934
rect 227786 193018 228022 193254
rect 227786 192698 228022 192934
rect 227786 157018 228022 157254
rect 227786 156698 228022 156934
rect 227786 121018 228022 121254
rect 227786 120698 228022 120934
rect 227786 85018 228022 85254
rect 227786 84698 228022 84934
rect 227786 49018 228022 49254
rect 227786 48698 228022 48934
rect 227786 13018 228022 13254
rect 227786 12698 228022 12934
rect 209786 -7162 210022 -6926
rect 209786 -7482 210022 -7246
rect 234986 308218 235222 308454
rect 234986 307898 235222 308134
rect 234986 272218 235222 272454
rect 234986 271898 235222 272134
rect 234986 236218 235222 236454
rect 234986 235898 235222 236134
rect 234986 200218 235222 200454
rect 234986 199898 235222 200134
rect 234986 164218 235222 164454
rect 234986 163898 235222 164134
rect 234986 128218 235222 128454
rect 234986 127898 235222 128134
rect 234986 92218 235222 92454
rect 234986 91898 235222 92134
rect 234986 56218 235222 56454
rect 234986 55898 235222 56134
rect 234986 20218 235222 20454
rect 234986 19898 235222 20134
rect 234986 -1522 235222 -1286
rect 234986 -1842 235222 -1606
rect 238586 311818 238822 312054
rect 238586 311498 238822 311734
rect 238586 275818 238822 276054
rect 238586 275498 238822 275734
rect 238586 239818 238822 240054
rect 238586 239498 238822 239734
rect 238586 203818 238822 204054
rect 238586 203498 238822 203734
rect 238586 167818 238822 168054
rect 238586 167498 238822 167734
rect 238586 131818 238822 132054
rect 238586 131498 238822 131734
rect 238586 95818 238822 96054
rect 238586 95498 238822 95734
rect 238586 59818 238822 60054
rect 238586 59498 238822 59734
rect 238586 23818 238822 24054
rect 238586 23498 238822 23734
rect 238586 -3402 238822 -3166
rect 238586 -3722 238822 -3486
rect 242186 315418 242422 315654
rect 242186 315098 242422 315334
rect 242186 279418 242422 279654
rect 242186 279098 242422 279334
rect 242186 243418 242422 243654
rect 242186 243098 242422 243334
rect 242186 207418 242422 207654
rect 242186 207098 242422 207334
rect 242186 171418 242422 171654
rect 242186 171098 242422 171334
rect 242186 135418 242422 135654
rect 242186 135098 242422 135334
rect 242186 99418 242422 99654
rect 242186 99098 242422 99334
rect 242186 63418 242422 63654
rect 242186 63098 242422 63334
rect 242186 27418 242422 27654
rect 242186 27098 242422 27334
rect 242186 -5282 242422 -5046
rect 242186 -5602 242422 -5366
rect 245786 283018 246022 283254
rect 245786 282698 246022 282934
rect 245786 247018 246022 247254
rect 245786 246698 246022 246934
rect 245786 211018 246022 211254
rect 245786 210698 246022 210934
rect 245786 175018 246022 175254
rect 245786 174698 246022 174934
rect 245786 139018 246022 139254
rect 245786 138698 246022 138934
rect 245786 103018 246022 103254
rect 245786 102698 246022 102934
rect 245786 67018 246022 67254
rect 245786 66698 246022 66934
rect 245786 31018 246022 31254
rect 245786 30698 246022 30934
rect 227786 -6222 228022 -5986
rect 227786 -6542 228022 -6306
rect 252986 290218 253222 290454
rect 252986 289898 253222 290134
rect 252986 254218 253222 254454
rect 252986 253898 253222 254134
rect 252986 218218 253222 218454
rect 252986 217898 253222 218134
rect 252986 182218 253222 182454
rect 252986 181898 253222 182134
rect 252986 146218 253222 146454
rect 252986 145898 253222 146134
rect 252986 110218 253222 110454
rect 252986 109898 253222 110134
rect 252986 74218 253222 74454
rect 252986 73898 253222 74134
rect 252986 38218 253222 38454
rect 252986 37898 253222 38134
rect 252986 2218 253222 2454
rect 252986 1898 253222 2134
rect 252986 -582 253222 -346
rect 252986 -902 253222 -666
rect 256586 293818 256822 294054
rect 256586 293498 256822 293734
rect 256586 257818 256822 258054
rect 256586 257498 256822 257734
rect 256586 221818 256822 222054
rect 256586 221498 256822 221734
rect 256586 185818 256822 186054
rect 256586 185498 256822 185734
rect 256586 149818 256822 150054
rect 256586 149498 256822 149734
rect 256586 113818 256822 114054
rect 256586 113498 256822 113734
rect 256586 77818 256822 78054
rect 256586 77498 256822 77734
rect 256586 41818 256822 42054
rect 256586 41498 256822 41734
rect 256586 5818 256822 6054
rect 256586 5498 256822 5734
rect 256586 -2462 256822 -2226
rect 256586 -2782 256822 -2546
rect 260186 297418 260422 297654
rect 260186 297098 260422 297334
rect 260186 261418 260422 261654
rect 260186 261098 260422 261334
rect 260186 225418 260422 225654
rect 260186 225098 260422 225334
rect 260186 189418 260422 189654
rect 260186 189098 260422 189334
rect 260186 153418 260422 153654
rect 260186 153098 260422 153334
rect 260186 117418 260422 117654
rect 260186 117098 260422 117334
rect 260186 81418 260422 81654
rect 260186 81098 260422 81334
rect 260186 45418 260422 45654
rect 260186 45098 260422 45334
rect 260186 9418 260422 9654
rect 260186 9098 260422 9334
rect 260186 -4342 260422 -4106
rect 260186 -4662 260422 -4426
rect 263786 301018 264022 301254
rect 263786 300698 264022 300934
rect 263786 265018 264022 265254
rect 263786 264698 264022 264934
rect 263786 229018 264022 229254
rect 263786 228698 264022 228934
rect 263786 193018 264022 193254
rect 263786 192698 264022 192934
rect 263786 157018 264022 157254
rect 263786 156698 264022 156934
rect 263786 121018 264022 121254
rect 263786 120698 264022 120934
rect 263786 85018 264022 85254
rect 263786 84698 264022 84934
rect 263786 49018 264022 49254
rect 263786 48698 264022 48934
rect 263786 13018 264022 13254
rect 263786 12698 264022 12934
rect 245786 -7162 246022 -6926
rect 245786 -7482 246022 -7246
rect 270986 308218 271222 308454
rect 270986 307898 271222 308134
rect 270986 272218 271222 272454
rect 270986 271898 271222 272134
rect 270986 236218 271222 236454
rect 270986 235898 271222 236134
rect 270986 200218 271222 200454
rect 270986 199898 271222 200134
rect 270986 164218 271222 164454
rect 270986 163898 271222 164134
rect 270986 128218 271222 128454
rect 270986 127898 271222 128134
rect 270986 92218 271222 92454
rect 270986 91898 271222 92134
rect 270986 56218 271222 56454
rect 270986 55898 271222 56134
rect 270986 20218 271222 20454
rect 270986 19898 271222 20134
rect 270986 -1522 271222 -1286
rect 270986 -1842 271222 -1606
rect 274586 311818 274822 312054
rect 274586 311498 274822 311734
rect 274586 275818 274822 276054
rect 274586 275498 274822 275734
rect 274586 239818 274822 240054
rect 274586 239498 274822 239734
rect 274586 203818 274822 204054
rect 274586 203498 274822 203734
rect 274586 167818 274822 168054
rect 274586 167498 274822 167734
rect 274586 131818 274822 132054
rect 274586 131498 274822 131734
rect 274586 95818 274822 96054
rect 274586 95498 274822 95734
rect 274586 59818 274822 60054
rect 274586 59498 274822 59734
rect 274586 23818 274822 24054
rect 274586 23498 274822 23734
rect 274586 -3402 274822 -3166
rect 274586 -3722 274822 -3486
rect 278186 315418 278422 315654
rect 278186 315098 278422 315334
rect 278186 279418 278422 279654
rect 278186 279098 278422 279334
rect 278186 243418 278422 243654
rect 278186 243098 278422 243334
rect 278186 207418 278422 207654
rect 278186 207098 278422 207334
rect 278186 171418 278422 171654
rect 278186 171098 278422 171334
rect 278186 135418 278422 135654
rect 278186 135098 278422 135334
rect 278186 99418 278422 99654
rect 278186 99098 278422 99334
rect 278186 63418 278422 63654
rect 278186 63098 278422 63334
rect 278186 27418 278422 27654
rect 278186 27098 278422 27334
rect 278186 -5282 278422 -5046
rect 278186 -5602 278422 -5366
rect 281786 283018 282022 283254
rect 281786 282698 282022 282934
rect 281786 247018 282022 247254
rect 281786 246698 282022 246934
rect 281786 211018 282022 211254
rect 281786 210698 282022 210934
rect 281786 175018 282022 175254
rect 281786 174698 282022 174934
rect 281786 139018 282022 139254
rect 281786 138698 282022 138934
rect 281786 103018 282022 103254
rect 281786 102698 282022 102934
rect 281786 67018 282022 67254
rect 281786 66698 282022 66934
rect 281786 31018 282022 31254
rect 281786 30698 282022 30934
rect 263786 -6222 264022 -5986
rect 263786 -6542 264022 -6306
rect 288986 290218 289222 290454
rect 288986 289898 289222 290134
rect 288986 254218 289222 254454
rect 288986 253898 289222 254134
rect 288986 218218 289222 218454
rect 288986 217898 289222 218134
rect 288986 182218 289222 182454
rect 288986 181898 289222 182134
rect 288986 146218 289222 146454
rect 288986 145898 289222 146134
rect 288986 110218 289222 110454
rect 288986 109898 289222 110134
rect 288986 74218 289222 74454
rect 288986 73898 289222 74134
rect 288986 38218 289222 38454
rect 288986 37898 289222 38134
rect 288986 2218 289222 2454
rect 288986 1898 289222 2134
rect 288986 -582 289222 -346
rect 288986 -902 289222 -666
rect 292586 689818 292822 690054
rect 292586 689498 292822 689734
rect 292586 653818 292822 654054
rect 292586 653498 292822 653734
rect 292586 617818 292822 618054
rect 292586 617498 292822 617734
rect 292586 581818 292822 582054
rect 292586 581498 292822 581734
rect 292586 545818 292822 546054
rect 292586 545498 292822 545734
rect 292586 509818 292822 510054
rect 292586 509498 292822 509734
rect 292586 473818 292822 474054
rect 292586 473498 292822 473734
rect 292586 437818 292822 438054
rect 292586 437498 292822 437734
rect 292586 401818 292822 402054
rect 292586 401498 292822 401734
rect 292586 365818 292822 366054
rect 292586 365498 292822 365734
rect 292586 329818 292822 330054
rect 292586 329498 292822 329734
rect 292586 293818 292822 294054
rect 292586 293498 292822 293734
rect 292586 257818 292822 258054
rect 292586 257498 292822 257734
rect 292586 221818 292822 222054
rect 292586 221498 292822 221734
rect 292586 185818 292822 186054
rect 292586 185498 292822 185734
rect 292586 149818 292822 150054
rect 292586 149498 292822 149734
rect 292586 113818 292822 114054
rect 292586 113498 292822 113734
rect 292586 77818 292822 78054
rect 292586 77498 292822 77734
rect 292586 41818 292822 42054
rect 292586 41498 292822 41734
rect 292586 5818 292822 6054
rect 292586 5498 292822 5734
rect 292586 -2462 292822 -2226
rect 292586 -2782 292822 -2546
rect 296186 693418 296422 693654
rect 296186 693098 296422 693334
rect 317786 711182 318022 711418
rect 317786 710862 318022 711098
rect 314186 709302 314422 709538
rect 314186 708982 314422 709218
rect 310586 707422 310822 707658
rect 310586 707102 310822 707338
rect 299786 697018 300022 697254
rect 299786 696698 300022 696934
rect 296186 657418 296422 657654
rect 296186 657098 296422 657334
rect 299786 661018 300022 661254
rect 299786 660698 300022 660934
rect 296186 621418 296422 621654
rect 296186 621098 296422 621334
rect 296186 585418 296422 585654
rect 296186 585098 296422 585334
rect 296186 549418 296422 549654
rect 296186 549098 296422 549334
rect 296186 513418 296422 513654
rect 296186 513098 296422 513334
rect 296186 477418 296422 477654
rect 296186 477098 296422 477334
rect 296186 441418 296422 441654
rect 296186 441098 296422 441334
rect 296186 405418 296422 405654
rect 296186 405098 296422 405334
rect 296186 369418 296422 369654
rect 296186 369098 296422 369334
rect 296186 333418 296422 333654
rect 296186 333098 296422 333334
rect 296186 297418 296422 297654
rect 296186 297098 296422 297334
rect 296186 261418 296422 261654
rect 296186 261098 296422 261334
rect 296186 225418 296422 225654
rect 296186 225098 296422 225334
rect 296186 189418 296422 189654
rect 296186 189098 296422 189334
rect 296186 153418 296422 153654
rect 296186 153098 296422 153334
rect 296186 117418 296422 117654
rect 296186 117098 296422 117334
rect 296186 81418 296422 81654
rect 296186 81098 296422 81334
rect 296186 45418 296422 45654
rect 296186 45098 296422 45334
rect 296186 9418 296422 9654
rect 296186 9098 296422 9334
rect 296186 -4342 296422 -4106
rect 296186 -4662 296422 -4426
rect 306986 705542 307222 705778
rect 306986 705222 307222 705458
rect 306986 668218 307222 668454
rect 306986 667898 307222 668134
rect 310586 671818 310822 672054
rect 310586 671498 310822 671734
rect 314186 675418 314422 675654
rect 314186 675098 314422 675334
rect 335786 710242 336022 710478
rect 335786 709922 336022 710158
rect 332186 708362 332422 708598
rect 332186 708042 332422 708278
rect 328586 706482 328822 706718
rect 328586 706162 328822 706398
rect 317786 679018 318022 679254
rect 317786 678698 318022 678934
rect 324986 704602 325222 704838
rect 324986 704282 325222 704518
rect 324986 686218 325222 686454
rect 324986 685898 325222 686134
rect 328586 689818 328822 690054
rect 328586 689498 328822 689734
rect 332186 693418 332422 693654
rect 332186 693098 332422 693334
rect 332186 657418 332422 657654
rect 332186 657098 332422 657334
rect 353786 711182 354022 711418
rect 353786 710862 354022 711098
rect 350186 709302 350422 709538
rect 350186 708982 350422 709218
rect 346586 707422 346822 707658
rect 346586 707102 346822 707338
rect 335786 697018 336022 697254
rect 335786 696698 336022 696934
rect 335786 661018 336022 661254
rect 335786 660698 336022 660934
rect 342986 705542 343222 705778
rect 342986 705222 343222 705458
rect 342986 668218 343222 668454
rect 342986 667898 343222 668134
rect 346586 671818 346822 672054
rect 346586 671498 346822 671734
rect 350186 675418 350422 675654
rect 350186 675098 350422 675334
rect 371786 710242 372022 710478
rect 371786 709922 372022 710158
rect 368186 708362 368422 708598
rect 368186 708042 368422 708278
rect 364586 706482 364822 706718
rect 364586 706162 364822 706398
rect 360986 704602 361222 704838
rect 360986 704282 361222 704518
rect 360986 686218 361222 686454
rect 360986 685898 361222 686134
rect 353786 679018 354022 679254
rect 353786 678698 354022 678934
rect 364586 689818 364822 690054
rect 364586 689498 364822 689734
rect 368186 693418 368422 693654
rect 368186 693098 368422 693334
rect 368186 657418 368422 657654
rect 368186 657098 368422 657334
rect 389786 711182 390022 711418
rect 389786 710862 390022 711098
rect 386186 709302 386422 709538
rect 386186 708982 386422 709218
rect 382586 707422 382822 707658
rect 382586 707102 382822 707338
rect 371786 697018 372022 697254
rect 371786 696698 372022 696934
rect 378986 705542 379222 705778
rect 378986 705222 379222 705458
rect 371786 661018 372022 661254
rect 371786 660698 372022 660934
rect 378986 668218 379222 668454
rect 378986 667898 379222 668134
rect 382586 671818 382822 672054
rect 382586 671498 382822 671734
rect 386186 675418 386422 675654
rect 386186 675098 386422 675334
rect 407786 710242 408022 710478
rect 407786 709922 408022 710158
rect 404186 708362 404422 708598
rect 404186 708042 404422 708278
rect 400586 706482 400822 706718
rect 400586 706162 400822 706398
rect 389786 679018 390022 679254
rect 389786 678698 390022 678934
rect 396986 704602 397222 704838
rect 396986 704282 397222 704518
rect 396986 686218 397222 686454
rect 396986 685898 397222 686134
rect 396986 650218 397222 650454
rect 396986 649898 397222 650134
rect 386982 643018 387218 643254
rect 386982 642698 387218 642934
rect 386982 639418 387218 639654
rect 386982 639098 387218 639334
rect 386982 635818 387218 636054
rect 386982 635498 387218 635734
rect 386982 632218 387218 632454
rect 386982 631898 387218 632134
rect 299786 625018 300022 625254
rect 299786 624698 300022 624934
rect 386536 625018 386772 625254
rect 386536 624698 386772 624934
rect 386536 621418 386772 621654
rect 386536 621098 386772 621334
rect 386536 617818 386772 618054
rect 386536 617498 386772 617734
rect 386536 614218 386772 614454
rect 386536 613898 386772 614134
rect 396986 614218 397222 614454
rect 396986 613898 397222 614134
rect 386982 607018 387218 607254
rect 386982 606698 387218 606934
rect 386982 603418 387218 603654
rect 386982 603098 387218 603334
rect 386982 599818 387218 600054
rect 386982 599498 387218 599734
rect 386982 596218 387218 596454
rect 386982 595898 387218 596134
rect 299786 589018 300022 589254
rect 299786 588698 300022 588934
rect 386536 589018 386772 589254
rect 386536 588698 386772 588934
rect 386536 585418 386772 585654
rect 386536 585098 386772 585334
rect 386536 581818 386772 582054
rect 386536 581498 386772 581734
rect 386536 578218 386772 578454
rect 386536 577898 386772 578134
rect 396986 578218 397222 578454
rect 396986 577898 397222 578134
rect 386982 571018 387218 571254
rect 386982 570698 387218 570934
rect 386982 567418 387218 567654
rect 386982 567098 387218 567334
rect 386982 563818 387218 564054
rect 386982 563498 387218 563734
rect 299786 553018 300022 553254
rect 299786 552698 300022 552934
rect 299786 517018 300022 517254
rect 299786 516698 300022 516934
rect 299786 481018 300022 481254
rect 299786 480698 300022 480934
rect 299786 445018 300022 445254
rect 299786 444698 300022 444934
rect 299786 409018 300022 409254
rect 299786 408698 300022 408934
rect 299786 373018 300022 373254
rect 299786 372698 300022 372934
rect 299786 337018 300022 337254
rect 299786 336698 300022 336934
rect 299786 301018 300022 301254
rect 299786 300698 300022 300934
rect 299786 265018 300022 265254
rect 299786 264698 300022 264934
rect 299786 229018 300022 229254
rect 299786 228698 300022 228934
rect 299786 193018 300022 193254
rect 299786 192698 300022 192934
rect 299786 157018 300022 157254
rect 299786 156698 300022 156934
rect 299786 121018 300022 121254
rect 299786 120698 300022 120934
rect 299786 85018 300022 85254
rect 299786 84698 300022 84934
rect 299786 49018 300022 49254
rect 299786 48698 300022 48934
rect 299786 13018 300022 13254
rect 299786 12698 300022 12934
rect 281786 -7162 282022 -6926
rect 281786 -7482 282022 -7246
rect 306986 524218 307222 524454
rect 306986 523898 307222 524134
rect 306986 488218 307222 488454
rect 306986 487898 307222 488134
rect 306986 452218 307222 452454
rect 306986 451898 307222 452134
rect 306986 416218 307222 416454
rect 306986 415898 307222 416134
rect 306986 380218 307222 380454
rect 306986 379898 307222 380134
rect 306986 344218 307222 344454
rect 306986 343898 307222 344134
rect 306986 308218 307222 308454
rect 306986 307898 307222 308134
rect 306986 272218 307222 272454
rect 306986 271898 307222 272134
rect 306986 236218 307222 236454
rect 306986 235898 307222 236134
rect 306986 200218 307222 200454
rect 306986 199898 307222 200134
rect 306986 164218 307222 164454
rect 306986 163898 307222 164134
rect 306986 128218 307222 128454
rect 306986 127898 307222 128134
rect 306986 92218 307222 92454
rect 306986 91898 307222 92134
rect 306986 56218 307222 56454
rect 306986 55898 307222 56134
rect 306986 20218 307222 20454
rect 306986 19898 307222 20134
rect 306986 -1522 307222 -1286
rect 306986 -1842 307222 -1606
rect 310586 527818 310822 528054
rect 310586 527498 310822 527734
rect 310586 491818 310822 492054
rect 310586 491498 310822 491734
rect 310586 455818 310822 456054
rect 310586 455498 310822 455734
rect 310586 419818 310822 420054
rect 310586 419498 310822 419734
rect 310586 383818 310822 384054
rect 310586 383498 310822 383734
rect 310586 347818 310822 348054
rect 310586 347498 310822 347734
rect 310586 311818 310822 312054
rect 310586 311498 310822 311734
rect 310586 275818 310822 276054
rect 310586 275498 310822 275734
rect 310586 239818 310822 240054
rect 310586 239498 310822 239734
rect 310586 203818 310822 204054
rect 310586 203498 310822 203734
rect 310586 167818 310822 168054
rect 310586 167498 310822 167734
rect 310586 131818 310822 132054
rect 310586 131498 310822 131734
rect 310586 95818 310822 96054
rect 310586 95498 310822 95734
rect 310586 59818 310822 60054
rect 310586 59498 310822 59734
rect 310586 23818 310822 24054
rect 310586 23498 310822 23734
rect 310586 -3402 310822 -3166
rect 310586 -3722 310822 -3486
rect 314186 531418 314422 531654
rect 314186 531098 314422 531334
rect 314186 495418 314422 495654
rect 314186 495098 314422 495334
rect 314186 459418 314422 459654
rect 314186 459098 314422 459334
rect 314186 423418 314422 423654
rect 314186 423098 314422 423334
rect 314186 387418 314422 387654
rect 314186 387098 314422 387334
rect 314186 351418 314422 351654
rect 314186 351098 314422 351334
rect 314186 315418 314422 315654
rect 314186 315098 314422 315334
rect 314186 279418 314422 279654
rect 314186 279098 314422 279334
rect 314186 243418 314422 243654
rect 314186 243098 314422 243334
rect 314186 207418 314422 207654
rect 314186 207098 314422 207334
rect 314186 171418 314422 171654
rect 314186 171098 314422 171334
rect 314186 135418 314422 135654
rect 314186 135098 314422 135334
rect 314186 99418 314422 99654
rect 314186 99098 314422 99334
rect 314186 63418 314422 63654
rect 314186 63098 314422 63334
rect 314186 27418 314422 27654
rect 314186 27098 314422 27334
rect 314186 -5282 314422 -5046
rect 314186 -5602 314422 -5366
rect 317786 535018 318022 535254
rect 317786 534698 318022 534934
rect 317786 499018 318022 499254
rect 317786 498698 318022 498934
rect 317786 463018 318022 463254
rect 317786 462698 318022 462934
rect 317786 427018 318022 427254
rect 317786 426698 318022 426934
rect 317786 391018 318022 391254
rect 317786 390698 318022 390934
rect 317786 355018 318022 355254
rect 317786 354698 318022 354934
rect 317786 319018 318022 319254
rect 317786 318698 318022 318934
rect 317786 283018 318022 283254
rect 317786 282698 318022 282934
rect 317786 247018 318022 247254
rect 317786 246698 318022 246934
rect 317786 211018 318022 211254
rect 317786 210698 318022 210934
rect 317786 175018 318022 175254
rect 317786 174698 318022 174934
rect 317786 139018 318022 139254
rect 317786 138698 318022 138934
rect 317786 103018 318022 103254
rect 317786 102698 318022 102934
rect 317786 67018 318022 67254
rect 317786 66698 318022 66934
rect 317786 31018 318022 31254
rect 317786 30698 318022 30934
rect 299786 -6222 300022 -5986
rect 299786 -6542 300022 -6306
rect 324986 542218 325222 542454
rect 324986 541898 325222 542134
rect 324986 506218 325222 506454
rect 324986 505898 325222 506134
rect 324986 470218 325222 470454
rect 324986 469898 325222 470134
rect 324986 434218 325222 434454
rect 324986 433898 325222 434134
rect 324986 398218 325222 398454
rect 324986 397898 325222 398134
rect 324986 362218 325222 362454
rect 324986 361898 325222 362134
rect 324986 326218 325222 326454
rect 324986 325898 325222 326134
rect 324986 290218 325222 290454
rect 324986 289898 325222 290134
rect 324986 254218 325222 254454
rect 324986 253898 325222 254134
rect 324986 218218 325222 218454
rect 324986 217898 325222 218134
rect 324986 182218 325222 182454
rect 324986 181898 325222 182134
rect 324986 146218 325222 146454
rect 324986 145898 325222 146134
rect 324986 110218 325222 110454
rect 324986 109898 325222 110134
rect 324986 74218 325222 74454
rect 324986 73898 325222 74134
rect 324986 38218 325222 38454
rect 324986 37898 325222 38134
rect 324986 2218 325222 2454
rect 324986 1898 325222 2134
rect 324986 -582 325222 -346
rect 324986 -902 325222 -666
rect 328586 545818 328822 546054
rect 328586 545498 328822 545734
rect 328586 509818 328822 510054
rect 328586 509498 328822 509734
rect 328586 473818 328822 474054
rect 328586 473498 328822 473734
rect 328586 437818 328822 438054
rect 328586 437498 328822 437734
rect 328586 401818 328822 402054
rect 328586 401498 328822 401734
rect 328586 365818 328822 366054
rect 328586 365498 328822 365734
rect 328586 329818 328822 330054
rect 328586 329498 328822 329734
rect 328586 293818 328822 294054
rect 328586 293498 328822 293734
rect 328586 257818 328822 258054
rect 328586 257498 328822 257734
rect 328586 221818 328822 222054
rect 328586 221498 328822 221734
rect 328586 185818 328822 186054
rect 328586 185498 328822 185734
rect 328586 149818 328822 150054
rect 328586 149498 328822 149734
rect 328586 113818 328822 114054
rect 328586 113498 328822 113734
rect 328586 77818 328822 78054
rect 328586 77498 328822 77734
rect 328586 41818 328822 42054
rect 328586 41498 328822 41734
rect 328586 5818 328822 6054
rect 328586 5498 328822 5734
rect 328586 -2462 328822 -2226
rect 328586 -2782 328822 -2546
rect 332186 549418 332422 549654
rect 332186 549098 332422 549334
rect 332186 513418 332422 513654
rect 332186 513098 332422 513334
rect 332186 477418 332422 477654
rect 332186 477098 332422 477334
rect 332186 441418 332422 441654
rect 332186 441098 332422 441334
rect 332186 405418 332422 405654
rect 332186 405098 332422 405334
rect 332186 369418 332422 369654
rect 332186 369098 332422 369334
rect 332186 333418 332422 333654
rect 332186 333098 332422 333334
rect 332186 297418 332422 297654
rect 332186 297098 332422 297334
rect 332186 261418 332422 261654
rect 332186 261098 332422 261334
rect 332186 225418 332422 225654
rect 332186 225098 332422 225334
rect 332186 189418 332422 189654
rect 332186 189098 332422 189334
rect 332186 153418 332422 153654
rect 332186 153098 332422 153334
rect 332186 117418 332422 117654
rect 332186 117098 332422 117334
rect 332186 81418 332422 81654
rect 332186 81098 332422 81334
rect 332186 45418 332422 45654
rect 332186 45098 332422 45334
rect 332186 9418 332422 9654
rect 332186 9098 332422 9334
rect 332186 -4342 332422 -4106
rect 332186 -4662 332422 -4426
rect 335786 553018 336022 553254
rect 335786 552698 336022 552934
rect 335786 517018 336022 517254
rect 335786 516698 336022 516934
rect 335786 481018 336022 481254
rect 335786 480698 336022 480934
rect 335786 445018 336022 445254
rect 335786 444698 336022 444934
rect 342986 524218 343222 524454
rect 342986 523898 343222 524134
rect 342986 488218 343222 488454
rect 342986 487898 343222 488134
rect 342986 452218 343222 452454
rect 342986 451898 343222 452134
rect 342986 416218 343222 416454
rect 342986 415898 343222 416134
rect 346586 527818 346822 528054
rect 346586 527498 346822 527734
rect 346586 491818 346822 492054
rect 346586 491498 346822 491734
rect 346586 455818 346822 456054
rect 346586 455498 346822 455734
rect 346586 419818 346822 420054
rect 346586 419498 346822 419734
rect 350186 531418 350422 531654
rect 350186 531098 350422 531334
rect 350186 495418 350422 495654
rect 350186 495098 350422 495334
rect 350186 459418 350422 459654
rect 350186 459098 350422 459334
rect 350186 423418 350422 423654
rect 350186 423098 350422 423334
rect 353786 535018 354022 535254
rect 353786 534698 354022 534934
rect 353786 499018 354022 499254
rect 353786 498698 354022 498934
rect 353786 463018 354022 463254
rect 353786 462698 354022 462934
rect 353786 427018 354022 427254
rect 353786 426698 354022 426934
rect 360986 542218 361222 542454
rect 360986 541898 361222 542134
rect 360986 506218 361222 506454
rect 360986 505898 361222 506134
rect 360986 470218 361222 470454
rect 360986 469898 361222 470134
rect 360986 434218 361222 434454
rect 360986 433898 361222 434134
rect 364586 545818 364822 546054
rect 364586 545498 364822 545734
rect 364586 509818 364822 510054
rect 364586 509498 364822 509734
rect 364586 473818 364822 474054
rect 364586 473498 364822 473734
rect 364586 437818 364822 438054
rect 364586 437498 364822 437734
rect 368186 549418 368422 549654
rect 368186 549098 368422 549334
rect 368186 513418 368422 513654
rect 368186 513098 368422 513334
rect 368186 477418 368422 477654
rect 368186 477098 368422 477334
rect 368186 441418 368422 441654
rect 368186 441098 368422 441334
rect 371786 553018 372022 553254
rect 371786 552698 372022 552934
rect 371786 517018 372022 517254
rect 371786 516698 372022 516934
rect 371786 481018 372022 481254
rect 371786 480698 372022 480934
rect 371786 445018 372022 445254
rect 371786 444698 372022 444934
rect 378986 524218 379222 524454
rect 378986 523898 379222 524134
rect 378986 488218 379222 488454
rect 378986 487898 379222 488134
rect 378986 452218 379222 452454
rect 378986 451898 379222 452134
rect 378986 416218 379222 416454
rect 378986 415898 379222 416134
rect 382586 527818 382822 528054
rect 382586 527498 382822 527734
rect 382586 491818 382822 492054
rect 382586 491498 382822 491734
rect 382586 455818 382822 456054
rect 382586 455498 382822 455734
rect 382586 419818 382822 420054
rect 382586 419498 382822 419734
rect 386186 531418 386422 531654
rect 386186 531098 386422 531334
rect 386186 495418 386422 495654
rect 386186 495098 386422 495334
rect 386186 459418 386422 459654
rect 386186 459098 386422 459334
rect 386186 423418 386422 423654
rect 386186 423098 386422 423334
rect 389786 535018 390022 535254
rect 389786 534698 390022 534934
rect 389786 499018 390022 499254
rect 389786 498698 390022 498934
rect 389786 463018 390022 463254
rect 389786 462698 390022 462934
rect 389786 427018 390022 427254
rect 389786 426698 390022 426934
rect 396986 542218 397222 542454
rect 396986 541898 397222 542134
rect 396986 506218 397222 506454
rect 396986 505898 397222 506134
rect 396986 470218 397222 470454
rect 396986 469898 397222 470134
rect 396986 434218 397222 434454
rect 396986 433898 397222 434134
rect 400586 689818 400822 690054
rect 400586 689498 400822 689734
rect 400586 653818 400822 654054
rect 400586 653498 400822 653734
rect 400586 617818 400822 618054
rect 400586 617498 400822 617734
rect 400586 581818 400822 582054
rect 400586 581498 400822 581734
rect 400586 545818 400822 546054
rect 400586 545498 400822 545734
rect 400586 509818 400822 510054
rect 400586 509498 400822 509734
rect 400586 473818 400822 474054
rect 400586 473498 400822 473734
rect 400586 437818 400822 438054
rect 400586 437498 400822 437734
rect 404186 693418 404422 693654
rect 404186 693098 404422 693334
rect 404186 657418 404422 657654
rect 404186 657098 404422 657334
rect 404186 621418 404422 621654
rect 404186 621098 404422 621334
rect 404186 585418 404422 585654
rect 404186 585098 404422 585334
rect 404186 549418 404422 549654
rect 404186 549098 404422 549334
rect 404186 513418 404422 513654
rect 404186 513098 404422 513334
rect 404186 477418 404422 477654
rect 404186 477098 404422 477334
rect 404186 441418 404422 441654
rect 404186 441098 404422 441334
rect 425786 711182 426022 711418
rect 425786 710862 426022 711098
rect 422186 709302 422422 709538
rect 422186 708982 422422 709218
rect 418586 707422 418822 707658
rect 418586 707102 418822 707338
rect 407786 697018 408022 697254
rect 407786 696698 408022 696934
rect 407786 661018 408022 661254
rect 407786 660698 408022 660934
rect 407786 625018 408022 625254
rect 407786 624698 408022 624934
rect 407786 589018 408022 589254
rect 407786 588698 408022 588934
rect 407786 553018 408022 553254
rect 407786 552698 408022 552934
rect 407786 517018 408022 517254
rect 407786 516698 408022 516934
rect 407786 481018 408022 481254
rect 407786 480698 408022 480934
rect 407786 445018 408022 445254
rect 407786 444698 408022 444934
rect 414986 705542 415222 705778
rect 414986 705222 415222 705458
rect 414986 668218 415222 668454
rect 414986 667898 415222 668134
rect 414986 632218 415222 632454
rect 414986 631898 415222 632134
rect 414986 596218 415222 596454
rect 414986 595898 415222 596134
rect 414986 560218 415222 560454
rect 414986 559898 415222 560134
rect 414986 524218 415222 524454
rect 414986 523898 415222 524134
rect 414986 488218 415222 488454
rect 414986 487898 415222 488134
rect 414986 452218 415222 452454
rect 414986 451898 415222 452134
rect 414986 416218 415222 416454
rect 414986 415898 415222 416134
rect 418586 671818 418822 672054
rect 418586 671498 418822 671734
rect 418586 635818 418822 636054
rect 418586 635498 418822 635734
rect 418586 599818 418822 600054
rect 418586 599498 418822 599734
rect 418586 563818 418822 564054
rect 418586 563498 418822 563734
rect 418586 527818 418822 528054
rect 418586 527498 418822 527734
rect 418586 491818 418822 492054
rect 418586 491498 418822 491734
rect 418586 455818 418822 456054
rect 418586 455498 418822 455734
rect 418586 419818 418822 420054
rect 418586 419498 418822 419734
rect 422186 675418 422422 675654
rect 422186 675098 422422 675334
rect 422186 639418 422422 639654
rect 422186 639098 422422 639334
rect 422186 603418 422422 603654
rect 422186 603098 422422 603334
rect 422186 567418 422422 567654
rect 422186 567098 422422 567334
rect 422186 531418 422422 531654
rect 422186 531098 422422 531334
rect 422186 495418 422422 495654
rect 422186 495098 422422 495334
rect 422186 459418 422422 459654
rect 422186 459098 422422 459334
rect 422186 423418 422422 423654
rect 422186 423098 422422 423334
rect 335786 409018 336022 409254
rect 335786 408698 336022 408934
rect 340524 409018 340760 409254
rect 340524 408698 340760 408934
rect 340524 405418 340760 405654
rect 340524 405098 340760 405334
rect 340524 401818 340760 402054
rect 340524 401498 340760 401734
rect 340524 398218 340760 398454
rect 340524 397898 340760 398134
rect 340078 391018 340314 391254
rect 340078 390698 340314 390934
rect 340078 387418 340314 387654
rect 340078 387098 340314 387334
rect 422186 387418 422422 387654
rect 422186 387098 422422 387334
rect 340078 383818 340314 384054
rect 340078 383498 340314 383734
rect 340078 380218 340314 380454
rect 340078 379898 340314 380134
rect 335786 373018 336022 373254
rect 335786 372698 336022 372934
rect 340524 373018 340760 373254
rect 340524 372698 340760 372934
rect 340524 369418 340760 369654
rect 340524 369098 340760 369334
rect 340524 365818 340760 366054
rect 340524 365498 340760 365734
rect 340524 362218 340760 362454
rect 340524 361898 340760 362134
rect 340078 355018 340314 355254
rect 340078 354698 340314 354934
rect 340078 351418 340314 351654
rect 340078 351098 340314 351334
rect 422186 351418 422422 351654
rect 422186 351098 422422 351334
rect 340078 347818 340314 348054
rect 340078 347498 340314 347734
rect 340078 344218 340314 344454
rect 340078 343898 340314 344134
rect 335786 337018 336022 337254
rect 335786 336698 336022 336934
rect 340524 337018 340760 337254
rect 340524 336698 340760 336934
rect 340524 333418 340760 333654
rect 340524 333098 340760 333334
rect 340524 329818 340760 330054
rect 340524 329498 340760 329734
rect 340524 326218 340760 326454
rect 340524 325898 340760 326134
rect 335786 301018 336022 301254
rect 335786 300698 336022 300934
rect 335786 265018 336022 265254
rect 335786 264698 336022 264934
rect 335786 229018 336022 229254
rect 335786 228698 336022 228934
rect 335786 193018 336022 193254
rect 335786 192698 336022 192934
rect 335786 157018 336022 157254
rect 335786 156698 336022 156934
rect 335786 121018 336022 121254
rect 335786 120698 336022 120934
rect 335786 85018 336022 85254
rect 335786 84698 336022 84934
rect 335786 49018 336022 49254
rect 335786 48698 336022 48934
rect 335786 13018 336022 13254
rect 335786 12698 336022 12934
rect 317786 -7162 318022 -6926
rect 317786 -7482 318022 -7246
rect 342986 308218 343222 308454
rect 342986 307898 343222 308134
rect 342986 272218 343222 272454
rect 342986 271898 343222 272134
rect 342986 236218 343222 236454
rect 342986 235898 343222 236134
rect 342986 200218 343222 200454
rect 342986 199898 343222 200134
rect 342986 164218 343222 164454
rect 342986 163898 343222 164134
rect 342986 128218 343222 128454
rect 342986 127898 343222 128134
rect 342986 92218 343222 92454
rect 342986 91898 343222 92134
rect 342986 56218 343222 56454
rect 342986 55898 343222 56134
rect 342986 20218 343222 20454
rect 342986 19898 343222 20134
rect 342986 -1522 343222 -1286
rect 342986 -1842 343222 -1606
rect 346586 311818 346822 312054
rect 346586 311498 346822 311734
rect 346586 275818 346822 276054
rect 346586 275498 346822 275734
rect 346586 239818 346822 240054
rect 346586 239498 346822 239734
rect 346586 203818 346822 204054
rect 346586 203498 346822 203734
rect 346586 167818 346822 168054
rect 346586 167498 346822 167734
rect 346586 131818 346822 132054
rect 346586 131498 346822 131734
rect 346586 95818 346822 96054
rect 346586 95498 346822 95734
rect 346586 59818 346822 60054
rect 346586 59498 346822 59734
rect 346586 23818 346822 24054
rect 346586 23498 346822 23734
rect 346586 -3402 346822 -3166
rect 346586 -3722 346822 -3486
rect 350186 315418 350422 315654
rect 350186 315098 350422 315334
rect 350186 279418 350422 279654
rect 350186 279098 350422 279334
rect 350186 243418 350422 243654
rect 350186 243098 350422 243334
rect 350186 207418 350422 207654
rect 350186 207098 350422 207334
rect 350186 171418 350422 171654
rect 350186 171098 350422 171334
rect 350186 135418 350422 135654
rect 350186 135098 350422 135334
rect 350186 99418 350422 99654
rect 350186 99098 350422 99334
rect 350186 63418 350422 63654
rect 350186 63098 350422 63334
rect 350186 27418 350422 27654
rect 350186 27098 350422 27334
rect 350186 -5282 350422 -5046
rect 350186 -5602 350422 -5366
rect 353786 283018 354022 283254
rect 353786 282698 354022 282934
rect 353786 247018 354022 247254
rect 353786 246698 354022 246934
rect 353786 211018 354022 211254
rect 353786 210698 354022 210934
rect 353786 175018 354022 175254
rect 353786 174698 354022 174934
rect 353786 139018 354022 139254
rect 353786 138698 354022 138934
rect 353786 103018 354022 103254
rect 353786 102698 354022 102934
rect 353786 67018 354022 67254
rect 353786 66698 354022 66934
rect 353786 31018 354022 31254
rect 353786 30698 354022 30934
rect 335786 -6222 336022 -5986
rect 335786 -6542 336022 -6306
rect 360986 290218 361222 290454
rect 360986 289898 361222 290134
rect 360986 254218 361222 254454
rect 360986 253898 361222 254134
rect 360986 218218 361222 218454
rect 360986 217898 361222 218134
rect 360986 182218 361222 182454
rect 360986 181898 361222 182134
rect 360986 146218 361222 146454
rect 360986 145898 361222 146134
rect 360986 110218 361222 110454
rect 360986 109898 361222 110134
rect 360986 74218 361222 74454
rect 360986 73898 361222 74134
rect 360986 38218 361222 38454
rect 360986 37898 361222 38134
rect 360986 2218 361222 2454
rect 360986 1898 361222 2134
rect 360986 -582 361222 -346
rect 360986 -902 361222 -666
rect 364586 293818 364822 294054
rect 364586 293498 364822 293734
rect 364586 257818 364822 258054
rect 364586 257498 364822 257734
rect 364586 221818 364822 222054
rect 364586 221498 364822 221734
rect 364586 185818 364822 186054
rect 364586 185498 364822 185734
rect 364586 149818 364822 150054
rect 364586 149498 364822 149734
rect 364586 113818 364822 114054
rect 364586 113498 364822 113734
rect 364586 77818 364822 78054
rect 364586 77498 364822 77734
rect 364586 41818 364822 42054
rect 364586 41498 364822 41734
rect 364586 5818 364822 6054
rect 364586 5498 364822 5734
rect 364586 -2462 364822 -2226
rect 364586 -2782 364822 -2546
rect 368186 297418 368422 297654
rect 368186 297098 368422 297334
rect 368186 261418 368422 261654
rect 368186 261098 368422 261334
rect 368186 225418 368422 225654
rect 368186 225098 368422 225334
rect 368186 189418 368422 189654
rect 368186 189098 368422 189334
rect 368186 153418 368422 153654
rect 368186 153098 368422 153334
rect 368186 117418 368422 117654
rect 368186 117098 368422 117334
rect 368186 81418 368422 81654
rect 368186 81098 368422 81334
rect 368186 45418 368422 45654
rect 368186 45098 368422 45334
rect 368186 9418 368422 9654
rect 368186 9098 368422 9334
rect 368186 -4342 368422 -4106
rect 368186 -4662 368422 -4426
rect 371786 301018 372022 301254
rect 371786 300698 372022 300934
rect 371786 265018 372022 265254
rect 371786 264698 372022 264934
rect 371786 229018 372022 229254
rect 371786 228698 372022 228934
rect 371786 193018 372022 193254
rect 371786 192698 372022 192934
rect 371786 157018 372022 157254
rect 371786 156698 372022 156934
rect 371786 121018 372022 121254
rect 371786 120698 372022 120934
rect 371786 85018 372022 85254
rect 371786 84698 372022 84934
rect 371786 49018 372022 49254
rect 371786 48698 372022 48934
rect 371786 13018 372022 13254
rect 371786 12698 372022 12934
rect 353786 -7162 354022 -6926
rect 353786 -7482 354022 -7246
rect 378986 308218 379222 308454
rect 378986 307898 379222 308134
rect 378986 272218 379222 272454
rect 378986 271898 379222 272134
rect 378986 236218 379222 236454
rect 378986 235898 379222 236134
rect 378986 200218 379222 200454
rect 378986 199898 379222 200134
rect 378986 164218 379222 164454
rect 378986 163898 379222 164134
rect 378986 128218 379222 128454
rect 378986 127898 379222 128134
rect 378986 92218 379222 92454
rect 378986 91898 379222 92134
rect 378986 56218 379222 56454
rect 378986 55898 379222 56134
rect 378986 20218 379222 20454
rect 378986 19898 379222 20134
rect 378986 -1522 379222 -1286
rect 378986 -1842 379222 -1606
rect 382586 311818 382822 312054
rect 382586 311498 382822 311734
rect 382586 275818 382822 276054
rect 382586 275498 382822 275734
rect 382586 239818 382822 240054
rect 382586 239498 382822 239734
rect 382586 203818 382822 204054
rect 382586 203498 382822 203734
rect 382586 167818 382822 168054
rect 382586 167498 382822 167734
rect 382586 131818 382822 132054
rect 382586 131498 382822 131734
rect 382586 95818 382822 96054
rect 382586 95498 382822 95734
rect 382586 59818 382822 60054
rect 382586 59498 382822 59734
rect 382586 23818 382822 24054
rect 382586 23498 382822 23734
rect 382586 -3402 382822 -3166
rect 382586 -3722 382822 -3486
rect 386186 315418 386422 315654
rect 386186 315098 386422 315334
rect 386186 279418 386422 279654
rect 386186 279098 386422 279334
rect 386186 243418 386422 243654
rect 386186 243098 386422 243334
rect 386186 207418 386422 207654
rect 386186 207098 386422 207334
rect 386186 171418 386422 171654
rect 386186 171098 386422 171334
rect 386186 135418 386422 135654
rect 386186 135098 386422 135334
rect 386186 99418 386422 99654
rect 386186 99098 386422 99334
rect 386186 63418 386422 63654
rect 386186 63098 386422 63334
rect 386186 27418 386422 27654
rect 386186 27098 386422 27334
rect 386186 -5282 386422 -5046
rect 386186 -5602 386422 -5366
rect 389786 283018 390022 283254
rect 389786 282698 390022 282934
rect 389786 247018 390022 247254
rect 389786 246698 390022 246934
rect 389786 211018 390022 211254
rect 389786 210698 390022 210934
rect 389786 175018 390022 175254
rect 389786 174698 390022 174934
rect 389786 139018 390022 139254
rect 389786 138698 390022 138934
rect 389786 103018 390022 103254
rect 389786 102698 390022 102934
rect 389786 67018 390022 67254
rect 389786 66698 390022 66934
rect 389786 31018 390022 31254
rect 389786 30698 390022 30934
rect 371786 -6222 372022 -5986
rect 371786 -6542 372022 -6306
rect 396986 290218 397222 290454
rect 396986 289898 397222 290134
rect 396986 254218 397222 254454
rect 396986 253898 397222 254134
rect 396986 218218 397222 218454
rect 396986 217898 397222 218134
rect 396986 182218 397222 182454
rect 396986 181898 397222 182134
rect 396986 146218 397222 146454
rect 396986 145898 397222 146134
rect 396986 110218 397222 110454
rect 396986 109898 397222 110134
rect 396986 74218 397222 74454
rect 396986 73898 397222 74134
rect 396986 38218 397222 38454
rect 396986 37898 397222 38134
rect 396986 2218 397222 2454
rect 396986 1898 397222 2134
rect 396986 -582 397222 -346
rect 396986 -902 397222 -666
rect 400586 293818 400822 294054
rect 400586 293498 400822 293734
rect 400586 257818 400822 258054
rect 400586 257498 400822 257734
rect 400586 221818 400822 222054
rect 400586 221498 400822 221734
rect 400586 185818 400822 186054
rect 400586 185498 400822 185734
rect 400586 149818 400822 150054
rect 400586 149498 400822 149734
rect 400586 113818 400822 114054
rect 400586 113498 400822 113734
rect 400586 77818 400822 78054
rect 400586 77498 400822 77734
rect 400586 41818 400822 42054
rect 400586 41498 400822 41734
rect 400586 5818 400822 6054
rect 400586 5498 400822 5734
rect 400586 -2462 400822 -2226
rect 400586 -2782 400822 -2546
rect 404186 297418 404422 297654
rect 404186 297098 404422 297334
rect 404186 261418 404422 261654
rect 404186 261098 404422 261334
rect 404186 225418 404422 225654
rect 404186 225098 404422 225334
rect 404186 189418 404422 189654
rect 404186 189098 404422 189334
rect 404186 153418 404422 153654
rect 404186 153098 404422 153334
rect 404186 117418 404422 117654
rect 404186 117098 404422 117334
rect 404186 81418 404422 81654
rect 404186 81098 404422 81334
rect 404186 45418 404422 45654
rect 404186 45098 404422 45334
rect 404186 9418 404422 9654
rect 404186 9098 404422 9334
rect 404186 -4342 404422 -4106
rect 404186 -4662 404422 -4426
rect 407786 301018 408022 301254
rect 407786 300698 408022 300934
rect 407786 265018 408022 265254
rect 407786 264698 408022 264934
rect 407786 229018 408022 229254
rect 407786 228698 408022 228934
rect 407786 193018 408022 193254
rect 407786 192698 408022 192934
rect 407786 157018 408022 157254
rect 407786 156698 408022 156934
rect 407786 121018 408022 121254
rect 407786 120698 408022 120934
rect 407786 85018 408022 85254
rect 407786 84698 408022 84934
rect 407786 49018 408022 49254
rect 407786 48698 408022 48934
rect 407786 13018 408022 13254
rect 407786 12698 408022 12934
rect 389786 -7162 390022 -6926
rect 389786 -7482 390022 -7246
rect 414986 308218 415222 308454
rect 414986 307898 415222 308134
rect 414986 272218 415222 272454
rect 414986 271898 415222 272134
rect 414986 236218 415222 236454
rect 414986 235898 415222 236134
rect 414986 200218 415222 200454
rect 414986 199898 415222 200134
rect 414986 164218 415222 164454
rect 414986 163898 415222 164134
rect 414986 128218 415222 128454
rect 414986 127898 415222 128134
rect 414986 92218 415222 92454
rect 414986 91898 415222 92134
rect 414986 56218 415222 56454
rect 414986 55898 415222 56134
rect 414986 20218 415222 20454
rect 414986 19898 415222 20134
rect 414986 -1522 415222 -1286
rect 414986 -1842 415222 -1606
rect 418586 311818 418822 312054
rect 418586 311498 418822 311734
rect 418586 275818 418822 276054
rect 418586 275498 418822 275734
rect 418586 239818 418822 240054
rect 418586 239498 418822 239734
rect 418586 203818 418822 204054
rect 418586 203498 418822 203734
rect 418586 167818 418822 168054
rect 418586 167498 418822 167734
rect 418586 131818 418822 132054
rect 418586 131498 418822 131734
rect 418586 95818 418822 96054
rect 418586 95498 418822 95734
rect 418586 59818 418822 60054
rect 418586 59498 418822 59734
rect 418586 23818 418822 24054
rect 418586 23498 418822 23734
rect 418586 -3402 418822 -3166
rect 418586 -3722 418822 -3486
rect 422186 315418 422422 315654
rect 422186 315098 422422 315334
rect 422186 279418 422422 279654
rect 422186 279098 422422 279334
rect 422186 243418 422422 243654
rect 422186 243098 422422 243334
rect 422186 207418 422422 207654
rect 422186 207098 422422 207334
rect 422186 171418 422422 171654
rect 422186 171098 422422 171334
rect 422186 135418 422422 135654
rect 422186 135098 422422 135334
rect 422186 99418 422422 99654
rect 422186 99098 422422 99334
rect 422186 63418 422422 63654
rect 422186 63098 422422 63334
rect 422186 27418 422422 27654
rect 422186 27098 422422 27334
rect 422186 -5282 422422 -5046
rect 422186 -5602 422422 -5366
rect 443786 710242 444022 710478
rect 443786 709922 444022 710158
rect 440186 708362 440422 708598
rect 440186 708042 440422 708278
rect 436586 706482 436822 706718
rect 436586 706162 436822 706398
rect 425786 679018 426022 679254
rect 425786 678698 426022 678934
rect 425786 643018 426022 643254
rect 425786 642698 426022 642934
rect 425786 607018 426022 607254
rect 425786 606698 426022 606934
rect 425786 571018 426022 571254
rect 425786 570698 426022 570934
rect 425786 535018 426022 535254
rect 425786 534698 426022 534934
rect 425786 499018 426022 499254
rect 425786 498698 426022 498934
rect 425786 463018 426022 463254
rect 425786 462698 426022 462934
rect 425786 427018 426022 427254
rect 425786 426698 426022 426934
rect 425786 391018 426022 391254
rect 425786 390698 426022 390934
rect 425786 355018 426022 355254
rect 425786 354698 426022 354934
rect 425786 319018 426022 319254
rect 425786 318698 426022 318934
rect 425786 283018 426022 283254
rect 425786 282698 426022 282934
rect 425786 247018 426022 247254
rect 425786 246698 426022 246934
rect 425786 211018 426022 211254
rect 425786 210698 426022 210934
rect 425786 175018 426022 175254
rect 425786 174698 426022 174934
rect 425786 139018 426022 139254
rect 425786 138698 426022 138934
rect 425786 103018 426022 103254
rect 425786 102698 426022 102934
rect 425786 67018 426022 67254
rect 425786 66698 426022 66934
rect 425786 31018 426022 31254
rect 425786 30698 426022 30934
rect 407786 -6222 408022 -5986
rect 407786 -6542 408022 -6306
rect 432986 704602 433222 704838
rect 432986 704282 433222 704518
rect 436586 689818 436822 690054
rect 436586 689498 436822 689734
rect 432986 686218 433222 686454
rect 432986 685898 433222 686134
rect 436586 653818 436822 654054
rect 436586 653498 436822 653734
rect 432986 650218 433222 650454
rect 432986 649898 433222 650134
rect 432986 614218 433222 614454
rect 432986 613898 433222 614134
rect 432986 578218 433222 578454
rect 432986 577898 433222 578134
rect 432986 542218 433222 542454
rect 432986 541898 433222 542134
rect 432986 506218 433222 506454
rect 432986 505898 433222 506134
rect 432986 470218 433222 470454
rect 432986 469898 433222 470134
rect 432986 434218 433222 434454
rect 432986 433898 433222 434134
rect 432986 398218 433222 398454
rect 432986 397898 433222 398134
rect 432986 362218 433222 362454
rect 432986 361898 433222 362134
rect 432986 326218 433222 326454
rect 432986 325898 433222 326134
rect 432986 290218 433222 290454
rect 432986 289898 433222 290134
rect 432986 254218 433222 254454
rect 432986 253898 433222 254134
rect 432986 218218 433222 218454
rect 432986 217898 433222 218134
rect 432986 182218 433222 182454
rect 432986 181898 433222 182134
rect 432986 146218 433222 146454
rect 432986 145898 433222 146134
rect 432986 110218 433222 110454
rect 432986 109898 433222 110134
rect 432986 74218 433222 74454
rect 432986 73898 433222 74134
rect 432986 38218 433222 38454
rect 432986 37898 433222 38134
rect 432986 2218 433222 2454
rect 432986 1898 433222 2134
rect 432986 -582 433222 -346
rect 432986 -902 433222 -666
rect 436586 617818 436822 618054
rect 436586 617498 436822 617734
rect 436586 581818 436822 582054
rect 436586 581498 436822 581734
rect 436586 545818 436822 546054
rect 436586 545498 436822 545734
rect 436586 509818 436822 510054
rect 436586 509498 436822 509734
rect 436586 473818 436822 474054
rect 436586 473498 436822 473734
rect 436586 437818 436822 438054
rect 436586 437498 436822 437734
rect 436586 401818 436822 402054
rect 436586 401498 436822 401734
rect 436586 365818 436822 366054
rect 436586 365498 436822 365734
rect 436586 329818 436822 330054
rect 436586 329498 436822 329734
rect 436586 293818 436822 294054
rect 436586 293498 436822 293734
rect 436586 257818 436822 258054
rect 436586 257498 436822 257734
rect 436586 221818 436822 222054
rect 436586 221498 436822 221734
rect 436586 185818 436822 186054
rect 436586 185498 436822 185734
rect 436586 149818 436822 150054
rect 436586 149498 436822 149734
rect 436586 113818 436822 114054
rect 436586 113498 436822 113734
rect 436586 77818 436822 78054
rect 436586 77498 436822 77734
rect 436586 41818 436822 42054
rect 436586 41498 436822 41734
rect 436586 5818 436822 6054
rect 436586 5498 436822 5734
rect 436586 -2462 436822 -2226
rect 436586 -2782 436822 -2546
rect 440186 693418 440422 693654
rect 440186 693098 440422 693334
rect 440186 657418 440422 657654
rect 440186 657098 440422 657334
rect 440186 621418 440422 621654
rect 440186 621098 440422 621334
rect 440186 585418 440422 585654
rect 440186 585098 440422 585334
rect 440186 549418 440422 549654
rect 440186 549098 440422 549334
rect 440186 513418 440422 513654
rect 440186 513098 440422 513334
rect 440186 477418 440422 477654
rect 440186 477098 440422 477334
rect 440186 441418 440422 441654
rect 440186 441098 440422 441334
rect 440186 405418 440422 405654
rect 440186 405098 440422 405334
rect 440186 369418 440422 369654
rect 440186 369098 440422 369334
rect 440186 333418 440422 333654
rect 440186 333098 440422 333334
rect 440186 297418 440422 297654
rect 440186 297098 440422 297334
rect 440186 261418 440422 261654
rect 440186 261098 440422 261334
rect 440186 225418 440422 225654
rect 440186 225098 440422 225334
rect 440186 189418 440422 189654
rect 440186 189098 440422 189334
rect 440186 153418 440422 153654
rect 440186 153098 440422 153334
rect 440186 117418 440422 117654
rect 440186 117098 440422 117334
rect 440186 81418 440422 81654
rect 440186 81098 440422 81334
rect 440186 45418 440422 45654
rect 440186 45098 440422 45334
rect 440186 9418 440422 9654
rect 440186 9098 440422 9334
rect 440186 -4342 440422 -4106
rect 440186 -4662 440422 -4426
rect 461786 711182 462022 711418
rect 461786 710862 462022 711098
rect 458186 709302 458422 709538
rect 458186 708982 458422 709218
rect 454586 707422 454822 707658
rect 454586 707102 454822 707338
rect 443786 697018 444022 697254
rect 443786 696698 444022 696934
rect 443786 661018 444022 661254
rect 443786 660698 444022 660934
rect 443786 625018 444022 625254
rect 443786 624698 444022 624934
rect 443786 589018 444022 589254
rect 443786 588698 444022 588934
rect 443786 553018 444022 553254
rect 443786 552698 444022 552934
rect 443786 517018 444022 517254
rect 443786 516698 444022 516934
rect 443786 481018 444022 481254
rect 443786 480698 444022 480934
rect 443786 445018 444022 445254
rect 443786 444698 444022 444934
rect 443786 409018 444022 409254
rect 443786 408698 444022 408934
rect 443786 373018 444022 373254
rect 443786 372698 444022 372934
rect 443786 337018 444022 337254
rect 443786 336698 444022 336934
rect 443786 301018 444022 301254
rect 443786 300698 444022 300934
rect 443786 265018 444022 265254
rect 443786 264698 444022 264934
rect 443786 229018 444022 229254
rect 443786 228698 444022 228934
rect 443786 193018 444022 193254
rect 443786 192698 444022 192934
rect 443786 157018 444022 157254
rect 443786 156698 444022 156934
rect 443786 121018 444022 121254
rect 443786 120698 444022 120934
rect 443786 85018 444022 85254
rect 443786 84698 444022 84934
rect 443786 49018 444022 49254
rect 443786 48698 444022 48934
rect 443786 13018 444022 13254
rect 443786 12698 444022 12934
rect 425786 -7162 426022 -6926
rect 425786 -7482 426022 -7246
rect 450986 705542 451222 705778
rect 450986 705222 451222 705458
rect 450986 668218 451222 668454
rect 450986 667898 451222 668134
rect 450986 632218 451222 632454
rect 450986 631898 451222 632134
rect 450986 596218 451222 596454
rect 450986 595898 451222 596134
rect 450986 560218 451222 560454
rect 450986 559898 451222 560134
rect 450986 524218 451222 524454
rect 450986 523898 451222 524134
rect 450986 488218 451222 488454
rect 450986 487898 451222 488134
rect 450986 452218 451222 452454
rect 450986 451898 451222 452134
rect 450986 416218 451222 416454
rect 450986 415898 451222 416134
rect 450986 380218 451222 380454
rect 450986 379898 451222 380134
rect 450986 344218 451222 344454
rect 450986 343898 451222 344134
rect 450986 308218 451222 308454
rect 450986 307898 451222 308134
rect 450986 272218 451222 272454
rect 450986 271898 451222 272134
rect 450986 236218 451222 236454
rect 450986 235898 451222 236134
rect 450986 200218 451222 200454
rect 450986 199898 451222 200134
rect 450986 164218 451222 164454
rect 450986 163898 451222 164134
rect 450986 128218 451222 128454
rect 450986 127898 451222 128134
rect 450986 92218 451222 92454
rect 450986 91898 451222 92134
rect 450986 56218 451222 56454
rect 450986 55898 451222 56134
rect 450986 20218 451222 20454
rect 450986 19898 451222 20134
rect 450986 -1522 451222 -1286
rect 450986 -1842 451222 -1606
rect 454586 671818 454822 672054
rect 454586 671498 454822 671734
rect 454586 635818 454822 636054
rect 454586 635498 454822 635734
rect 454586 599818 454822 600054
rect 454586 599498 454822 599734
rect 454586 563818 454822 564054
rect 454586 563498 454822 563734
rect 454586 527818 454822 528054
rect 454586 527498 454822 527734
rect 454586 491818 454822 492054
rect 454586 491498 454822 491734
rect 454586 455818 454822 456054
rect 454586 455498 454822 455734
rect 454586 419818 454822 420054
rect 454586 419498 454822 419734
rect 454586 383818 454822 384054
rect 454586 383498 454822 383734
rect 454586 347818 454822 348054
rect 454586 347498 454822 347734
rect 454586 311818 454822 312054
rect 454586 311498 454822 311734
rect 454586 275818 454822 276054
rect 454586 275498 454822 275734
rect 454586 239818 454822 240054
rect 454586 239498 454822 239734
rect 454586 203818 454822 204054
rect 454586 203498 454822 203734
rect 454586 167818 454822 168054
rect 454586 167498 454822 167734
rect 454586 131818 454822 132054
rect 454586 131498 454822 131734
rect 454586 95818 454822 96054
rect 454586 95498 454822 95734
rect 454586 59818 454822 60054
rect 454586 59498 454822 59734
rect 454586 23818 454822 24054
rect 454586 23498 454822 23734
rect 454586 -3402 454822 -3166
rect 454586 -3722 454822 -3486
rect 458186 675418 458422 675654
rect 458186 675098 458422 675334
rect 458186 639418 458422 639654
rect 458186 639098 458422 639334
rect 458186 603418 458422 603654
rect 458186 603098 458422 603334
rect 458186 567418 458422 567654
rect 458186 567098 458422 567334
rect 458186 531418 458422 531654
rect 458186 531098 458422 531334
rect 458186 495418 458422 495654
rect 458186 495098 458422 495334
rect 458186 459418 458422 459654
rect 458186 459098 458422 459334
rect 458186 423418 458422 423654
rect 458186 423098 458422 423334
rect 458186 387418 458422 387654
rect 458186 387098 458422 387334
rect 458186 351418 458422 351654
rect 458186 351098 458422 351334
rect 458186 315418 458422 315654
rect 458186 315098 458422 315334
rect 458186 279418 458422 279654
rect 458186 279098 458422 279334
rect 458186 243418 458422 243654
rect 458186 243098 458422 243334
rect 458186 207418 458422 207654
rect 458186 207098 458422 207334
rect 458186 171418 458422 171654
rect 458186 171098 458422 171334
rect 458186 135418 458422 135654
rect 458186 135098 458422 135334
rect 458186 99418 458422 99654
rect 458186 99098 458422 99334
rect 458186 63418 458422 63654
rect 458186 63098 458422 63334
rect 458186 27418 458422 27654
rect 458186 27098 458422 27334
rect 458186 -5282 458422 -5046
rect 458186 -5602 458422 -5366
rect 479786 710242 480022 710478
rect 479786 709922 480022 710158
rect 476186 708362 476422 708598
rect 476186 708042 476422 708278
rect 472586 706482 472822 706718
rect 472586 706162 472822 706398
rect 461786 679018 462022 679254
rect 461786 678698 462022 678934
rect 461786 643018 462022 643254
rect 461786 642698 462022 642934
rect 461786 607018 462022 607254
rect 461786 606698 462022 606934
rect 461786 571018 462022 571254
rect 461786 570698 462022 570934
rect 461786 535018 462022 535254
rect 461786 534698 462022 534934
rect 461786 499018 462022 499254
rect 461786 498698 462022 498934
rect 461786 463018 462022 463254
rect 461786 462698 462022 462934
rect 461786 427018 462022 427254
rect 461786 426698 462022 426934
rect 461786 391018 462022 391254
rect 461786 390698 462022 390934
rect 461786 355018 462022 355254
rect 461786 354698 462022 354934
rect 461786 319018 462022 319254
rect 461786 318698 462022 318934
rect 461786 283018 462022 283254
rect 461786 282698 462022 282934
rect 461786 247018 462022 247254
rect 461786 246698 462022 246934
rect 461786 211018 462022 211254
rect 461786 210698 462022 210934
rect 461786 175018 462022 175254
rect 461786 174698 462022 174934
rect 461786 139018 462022 139254
rect 461786 138698 462022 138934
rect 461786 103018 462022 103254
rect 461786 102698 462022 102934
rect 461786 67018 462022 67254
rect 461786 66698 462022 66934
rect 461786 31018 462022 31254
rect 461786 30698 462022 30934
rect 443786 -6222 444022 -5986
rect 443786 -6542 444022 -6306
rect 468986 704602 469222 704838
rect 468986 704282 469222 704518
rect 468986 686218 469222 686454
rect 468986 685898 469222 686134
rect 468986 650218 469222 650454
rect 468986 649898 469222 650134
rect 468986 614218 469222 614454
rect 468986 613898 469222 614134
rect 468986 578218 469222 578454
rect 468986 577898 469222 578134
rect 468986 542218 469222 542454
rect 468986 541898 469222 542134
rect 468986 506218 469222 506454
rect 468986 505898 469222 506134
rect 468986 470218 469222 470454
rect 468986 469898 469222 470134
rect 468986 434218 469222 434454
rect 468986 433898 469222 434134
rect 468986 398218 469222 398454
rect 468986 397898 469222 398134
rect 468986 362218 469222 362454
rect 468986 361898 469222 362134
rect 468986 326218 469222 326454
rect 468986 325898 469222 326134
rect 468986 290218 469222 290454
rect 468986 289898 469222 290134
rect 468986 254218 469222 254454
rect 468986 253898 469222 254134
rect 468986 218218 469222 218454
rect 468986 217898 469222 218134
rect 468986 182218 469222 182454
rect 468986 181898 469222 182134
rect 468986 146218 469222 146454
rect 468986 145898 469222 146134
rect 468986 110218 469222 110454
rect 468986 109898 469222 110134
rect 468986 74218 469222 74454
rect 468986 73898 469222 74134
rect 468986 38218 469222 38454
rect 468986 37898 469222 38134
rect 468986 2218 469222 2454
rect 468986 1898 469222 2134
rect 468986 -582 469222 -346
rect 468986 -902 469222 -666
rect 472586 689818 472822 690054
rect 472586 689498 472822 689734
rect 472586 653818 472822 654054
rect 472586 653498 472822 653734
rect 472586 617818 472822 618054
rect 472586 617498 472822 617734
rect 472586 581818 472822 582054
rect 472586 581498 472822 581734
rect 472586 545818 472822 546054
rect 472586 545498 472822 545734
rect 472586 509818 472822 510054
rect 472586 509498 472822 509734
rect 472586 473818 472822 474054
rect 472586 473498 472822 473734
rect 472586 437818 472822 438054
rect 472586 437498 472822 437734
rect 472586 401818 472822 402054
rect 472586 401498 472822 401734
rect 472586 365818 472822 366054
rect 472586 365498 472822 365734
rect 472586 329818 472822 330054
rect 472586 329498 472822 329734
rect 472586 293818 472822 294054
rect 472586 293498 472822 293734
rect 472586 257818 472822 258054
rect 472586 257498 472822 257734
rect 472586 221818 472822 222054
rect 472586 221498 472822 221734
rect 472586 185818 472822 186054
rect 472586 185498 472822 185734
rect 472586 149818 472822 150054
rect 472586 149498 472822 149734
rect 472586 113818 472822 114054
rect 472586 113498 472822 113734
rect 472586 77818 472822 78054
rect 472586 77498 472822 77734
rect 472586 41818 472822 42054
rect 472586 41498 472822 41734
rect 472586 5818 472822 6054
rect 472586 5498 472822 5734
rect 472586 -2462 472822 -2226
rect 472586 -2782 472822 -2546
rect 476186 693418 476422 693654
rect 476186 693098 476422 693334
rect 476186 657418 476422 657654
rect 476186 657098 476422 657334
rect 476186 621418 476422 621654
rect 476186 621098 476422 621334
rect 476186 585418 476422 585654
rect 476186 585098 476422 585334
rect 476186 549418 476422 549654
rect 476186 549098 476422 549334
rect 476186 513418 476422 513654
rect 476186 513098 476422 513334
rect 476186 477418 476422 477654
rect 476186 477098 476422 477334
rect 476186 441418 476422 441654
rect 476186 441098 476422 441334
rect 476186 405418 476422 405654
rect 476186 405098 476422 405334
rect 476186 369418 476422 369654
rect 476186 369098 476422 369334
rect 476186 333418 476422 333654
rect 476186 333098 476422 333334
rect 476186 297418 476422 297654
rect 476186 297098 476422 297334
rect 476186 261418 476422 261654
rect 476186 261098 476422 261334
rect 476186 225418 476422 225654
rect 476186 225098 476422 225334
rect 476186 189418 476422 189654
rect 476186 189098 476422 189334
rect 476186 153418 476422 153654
rect 476186 153098 476422 153334
rect 476186 117418 476422 117654
rect 476186 117098 476422 117334
rect 476186 81418 476422 81654
rect 476186 81098 476422 81334
rect 476186 45418 476422 45654
rect 476186 45098 476422 45334
rect 476186 9418 476422 9654
rect 476186 9098 476422 9334
rect 476186 -4342 476422 -4106
rect 476186 -4662 476422 -4426
rect 497786 711182 498022 711418
rect 497786 710862 498022 711098
rect 494186 709302 494422 709538
rect 494186 708982 494422 709218
rect 490586 707422 490822 707658
rect 490586 707102 490822 707338
rect 479786 697018 480022 697254
rect 479786 696698 480022 696934
rect 479786 661018 480022 661254
rect 479786 660698 480022 660934
rect 479786 625018 480022 625254
rect 479786 624698 480022 624934
rect 479786 589018 480022 589254
rect 479786 588698 480022 588934
rect 479786 553018 480022 553254
rect 479786 552698 480022 552934
rect 479786 517018 480022 517254
rect 479786 516698 480022 516934
rect 479786 481018 480022 481254
rect 479786 480698 480022 480934
rect 479786 445018 480022 445254
rect 479786 444698 480022 444934
rect 479786 409018 480022 409254
rect 479786 408698 480022 408934
rect 479786 373018 480022 373254
rect 479786 372698 480022 372934
rect 479786 337018 480022 337254
rect 479786 336698 480022 336934
rect 479786 301018 480022 301254
rect 479786 300698 480022 300934
rect 479786 265018 480022 265254
rect 479786 264698 480022 264934
rect 479786 229018 480022 229254
rect 479786 228698 480022 228934
rect 479786 193018 480022 193254
rect 479786 192698 480022 192934
rect 479786 157018 480022 157254
rect 479786 156698 480022 156934
rect 479786 121018 480022 121254
rect 479786 120698 480022 120934
rect 479786 85018 480022 85254
rect 479786 84698 480022 84934
rect 479786 49018 480022 49254
rect 479786 48698 480022 48934
rect 479786 13018 480022 13254
rect 479786 12698 480022 12934
rect 461786 -7162 462022 -6926
rect 461786 -7482 462022 -7246
rect 486986 705542 487222 705778
rect 486986 705222 487222 705458
rect 486986 668218 487222 668454
rect 486986 667898 487222 668134
rect 486986 632218 487222 632454
rect 486986 631898 487222 632134
rect 486986 596218 487222 596454
rect 486986 595898 487222 596134
rect 486986 560218 487222 560454
rect 486986 559898 487222 560134
rect 486986 524218 487222 524454
rect 486986 523898 487222 524134
rect 486986 488218 487222 488454
rect 486986 487898 487222 488134
rect 486986 452218 487222 452454
rect 486986 451898 487222 452134
rect 486986 416218 487222 416454
rect 486986 415898 487222 416134
rect 486986 380218 487222 380454
rect 486986 379898 487222 380134
rect 486986 344218 487222 344454
rect 486986 343898 487222 344134
rect 486986 308218 487222 308454
rect 486986 307898 487222 308134
rect 486986 272218 487222 272454
rect 486986 271898 487222 272134
rect 486986 236218 487222 236454
rect 486986 235898 487222 236134
rect 486986 200218 487222 200454
rect 486986 199898 487222 200134
rect 486986 164218 487222 164454
rect 486986 163898 487222 164134
rect 486986 128218 487222 128454
rect 486986 127898 487222 128134
rect 486986 92218 487222 92454
rect 486986 91898 487222 92134
rect 486986 56218 487222 56454
rect 486986 55898 487222 56134
rect 486986 20218 487222 20454
rect 486986 19898 487222 20134
rect 486986 -1522 487222 -1286
rect 486986 -1842 487222 -1606
rect 490586 671818 490822 672054
rect 490586 671498 490822 671734
rect 490586 635818 490822 636054
rect 490586 635498 490822 635734
rect 490586 599818 490822 600054
rect 490586 599498 490822 599734
rect 490586 563818 490822 564054
rect 490586 563498 490822 563734
rect 494186 675418 494422 675654
rect 494186 675098 494422 675334
rect 494186 639418 494422 639654
rect 494186 639098 494422 639334
rect 494186 603418 494422 603654
rect 494186 603098 494422 603334
rect 494186 567418 494422 567654
rect 494186 567098 494422 567334
rect 490586 527818 490822 528054
rect 490586 527498 490822 527734
rect 490586 491818 490822 492054
rect 490586 491498 490822 491734
rect 490586 455818 490822 456054
rect 490586 455498 490822 455734
rect 490586 419818 490822 420054
rect 490586 419498 490822 419734
rect 490586 383818 490822 384054
rect 490586 383498 490822 383734
rect 490586 347818 490822 348054
rect 490586 347498 490822 347734
rect 490586 311818 490822 312054
rect 490586 311498 490822 311734
rect 490586 275818 490822 276054
rect 490586 275498 490822 275734
rect 490586 239818 490822 240054
rect 490586 239498 490822 239734
rect 490586 203818 490822 204054
rect 490586 203498 490822 203734
rect 490586 167818 490822 168054
rect 490586 167498 490822 167734
rect 490586 131818 490822 132054
rect 490586 131498 490822 131734
rect 490586 95818 490822 96054
rect 490586 95498 490822 95734
rect 490586 59818 490822 60054
rect 490586 59498 490822 59734
rect 490586 23818 490822 24054
rect 490586 23498 490822 23734
rect 490586 -3402 490822 -3166
rect 490586 -3722 490822 -3486
rect 494186 531418 494422 531654
rect 494186 531098 494422 531334
rect 494186 495418 494422 495654
rect 494186 495098 494422 495334
rect 494186 459418 494422 459654
rect 494186 459098 494422 459334
rect 494186 423418 494422 423654
rect 494186 423098 494422 423334
rect 494186 387418 494422 387654
rect 494186 387098 494422 387334
rect 494186 351418 494422 351654
rect 494186 351098 494422 351334
rect 494186 315418 494422 315654
rect 494186 315098 494422 315334
rect 494186 279418 494422 279654
rect 494186 279098 494422 279334
rect 494186 243418 494422 243654
rect 494186 243098 494422 243334
rect 494186 207418 494422 207654
rect 494186 207098 494422 207334
rect 494186 171418 494422 171654
rect 494186 171098 494422 171334
rect 494186 135418 494422 135654
rect 494186 135098 494422 135334
rect 494186 99418 494422 99654
rect 494186 99098 494422 99334
rect 494186 63418 494422 63654
rect 494186 63098 494422 63334
rect 494186 27418 494422 27654
rect 494186 27098 494422 27334
rect 494186 -5282 494422 -5046
rect 494186 -5602 494422 -5366
rect 515786 710242 516022 710478
rect 515786 709922 516022 710158
rect 512186 708362 512422 708598
rect 512186 708042 512422 708278
rect 508586 706482 508822 706718
rect 508586 706162 508822 706398
rect 497786 679018 498022 679254
rect 497786 678698 498022 678934
rect 497786 643018 498022 643254
rect 497786 642698 498022 642934
rect 497786 607018 498022 607254
rect 497786 606698 498022 606934
rect 497786 571018 498022 571254
rect 497786 570698 498022 570934
rect 497786 535018 498022 535254
rect 497786 534698 498022 534934
rect 497786 499018 498022 499254
rect 497786 498698 498022 498934
rect 497786 463018 498022 463254
rect 497786 462698 498022 462934
rect 497786 427018 498022 427254
rect 497786 426698 498022 426934
rect 497786 391018 498022 391254
rect 497786 390698 498022 390934
rect 497786 355018 498022 355254
rect 497786 354698 498022 354934
rect 497786 319018 498022 319254
rect 497786 318698 498022 318934
rect 497786 283018 498022 283254
rect 497786 282698 498022 282934
rect 497786 247018 498022 247254
rect 497786 246698 498022 246934
rect 497786 211018 498022 211254
rect 497786 210698 498022 210934
rect 497786 175018 498022 175254
rect 497786 174698 498022 174934
rect 497786 139018 498022 139254
rect 497786 138698 498022 138934
rect 497786 103018 498022 103254
rect 497786 102698 498022 102934
rect 497786 67018 498022 67254
rect 497786 66698 498022 66934
rect 497786 31018 498022 31254
rect 497786 30698 498022 30934
rect 479786 -6222 480022 -5986
rect 479786 -6542 480022 -6306
rect 504986 704602 505222 704838
rect 504986 704282 505222 704518
rect 504986 686218 505222 686454
rect 504986 685898 505222 686134
rect 504986 650218 505222 650454
rect 504986 649898 505222 650134
rect 504986 614218 505222 614454
rect 504986 613898 505222 614134
rect 504986 578218 505222 578454
rect 504986 577898 505222 578134
rect 504986 542218 505222 542454
rect 504986 541898 505222 542134
rect 504986 506218 505222 506454
rect 504986 505898 505222 506134
rect 504986 470218 505222 470454
rect 504986 469898 505222 470134
rect 504986 434218 505222 434454
rect 504986 433898 505222 434134
rect 504986 398218 505222 398454
rect 504986 397898 505222 398134
rect 504986 362218 505222 362454
rect 504986 361898 505222 362134
rect 504986 326218 505222 326454
rect 504986 325898 505222 326134
rect 504986 290218 505222 290454
rect 504986 289898 505222 290134
rect 504986 254218 505222 254454
rect 504986 253898 505222 254134
rect 504986 218218 505222 218454
rect 504986 217898 505222 218134
rect 504986 182218 505222 182454
rect 504986 181898 505222 182134
rect 504986 146218 505222 146454
rect 504986 145898 505222 146134
rect 504986 110218 505222 110454
rect 504986 109898 505222 110134
rect 504986 74218 505222 74454
rect 504986 73898 505222 74134
rect 504986 38218 505222 38454
rect 504986 37898 505222 38134
rect 504986 2218 505222 2454
rect 504986 1898 505222 2134
rect 504986 -582 505222 -346
rect 504986 -902 505222 -666
rect 508586 689818 508822 690054
rect 508586 689498 508822 689734
rect 508586 653818 508822 654054
rect 508586 653498 508822 653734
rect 508586 617818 508822 618054
rect 508586 617498 508822 617734
rect 508586 581818 508822 582054
rect 508586 581498 508822 581734
rect 508586 545818 508822 546054
rect 508586 545498 508822 545734
rect 508586 509818 508822 510054
rect 508586 509498 508822 509734
rect 508586 473818 508822 474054
rect 508586 473498 508822 473734
rect 508586 437818 508822 438054
rect 508586 437498 508822 437734
rect 508586 401818 508822 402054
rect 508586 401498 508822 401734
rect 508586 365818 508822 366054
rect 508586 365498 508822 365734
rect 508586 329818 508822 330054
rect 508586 329498 508822 329734
rect 508586 293818 508822 294054
rect 508586 293498 508822 293734
rect 508586 257818 508822 258054
rect 508586 257498 508822 257734
rect 508586 221818 508822 222054
rect 508586 221498 508822 221734
rect 508586 185818 508822 186054
rect 508586 185498 508822 185734
rect 508586 149818 508822 150054
rect 508586 149498 508822 149734
rect 508586 113818 508822 114054
rect 508586 113498 508822 113734
rect 508586 77818 508822 78054
rect 508586 77498 508822 77734
rect 508586 41818 508822 42054
rect 508586 41498 508822 41734
rect 508586 5818 508822 6054
rect 508586 5498 508822 5734
rect 508586 -2462 508822 -2226
rect 508586 -2782 508822 -2546
rect 512186 693418 512422 693654
rect 512186 693098 512422 693334
rect 512186 657418 512422 657654
rect 512186 657098 512422 657334
rect 512186 621418 512422 621654
rect 512186 621098 512422 621334
rect 512186 585418 512422 585654
rect 512186 585098 512422 585334
rect 512186 549418 512422 549654
rect 512186 549098 512422 549334
rect 512186 513418 512422 513654
rect 512186 513098 512422 513334
rect 512186 477418 512422 477654
rect 512186 477098 512422 477334
rect 512186 441418 512422 441654
rect 512186 441098 512422 441334
rect 512186 405418 512422 405654
rect 512186 405098 512422 405334
rect 512186 369418 512422 369654
rect 512186 369098 512422 369334
rect 512186 333418 512422 333654
rect 512186 333098 512422 333334
rect 512186 297418 512422 297654
rect 512186 297098 512422 297334
rect 512186 261418 512422 261654
rect 512186 261098 512422 261334
rect 512186 225418 512422 225654
rect 512186 225098 512422 225334
rect 512186 189418 512422 189654
rect 512186 189098 512422 189334
rect 512186 153418 512422 153654
rect 512186 153098 512422 153334
rect 512186 117418 512422 117654
rect 512186 117098 512422 117334
rect 512186 81418 512422 81654
rect 512186 81098 512422 81334
rect 512186 45418 512422 45654
rect 512186 45098 512422 45334
rect 512186 9418 512422 9654
rect 512186 9098 512422 9334
rect 512186 -4342 512422 -4106
rect 512186 -4662 512422 -4426
rect 533786 711182 534022 711418
rect 533786 710862 534022 711098
rect 530186 709302 530422 709538
rect 530186 708982 530422 709218
rect 526586 707422 526822 707658
rect 526586 707102 526822 707338
rect 515786 697018 516022 697254
rect 515786 696698 516022 696934
rect 515786 661018 516022 661254
rect 515786 660698 516022 660934
rect 515786 625018 516022 625254
rect 515786 624698 516022 624934
rect 515786 589018 516022 589254
rect 515786 588698 516022 588934
rect 515786 553018 516022 553254
rect 515786 552698 516022 552934
rect 515786 517018 516022 517254
rect 515786 516698 516022 516934
rect 515786 481018 516022 481254
rect 515786 480698 516022 480934
rect 515786 445018 516022 445254
rect 515786 444698 516022 444934
rect 515786 409018 516022 409254
rect 515786 408698 516022 408934
rect 515786 373018 516022 373254
rect 515786 372698 516022 372934
rect 515786 337018 516022 337254
rect 515786 336698 516022 336934
rect 515786 301018 516022 301254
rect 515786 300698 516022 300934
rect 515786 265018 516022 265254
rect 515786 264698 516022 264934
rect 515786 229018 516022 229254
rect 515786 228698 516022 228934
rect 515786 193018 516022 193254
rect 515786 192698 516022 192934
rect 515786 157018 516022 157254
rect 515786 156698 516022 156934
rect 515786 121018 516022 121254
rect 515786 120698 516022 120934
rect 515786 85018 516022 85254
rect 515786 84698 516022 84934
rect 515786 49018 516022 49254
rect 515786 48698 516022 48934
rect 515786 13018 516022 13254
rect 515786 12698 516022 12934
rect 497786 -7162 498022 -6926
rect 497786 -7482 498022 -7246
rect 522986 705542 523222 705778
rect 522986 705222 523222 705458
rect 522986 668218 523222 668454
rect 522986 667898 523222 668134
rect 522986 632218 523222 632454
rect 522986 631898 523222 632134
rect 522986 596218 523222 596454
rect 522986 595898 523222 596134
rect 522986 560218 523222 560454
rect 522986 559898 523222 560134
rect 522986 524218 523222 524454
rect 522986 523898 523222 524134
rect 522986 488218 523222 488454
rect 522986 487898 523222 488134
rect 522986 452218 523222 452454
rect 522986 451898 523222 452134
rect 522986 416218 523222 416454
rect 522986 415898 523222 416134
rect 522986 380218 523222 380454
rect 522986 379898 523222 380134
rect 522986 344218 523222 344454
rect 522986 343898 523222 344134
rect 522986 308218 523222 308454
rect 522986 307898 523222 308134
rect 522986 272218 523222 272454
rect 522986 271898 523222 272134
rect 522986 236218 523222 236454
rect 522986 235898 523222 236134
rect 522986 200218 523222 200454
rect 522986 199898 523222 200134
rect 522986 164218 523222 164454
rect 522986 163898 523222 164134
rect 522986 128218 523222 128454
rect 522986 127898 523222 128134
rect 522986 92218 523222 92454
rect 522986 91898 523222 92134
rect 522986 56218 523222 56454
rect 522986 55898 523222 56134
rect 522986 20218 523222 20454
rect 522986 19898 523222 20134
rect 522986 -1522 523222 -1286
rect 522986 -1842 523222 -1606
rect 526586 671818 526822 672054
rect 526586 671498 526822 671734
rect 526586 635818 526822 636054
rect 526586 635498 526822 635734
rect 526586 599818 526822 600054
rect 526586 599498 526822 599734
rect 526586 563818 526822 564054
rect 526586 563498 526822 563734
rect 526586 527818 526822 528054
rect 526586 527498 526822 527734
rect 526586 491818 526822 492054
rect 526586 491498 526822 491734
rect 526586 455818 526822 456054
rect 526586 455498 526822 455734
rect 526586 419818 526822 420054
rect 526586 419498 526822 419734
rect 526586 383818 526822 384054
rect 526586 383498 526822 383734
rect 526586 347818 526822 348054
rect 526586 347498 526822 347734
rect 526586 311818 526822 312054
rect 526586 311498 526822 311734
rect 526586 275818 526822 276054
rect 526586 275498 526822 275734
rect 526586 239818 526822 240054
rect 526586 239498 526822 239734
rect 526586 203818 526822 204054
rect 526586 203498 526822 203734
rect 526586 167818 526822 168054
rect 526586 167498 526822 167734
rect 526586 131818 526822 132054
rect 526586 131498 526822 131734
rect 526586 95818 526822 96054
rect 526586 95498 526822 95734
rect 526586 59818 526822 60054
rect 526586 59498 526822 59734
rect 526586 23818 526822 24054
rect 526586 23498 526822 23734
rect 526586 -3402 526822 -3166
rect 526586 -3722 526822 -3486
rect 530186 675418 530422 675654
rect 530186 675098 530422 675334
rect 530186 639418 530422 639654
rect 530186 639098 530422 639334
rect 530186 603418 530422 603654
rect 530186 603098 530422 603334
rect 530186 567418 530422 567654
rect 530186 567098 530422 567334
rect 530186 531418 530422 531654
rect 530186 531098 530422 531334
rect 530186 495418 530422 495654
rect 530186 495098 530422 495334
rect 530186 459418 530422 459654
rect 530186 459098 530422 459334
rect 530186 423418 530422 423654
rect 530186 423098 530422 423334
rect 530186 387418 530422 387654
rect 530186 387098 530422 387334
rect 530186 351418 530422 351654
rect 530186 351098 530422 351334
rect 530186 315418 530422 315654
rect 530186 315098 530422 315334
rect 530186 279418 530422 279654
rect 530186 279098 530422 279334
rect 530186 243418 530422 243654
rect 530186 243098 530422 243334
rect 530186 207418 530422 207654
rect 530186 207098 530422 207334
rect 530186 171418 530422 171654
rect 530186 171098 530422 171334
rect 530186 135418 530422 135654
rect 530186 135098 530422 135334
rect 530186 99418 530422 99654
rect 530186 99098 530422 99334
rect 530186 63418 530422 63654
rect 530186 63098 530422 63334
rect 530186 27418 530422 27654
rect 530186 27098 530422 27334
rect 530186 -5282 530422 -5046
rect 530186 -5602 530422 -5366
rect 551786 710242 552022 710478
rect 551786 709922 552022 710158
rect 548186 708362 548422 708598
rect 548186 708042 548422 708278
rect 544586 706482 544822 706718
rect 544586 706162 544822 706398
rect 533786 679018 534022 679254
rect 533786 678698 534022 678934
rect 533786 643018 534022 643254
rect 533786 642698 534022 642934
rect 533786 607018 534022 607254
rect 533786 606698 534022 606934
rect 533786 571018 534022 571254
rect 533786 570698 534022 570934
rect 533786 535018 534022 535254
rect 533786 534698 534022 534934
rect 533786 499018 534022 499254
rect 533786 498698 534022 498934
rect 533786 463018 534022 463254
rect 533786 462698 534022 462934
rect 533786 427018 534022 427254
rect 533786 426698 534022 426934
rect 533786 391018 534022 391254
rect 533786 390698 534022 390934
rect 533786 355018 534022 355254
rect 533786 354698 534022 354934
rect 533786 319018 534022 319254
rect 533786 318698 534022 318934
rect 533786 283018 534022 283254
rect 533786 282698 534022 282934
rect 533786 247018 534022 247254
rect 533786 246698 534022 246934
rect 533786 211018 534022 211254
rect 533786 210698 534022 210934
rect 533786 175018 534022 175254
rect 533786 174698 534022 174934
rect 533786 139018 534022 139254
rect 533786 138698 534022 138934
rect 533786 103018 534022 103254
rect 533786 102698 534022 102934
rect 533786 67018 534022 67254
rect 533786 66698 534022 66934
rect 533786 31018 534022 31254
rect 533786 30698 534022 30934
rect 515786 -6222 516022 -5986
rect 515786 -6542 516022 -6306
rect 540986 704602 541222 704838
rect 540986 704282 541222 704518
rect 540986 686218 541222 686454
rect 540986 685898 541222 686134
rect 540986 650218 541222 650454
rect 540986 649898 541222 650134
rect 540986 614218 541222 614454
rect 540986 613898 541222 614134
rect 540986 578218 541222 578454
rect 540986 577898 541222 578134
rect 540986 542218 541222 542454
rect 540986 541898 541222 542134
rect 540986 506218 541222 506454
rect 540986 505898 541222 506134
rect 540986 470218 541222 470454
rect 540986 469898 541222 470134
rect 540986 434218 541222 434454
rect 540986 433898 541222 434134
rect 540986 398218 541222 398454
rect 540986 397898 541222 398134
rect 540986 362218 541222 362454
rect 540986 361898 541222 362134
rect 540986 326218 541222 326454
rect 540986 325898 541222 326134
rect 540986 290218 541222 290454
rect 540986 289898 541222 290134
rect 540986 254218 541222 254454
rect 540986 253898 541222 254134
rect 540986 218218 541222 218454
rect 540986 217898 541222 218134
rect 540986 182218 541222 182454
rect 540986 181898 541222 182134
rect 540986 146218 541222 146454
rect 540986 145898 541222 146134
rect 540986 110218 541222 110454
rect 540986 109898 541222 110134
rect 540986 74218 541222 74454
rect 540986 73898 541222 74134
rect 540986 38218 541222 38454
rect 540986 37898 541222 38134
rect 540986 2218 541222 2454
rect 540986 1898 541222 2134
rect 540986 -582 541222 -346
rect 540986 -902 541222 -666
rect 544586 689818 544822 690054
rect 544586 689498 544822 689734
rect 544586 653818 544822 654054
rect 544586 653498 544822 653734
rect 544586 617818 544822 618054
rect 544586 617498 544822 617734
rect 544586 581818 544822 582054
rect 544586 581498 544822 581734
rect 544586 545818 544822 546054
rect 544586 545498 544822 545734
rect 544586 509818 544822 510054
rect 544586 509498 544822 509734
rect 544586 473818 544822 474054
rect 544586 473498 544822 473734
rect 544586 437818 544822 438054
rect 544586 437498 544822 437734
rect 544586 401818 544822 402054
rect 544586 401498 544822 401734
rect 544586 365818 544822 366054
rect 544586 365498 544822 365734
rect 544586 329818 544822 330054
rect 544586 329498 544822 329734
rect 544586 293818 544822 294054
rect 544586 293498 544822 293734
rect 544586 257818 544822 258054
rect 544586 257498 544822 257734
rect 544586 221818 544822 222054
rect 544586 221498 544822 221734
rect 544586 185818 544822 186054
rect 544586 185498 544822 185734
rect 544586 149818 544822 150054
rect 544586 149498 544822 149734
rect 544586 113818 544822 114054
rect 544586 113498 544822 113734
rect 544586 77818 544822 78054
rect 544586 77498 544822 77734
rect 544586 41818 544822 42054
rect 544586 41498 544822 41734
rect 544586 5818 544822 6054
rect 544586 5498 544822 5734
rect 544586 -2462 544822 -2226
rect 544586 -2782 544822 -2546
rect 569786 711182 570022 711418
rect 569786 710862 570022 711098
rect 566186 709302 566422 709538
rect 566186 708982 566422 709218
rect 562586 707422 562822 707658
rect 562586 707102 562822 707338
rect 551786 697018 552022 697254
rect 548186 693418 548422 693654
rect 548186 693098 548422 693334
rect 551786 696698 552022 696934
rect 548186 657418 548422 657654
rect 548186 657098 548422 657334
rect 548186 621418 548422 621654
rect 548186 621098 548422 621334
rect 548186 585418 548422 585654
rect 548186 585098 548422 585334
rect 548186 549418 548422 549654
rect 548186 549098 548422 549334
rect 551786 661018 552022 661254
rect 551786 660698 552022 660934
rect 551786 625018 552022 625254
rect 551786 624698 552022 624934
rect 551786 589018 552022 589254
rect 551786 588698 552022 588934
rect 551786 553018 552022 553254
rect 551786 552698 552022 552934
rect 548186 513418 548422 513654
rect 548186 513098 548422 513334
rect 548186 477418 548422 477654
rect 548186 477098 548422 477334
rect 548186 441418 548422 441654
rect 548186 441098 548422 441334
rect 548186 405418 548422 405654
rect 548186 405098 548422 405334
rect 548186 369418 548422 369654
rect 548186 369098 548422 369334
rect 548186 333418 548422 333654
rect 548186 333098 548422 333334
rect 548186 297418 548422 297654
rect 548186 297098 548422 297334
rect 548186 261418 548422 261654
rect 548186 261098 548422 261334
rect 548186 225418 548422 225654
rect 548186 225098 548422 225334
rect 548186 189418 548422 189654
rect 548186 189098 548422 189334
rect 548186 153418 548422 153654
rect 548186 153098 548422 153334
rect 548186 117418 548422 117654
rect 548186 117098 548422 117334
rect 548186 81418 548422 81654
rect 548186 81098 548422 81334
rect 548186 45418 548422 45654
rect 548186 45098 548422 45334
rect 548186 9418 548422 9654
rect 548186 9098 548422 9334
rect 548186 -4342 548422 -4106
rect 548186 -4662 548422 -4426
rect 551786 517018 552022 517254
rect 551786 516698 552022 516934
rect 551786 481018 552022 481254
rect 551786 480698 552022 480934
rect 551786 445018 552022 445254
rect 551786 444698 552022 444934
rect 551786 409018 552022 409254
rect 551786 408698 552022 408934
rect 551786 373018 552022 373254
rect 551786 372698 552022 372934
rect 551786 337018 552022 337254
rect 551786 336698 552022 336934
rect 551786 301018 552022 301254
rect 551786 300698 552022 300934
rect 551786 265018 552022 265254
rect 551786 264698 552022 264934
rect 551786 229018 552022 229254
rect 551786 228698 552022 228934
rect 551786 193018 552022 193254
rect 551786 192698 552022 192934
rect 551786 157018 552022 157254
rect 551786 156698 552022 156934
rect 551786 121018 552022 121254
rect 551786 120698 552022 120934
rect 551786 85018 552022 85254
rect 551786 84698 552022 84934
rect 551786 49018 552022 49254
rect 551786 48698 552022 48934
rect 551786 13018 552022 13254
rect 551786 12698 552022 12934
rect 533786 -7162 534022 -6926
rect 533786 -7482 534022 -7246
rect 558986 705542 559222 705778
rect 558986 705222 559222 705458
rect 558986 668218 559222 668454
rect 558986 667898 559222 668134
rect 558986 632218 559222 632454
rect 558986 631898 559222 632134
rect 558986 596218 559222 596454
rect 558986 595898 559222 596134
rect 558986 560218 559222 560454
rect 558986 559898 559222 560134
rect 558986 524218 559222 524454
rect 558986 523898 559222 524134
rect 558986 488218 559222 488454
rect 558986 487898 559222 488134
rect 558986 452218 559222 452454
rect 558986 451898 559222 452134
rect 558986 416218 559222 416454
rect 558986 415898 559222 416134
rect 558986 380218 559222 380454
rect 558986 379898 559222 380134
rect 558986 344218 559222 344454
rect 558986 343898 559222 344134
rect 558986 308218 559222 308454
rect 558986 307898 559222 308134
rect 558986 272218 559222 272454
rect 558986 271898 559222 272134
rect 558986 236218 559222 236454
rect 558986 235898 559222 236134
rect 558986 200218 559222 200454
rect 558986 199898 559222 200134
rect 558986 164218 559222 164454
rect 558986 163898 559222 164134
rect 558986 128218 559222 128454
rect 558986 127898 559222 128134
rect 558986 92218 559222 92454
rect 558986 91898 559222 92134
rect 558986 56218 559222 56454
rect 558986 55898 559222 56134
rect 558986 20218 559222 20454
rect 558986 19898 559222 20134
rect 558986 -1522 559222 -1286
rect 558986 -1842 559222 -1606
rect 562586 671818 562822 672054
rect 562586 671498 562822 671734
rect 562586 635818 562822 636054
rect 562586 635498 562822 635734
rect 562586 599818 562822 600054
rect 562586 599498 562822 599734
rect 562586 563818 562822 564054
rect 562586 563498 562822 563734
rect 562586 527818 562822 528054
rect 562586 527498 562822 527734
rect 562586 491818 562822 492054
rect 562586 491498 562822 491734
rect 562586 455818 562822 456054
rect 562586 455498 562822 455734
rect 562586 419818 562822 420054
rect 562586 419498 562822 419734
rect 562586 383818 562822 384054
rect 562586 383498 562822 383734
rect 562586 347818 562822 348054
rect 562586 347498 562822 347734
rect 562586 311818 562822 312054
rect 562586 311498 562822 311734
rect 562586 275818 562822 276054
rect 562586 275498 562822 275734
rect 562586 239818 562822 240054
rect 562586 239498 562822 239734
rect 562586 203818 562822 204054
rect 562586 203498 562822 203734
rect 562586 167818 562822 168054
rect 562586 167498 562822 167734
rect 562586 131818 562822 132054
rect 562586 131498 562822 131734
rect 562586 95818 562822 96054
rect 562586 95498 562822 95734
rect 562586 59818 562822 60054
rect 562586 59498 562822 59734
rect 562586 23818 562822 24054
rect 562586 23498 562822 23734
rect 562586 -3402 562822 -3166
rect 562586 -3722 562822 -3486
rect 566186 675418 566422 675654
rect 566186 675098 566422 675334
rect 566186 639418 566422 639654
rect 566186 639098 566422 639334
rect 566186 603418 566422 603654
rect 566186 603098 566422 603334
rect 566186 567418 566422 567654
rect 566186 567098 566422 567334
rect 566186 531418 566422 531654
rect 566186 531098 566422 531334
rect 566186 495418 566422 495654
rect 566186 495098 566422 495334
rect 566186 459418 566422 459654
rect 566186 459098 566422 459334
rect 566186 423418 566422 423654
rect 566186 423098 566422 423334
rect 566186 387418 566422 387654
rect 566186 387098 566422 387334
rect 566186 351418 566422 351654
rect 566186 351098 566422 351334
rect 566186 315418 566422 315654
rect 566186 315098 566422 315334
rect 566186 279418 566422 279654
rect 566186 279098 566422 279334
rect 566186 243418 566422 243654
rect 566186 243098 566422 243334
rect 566186 207418 566422 207654
rect 566186 207098 566422 207334
rect 566186 171418 566422 171654
rect 566186 171098 566422 171334
rect 566186 135418 566422 135654
rect 566186 135098 566422 135334
rect 566186 99418 566422 99654
rect 566186 99098 566422 99334
rect 566186 63418 566422 63654
rect 566186 63098 566422 63334
rect 566186 27418 566422 27654
rect 566186 27098 566422 27334
rect 566186 -5282 566422 -5046
rect 566186 -5602 566422 -5366
rect 592082 711182 592318 711418
rect 592082 710862 592318 711098
rect 591142 710242 591378 710478
rect 591142 709922 591378 710158
rect 590202 709302 590438 709538
rect 590202 708982 590438 709218
rect 589262 708362 589498 708598
rect 589262 708042 589498 708278
rect 588322 707422 588558 707658
rect 588322 707102 588558 707338
rect 580586 706482 580822 706718
rect 580586 706162 580822 706398
rect 569786 679018 570022 679254
rect 569786 678698 570022 678934
rect 569786 643018 570022 643254
rect 569786 642698 570022 642934
rect 569786 607018 570022 607254
rect 569786 606698 570022 606934
rect 569786 571018 570022 571254
rect 569786 570698 570022 570934
rect 569786 535018 570022 535254
rect 569786 534698 570022 534934
rect 569786 499018 570022 499254
rect 569786 498698 570022 498934
rect 569786 463018 570022 463254
rect 569786 462698 570022 462934
rect 569786 427018 570022 427254
rect 569786 426698 570022 426934
rect 569786 391018 570022 391254
rect 569786 390698 570022 390934
rect 569786 355018 570022 355254
rect 569786 354698 570022 354934
rect 569786 319018 570022 319254
rect 569786 318698 570022 318934
rect 569786 283018 570022 283254
rect 569786 282698 570022 282934
rect 569786 247018 570022 247254
rect 569786 246698 570022 246934
rect 569786 211018 570022 211254
rect 569786 210698 570022 210934
rect 569786 175018 570022 175254
rect 569786 174698 570022 174934
rect 569786 139018 570022 139254
rect 569786 138698 570022 138934
rect 569786 103018 570022 103254
rect 569786 102698 570022 102934
rect 569786 67018 570022 67254
rect 569786 66698 570022 66934
rect 569786 31018 570022 31254
rect 569786 30698 570022 30934
rect 551786 -6222 552022 -5986
rect 551786 -6542 552022 -6306
rect 576986 704602 577222 704838
rect 576986 704282 577222 704518
rect 576986 686218 577222 686454
rect 576986 685898 577222 686134
rect 587382 706482 587618 706718
rect 587382 706162 587618 706398
rect 586442 705542 586678 705778
rect 586442 705222 586678 705458
rect 580586 689818 580822 690054
rect 580586 689498 580822 689734
rect 580586 653818 580822 654054
rect 580586 653498 580822 653734
rect 576986 650218 577222 650454
rect 576986 649898 577222 650134
rect 576986 614218 577222 614454
rect 576986 613898 577222 614134
rect 576986 578218 577222 578454
rect 576986 577898 577222 578134
rect 576986 542218 577222 542454
rect 576986 541898 577222 542134
rect 576986 506218 577222 506454
rect 576986 505898 577222 506134
rect 576986 470218 577222 470454
rect 576986 469898 577222 470134
rect 576986 434218 577222 434454
rect 576986 433898 577222 434134
rect 576986 398218 577222 398454
rect 576986 397898 577222 398134
rect 576986 362218 577222 362454
rect 576986 361898 577222 362134
rect 576986 326218 577222 326454
rect 576986 325898 577222 326134
rect 576986 290218 577222 290454
rect 576986 289898 577222 290134
rect 576986 254218 577222 254454
rect 576986 253898 577222 254134
rect 576986 218218 577222 218454
rect 576986 217898 577222 218134
rect 576986 182218 577222 182454
rect 576986 181898 577222 182134
rect 576986 146218 577222 146454
rect 576986 145898 577222 146134
rect 576986 110218 577222 110454
rect 576986 109898 577222 110134
rect 576986 74218 577222 74454
rect 576986 73898 577222 74134
rect 576986 38218 577222 38454
rect 576986 37898 577222 38134
rect 576986 2218 577222 2454
rect 576986 1898 577222 2134
rect 576986 -582 577222 -346
rect 576986 -902 577222 -666
rect 580586 617818 580822 618054
rect 580586 617498 580822 617734
rect 580586 581818 580822 582054
rect 580586 581498 580822 581734
rect 580586 545818 580822 546054
rect 580586 545498 580822 545734
rect 580586 509818 580822 510054
rect 580586 509498 580822 509734
rect 580586 473818 580822 474054
rect 580586 473498 580822 473734
rect 580586 437818 580822 438054
rect 580586 437498 580822 437734
rect 580586 401818 580822 402054
rect 580586 401498 580822 401734
rect 580586 365818 580822 366054
rect 580586 365498 580822 365734
rect 580586 329818 580822 330054
rect 580586 329498 580822 329734
rect 580586 293818 580822 294054
rect 580586 293498 580822 293734
rect 580586 257818 580822 258054
rect 580586 257498 580822 257734
rect 580586 221818 580822 222054
rect 580586 221498 580822 221734
rect 580586 185818 580822 186054
rect 580586 185498 580822 185734
rect 580586 149818 580822 150054
rect 580586 149498 580822 149734
rect 580586 113818 580822 114054
rect 580586 113498 580822 113734
rect 580586 77818 580822 78054
rect 580586 77498 580822 77734
rect 580586 41818 580822 42054
rect 580586 41498 580822 41734
rect 580586 5818 580822 6054
rect 580586 5498 580822 5734
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 686218 585738 686454
rect 585502 685898 585738 686134
rect 585502 650218 585738 650454
rect 585502 649898 585738 650134
rect 585502 614218 585738 614454
rect 585502 613898 585738 614134
rect 585502 578218 585738 578454
rect 585502 577898 585738 578134
rect 585502 542218 585738 542454
rect 585502 541898 585738 542134
rect 585502 506218 585738 506454
rect 585502 505898 585738 506134
rect 585502 470218 585738 470454
rect 585502 469898 585738 470134
rect 585502 434218 585738 434454
rect 585502 433898 585738 434134
rect 585502 398218 585738 398454
rect 585502 397898 585738 398134
rect 585502 362218 585738 362454
rect 585502 361898 585738 362134
rect 585502 326218 585738 326454
rect 585502 325898 585738 326134
rect 585502 290218 585738 290454
rect 585502 289898 585738 290134
rect 585502 254218 585738 254454
rect 585502 253898 585738 254134
rect 585502 218218 585738 218454
rect 585502 217898 585738 218134
rect 585502 182218 585738 182454
rect 585502 181898 585738 182134
rect 585502 146218 585738 146454
rect 585502 145898 585738 146134
rect 585502 110218 585738 110454
rect 585502 109898 585738 110134
rect 585502 74218 585738 74454
rect 585502 73898 585738 74134
rect 585502 38218 585738 38454
rect 585502 37898 585738 38134
rect 585502 2218 585738 2454
rect 585502 1898 585738 2134
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586442 668218 586678 668454
rect 586442 667898 586678 668134
rect 586442 632218 586678 632454
rect 586442 631898 586678 632134
rect 586442 596218 586678 596454
rect 586442 595898 586678 596134
rect 586442 560218 586678 560454
rect 586442 559898 586678 560134
rect 586442 524218 586678 524454
rect 586442 523898 586678 524134
rect 586442 488218 586678 488454
rect 586442 487898 586678 488134
rect 586442 452218 586678 452454
rect 586442 451898 586678 452134
rect 586442 416218 586678 416454
rect 586442 415898 586678 416134
rect 586442 380218 586678 380454
rect 586442 379898 586678 380134
rect 586442 344218 586678 344454
rect 586442 343898 586678 344134
rect 586442 308218 586678 308454
rect 586442 307898 586678 308134
rect 586442 272218 586678 272454
rect 586442 271898 586678 272134
rect 586442 236218 586678 236454
rect 586442 235898 586678 236134
rect 586442 200218 586678 200454
rect 586442 199898 586678 200134
rect 586442 164218 586678 164454
rect 586442 163898 586678 164134
rect 586442 128218 586678 128454
rect 586442 127898 586678 128134
rect 586442 92218 586678 92454
rect 586442 91898 586678 92134
rect 586442 56218 586678 56454
rect 586442 55898 586678 56134
rect 586442 20218 586678 20454
rect 586442 19898 586678 20134
rect 586442 -1522 586678 -1286
rect 586442 -1842 586678 -1606
rect 587382 689818 587618 690054
rect 587382 689498 587618 689734
rect 587382 653818 587618 654054
rect 587382 653498 587618 653734
rect 587382 617818 587618 618054
rect 587382 617498 587618 617734
rect 587382 581818 587618 582054
rect 587382 581498 587618 581734
rect 587382 545818 587618 546054
rect 587382 545498 587618 545734
rect 587382 509818 587618 510054
rect 587382 509498 587618 509734
rect 587382 473818 587618 474054
rect 587382 473498 587618 473734
rect 587382 437818 587618 438054
rect 587382 437498 587618 437734
rect 587382 401818 587618 402054
rect 587382 401498 587618 401734
rect 587382 365818 587618 366054
rect 587382 365498 587618 365734
rect 587382 329818 587618 330054
rect 587382 329498 587618 329734
rect 587382 293818 587618 294054
rect 587382 293498 587618 293734
rect 587382 257818 587618 258054
rect 587382 257498 587618 257734
rect 587382 221818 587618 222054
rect 587382 221498 587618 221734
rect 587382 185818 587618 186054
rect 587382 185498 587618 185734
rect 587382 149818 587618 150054
rect 587382 149498 587618 149734
rect 587382 113818 587618 114054
rect 587382 113498 587618 113734
rect 587382 77818 587618 78054
rect 587382 77498 587618 77734
rect 587382 41818 587618 42054
rect 587382 41498 587618 41734
rect 587382 5818 587618 6054
rect 587382 5498 587618 5734
rect 580586 -2462 580822 -2226
rect 580586 -2782 580822 -2546
rect 587382 -2462 587618 -2226
rect 587382 -2782 587618 -2546
rect 588322 671818 588558 672054
rect 588322 671498 588558 671734
rect 588322 635818 588558 636054
rect 588322 635498 588558 635734
rect 588322 599818 588558 600054
rect 588322 599498 588558 599734
rect 588322 563818 588558 564054
rect 588322 563498 588558 563734
rect 588322 527818 588558 528054
rect 588322 527498 588558 527734
rect 588322 491818 588558 492054
rect 588322 491498 588558 491734
rect 588322 455818 588558 456054
rect 588322 455498 588558 455734
rect 588322 419818 588558 420054
rect 588322 419498 588558 419734
rect 588322 383818 588558 384054
rect 588322 383498 588558 383734
rect 588322 347818 588558 348054
rect 588322 347498 588558 347734
rect 588322 311818 588558 312054
rect 588322 311498 588558 311734
rect 588322 275818 588558 276054
rect 588322 275498 588558 275734
rect 588322 239818 588558 240054
rect 588322 239498 588558 239734
rect 588322 203818 588558 204054
rect 588322 203498 588558 203734
rect 588322 167818 588558 168054
rect 588322 167498 588558 167734
rect 588322 131818 588558 132054
rect 588322 131498 588558 131734
rect 588322 95818 588558 96054
rect 588322 95498 588558 95734
rect 588322 59818 588558 60054
rect 588322 59498 588558 59734
rect 588322 23818 588558 24054
rect 588322 23498 588558 23734
rect 588322 -3402 588558 -3166
rect 588322 -3722 588558 -3486
rect 589262 693418 589498 693654
rect 589262 693098 589498 693334
rect 589262 657418 589498 657654
rect 589262 657098 589498 657334
rect 589262 621418 589498 621654
rect 589262 621098 589498 621334
rect 589262 585418 589498 585654
rect 589262 585098 589498 585334
rect 589262 549418 589498 549654
rect 589262 549098 589498 549334
rect 589262 513418 589498 513654
rect 589262 513098 589498 513334
rect 589262 477418 589498 477654
rect 589262 477098 589498 477334
rect 589262 441418 589498 441654
rect 589262 441098 589498 441334
rect 589262 405418 589498 405654
rect 589262 405098 589498 405334
rect 589262 369418 589498 369654
rect 589262 369098 589498 369334
rect 589262 333418 589498 333654
rect 589262 333098 589498 333334
rect 589262 297418 589498 297654
rect 589262 297098 589498 297334
rect 589262 261418 589498 261654
rect 589262 261098 589498 261334
rect 589262 225418 589498 225654
rect 589262 225098 589498 225334
rect 589262 189418 589498 189654
rect 589262 189098 589498 189334
rect 589262 153418 589498 153654
rect 589262 153098 589498 153334
rect 589262 117418 589498 117654
rect 589262 117098 589498 117334
rect 589262 81418 589498 81654
rect 589262 81098 589498 81334
rect 589262 45418 589498 45654
rect 589262 45098 589498 45334
rect 589262 9418 589498 9654
rect 589262 9098 589498 9334
rect 589262 -4342 589498 -4106
rect 589262 -4662 589498 -4426
rect 590202 675418 590438 675654
rect 590202 675098 590438 675334
rect 590202 639418 590438 639654
rect 590202 639098 590438 639334
rect 590202 603418 590438 603654
rect 590202 603098 590438 603334
rect 590202 567418 590438 567654
rect 590202 567098 590438 567334
rect 590202 531418 590438 531654
rect 590202 531098 590438 531334
rect 590202 495418 590438 495654
rect 590202 495098 590438 495334
rect 590202 459418 590438 459654
rect 590202 459098 590438 459334
rect 590202 423418 590438 423654
rect 590202 423098 590438 423334
rect 590202 387418 590438 387654
rect 590202 387098 590438 387334
rect 590202 351418 590438 351654
rect 590202 351098 590438 351334
rect 590202 315418 590438 315654
rect 590202 315098 590438 315334
rect 590202 279418 590438 279654
rect 590202 279098 590438 279334
rect 590202 243418 590438 243654
rect 590202 243098 590438 243334
rect 590202 207418 590438 207654
rect 590202 207098 590438 207334
rect 590202 171418 590438 171654
rect 590202 171098 590438 171334
rect 590202 135418 590438 135654
rect 590202 135098 590438 135334
rect 590202 99418 590438 99654
rect 590202 99098 590438 99334
rect 590202 63418 590438 63654
rect 590202 63098 590438 63334
rect 590202 27418 590438 27654
rect 590202 27098 590438 27334
rect 590202 -5282 590438 -5046
rect 590202 -5602 590438 -5366
rect 591142 697018 591378 697254
rect 591142 696698 591378 696934
rect 591142 661018 591378 661254
rect 591142 660698 591378 660934
rect 591142 625018 591378 625254
rect 591142 624698 591378 624934
rect 591142 589018 591378 589254
rect 591142 588698 591378 588934
rect 591142 553018 591378 553254
rect 591142 552698 591378 552934
rect 591142 517018 591378 517254
rect 591142 516698 591378 516934
rect 591142 481018 591378 481254
rect 591142 480698 591378 480934
rect 591142 445018 591378 445254
rect 591142 444698 591378 444934
rect 591142 409018 591378 409254
rect 591142 408698 591378 408934
rect 591142 373018 591378 373254
rect 591142 372698 591378 372934
rect 591142 337018 591378 337254
rect 591142 336698 591378 336934
rect 591142 301018 591378 301254
rect 591142 300698 591378 300934
rect 591142 265018 591378 265254
rect 591142 264698 591378 264934
rect 591142 229018 591378 229254
rect 591142 228698 591378 228934
rect 591142 193018 591378 193254
rect 591142 192698 591378 192934
rect 591142 157018 591378 157254
rect 591142 156698 591378 156934
rect 591142 121018 591378 121254
rect 591142 120698 591378 120934
rect 591142 85018 591378 85254
rect 591142 84698 591378 84934
rect 591142 49018 591378 49254
rect 591142 48698 591378 48934
rect 591142 13018 591378 13254
rect 591142 12698 591378 12934
rect 591142 -6222 591378 -5986
rect 591142 -6542 591378 -6306
rect 592082 679018 592318 679254
rect 592082 678698 592318 678934
rect 592082 643018 592318 643254
rect 592082 642698 592318 642934
rect 592082 607018 592318 607254
rect 592082 606698 592318 606934
rect 592082 571018 592318 571254
rect 592082 570698 592318 570934
rect 592082 535018 592318 535254
rect 592082 534698 592318 534934
rect 592082 499018 592318 499254
rect 592082 498698 592318 498934
rect 592082 463018 592318 463254
rect 592082 462698 592318 462934
rect 592082 427018 592318 427254
rect 592082 426698 592318 426934
rect 592082 391018 592318 391254
rect 592082 390698 592318 390934
rect 592082 355018 592318 355254
rect 592082 354698 592318 354934
rect 592082 319018 592318 319254
rect 592082 318698 592318 318934
rect 592082 283018 592318 283254
rect 592082 282698 592318 282934
rect 592082 247018 592318 247254
rect 592082 246698 592318 246934
rect 592082 211018 592318 211254
rect 592082 210698 592318 210934
rect 592082 175018 592318 175254
rect 592082 174698 592318 174934
rect 592082 139018 592318 139254
rect 592082 138698 592318 138934
rect 592082 103018 592318 103254
rect 592082 102698 592318 102934
rect 592082 67018 592318 67254
rect 592082 66698 592318 66934
rect 592082 31018 592318 31254
rect 592082 30698 592318 30934
rect 569786 -7162 570022 -6926
rect 569786 -7482 570022 -7246
rect 592082 -7162 592318 -6926
rect 592082 -7482 592318 -7246
<< metal5 >>
rect -8576 711440 -7976 711442
rect 29604 711440 30204 711442
rect 65604 711440 66204 711442
rect 101604 711440 102204 711442
rect 137604 711440 138204 711442
rect 173604 711440 174204 711442
rect 209604 711440 210204 711442
rect 245604 711440 246204 711442
rect 281604 711440 282204 711442
rect 317604 711440 318204 711442
rect 353604 711440 354204 711442
rect 389604 711440 390204 711442
rect 425604 711440 426204 711442
rect 461604 711440 462204 711442
rect 497604 711440 498204 711442
rect 533604 711440 534204 711442
rect 569604 711440 570204 711442
rect 591900 711440 592500 711442
rect -8576 711418 592500 711440
rect -8576 711182 -8394 711418
rect -8158 711182 29786 711418
rect 30022 711182 65786 711418
rect 66022 711182 101786 711418
rect 102022 711182 137786 711418
rect 138022 711182 173786 711418
rect 174022 711182 209786 711418
rect 210022 711182 245786 711418
rect 246022 711182 281786 711418
rect 282022 711182 317786 711418
rect 318022 711182 353786 711418
rect 354022 711182 389786 711418
rect 390022 711182 425786 711418
rect 426022 711182 461786 711418
rect 462022 711182 497786 711418
rect 498022 711182 533786 711418
rect 534022 711182 569786 711418
rect 570022 711182 592082 711418
rect 592318 711182 592500 711418
rect -8576 711098 592500 711182
rect -8576 710862 -8394 711098
rect -8158 710862 29786 711098
rect 30022 710862 65786 711098
rect 66022 710862 101786 711098
rect 102022 710862 137786 711098
rect 138022 710862 173786 711098
rect 174022 710862 209786 711098
rect 210022 710862 245786 711098
rect 246022 710862 281786 711098
rect 282022 710862 317786 711098
rect 318022 710862 353786 711098
rect 354022 710862 389786 711098
rect 390022 710862 425786 711098
rect 426022 710862 461786 711098
rect 462022 710862 497786 711098
rect 498022 710862 533786 711098
rect 534022 710862 569786 711098
rect 570022 710862 592082 711098
rect 592318 710862 592500 711098
rect -8576 710840 592500 710862
rect -8576 710838 -7976 710840
rect 29604 710838 30204 710840
rect 65604 710838 66204 710840
rect 101604 710838 102204 710840
rect 137604 710838 138204 710840
rect 173604 710838 174204 710840
rect 209604 710838 210204 710840
rect 245604 710838 246204 710840
rect 281604 710838 282204 710840
rect 317604 710838 318204 710840
rect 353604 710838 354204 710840
rect 389604 710838 390204 710840
rect 425604 710838 426204 710840
rect 461604 710838 462204 710840
rect 497604 710838 498204 710840
rect 533604 710838 534204 710840
rect 569604 710838 570204 710840
rect 591900 710838 592500 710840
rect -7636 710500 -7036 710502
rect 11604 710500 12204 710502
rect 47604 710500 48204 710502
rect 83604 710500 84204 710502
rect 119604 710500 120204 710502
rect 155604 710500 156204 710502
rect 191604 710500 192204 710502
rect 227604 710500 228204 710502
rect 263604 710500 264204 710502
rect 299604 710500 300204 710502
rect 335604 710500 336204 710502
rect 371604 710500 372204 710502
rect 407604 710500 408204 710502
rect 443604 710500 444204 710502
rect 479604 710500 480204 710502
rect 515604 710500 516204 710502
rect 551604 710500 552204 710502
rect 590960 710500 591560 710502
rect -7636 710478 591560 710500
rect -7636 710242 -7454 710478
rect -7218 710242 11786 710478
rect 12022 710242 47786 710478
rect 48022 710242 83786 710478
rect 84022 710242 119786 710478
rect 120022 710242 155786 710478
rect 156022 710242 191786 710478
rect 192022 710242 227786 710478
rect 228022 710242 263786 710478
rect 264022 710242 299786 710478
rect 300022 710242 335786 710478
rect 336022 710242 371786 710478
rect 372022 710242 407786 710478
rect 408022 710242 443786 710478
rect 444022 710242 479786 710478
rect 480022 710242 515786 710478
rect 516022 710242 551786 710478
rect 552022 710242 591142 710478
rect 591378 710242 591560 710478
rect -7636 710158 591560 710242
rect -7636 709922 -7454 710158
rect -7218 709922 11786 710158
rect 12022 709922 47786 710158
rect 48022 709922 83786 710158
rect 84022 709922 119786 710158
rect 120022 709922 155786 710158
rect 156022 709922 191786 710158
rect 192022 709922 227786 710158
rect 228022 709922 263786 710158
rect 264022 709922 299786 710158
rect 300022 709922 335786 710158
rect 336022 709922 371786 710158
rect 372022 709922 407786 710158
rect 408022 709922 443786 710158
rect 444022 709922 479786 710158
rect 480022 709922 515786 710158
rect 516022 709922 551786 710158
rect 552022 709922 591142 710158
rect 591378 709922 591560 710158
rect -7636 709900 591560 709922
rect -7636 709898 -7036 709900
rect 11604 709898 12204 709900
rect 47604 709898 48204 709900
rect 83604 709898 84204 709900
rect 119604 709898 120204 709900
rect 155604 709898 156204 709900
rect 191604 709898 192204 709900
rect 227604 709898 228204 709900
rect 263604 709898 264204 709900
rect 299604 709898 300204 709900
rect 335604 709898 336204 709900
rect 371604 709898 372204 709900
rect 407604 709898 408204 709900
rect 443604 709898 444204 709900
rect 479604 709898 480204 709900
rect 515604 709898 516204 709900
rect 551604 709898 552204 709900
rect 590960 709898 591560 709900
rect -6696 709560 -6096 709562
rect 26004 709560 26604 709562
rect 62004 709560 62604 709562
rect 98004 709560 98604 709562
rect 134004 709560 134604 709562
rect 170004 709560 170604 709562
rect 206004 709560 206604 709562
rect 242004 709560 242604 709562
rect 278004 709560 278604 709562
rect 314004 709560 314604 709562
rect 350004 709560 350604 709562
rect 386004 709560 386604 709562
rect 422004 709560 422604 709562
rect 458004 709560 458604 709562
rect 494004 709560 494604 709562
rect 530004 709560 530604 709562
rect 566004 709560 566604 709562
rect 590020 709560 590620 709562
rect -6696 709538 590620 709560
rect -6696 709302 -6514 709538
rect -6278 709302 26186 709538
rect 26422 709302 62186 709538
rect 62422 709302 98186 709538
rect 98422 709302 134186 709538
rect 134422 709302 170186 709538
rect 170422 709302 206186 709538
rect 206422 709302 242186 709538
rect 242422 709302 278186 709538
rect 278422 709302 314186 709538
rect 314422 709302 350186 709538
rect 350422 709302 386186 709538
rect 386422 709302 422186 709538
rect 422422 709302 458186 709538
rect 458422 709302 494186 709538
rect 494422 709302 530186 709538
rect 530422 709302 566186 709538
rect 566422 709302 590202 709538
rect 590438 709302 590620 709538
rect -6696 709218 590620 709302
rect -6696 708982 -6514 709218
rect -6278 708982 26186 709218
rect 26422 708982 62186 709218
rect 62422 708982 98186 709218
rect 98422 708982 134186 709218
rect 134422 708982 170186 709218
rect 170422 708982 206186 709218
rect 206422 708982 242186 709218
rect 242422 708982 278186 709218
rect 278422 708982 314186 709218
rect 314422 708982 350186 709218
rect 350422 708982 386186 709218
rect 386422 708982 422186 709218
rect 422422 708982 458186 709218
rect 458422 708982 494186 709218
rect 494422 708982 530186 709218
rect 530422 708982 566186 709218
rect 566422 708982 590202 709218
rect 590438 708982 590620 709218
rect -6696 708960 590620 708982
rect -6696 708958 -6096 708960
rect 26004 708958 26604 708960
rect 62004 708958 62604 708960
rect 98004 708958 98604 708960
rect 134004 708958 134604 708960
rect 170004 708958 170604 708960
rect 206004 708958 206604 708960
rect 242004 708958 242604 708960
rect 278004 708958 278604 708960
rect 314004 708958 314604 708960
rect 350004 708958 350604 708960
rect 386004 708958 386604 708960
rect 422004 708958 422604 708960
rect 458004 708958 458604 708960
rect 494004 708958 494604 708960
rect 530004 708958 530604 708960
rect 566004 708958 566604 708960
rect 590020 708958 590620 708960
rect -5756 708620 -5156 708622
rect 8004 708620 8604 708622
rect 44004 708620 44604 708622
rect 80004 708620 80604 708622
rect 116004 708620 116604 708622
rect 152004 708620 152604 708622
rect 188004 708620 188604 708622
rect 224004 708620 224604 708622
rect 260004 708620 260604 708622
rect 296004 708620 296604 708622
rect 332004 708620 332604 708622
rect 368004 708620 368604 708622
rect 404004 708620 404604 708622
rect 440004 708620 440604 708622
rect 476004 708620 476604 708622
rect 512004 708620 512604 708622
rect 548004 708620 548604 708622
rect 589080 708620 589680 708622
rect -5756 708598 589680 708620
rect -5756 708362 -5574 708598
rect -5338 708362 8186 708598
rect 8422 708362 44186 708598
rect 44422 708362 80186 708598
rect 80422 708362 116186 708598
rect 116422 708362 152186 708598
rect 152422 708362 188186 708598
rect 188422 708362 224186 708598
rect 224422 708362 260186 708598
rect 260422 708362 296186 708598
rect 296422 708362 332186 708598
rect 332422 708362 368186 708598
rect 368422 708362 404186 708598
rect 404422 708362 440186 708598
rect 440422 708362 476186 708598
rect 476422 708362 512186 708598
rect 512422 708362 548186 708598
rect 548422 708362 589262 708598
rect 589498 708362 589680 708598
rect -5756 708278 589680 708362
rect -5756 708042 -5574 708278
rect -5338 708042 8186 708278
rect 8422 708042 44186 708278
rect 44422 708042 80186 708278
rect 80422 708042 116186 708278
rect 116422 708042 152186 708278
rect 152422 708042 188186 708278
rect 188422 708042 224186 708278
rect 224422 708042 260186 708278
rect 260422 708042 296186 708278
rect 296422 708042 332186 708278
rect 332422 708042 368186 708278
rect 368422 708042 404186 708278
rect 404422 708042 440186 708278
rect 440422 708042 476186 708278
rect 476422 708042 512186 708278
rect 512422 708042 548186 708278
rect 548422 708042 589262 708278
rect 589498 708042 589680 708278
rect -5756 708020 589680 708042
rect -5756 708018 -5156 708020
rect 8004 708018 8604 708020
rect 44004 708018 44604 708020
rect 80004 708018 80604 708020
rect 116004 708018 116604 708020
rect 152004 708018 152604 708020
rect 188004 708018 188604 708020
rect 224004 708018 224604 708020
rect 260004 708018 260604 708020
rect 296004 708018 296604 708020
rect 332004 708018 332604 708020
rect 368004 708018 368604 708020
rect 404004 708018 404604 708020
rect 440004 708018 440604 708020
rect 476004 708018 476604 708020
rect 512004 708018 512604 708020
rect 548004 708018 548604 708020
rect 589080 708018 589680 708020
rect -4816 707680 -4216 707682
rect 22404 707680 23004 707682
rect 58404 707680 59004 707682
rect 94404 707680 95004 707682
rect 130404 707680 131004 707682
rect 166404 707680 167004 707682
rect 202404 707680 203004 707682
rect 238404 707680 239004 707682
rect 274404 707680 275004 707682
rect 310404 707680 311004 707682
rect 346404 707680 347004 707682
rect 382404 707680 383004 707682
rect 418404 707680 419004 707682
rect 454404 707680 455004 707682
rect 490404 707680 491004 707682
rect 526404 707680 527004 707682
rect 562404 707680 563004 707682
rect 588140 707680 588740 707682
rect -4816 707658 588740 707680
rect -4816 707422 -4634 707658
rect -4398 707422 22586 707658
rect 22822 707422 58586 707658
rect 58822 707422 94586 707658
rect 94822 707422 130586 707658
rect 130822 707422 166586 707658
rect 166822 707422 202586 707658
rect 202822 707422 238586 707658
rect 238822 707422 274586 707658
rect 274822 707422 310586 707658
rect 310822 707422 346586 707658
rect 346822 707422 382586 707658
rect 382822 707422 418586 707658
rect 418822 707422 454586 707658
rect 454822 707422 490586 707658
rect 490822 707422 526586 707658
rect 526822 707422 562586 707658
rect 562822 707422 588322 707658
rect 588558 707422 588740 707658
rect -4816 707338 588740 707422
rect -4816 707102 -4634 707338
rect -4398 707102 22586 707338
rect 22822 707102 58586 707338
rect 58822 707102 94586 707338
rect 94822 707102 130586 707338
rect 130822 707102 166586 707338
rect 166822 707102 202586 707338
rect 202822 707102 238586 707338
rect 238822 707102 274586 707338
rect 274822 707102 310586 707338
rect 310822 707102 346586 707338
rect 346822 707102 382586 707338
rect 382822 707102 418586 707338
rect 418822 707102 454586 707338
rect 454822 707102 490586 707338
rect 490822 707102 526586 707338
rect 526822 707102 562586 707338
rect 562822 707102 588322 707338
rect 588558 707102 588740 707338
rect -4816 707080 588740 707102
rect -4816 707078 -4216 707080
rect 22404 707078 23004 707080
rect 58404 707078 59004 707080
rect 94404 707078 95004 707080
rect 130404 707078 131004 707080
rect 166404 707078 167004 707080
rect 202404 707078 203004 707080
rect 238404 707078 239004 707080
rect 274404 707078 275004 707080
rect 310404 707078 311004 707080
rect 346404 707078 347004 707080
rect 382404 707078 383004 707080
rect 418404 707078 419004 707080
rect 454404 707078 455004 707080
rect 490404 707078 491004 707080
rect 526404 707078 527004 707080
rect 562404 707078 563004 707080
rect 588140 707078 588740 707080
rect -3876 706740 -3276 706742
rect 4404 706740 5004 706742
rect 40404 706740 41004 706742
rect 76404 706740 77004 706742
rect 112404 706740 113004 706742
rect 148404 706740 149004 706742
rect 184404 706740 185004 706742
rect 220404 706740 221004 706742
rect 256404 706740 257004 706742
rect 292404 706740 293004 706742
rect 328404 706740 329004 706742
rect 364404 706740 365004 706742
rect 400404 706740 401004 706742
rect 436404 706740 437004 706742
rect 472404 706740 473004 706742
rect 508404 706740 509004 706742
rect 544404 706740 545004 706742
rect 580404 706740 581004 706742
rect 587200 706740 587800 706742
rect -3876 706718 587800 706740
rect -3876 706482 -3694 706718
rect -3458 706482 4586 706718
rect 4822 706482 40586 706718
rect 40822 706482 76586 706718
rect 76822 706482 112586 706718
rect 112822 706482 148586 706718
rect 148822 706482 184586 706718
rect 184822 706482 220586 706718
rect 220822 706482 256586 706718
rect 256822 706482 292586 706718
rect 292822 706482 328586 706718
rect 328822 706482 364586 706718
rect 364822 706482 400586 706718
rect 400822 706482 436586 706718
rect 436822 706482 472586 706718
rect 472822 706482 508586 706718
rect 508822 706482 544586 706718
rect 544822 706482 580586 706718
rect 580822 706482 587382 706718
rect 587618 706482 587800 706718
rect -3876 706398 587800 706482
rect -3876 706162 -3694 706398
rect -3458 706162 4586 706398
rect 4822 706162 40586 706398
rect 40822 706162 76586 706398
rect 76822 706162 112586 706398
rect 112822 706162 148586 706398
rect 148822 706162 184586 706398
rect 184822 706162 220586 706398
rect 220822 706162 256586 706398
rect 256822 706162 292586 706398
rect 292822 706162 328586 706398
rect 328822 706162 364586 706398
rect 364822 706162 400586 706398
rect 400822 706162 436586 706398
rect 436822 706162 472586 706398
rect 472822 706162 508586 706398
rect 508822 706162 544586 706398
rect 544822 706162 580586 706398
rect 580822 706162 587382 706398
rect 587618 706162 587800 706398
rect -3876 706140 587800 706162
rect -3876 706138 -3276 706140
rect 4404 706138 5004 706140
rect 40404 706138 41004 706140
rect 76404 706138 77004 706140
rect 112404 706138 113004 706140
rect 148404 706138 149004 706140
rect 184404 706138 185004 706140
rect 220404 706138 221004 706140
rect 256404 706138 257004 706140
rect 292404 706138 293004 706140
rect 328404 706138 329004 706140
rect 364404 706138 365004 706140
rect 400404 706138 401004 706140
rect 436404 706138 437004 706140
rect 472404 706138 473004 706140
rect 508404 706138 509004 706140
rect 544404 706138 545004 706140
rect 580404 706138 581004 706140
rect 587200 706138 587800 706140
rect -2936 705800 -2336 705802
rect 18804 705800 19404 705802
rect 54804 705800 55404 705802
rect 90804 705800 91404 705802
rect 126804 705800 127404 705802
rect 162804 705800 163404 705802
rect 198804 705800 199404 705802
rect 234804 705800 235404 705802
rect 270804 705800 271404 705802
rect 306804 705800 307404 705802
rect 342804 705800 343404 705802
rect 378804 705800 379404 705802
rect 414804 705800 415404 705802
rect 450804 705800 451404 705802
rect 486804 705800 487404 705802
rect 522804 705800 523404 705802
rect 558804 705800 559404 705802
rect 586260 705800 586860 705802
rect -2936 705778 586860 705800
rect -2936 705542 -2754 705778
rect -2518 705542 18986 705778
rect 19222 705542 54986 705778
rect 55222 705542 90986 705778
rect 91222 705542 126986 705778
rect 127222 705542 162986 705778
rect 163222 705542 198986 705778
rect 199222 705542 234986 705778
rect 235222 705542 270986 705778
rect 271222 705542 306986 705778
rect 307222 705542 342986 705778
rect 343222 705542 378986 705778
rect 379222 705542 414986 705778
rect 415222 705542 450986 705778
rect 451222 705542 486986 705778
rect 487222 705542 522986 705778
rect 523222 705542 558986 705778
rect 559222 705542 586442 705778
rect 586678 705542 586860 705778
rect -2936 705458 586860 705542
rect -2936 705222 -2754 705458
rect -2518 705222 18986 705458
rect 19222 705222 54986 705458
rect 55222 705222 90986 705458
rect 91222 705222 126986 705458
rect 127222 705222 162986 705458
rect 163222 705222 198986 705458
rect 199222 705222 234986 705458
rect 235222 705222 270986 705458
rect 271222 705222 306986 705458
rect 307222 705222 342986 705458
rect 343222 705222 378986 705458
rect 379222 705222 414986 705458
rect 415222 705222 450986 705458
rect 451222 705222 486986 705458
rect 487222 705222 522986 705458
rect 523222 705222 558986 705458
rect 559222 705222 586442 705458
rect 586678 705222 586860 705458
rect -2936 705200 586860 705222
rect -2936 705198 -2336 705200
rect 18804 705198 19404 705200
rect 54804 705198 55404 705200
rect 90804 705198 91404 705200
rect 126804 705198 127404 705200
rect 162804 705198 163404 705200
rect 198804 705198 199404 705200
rect 234804 705198 235404 705200
rect 270804 705198 271404 705200
rect 306804 705198 307404 705200
rect 342804 705198 343404 705200
rect 378804 705198 379404 705200
rect 414804 705198 415404 705200
rect 450804 705198 451404 705200
rect 486804 705198 487404 705200
rect 522804 705198 523404 705200
rect 558804 705198 559404 705200
rect 586260 705198 586860 705200
rect -1996 704860 -1396 704862
rect 804 704860 1404 704862
rect 36804 704860 37404 704862
rect 72804 704860 73404 704862
rect 108804 704860 109404 704862
rect 144804 704860 145404 704862
rect 180804 704860 181404 704862
rect 216804 704860 217404 704862
rect 252804 704860 253404 704862
rect 288804 704860 289404 704862
rect 324804 704860 325404 704862
rect 360804 704860 361404 704862
rect 396804 704860 397404 704862
rect 432804 704860 433404 704862
rect 468804 704860 469404 704862
rect 504804 704860 505404 704862
rect 540804 704860 541404 704862
rect 576804 704860 577404 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 986 704838
rect 1222 704602 36986 704838
rect 37222 704602 72986 704838
rect 73222 704602 108986 704838
rect 109222 704602 144986 704838
rect 145222 704602 180986 704838
rect 181222 704602 216986 704838
rect 217222 704602 252986 704838
rect 253222 704602 288986 704838
rect 289222 704602 324986 704838
rect 325222 704602 360986 704838
rect 361222 704602 396986 704838
rect 397222 704602 432986 704838
rect 433222 704602 468986 704838
rect 469222 704602 504986 704838
rect 505222 704602 540986 704838
rect 541222 704602 576986 704838
rect 577222 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 986 704518
rect 1222 704282 36986 704518
rect 37222 704282 72986 704518
rect 73222 704282 108986 704518
rect 109222 704282 144986 704518
rect 145222 704282 180986 704518
rect 181222 704282 216986 704518
rect 217222 704282 252986 704518
rect 253222 704282 288986 704518
rect 289222 704282 324986 704518
rect 325222 704282 360986 704518
rect 361222 704282 396986 704518
rect 397222 704282 432986 704518
rect 433222 704282 468986 704518
rect 469222 704282 504986 704518
rect 505222 704282 540986 704518
rect 541222 704282 576986 704518
rect 577222 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 804 704258 1404 704260
rect 36804 704258 37404 704260
rect 72804 704258 73404 704260
rect 108804 704258 109404 704260
rect 144804 704258 145404 704260
rect 180804 704258 181404 704260
rect 216804 704258 217404 704260
rect 252804 704258 253404 704260
rect 288804 704258 289404 704260
rect 324804 704258 325404 704260
rect 360804 704258 361404 704260
rect 396804 704258 397404 704260
rect 432804 704258 433404 704260
rect 468804 704258 469404 704260
rect 504804 704258 505404 704260
rect 540804 704258 541404 704260
rect 576804 704258 577404 704260
rect 585320 704258 585920 704260
rect -7636 697276 -7036 697278
rect 11604 697276 12204 697278
rect 47604 697276 48204 697278
rect 83604 697276 84204 697278
rect 119604 697276 120204 697278
rect 155604 697276 156204 697278
rect 191604 697276 192204 697278
rect 227604 697276 228204 697278
rect 263604 697276 264204 697278
rect 299604 697276 300204 697278
rect 335604 697276 336204 697278
rect 371604 697276 372204 697278
rect 407604 697276 408204 697278
rect 443604 697276 444204 697278
rect 479604 697276 480204 697278
rect 515604 697276 516204 697278
rect 551604 697276 552204 697278
rect 590960 697276 591560 697278
rect -8576 697254 592500 697276
rect -8576 697018 -7454 697254
rect -7218 697018 11786 697254
rect 12022 697018 47786 697254
rect 48022 697018 83786 697254
rect 84022 697018 119786 697254
rect 120022 697018 155786 697254
rect 156022 697018 191786 697254
rect 192022 697018 227786 697254
rect 228022 697018 263786 697254
rect 264022 697018 299786 697254
rect 300022 697018 335786 697254
rect 336022 697018 371786 697254
rect 372022 697018 407786 697254
rect 408022 697018 443786 697254
rect 444022 697018 479786 697254
rect 480022 697018 515786 697254
rect 516022 697018 551786 697254
rect 552022 697018 591142 697254
rect 591378 697018 592500 697254
rect -8576 696934 592500 697018
rect -8576 696698 -7454 696934
rect -7218 696698 11786 696934
rect 12022 696698 47786 696934
rect 48022 696698 83786 696934
rect 84022 696698 119786 696934
rect 120022 696698 155786 696934
rect 156022 696698 191786 696934
rect 192022 696698 227786 696934
rect 228022 696698 263786 696934
rect 264022 696698 299786 696934
rect 300022 696698 335786 696934
rect 336022 696698 371786 696934
rect 372022 696698 407786 696934
rect 408022 696698 443786 696934
rect 444022 696698 479786 696934
rect 480022 696698 515786 696934
rect 516022 696698 551786 696934
rect 552022 696698 591142 696934
rect 591378 696698 592500 696934
rect -8576 696676 592500 696698
rect -7636 696674 -7036 696676
rect 11604 696674 12204 696676
rect 47604 696674 48204 696676
rect 83604 696674 84204 696676
rect 119604 696674 120204 696676
rect 155604 696674 156204 696676
rect 191604 696674 192204 696676
rect 227604 696674 228204 696676
rect 263604 696674 264204 696676
rect 299604 696674 300204 696676
rect 335604 696674 336204 696676
rect 371604 696674 372204 696676
rect 407604 696674 408204 696676
rect 443604 696674 444204 696676
rect 479604 696674 480204 696676
rect 515604 696674 516204 696676
rect 551604 696674 552204 696676
rect 590960 696674 591560 696676
rect -5756 693676 -5156 693678
rect 8004 693676 8604 693678
rect 44004 693676 44604 693678
rect 80004 693676 80604 693678
rect 116004 693676 116604 693678
rect 152004 693676 152604 693678
rect 188004 693676 188604 693678
rect 224004 693676 224604 693678
rect 260004 693676 260604 693678
rect 296004 693676 296604 693678
rect 332004 693676 332604 693678
rect 368004 693676 368604 693678
rect 404004 693676 404604 693678
rect 440004 693676 440604 693678
rect 476004 693676 476604 693678
rect 512004 693676 512604 693678
rect 548004 693676 548604 693678
rect 589080 693676 589680 693678
rect -6696 693654 590620 693676
rect -6696 693418 -5574 693654
rect -5338 693418 8186 693654
rect 8422 693418 44186 693654
rect 44422 693418 80186 693654
rect 80422 693418 116186 693654
rect 116422 693418 152186 693654
rect 152422 693418 188186 693654
rect 188422 693418 224186 693654
rect 224422 693418 260186 693654
rect 260422 693418 296186 693654
rect 296422 693418 332186 693654
rect 332422 693418 368186 693654
rect 368422 693418 404186 693654
rect 404422 693418 440186 693654
rect 440422 693418 476186 693654
rect 476422 693418 512186 693654
rect 512422 693418 548186 693654
rect 548422 693418 589262 693654
rect 589498 693418 590620 693654
rect -6696 693334 590620 693418
rect -6696 693098 -5574 693334
rect -5338 693098 8186 693334
rect 8422 693098 44186 693334
rect 44422 693098 80186 693334
rect 80422 693098 116186 693334
rect 116422 693098 152186 693334
rect 152422 693098 188186 693334
rect 188422 693098 224186 693334
rect 224422 693098 260186 693334
rect 260422 693098 296186 693334
rect 296422 693098 332186 693334
rect 332422 693098 368186 693334
rect 368422 693098 404186 693334
rect 404422 693098 440186 693334
rect 440422 693098 476186 693334
rect 476422 693098 512186 693334
rect 512422 693098 548186 693334
rect 548422 693098 589262 693334
rect 589498 693098 590620 693334
rect -6696 693076 590620 693098
rect -5756 693074 -5156 693076
rect 8004 693074 8604 693076
rect 44004 693074 44604 693076
rect 80004 693074 80604 693076
rect 116004 693074 116604 693076
rect 152004 693074 152604 693076
rect 188004 693074 188604 693076
rect 224004 693074 224604 693076
rect 260004 693074 260604 693076
rect 296004 693074 296604 693076
rect 332004 693074 332604 693076
rect 368004 693074 368604 693076
rect 404004 693074 404604 693076
rect 440004 693074 440604 693076
rect 476004 693074 476604 693076
rect 512004 693074 512604 693076
rect 548004 693074 548604 693076
rect 589080 693074 589680 693076
rect -3876 690076 -3276 690078
rect 4404 690076 5004 690078
rect 40404 690076 41004 690078
rect 76404 690076 77004 690078
rect 112404 690076 113004 690078
rect 148404 690076 149004 690078
rect 184404 690076 185004 690078
rect 220404 690076 221004 690078
rect 256404 690076 257004 690078
rect 292404 690076 293004 690078
rect 328404 690076 329004 690078
rect 364404 690076 365004 690078
rect 400404 690076 401004 690078
rect 436404 690076 437004 690078
rect 472404 690076 473004 690078
rect 508404 690076 509004 690078
rect 544404 690076 545004 690078
rect 580404 690076 581004 690078
rect 587200 690076 587800 690078
rect -4816 690054 588740 690076
rect -4816 689818 -3694 690054
rect -3458 689818 4586 690054
rect 4822 689818 40586 690054
rect 40822 689818 76586 690054
rect 76822 689818 112586 690054
rect 112822 689818 148586 690054
rect 148822 689818 184586 690054
rect 184822 689818 220586 690054
rect 220822 689818 256586 690054
rect 256822 689818 292586 690054
rect 292822 689818 328586 690054
rect 328822 689818 364586 690054
rect 364822 689818 400586 690054
rect 400822 689818 436586 690054
rect 436822 689818 472586 690054
rect 472822 689818 508586 690054
rect 508822 689818 544586 690054
rect 544822 689818 580586 690054
rect 580822 689818 587382 690054
rect 587618 689818 588740 690054
rect -4816 689734 588740 689818
rect -4816 689498 -3694 689734
rect -3458 689498 4586 689734
rect 4822 689498 40586 689734
rect 40822 689498 76586 689734
rect 76822 689498 112586 689734
rect 112822 689498 148586 689734
rect 148822 689498 184586 689734
rect 184822 689498 220586 689734
rect 220822 689498 256586 689734
rect 256822 689498 292586 689734
rect 292822 689498 328586 689734
rect 328822 689498 364586 689734
rect 364822 689498 400586 689734
rect 400822 689498 436586 689734
rect 436822 689498 472586 689734
rect 472822 689498 508586 689734
rect 508822 689498 544586 689734
rect 544822 689498 580586 689734
rect 580822 689498 587382 689734
rect 587618 689498 588740 689734
rect -4816 689476 588740 689498
rect -3876 689474 -3276 689476
rect 4404 689474 5004 689476
rect 40404 689474 41004 689476
rect 76404 689474 77004 689476
rect 112404 689474 113004 689476
rect 148404 689474 149004 689476
rect 184404 689474 185004 689476
rect 220404 689474 221004 689476
rect 256404 689474 257004 689476
rect 292404 689474 293004 689476
rect 328404 689474 329004 689476
rect 364404 689474 365004 689476
rect 400404 689474 401004 689476
rect 436404 689474 437004 689476
rect 472404 689474 473004 689476
rect 508404 689474 509004 689476
rect 544404 689474 545004 689476
rect 580404 689474 581004 689476
rect 587200 689474 587800 689476
rect -1996 686476 -1396 686478
rect 804 686476 1404 686478
rect 36804 686476 37404 686478
rect 72804 686476 73404 686478
rect 108804 686476 109404 686478
rect 144804 686476 145404 686478
rect 180804 686476 181404 686478
rect 216804 686476 217404 686478
rect 252804 686476 253404 686478
rect 288804 686476 289404 686478
rect 324804 686476 325404 686478
rect 360804 686476 361404 686478
rect 396804 686476 397404 686478
rect 432804 686476 433404 686478
rect 468804 686476 469404 686478
rect 504804 686476 505404 686478
rect 540804 686476 541404 686478
rect 576804 686476 577404 686478
rect 585320 686476 585920 686478
rect -2936 686454 586860 686476
rect -2936 686218 -1814 686454
rect -1578 686218 986 686454
rect 1222 686218 36986 686454
rect 37222 686218 72986 686454
rect 73222 686218 108986 686454
rect 109222 686218 144986 686454
rect 145222 686218 180986 686454
rect 181222 686218 216986 686454
rect 217222 686218 252986 686454
rect 253222 686218 288986 686454
rect 289222 686218 324986 686454
rect 325222 686218 360986 686454
rect 361222 686218 396986 686454
rect 397222 686218 432986 686454
rect 433222 686218 468986 686454
rect 469222 686218 504986 686454
rect 505222 686218 540986 686454
rect 541222 686218 576986 686454
rect 577222 686218 585502 686454
rect 585738 686218 586860 686454
rect -2936 686134 586860 686218
rect -2936 685898 -1814 686134
rect -1578 685898 986 686134
rect 1222 685898 36986 686134
rect 37222 685898 72986 686134
rect 73222 685898 108986 686134
rect 109222 685898 144986 686134
rect 145222 685898 180986 686134
rect 181222 685898 216986 686134
rect 217222 685898 252986 686134
rect 253222 685898 288986 686134
rect 289222 685898 324986 686134
rect 325222 685898 360986 686134
rect 361222 685898 396986 686134
rect 397222 685898 432986 686134
rect 433222 685898 468986 686134
rect 469222 685898 504986 686134
rect 505222 685898 540986 686134
rect 541222 685898 576986 686134
rect 577222 685898 585502 686134
rect 585738 685898 586860 686134
rect -2936 685876 586860 685898
rect -1996 685874 -1396 685876
rect 804 685874 1404 685876
rect 36804 685874 37404 685876
rect 72804 685874 73404 685876
rect 108804 685874 109404 685876
rect 144804 685874 145404 685876
rect 180804 685874 181404 685876
rect 216804 685874 217404 685876
rect 252804 685874 253404 685876
rect 288804 685874 289404 685876
rect 324804 685874 325404 685876
rect 360804 685874 361404 685876
rect 396804 685874 397404 685876
rect 432804 685874 433404 685876
rect 468804 685874 469404 685876
rect 504804 685874 505404 685876
rect 540804 685874 541404 685876
rect 576804 685874 577404 685876
rect 585320 685874 585920 685876
rect -8576 679276 -7976 679278
rect 29604 679276 30204 679278
rect 65604 679276 66204 679278
rect 101604 679276 102204 679278
rect 137604 679276 138204 679278
rect 173604 679276 174204 679278
rect 209604 679276 210204 679278
rect 245604 679276 246204 679278
rect 281604 679276 282204 679278
rect 317604 679276 318204 679278
rect 353604 679276 354204 679278
rect 389604 679276 390204 679278
rect 425604 679276 426204 679278
rect 461604 679276 462204 679278
rect 497604 679276 498204 679278
rect 533604 679276 534204 679278
rect 569604 679276 570204 679278
rect 591900 679276 592500 679278
rect -8576 679254 592500 679276
rect -8576 679018 -8394 679254
rect -8158 679018 29786 679254
rect 30022 679018 65786 679254
rect 66022 679018 101786 679254
rect 102022 679018 137786 679254
rect 138022 679018 173786 679254
rect 174022 679018 209786 679254
rect 210022 679018 245786 679254
rect 246022 679018 281786 679254
rect 282022 679018 317786 679254
rect 318022 679018 353786 679254
rect 354022 679018 389786 679254
rect 390022 679018 425786 679254
rect 426022 679018 461786 679254
rect 462022 679018 497786 679254
rect 498022 679018 533786 679254
rect 534022 679018 569786 679254
rect 570022 679018 592082 679254
rect 592318 679018 592500 679254
rect -8576 678934 592500 679018
rect -8576 678698 -8394 678934
rect -8158 678698 29786 678934
rect 30022 678698 65786 678934
rect 66022 678698 101786 678934
rect 102022 678698 137786 678934
rect 138022 678698 173786 678934
rect 174022 678698 209786 678934
rect 210022 678698 245786 678934
rect 246022 678698 281786 678934
rect 282022 678698 317786 678934
rect 318022 678698 353786 678934
rect 354022 678698 389786 678934
rect 390022 678698 425786 678934
rect 426022 678698 461786 678934
rect 462022 678698 497786 678934
rect 498022 678698 533786 678934
rect 534022 678698 569786 678934
rect 570022 678698 592082 678934
rect 592318 678698 592500 678934
rect -8576 678676 592500 678698
rect -8576 678674 -7976 678676
rect 29604 678674 30204 678676
rect 65604 678674 66204 678676
rect 101604 678674 102204 678676
rect 137604 678674 138204 678676
rect 173604 678674 174204 678676
rect 209604 678674 210204 678676
rect 245604 678674 246204 678676
rect 281604 678674 282204 678676
rect 317604 678674 318204 678676
rect 353604 678674 354204 678676
rect 389604 678674 390204 678676
rect 425604 678674 426204 678676
rect 461604 678674 462204 678676
rect 497604 678674 498204 678676
rect 533604 678674 534204 678676
rect 569604 678674 570204 678676
rect 591900 678674 592500 678676
rect -6696 675676 -6096 675678
rect 26004 675676 26604 675678
rect 62004 675676 62604 675678
rect 98004 675676 98604 675678
rect 134004 675676 134604 675678
rect 170004 675676 170604 675678
rect 206004 675676 206604 675678
rect 242004 675676 242604 675678
rect 278004 675676 278604 675678
rect 314004 675676 314604 675678
rect 350004 675676 350604 675678
rect 386004 675676 386604 675678
rect 422004 675676 422604 675678
rect 458004 675676 458604 675678
rect 494004 675676 494604 675678
rect 530004 675676 530604 675678
rect 566004 675676 566604 675678
rect 590020 675676 590620 675678
rect -6696 675654 590620 675676
rect -6696 675418 -6514 675654
rect -6278 675418 26186 675654
rect 26422 675418 62186 675654
rect 62422 675418 98186 675654
rect 98422 675418 134186 675654
rect 134422 675418 170186 675654
rect 170422 675418 206186 675654
rect 206422 675418 242186 675654
rect 242422 675418 278186 675654
rect 278422 675418 314186 675654
rect 314422 675418 350186 675654
rect 350422 675418 386186 675654
rect 386422 675418 422186 675654
rect 422422 675418 458186 675654
rect 458422 675418 494186 675654
rect 494422 675418 530186 675654
rect 530422 675418 566186 675654
rect 566422 675418 590202 675654
rect 590438 675418 590620 675654
rect -6696 675334 590620 675418
rect -6696 675098 -6514 675334
rect -6278 675098 26186 675334
rect 26422 675098 62186 675334
rect 62422 675098 98186 675334
rect 98422 675098 134186 675334
rect 134422 675098 170186 675334
rect 170422 675098 206186 675334
rect 206422 675098 242186 675334
rect 242422 675098 278186 675334
rect 278422 675098 314186 675334
rect 314422 675098 350186 675334
rect 350422 675098 386186 675334
rect 386422 675098 422186 675334
rect 422422 675098 458186 675334
rect 458422 675098 494186 675334
rect 494422 675098 530186 675334
rect 530422 675098 566186 675334
rect 566422 675098 590202 675334
rect 590438 675098 590620 675334
rect -6696 675076 590620 675098
rect -6696 675074 -6096 675076
rect 26004 675074 26604 675076
rect 62004 675074 62604 675076
rect 98004 675074 98604 675076
rect 134004 675074 134604 675076
rect 170004 675074 170604 675076
rect 206004 675074 206604 675076
rect 242004 675074 242604 675076
rect 278004 675074 278604 675076
rect 314004 675074 314604 675076
rect 350004 675074 350604 675076
rect 386004 675074 386604 675076
rect 422004 675074 422604 675076
rect 458004 675074 458604 675076
rect 494004 675074 494604 675076
rect 530004 675074 530604 675076
rect 566004 675074 566604 675076
rect 590020 675074 590620 675076
rect -4816 672076 -4216 672078
rect 22404 672076 23004 672078
rect 58404 672076 59004 672078
rect 94404 672076 95004 672078
rect 130404 672076 131004 672078
rect 166404 672076 167004 672078
rect 202404 672076 203004 672078
rect 238404 672076 239004 672078
rect 274404 672076 275004 672078
rect 310404 672076 311004 672078
rect 346404 672076 347004 672078
rect 382404 672076 383004 672078
rect 418404 672076 419004 672078
rect 454404 672076 455004 672078
rect 490404 672076 491004 672078
rect 526404 672076 527004 672078
rect 562404 672076 563004 672078
rect 588140 672076 588740 672078
rect -4816 672054 588740 672076
rect -4816 671818 -4634 672054
rect -4398 671818 22586 672054
rect 22822 671818 58586 672054
rect 58822 671818 94586 672054
rect 94822 671818 130586 672054
rect 130822 671818 166586 672054
rect 166822 671818 202586 672054
rect 202822 671818 238586 672054
rect 238822 671818 274586 672054
rect 274822 671818 310586 672054
rect 310822 671818 346586 672054
rect 346822 671818 382586 672054
rect 382822 671818 418586 672054
rect 418822 671818 454586 672054
rect 454822 671818 490586 672054
rect 490822 671818 526586 672054
rect 526822 671818 562586 672054
rect 562822 671818 588322 672054
rect 588558 671818 588740 672054
rect -4816 671734 588740 671818
rect -4816 671498 -4634 671734
rect -4398 671498 22586 671734
rect 22822 671498 58586 671734
rect 58822 671498 94586 671734
rect 94822 671498 130586 671734
rect 130822 671498 166586 671734
rect 166822 671498 202586 671734
rect 202822 671498 238586 671734
rect 238822 671498 274586 671734
rect 274822 671498 310586 671734
rect 310822 671498 346586 671734
rect 346822 671498 382586 671734
rect 382822 671498 418586 671734
rect 418822 671498 454586 671734
rect 454822 671498 490586 671734
rect 490822 671498 526586 671734
rect 526822 671498 562586 671734
rect 562822 671498 588322 671734
rect 588558 671498 588740 671734
rect -4816 671476 588740 671498
rect -4816 671474 -4216 671476
rect 22404 671474 23004 671476
rect 58404 671474 59004 671476
rect 94404 671474 95004 671476
rect 130404 671474 131004 671476
rect 166404 671474 167004 671476
rect 202404 671474 203004 671476
rect 238404 671474 239004 671476
rect 274404 671474 275004 671476
rect 310404 671474 311004 671476
rect 346404 671474 347004 671476
rect 382404 671474 383004 671476
rect 418404 671474 419004 671476
rect 454404 671474 455004 671476
rect 490404 671474 491004 671476
rect 526404 671474 527004 671476
rect 562404 671474 563004 671476
rect 588140 671474 588740 671476
rect -2936 668476 -2336 668478
rect 18804 668476 19404 668478
rect 54804 668476 55404 668478
rect 90804 668476 91404 668478
rect 126804 668476 127404 668478
rect 162804 668476 163404 668478
rect 198804 668476 199404 668478
rect 234804 668476 235404 668478
rect 270804 668476 271404 668478
rect 306804 668476 307404 668478
rect 342804 668476 343404 668478
rect 378804 668476 379404 668478
rect 414804 668476 415404 668478
rect 450804 668476 451404 668478
rect 486804 668476 487404 668478
rect 522804 668476 523404 668478
rect 558804 668476 559404 668478
rect 586260 668476 586860 668478
rect -2936 668454 586860 668476
rect -2936 668218 -2754 668454
rect -2518 668218 18986 668454
rect 19222 668218 54986 668454
rect 55222 668218 90986 668454
rect 91222 668218 126986 668454
rect 127222 668218 162986 668454
rect 163222 668218 198986 668454
rect 199222 668218 234986 668454
rect 235222 668218 270986 668454
rect 271222 668218 306986 668454
rect 307222 668218 342986 668454
rect 343222 668218 378986 668454
rect 379222 668218 414986 668454
rect 415222 668218 450986 668454
rect 451222 668218 486986 668454
rect 487222 668218 522986 668454
rect 523222 668218 558986 668454
rect 559222 668218 586442 668454
rect 586678 668218 586860 668454
rect -2936 668134 586860 668218
rect -2936 667898 -2754 668134
rect -2518 667898 18986 668134
rect 19222 667898 54986 668134
rect 55222 667898 90986 668134
rect 91222 667898 126986 668134
rect 127222 667898 162986 668134
rect 163222 667898 198986 668134
rect 199222 667898 234986 668134
rect 235222 667898 270986 668134
rect 271222 667898 306986 668134
rect 307222 667898 342986 668134
rect 343222 667898 378986 668134
rect 379222 667898 414986 668134
rect 415222 667898 450986 668134
rect 451222 667898 486986 668134
rect 487222 667898 522986 668134
rect 523222 667898 558986 668134
rect 559222 667898 586442 668134
rect 586678 667898 586860 668134
rect -2936 667876 586860 667898
rect -2936 667874 -2336 667876
rect 18804 667874 19404 667876
rect 54804 667874 55404 667876
rect 90804 667874 91404 667876
rect 126804 667874 127404 667876
rect 162804 667874 163404 667876
rect 198804 667874 199404 667876
rect 234804 667874 235404 667876
rect 270804 667874 271404 667876
rect 306804 667874 307404 667876
rect 342804 667874 343404 667876
rect 378804 667874 379404 667876
rect 414804 667874 415404 667876
rect 450804 667874 451404 667876
rect 486804 667874 487404 667876
rect 522804 667874 523404 667876
rect 558804 667874 559404 667876
rect 586260 667874 586860 667876
rect -7636 661276 -7036 661278
rect 11604 661276 12204 661278
rect 47604 661276 48204 661278
rect 83604 661276 84204 661278
rect 119604 661276 120204 661278
rect 155604 661276 156204 661278
rect 191604 661276 192204 661278
rect 227604 661276 228204 661278
rect 263604 661276 264204 661278
rect 299604 661276 300204 661278
rect 335604 661276 336204 661278
rect 371604 661276 372204 661278
rect 407604 661276 408204 661278
rect 443604 661276 444204 661278
rect 479604 661276 480204 661278
rect 515604 661276 516204 661278
rect 551604 661276 552204 661278
rect 590960 661276 591560 661278
rect -8576 661254 592500 661276
rect -8576 661018 -7454 661254
rect -7218 661018 11786 661254
rect 12022 661018 47786 661254
rect 48022 661018 83786 661254
rect 84022 661018 119786 661254
rect 120022 661018 155786 661254
rect 156022 661018 191786 661254
rect 192022 661018 227786 661254
rect 228022 661018 263786 661254
rect 264022 661018 299786 661254
rect 300022 661018 335786 661254
rect 336022 661018 371786 661254
rect 372022 661018 407786 661254
rect 408022 661018 443786 661254
rect 444022 661018 479786 661254
rect 480022 661018 515786 661254
rect 516022 661018 551786 661254
rect 552022 661018 591142 661254
rect 591378 661018 592500 661254
rect -8576 660934 592500 661018
rect -8576 660698 -7454 660934
rect -7218 660698 11786 660934
rect 12022 660698 47786 660934
rect 48022 660698 83786 660934
rect 84022 660698 119786 660934
rect 120022 660698 155786 660934
rect 156022 660698 191786 660934
rect 192022 660698 227786 660934
rect 228022 660698 263786 660934
rect 264022 660698 299786 660934
rect 300022 660698 335786 660934
rect 336022 660698 371786 660934
rect 372022 660698 407786 660934
rect 408022 660698 443786 660934
rect 444022 660698 479786 660934
rect 480022 660698 515786 660934
rect 516022 660698 551786 660934
rect 552022 660698 591142 660934
rect 591378 660698 592500 660934
rect -8576 660676 592500 660698
rect -7636 660674 -7036 660676
rect 11604 660674 12204 660676
rect 47604 660674 48204 660676
rect 83604 660674 84204 660676
rect 119604 660674 120204 660676
rect 155604 660674 156204 660676
rect 191604 660674 192204 660676
rect 227604 660674 228204 660676
rect 263604 660674 264204 660676
rect 299604 660674 300204 660676
rect 335604 660674 336204 660676
rect 371604 660674 372204 660676
rect 407604 660674 408204 660676
rect 443604 660674 444204 660676
rect 479604 660674 480204 660676
rect 515604 660674 516204 660676
rect 551604 660674 552204 660676
rect 590960 660674 591560 660676
rect -5756 657676 -5156 657678
rect 8004 657676 8604 657678
rect 44004 657676 44604 657678
rect 80004 657676 80604 657678
rect 116004 657676 116604 657678
rect 152004 657676 152604 657678
rect 188004 657676 188604 657678
rect 224004 657676 224604 657678
rect 260004 657676 260604 657678
rect 296004 657676 296604 657678
rect 332004 657676 332604 657678
rect 368004 657676 368604 657678
rect 404004 657676 404604 657678
rect 440004 657676 440604 657678
rect 476004 657676 476604 657678
rect 512004 657676 512604 657678
rect 548004 657676 548604 657678
rect 589080 657676 589680 657678
rect -6696 657654 590620 657676
rect -6696 657418 -5574 657654
rect -5338 657418 8186 657654
rect 8422 657418 44186 657654
rect 44422 657418 80186 657654
rect 80422 657418 116186 657654
rect 116422 657418 152186 657654
rect 152422 657418 188186 657654
rect 188422 657418 224186 657654
rect 224422 657418 260186 657654
rect 260422 657418 296186 657654
rect 296422 657418 332186 657654
rect 332422 657418 368186 657654
rect 368422 657418 404186 657654
rect 404422 657418 440186 657654
rect 440422 657418 476186 657654
rect 476422 657418 512186 657654
rect 512422 657418 548186 657654
rect 548422 657418 589262 657654
rect 589498 657418 590620 657654
rect -6696 657334 590620 657418
rect -6696 657098 -5574 657334
rect -5338 657098 8186 657334
rect 8422 657098 44186 657334
rect 44422 657098 80186 657334
rect 80422 657098 116186 657334
rect 116422 657098 152186 657334
rect 152422 657098 188186 657334
rect 188422 657098 224186 657334
rect 224422 657098 260186 657334
rect 260422 657098 296186 657334
rect 296422 657098 332186 657334
rect 332422 657098 368186 657334
rect 368422 657098 404186 657334
rect 404422 657098 440186 657334
rect 440422 657098 476186 657334
rect 476422 657098 512186 657334
rect 512422 657098 548186 657334
rect 548422 657098 589262 657334
rect 589498 657098 590620 657334
rect -6696 657076 590620 657098
rect -5756 657074 -5156 657076
rect 8004 657074 8604 657076
rect 44004 657074 44604 657076
rect 80004 657074 80604 657076
rect 116004 657074 116604 657076
rect 152004 657074 152604 657076
rect 188004 657074 188604 657076
rect 224004 657074 224604 657076
rect 260004 657074 260604 657076
rect 296004 657074 296604 657076
rect 332004 657074 332604 657076
rect 368004 657074 368604 657076
rect 404004 657074 404604 657076
rect 440004 657074 440604 657076
rect 476004 657074 476604 657076
rect 512004 657074 512604 657076
rect 548004 657074 548604 657076
rect 589080 657074 589680 657076
rect -3876 654076 -3276 654078
rect 4404 654076 5004 654078
rect 40404 654076 41004 654078
rect 148404 654076 149004 654078
rect 184404 654076 185004 654078
rect 292404 654076 293004 654078
rect 400404 654076 401004 654078
rect 436404 654076 437004 654078
rect 472404 654076 473004 654078
rect 508404 654076 509004 654078
rect 544404 654076 545004 654078
rect 580404 654076 581004 654078
rect 587200 654076 587800 654078
rect -4816 654054 588740 654076
rect -4816 653818 -3694 654054
rect -3458 653818 4586 654054
rect 4822 653818 40586 654054
rect 40822 653818 148586 654054
rect 148822 653818 184586 654054
rect 184822 653818 292586 654054
rect 292822 653818 400586 654054
rect 400822 653818 436586 654054
rect 436822 653818 472586 654054
rect 472822 653818 508586 654054
rect 508822 653818 544586 654054
rect 544822 653818 580586 654054
rect 580822 653818 587382 654054
rect 587618 653818 588740 654054
rect -4816 653734 588740 653818
rect -4816 653498 -3694 653734
rect -3458 653498 4586 653734
rect 4822 653498 40586 653734
rect 40822 653498 148586 653734
rect 148822 653498 184586 653734
rect 184822 653498 292586 653734
rect 292822 653498 400586 653734
rect 400822 653498 436586 653734
rect 436822 653498 472586 653734
rect 472822 653498 508586 653734
rect 508822 653498 544586 653734
rect 544822 653498 580586 653734
rect 580822 653498 587382 653734
rect 587618 653498 588740 653734
rect -4816 653476 588740 653498
rect -3876 653474 -3276 653476
rect 4404 653474 5004 653476
rect 40404 653474 41004 653476
rect 148404 653474 149004 653476
rect 184404 653474 185004 653476
rect 292404 653474 293004 653476
rect 400404 653474 401004 653476
rect 436404 653474 437004 653476
rect 472404 653474 473004 653476
rect 508404 653474 509004 653476
rect 544404 653474 545004 653476
rect 580404 653474 581004 653476
rect 587200 653474 587800 653476
rect -1996 650476 -1396 650478
rect 804 650476 1404 650478
rect 36804 650476 37404 650478
rect 144804 650476 145404 650478
rect 180804 650476 181404 650478
rect 288804 650476 289404 650478
rect 396804 650476 397404 650478
rect 432804 650476 433404 650478
rect 468804 650476 469404 650478
rect 504804 650476 505404 650478
rect 540804 650476 541404 650478
rect 576804 650476 577404 650478
rect 585320 650476 585920 650478
rect -2936 650454 586860 650476
rect -2936 650218 -1814 650454
rect -1578 650218 986 650454
rect 1222 650218 36986 650454
rect 37222 650218 144986 650454
rect 145222 650218 180986 650454
rect 181222 650218 288986 650454
rect 289222 650218 396986 650454
rect 397222 650218 432986 650454
rect 433222 650218 468986 650454
rect 469222 650218 504986 650454
rect 505222 650218 540986 650454
rect 541222 650218 576986 650454
rect 577222 650218 585502 650454
rect 585738 650218 586860 650454
rect -2936 650134 586860 650218
rect -2936 649898 -1814 650134
rect -1578 649898 986 650134
rect 1222 649898 36986 650134
rect 37222 649898 144986 650134
rect 145222 649898 180986 650134
rect 181222 649898 288986 650134
rect 289222 649898 396986 650134
rect 397222 649898 432986 650134
rect 433222 649898 468986 650134
rect 469222 649898 504986 650134
rect 505222 649898 540986 650134
rect 541222 649898 576986 650134
rect 577222 649898 585502 650134
rect 585738 649898 586860 650134
rect -2936 649876 586860 649898
rect -1996 649874 -1396 649876
rect 804 649874 1404 649876
rect 36804 649874 37404 649876
rect 144804 649874 145404 649876
rect 180804 649874 181404 649876
rect 288804 649874 289404 649876
rect 396804 649874 397404 649876
rect 432804 649874 433404 649876
rect 468804 649874 469404 649876
rect 504804 649874 505404 649876
rect 540804 649874 541404 649876
rect 576804 649874 577404 649876
rect 585320 649874 585920 649876
rect -8576 643276 -7976 643278
rect 29604 643276 30204 643278
rect 136938 643276 137262 643278
rect 173604 643276 174204 643278
rect 266938 643276 267262 643278
rect 281604 643276 282204 643278
rect 386938 643276 387262 643278
rect 425604 643276 426204 643278
rect 461604 643276 462204 643278
rect 497604 643276 498204 643278
rect 533604 643276 534204 643278
rect 569604 643276 570204 643278
rect 591900 643276 592500 643278
rect -8576 643254 592500 643276
rect -8576 643018 -8394 643254
rect -8158 643018 29786 643254
rect 30022 643018 136982 643254
rect 137218 643018 173786 643254
rect 174022 643018 266982 643254
rect 267218 643018 281786 643254
rect 282022 643018 386982 643254
rect 387218 643018 425786 643254
rect 426022 643018 461786 643254
rect 462022 643018 497786 643254
rect 498022 643018 533786 643254
rect 534022 643018 569786 643254
rect 570022 643018 592082 643254
rect 592318 643018 592500 643254
rect -8576 642934 592500 643018
rect -8576 642698 -8394 642934
rect -8158 642698 29786 642934
rect 30022 642698 136982 642934
rect 137218 642698 173786 642934
rect 174022 642698 266982 642934
rect 267218 642698 281786 642934
rect 282022 642698 386982 642934
rect 387218 642698 425786 642934
rect 426022 642698 461786 642934
rect 462022 642698 497786 642934
rect 498022 642698 533786 642934
rect 534022 642698 569786 642934
rect 570022 642698 592082 642934
rect 592318 642698 592500 642934
rect -8576 642676 592500 642698
rect -8576 642674 -7976 642676
rect 29604 642674 30204 642676
rect 136938 642674 137262 642676
rect 173604 642674 174204 642676
rect 266938 642674 267262 642676
rect 281604 642674 282204 642676
rect 386938 642674 387262 642676
rect 425604 642674 426204 642676
rect 461604 642674 462204 642676
rect 497604 642674 498204 642676
rect 533604 642674 534204 642676
rect 569604 642674 570204 642676
rect 591900 642674 592500 642676
rect -6696 639676 -6096 639678
rect 26004 639676 26604 639678
rect 136938 639676 137262 639678
rect 170004 639676 170604 639678
rect 266938 639676 267262 639678
rect 278004 639676 278604 639678
rect 386938 639676 387262 639678
rect 422004 639676 422604 639678
rect 458004 639676 458604 639678
rect 494004 639676 494604 639678
rect 530004 639676 530604 639678
rect 566004 639676 566604 639678
rect 590020 639676 590620 639678
rect -6696 639654 590620 639676
rect -6696 639418 -6514 639654
rect -6278 639418 26186 639654
rect 26422 639418 136982 639654
rect 137218 639418 170186 639654
rect 170422 639418 266982 639654
rect 267218 639418 278186 639654
rect 278422 639418 386982 639654
rect 387218 639418 422186 639654
rect 422422 639418 458186 639654
rect 458422 639418 494186 639654
rect 494422 639418 530186 639654
rect 530422 639418 566186 639654
rect 566422 639418 590202 639654
rect 590438 639418 590620 639654
rect -6696 639334 590620 639418
rect -6696 639098 -6514 639334
rect -6278 639098 26186 639334
rect 26422 639098 136982 639334
rect 137218 639098 170186 639334
rect 170422 639098 266982 639334
rect 267218 639098 278186 639334
rect 278422 639098 386982 639334
rect 387218 639098 422186 639334
rect 422422 639098 458186 639334
rect 458422 639098 494186 639334
rect 494422 639098 530186 639334
rect 530422 639098 566186 639334
rect 566422 639098 590202 639334
rect 590438 639098 590620 639334
rect -6696 639076 590620 639098
rect -6696 639074 -6096 639076
rect 26004 639074 26604 639076
rect 136938 639074 137262 639076
rect 170004 639074 170604 639076
rect 266938 639074 267262 639076
rect 278004 639074 278604 639076
rect 386938 639074 387262 639076
rect 422004 639074 422604 639076
rect 458004 639074 458604 639076
rect 494004 639074 494604 639076
rect 530004 639074 530604 639076
rect 566004 639074 566604 639076
rect 590020 639074 590620 639076
rect -4816 636076 -4216 636078
rect 22404 636076 23004 636078
rect 136938 636076 137262 636078
rect 166404 636076 167004 636078
rect 266938 636076 267262 636078
rect 274404 636076 275004 636078
rect 386938 636076 387262 636078
rect 418404 636076 419004 636078
rect 454404 636076 455004 636078
rect 490404 636076 491004 636078
rect 526404 636076 527004 636078
rect 562404 636076 563004 636078
rect 588140 636076 588740 636078
rect -4816 636054 588740 636076
rect -4816 635818 -4634 636054
rect -4398 635818 22586 636054
rect 22822 635818 136982 636054
rect 137218 635818 166586 636054
rect 166822 635818 266982 636054
rect 267218 635818 274586 636054
rect 274822 635818 386982 636054
rect 387218 635818 418586 636054
rect 418822 635818 454586 636054
rect 454822 635818 490586 636054
rect 490822 635818 526586 636054
rect 526822 635818 562586 636054
rect 562822 635818 588322 636054
rect 588558 635818 588740 636054
rect -4816 635734 588740 635818
rect -4816 635498 -4634 635734
rect -4398 635498 22586 635734
rect 22822 635498 136982 635734
rect 137218 635498 166586 635734
rect 166822 635498 266982 635734
rect 267218 635498 274586 635734
rect 274822 635498 386982 635734
rect 387218 635498 418586 635734
rect 418822 635498 454586 635734
rect 454822 635498 490586 635734
rect 490822 635498 526586 635734
rect 526822 635498 562586 635734
rect 562822 635498 588322 635734
rect 588558 635498 588740 635734
rect -4816 635476 588740 635498
rect -4816 635474 -4216 635476
rect 22404 635474 23004 635476
rect 136938 635474 137262 635476
rect 166404 635474 167004 635476
rect 266938 635474 267262 635476
rect 274404 635474 275004 635476
rect 386938 635474 387262 635476
rect 418404 635474 419004 635476
rect 454404 635474 455004 635476
rect 490404 635474 491004 635476
rect 526404 635474 527004 635476
rect 562404 635474 563004 635476
rect 588140 635474 588740 635476
rect -2936 632476 -2336 632478
rect 18804 632476 19404 632478
rect 54804 632476 55404 632478
rect 136938 632476 137262 632478
rect 162804 632476 163404 632478
rect 266938 632476 267262 632478
rect 270804 632476 271404 632478
rect 386938 632476 387262 632478
rect 414804 632476 415404 632478
rect 450804 632476 451404 632478
rect 486804 632476 487404 632478
rect 522804 632476 523404 632478
rect 558804 632476 559404 632478
rect 586260 632476 586860 632478
rect -2936 632454 586860 632476
rect -2936 632218 -2754 632454
rect -2518 632218 18986 632454
rect 19222 632218 54986 632454
rect 55222 632218 136982 632454
rect 137218 632218 162986 632454
rect 163222 632218 266982 632454
rect 267218 632218 270986 632454
rect 271222 632218 386982 632454
rect 387218 632218 414986 632454
rect 415222 632218 450986 632454
rect 451222 632218 486986 632454
rect 487222 632218 522986 632454
rect 523222 632218 558986 632454
rect 559222 632218 586442 632454
rect 586678 632218 586860 632454
rect -2936 632134 586860 632218
rect -2936 631898 -2754 632134
rect -2518 631898 18986 632134
rect 19222 631898 54986 632134
rect 55222 631898 136982 632134
rect 137218 631898 162986 632134
rect 163222 631898 266982 632134
rect 267218 631898 270986 632134
rect 271222 631898 386982 632134
rect 387218 631898 414986 632134
rect 415222 631898 450986 632134
rect 451222 631898 486986 632134
rect 487222 631898 522986 632134
rect 523222 631898 558986 632134
rect 559222 631898 586442 632134
rect 586678 631898 586860 632134
rect -2936 631876 586860 631898
rect -2936 631874 -2336 631876
rect 18804 631874 19404 631876
rect 54804 631874 55404 631876
rect 136938 631874 137262 631876
rect 162804 631874 163404 631876
rect 266938 631874 267262 631876
rect 270804 631874 271404 631876
rect 386938 631874 387262 631876
rect 414804 631874 415404 631876
rect 450804 631874 451404 631876
rect 486804 631874 487404 631876
rect 522804 631874 523404 631876
rect 558804 631874 559404 631876
rect 586260 631874 586860 631876
rect -7636 625276 -7036 625278
rect 11604 625276 12204 625278
rect 47604 625276 48204 625278
rect 136494 625276 136814 625278
rect 155604 625276 156204 625278
rect 266494 625276 266814 625278
rect 299604 625276 300204 625278
rect 386494 625276 386814 625278
rect 407604 625276 408204 625278
rect 443604 625276 444204 625278
rect 479604 625276 480204 625278
rect 515604 625276 516204 625278
rect 551604 625276 552204 625278
rect 590960 625276 591560 625278
rect -8576 625254 592500 625276
rect -8576 625018 -7454 625254
rect -7218 625018 11786 625254
rect 12022 625018 47786 625254
rect 48022 625018 136536 625254
rect 136772 625018 155786 625254
rect 156022 625018 266536 625254
rect 266772 625018 299786 625254
rect 300022 625018 386536 625254
rect 386772 625018 407786 625254
rect 408022 625018 443786 625254
rect 444022 625018 479786 625254
rect 480022 625018 515786 625254
rect 516022 625018 551786 625254
rect 552022 625018 591142 625254
rect 591378 625018 592500 625254
rect -8576 624934 592500 625018
rect -8576 624698 -7454 624934
rect -7218 624698 11786 624934
rect 12022 624698 47786 624934
rect 48022 624698 136536 624934
rect 136772 624698 155786 624934
rect 156022 624698 266536 624934
rect 266772 624698 299786 624934
rect 300022 624698 386536 624934
rect 386772 624698 407786 624934
rect 408022 624698 443786 624934
rect 444022 624698 479786 624934
rect 480022 624698 515786 624934
rect 516022 624698 551786 624934
rect 552022 624698 591142 624934
rect 591378 624698 592500 624934
rect -8576 624676 592500 624698
rect -7636 624674 -7036 624676
rect 11604 624674 12204 624676
rect 47604 624674 48204 624676
rect 136494 624674 136814 624676
rect 155604 624674 156204 624676
rect 266494 624674 266814 624676
rect 299604 624674 300204 624676
rect 386494 624674 386814 624676
rect 407604 624674 408204 624676
rect 443604 624674 444204 624676
rect 479604 624674 480204 624676
rect 515604 624674 516204 624676
rect 551604 624674 552204 624676
rect 590960 624674 591560 624676
rect -5756 621676 -5156 621678
rect 8004 621676 8604 621678
rect 44004 621676 44604 621678
rect 136494 621676 136814 621678
rect 152004 621676 152604 621678
rect 266494 621676 266814 621678
rect 296004 621676 296604 621678
rect 386494 621676 386814 621678
rect 404004 621676 404604 621678
rect 440004 621676 440604 621678
rect 476004 621676 476604 621678
rect 512004 621676 512604 621678
rect 548004 621676 548604 621678
rect 589080 621676 589680 621678
rect -6696 621654 590620 621676
rect -6696 621418 -5574 621654
rect -5338 621418 8186 621654
rect 8422 621418 44186 621654
rect 44422 621418 136536 621654
rect 136772 621418 152186 621654
rect 152422 621418 266536 621654
rect 266772 621418 296186 621654
rect 296422 621418 386536 621654
rect 386772 621418 404186 621654
rect 404422 621418 440186 621654
rect 440422 621418 476186 621654
rect 476422 621418 512186 621654
rect 512422 621418 548186 621654
rect 548422 621418 589262 621654
rect 589498 621418 590620 621654
rect -6696 621334 590620 621418
rect -6696 621098 -5574 621334
rect -5338 621098 8186 621334
rect 8422 621098 44186 621334
rect 44422 621098 136536 621334
rect 136772 621098 152186 621334
rect 152422 621098 266536 621334
rect 266772 621098 296186 621334
rect 296422 621098 386536 621334
rect 386772 621098 404186 621334
rect 404422 621098 440186 621334
rect 440422 621098 476186 621334
rect 476422 621098 512186 621334
rect 512422 621098 548186 621334
rect 548422 621098 589262 621334
rect 589498 621098 590620 621334
rect -6696 621076 590620 621098
rect -5756 621074 -5156 621076
rect 8004 621074 8604 621076
rect 44004 621074 44604 621076
rect 136494 621074 136814 621076
rect 152004 621074 152604 621076
rect 266494 621074 266814 621076
rect 296004 621074 296604 621076
rect 386494 621074 386814 621076
rect 404004 621074 404604 621076
rect 440004 621074 440604 621076
rect 476004 621074 476604 621076
rect 512004 621074 512604 621076
rect 548004 621074 548604 621076
rect 589080 621074 589680 621076
rect -3876 618076 -3276 618078
rect 4404 618076 5004 618078
rect 40404 618076 41004 618078
rect 136494 618076 136814 618078
rect 148404 618076 149004 618078
rect 184404 618076 185004 618078
rect 266494 618076 266814 618078
rect 292404 618076 293004 618078
rect 386494 618076 386814 618078
rect 400404 618076 401004 618078
rect 436404 618076 437004 618078
rect 472404 618076 473004 618078
rect 508404 618076 509004 618078
rect 544404 618076 545004 618078
rect 580404 618076 581004 618078
rect 587200 618076 587800 618078
rect -4816 618054 588740 618076
rect -4816 617818 -3694 618054
rect -3458 617818 4586 618054
rect 4822 617818 40586 618054
rect 40822 617818 136536 618054
rect 136772 617818 148586 618054
rect 148822 617818 184586 618054
rect 184822 617818 266536 618054
rect 266772 617818 292586 618054
rect 292822 617818 386536 618054
rect 386772 617818 400586 618054
rect 400822 617818 436586 618054
rect 436822 617818 472586 618054
rect 472822 617818 508586 618054
rect 508822 617818 544586 618054
rect 544822 617818 580586 618054
rect 580822 617818 587382 618054
rect 587618 617818 588740 618054
rect -4816 617734 588740 617818
rect -4816 617498 -3694 617734
rect -3458 617498 4586 617734
rect 4822 617498 40586 617734
rect 40822 617498 136536 617734
rect 136772 617498 148586 617734
rect 148822 617498 184586 617734
rect 184822 617498 266536 617734
rect 266772 617498 292586 617734
rect 292822 617498 386536 617734
rect 386772 617498 400586 617734
rect 400822 617498 436586 617734
rect 436822 617498 472586 617734
rect 472822 617498 508586 617734
rect 508822 617498 544586 617734
rect 544822 617498 580586 617734
rect 580822 617498 587382 617734
rect 587618 617498 588740 617734
rect -4816 617476 588740 617498
rect -3876 617474 -3276 617476
rect 4404 617474 5004 617476
rect 40404 617474 41004 617476
rect 136494 617474 136814 617476
rect 148404 617474 149004 617476
rect 184404 617474 185004 617476
rect 266494 617474 266814 617476
rect 292404 617474 293004 617476
rect 386494 617474 386814 617476
rect 400404 617474 401004 617476
rect 436404 617474 437004 617476
rect 472404 617474 473004 617476
rect 508404 617474 509004 617476
rect 544404 617474 545004 617476
rect 580404 617474 581004 617476
rect 587200 617474 587800 617476
rect -1996 614476 -1396 614478
rect 804 614476 1404 614478
rect 36804 614476 37404 614478
rect 136494 614476 136814 614478
rect 144804 614476 145404 614478
rect 180804 614476 181404 614478
rect 266494 614476 266814 614478
rect 288804 614476 289404 614478
rect 386494 614476 386814 614478
rect 396804 614476 397404 614478
rect 432804 614476 433404 614478
rect 468804 614476 469404 614478
rect 504804 614476 505404 614478
rect 540804 614476 541404 614478
rect 576804 614476 577404 614478
rect 585320 614476 585920 614478
rect -2936 614454 586860 614476
rect -2936 614218 -1814 614454
rect -1578 614218 986 614454
rect 1222 614218 36986 614454
rect 37222 614218 136536 614454
rect 136772 614218 144986 614454
rect 145222 614218 180986 614454
rect 181222 614218 266536 614454
rect 266772 614218 288986 614454
rect 289222 614218 386536 614454
rect 386772 614218 396986 614454
rect 397222 614218 432986 614454
rect 433222 614218 468986 614454
rect 469222 614218 504986 614454
rect 505222 614218 540986 614454
rect 541222 614218 576986 614454
rect 577222 614218 585502 614454
rect 585738 614218 586860 614454
rect -2936 614134 586860 614218
rect -2936 613898 -1814 614134
rect -1578 613898 986 614134
rect 1222 613898 36986 614134
rect 37222 613898 136536 614134
rect 136772 613898 144986 614134
rect 145222 613898 180986 614134
rect 181222 613898 266536 614134
rect 266772 613898 288986 614134
rect 289222 613898 386536 614134
rect 386772 613898 396986 614134
rect 397222 613898 432986 614134
rect 433222 613898 468986 614134
rect 469222 613898 504986 614134
rect 505222 613898 540986 614134
rect 541222 613898 576986 614134
rect 577222 613898 585502 614134
rect 585738 613898 586860 614134
rect -2936 613876 586860 613898
rect -1996 613874 -1396 613876
rect 804 613874 1404 613876
rect 36804 613874 37404 613876
rect 136494 613874 136814 613876
rect 144804 613874 145404 613876
rect 180804 613874 181404 613876
rect 266494 613874 266814 613876
rect 288804 613874 289404 613876
rect 386494 613874 386814 613876
rect 396804 613874 397404 613876
rect 432804 613874 433404 613876
rect 468804 613874 469404 613876
rect 504804 613874 505404 613876
rect 540804 613874 541404 613876
rect 576804 613874 577404 613876
rect 585320 613874 585920 613876
rect -8576 607276 -7976 607278
rect 29604 607276 30204 607278
rect 136938 607276 137262 607278
rect 173604 607276 174204 607278
rect 266938 607276 267262 607278
rect 281604 607276 282204 607278
rect 386938 607276 387262 607278
rect 425604 607276 426204 607278
rect 461604 607276 462204 607278
rect 497604 607276 498204 607278
rect 533604 607276 534204 607278
rect 569604 607276 570204 607278
rect 591900 607276 592500 607278
rect -8576 607254 592500 607276
rect -8576 607018 -8394 607254
rect -8158 607018 29786 607254
rect 30022 607018 136982 607254
rect 137218 607018 173786 607254
rect 174022 607018 266982 607254
rect 267218 607018 281786 607254
rect 282022 607018 386982 607254
rect 387218 607018 425786 607254
rect 426022 607018 461786 607254
rect 462022 607018 497786 607254
rect 498022 607018 533786 607254
rect 534022 607018 569786 607254
rect 570022 607018 592082 607254
rect 592318 607018 592500 607254
rect -8576 606934 592500 607018
rect -8576 606698 -8394 606934
rect -8158 606698 29786 606934
rect 30022 606698 136982 606934
rect 137218 606698 173786 606934
rect 174022 606698 266982 606934
rect 267218 606698 281786 606934
rect 282022 606698 386982 606934
rect 387218 606698 425786 606934
rect 426022 606698 461786 606934
rect 462022 606698 497786 606934
rect 498022 606698 533786 606934
rect 534022 606698 569786 606934
rect 570022 606698 592082 606934
rect 592318 606698 592500 606934
rect -8576 606676 592500 606698
rect -8576 606674 -7976 606676
rect 29604 606674 30204 606676
rect 136938 606674 137262 606676
rect 173604 606674 174204 606676
rect 266938 606674 267262 606676
rect 281604 606674 282204 606676
rect 386938 606674 387262 606676
rect 425604 606674 426204 606676
rect 461604 606674 462204 606676
rect 497604 606674 498204 606676
rect 533604 606674 534204 606676
rect 569604 606674 570204 606676
rect 591900 606674 592500 606676
rect -6696 603676 -6096 603678
rect 26004 603676 26604 603678
rect 136938 603676 137262 603678
rect 170004 603676 170604 603678
rect 266938 603676 267262 603678
rect 278004 603676 278604 603678
rect 386938 603676 387262 603678
rect 422004 603676 422604 603678
rect 458004 603676 458604 603678
rect 494004 603676 494604 603678
rect 530004 603676 530604 603678
rect 566004 603676 566604 603678
rect 590020 603676 590620 603678
rect -6696 603654 590620 603676
rect -6696 603418 -6514 603654
rect -6278 603418 26186 603654
rect 26422 603418 136982 603654
rect 137218 603418 170186 603654
rect 170422 603418 266982 603654
rect 267218 603418 278186 603654
rect 278422 603418 386982 603654
rect 387218 603418 422186 603654
rect 422422 603418 458186 603654
rect 458422 603418 494186 603654
rect 494422 603418 530186 603654
rect 530422 603418 566186 603654
rect 566422 603418 590202 603654
rect 590438 603418 590620 603654
rect -6696 603334 590620 603418
rect -6696 603098 -6514 603334
rect -6278 603098 26186 603334
rect 26422 603098 136982 603334
rect 137218 603098 170186 603334
rect 170422 603098 266982 603334
rect 267218 603098 278186 603334
rect 278422 603098 386982 603334
rect 387218 603098 422186 603334
rect 422422 603098 458186 603334
rect 458422 603098 494186 603334
rect 494422 603098 530186 603334
rect 530422 603098 566186 603334
rect 566422 603098 590202 603334
rect 590438 603098 590620 603334
rect -6696 603076 590620 603098
rect -6696 603074 -6096 603076
rect 26004 603074 26604 603076
rect 136938 603074 137262 603076
rect 170004 603074 170604 603076
rect 266938 603074 267262 603076
rect 278004 603074 278604 603076
rect 386938 603074 387262 603076
rect 422004 603074 422604 603076
rect 458004 603074 458604 603076
rect 494004 603074 494604 603076
rect 530004 603074 530604 603076
rect 566004 603074 566604 603076
rect 590020 603074 590620 603076
rect -4816 600076 -4216 600078
rect 22404 600076 23004 600078
rect 136938 600076 137262 600078
rect 166404 600076 167004 600078
rect 266938 600076 267262 600078
rect 274404 600076 275004 600078
rect 386938 600076 387262 600078
rect 418404 600076 419004 600078
rect 454404 600076 455004 600078
rect 490404 600076 491004 600078
rect 526404 600076 527004 600078
rect 562404 600076 563004 600078
rect 588140 600076 588740 600078
rect -4816 600054 588740 600076
rect -4816 599818 -4634 600054
rect -4398 599818 22586 600054
rect 22822 599818 136982 600054
rect 137218 599818 166586 600054
rect 166822 599818 266982 600054
rect 267218 599818 274586 600054
rect 274822 599818 386982 600054
rect 387218 599818 418586 600054
rect 418822 599818 454586 600054
rect 454822 599818 490586 600054
rect 490822 599818 526586 600054
rect 526822 599818 562586 600054
rect 562822 599818 588322 600054
rect 588558 599818 588740 600054
rect -4816 599734 588740 599818
rect -4816 599498 -4634 599734
rect -4398 599498 22586 599734
rect 22822 599498 136982 599734
rect 137218 599498 166586 599734
rect 166822 599498 266982 599734
rect 267218 599498 274586 599734
rect 274822 599498 386982 599734
rect 387218 599498 418586 599734
rect 418822 599498 454586 599734
rect 454822 599498 490586 599734
rect 490822 599498 526586 599734
rect 526822 599498 562586 599734
rect 562822 599498 588322 599734
rect 588558 599498 588740 599734
rect -4816 599476 588740 599498
rect -4816 599474 -4216 599476
rect 22404 599474 23004 599476
rect 136938 599474 137262 599476
rect 166404 599474 167004 599476
rect 266938 599474 267262 599476
rect 274404 599474 275004 599476
rect 386938 599474 387262 599476
rect 418404 599474 419004 599476
rect 454404 599474 455004 599476
rect 490404 599474 491004 599476
rect 526404 599474 527004 599476
rect 562404 599474 563004 599476
rect 588140 599474 588740 599476
rect -2936 596476 -2336 596478
rect 18804 596476 19404 596478
rect 54804 596476 55404 596478
rect 136938 596476 137262 596478
rect 162804 596476 163404 596478
rect 266938 596476 267262 596478
rect 270804 596476 271404 596478
rect 386938 596476 387262 596478
rect 414804 596476 415404 596478
rect 450804 596476 451404 596478
rect 486804 596476 487404 596478
rect 522804 596476 523404 596478
rect 558804 596476 559404 596478
rect 586260 596476 586860 596478
rect -2936 596454 586860 596476
rect -2936 596218 -2754 596454
rect -2518 596218 18986 596454
rect 19222 596218 54986 596454
rect 55222 596218 136982 596454
rect 137218 596218 162986 596454
rect 163222 596218 266982 596454
rect 267218 596218 270986 596454
rect 271222 596218 386982 596454
rect 387218 596218 414986 596454
rect 415222 596218 450986 596454
rect 451222 596218 486986 596454
rect 487222 596218 522986 596454
rect 523222 596218 558986 596454
rect 559222 596218 586442 596454
rect 586678 596218 586860 596454
rect -2936 596134 586860 596218
rect -2936 595898 -2754 596134
rect -2518 595898 18986 596134
rect 19222 595898 54986 596134
rect 55222 595898 136982 596134
rect 137218 595898 162986 596134
rect 163222 595898 266982 596134
rect 267218 595898 270986 596134
rect 271222 595898 386982 596134
rect 387218 595898 414986 596134
rect 415222 595898 450986 596134
rect 451222 595898 486986 596134
rect 487222 595898 522986 596134
rect 523222 595898 558986 596134
rect 559222 595898 586442 596134
rect 586678 595898 586860 596134
rect -2936 595876 586860 595898
rect -2936 595874 -2336 595876
rect 18804 595874 19404 595876
rect 54804 595874 55404 595876
rect 136938 595874 137262 595876
rect 162804 595874 163404 595876
rect 266938 595874 267262 595876
rect 270804 595874 271404 595876
rect 386938 595874 387262 595876
rect 414804 595874 415404 595876
rect 450804 595874 451404 595876
rect 486804 595874 487404 595876
rect 522804 595874 523404 595876
rect 558804 595874 559404 595876
rect 586260 595874 586860 595876
rect -7636 589276 -7036 589278
rect 11604 589276 12204 589278
rect 47604 589276 48204 589278
rect 136494 589276 136814 589278
rect 155604 589276 156204 589278
rect 266494 589276 266814 589278
rect 299604 589276 300204 589278
rect 386494 589276 386814 589278
rect 407604 589276 408204 589278
rect 443604 589276 444204 589278
rect 479604 589276 480204 589278
rect 515604 589276 516204 589278
rect 551604 589276 552204 589278
rect 590960 589276 591560 589278
rect -8576 589254 592500 589276
rect -8576 589018 -7454 589254
rect -7218 589018 11786 589254
rect 12022 589018 47786 589254
rect 48022 589018 136536 589254
rect 136772 589018 155786 589254
rect 156022 589018 266536 589254
rect 266772 589018 299786 589254
rect 300022 589018 386536 589254
rect 386772 589018 407786 589254
rect 408022 589018 443786 589254
rect 444022 589018 479786 589254
rect 480022 589018 515786 589254
rect 516022 589018 551786 589254
rect 552022 589018 591142 589254
rect 591378 589018 592500 589254
rect -8576 588934 592500 589018
rect -8576 588698 -7454 588934
rect -7218 588698 11786 588934
rect 12022 588698 47786 588934
rect 48022 588698 136536 588934
rect 136772 588698 155786 588934
rect 156022 588698 266536 588934
rect 266772 588698 299786 588934
rect 300022 588698 386536 588934
rect 386772 588698 407786 588934
rect 408022 588698 443786 588934
rect 444022 588698 479786 588934
rect 480022 588698 515786 588934
rect 516022 588698 551786 588934
rect 552022 588698 591142 588934
rect 591378 588698 592500 588934
rect -8576 588676 592500 588698
rect -7636 588674 -7036 588676
rect 11604 588674 12204 588676
rect 47604 588674 48204 588676
rect 136494 588674 136814 588676
rect 155604 588674 156204 588676
rect 266494 588674 266814 588676
rect 299604 588674 300204 588676
rect 386494 588674 386814 588676
rect 407604 588674 408204 588676
rect 443604 588674 444204 588676
rect 479604 588674 480204 588676
rect 515604 588674 516204 588676
rect 551604 588674 552204 588676
rect 590960 588674 591560 588676
rect -5756 585676 -5156 585678
rect 8004 585676 8604 585678
rect 44004 585676 44604 585678
rect 136494 585676 136814 585678
rect 152004 585676 152604 585678
rect 266494 585676 266814 585678
rect 296004 585676 296604 585678
rect 386494 585676 386814 585678
rect 404004 585676 404604 585678
rect 440004 585676 440604 585678
rect 476004 585676 476604 585678
rect 512004 585676 512604 585678
rect 548004 585676 548604 585678
rect 589080 585676 589680 585678
rect -6696 585654 590620 585676
rect -6696 585418 -5574 585654
rect -5338 585418 8186 585654
rect 8422 585418 44186 585654
rect 44422 585418 136536 585654
rect 136772 585418 152186 585654
rect 152422 585418 266536 585654
rect 266772 585418 296186 585654
rect 296422 585418 386536 585654
rect 386772 585418 404186 585654
rect 404422 585418 440186 585654
rect 440422 585418 476186 585654
rect 476422 585418 512186 585654
rect 512422 585418 548186 585654
rect 548422 585418 589262 585654
rect 589498 585418 590620 585654
rect -6696 585334 590620 585418
rect -6696 585098 -5574 585334
rect -5338 585098 8186 585334
rect 8422 585098 44186 585334
rect 44422 585098 136536 585334
rect 136772 585098 152186 585334
rect 152422 585098 266536 585334
rect 266772 585098 296186 585334
rect 296422 585098 386536 585334
rect 386772 585098 404186 585334
rect 404422 585098 440186 585334
rect 440422 585098 476186 585334
rect 476422 585098 512186 585334
rect 512422 585098 548186 585334
rect 548422 585098 589262 585334
rect 589498 585098 590620 585334
rect -6696 585076 590620 585098
rect -5756 585074 -5156 585076
rect 8004 585074 8604 585076
rect 44004 585074 44604 585076
rect 136494 585074 136814 585076
rect 152004 585074 152604 585076
rect 266494 585074 266814 585076
rect 296004 585074 296604 585076
rect 386494 585074 386814 585076
rect 404004 585074 404604 585076
rect 440004 585074 440604 585076
rect 476004 585074 476604 585076
rect 512004 585074 512604 585076
rect 548004 585074 548604 585076
rect 589080 585074 589680 585076
rect -3876 582076 -3276 582078
rect 4404 582076 5004 582078
rect 40404 582076 41004 582078
rect 136494 582076 136814 582078
rect 148404 582076 149004 582078
rect 184404 582076 185004 582078
rect 266494 582076 266814 582078
rect 292404 582076 293004 582078
rect 386494 582076 386814 582078
rect 400404 582076 401004 582078
rect 436404 582076 437004 582078
rect 472404 582076 473004 582078
rect 508404 582076 509004 582078
rect 544404 582076 545004 582078
rect 580404 582076 581004 582078
rect 587200 582076 587800 582078
rect -4816 582054 588740 582076
rect -4816 581818 -3694 582054
rect -3458 581818 4586 582054
rect 4822 581818 40586 582054
rect 40822 581818 136536 582054
rect 136772 581818 148586 582054
rect 148822 581818 184586 582054
rect 184822 581818 266536 582054
rect 266772 581818 292586 582054
rect 292822 581818 386536 582054
rect 386772 581818 400586 582054
rect 400822 581818 436586 582054
rect 436822 581818 472586 582054
rect 472822 581818 508586 582054
rect 508822 581818 544586 582054
rect 544822 581818 580586 582054
rect 580822 581818 587382 582054
rect 587618 581818 588740 582054
rect -4816 581734 588740 581818
rect -4816 581498 -3694 581734
rect -3458 581498 4586 581734
rect 4822 581498 40586 581734
rect 40822 581498 136536 581734
rect 136772 581498 148586 581734
rect 148822 581498 184586 581734
rect 184822 581498 266536 581734
rect 266772 581498 292586 581734
rect 292822 581498 386536 581734
rect 386772 581498 400586 581734
rect 400822 581498 436586 581734
rect 436822 581498 472586 581734
rect 472822 581498 508586 581734
rect 508822 581498 544586 581734
rect 544822 581498 580586 581734
rect 580822 581498 587382 581734
rect 587618 581498 588740 581734
rect -4816 581476 588740 581498
rect -3876 581474 -3276 581476
rect 4404 581474 5004 581476
rect 40404 581474 41004 581476
rect 136494 581474 136814 581476
rect 148404 581474 149004 581476
rect 184404 581474 185004 581476
rect 266494 581474 266814 581476
rect 292404 581474 293004 581476
rect 386494 581474 386814 581476
rect 400404 581474 401004 581476
rect 436404 581474 437004 581476
rect 472404 581474 473004 581476
rect 508404 581474 509004 581476
rect 544404 581474 545004 581476
rect 580404 581474 581004 581476
rect 587200 581474 587800 581476
rect -1996 578476 -1396 578478
rect 804 578476 1404 578478
rect 36804 578476 37404 578478
rect 136494 578476 136814 578478
rect 144804 578476 145404 578478
rect 180804 578476 181404 578478
rect 266494 578476 266814 578478
rect 288804 578476 289404 578478
rect 386494 578476 386814 578478
rect 396804 578476 397404 578478
rect 432804 578476 433404 578478
rect 468804 578476 469404 578478
rect 504804 578476 505404 578478
rect 540804 578476 541404 578478
rect 576804 578476 577404 578478
rect 585320 578476 585920 578478
rect -2936 578454 586860 578476
rect -2936 578218 -1814 578454
rect -1578 578218 986 578454
rect 1222 578218 36986 578454
rect 37222 578218 136536 578454
rect 136772 578218 144986 578454
rect 145222 578218 180986 578454
rect 181222 578218 266536 578454
rect 266772 578218 288986 578454
rect 289222 578218 386536 578454
rect 386772 578218 396986 578454
rect 397222 578218 432986 578454
rect 433222 578218 468986 578454
rect 469222 578218 504986 578454
rect 505222 578218 540986 578454
rect 541222 578218 576986 578454
rect 577222 578218 585502 578454
rect 585738 578218 586860 578454
rect -2936 578134 586860 578218
rect -2936 577898 -1814 578134
rect -1578 577898 986 578134
rect 1222 577898 36986 578134
rect 37222 577898 136536 578134
rect 136772 577898 144986 578134
rect 145222 577898 180986 578134
rect 181222 577898 266536 578134
rect 266772 577898 288986 578134
rect 289222 577898 386536 578134
rect 386772 577898 396986 578134
rect 397222 577898 432986 578134
rect 433222 577898 468986 578134
rect 469222 577898 504986 578134
rect 505222 577898 540986 578134
rect 541222 577898 576986 578134
rect 577222 577898 585502 578134
rect 585738 577898 586860 578134
rect -2936 577876 586860 577898
rect -1996 577874 -1396 577876
rect 804 577874 1404 577876
rect 36804 577874 37404 577876
rect 136494 577874 136814 577876
rect 144804 577874 145404 577876
rect 180804 577874 181404 577876
rect 266494 577874 266814 577876
rect 288804 577874 289404 577876
rect 386494 577874 386814 577876
rect 396804 577874 397404 577876
rect 432804 577874 433404 577876
rect 468804 577874 469404 577876
rect 504804 577874 505404 577876
rect 540804 577874 541404 577876
rect 576804 577874 577404 577876
rect 585320 577874 585920 577876
rect -8576 571276 -7976 571278
rect 29604 571276 30204 571278
rect 136938 571276 137262 571278
rect 173604 571276 174204 571278
rect 266938 571276 267262 571278
rect 281604 571276 282204 571278
rect 386938 571276 387262 571278
rect 425604 571276 426204 571278
rect 461604 571276 462204 571278
rect 497604 571276 498204 571278
rect 533604 571276 534204 571278
rect 569604 571276 570204 571278
rect 591900 571276 592500 571278
rect -8576 571254 592500 571276
rect -8576 571018 -8394 571254
rect -8158 571018 29786 571254
rect 30022 571018 136982 571254
rect 137218 571018 173786 571254
rect 174022 571018 266982 571254
rect 267218 571018 281786 571254
rect 282022 571018 386982 571254
rect 387218 571018 425786 571254
rect 426022 571018 461786 571254
rect 462022 571018 497786 571254
rect 498022 571018 533786 571254
rect 534022 571018 569786 571254
rect 570022 571018 592082 571254
rect 592318 571018 592500 571254
rect -8576 570934 592500 571018
rect -8576 570698 -8394 570934
rect -8158 570698 29786 570934
rect 30022 570698 136982 570934
rect 137218 570698 173786 570934
rect 174022 570698 266982 570934
rect 267218 570698 281786 570934
rect 282022 570698 386982 570934
rect 387218 570698 425786 570934
rect 426022 570698 461786 570934
rect 462022 570698 497786 570934
rect 498022 570698 533786 570934
rect 534022 570698 569786 570934
rect 570022 570698 592082 570934
rect 592318 570698 592500 570934
rect -8576 570676 592500 570698
rect -8576 570674 -7976 570676
rect 29604 570674 30204 570676
rect 136938 570674 137262 570676
rect 173604 570674 174204 570676
rect 266938 570674 267262 570676
rect 281604 570674 282204 570676
rect 386938 570674 387262 570676
rect 425604 570674 426204 570676
rect 461604 570674 462204 570676
rect 497604 570674 498204 570676
rect 533604 570674 534204 570676
rect 569604 570674 570204 570676
rect 591900 570674 592500 570676
rect -6696 567676 -6096 567678
rect 26004 567676 26604 567678
rect 136938 567676 137262 567678
rect 170004 567676 170604 567678
rect 266938 567676 267262 567678
rect 278004 567676 278604 567678
rect 386938 567676 387262 567678
rect 422004 567676 422604 567678
rect 458004 567676 458604 567678
rect 494004 567676 494604 567678
rect 530004 567676 530604 567678
rect 566004 567676 566604 567678
rect 590020 567676 590620 567678
rect -6696 567654 590620 567676
rect -6696 567418 -6514 567654
rect -6278 567418 26186 567654
rect 26422 567418 136982 567654
rect 137218 567418 170186 567654
rect 170422 567418 266982 567654
rect 267218 567418 278186 567654
rect 278422 567418 386982 567654
rect 387218 567418 422186 567654
rect 422422 567418 458186 567654
rect 458422 567418 494186 567654
rect 494422 567418 530186 567654
rect 530422 567418 566186 567654
rect 566422 567418 590202 567654
rect 590438 567418 590620 567654
rect -6696 567334 590620 567418
rect -6696 567098 -6514 567334
rect -6278 567098 26186 567334
rect 26422 567098 136982 567334
rect 137218 567098 170186 567334
rect 170422 567098 266982 567334
rect 267218 567098 278186 567334
rect 278422 567098 386982 567334
rect 387218 567098 422186 567334
rect 422422 567098 458186 567334
rect 458422 567098 494186 567334
rect 494422 567098 530186 567334
rect 530422 567098 566186 567334
rect 566422 567098 590202 567334
rect 590438 567098 590620 567334
rect -6696 567076 590620 567098
rect -6696 567074 -6096 567076
rect 26004 567074 26604 567076
rect 136938 567074 137262 567076
rect 170004 567074 170604 567076
rect 266938 567074 267262 567076
rect 278004 567074 278604 567076
rect 386938 567074 387262 567076
rect 422004 567074 422604 567076
rect 458004 567074 458604 567076
rect 494004 567074 494604 567076
rect 530004 567074 530604 567076
rect 566004 567074 566604 567076
rect 590020 567074 590620 567076
rect -4816 564076 -4216 564078
rect 22404 564076 23004 564078
rect 136938 564076 137262 564078
rect 166404 564076 167004 564078
rect 266938 564076 267262 564078
rect 274404 564076 275004 564078
rect 386938 564076 387262 564078
rect 418404 564076 419004 564078
rect 454404 564076 455004 564078
rect 490404 564076 491004 564078
rect 526404 564076 527004 564078
rect 562404 564076 563004 564078
rect 588140 564076 588740 564078
rect -4816 564054 588740 564076
rect -4816 563818 -4634 564054
rect -4398 563818 22586 564054
rect 22822 563818 136982 564054
rect 137218 563818 166586 564054
rect 166822 563818 266982 564054
rect 267218 563818 274586 564054
rect 274822 563818 386982 564054
rect 387218 563818 418586 564054
rect 418822 563818 454586 564054
rect 454822 563818 490586 564054
rect 490822 563818 526586 564054
rect 526822 563818 562586 564054
rect 562822 563818 588322 564054
rect 588558 563818 588740 564054
rect -4816 563734 588740 563818
rect -4816 563498 -4634 563734
rect -4398 563498 22586 563734
rect 22822 563498 136982 563734
rect 137218 563498 166586 563734
rect 166822 563498 266982 563734
rect 267218 563498 274586 563734
rect 274822 563498 386982 563734
rect 387218 563498 418586 563734
rect 418822 563498 454586 563734
rect 454822 563498 490586 563734
rect 490822 563498 526586 563734
rect 526822 563498 562586 563734
rect 562822 563498 588322 563734
rect 588558 563498 588740 563734
rect -4816 563476 588740 563498
rect -4816 563474 -4216 563476
rect 22404 563474 23004 563476
rect 136938 563474 137262 563476
rect 166404 563474 167004 563476
rect 266938 563474 267262 563476
rect 274404 563474 275004 563476
rect 386938 563474 387262 563476
rect 418404 563474 419004 563476
rect 454404 563474 455004 563476
rect 490404 563474 491004 563476
rect 526404 563474 527004 563476
rect 562404 563474 563004 563476
rect 588140 563474 588740 563476
rect -2936 560476 -2336 560478
rect 18804 560476 19404 560478
rect 54804 560476 55404 560478
rect 162804 560476 163404 560478
rect 270804 560476 271404 560478
rect 414804 560476 415404 560478
rect 450804 560476 451404 560478
rect 486804 560476 487404 560478
rect 522804 560476 523404 560478
rect 558804 560476 559404 560478
rect 586260 560476 586860 560478
rect -2936 560454 586860 560476
rect -2936 560218 -2754 560454
rect -2518 560218 18986 560454
rect 19222 560218 54986 560454
rect 55222 560218 162986 560454
rect 163222 560218 270986 560454
rect 271222 560218 414986 560454
rect 415222 560218 450986 560454
rect 451222 560218 486986 560454
rect 487222 560218 522986 560454
rect 523222 560218 558986 560454
rect 559222 560218 586442 560454
rect 586678 560218 586860 560454
rect -2936 560134 586860 560218
rect -2936 559898 -2754 560134
rect -2518 559898 18986 560134
rect 19222 559898 54986 560134
rect 55222 559898 162986 560134
rect 163222 559898 270986 560134
rect 271222 559898 414986 560134
rect 415222 559898 450986 560134
rect 451222 559898 486986 560134
rect 487222 559898 522986 560134
rect 523222 559898 558986 560134
rect 559222 559898 586442 560134
rect 586678 559898 586860 560134
rect -2936 559876 586860 559898
rect -2936 559874 -2336 559876
rect 18804 559874 19404 559876
rect 54804 559874 55404 559876
rect 162804 559874 163404 559876
rect 270804 559874 271404 559876
rect 414804 559874 415404 559876
rect 450804 559874 451404 559876
rect 486804 559874 487404 559876
rect 522804 559874 523404 559876
rect 558804 559874 559404 559876
rect 586260 559874 586860 559876
rect -7636 553276 -7036 553278
rect 11604 553276 12204 553278
rect 47604 553276 48204 553278
rect 83604 553276 84204 553278
rect 119604 553276 120204 553278
rect 155604 553276 156204 553278
rect 191604 553276 192204 553278
rect 227604 553276 228204 553278
rect 263604 553276 264204 553278
rect 299604 553276 300204 553278
rect 335604 553276 336204 553278
rect 371604 553276 372204 553278
rect 407604 553276 408204 553278
rect 443604 553276 444204 553278
rect 479604 553276 480204 553278
rect 515604 553276 516204 553278
rect 551604 553276 552204 553278
rect 590960 553276 591560 553278
rect -8576 553254 592500 553276
rect -8576 553018 -7454 553254
rect -7218 553018 11786 553254
rect 12022 553018 47786 553254
rect 48022 553018 83786 553254
rect 84022 553018 119786 553254
rect 120022 553018 155786 553254
rect 156022 553018 191786 553254
rect 192022 553018 227786 553254
rect 228022 553018 263786 553254
rect 264022 553018 299786 553254
rect 300022 553018 335786 553254
rect 336022 553018 371786 553254
rect 372022 553018 407786 553254
rect 408022 553018 443786 553254
rect 444022 553018 479786 553254
rect 480022 553018 515786 553254
rect 516022 553018 551786 553254
rect 552022 553018 591142 553254
rect 591378 553018 592500 553254
rect -8576 552934 592500 553018
rect -8576 552698 -7454 552934
rect -7218 552698 11786 552934
rect 12022 552698 47786 552934
rect 48022 552698 83786 552934
rect 84022 552698 119786 552934
rect 120022 552698 155786 552934
rect 156022 552698 191786 552934
rect 192022 552698 227786 552934
rect 228022 552698 263786 552934
rect 264022 552698 299786 552934
rect 300022 552698 335786 552934
rect 336022 552698 371786 552934
rect 372022 552698 407786 552934
rect 408022 552698 443786 552934
rect 444022 552698 479786 552934
rect 480022 552698 515786 552934
rect 516022 552698 551786 552934
rect 552022 552698 591142 552934
rect 591378 552698 592500 552934
rect -8576 552676 592500 552698
rect -7636 552674 -7036 552676
rect 11604 552674 12204 552676
rect 47604 552674 48204 552676
rect 83604 552674 84204 552676
rect 119604 552674 120204 552676
rect 155604 552674 156204 552676
rect 191604 552674 192204 552676
rect 227604 552674 228204 552676
rect 263604 552674 264204 552676
rect 299604 552674 300204 552676
rect 335604 552674 336204 552676
rect 371604 552674 372204 552676
rect 407604 552674 408204 552676
rect 443604 552674 444204 552676
rect 479604 552674 480204 552676
rect 515604 552674 516204 552676
rect 551604 552674 552204 552676
rect 590960 552674 591560 552676
rect -5756 549676 -5156 549678
rect 8004 549676 8604 549678
rect 44004 549676 44604 549678
rect 80004 549676 80604 549678
rect 116004 549676 116604 549678
rect 152004 549676 152604 549678
rect 188004 549676 188604 549678
rect 224004 549676 224604 549678
rect 260004 549676 260604 549678
rect 296004 549676 296604 549678
rect 332004 549676 332604 549678
rect 368004 549676 368604 549678
rect 404004 549676 404604 549678
rect 440004 549676 440604 549678
rect 476004 549676 476604 549678
rect 512004 549676 512604 549678
rect 548004 549676 548604 549678
rect 589080 549676 589680 549678
rect -6696 549654 590620 549676
rect -6696 549418 -5574 549654
rect -5338 549418 8186 549654
rect 8422 549418 44186 549654
rect 44422 549418 80186 549654
rect 80422 549418 116186 549654
rect 116422 549418 152186 549654
rect 152422 549418 188186 549654
rect 188422 549418 224186 549654
rect 224422 549418 260186 549654
rect 260422 549418 296186 549654
rect 296422 549418 332186 549654
rect 332422 549418 368186 549654
rect 368422 549418 404186 549654
rect 404422 549418 440186 549654
rect 440422 549418 476186 549654
rect 476422 549418 512186 549654
rect 512422 549418 548186 549654
rect 548422 549418 589262 549654
rect 589498 549418 590620 549654
rect -6696 549334 590620 549418
rect -6696 549098 -5574 549334
rect -5338 549098 8186 549334
rect 8422 549098 44186 549334
rect 44422 549098 80186 549334
rect 80422 549098 116186 549334
rect 116422 549098 152186 549334
rect 152422 549098 188186 549334
rect 188422 549098 224186 549334
rect 224422 549098 260186 549334
rect 260422 549098 296186 549334
rect 296422 549098 332186 549334
rect 332422 549098 368186 549334
rect 368422 549098 404186 549334
rect 404422 549098 440186 549334
rect 440422 549098 476186 549334
rect 476422 549098 512186 549334
rect 512422 549098 548186 549334
rect 548422 549098 589262 549334
rect 589498 549098 590620 549334
rect -6696 549076 590620 549098
rect -5756 549074 -5156 549076
rect 8004 549074 8604 549076
rect 44004 549074 44604 549076
rect 80004 549074 80604 549076
rect 116004 549074 116604 549076
rect 152004 549074 152604 549076
rect 188004 549074 188604 549076
rect 224004 549074 224604 549076
rect 260004 549074 260604 549076
rect 296004 549074 296604 549076
rect 332004 549074 332604 549076
rect 368004 549074 368604 549076
rect 404004 549074 404604 549076
rect 440004 549074 440604 549076
rect 476004 549074 476604 549076
rect 512004 549074 512604 549076
rect 548004 549074 548604 549076
rect 589080 549074 589680 549076
rect -3876 546076 -3276 546078
rect 4404 546076 5004 546078
rect 40404 546076 41004 546078
rect 76404 546076 77004 546078
rect 112404 546076 113004 546078
rect 148404 546076 149004 546078
rect 184404 546076 185004 546078
rect 220404 546076 221004 546078
rect 256404 546076 257004 546078
rect 292404 546076 293004 546078
rect 328404 546076 329004 546078
rect 364404 546076 365004 546078
rect 400404 546076 401004 546078
rect 436404 546076 437004 546078
rect 472404 546076 473004 546078
rect 508404 546076 509004 546078
rect 544404 546076 545004 546078
rect 580404 546076 581004 546078
rect 587200 546076 587800 546078
rect -4816 546054 588740 546076
rect -4816 545818 -3694 546054
rect -3458 545818 4586 546054
rect 4822 545818 40586 546054
rect 40822 545818 76586 546054
rect 76822 545818 112586 546054
rect 112822 545818 148586 546054
rect 148822 545818 184586 546054
rect 184822 545818 220586 546054
rect 220822 545818 256586 546054
rect 256822 545818 292586 546054
rect 292822 545818 328586 546054
rect 328822 545818 364586 546054
rect 364822 545818 400586 546054
rect 400822 545818 436586 546054
rect 436822 545818 472586 546054
rect 472822 545818 508586 546054
rect 508822 545818 544586 546054
rect 544822 545818 580586 546054
rect 580822 545818 587382 546054
rect 587618 545818 588740 546054
rect -4816 545734 588740 545818
rect -4816 545498 -3694 545734
rect -3458 545498 4586 545734
rect 4822 545498 40586 545734
rect 40822 545498 76586 545734
rect 76822 545498 112586 545734
rect 112822 545498 148586 545734
rect 148822 545498 184586 545734
rect 184822 545498 220586 545734
rect 220822 545498 256586 545734
rect 256822 545498 292586 545734
rect 292822 545498 328586 545734
rect 328822 545498 364586 545734
rect 364822 545498 400586 545734
rect 400822 545498 436586 545734
rect 436822 545498 472586 545734
rect 472822 545498 508586 545734
rect 508822 545498 544586 545734
rect 544822 545498 580586 545734
rect 580822 545498 587382 545734
rect 587618 545498 588740 545734
rect -4816 545476 588740 545498
rect -3876 545474 -3276 545476
rect 4404 545474 5004 545476
rect 40404 545474 41004 545476
rect 76404 545474 77004 545476
rect 112404 545474 113004 545476
rect 148404 545474 149004 545476
rect 184404 545474 185004 545476
rect 220404 545474 221004 545476
rect 256404 545474 257004 545476
rect 292404 545474 293004 545476
rect 328404 545474 329004 545476
rect 364404 545474 365004 545476
rect 400404 545474 401004 545476
rect 436404 545474 437004 545476
rect 472404 545474 473004 545476
rect 508404 545474 509004 545476
rect 544404 545474 545004 545476
rect 580404 545474 581004 545476
rect 587200 545474 587800 545476
rect -1996 542476 -1396 542478
rect 804 542476 1404 542478
rect 36804 542476 37404 542478
rect 288804 542476 289404 542478
rect 324804 542476 325404 542478
rect 360804 542476 361404 542478
rect 396804 542476 397404 542478
rect 432804 542476 433404 542478
rect 468804 542476 469404 542478
rect 504804 542476 505404 542478
rect 540804 542476 541404 542478
rect 576804 542476 577404 542478
rect 585320 542476 585920 542478
rect -2936 542454 586860 542476
rect -2936 542218 -1814 542454
rect -1578 542218 986 542454
rect 1222 542218 36986 542454
rect 37222 542218 288986 542454
rect 289222 542218 324986 542454
rect 325222 542218 360986 542454
rect 361222 542218 396986 542454
rect 397222 542218 432986 542454
rect 433222 542218 468986 542454
rect 469222 542218 504986 542454
rect 505222 542218 540986 542454
rect 541222 542218 576986 542454
rect 577222 542218 585502 542454
rect 585738 542218 586860 542454
rect -2936 542134 586860 542218
rect -2936 541898 -1814 542134
rect -1578 541898 986 542134
rect 1222 541898 36986 542134
rect 37222 541898 288986 542134
rect 289222 541898 324986 542134
rect 325222 541898 360986 542134
rect 361222 541898 396986 542134
rect 397222 541898 432986 542134
rect 433222 541898 468986 542134
rect 469222 541898 504986 542134
rect 505222 541898 540986 542134
rect 541222 541898 576986 542134
rect 577222 541898 585502 542134
rect 585738 541898 586860 542134
rect -2936 541876 586860 541898
rect -1996 541874 -1396 541876
rect 804 541874 1404 541876
rect 36804 541874 37404 541876
rect 288804 541874 289404 541876
rect 324804 541874 325404 541876
rect 360804 541874 361404 541876
rect 396804 541874 397404 541876
rect 432804 541874 433404 541876
rect 468804 541874 469404 541876
rect 504804 541874 505404 541876
rect 540804 541874 541404 541876
rect 576804 541874 577404 541876
rect 585320 541874 585920 541876
rect -8576 535276 -7976 535278
rect 29604 535276 30204 535278
rect 79568 535276 79888 535278
rect 317604 535276 318204 535278
rect 353604 535276 354204 535278
rect 389604 535276 390204 535278
rect 425604 535276 426204 535278
rect 461604 535276 462204 535278
rect 497604 535276 498204 535278
rect 533604 535276 534204 535278
rect 569604 535276 570204 535278
rect 591900 535276 592500 535278
rect -8576 535254 592500 535276
rect -8576 535018 -8394 535254
rect -8158 535018 29786 535254
rect 30022 535018 79610 535254
rect 79846 535018 317786 535254
rect 318022 535018 353786 535254
rect 354022 535018 389786 535254
rect 390022 535018 425786 535254
rect 426022 535018 461786 535254
rect 462022 535018 497786 535254
rect 498022 535018 533786 535254
rect 534022 535018 569786 535254
rect 570022 535018 592082 535254
rect 592318 535018 592500 535254
rect -8576 534934 592500 535018
rect -8576 534698 -8394 534934
rect -8158 534698 29786 534934
rect 30022 534698 79610 534934
rect 79846 534698 317786 534934
rect 318022 534698 353786 534934
rect 354022 534698 389786 534934
rect 390022 534698 425786 534934
rect 426022 534698 461786 534934
rect 462022 534698 497786 534934
rect 498022 534698 533786 534934
rect 534022 534698 569786 534934
rect 570022 534698 592082 534934
rect 592318 534698 592500 534934
rect -8576 534676 592500 534698
rect -8576 534674 -7976 534676
rect 29604 534674 30204 534676
rect 79568 534674 79888 534676
rect 317604 534674 318204 534676
rect 353604 534674 354204 534676
rect 389604 534674 390204 534676
rect 425604 534674 426204 534676
rect 461604 534674 462204 534676
rect 497604 534674 498204 534676
rect 533604 534674 534204 534676
rect 569604 534674 570204 534676
rect 591900 534674 592500 534676
rect -6696 531676 -6096 531678
rect 26004 531676 26604 531678
rect 79568 531676 79888 531678
rect 314004 531676 314604 531678
rect 350004 531676 350604 531678
rect 386004 531676 386604 531678
rect 422004 531676 422604 531678
rect 458004 531676 458604 531678
rect 494004 531676 494604 531678
rect 530004 531676 530604 531678
rect 566004 531676 566604 531678
rect 590020 531676 590620 531678
rect -6696 531654 590620 531676
rect -6696 531418 -6514 531654
rect -6278 531418 26186 531654
rect 26422 531418 79610 531654
rect 79846 531418 314186 531654
rect 314422 531418 350186 531654
rect 350422 531418 386186 531654
rect 386422 531418 422186 531654
rect 422422 531418 458186 531654
rect 458422 531418 494186 531654
rect 494422 531418 530186 531654
rect 530422 531418 566186 531654
rect 566422 531418 590202 531654
rect 590438 531418 590620 531654
rect -6696 531334 590620 531418
rect -6696 531098 -6514 531334
rect -6278 531098 26186 531334
rect 26422 531098 79610 531334
rect 79846 531098 314186 531334
rect 314422 531098 350186 531334
rect 350422 531098 386186 531334
rect 386422 531098 422186 531334
rect 422422 531098 458186 531334
rect 458422 531098 494186 531334
rect 494422 531098 530186 531334
rect 530422 531098 566186 531334
rect 566422 531098 590202 531334
rect 590438 531098 590620 531334
rect -6696 531076 590620 531098
rect -6696 531074 -6096 531076
rect 26004 531074 26604 531076
rect 79568 531074 79888 531076
rect 314004 531074 314604 531076
rect 350004 531074 350604 531076
rect 386004 531074 386604 531076
rect 422004 531074 422604 531076
rect 458004 531074 458604 531076
rect 494004 531074 494604 531076
rect 530004 531074 530604 531076
rect 566004 531074 566604 531076
rect 590020 531074 590620 531076
rect -4816 528076 -4216 528078
rect 22404 528076 23004 528078
rect 79568 528076 79888 528078
rect 310404 528076 311004 528078
rect 346404 528076 347004 528078
rect 382404 528076 383004 528078
rect 418404 528076 419004 528078
rect 454404 528076 455004 528078
rect 490404 528076 491004 528078
rect 526404 528076 527004 528078
rect 562404 528076 563004 528078
rect 588140 528076 588740 528078
rect -4816 528054 588740 528076
rect -4816 527818 -4634 528054
rect -4398 527818 22586 528054
rect 22822 527818 79610 528054
rect 79846 527818 310586 528054
rect 310822 527818 346586 528054
rect 346822 527818 382586 528054
rect 382822 527818 418586 528054
rect 418822 527818 454586 528054
rect 454822 527818 490586 528054
rect 490822 527818 526586 528054
rect 526822 527818 562586 528054
rect 562822 527818 588322 528054
rect 588558 527818 588740 528054
rect -4816 527734 588740 527818
rect -4816 527498 -4634 527734
rect -4398 527498 22586 527734
rect 22822 527498 79610 527734
rect 79846 527498 310586 527734
rect 310822 527498 346586 527734
rect 346822 527498 382586 527734
rect 382822 527498 418586 527734
rect 418822 527498 454586 527734
rect 454822 527498 490586 527734
rect 490822 527498 526586 527734
rect 526822 527498 562586 527734
rect 562822 527498 588322 527734
rect 588558 527498 588740 527734
rect -4816 527476 588740 527498
rect -4816 527474 -4216 527476
rect 22404 527474 23004 527476
rect 79568 527474 79888 527476
rect 310404 527474 311004 527476
rect 346404 527474 347004 527476
rect 382404 527474 383004 527476
rect 418404 527474 419004 527476
rect 454404 527474 455004 527476
rect 490404 527474 491004 527476
rect 526404 527474 527004 527476
rect 562404 527474 563004 527476
rect 588140 527474 588740 527476
rect -2936 524476 -2336 524478
rect 18804 524476 19404 524478
rect 54804 524476 55404 524478
rect 79568 524476 79888 524478
rect 306804 524476 307404 524478
rect 342804 524476 343404 524478
rect 378804 524476 379404 524478
rect 414804 524476 415404 524478
rect 450804 524476 451404 524478
rect 486804 524476 487404 524478
rect 522804 524476 523404 524478
rect 558804 524476 559404 524478
rect 586260 524476 586860 524478
rect -2936 524454 586860 524476
rect -2936 524218 -2754 524454
rect -2518 524218 18986 524454
rect 19222 524218 54986 524454
rect 55222 524218 79610 524454
rect 79846 524218 306986 524454
rect 307222 524218 342986 524454
rect 343222 524218 378986 524454
rect 379222 524218 414986 524454
rect 415222 524218 450986 524454
rect 451222 524218 486986 524454
rect 487222 524218 522986 524454
rect 523222 524218 558986 524454
rect 559222 524218 586442 524454
rect 586678 524218 586860 524454
rect -2936 524134 586860 524218
rect -2936 523898 -2754 524134
rect -2518 523898 18986 524134
rect 19222 523898 54986 524134
rect 55222 523898 79610 524134
rect 79846 523898 306986 524134
rect 307222 523898 342986 524134
rect 343222 523898 378986 524134
rect 379222 523898 414986 524134
rect 415222 523898 450986 524134
rect 451222 523898 486986 524134
rect 487222 523898 522986 524134
rect 523222 523898 558986 524134
rect 559222 523898 586442 524134
rect 586678 523898 586860 524134
rect -2936 523876 586860 523898
rect -2936 523874 -2336 523876
rect 18804 523874 19404 523876
rect 54804 523874 55404 523876
rect 79568 523874 79888 523876
rect 306804 523874 307404 523876
rect 342804 523874 343404 523876
rect 378804 523874 379404 523876
rect 414804 523874 415404 523876
rect 450804 523874 451404 523876
rect 486804 523874 487404 523876
rect 522804 523874 523404 523876
rect 558804 523874 559404 523876
rect 586260 523874 586860 523876
rect -7636 517276 -7036 517278
rect 11604 517276 12204 517278
rect 47604 517276 48204 517278
rect 64208 517276 64528 517278
rect 299604 517276 300204 517278
rect 335604 517276 336204 517278
rect 371604 517276 372204 517278
rect 407604 517276 408204 517278
rect 443604 517276 444204 517278
rect 479604 517276 480204 517278
rect 515604 517276 516204 517278
rect 551604 517276 552204 517278
rect 590960 517276 591560 517278
rect -8576 517254 592500 517276
rect -8576 517018 -7454 517254
rect -7218 517018 11786 517254
rect 12022 517018 47786 517254
rect 48022 517018 64250 517254
rect 64486 517018 299786 517254
rect 300022 517018 335786 517254
rect 336022 517018 371786 517254
rect 372022 517018 407786 517254
rect 408022 517018 443786 517254
rect 444022 517018 479786 517254
rect 480022 517018 515786 517254
rect 516022 517018 551786 517254
rect 552022 517018 591142 517254
rect 591378 517018 592500 517254
rect -8576 516934 592500 517018
rect -8576 516698 -7454 516934
rect -7218 516698 11786 516934
rect 12022 516698 47786 516934
rect 48022 516698 64250 516934
rect 64486 516698 299786 516934
rect 300022 516698 335786 516934
rect 336022 516698 371786 516934
rect 372022 516698 407786 516934
rect 408022 516698 443786 516934
rect 444022 516698 479786 516934
rect 480022 516698 515786 516934
rect 516022 516698 551786 516934
rect 552022 516698 591142 516934
rect 591378 516698 592500 516934
rect -8576 516676 592500 516698
rect -7636 516674 -7036 516676
rect 11604 516674 12204 516676
rect 47604 516674 48204 516676
rect 64208 516674 64528 516676
rect 299604 516674 300204 516676
rect 335604 516674 336204 516676
rect 371604 516674 372204 516676
rect 407604 516674 408204 516676
rect 443604 516674 444204 516676
rect 479604 516674 480204 516676
rect 515604 516674 516204 516676
rect 551604 516674 552204 516676
rect 590960 516674 591560 516676
rect -5756 513676 -5156 513678
rect 8004 513676 8604 513678
rect 44004 513676 44604 513678
rect 64208 513676 64528 513678
rect 296004 513676 296604 513678
rect 332004 513676 332604 513678
rect 368004 513676 368604 513678
rect 404004 513676 404604 513678
rect 440004 513676 440604 513678
rect 476004 513676 476604 513678
rect 512004 513676 512604 513678
rect 548004 513676 548604 513678
rect 589080 513676 589680 513678
rect -6696 513654 590620 513676
rect -6696 513418 -5574 513654
rect -5338 513418 8186 513654
rect 8422 513418 44186 513654
rect 44422 513418 64250 513654
rect 64486 513418 296186 513654
rect 296422 513418 332186 513654
rect 332422 513418 368186 513654
rect 368422 513418 404186 513654
rect 404422 513418 440186 513654
rect 440422 513418 476186 513654
rect 476422 513418 512186 513654
rect 512422 513418 548186 513654
rect 548422 513418 589262 513654
rect 589498 513418 590620 513654
rect -6696 513334 590620 513418
rect -6696 513098 -5574 513334
rect -5338 513098 8186 513334
rect 8422 513098 44186 513334
rect 44422 513098 64250 513334
rect 64486 513098 296186 513334
rect 296422 513098 332186 513334
rect 332422 513098 368186 513334
rect 368422 513098 404186 513334
rect 404422 513098 440186 513334
rect 440422 513098 476186 513334
rect 476422 513098 512186 513334
rect 512422 513098 548186 513334
rect 548422 513098 589262 513334
rect 589498 513098 590620 513334
rect -6696 513076 590620 513098
rect -5756 513074 -5156 513076
rect 8004 513074 8604 513076
rect 44004 513074 44604 513076
rect 64208 513074 64528 513076
rect 296004 513074 296604 513076
rect 332004 513074 332604 513076
rect 368004 513074 368604 513076
rect 404004 513074 404604 513076
rect 440004 513074 440604 513076
rect 476004 513074 476604 513076
rect 512004 513074 512604 513076
rect 548004 513074 548604 513076
rect 589080 513074 589680 513076
rect -3876 510076 -3276 510078
rect 4404 510076 5004 510078
rect 40404 510076 41004 510078
rect 64208 510076 64528 510078
rect 292404 510076 293004 510078
rect 328404 510076 329004 510078
rect 364404 510076 365004 510078
rect 400404 510076 401004 510078
rect 436404 510076 437004 510078
rect 472404 510076 473004 510078
rect 508404 510076 509004 510078
rect 544404 510076 545004 510078
rect 580404 510076 581004 510078
rect 587200 510076 587800 510078
rect -4816 510054 588740 510076
rect -4816 509818 -3694 510054
rect -3458 509818 4586 510054
rect 4822 509818 40586 510054
rect 40822 509818 64250 510054
rect 64486 509818 292586 510054
rect 292822 509818 328586 510054
rect 328822 509818 364586 510054
rect 364822 509818 400586 510054
rect 400822 509818 436586 510054
rect 436822 509818 472586 510054
rect 472822 509818 508586 510054
rect 508822 509818 544586 510054
rect 544822 509818 580586 510054
rect 580822 509818 587382 510054
rect 587618 509818 588740 510054
rect -4816 509734 588740 509818
rect -4816 509498 -3694 509734
rect -3458 509498 4586 509734
rect 4822 509498 40586 509734
rect 40822 509498 64250 509734
rect 64486 509498 292586 509734
rect 292822 509498 328586 509734
rect 328822 509498 364586 509734
rect 364822 509498 400586 509734
rect 400822 509498 436586 509734
rect 436822 509498 472586 509734
rect 472822 509498 508586 509734
rect 508822 509498 544586 509734
rect 544822 509498 580586 509734
rect 580822 509498 587382 509734
rect 587618 509498 588740 509734
rect -4816 509476 588740 509498
rect -3876 509474 -3276 509476
rect 4404 509474 5004 509476
rect 40404 509474 41004 509476
rect 64208 509474 64528 509476
rect 292404 509474 293004 509476
rect 328404 509474 329004 509476
rect 364404 509474 365004 509476
rect 400404 509474 401004 509476
rect 436404 509474 437004 509476
rect 472404 509474 473004 509476
rect 508404 509474 509004 509476
rect 544404 509474 545004 509476
rect 580404 509474 581004 509476
rect 587200 509474 587800 509476
rect -1996 506476 -1396 506478
rect 804 506476 1404 506478
rect 36804 506476 37404 506478
rect 64208 506476 64528 506478
rect 288804 506476 289404 506478
rect 324804 506476 325404 506478
rect 360804 506476 361404 506478
rect 396804 506476 397404 506478
rect 432804 506476 433404 506478
rect 468804 506476 469404 506478
rect 504804 506476 505404 506478
rect 540804 506476 541404 506478
rect 576804 506476 577404 506478
rect 585320 506476 585920 506478
rect -2936 506454 586860 506476
rect -2936 506218 -1814 506454
rect -1578 506218 986 506454
rect 1222 506218 36986 506454
rect 37222 506218 64250 506454
rect 64486 506218 288986 506454
rect 289222 506218 324986 506454
rect 325222 506218 360986 506454
rect 361222 506218 396986 506454
rect 397222 506218 432986 506454
rect 433222 506218 468986 506454
rect 469222 506218 504986 506454
rect 505222 506218 540986 506454
rect 541222 506218 576986 506454
rect 577222 506218 585502 506454
rect 585738 506218 586860 506454
rect -2936 506134 586860 506218
rect -2936 505898 -1814 506134
rect -1578 505898 986 506134
rect 1222 505898 36986 506134
rect 37222 505898 64250 506134
rect 64486 505898 288986 506134
rect 289222 505898 324986 506134
rect 325222 505898 360986 506134
rect 361222 505898 396986 506134
rect 397222 505898 432986 506134
rect 433222 505898 468986 506134
rect 469222 505898 504986 506134
rect 505222 505898 540986 506134
rect 541222 505898 576986 506134
rect 577222 505898 585502 506134
rect 585738 505898 586860 506134
rect -2936 505876 586860 505898
rect -1996 505874 -1396 505876
rect 804 505874 1404 505876
rect 36804 505874 37404 505876
rect 64208 505874 64528 505876
rect 288804 505874 289404 505876
rect 324804 505874 325404 505876
rect 360804 505874 361404 505876
rect 396804 505874 397404 505876
rect 432804 505874 433404 505876
rect 468804 505874 469404 505876
rect 504804 505874 505404 505876
rect 540804 505874 541404 505876
rect 576804 505874 577404 505876
rect 585320 505874 585920 505876
rect -8576 499276 -7976 499278
rect 29604 499276 30204 499278
rect 79568 499276 79888 499278
rect 317604 499276 318204 499278
rect 353604 499276 354204 499278
rect 389604 499276 390204 499278
rect 425604 499276 426204 499278
rect 461604 499276 462204 499278
rect 497604 499276 498204 499278
rect 533604 499276 534204 499278
rect 569604 499276 570204 499278
rect 591900 499276 592500 499278
rect -8576 499254 592500 499276
rect -8576 499018 -8394 499254
rect -8158 499018 29786 499254
rect 30022 499018 79610 499254
rect 79846 499018 317786 499254
rect 318022 499018 353786 499254
rect 354022 499018 389786 499254
rect 390022 499018 425786 499254
rect 426022 499018 461786 499254
rect 462022 499018 497786 499254
rect 498022 499018 533786 499254
rect 534022 499018 569786 499254
rect 570022 499018 592082 499254
rect 592318 499018 592500 499254
rect -8576 498934 592500 499018
rect -8576 498698 -8394 498934
rect -8158 498698 29786 498934
rect 30022 498698 79610 498934
rect 79846 498698 317786 498934
rect 318022 498698 353786 498934
rect 354022 498698 389786 498934
rect 390022 498698 425786 498934
rect 426022 498698 461786 498934
rect 462022 498698 497786 498934
rect 498022 498698 533786 498934
rect 534022 498698 569786 498934
rect 570022 498698 592082 498934
rect 592318 498698 592500 498934
rect -8576 498676 592500 498698
rect -8576 498674 -7976 498676
rect 29604 498674 30204 498676
rect 79568 498674 79888 498676
rect 317604 498674 318204 498676
rect 353604 498674 354204 498676
rect 389604 498674 390204 498676
rect 425604 498674 426204 498676
rect 461604 498674 462204 498676
rect 497604 498674 498204 498676
rect 533604 498674 534204 498676
rect 569604 498674 570204 498676
rect 591900 498674 592500 498676
rect -6696 495676 -6096 495678
rect 26004 495676 26604 495678
rect 79568 495676 79888 495678
rect 314004 495676 314604 495678
rect 350004 495676 350604 495678
rect 386004 495676 386604 495678
rect 422004 495676 422604 495678
rect 458004 495676 458604 495678
rect 494004 495676 494604 495678
rect 530004 495676 530604 495678
rect 566004 495676 566604 495678
rect 590020 495676 590620 495678
rect -6696 495654 590620 495676
rect -6696 495418 -6514 495654
rect -6278 495418 26186 495654
rect 26422 495418 79610 495654
rect 79846 495418 314186 495654
rect 314422 495418 350186 495654
rect 350422 495418 386186 495654
rect 386422 495418 422186 495654
rect 422422 495418 458186 495654
rect 458422 495418 494186 495654
rect 494422 495418 530186 495654
rect 530422 495418 566186 495654
rect 566422 495418 590202 495654
rect 590438 495418 590620 495654
rect -6696 495334 590620 495418
rect -6696 495098 -6514 495334
rect -6278 495098 26186 495334
rect 26422 495098 79610 495334
rect 79846 495098 314186 495334
rect 314422 495098 350186 495334
rect 350422 495098 386186 495334
rect 386422 495098 422186 495334
rect 422422 495098 458186 495334
rect 458422 495098 494186 495334
rect 494422 495098 530186 495334
rect 530422 495098 566186 495334
rect 566422 495098 590202 495334
rect 590438 495098 590620 495334
rect -6696 495076 590620 495098
rect -6696 495074 -6096 495076
rect 26004 495074 26604 495076
rect 79568 495074 79888 495076
rect 314004 495074 314604 495076
rect 350004 495074 350604 495076
rect 386004 495074 386604 495076
rect 422004 495074 422604 495076
rect 458004 495074 458604 495076
rect 494004 495074 494604 495076
rect 530004 495074 530604 495076
rect 566004 495074 566604 495076
rect 590020 495074 590620 495076
rect -4816 492076 -4216 492078
rect 22404 492076 23004 492078
rect 79568 492076 79888 492078
rect 310404 492076 311004 492078
rect 346404 492076 347004 492078
rect 382404 492076 383004 492078
rect 418404 492076 419004 492078
rect 454404 492076 455004 492078
rect 490404 492076 491004 492078
rect 526404 492076 527004 492078
rect 562404 492076 563004 492078
rect 588140 492076 588740 492078
rect -4816 492054 588740 492076
rect -4816 491818 -4634 492054
rect -4398 491818 22586 492054
rect 22822 491818 79610 492054
rect 79846 491818 310586 492054
rect 310822 491818 346586 492054
rect 346822 491818 382586 492054
rect 382822 491818 418586 492054
rect 418822 491818 454586 492054
rect 454822 491818 490586 492054
rect 490822 491818 526586 492054
rect 526822 491818 562586 492054
rect 562822 491818 588322 492054
rect 588558 491818 588740 492054
rect -4816 491734 588740 491818
rect -4816 491498 -4634 491734
rect -4398 491498 22586 491734
rect 22822 491498 79610 491734
rect 79846 491498 310586 491734
rect 310822 491498 346586 491734
rect 346822 491498 382586 491734
rect 382822 491498 418586 491734
rect 418822 491498 454586 491734
rect 454822 491498 490586 491734
rect 490822 491498 526586 491734
rect 526822 491498 562586 491734
rect 562822 491498 588322 491734
rect 588558 491498 588740 491734
rect -4816 491476 588740 491498
rect -4816 491474 -4216 491476
rect 22404 491474 23004 491476
rect 79568 491474 79888 491476
rect 310404 491474 311004 491476
rect 346404 491474 347004 491476
rect 382404 491474 383004 491476
rect 418404 491474 419004 491476
rect 454404 491474 455004 491476
rect 490404 491474 491004 491476
rect 526404 491474 527004 491476
rect 562404 491474 563004 491476
rect 588140 491474 588740 491476
rect -2936 488476 -2336 488478
rect 18804 488476 19404 488478
rect 54804 488476 55404 488478
rect 79568 488476 79888 488478
rect 306804 488476 307404 488478
rect 342804 488476 343404 488478
rect 378804 488476 379404 488478
rect 414804 488476 415404 488478
rect 450804 488476 451404 488478
rect 486804 488476 487404 488478
rect 522804 488476 523404 488478
rect 558804 488476 559404 488478
rect 586260 488476 586860 488478
rect -2936 488454 586860 488476
rect -2936 488218 -2754 488454
rect -2518 488218 18986 488454
rect 19222 488218 54986 488454
rect 55222 488218 79610 488454
rect 79846 488218 306986 488454
rect 307222 488218 342986 488454
rect 343222 488218 378986 488454
rect 379222 488218 414986 488454
rect 415222 488218 450986 488454
rect 451222 488218 486986 488454
rect 487222 488218 522986 488454
rect 523222 488218 558986 488454
rect 559222 488218 586442 488454
rect 586678 488218 586860 488454
rect -2936 488134 586860 488218
rect -2936 487898 -2754 488134
rect -2518 487898 18986 488134
rect 19222 487898 54986 488134
rect 55222 487898 79610 488134
rect 79846 487898 306986 488134
rect 307222 487898 342986 488134
rect 343222 487898 378986 488134
rect 379222 487898 414986 488134
rect 415222 487898 450986 488134
rect 451222 487898 486986 488134
rect 487222 487898 522986 488134
rect 523222 487898 558986 488134
rect 559222 487898 586442 488134
rect 586678 487898 586860 488134
rect -2936 487876 586860 487898
rect -2936 487874 -2336 487876
rect 18804 487874 19404 487876
rect 54804 487874 55404 487876
rect 79568 487874 79888 487876
rect 306804 487874 307404 487876
rect 342804 487874 343404 487876
rect 378804 487874 379404 487876
rect 414804 487874 415404 487876
rect 450804 487874 451404 487876
rect 486804 487874 487404 487876
rect 522804 487874 523404 487876
rect 558804 487874 559404 487876
rect 586260 487874 586860 487876
rect -7636 481276 -7036 481278
rect 11604 481276 12204 481278
rect 47604 481276 48204 481278
rect 64208 481276 64528 481278
rect 299604 481276 300204 481278
rect 335604 481276 336204 481278
rect 371604 481276 372204 481278
rect 407604 481276 408204 481278
rect 443604 481276 444204 481278
rect 479604 481276 480204 481278
rect 515604 481276 516204 481278
rect 551604 481276 552204 481278
rect 590960 481276 591560 481278
rect -8576 481254 592500 481276
rect -8576 481018 -7454 481254
rect -7218 481018 11786 481254
rect 12022 481018 47786 481254
rect 48022 481018 64250 481254
rect 64486 481018 299786 481254
rect 300022 481018 335786 481254
rect 336022 481018 371786 481254
rect 372022 481018 407786 481254
rect 408022 481018 443786 481254
rect 444022 481018 479786 481254
rect 480022 481018 515786 481254
rect 516022 481018 551786 481254
rect 552022 481018 591142 481254
rect 591378 481018 592500 481254
rect -8576 480934 592500 481018
rect -8576 480698 -7454 480934
rect -7218 480698 11786 480934
rect 12022 480698 47786 480934
rect 48022 480698 64250 480934
rect 64486 480698 299786 480934
rect 300022 480698 335786 480934
rect 336022 480698 371786 480934
rect 372022 480698 407786 480934
rect 408022 480698 443786 480934
rect 444022 480698 479786 480934
rect 480022 480698 515786 480934
rect 516022 480698 551786 480934
rect 552022 480698 591142 480934
rect 591378 480698 592500 480934
rect -8576 480676 592500 480698
rect -7636 480674 -7036 480676
rect 11604 480674 12204 480676
rect 47604 480674 48204 480676
rect 64208 480674 64528 480676
rect 299604 480674 300204 480676
rect 335604 480674 336204 480676
rect 371604 480674 372204 480676
rect 407604 480674 408204 480676
rect 443604 480674 444204 480676
rect 479604 480674 480204 480676
rect 515604 480674 516204 480676
rect 551604 480674 552204 480676
rect 590960 480674 591560 480676
rect -5756 477676 -5156 477678
rect 8004 477676 8604 477678
rect 44004 477676 44604 477678
rect 64208 477676 64528 477678
rect 296004 477676 296604 477678
rect 332004 477676 332604 477678
rect 368004 477676 368604 477678
rect 404004 477676 404604 477678
rect 440004 477676 440604 477678
rect 476004 477676 476604 477678
rect 512004 477676 512604 477678
rect 548004 477676 548604 477678
rect 589080 477676 589680 477678
rect -6696 477654 590620 477676
rect -6696 477418 -5574 477654
rect -5338 477418 8186 477654
rect 8422 477418 44186 477654
rect 44422 477418 64250 477654
rect 64486 477418 296186 477654
rect 296422 477418 332186 477654
rect 332422 477418 368186 477654
rect 368422 477418 404186 477654
rect 404422 477418 440186 477654
rect 440422 477418 476186 477654
rect 476422 477418 512186 477654
rect 512422 477418 548186 477654
rect 548422 477418 589262 477654
rect 589498 477418 590620 477654
rect -6696 477334 590620 477418
rect -6696 477098 -5574 477334
rect -5338 477098 8186 477334
rect 8422 477098 44186 477334
rect 44422 477098 64250 477334
rect 64486 477098 296186 477334
rect 296422 477098 332186 477334
rect 332422 477098 368186 477334
rect 368422 477098 404186 477334
rect 404422 477098 440186 477334
rect 440422 477098 476186 477334
rect 476422 477098 512186 477334
rect 512422 477098 548186 477334
rect 548422 477098 589262 477334
rect 589498 477098 590620 477334
rect -6696 477076 590620 477098
rect -5756 477074 -5156 477076
rect 8004 477074 8604 477076
rect 44004 477074 44604 477076
rect 64208 477074 64528 477076
rect 296004 477074 296604 477076
rect 332004 477074 332604 477076
rect 368004 477074 368604 477076
rect 404004 477074 404604 477076
rect 440004 477074 440604 477076
rect 476004 477074 476604 477076
rect 512004 477074 512604 477076
rect 548004 477074 548604 477076
rect 589080 477074 589680 477076
rect -3876 474076 -3276 474078
rect 4404 474076 5004 474078
rect 40404 474076 41004 474078
rect 64208 474076 64528 474078
rect 292404 474076 293004 474078
rect 328404 474076 329004 474078
rect 364404 474076 365004 474078
rect 400404 474076 401004 474078
rect 436404 474076 437004 474078
rect 472404 474076 473004 474078
rect 508404 474076 509004 474078
rect 544404 474076 545004 474078
rect 580404 474076 581004 474078
rect 587200 474076 587800 474078
rect -4816 474054 588740 474076
rect -4816 473818 -3694 474054
rect -3458 473818 4586 474054
rect 4822 473818 40586 474054
rect 40822 473818 64250 474054
rect 64486 473818 292586 474054
rect 292822 473818 328586 474054
rect 328822 473818 364586 474054
rect 364822 473818 400586 474054
rect 400822 473818 436586 474054
rect 436822 473818 472586 474054
rect 472822 473818 508586 474054
rect 508822 473818 544586 474054
rect 544822 473818 580586 474054
rect 580822 473818 587382 474054
rect 587618 473818 588740 474054
rect -4816 473734 588740 473818
rect -4816 473498 -3694 473734
rect -3458 473498 4586 473734
rect 4822 473498 40586 473734
rect 40822 473498 64250 473734
rect 64486 473498 292586 473734
rect 292822 473498 328586 473734
rect 328822 473498 364586 473734
rect 364822 473498 400586 473734
rect 400822 473498 436586 473734
rect 436822 473498 472586 473734
rect 472822 473498 508586 473734
rect 508822 473498 544586 473734
rect 544822 473498 580586 473734
rect 580822 473498 587382 473734
rect 587618 473498 588740 473734
rect -4816 473476 588740 473498
rect -3876 473474 -3276 473476
rect 4404 473474 5004 473476
rect 40404 473474 41004 473476
rect 64208 473474 64528 473476
rect 292404 473474 293004 473476
rect 328404 473474 329004 473476
rect 364404 473474 365004 473476
rect 400404 473474 401004 473476
rect 436404 473474 437004 473476
rect 472404 473474 473004 473476
rect 508404 473474 509004 473476
rect 544404 473474 545004 473476
rect 580404 473474 581004 473476
rect 587200 473474 587800 473476
rect -1996 470476 -1396 470478
rect 804 470476 1404 470478
rect 36804 470476 37404 470478
rect 64208 470476 64528 470478
rect 288804 470476 289404 470478
rect 324804 470476 325404 470478
rect 360804 470476 361404 470478
rect 396804 470476 397404 470478
rect 432804 470476 433404 470478
rect 468804 470476 469404 470478
rect 504804 470476 505404 470478
rect 540804 470476 541404 470478
rect 576804 470476 577404 470478
rect 585320 470476 585920 470478
rect -2936 470454 586860 470476
rect -2936 470218 -1814 470454
rect -1578 470218 986 470454
rect 1222 470218 36986 470454
rect 37222 470218 64250 470454
rect 64486 470218 288986 470454
rect 289222 470218 324986 470454
rect 325222 470218 360986 470454
rect 361222 470218 396986 470454
rect 397222 470218 432986 470454
rect 433222 470218 468986 470454
rect 469222 470218 504986 470454
rect 505222 470218 540986 470454
rect 541222 470218 576986 470454
rect 577222 470218 585502 470454
rect 585738 470218 586860 470454
rect -2936 470134 586860 470218
rect -2936 469898 -1814 470134
rect -1578 469898 986 470134
rect 1222 469898 36986 470134
rect 37222 469898 64250 470134
rect 64486 469898 288986 470134
rect 289222 469898 324986 470134
rect 325222 469898 360986 470134
rect 361222 469898 396986 470134
rect 397222 469898 432986 470134
rect 433222 469898 468986 470134
rect 469222 469898 504986 470134
rect 505222 469898 540986 470134
rect 541222 469898 576986 470134
rect 577222 469898 585502 470134
rect 585738 469898 586860 470134
rect -2936 469876 586860 469898
rect -1996 469874 -1396 469876
rect 804 469874 1404 469876
rect 36804 469874 37404 469876
rect 64208 469874 64528 469876
rect 288804 469874 289404 469876
rect 324804 469874 325404 469876
rect 360804 469874 361404 469876
rect 396804 469874 397404 469876
rect 432804 469874 433404 469876
rect 468804 469874 469404 469876
rect 504804 469874 505404 469876
rect 540804 469874 541404 469876
rect 576804 469874 577404 469876
rect 585320 469874 585920 469876
rect -8576 463276 -7976 463278
rect 29604 463276 30204 463278
rect 79568 463276 79888 463278
rect 317604 463276 318204 463278
rect 353604 463276 354204 463278
rect 389604 463276 390204 463278
rect 425604 463276 426204 463278
rect 461604 463276 462204 463278
rect 497604 463276 498204 463278
rect 533604 463276 534204 463278
rect 569604 463276 570204 463278
rect 591900 463276 592500 463278
rect -8576 463254 592500 463276
rect -8576 463018 -8394 463254
rect -8158 463018 29786 463254
rect 30022 463018 79610 463254
rect 79846 463018 317786 463254
rect 318022 463018 353786 463254
rect 354022 463018 389786 463254
rect 390022 463018 425786 463254
rect 426022 463018 461786 463254
rect 462022 463018 497786 463254
rect 498022 463018 533786 463254
rect 534022 463018 569786 463254
rect 570022 463018 592082 463254
rect 592318 463018 592500 463254
rect -8576 462934 592500 463018
rect -8576 462698 -8394 462934
rect -8158 462698 29786 462934
rect 30022 462698 79610 462934
rect 79846 462698 317786 462934
rect 318022 462698 353786 462934
rect 354022 462698 389786 462934
rect 390022 462698 425786 462934
rect 426022 462698 461786 462934
rect 462022 462698 497786 462934
rect 498022 462698 533786 462934
rect 534022 462698 569786 462934
rect 570022 462698 592082 462934
rect 592318 462698 592500 462934
rect -8576 462676 592500 462698
rect -8576 462674 -7976 462676
rect 29604 462674 30204 462676
rect 79568 462674 79888 462676
rect 317604 462674 318204 462676
rect 353604 462674 354204 462676
rect 389604 462674 390204 462676
rect 425604 462674 426204 462676
rect 461604 462674 462204 462676
rect 497604 462674 498204 462676
rect 533604 462674 534204 462676
rect 569604 462674 570204 462676
rect 591900 462674 592500 462676
rect -6696 459676 -6096 459678
rect 26004 459676 26604 459678
rect 79568 459676 79888 459678
rect 314004 459676 314604 459678
rect 350004 459676 350604 459678
rect 386004 459676 386604 459678
rect 422004 459676 422604 459678
rect 458004 459676 458604 459678
rect 494004 459676 494604 459678
rect 530004 459676 530604 459678
rect 566004 459676 566604 459678
rect 590020 459676 590620 459678
rect -6696 459654 590620 459676
rect -6696 459418 -6514 459654
rect -6278 459418 26186 459654
rect 26422 459418 79610 459654
rect 79846 459418 314186 459654
rect 314422 459418 350186 459654
rect 350422 459418 386186 459654
rect 386422 459418 422186 459654
rect 422422 459418 458186 459654
rect 458422 459418 494186 459654
rect 494422 459418 530186 459654
rect 530422 459418 566186 459654
rect 566422 459418 590202 459654
rect 590438 459418 590620 459654
rect -6696 459334 590620 459418
rect -6696 459098 -6514 459334
rect -6278 459098 26186 459334
rect 26422 459098 79610 459334
rect 79846 459098 314186 459334
rect 314422 459098 350186 459334
rect 350422 459098 386186 459334
rect 386422 459098 422186 459334
rect 422422 459098 458186 459334
rect 458422 459098 494186 459334
rect 494422 459098 530186 459334
rect 530422 459098 566186 459334
rect 566422 459098 590202 459334
rect 590438 459098 590620 459334
rect -6696 459076 590620 459098
rect -6696 459074 -6096 459076
rect 26004 459074 26604 459076
rect 79568 459074 79888 459076
rect 314004 459074 314604 459076
rect 350004 459074 350604 459076
rect 386004 459074 386604 459076
rect 422004 459074 422604 459076
rect 458004 459074 458604 459076
rect 494004 459074 494604 459076
rect 530004 459074 530604 459076
rect 566004 459074 566604 459076
rect 590020 459074 590620 459076
rect -4816 456076 -4216 456078
rect 22404 456076 23004 456078
rect 79568 456076 79888 456078
rect 310404 456076 311004 456078
rect 346404 456076 347004 456078
rect 382404 456076 383004 456078
rect 418404 456076 419004 456078
rect 454404 456076 455004 456078
rect 490404 456076 491004 456078
rect 526404 456076 527004 456078
rect 562404 456076 563004 456078
rect 588140 456076 588740 456078
rect -4816 456054 588740 456076
rect -4816 455818 -4634 456054
rect -4398 455818 22586 456054
rect 22822 455818 79610 456054
rect 79846 455818 310586 456054
rect 310822 455818 346586 456054
rect 346822 455818 382586 456054
rect 382822 455818 418586 456054
rect 418822 455818 454586 456054
rect 454822 455818 490586 456054
rect 490822 455818 526586 456054
rect 526822 455818 562586 456054
rect 562822 455818 588322 456054
rect 588558 455818 588740 456054
rect -4816 455734 588740 455818
rect -4816 455498 -4634 455734
rect -4398 455498 22586 455734
rect 22822 455498 79610 455734
rect 79846 455498 310586 455734
rect 310822 455498 346586 455734
rect 346822 455498 382586 455734
rect 382822 455498 418586 455734
rect 418822 455498 454586 455734
rect 454822 455498 490586 455734
rect 490822 455498 526586 455734
rect 526822 455498 562586 455734
rect 562822 455498 588322 455734
rect 588558 455498 588740 455734
rect -4816 455476 588740 455498
rect -4816 455474 -4216 455476
rect 22404 455474 23004 455476
rect 79568 455474 79888 455476
rect 310404 455474 311004 455476
rect 346404 455474 347004 455476
rect 382404 455474 383004 455476
rect 418404 455474 419004 455476
rect 454404 455474 455004 455476
rect 490404 455474 491004 455476
rect 526404 455474 527004 455476
rect 562404 455474 563004 455476
rect 588140 455474 588740 455476
rect -2936 452476 -2336 452478
rect 18804 452476 19404 452478
rect 54804 452476 55404 452478
rect 79568 452476 79888 452478
rect 306804 452476 307404 452478
rect 342804 452476 343404 452478
rect 378804 452476 379404 452478
rect 414804 452476 415404 452478
rect 450804 452476 451404 452478
rect 486804 452476 487404 452478
rect 522804 452476 523404 452478
rect 558804 452476 559404 452478
rect 586260 452476 586860 452478
rect -2936 452454 586860 452476
rect -2936 452218 -2754 452454
rect -2518 452218 18986 452454
rect 19222 452218 54986 452454
rect 55222 452218 79610 452454
rect 79846 452218 306986 452454
rect 307222 452218 342986 452454
rect 343222 452218 378986 452454
rect 379222 452218 414986 452454
rect 415222 452218 450986 452454
rect 451222 452218 486986 452454
rect 487222 452218 522986 452454
rect 523222 452218 558986 452454
rect 559222 452218 586442 452454
rect 586678 452218 586860 452454
rect -2936 452134 586860 452218
rect -2936 451898 -2754 452134
rect -2518 451898 18986 452134
rect 19222 451898 54986 452134
rect 55222 451898 79610 452134
rect 79846 451898 306986 452134
rect 307222 451898 342986 452134
rect 343222 451898 378986 452134
rect 379222 451898 414986 452134
rect 415222 451898 450986 452134
rect 451222 451898 486986 452134
rect 487222 451898 522986 452134
rect 523222 451898 558986 452134
rect 559222 451898 586442 452134
rect 586678 451898 586860 452134
rect -2936 451876 586860 451898
rect -2936 451874 -2336 451876
rect 18804 451874 19404 451876
rect 54804 451874 55404 451876
rect 79568 451874 79888 451876
rect 306804 451874 307404 451876
rect 342804 451874 343404 451876
rect 378804 451874 379404 451876
rect 414804 451874 415404 451876
rect 450804 451874 451404 451876
rect 486804 451874 487404 451876
rect 522804 451874 523404 451876
rect 558804 451874 559404 451876
rect 586260 451874 586860 451876
rect -7636 445276 -7036 445278
rect 11604 445276 12204 445278
rect 47604 445276 48204 445278
rect 64208 445276 64528 445278
rect 299604 445276 300204 445278
rect 335604 445276 336204 445278
rect 371604 445276 372204 445278
rect 407604 445276 408204 445278
rect 443604 445276 444204 445278
rect 479604 445276 480204 445278
rect 515604 445276 516204 445278
rect 551604 445276 552204 445278
rect 590960 445276 591560 445278
rect -8576 445254 592500 445276
rect -8576 445018 -7454 445254
rect -7218 445018 11786 445254
rect 12022 445018 47786 445254
rect 48022 445018 64250 445254
rect 64486 445018 299786 445254
rect 300022 445018 335786 445254
rect 336022 445018 371786 445254
rect 372022 445018 407786 445254
rect 408022 445018 443786 445254
rect 444022 445018 479786 445254
rect 480022 445018 515786 445254
rect 516022 445018 551786 445254
rect 552022 445018 591142 445254
rect 591378 445018 592500 445254
rect -8576 444934 592500 445018
rect -8576 444698 -7454 444934
rect -7218 444698 11786 444934
rect 12022 444698 47786 444934
rect 48022 444698 64250 444934
rect 64486 444698 299786 444934
rect 300022 444698 335786 444934
rect 336022 444698 371786 444934
rect 372022 444698 407786 444934
rect 408022 444698 443786 444934
rect 444022 444698 479786 444934
rect 480022 444698 515786 444934
rect 516022 444698 551786 444934
rect 552022 444698 591142 444934
rect 591378 444698 592500 444934
rect -8576 444676 592500 444698
rect -7636 444674 -7036 444676
rect 11604 444674 12204 444676
rect 47604 444674 48204 444676
rect 64208 444674 64528 444676
rect 299604 444674 300204 444676
rect 335604 444674 336204 444676
rect 371604 444674 372204 444676
rect 407604 444674 408204 444676
rect 443604 444674 444204 444676
rect 479604 444674 480204 444676
rect 515604 444674 516204 444676
rect 551604 444674 552204 444676
rect 590960 444674 591560 444676
rect -5756 441676 -5156 441678
rect 8004 441676 8604 441678
rect 44004 441676 44604 441678
rect 64208 441676 64528 441678
rect 296004 441676 296604 441678
rect 332004 441676 332604 441678
rect 368004 441676 368604 441678
rect 404004 441676 404604 441678
rect 440004 441676 440604 441678
rect 476004 441676 476604 441678
rect 512004 441676 512604 441678
rect 548004 441676 548604 441678
rect 589080 441676 589680 441678
rect -6696 441654 590620 441676
rect -6696 441418 -5574 441654
rect -5338 441418 8186 441654
rect 8422 441418 44186 441654
rect 44422 441418 64250 441654
rect 64486 441418 296186 441654
rect 296422 441418 332186 441654
rect 332422 441418 368186 441654
rect 368422 441418 404186 441654
rect 404422 441418 440186 441654
rect 440422 441418 476186 441654
rect 476422 441418 512186 441654
rect 512422 441418 548186 441654
rect 548422 441418 589262 441654
rect 589498 441418 590620 441654
rect -6696 441334 590620 441418
rect -6696 441098 -5574 441334
rect -5338 441098 8186 441334
rect 8422 441098 44186 441334
rect 44422 441098 64250 441334
rect 64486 441098 296186 441334
rect 296422 441098 332186 441334
rect 332422 441098 368186 441334
rect 368422 441098 404186 441334
rect 404422 441098 440186 441334
rect 440422 441098 476186 441334
rect 476422 441098 512186 441334
rect 512422 441098 548186 441334
rect 548422 441098 589262 441334
rect 589498 441098 590620 441334
rect -6696 441076 590620 441098
rect -5756 441074 -5156 441076
rect 8004 441074 8604 441076
rect 44004 441074 44604 441076
rect 64208 441074 64528 441076
rect 296004 441074 296604 441076
rect 332004 441074 332604 441076
rect 368004 441074 368604 441076
rect 404004 441074 404604 441076
rect 440004 441074 440604 441076
rect 476004 441074 476604 441076
rect 512004 441074 512604 441076
rect 548004 441074 548604 441076
rect 589080 441074 589680 441076
rect -3876 438076 -3276 438078
rect 4404 438076 5004 438078
rect 40404 438076 41004 438078
rect 64208 438076 64528 438078
rect 292404 438076 293004 438078
rect 328404 438076 329004 438078
rect 364404 438076 365004 438078
rect 400404 438076 401004 438078
rect 436404 438076 437004 438078
rect 472404 438076 473004 438078
rect 508404 438076 509004 438078
rect 544404 438076 545004 438078
rect 580404 438076 581004 438078
rect 587200 438076 587800 438078
rect -4816 438054 588740 438076
rect -4816 437818 -3694 438054
rect -3458 437818 4586 438054
rect 4822 437818 40586 438054
rect 40822 437818 64250 438054
rect 64486 437818 292586 438054
rect 292822 437818 328586 438054
rect 328822 437818 364586 438054
rect 364822 437818 400586 438054
rect 400822 437818 436586 438054
rect 436822 437818 472586 438054
rect 472822 437818 508586 438054
rect 508822 437818 544586 438054
rect 544822 437818 580586 438054
rect 580822 437818 587382 438054
rect 587618 437818 588740 438054
rect -4816 437734 588740 437818
rect -4816 437498 -3694 437734
rect -3458 437498 4586 437734
rect 4822 437498 40586 437734
rect 40822 437498 64250 437734
rect 64486 437498 292586 437734
rect 292822 437498 328586 437734
rect 328822 437498 364586 437734
rect 364822 437498 400586 437734
rect 400822 437498 436586 437734
rect 436822 437498 472586 437734
rect 472822 437498 508586 437734
rect 508822 437498 544586 437734
rect 544822 437498 580586 437734
rect 580822 437498 587382 437734
rect 587618 437498 588740 437734
rect -4816 437476 588740 437498
rect -3876 437474 -3276 437476
rect 4404 437474 5004 437476
rect 40404 437474 41004 437476
rect 64208 437474 64528 437476
rect 292404 437474 293004 437476
rect 328404 437474 329004 437476
rect 364404 437474 365004 437476
rect 400404 437474 401004 437476
rect 436404 437474 437004 437476
rect 472404 437474 473004 437476
rect 508404 437474 509004 437476
rect 544404 437474 545004 437476
rect 580404 437474 581004 437476
rect 587200 437474 587800 437476
rect -1996 434476 -1396 434478
rect 804 434476 1404 434478
rect 36804 434476 37404 434478
rect 64208 434476 64528 434478
rect 288804 434476 289404 434478
rect 324804 434476 325404 434478
rect 360804 434476 361404 434478
rect 396804 434476 397404 434478
rect 432804 434476 433404 434478
rect 468804 434476 469404 434478
rect 504804 434476 505404 434478
rect 540804 434476 541404 434478
rect 576804 434476 577404 434478
rect 585320 434476 585920 434478
rect -2936 434454 586860 434476
rect -2936 434218 -1814 434454
rect -1578 434218 986 434454
rect 1222 434218 36986 434454
rect 37222 434218 64250 434454
rect 64486 434218 288986 434454
rect 289222 434218 324986 434454
rect 325222 434218 360986 434454
rect 361222 434218 396986 434454
rect 397222 434218 432986 434454
rect 433222 434218 468986 434454
rect 469222 434218 504986 434454
rect 505222 434218 540986 434454
rect 541222 434218 576986 434454
rect 577222 434218 585502 434454
rect 585738 434218 586860 434454
rect -2936 434134 586860 434218
rect -2936 433898 -1814 434134
rect -1578 433898 986 434134
rect 1222 433898 36986 434134
rect 37222 433898 64250 434134
rect 64486 433898 288986 434134
rect 289222 433898 324986 434134
rect 325222 433898 360986 434134
rect 361222 433898 396986 434134
rect 397222 433898 432986 434134
rect 433222 433898 468986 434134
rect 469222 433898 504986 434134
rect 505222 433898 540986 434134
rect 541222 433898 576986 434134
rect 577222 433898 585502 434134
rect 585738 433898 586860 434134
rect -2936 433876 586860 433898
rect -1996 433874 -1396 433876
rect 804 433874 1404 433876
rect 36804 433874 37404 433876
rect 64208 433874 64528 433876
rect 288804 433874 289404 433876
rect 324804 433874 325404 433876
rect 360804 433874 361404 433876
rect 396804 433874 397404 433876
rect 432804 433874 433404 433876
rect 468804 433874 469404 433876
rect 504804 433874 505404 433876
rect 540804 433874 541404 433876
rect 576804 433874 577404 433876
rect 585320 433874 585920 433876
rect -8576 427276 -7976 427278
rect 29604 427276 30204 427278
rect 79568 427276 79888 427278
rect 317604 427276 318204 427278
rect 353604 427276 354204 427278
rect 389604 427276 390204 427278
rect 425604 427276 426204 427278
rect 461604 427276 462204 427278
rect 497604 427276 498204 427278
rect 533604 427276 534204 427278
rect 569604 427276 570204 427278
rect 591900 427276 592500 427278
rect -8576 427254 592500 427276
rect -8576 427018 -8394 427254
rect -8158 427018 29786 427254
rect 30022 427018 79610 427254
rect 79846 427018 317786 427254
rect 318022 427018 353786 427254
rect 354022 427018 389786 427254
rect 390022 427018 425786 427254
rect 426022 427018 461786 427254
rect 462022 427018 497786 427254
rect 498022 427018 533786 427254
rect 534022 427018 569786 427254
rect 570022 427018 592082 427254
rect 592318 427018 592500 427254
rect -8576 426934 592500 427018
rect -8576 426698 -8394 426934
rect -8158 426698 29786 426934
rect 30022 426698 79610 426934
rect 79846 426698 317786 426934
rect 318022 426698 353786 426934
rect 354022 426698 389786 426934
rect 390022 426698 425786 426934
rect 426022 426698 461786 426934
rect 462022 426698 497786 426934
rect 498022 426698 533786 426934
rect 534022 426698 569786 426934
rect 570022 426698 592082 426934
rect 592318 426698 592500 426934
rect -8576 426676 592500 426698
rect -8576 426674 -7976 426676
rect 29604 426674 30204 426676
rect 79568 426674 79888 426676
rect 317604 426674 318204 426676
rect 353604 426674 354204 426676
rect 389604 426674 390204 426676
rect 425604 426674 426204 426676
rect 461604 426674 462204 426676
rect 497604 426674 498204 426676
rect 533604 426674 534204 426676
rect 569604 426674 570204 426676
rect 591900 426674 592500 426676
rect -6696 423676 -6096 423678
rect 26004 423676 26604 423678
rect 79568 423676 79888 423678
rect 314004 423676 314604 423678
rect 350004 423676 350604 423678
rect 386004 423676 386604 423678
rect 422004 423676 422604 423678
rect 458004 423676 458604 423678
rect 494004 423676 494604 423678
rect 530004 423676 530604 423678
rect 566004 423676 566604 423678
rect 590020 423676 590620 423678
rect -6696 423654 590620 423676
rect -6696 423418 -6514 423654
rect -6278 423418 26186 423654
rect 26422 423418 79610 423654
rect 79846 423418 314186 423654
rect 314422 423418 350186 423654
rect 350422 423418 386186 423654
rect 386422 423418 422186 423654
rect 422422 423418 458186 423654
rect 458422 423418 494186 423654
rect 494422 423418 530186 423654
rect 530422 423418 566186 423654
rect 566422 423418 590202 423654
rect 590438 423418 590620 423654
rect -6696 423334 590620 423418
rect -6696 423098 -6514 423334
rect -6278 423098 26186 423334
rect 26422 423098 79610 423334
rect 79846 423098 314186 423334
rect 314422 423098 350186 423334
rect 350422 423098 386186 423334
rect 386422 423098 422186 423334
rect 422422 423098 458186 423334
rect 458422 423098 494186 423334
rect 494422 423098 530186 423334
rect 530422 423098 566186 423334
rect 566422 423098 590202 423334
rect 590438 423098 590620 423334
rect -6696 423076 590620 423098
rect -6696 423074 -6096 423076
rect 26004 423074 26604 423076
rect 79568 423074 79888 423076
rect 314004 423074 314604 423076
rect 350004 423074 350604 423076
rect 386004 423074 386604 423076
rect 422004 423074 422604 423076
rect 458004 423074 458604 423076
rect 494004 423074 494604 423076
rect 530004 423074 530604 423076
rect 566004 423074 566604 423076
rect 590020 423074 590620 423076
rect -4816 420076 -4216 420078
rect 22404 420076 23004 420078
rect 79568 420076 79888 420078
rect 310404 420076 311004 420078
rect 346404 420076 347004 420078
rect 382404 420076 383004 420078
rect 418404 420076 419004 420078
rect 454404 420076 455004 420078
rect 490404 420076 491004 420078
rect 526404 420076 527004 420078
rect 562404 420076 563004 420078
rect 588140 420076 588740 420078
rect -4816 420054 588740 420076
rect -4816 419818 -4634 420054
rect -4398 419818 22586 420054
rect 22822 419818 79610 420054
rect 79846 419818 310586 420054
rect 310822 419818 346586 420054
rect 346822 419818 382586 420054
rect 382822 419818 418586 420054
rect 418822 419818 454586 420054
rect 454822 419818 490586 420054
rect 490822 419818 526586 420054
rect 526822 419818 562586 420054
rect 562822 419818 588322 420054
rect 588558 419818 588740 420054
rect -4816 419734 588740 419818
rect -4816 419498 -4634 419734
rect -4398 419498 22586 419734
rect 22822 419498 79610 419734
rect 79846 419498 310586 419734
rect 310822 419498 346586 419734
rect 346822 419498 382586 419734
rect 382822 419498 418586 419734
rect 418822 419498 454586 419734
rect 454822 419498 490586 419734
rect 490822 419498 526586 419734
rect 526822 419498 562586 419734
rect 562822 419498 588322 419734
rect 588558 419498 588740 419734
rect -4816 419476 588740 419498
rect -4816 419474 -4216 419476
rect 22404 419474 23004 419476
rect 79568 419474 79888 419476
rect 310404 419474 311004 419476
rect 346404 419474 347004 419476
rect 382404 419474 383004 419476
rect 418404 419474 419004 419476
rect 454404 419474 455004 419476
rect 490404 419474 491004 419476
rect 526404 419474 527004 419476
rect 562404 419474 563004 419476
rect 588140 419474 588740 419476
rect -2936 416476 -2336 416478
rect 18804 416476 19404 416478
rect 54804 416476 55404 416478
rect 79568 416476 79888 416478
rect 306804 416476 307404 416478
rect 342804 416476 343404 416478
rect 378804 416476 379404 416478
rect 414804 416476 415404 416478
rect 450804 416476 451404 416478
rect 486804 416476 487404 416478
rect 522804 416476 523404 416478
rect 558804 416476 559404 416478
rect 586260 416476 586860 416478
rect -2936 416454 586860 416476
rect -2936 416218 -2754 416454
rect -2518 416218 18986 416454
rect 19222 416218 54986 416454
rect 55222 416218 79610 416454
rect 79846 416218 306986 416454
rect 307222 416218 342986 416454
rect 343222 416218 378986 416454
rect 379222 416218 414986 416454
rect 415222 416218 450986 416454
rect 451222 416218 486986 416454
rect 487222 416218 522986 416454
rect 523222 416218 558986 416454
rect 559222 416218 586442 416454
rect 586678 416218 586860 416454
rect -2936 416134 586860 416218
rect -2936 415898 -2754 416134
rect -2518 415898 18986 416134
rect 19222 415898 54986 416134
rect 55222 415898 79610 416134
rect 79846 415898 306986 416134
rect 307222 415898 342986 416134
rect 343222 415898 378986 416134
rect 379222 415898 414986 416134
rect 415222 415898 450986 416134
rect 451222 415898 486986 416134
rect 487222 415898 522986 416134
rect 523222 415898 558986 416134
rect 559222 415898 586442 416134
rect 586678 415898 586860 416134
rect -2936 415876 586860 415898
rect -2936 415874 -2336 415876
rect 18804 415874 19404 415876
rect 54804 415874 55404 415876
rect 79568 415874 79888 415876
rect 306804 415874 307404 415876
rect 342804 415874 343404 415876
rect 378804 415874 379404 415876
rect 414804 415874 415404 415876
rect 450804 415874 451404 415876
rect 486804 415874 487404 415876
rect 522804 415874 523404 415876
rect 558804 415874 559404 415876
rect 586260 415874 586860 415876
rect -7636 409276 -7036 409278
rect 11604 409276 12204 409278
rect 47604 409276 48204 409278
rect 64208 409276 64528 409278
rect 299604 409276 300204 409278
rect 335604 409276 336204 409278
rect 340482 409276 340802 409278
rect 443604 409276 444204 409278
rect 479604 409276 480204 409278
rect 515604 409276 516204 409278
rect 551604 409276 552204 409278
rect 590960 409276 591560 409278
rect -8576 409254 592500 409276
rect -8576 409018 -7454 409254
rect -7218 409018 11786 409254
rect 12022 409018 47786 409254
rect 48022 409018 64250 409254
rect 64486 409018 299786 409254
rect 300022 409018 335786 409254
rect 336022 409018 340524 409254
rect 340760 409018 443786 409254
rect 444022 409018 479786 409254
rect 480022 409018 515786 409254
rect 516022 409018 551786 409254
rect 552022 409018 591142 409254
rect 591378 409018 592500 409254
rect -8576 408934 592500 409018
rect -8576 408698 -7454 408934
rect -7218 408698 11786 408934
rect 12022 408698 47786 408934
rect 48022 408698 64250 408934
rect 64486 408698 299786 408934
rect 300022 408698 335786 408934
rect 336022 408698 340524 408934
rect 340760 408698 443786 408934
rect 444022 408698 479786 408934
rect 480022 408698 515786 408934
rect 516022 408698 551786 408934
rect 552022 408698 591142 408934
rect 591378 408698 592500 408934
rect -8576 408676 592500 408698
rect -7636 408674 -7036 408676
rect 11604 408674 12204 408676
rect 47604 408674 48204 408676
rect 64208 408674 64528 408676
rect 299604 408674 300204 408676
rect 335604 408674 336204 408676
rect 340482 408674 340802 408676
rect 443604 408674 444204 408676
rect 479604 408674 480204 408676
rect 515604 408674 516204 408676
rect 551604 408674 552204 408676
rect 590960 408674 591560 408676
rect -5756 405676 -5156 405678
rect 8004 405676 8604 405678
rect 44004 405676 44604 405678
rect 64208 405676 64528 405678
rect 296004 405676 296604 405678
rect 332004 405676 332604 405678
rect 340482 405676 340802 405678
rect 440004 405676 440604 405678
rect 476004 405676 476604 405678
rect 512004 405676 512604 405678
rect 548004 405676 548604 405678
rect 589080 405676 589680 405678
rect -6696 405654 590620 405676
rect -6696 405418 -5574 405654
rect -5338 405418 8186 405654
rect 8422 405418 44186 405654
rect 44422 405418 64250 405654
rect 64486 405418 296186 405654
rect 296422 405418 332186 405654
rect 332422 405418 340524 405654
rect 340760 405418 440186 405654
rect 440422 405418 476186 405654
rect 476422 405418 512186 405654
rect 512422 405418 548186 405654
rect 548422 405418 589262 405654
rect 589498 405418 590620 405654
rect -6696 405334 590620 405418
rect -6696 405098 -5574 405334
rect -5338 405098 8186 405334
rect 8422 405098 44186 405334
rect 44422 405098 64250 405334
rect 64486 405098 296186 405334
rect 296422 405098 332186 405334
rect 332422 405098 340524 405334
rect 340760 405098 440186 405334
rect 440422 405098 476186 405334
rect 476422 405098 512186 405334
rect 512422 405098 548186 405334
rect 548422 405098 589262 405334
rect 589498 405098 590620 405334
rect -6696 405076 590620 405098
rect -5756 405074 -5156 405076
rect 8004 405074 8604 405076
rect 44004 405074 44604 405076
rect 64208 405074 64528 405076
rect 296004 405074 296604 405076
rect 332004 405074 332604 405076
rect 340482 405074 340802 405076
rect 440004 405074 440604 405076
rect 476004 405074 476604 405076
rect 512004 405074 512604 405076
rect 548004 405074 548604 405076
rect 589080 405074 589680 405076
rect -3876 402076 -3276 402078
rect 4404 402076 5004 402078
rect 40404 402076 41004 402078
rect 64208 402076 64528 402078
rect 292404 402076 293004 402078
rect 328404 402076 329004 402078
rect 340482 402076 340802 402078
rect 436404 402076 437004 402078
rect 472404 402076 473004 402078
rect 508404 402076 509004 402078
rect 544404 402076 545004 402078
rect 580404 402076 581004 402078
rect 587200 402076 587800 402078
rect -4816 402054 588740 402076
rect -4816 401818 -3694 402054
rect -3458 401818 4586 402054
rect 4822 401818 40586 402054
rect 40822 401818 64250 402054
rect 64486 401818 292586 402054
rect 292822 401818 328586 402054
rect 328822 401818 340524 402054
rect 340760 401818 436586 402054
rect 436822 401818 472586 402054
rect 472822 401818 508586 402054
rect 508822 401818 544586 402054
rect 544822 401818 580586 402054
rect 580822 401818 587382 402054
rect 587618 401818 588740 402054
rect -4816 401734 588740 401818
rect -4816 401498 -3694 401734
rect -3458 401498 4586 401734
rect 4822 401498 40586 401734
rect 40822 401498 64250 401734
rect 64486 401498 292586 401734
rect 292822 401498 328586 401734
rect 328822 401498 340524 401734
rect 340760 401498 436586 401734
rect 436822 401498 472586 401734
rect 472822 401498 508586 401734
rect 508822 401498 544586 401734
rect 544822 401498 580586 401734
rect 580822 401498 587382 401734
rect 587618 401498 588740 401734
rect -4816 401476 588740 401498
rect -3876 401474 -3276 401476
rect 4404 401474 5004 401476
rect 40404 401474 41004 401476
rect 64208 401474 64528 401476
rect 292404 401474 293004 401476
rect 328404 401474 329004 401476
rect 340482 401474 340802 401476
rect 436404 401474 437004 401476
rect 472404 401474 473004 401476
rect 508404 401474 509004 401476
rect 544404 401474 545004 401476
rect 580404 401474 581004 401476
rect 587200 401474 587800 401476
rect -1996 398476 -1396 398478
rect 804 398476 1404 398478
rect 36804 398476 37404 398478
rect 64208 398476 64528 398478
rect 288804 398476 289404 398478
rect 324804 398476 325404 398478
rect 340482 398476 340802 398478
rect 432804 398476 433404 398478
rect 468804 398476 469404 398478
rect 504804 398476 505404 398478
rect 540804 398476 541404 398478
rect 576804 398476 577404 398478
rect 585320 398476 585920 398478
rect -2936 398454 586860 398476
rect -2936 398218 -1814 398454
rect -1578 398218 986 398454
rect 1222 398218 36986 398454
rect 37222 398218 64250 398454
rect 64486 398218 288986 398454
rect 289222 398218 324986 398454
rect 325222 398218 340524 398454
rect 340760 398218 432986 398454
rect 433222 398218 468986 398454
rect 469222 398218 504986 398454
rect 505222 398218 540986 398454
rect 541222 398218 576986 398454
rect 577222 398218 585502 398454
rect 585738 398218 586860 398454
rect -2936 398134 586860 398218
rect -2936 397898 -1814 398134
rect -1578 397898 986 398134
rect 1222 397898 36986 398134
rect 37222 397898 64250 398134
rect 64486 397898 288986 398134
rect 289222 397898 324986 398134
rect 325222 397898 340524 398134
rect 340760 397898 432986 398134
rect 433222 397898 468986 398134
rect 469222 397898 504986 398134
rect 505222 397898 540986 398134
rect 541222 397898 576986 398134
rect 577222 397898 585502 398134
rect 585738 397898 586860 398134
rect -2936 397876 586860 397898
rect -1996 397874 -1396 397876
rect 804 397874 1404 397876
rect 36804 397874 37404 397876
rect 64208 397874 64528 397876
rect 288804 397874 289404 397876
rect 324804 397874 325404 397876
rect 340482 397874 340802 397876
rect 432804 397874 433404 397876
rect 468804 397874 469404 397876
rect 504804 397874 505404 397876
rect 540804 397874 541404 397876
rect 576804 397874 577404 397876
rect 585320 397874 585920 397876
rect -8576 391276 -7976 391278
rect 29604 391276 30204 391278
rect 79568 391276 79888 391278
rect 317604 391276 318204 391278
rect 340034 391276 340358 391278
rect 425604 391276 426204 391278
rect 461604 391276 462204 391278
rect 497604 391276 498204 391278
rect 533604 391276 534204 391278
rect 569604 391276 570204 391278
rect 591900 391276 592500 391278
rect -8576 391254 592500 391276
rect -8576 391018 -8394 391254
rect -8158 391018 29786 391254
rect 30022 391018 79610 391254
rect 79846 391018 317786 391254
rect 318022 391018 340078 391254
rect 340314 391018 425786 391254
rect 426022 391018 461786 391254
rect 462022 391018 497786 391254
rect 498022 391018 533786 391254
rect 534022 391018 569786 391254
rect 570022 391018 592082 391254
rect 592318 391018 592500 391254
rect -8576 390934 592500 391018
rect -8576 390698 -8394 390934
rect -8158 390698 29786 390934
rect 30022 390698 79610 390934
rect 79846 390698 317786 390934
rect 318022 390698 340078 390934
rect 340314 390698 425786 390934
rect 426022 390698 461786 390934
rect 462022 390698 497786 390934
rect 498022 390698 533786 390934
rect 534022 390698 569786 390934
rect 570022 390698 592082 390934
rect 592318 390698 592500 390934
rect -8576 390676 592500 390698
rect -8576 390674 -7976 390676
rect 29604 390674 30204 390676
rect 79568 390674 79888 390676
rect 317604 390674 318204 390676
rect 340034 390674 340358 390676
rect 425604 390674 426204 390676
rect 461604 390674 462204 390676
rect 497604 390674 498204 390676
rect 533604 390674 534204 390676
rect 569604 390674 570204 390676
rect 591900 390674 592500 390676
rect -6696 387676 -6096 387678
rect 26004 387676 26604 387678
rect 79568 387676 79888 387678
rect 314004 387676 314604 387678
rect 340034 387676 340358 387678
rect 422004 387676 422604 387678
rect 458004 387676 458604 387678
rect 494004 387676 494604 387678
rect 530004 387676 530604 387678
rect 566004 387676 566604 387678
rect 590020 387676 590620 387678
rect -6696 387654 590620 387676
rect -6696 387418 -6514 387654
rect -6278 387418 26186 387654
rect 26422 387418 79610 387654
rect 79846 387418 314186 387654
rect 314422 387418 340078 387654
rect 340314 387418 422186 387654
rect 422422 387418 458186 387654
rect 458422 387418 494186 387654
rect 494422 387418 530186 387654
rect 530422 387418 566186 387654
rect 566422 387418 590202 387654
rect 590438 387418 590620 387654
rect -6696 387334 590620 387418
rect -6696 387098 -6514 387334
rect -6278 387098 26186 387334
rect 26422 387098 79610 387334
rect 79846 387098 314186 387334
rect 314422 387098 340078 387334
rect 340314 387098 422186 387334
rect 422422 387098 458186 387334
rect 458422 387098 494186 387334
rect 494422 387098 530186 387334
rect 530422 387098 566186 387334
rect 566422 387098 590202 387334
rect 590438 387098 590620 387334
rect -6696 387076 590620 387098
rect -6696 387074 -6096 387076
rect 26004 387074 26604 387076
rect 79568 387074 79888 387076
rect 314004 387074 314604 387076
rect 340034 387074 340358 387076
rect 422004 387074 422604 387076
rect 458004 387074 458604 387076
rect 494004 387074 494604 387076
rect 530004 387074 530604 387076
rect 566004 387074 566604 387076
rect 590020 387074 590620 387076
rect -4816 384076 -4216 384078
rect 22404 384076 23004 384078
rect 79568 384076 79888 384078
rect 310404 384076 311004 384078
rect 340034 384076 340358 384078
rect 454404 384076 455004 384078
rect 490404 384076 491004 384078
rect 526404 384076 527004 384078
rect 562404 384076 563004 384078
rect 588140 384076 588740 384078
rect -4816 384054 588740 384076
rect -4816 383818 -4634 384054
rect -4398 383818 22586 384054
rect 22822 383818 79610 384054
rect 79846 383818 310586 384054
rect 310822 383818 340078 384054
rect 340314 383818 454586 384054
rect 454822 383818 490586 384054
rect 490822 383818 526586 384054
rect 526822 383818 562586 384054
rect 562822 383818 588322 384054
rect 588558 383818 588740 384054
rect -4816 383734 588740 383818
rect -4816 383498 -4634 383734
rect -4398 383498 22586 383734
rect 22822 383498 79610 383734
rect 79846 383498 310586 383734
rect 310822 383498 340078 383734
rect 340314 383498 454586 383734
rect 454822 383498 490586 383734
rect 490822 383498 526586 383734
rect 526822 383498 562586 383734
rect 562822 383498 588322 383734
rect 588558 383498 588740 383734
rect -4816 383476 588740 383498
rect -4816 383474 -4216 383476
rect 22404 383474 23004 383476
rect 79568 383474 79888 383476
rect 310404 383474 311004 383476
rect 340034 383474 340358 383476
rect 454404 383474 455004 383476
rect 490404 383474 491004 383476
rect 526404 383474 527004 383476
rect 562404 383474 563004 383476
rect 588140 383474 588740 383476
rect -2936 380476 -2336 380478
rect 18804 380476 19404 380478
rect 54804 380476 55404 380478
rect 79568 380476 79888 380478
rect 306804 380476 307404 380478
rect 340034 380476 340358 380478
rect 450804 380476 451404 380478
rect 486804 380476 487404 380478
rect 522804 380476 523404 380478
rect 558804 380476 559404 380478
rect 586260 380476 586860 380478
rect -2936 380454 586860 380476
rect -2936 380218 -2754 380454
rect -2518 380218 18986 380454
rect 19222 380218 54986 380454
rect 55222 380218 79610 380454
rect 79846 380218 306986 380454
rect 307222 380218 340078 380454
rect 340314 380218 450986 380454
rect 451222 380218 486986 380454
rect 487222 380218 522986 380454
rect 523222 380218 558986 380454
rect 559222 380218 586442 380454
rect 586678 380218 586860 380454
rect -2936 380134 586860 380218
rect -2936 379898 -2754 380134
rect -2518 379898 18986 380134
rect 19222 379898 54986 380134
rect 55222 379898 79610 380134
rect 79846 379898 306986 380134
rect 307222 379898 340078 380134
rect 340314 379898 450986 380134
rect 451222 379898 486986 380134
rect 487222 379898 522986 380134
rect 523222 379898 558986 380134
rect 559222 379898 586442 380134
rect 586678 379898 586860 380134
rect -2936 379876 586860 379898
rect -2936 379874 -2336 379876
rect 18804 379874 19404 379876
rect 54804 379874 55404 379876
rect 79568 379874 79888 379876
rect 306804 379874 307404 379876
rect 340034 379874 340358 379876
rect 450804 379874 451404 379876
rect 486804 379874 487404 379876
rect 522804 379874 523404 379876
rect 558804 379874 559404 379876
rect 586260 379874 586860 379876
rect -7636 373276 -7036 373278
rect 11604 373276 12204 373278
rect 47604 373276 48204 373278
rect 64208 373276 64528 373278
rect 299604 373276 300204 373278
rect 335604 373276 336204 373278
rect 340482 373276 340802 373278
rect 443604 373276 444204 373278
rect 479604 373276 480204 373278
rect 515604 373276 516204 373278
rect 551604 373276 552204 373278
rect 590960 373276 591560 373278
rect -8576 373254 592500 373276
rect -8576 373018 -7454 373254
rect -7218 373018 11786 373254
rect 12022 373018 47786 373254
rect 48022 373018 64250 373254
rect 64486 373018 299786 373254
rect 300022 373018 335786 373254
rect 336022 373018 340524 373254
rect 340760 373018 443786 373254
rect 444022 373018 479786 373254
rect 480022 373018 515786 373254
rect 516022 373018 551786 373254
rect 552022 373018 591142 373254
rect 591378 373018 592500 373254
rect -8576 372934 592500 373018
rect -8576 372698 -7454 372934
rect -7218 372698 11786 372934
rect 12022 372698 47786 372934
rect 48022 372698 64250 372934
rect 64486 372698 299786 372934
rect 300022 372698 335786 372934
rect 336022 372698 340524 372934
rect 340760 372698 443786 372934
rect 444022 372698 479786 372934
rect 480022 372698 515786 372934
rect 516022 372698 551786 372934
rect 552022 372698 591142 372934
rect 591378 372698 592500 372934
rect -8576 372676 592500 372698
rect -7636 372674 -7036 372676
rect 11604 372674 12204 372676
rect 47604 372674 48204 372676
rect 64208 372674 64528 372676
rect 299604 372674 300204 372676
rect 335604 372674 336204 372676
rect 340482 372674 340802 372676
rect 443604 372674 444204 372676
rect 479604 372674 480204 372676
rect 515604 372674 516204 372676
rect 551604 372674 552204 372676
rect 590960 372674 591560 372676
rect -5756 369676 -5156 369678
rect 8004 369676 8604 369678
rect 44004 369676 44604 369678
rect 64208 369676 64528 369678
rect 296004 369676 296604 369678
rect 332004 369676 332604 369678
rect 340482 369676 340802 369678
rect 440004 369676 440604 369678
rect 476004 369676 476604 369678
rect 512004 369676 512604 369678
rect 548004 369676 548604 369678
rect 589080 369676 589680 369678
rect -6696 369654 590620 369676
rect -6696 369418 -5574 369654
rect -5338 369418 8186 369654
rect 8422 369418 44186 369654
rect 44422 369418 64250 369654
rect 64486 369418 296186 369654
rect 296422 369418 332186 369654
rect 332422 369418 340524 369654
rect 340760 369418 440186 369654
rect 440422 369418 476186 369654
rect 476422 369418 512186 369654
rect 512422 369418 548186 369654
rect 548422 369418 589262 369654
rect 589498 369418 590620 369654
rect -6696 369334 590620 369418
rect -6696 369098 -5574 369334
rect -5338 369098 8186 369334
rect 8422 369098 44186 369334
rect 44422 369098 64250 369334
rect 64486 369098 296186 369334
rect 296422 369098 332186 369334
rect 332422 369098 340524 369334
rect 340760 369098 440186 369334
rect 440422 369098 476186 369334
rect 476422 369098 512186 369334
rect 512422 369098 548186 369334
rect 548422 369098 589262 369334
rect 589498 369098 590620 369334
rect -6696 369076 590620 369098
rect -5756 369074 -5156 369076
rect 8004 369074 8604 369076
rect 44004 369074 44604 369076
rect 64208 369074 64528 369076
rect 296004 369074 296604 369076
rect 332004 369074 332604 369076
rect 340482 369074 340802 369076
rect 440004 369074 440604 369076
rect 476004 369074 476604 369076
rect 512004 369074 512604 369076
rect 548004 369074 548604 369076
rect 589080 369074 589680 369076
rect -3876 366076 -3276 366078
rect 4404 366076 5004 366078
rect 40404 366076 41004 366078
rect 64208 366076 64528 366078
rect 292404 366076 293004 366078
rect 328404 366076 329004 366078
rect 340482 366076 340802 366078
rect 436404 366076 437004 366078
rect 472404 366076 473004 366078
rect 508404 366076 509004 366078
rect 544404 366076 545004 366078
rect 580404 366076 581004 366078
rect 587200 366076 587800 366078
rect -4816 366054 588740 366076
rect -4816 365818 -3694 366054
rect -3458 365818 4586 366054
rect 4822 365818 40586 366054
rect 40822 365818 64250 366054
rect 64486 365818 292586 366054
rect 292822 365818 328586 366054
rect 328822 365818 340524 366054
rect 340760 365818 436586 366054
rect 436822 365818 472586 366054
rect 472822 365818 508586 366054
rect 508822 365818 544586 366054
rect 544822 365818 580586 366054
rect 580822 365818 587382 366054
rect 587618 365818 588740 366054
rect -4816 365734 588740 365818
rect -4816 365498 -3694 365734
rect -3458 365498 4586 365734
rect 4822 365498 40586 365734
rect 40822 365498 64250 365734
rect 64486 365498 292586 365734
rect 292822 365498 328586 365734
rect 328822 365498 340524 365734
rect 340760 365498 436586 365734
rect 436822 365498 472586 365734
rect 472822 365498 508586 365734
rect 508822 365498 544586 365734
rect 544822 365498 580586 365734
rect 580822 365498 587382 365734
rect 587618 365498 588740 365734
rect -4816 365476 588740 365498
rect -3876 365474 -3276 365476
rect 4404 365474 5004 365476
rect 40404 365474 41004 365476
rect 64208 365474 64528 365476
rect 292404 365474 293004 365476
rect 328404 365474 329004 365476
rect 340482 365474 340802 365476
rect 436404 365474 437004 365476
rect 472404 365474 473004 365476
rect 508404 365474 509004 365476
rect 544404 365474 545004 365476
rect 580404 365474 581004 365476
rect 587200 365474 587800 365476
rect -1996 362476 -1396 362478
rect 804 362476 1404 362478
rect 36804 362476 37404 362478
rect 64208 362476 64528 362478
rect 288804 362476 289404 362478
rect 324804 362476 325404 362478
rect 340482 362476 340802 362478
rect 432804 362476 433404 362478
rect 468804 362476 469404 362478
rect 504804 362476 505404 362478
rect 540804 362476 541404 362478
rect 576804 362476 577404 362478
rect 585320 362476 585920 362478
rect -2936 362454 586860 362476
rect -2936 362218 -1814 362454
rect -1578 362218 986 362454
rect 1222 362218 36986 362454
rect 37222 362218 64250 362454
rect 64486 362218 288986 362454
rect 289222 362218 324986 362454
rect 325222 362218 340524 362454
rect 340760 362218 432986 362454
rect 433222 362218 468986 362454
rect 469222 362218 504986 362454
rect 505222 362218 540986 362454
rect 541222 362218 576986 362454
rect 577222 362218 585502 362454
rect 585738 362218 586860 362454
rect -2936 362134 586860 362218
rect -2936 361898 -1814 362134
rect -1578 361898 986 362134
rect 1222 361898 36986 362134
rect 37222 361898 64250 362134
rect 64486 361898 288986 362134
rect 289222 361898 324986 362134
rect 325222 361898 340524 362134
rect 340760 361898 432986 362134
rect 433222 361898 468986 362134
rect 469222 361898 504986 362134
rect 505222 361898 540986 362134
rect 541222 361898 576986 362134
rect 577222 361898 585502 362134
rect 585738 361898 586860 362134
rect -2936 361876 586860 361898
rect -1996 361874 -1396 361876
rect 804 361874 1404 361876
rect 36804 361874 37404 361876
rect 64208 361874 64528 361876
rect 288804 361874 289404 361876
rect 324804 361874 325404 361876
rect 340482 361874 340802 361876
rect 432804 361874 433404 361876
rect 468804 361874 469404 361876
rect 504804 361874 505404 361876
rect 540804 361874 541404 361876
rect 576804 361874 577404 361876
rect 585320 361874 585920 361876
rect -8576 355276 -7976 355278
rect 29604 355276 30204 355278
rect 79568 355276 79888 355278
rect 317604 355276 318204 355278
rect 340034 355276 340358 355278
rect 425604 355276 426204 355278
rect 461604 355276 462204 355278
rect 497604 355276 498204 355278
rect 533604 355276 534204 355278
rect 569604 355276 570204 355278
rect 591900 355276 592500 355278
rect -8576 355254 592500 355276
rect -8576 355018 -8394 355254
rect -8158 355018 29786 355254
rect 30022 355018 79610 355254
rect 79846 355018 317786 355254
rect 318022 355018 340078 355254
rect 340314 355018 425786 355254
rect 426022 355018 461786 355254
rect 462022 355018 497786 355254
rect 498022 355018 533786 355254
rect 534022 355018 569786 355254
rect 570022 355018 592082 355254
rect 592318 355018 592500 355254
rect -8576 354934 592500 355018
rect -8576 354698 -8394 354934
rect -8158 354698 29786 354934
rect 30022 354698 79610 354934
rect 79846 354698 317786 354934
rect 318022 354698 340078 354934
rect 340314 354698 425786 354934
rect 426022 354698 461786 354934
rect 462022 354698 497786 354934
rect 498022 354698 533786 354934
rect 534022 354698 569786 354934
rect 570022 354698 592082 354934
rect 592318 354698 592500 354934
rect -8576 354676 592500 354698
rect -8576 354674 -7976 354676
rect 29604 354674 30204 354676
rect 79568 354674 79888 354676
rect 317604 354674 318204 354676
rect 340034 354674 340358 354676
rect 425604 354674 426204 354676
rect 461604 354674 462204 354676
rect 497604 354674 498204 354676
rect 533604 354674 534204 354676
rect 569604 354674 570204 354676
rect 591900 354674 592500 354676
rect -6696 351676 -6096 351678
rect 26004 351676 26604 351678
rect 79568 351676 79888 351678
rect 314004 351676 314604 351678
rect 340034 351676 340358 351678
rect 422004 351676 422604 351678
rect 458004 351676 458604 351678
rect 494004 351676 494604 351678
rect 530004 351676 530604 351678
rect 566004 351676 566604 351678
rect 590020 351676 590620 351678
rect -6696 351654 590620 351676
rect -6696 351418 -6514 351654
rect -6278 351418 26186 351654
rect 26422 351418 79610 351654
rect 79846 351418 314186 351654
rect 314422 351418 340078 351654
rect 340314 351418 422186 351654
rect 422422 351418 458186 351654
rect 458422 351418 494186 351654
rect 494422 351418 530186 351654
rect 530422 351418 566186 351654
rect 566422 351418 590202 351654
rect 590438 351418 590620 351654
rect -6696 351334 590620 351418
rect -6696 351098 -6514 351334
rect -6278 351098 26186 351334
rect 26422 351098 79610 351334
rect 79846 351098 314186 351334
rect 314422 351098 340078 351334
rect 340314 351098 422186 351334
rect 422422 351098 458186 351334
rect 458422 351098 494186 351334
rect 494422 351098 530186 351334
rect 530422 351098 566186 351334
rect 566422 351098 590202 351334
rect 590438 351098 590620 351334
rect -6696 351076 590620 351098
rect -6696 351074 -6096 351076
rect 26004 351074 26604 351076
rect 79568 351074 79888 351076
rect 314004 351074 314604 351076
rect 340034 351074 340358 351076
rect 422004 351074 422604 351076
rect 458004 351074 458604 351076
rect 494004 351074 494604 351076
rect 530004 351074 530604 351076
rect 566004 351074 566604 351076
rect 590020 351074 590620 351076
rect -4816 348076 -4216 348078
rect 22404 348076 23004 348078
rect 79568 348076 79888 348078
rect 310404 348076 311004 348078
rect 340034 348076 340358 348078
rect 454404 348076 455004 348078
rect 490404 348076 491004 348078
rect 526404 348076 527004 348078
rect 562404 348076 563004 348078
rect 588140 348076 588740 348078
rect -4816 348054 588740 348076
rect -4816 347818 -4634 348054
rect -4398 347818 22586 348054
rect 22822 347818 79610 348054
rect 79846 347818 310586 348054
rect 310822 347818 340078 348054
rect 340314 347818 454586 348054
rect 454822 347818 490586 348054
rect 490822 347818 526586 348054
rect 526822 347818 562586 348054
rect 562822 347818 588322 348054
rect 588558 347818 588740 348054
rect -4816 347734 588740 347818
rect -4816 347498 -4634 347734
rect -4398 347498 22586 347734
rect 22822 347498 79610 347734
rect 79846 347498 310586 347734
rect 310822 347498 340078 347734
rect 340314 347498 454586 347734
rect 454822 347498 490586 347734
rect 490822 347498 526586 347734
rect 526822 347498 562586 347734
rect 562822 347498 588322 347734
rect 588558 347498 588740 347734
rect -4816 347476 588740 347498
rect -4816 347474 -4216 347476
rect 22404 347474 23004 347476
rect 79568 347474 79888 347476
rect 310404 347474 311004 347476
rect 340034 347474 340358 347476
rect 454404 347474 455004 347476
rect 490404 347474 491004 347476
rect 526404 347474 527004 347476
rect 562404 347474 563004 347476
rect 588140 347474 588740 347476
rect -2936 344476 -2336 344478
rect 18804 344476 19404 344478
rect 54804 344476 55404 344478
rect 79568 344476 79888 344478
rect 306804 344476 307404 344478
rect 340034 344476 340358 344478
rect 450804 344476 451404 344478
rect 486804 344476 487404 344478
rect 522804 344476 523404 344478
rect 558804 344476 559404 344478
rect 586260 344476 586860 344478
rect -2936 344454 586860 344476
rect -2936 344218 -2754 344454
rect -2518 344218 18986 344454
rect 19222 344218 54986 344454
rect 55222 344218 79610 344454
rect 79846 344218 306986 344454
rect 307222 344218 340078 344454
rect 340314 344218 450986 344454
rect 451222 344218 486986 344454
rect 487222 344218 522986 344454
rect 523222 344218 558986 344454
rect 559222 344218 586442 344454
rect 586678 344218 586860 344454
rect -2936 344134 586860 344218
rect -2936 343898 -2754 344134
rect -2518 343898 18986 344134
rect 19222 343898 54986 344134
rect 55222 343898 79610 344134
rect 79846 343898 306986 344134
rect 307222 343898 340078 344134
rect 340314 343898 450986 344134
rect 451222 343898 486986 344134
rect 487222 343898 522986 344134
rect 523222 343898 558986 344134
rect 559222 343898 586442 344134
rect 586678 343898 586860 344134
rect -2936 343876 586860 343898
rect -2936 343874 -2336 343876
rect 18804 343874 19404 343876
rect 54804 343874 55404 343876
rect 79568 343874 79888 343876
rect 306804 343874 307404 343876
rect 340034 343874 340358 343876
rect 450804 343874 451404 343876
rect 486804 343874 487404 343876
rect 522804 343874 523404 343876
rect 558804 343874 559404 343876
rect 586260 343874 586860 343876
rect -7636 337276 -7036 337278
rect 11604 337276 12204 337278
rect 47604 337276 48204 337278
rect 64208 337276 64528 337278
rect 299604 337276 300204 337278
rect 335604 337276 336204 337278
rect 340482 337276 340802 337278
rect 443604 337276 444204 337278
rect 479604 337276 480204 337278
rect 515604 337276 516204 337278
rect 551604 337276 552204 337278
rect 590960 337276 591560 337278
rect -8576 337254 592500 337276
rect -8576 337018 -7454 337254
rect -7218 337018 11786 337254
rect 12022 337018 47786 337254
rect 48022 337018 64250 337254
rect 64486 337018 299786 337254
rect 300022 337018 335786 337254
rect 336022 337018 340524 337254
rect 340760 337018 443786 337254
rect 444022 337018 479786 337254
rect 480022 337018 515786 337254
rect 516022 337018 551786 337254
rect 552022 337018 591142 337254
rect 591378 337018 592500 337254
rect -8576 336934 592500 337018
rect -8576 336698 -7454 336934
rect -7218 336698 11786 336934
rect 12022 336698 47786 336934
rect 48022 336698 64250 336934
rect 64486 336698 299786 336934
rect 300022 336698 335786 336934
rect 336022 336698 340524 336934
rect 340760 336698 443786 336934
rect 444022 336698 479786 336934
rect 480022 336698 515786 336934
rect 516022 336698 551786 336934
rect 552022 336698 591142 336934
rect 591378 336698 592500 336934
rect -8576 336676 592500 336698
rect -7636 336674 -7036 336676
rect 11604 336674 12204 336676
rect 47604 336674 48204 336676
rect 64208 336674 64528 336676
rect 299604 336674 300204 336676
rect 335604 336674 336204 336676
rect 340482 336674 340802 336676
rect 443604 336674 444204 336676
rect 479604 336674 480204 336676
rect 515604 336674 516204 336676
rect 551604 336674 552204 336676
rect 590960 336674 591560 336676
rect -5756 333676 -5156 333678
rect 8004 333676 8604 333678
rect 44004 333676 44604 333678
rect 64208 333676 64528 333678
rect 296004 333676 296604 333678
rect 332004 333676 332604 333678
rect 340482 333676 340802 333678
rect 440004 333676 440604 333678
rect 476004 333676 476604 333678
rect 512004 333676 512604 333678
rect 548004 333676 548604 333678
rect 589080 333676 589680 333678
rect -6696 333654 590620 333676
rect -6696 333418 -5574 333654
rect -5338 333418 8186 333654
rect 8422 333418 44186 333654
rect 44422 333418 64250 333654
rect 64486 333418 296186 333654
rect 296422 333418 332186 333654
rect 332422 333418 340524 333654
rect 340760 333418 440186 333654
rect 440422 333418 476186 333654
rect 476422 333418 512186 333654
rect 512422 333418 548186 333654
rect 548422 333418 589262 333654
rect 589498 333418 590620 333654
rect -6696 333334 590620 333418
rect -6696 333098 -5574 333334
rect -5338 333098 8186 333334
rect 8422 333098 44186 333334
rect 44422 333098 64250 333334
rect 64486 333098 296186 333334
rect 296422 333098 332186 333334
rect 332422 333098 340524 333334
rect 340760 333098 440186 333334
rect 440422 333098 476186 333334
rect 476422 333098 512186 333334
rect 512422 333098 548186 333334
rect 548422 333098 589262 333334
rect 589498 333098 590620 333334
rect -6696 333076 590620 333098
rect -5756 333074 -5156 333076
rect 8004 333074 8604 333076
rect 44004 333074 44604 333076
rect 64208 333074 64528 333076
rect 296004 333074 296604 333076
rect 332004 333074 332604 333076
rect 340482 333074 340802 333076
rect 440004 333074 440604 333076
rect 476004 333074 476604 333076
rect 512004 333074 512604 333076
rect 548004 333074 548604 333076
rect 589080 333074 589680 333076
rect -3876 330076 -3276 330078
rect 4404 330076 5004 330078
rect 40404 330076 41004 330078
rect 64208 330076 64528 330078
rect 292404 330076 293004 330078
rect 328404 330076 329004 330078
rect 340482 330076 340802 330078
rect 436404 330076 437004 330078
rect 472404 330076 473004 330078
rect 508404 330076 509004 330078
rect 544404 330076 545004 330078
rect 580404 330076 581004 330078
rect 587200 330076 587800 330078
rect -4816 330054 588740 330076
rect -4816 329818 -3694 330054
rect -3458 329818 4586 330054
rect 4822 329818 40586 330054
rect 40822 329818 64250 330054
rect 64486 329818 292586 330054
rect 292822 329818 328586 330054
rect 328822 329818 340524 330054
rect 340760 329818 436586 330054
rect 436822 329818 472586 330054
rect 472822 329818 508586 330054
rect 508822 329818 544586 330054
rect 544822 329818 580586 330054
rect 580822 329818 587382 330054
rect 587618 329818 588740 330054
rect -4816 329734 588740 329818
rect -4816 329498 -3694 329734
rect -3458 329498 4586 329734
rect 4822 329498 40586 329734
rect 40822 329498 64250 329734
rect 64486 329498 292586 329734
rect 292822 329498 328586 329734
rect 328822 329498 340524 329734
rect 340760 329498 436586 329734
rect 436822 329498 472586 329734
rect 472822 329498 508586 329734
rect 508822 329498 544586 329734
rect 544822 329498 580586 329734
rect 580822 329498 587382 329734
rect 587618 329498 588740 329734
rect -4816 329476 588740 329498
rect -3876 329474 -3276 329476
rect 4404 329474 5004 329476
rect 40404 329474 41004 329476
rect 64208 329474 64528 329476
rect 292404 329474 293004 329476
rect 328404 329474 329004 329476
rect 340482 329474 340802 329476
rect 436404 329474 437004 329476
rect 472404 329474 473004 329476
rect 508404 329474 509004 329476
rect 544404 329474 545004 329476
rect 580404 329474 581004 329476
rect 587200 329474 587800 329476
rect -1996 326476 -1396 326478
rect 804 326476 1404 326478
rect 36804 326476 37404 326478
rect 64208 326476 64528 326478
rect 288804 326476 289404 326478
rect 324804 326476 325404 326478
rect 340482 326476 340802 326478
rect 432804 326476 433404 326478
rect 468804 326476 469404 326478
rect 504804 326476 505404 326478
rect 540804 326476 541404 326478
rect 576804 326476 577404 326478
rect 585320 326476 585920 326478
rect -2936 326454 586860 326476
rect -2936 326218 -1814 326454
rect -1578 326218 986 326454
rect 1222 326218 36986 326454
rect 37222 326218 64250 326454
rect 64486 326218 288986 326454
rect 289222 326218 324986 326454
rect 325222 326218 340524 326454
rect 340760 326218 432986 326454
rect 433222 326218 468986 326454
rect 469222 326218 504986 326454
rect 505222 326218 540986 326454
rect 541222 326218 576986 326454
rect 577222 326218 585502 326454
rect 585738 326218 586860 326454
rect -2936 326134 586860 326218
rect -2936 325898 -1814 326134
rect -1578 325898 986 326134
rect 1222 325898 36986 326134
rect 37222 325898 64250 326134
rect 64486 325898 288986 326134
rect 289222 325898 324986 326134
rect 325222 325898 340524 326134
rect 340760 325898 432986 326134
rect 433222 325898 468986 326134
rect 469222 325898 504986 326134
rect 505222 325898 540986 326134
rect 541222 325898 576986 326134
rect 577222 325898 585502 326134
rect 585738 325898 586860 326134
rect -2936 325876 586860 325898
rect -1996 325874 -1396 325876
rect 804 325874 1404 325876
rect 36804 325874 37404 325876
rect 64208 325874 64528 325876
rect 288804 325874 289404 325876
rect 324804 325874 325404 325876
rect 340482 325874 340802 325876
rect 432804 325874 433404 325876
rect 468804 325874 469404 325876
rect 504804 325874 505404 325876
rect 540804 325874 541404 325876
rect 576804 325874 577404 325876
rect 585320 325874 585920 325876
rect -8576 319276 -7976 319278
rect 29604 319276 30204 319278
rect 317604 319276 318204 319278
rect 425604 319276 426204 319278
rect 461604 319276 462204 319278
rect 497604 319276 498204 319278
rect 533604 319276 534204 319278
rect 569604 319276 570204 319278
rect 591900 319276 592500 319278
rect -8576 319254 592500 319276
rect -8576 319018 -8394 319254
rect -8158 319018 29786 319254
rect 30022 319018 317786 319254
rect 318022 319018 425786 319254
rect 426022 319018 461786 319254
rect 462022 319018 497786 319254
rect 498022 319018 533786 319254
rect 534022 319018 569786 319254
rect 570022 319018 592082 319254
rect 592318 319018 592500 319254
rect -8576 318934 592500 319018
rect -8576 318698 -8394 318934
rect -8158 318698 29786 318934
rect 30022 318698 317786 318934
rect 318022 318698 425786 318934
rect 426022 318698 461786 318934
rect 462022 318698 497786 318934
rect 498022 318698 533786 318934
rect 534022 318698 569786 318934
rect 570022 318698 592082 318934
rect 592318 318698 592500 318934
rect -8576 318676 592500 318698
rect -8576 318674 -7976 318676
rect 29604 318674 30204 318676
rect 317604 318674 318204 318676
rect 425604 318674 426204 318676
rect 461604 318674 462204 318676
rect 497604 318674 498204 318676
rect 533604 318674 534204 318676
rect 569604 318674 570204 318676
rect 591900 318674 592500 318676
rect -6696 315676 -6096 315678
rect 26004 315676 26604 315678
rect 62004 315676 62604 315678
rect 98004 315676 98604 315678
rect 134004 315676 134604 315678
rect 170004 315676 170604 315678
rect 206004 315676 206604 315678
rect 242004 315676 242604 315678
rect 278004 315676 278604 315678
rect 314004 315676 314604 315678
rect 350004 315676 350604 315678
rect 386004 315676 386604 315678
rect 422004 315676 422604 315678
rect 458004 315676 458604 315678
rect 494004 315676 494604 315678
rect 530004 315676 530604 315678
rect 566004 315676 566604 315678
rect 590020 315676 590620 315678
rect -6696 315654 590620 315676
rect -6696 315418 -6514 315654
rect -6278 315418 26186 315654
rect 26422 315418 62186 315654
rect 62422 315418 98186 315654
rect 98422 315418 134186 315654
rect 134422 315418 170186 315654
rect 170422 315418 206186 315654
rect 206422 315418 242186 315654
rect 242422 315418 278186 315654
rect 278422 315418 314186 315654
rect 314422 315418 350186 315654
rect 350422 315418 386186 315654
rect 386422 315418 422186 315654
rect 422422 315418 458186 315654
rect 458422 315418 494186 315654
rect 494422 315418 530186 315654
rect 530422 315418 566186 315654
rect 566422 315418 590202 315654
rect 590438 315418 590620 315654
rect -6696 315334 590620 315418
rect -6696 315098 -6514 315334
rect -6278 315098 26186 315334
rect 26422 315098 62186 315334
rect 62422 315098 98186 315334
rect 98422 315098 134186 315334
rect 134422 315098 170186 315334
rect 170422 315098 206186 315334
rect 206422 315098 242186 315334
rect 242422 315098 278186 315334
rect 278422 315098 314186 315334
rect 314422 315098 350186 315334
rect 350422 315098 386186 315334
rect 386422 315098 422186 315334
rect 422422 315098 458186 315334
rect 458422 315098 494186 315334
rect 494422 315098 530186 315334
rect 530422 315098 566186 315334
rect 566422 315098 590202 315334
rect 590438 315098 590620 315334
rect -6696 315076 590620 315098
rect -6696 315074 -6096 315076
rect 26004 315074 26604 315076
rect 62004 315074 62604 315076
rect 98004 315074 98604 315076
rect 134004 315074 134604 315076
rect 170004 315074 170604 315076
rect 206004 315074 206604 315076
rect 242004 315074 242604 315076
rect 278004 315074 278604 315076
rect 314004 315074 314604 315076
rect 350004 315074 350604 315076
rect 386004 315074 386604 315076
rect 422004 315074 422604 315076
rect 458004 315074 458604 315076
rect 494004 315074 494604 315076
rect 530004 315074 530604 315076
rect 566004 315074 566604 315076
rect 590020 315074 590620 315076
rect -4816 312076 -4216 312078
rect 22404 312076 23004 312078
rect 58404 312076 59004 312078
rect 94404 312076 95004 312078
rect 130404 312076 131004 312078
rect 166404 312076 167004 312078
rect 202404 312076 203004 312078
rect 238404 312076 239004 312078
rect 274404 312076 275004 312078
rect 310404 312076 311004 312078
rect 346404 312076 347004 312078
rect 382404 312076 383004 312078
rect 418404 312076 419004 312078
rect 454404 312076 455004 312078
rect 490404 312076 491004 312078
rect 526404 312076 527004 312078
rect 562404 312076 563004 312078
rect 588140 312076 588740 312078
rect -4816 312054 588740 312076
rect -4816 311818 -4634 312054
rect -4398 311818 22586 312054
rect 22822 311818 58586 312054
rect 58822 311818 94586 312054
rect 94822 311818 130586 312054
rect 130822 311818 166586 312054
rect 166822 311818 202586 312054
rect 202822 311818 238586 312054
rect 238822 311818 274586 312054
rect 274822 311818 310586 312054
rect 310822 311818 346586 312054
rect 346822 311818 382586 312054
rect 382822 311818 418586 312054
rect 418822 311818 454586 312054
rect 454822 311818 490586 312054
rect 490822 311818 526586 312054
rect 526822 311818 562586 312054
rect 562822 311818 588322 312054
rect 588558 311818 588740 312054
rect -4816 311734 588740 311818
rect -4816 311498 -4634 311734
rect -4398 311498 22586 311734
rect 22822 311498 58586 311734
rect 58822 311498 94586 311734
rect 94822 311498 130586 311734
rect 130822 311498 166586 311734
rect 166822 311498 202586 311734
rect 202822 311498 238586 311734
rect 238822 311498 274586 311734
rect 274822 311498 310586 311734
rect 310822 311498 346586 311734
rect 346822 311498 382586 311734
rect 382822 311498 418586 311734
rect 418822 311498 454586 311734
rect 454822 311498 490586 311734
rect 490822 311498 526586 311734
rect 526822 311498 562586 311734
rect 562822 311498 588322 311734
rect 588558 311498 588740 311734
rect -4816 311476 588740 311498
rect -4816 311474 -4216 311476
rect 22404 311474 23004 311476
rect 58404 311474 59004 311476
rect 94404 311474 95004 311476
rect 130404 311474 131004 311476
rect 166404 311474 167004 311476
rect 202404 311474 203004 311476
rect 238404 311474 239004 311476
rect 274404 311474 275004 311476
rect 310404 311474 311004 311476
rect 346404 311474 347004 311476
rect 382404 311474 383004 311476
rect 418404 311474 419004 311476
rect 454404 311474 455004 311476
rect 490404 311474 491004 311476
rect 526404 311474 527004 311476
rect 562404 311474 563004 311476
rect 588140 311474 588740 311476
rect -2936 308476 -2336 308478
rect 18804 308476 19404 308478
rect 54804 308476 55404 308478
rect 90804 308476 91404 308478
rect 126804 308476 127404 308478
rect 162804 308476 163404 308478
rect 198804 308476 199404 308478
rect 234804 308476 235404 308478
rect 270804 308476 271404 308478
rect 306804 308476 307404 308478
rect 342804 308476 343404 308478
rect 378804 308476 379404 308478
rect 414804 308476 415404 308478
rect 450804 308476 451404 308478
rect 486804 308476 487404 308478
rect 522804 308476 523404 308478
rect 558804 308476 559404 308478
rect 586260 308476 586860 308478
rect -2936 308454 586860 308476
rect -2936 308218 -2754 308454
rect -2518 308218 18986 308454
rect 19222 308218 54986 308454
rect 55222 308218 90986 308454
rect 91222 308218 126986 308454
rect 127222 308218 162986 308454
rect 163222 308218 198986 308454
rect 199222 308218 234986 308454
rect 235222 308218 270986 308454
rect 271222 308218 306986 308454
rect 307222 308218 342986 308454
rect 343222 308218 378986 308454
rect 379222 308218 414986 308454
rect 415222 308218 450986 308454
rect 451222 308218 486986 308454
rect 487222 308218 522986 308454
rect 523222 308218 558986 308454
rect 559222 308218 586442 308454
rect 586678 308218 586860 308454
rect -2936 308134 586860 308218
rect -2936 307898 -2754 308134
rect -2518 307898 18986 308134
rect 19222 307898 54986 308134
rect 55222 307898 90986 308134
rect 91222 307898 126986 308134
rect 127222 307898 162986 308134
rect 163222 307898 198986 308134
rect 199222 307898 234986 308134
rect 235222 307898 270986 308134
rect 271222 307898 306986 308134
rect 307222 307898 342986 308134
rect 343222 307898 378986 308134
rect 379222 307898 414986 308134
rect 415222 307898 450986 308134
rect 451222 307898 486986 308134
rect 487222 307898 522986 308134
rect 523222 307898 558986 308134
rect 559222 307898 586442 308134
rect 586678 307898 586860 308134
rect -2936 307876 586860 307898
rect -2936 307874 -2336 307876
rect 18804 307874 19404 307876
rect 54804 307874 55404 307876
rect 90804 307874 91404 307876
rect 126804 307874 127404 307876
rect 162804 307874 163404 307876
rect 198804 307874 199404 307876
rect 234804 307874 235404 307876
rect 270804 307874 271404 307876
rect 306804 307874 307404 307876
rect 342804 307874 343404 307876
rect 378804 307874 379404 307876
rect 414804 307874 415404 307876
rect 450804 307874 451404 307876
rect 486804 307874 487404 307876
rect 522804 307874 523404 307876
rect 558804 307874 559404 307876
rect 586260 307874 586860 307876
rect -7636 301276 -7036 301278
rect 11604 301276 12204 301278
rect 47604 301276 48204 301278
rect 83604 301276 84204 301278
rect 119604 301276 120204 301278
rect 155604 301276 156204 301278
rect 191604 301276 192204 301278
rect 227604 301276 228204 301278
rect 263604 301276 264204 301278
rect 299604 301276 300204 301278
rect 335604 301276 336204 301278
rect 371604 301276 372204 301278
rect 407604 301276 408204 301278
rect 443604 301276 444204 301278
rect 479604 301276 480204 301278
rect 515604 301276 516204 301278
rect 551604 301276 552204 301278
rect 590960 301276 591560 301278
rect -8576 301254 592500 301276
rect -8576 301018 -7454 301254
rect -7218 301018 11786 301254
rect 12022 301018 47786 301254
rect 48022 301018 83786 301254
rect 84022 301018 119786 301254
rect 120022 301018 155786 301254
rect 156022 301018 191786 301254
rect 192022 301018 227786 301254
rect 228022 301018 263786 301254
rect 264022 301018 299786 301254
rect 300022 301018 335786 301254
rect 336022 301018 371786 301254
rect 372022 301018 407786 301254
rect 408022 301018 443786 301254
rect 444022 301018 479786 301254
rect 480022 301018 515786 301254
rect 516022 301018 551786 301254
rect 552022 301018 591142 301254
rect 591378 301018 592500 301254
rect -8576 300934 592500 301018
rect -8576 300698 -7454 300934
rect -7218 300698 11786 300934
rect 12022 300698 47786 300934
rect 48022 300698 83786 300934
rect 84022 300698 119786 300934
rect 120022 300698 155786 300934
rect 156022 300698 191786 300934
rect 192022 300698 227786 300934
rect 228022 300698 263786 300934
rect 264022 300698 299786 300934
rect 300022 300698 335786 300934
rect 336022 300698 371786 300934
rect 372022 300698 407786 300934
rect 408022 300698 443786 300934
rect 444022 300698 479786 300934
rect 480022 300698 515786 300934
rect 516022 300698 551786 300934
rect 552022 300698 591142 300934
rect 591378 300698 592500 300934
rect -8576 300676 592500 300698
rect -7636 300674 -7036 300676
rect 11604 300674 12204 300676
rect 47604 300674 48204 300676
rect 83604 300674 84204 300676
rect 119604 300674 120204 300676
rect 155604 300674 156204 300676
rect 191604 300674 192204 300676
rect 227604 300674 228204 300676
rect 263604 300674 264204 300676
rect 299604 300674 300204 300676
rect 335604 300674 336204 300676
rect 371604 300674 372204 300676
rect 407604 300674 408204 300676
rect 443604 300674 444204 300676
rect 479604 300674 480204 300676
rect 515604 300674 516204 300676
rect 551604 300674 552204 300676
rect 590960 300674 591560 300676
rect -5756 297676 -5156 297678
rect 8004 297676 8604 297678
rect 44004 297676 44604 297678
rect 80004 297676 80604 297678
rect 116004 297676 116604 297678
rect 152004 297676 152604 297678
rect 188004 297676 188604 297678
rect 224004 297676 224604 297678
rect 260004 297676 260604 297678
rect 296004 297676 296604 297678
rect 332004 297676 332604 297678
rect 368004 297676 368604 297678
rect 404004 297676 404604 297678
rect 440004 297676 440604 297678
rect 476004 297676 476604 297678
rect 512004 297676 512604 297678
rect 548004 297676 548604 297678
rect 589080 297676 589680 297678
rect -6696 297654 590620 297676
rect -6696 297418 -5574 297654
rect -5338 297418 8186 297654
rect 8422 297418 44186 297654
rect 44422 297418 80186 297654
rect 80422 297418 116186 297654
rect 116422 297418 152186 297654
rect 152422 297418 188186 297654
rect 188422 297418 224186 297654
rect 224422 297418 260186 297654
rect 260422 297418 296186 297654
rect 296422 297418 332186 297654
rect 332422 297418 368186 297654
rect 368422 297418 404186 297654
rect 404422 297418 440186 297654
rect 440422 297418 476186 297654
rect 476422 297418 512186 297654
rect 512422 297418 548186 297654
rect 548422 297418 589262 297654
rect 589498 297418 590620 297654
rect -6696 297334 590620 297418
rect -6696 297098 -5574 297334
rect -5338 297098 8186 297334
rect 8422 297098 44186 297334
rect 44422 297098 80186 297334
rect 80422 297098 116186 297334
rect 116422 297098 152186 297334
rect 152422 297098 188186 297334
rect 188422 297098 224186 297334
rect 224422 297098 260186 297334
rect 260422 297098 296186 297334
rect 296422 297098 332186 297334
rect 332422 297098 368186 297334
rect 368422 297098 404186 297334
rect 404422 297098 440186 297334
rect 440422 297098 476186 297334
rect 476422 297098 512186 297334
rect 512422 297098 548186 297334
rect 548422 297098 589262 297334
rect 589498 297098 590620 297334
rect -6696 297076 590620 297098
rect -5756 297074 -5156 297076
rect 8004 297074 8604 297076
rect 44004 297074 44604 297076
rect 80004 297074 80604 297076
rect 116004 297074 116604 297076
rect 152004 297074 152604 297076
rect 188004 297074 188604 297076
rect 224004 297074 224604 297076
rect 260004 297074 260604 297076
rect 296004 297074 296604 297076
rect 332004 297074 332604 297076
rect 368004 297074 368604 297076
rect 404004 297074 404604 297076
rect 440004 297074 440604 297076
rect 476004 297074 476604 297076
rect 512004 297074 512604 297076
rect 548004 297074 548604 297076
rect 589080 297074 589680 297076
rect -3876 294076 -3276 294078
rect 4404 294076 5004 294078
rect 40404 294076 41004 294078
rect 76404 294076 77004 294078
rect 112404 294076 113004 294078
rect 148404 294076 149004 294078
rect 184404 294076 185004 294078
rect 220404 294076 221004 294078
rect 256404 294076 257004 294078
rect 292404 294076 293004 294078
rect 328404 294076 329004 294078
rect 364404 294076 365004 294078
rect 400404 294076 401004 294078
rect 436404 294076 437004 294078
rect 472404 294076 473004 294078
rect 508404 294076 509004 294078
rect 544404 294076 545004 294078
rect 580404 294076 581004 294078
rect 587200 294076 587800 294078
rect -4816 294054 588740 294076
rect -4816 293818 -3694 294054
rect -3458 293818 4586 294054
rect 4822 293818 40586 294054
rect 40822 293818 76586 294054
rect 76822 293818 112586 294054
rect 112822 293818 148586 294054
rect 148822 293818 184586 294054
rect 184822 293818 220586 294054
rect 220822 293818 256586 294054
rect 256822 293818 292586 294054
rect 292822 293818 328586 294054
rect 328822 293818 364586 294054
rect 364822 293818 400586 294054
rect 400822 293818 436586 294054
rect 436822 293818 472586 294054
rect 472822 293818 508586 294054
rect 508822 293818 544586 294054
rect 544822 293818 580586 294054
rect 580822 293818 587382 294054
rect 587618 293818 588740 294054
rect -4816 293734 588740 293818
rect -4816 293498 -3694 293734
rect -3458 293498 4586 293734
rect 4822 293498 40586 293734
rect 40822 293498 76586 293734
rect 76822 293498 112586 293734
rect 112822 293498 148586 293734
rect 148822 293498 184586 293734
rect 184822 293498 220586 293734
rect 220822 293498 256586 293734
rect 256822 293498 292586 293734
rect 292822 293498 328586 293734
rect 328822 293498 364586 293734
rect 364822 293498 400586 293734
rect 400822 293498 436586 293734
rect 436822 293498 472586 293734
rect 472822 293498 508586 293734
rect 508822 293498 544586 293734
rect 544822 293498 580586 293734
rect 580822 293498 587382 293734
rect 587618 293498 588740 293734
rect -4816 293476 588740 293498
rect -3876 293474 -3276 293476
rect 4404 293474 5004 293476
rect 40404 293474 41004 293476
rect 76404 293474 77004 293476
rect 112404 293474 113004 293476
rect 148404 293474 149004 293476
rect 184404 293474 185004 293476
rect 220404 293474 221004 293476
rect 256404 293474 257004 293476
rect 292404 293474 293004 293476
rect 328404 293474 329004 293476
rect 364404 293474 365004 293476
rect 400404 293474 401004 293476
rect 436404 293474 437004 293476
rect 472404 293474 473004 293476
rect 508404 293474 509004 293476
rect 544404 293474 545004 293476
rect 580404 293474 581004 293476
rect 587200 293474 587800 293476
rect -1996 290476 -1396 290478
rect 804 290476 1404 290478
rect 36804 290476 37404 290478
rect 72804 290476 73404 290478
rect 108804 290476 109404 290478
rect 144804 290476 145404 290478
rect 180804 290476 181404 290478
rect 216804 290476 217404 290478
rect 252804 290476 253404 290478
rect 288804 290476 289404 290478
rect 324804 290476 325404 290478
rect 360804 290476 361404 290478
rect 396804 290476 397404 290478
rect 432804 290476 433404 290478
rect 468804 290476 469404 290478
rect 504804 290476 505404 290478
rect 540804 290476 541404 290478
rect 576804 290476 577404 290478
rect 585320 290476 585920 290478
rect -2936 290454 586860 290476
rect -2936 290218 -1814 290454
rect -1578 290218 986 290454
rect 1222 290218 36986 290454
rect 37222 290218 72986 290454
rect 73222 290218 108986 290454
rect 109222 290218 144986 290454
rect 145222 290218 180986 290454
rect 181222 290218 216986 290454
rect 217222 290218 252986 290454
rect 253222 290218 288986 290454
rect 289222 290218 324986 290454
rect 325222 290218 360986 290454
rect 361222 290218 396986 290454
rect 397222 290218 432986 290454
rect 433222 290218 468986 290454
rect 469222 290218 504986 290454
rect 505222 290218 540986 290454
rect 541222 290218 576986 290454
rect 577222 290218 585502 290454
rect 585738 290218 586860 290454
rect -2936 290134 586860 290218
rect -2936 289898 -1814 290134
rect -1578 289898 986 290134
rect 1222 289898 36986 290134
rect 37222 289898 72986 290134
rect 73222 289898 108986 290134
rect 109222 289898 144986 290134
rect 145222 289898 180986 290134
rect 181222 289898 216986 290134
rect 217222 289898 252986 290134
rect 253222 289898 288986 290134
rect 289222 289898 324986 290134
rect 325222 289898 360986 290134
rect 361222 289898 396986 290134
rect 397222 289898 432986 290134
rect 433222 289898 468986 290134
rect 469222 289898 504986 290134
rect 505222 289898 540986 290134
rect 541222 289898 576986 290134
rect 577222 289898 585502 290134
rect 585738 289898 586860 290134
rect -2936 289876 586860 289898
rect -1996 289874 -1396 289876
rect 804 289874 1404 289876
rect 36804 289874 37404 289876
rect 72804 289874 73404 289876
rect 108804 289874 109404 289876
rect 144804 289874 145404 289876
rect 180804 289874 181404 289876
rect 216804 289874 217404 289876
rect 252804 289874 253404 289876
rect 288804 289874 289404 289876
rect 324804 289874 325404 289876
rect 360804 289874 361404 289876
rect 396804 289874 397404 289876
rect 432804 289874 433404 289876
rect 468804 289874 469404 289876
rect 504804 289874 505404 289876
rect 540804 289874 541404 289876
rect 576804 289874 577404 289876
rect 585320 289874 585920 289876
rect -8576 283276 -7976 283278
rect 29604 283276 30204 283278
rect 65604 283276 66204 283278
rect 101604 283276 102204 283278
rect 137604 283276 138204 283278
rect 173604 283276 174204 283278
rect 209604 283276 210204 283278
rect 245604 283276 246204 283278
rect 281604 283276 282204 283278
rect 317604 283276 318204 283278
rect 353604 283276 354204 283278
rect 389604 283276 390204 283278
rect 425604 283276 426204 283278
rect 461604 283276 462204 283278
rect 497604 283276 498204 283278
rect 533604 283276 534204 283278
rect 569604 283276 570204 283278
rect 591900 283276 592500 283278
rect -8576 283254 592500 283276
rect -8576 283018 -8394 283254
rect -8158 283018 29786 283254
rect 30022 283018 65786 283254
rect 66022 283018 101786 283254
rect 102022 283018 137786 283254
rect 138022 283018 173786 283254
rect 174022 283018 209786 283254
rect 210022 283018 245786 283254
rect 246022 283018 281786 283254
rect 282022 283018 317786 283254
rect 318022 283018 353786 283254
rect 354022 283018 389786 283254
rect 390022 283018 425786 283254
rect 426022 283018 461786 283254
rect 462022 283018 497786 283254
rect 498022 283018 533786 283254
rect 534022 283018 569786 283254
rect 570022 283018 592082 283254
rect 592318 283018 592500 283254
rect -8576 282934 592500 283018
rect -8576 282698 -8394 282934
rect -8158 282698 29786 282934
rect 30022 282698 65786 282934
rect 66022 282698 101786 282934
rect 102022 282698 137786 282934
rect 138022 282698 173786 282934
rect 174022 282698 209786 282934
rect 210022 282698 245786 282934
rect 246022 282698 281786 282934
rect 282022 282698 317786 282934
rect 318022 282698 353786 282934
rect 354022 282698 389786 282934
rect 390022 282698 425786 282934
rect 426022 282698 461786 282934
rect 462022 282698 497786 282934
rect 498022 282698 533786 282934
rect 534022 282698 569786 282934
rect 570022 282698 592082 282934
rect 592318 282698 592500 282934
rect -8576 282676 592500 282698
rect -8576 282674 -7976 282676
rect 29604 282674 30204 282676
rect 65604 282674 66204 282676
rect 101604 282674 102204 282676
rect 137604 282674 138204 282676
rect 173604 282674 174204 282676
rect 209604 282674 210204 282676
rect 245604 282674 246204 282676
rect 281604 282674 282204 282676
rect 317604 282674 318204 282676
rect 353604 282674 354204 282676
rect 389604 282674 390204 282676
rect 425604 282674 426204 282676
rect 461604 282674 462204 282676
rect 497604 282674 498204 282676
rect 533604 282674 534204 282676
rect 569604 282674 570204 282676
rect 591900 282674 592500 282676
rect -6696 279676 -6096 279678
rect 26004 279676 26604 279678
rect 62004 279676 62604 279678
rect 98004 279676 98604 279678
rect 134004 279676 134604 279678
rect 170004 279676 170604 279678
rect 206004 279676 206604 279678
rect 242004 279676 242604 279678
rect 278004 279676 278604 279678
rect 314004 279676 314604 279678
rect 350004 279676 350604 279678
rect 386004 279676 386604 279678
rect 422004 279676 422604 279678
rect 458004 279676 458604 279678
rect 494004 279676 494604 279678
rect 530004 279676 530604 279678
rect 566004 279676 566604 279678
rect 590020 279676 590620 279678
rect -6696 279654 590620 279676
rect -6696 279418 -6514 279654
rect -6278 279418 26186 279654
rect 26422 279418 62186 279654
rect 62422 279418 98186 279654
rect 98422 279418 134186 279654
rect 134422 279418 170186 279654
rect 170422 279418 206186 279654
rect 206422 279418 242186 279654
rect 242422 279418 278186 279654
rect 278422 279418 314186 279654
rect 314422 279418 350186 279654
rect 350422 279418 386186 279654
rect 386422 279418 422186 279654
rect 422422 279418 458186 279654
rect 458422 279418 494186 279654
rect 494422 279418 530186 279654
rect 530422 279418 566186 279654
rect 566422 279418 590202 279654
rect 590438 279418 590620 279654
rect -6696 279334 590620 279418
rect -6696 279098 -6514 279334
rect -6278 279098 26186 279334
rect 26422 279098 62186 279334
rect 62422 279098 98186 279334
rect 98422 279098 134186 279334
rect 134422 279098 170186 279334
rect 170422 279098 206186 279334
rect 206422 279098 242186 279334
rect 242422 279098 278186 279334
rect 278422 279098 314186 279334
rect 314422 279098 350186 279334
rect 350422 279098 386186 279334
rect 386422 279098 422186 279334
rect 422422 279098 458186 279334
rect 458422 279098 494186 279334
rect 494422 279098 530186 279334
rect 530422 279098 566186 279334
rect 566422 279098 590202 279334
rect 590438 279098 590620 279334
rect -6696 279076 590620 279098
rect -6696 279074 -6096 279076
rect 26004 279074 26604 279076
rect 62004 279074 62604 279076
rect 98004 279074 98604 279076
rect 134004 279074 134604 279076
rect 170004 279074 170604 279076
rect 206004 279074 206604 279076
rect 242004 279074 242604 279076
rect 278004 279074 278604 279076
rect 314004 279074 314604 279076
rect 350004 279074 350604 279076
rect 386004 279074 386604 279076
rect 422004 279074 422604 279076
rect 458004 279074 458604 279076
rect 494004 279074 494604 279076
rect 530004 279074 530604 279076
rect 566004 279074 566604 279076
rect 590020 279074 590620 279076
rect -4816 276076 -4216 276078
rect 22404 276076 23004 276078
rect 58404 276076 59004 276078
rect 94404 276076 95004 276078
rect 130404 276076 131004 276078
rect 166404 276076 167004 276078
rect 202404 276076 203004 276078
rect 238404 276076 239004 276078
rect 274404 276076 275004 276078
rect 310404 276076 311004 276078
rect 346404 276076 347004 276078
rect 382404 276076 383004 276078
rect 418404 276076 419004 276078
rect 454404 276076 455004 276078
rect 490404 276076 491004 276078
rect 526404 276076 527004 276078
rect 562404 276076 563004 276078
rect 588140 276076 588740 276078
rect -4816 276054 588740 276076
rect -4816 275818 -4634 276054
rect -4398 275818 22586 276054
rect 22822 275818 58586 276054
rect 58822 275818 94586 276054
rect 94822 275818 130586 276054
rect 130822 275818 166586 276054
rect 166822 275818 202586 276054
rect 202822 275818 238586 276054
rect 238822 275818 274586 276054
rect 274822 275818 310586 276054
rect 310822 275818 346586 276054
rect 346822 275818 382586 276054
rect 382822 275818 418586 276054
rect 418822 275818 454586 276054
rect 454822 275818 490586 276054
rect 490822 275818 526586 276054
rect 526822 275818 562586 276054
rect 562822 275818 588322 276054
rect 588558 275818 588740 276054
rect -4816 275734 588740 275818
rect -4816 275498 -4634 275734
rect -4398 275498 22586 275734
rect 22822 275498 58586 275734
rect 58822 275498 94586 275734
rect 94822 275498 130586 275734
rect 130822 275498 166586 275734
rect 166822 275498 202586 275734
rect 202822 275498 238586 275734
rect 238822 275498 274586 275734
rect 274822 275498 310586 275734
rect 310822 275498 346586 275734
rect 346822 275498 382586 275734
rect 382822 275498 418586 275734
rect 418822 275498 454586 275734
rect 454822 275498 490586 275734
rect 490822 275498 526586 275734
rect 526822 275498 562586 275734
rect 562822 275498 588322 275734
rect 588558 275498 588740 275734
rect -4816 275476 588740 275498
rect -4816 275474 -4216 275476
rect 22404 275474 23004 275476
rect 58404 275474 59004 275476
rect 94404 275474 95004 275476
rect 130404 275474 131004 275476
rect 166404 275474 167004 275476
rect 202404 275474 203004 275476
rect 238404 275474 239004 275476
rect 274404 275474 275004 275476
rect 310404 275474 311004 275476
rect 346404 275474 347004 275476
rect 382404 275474 383004 275476
rect 418404 275474 419004 275476
rect 454404 275474 455004 275476
rect 490404 275474 491004 275476
rect 526404 275474 527004 275476
rect 562404 275474 563004 275476
rect 588140 275474 588740 275476
rect -2936 272476 -2336 272478
rect 18804 272476 19404 272478
rect 54804 272476 55404 272478
rect 90804 272476 91404 272478
rect 126804 272476 127404 272478
rect 162804 272476 163404 272478
rect 198804 272476 199404 272478
rect 234804 272476 235404 272478
rect 270804 272476 271404 272478
rect 306804 272476 307404 272478
rect 342804 272476 343404 272478
rect 378804 272476 379404 272478
rect 414804 272476 415404 272478
rect 450804 272476 451404 272478
rect 486804 272476 487404 272478
rect 522804 272476 523404 272478
rect 558804 272476 559404 272478
rect 586260 272476 586860 272478
rect -2936 272454 586860 272476
rect -2936 272218 -2754 272454
rect -2518 272218 18986 272454
rect 19222 272218 54986 272454
rect 55222 272218 90986 272454
rect 91222 272218 126986 272454
rect 127222 272218 162986 272454
rect 163222 272218 198986 272454
rect 199222 272218 234986 272454
rect 235222 272218 270986 272454
rect 271222 272218 306986 272454
rect 307222 272218 342986 272454
rect 343222 272218 378986 272454
rect 379222 272218 414986 272454
rect 415222 272218 450986 272454
rect 451222 272218 486986 272454
rect 487222 272218 522986 272454
rect 523222 272218 558986 272454
rect 559222 272218 586442 272454
rect 586678 272218 586860 272454
rect -2936 272134 586860 272218
rect -2936 271898 -2754 272134
rect -2518 271898 18986 272134
rect 19222 271898 54986 272134
rect 55222 271898 90986 272134
rect 91222 271898 126986 272134
rect 127222 271898 162986 272134
rect 163222 271898 198986 272134
rect 199222 271898 234986 272134
rect 235222 271898 270986 272134
rect 271222 271898 306986 272134
rect 307222 271898 342986 272134
rect 343222 271898 378986 272134
rect 379222 271898 414986 272134
rect 415222 271898 450986 272134
rect 451222 271898 486986 272134
rect 487222 271898 522986 272134
rect 523222 271898 558986 272134
rect 559222 271898 586442 272134
rect 586678 271898 586860 272134
rect -2936 271876 586860 271898
rect -2936 271874 -2336 271876
rect 18804 271874 19404 271876
rect 54804 271874 55404 271876
rect 90804 271874 91404 271876
rect 126804 271874 127404 271876
rect 162804 271874 163404 271876
rect 198804 271874 199404 271876
rect 234804 271874 235404 271876
rect 270804 271874 271404 271876
rect 306804 271874 307404 271876
rect 342804 271874 343404 271876
rect 378804 271874 379404 271876
rect 414804 271874 415404 271876
rect 450804 271874 451404 271876
rect 486804 271874 487404 271876
rect 522804 271874 523404 271876
rect 558804 271874 559404 271876
rect 586260 271874 586860 271876
rect -7636 265276 -7036 265278
rect 11604 265276 12204 265278
rect 47604 265276 48204 265278
rect 83604 265276 84204 265278
rect 119604 265276 120204 265278
rect 155604 265276 156204 265278
rect 191604 265276 192204 265278
rect 227604 265276 228204 265278
rect 263604 265276 264204 265278
rect 299604 265276 300204 265278
rect 335604 265276 336204 265278
rect 371604 265276 372204 265278
rect 407604 265276 408204 265278
rect 443604 265276 444204 265278
rect 479604 265276 480204 265278
rect 515604 265276 516204 265278
rect 551604 265276 552204 265278
rect 590960 265276 591560 265278
rect -8576 265254 592500 265276
rect -8576 265018 -7454 265254
rect -7218 265018 11786 265254
rect 12022 265018 47786 265254
rect 48022 265018 83786 265254
rect 84022 265018 119786 265254
rect 120022 265018 155786 265254
rect 156022 265018 191786 265254
rect 192022 265018 227786 265254
rect 228022 265018 263786 265254
rect 264022 265018 299786 265254
rect 300022 265018 335786 265254
rect 336022 265018 371786 265254
rect 372022 265018 407786 265254
rect 408022 265018 443786 265254
rect 444022 265018 479786 265254
rect 480022 265018 515786 265254
rect 516022 265018 551786 265254
rect 552022 265018 591142 265254
rect 591378 265018 592500 265254
rect -8576 264934 592500 265018
rect -8576 264698 -7454 264934
rect -7218 264698 11786 264934
rect 12022 264698 47786 264934
rect 48022 264698 83786 264934
rect 84022 264698 119786 264934
rect 120022 264698 155786 264934
rect 156022 264698 191786 264934
rect 192022 264698 227786 264934
rect 228022 264698 263786 264934
rect 264022 264698 299786 264934
rect 300022 264698 335786 264934
rect 336022 264698 371786 264934
rect 372022 264698 407786 264934
rect 408022 264698 443786 264934
rect 444022 264698 479786 264934
rect 480022 264698 515786 264934
rect 516022 264698 551786 264934
rect 552022 264698 591142 264934
rect 591378 264698 592500 264934
rect -8576 264676 592500 264698
rect -7636 264674 -7036 264676
rect 11604 264674 12204 264676
rect 47604 264674 48204 264676
rect 83604 264674 84204 264676
rect 119604 264674 120204 264676
rect 155604 264674 156204 264676
rect 191604 264674 192204 264676
rect 227604 264674 228204 264676
rect 263604 264674 264204 264676
rect 299604 264674 300204 264676
rect 335604 264674 336204 264676
rect 371604 264674 372204 264676
rect 407604 264674 408204 264676
rect 443604 264674 444204 264676
rect 479604 264674 480204 264676
rect 515604 264674 516204 264676
rect 551604 264674 552204 264676
rect 590960 264674 591560 264676
rect -5756 261676 -5156 261678
rect 8004 261676 8604 261678
rect 44004 261676 44604 261678
rect 80004 261676 80604 261678
rect 116004 261676 116604 261678
rect 152004 261676 152604 261678
rect 188004 261676 188604 261678
rect 224004 261676 224604 261678
rect 260004 261676 260604 261678
rect 296004 261676 296604 261678
rect 332004 261676 332604 261678
rect 368004 261676 368604 261678
rect 404004 261676 404604 261678
rect 440004 261676 440604 261678
rect 476004 261676 476604 261678
rect 512004 261676 512604 261678
rect 548004 261676 548604 261678
rect 589080 261676 589680 261678
rect -6696 261654 590620 261676
rect -6696 261418 -5574 261654
rect -5338 261418 8186 261654
rect 8422 261418 44186 261654
rect 44422 261418 80186 261654
rect 80422 261418 116186 261654
rect 116422 261418 152186 261654
rect 152422 261418 188186 261654
rect 188422 261418 224186 261654
rect 224422 261418 260186 261654
rect 260422 261418 296186 261654
rect 296422 261418 332186 261654
rect 332422 261418 368186 261654
rect 368422 261418 404186 261654
rect 404422 261418 440186 261654
rect 440422 261418 476186 261654
rect 476422 261418 512186 261654
rect 512422 261418 548186 261654
rect 548422 261418 589262 261654
rect 589498 261418 590620 261654
rect -6696 261334 590620 261418
rect -6696 261098 -5574 261334
rect -5338 261098 8186 261334
rect 8422 261098 44186 261334
rect 44422 261098 80186 261334
rect 80422 261098 116186 261334
rect 116422 261098 152186 261334
rect 152422 261098 188186 261334
rect 188422 261098 224186 261334
rect 224422 261098 260186 261334
rect 260422 261098 296186 261334
rect 296422 261098 332186 261334
rect 332422 261098 368186 261334
rect 368422 261098 404186 261334
rect 404422 261098 440186 261334
rect 440422 261098 476186 261334
rect 476422 261098 512186 261334
rect 512422 261098 548186 261334
rect 548422 261098 589262 261334
rect 589498 261098 590620 261334
rect -6696 261076 590620 261098
rect -5756 261074 -5156 261076
rect 8004 261074 8604 261076
rect 44004 261074 44604 261076
rect 80004 261074 80604 261076
rect 116004 261074 116604 261076
rect 152004 261074 152604 261076
rect 188004 261074 188604 261076
rect 224004 261074 224604 261076
rect 260004 261074 260604 261076
rect 296004 261074 296604 261076
rect 332004 261074 332604 261076
rect 368004 261074 368604 261076
rect 404004 261074 404604 261076
rect 440004 261074 440604 261076
rect 476004 261074 476604 261076
rect 512004 261074 512604 261076
rect 548004 261074 548604 261076
rect 589080 261074 589680 261076
rect -3876 258076 -3276 258078
rect 4404 258076 5004 258078
rect 40404 258076 41004 258078
rect 76404 258076 77004 258078
rect 112404 258076 113004 258078
rect 148404 258076 149004 258078
rect 184404 258076 185004 258078
rect 220404 258076 221004 258078
rect 256404 258076 257004 258078
rect 292404 258076 293004 258078
rect 328404 258076 329004 258078
rect 364404 258076 365004 258078
rect 400404 258076 401004 258078
rect 436404 258076 437004 258078
rect 472404 258076 473004 258078
rect 508404 258076 509004 258078
rect 544404 258076 545004 258078
rect 580404 258076 581004 258078
rect 587200 258076 587800 258078
rect -4816 258054 588740 258076
rect -4816 257818 -3694 258054
rect -3458 257818 4586 258054
rect 4822 257818 40586 258054
rect 40822 257818 76586 258054
rect 76822 257818 112586 258054
rect 112822 257818 148586 258054
rect 148822 257818 184586 258054
rect 184822 257818 220586 258054
rect 220822 257818 256586 258054
rect 256822 257818 292586 258054
rect 292822 257818 328586 258054
rect 328822 257818 364586 258054
rect 364822 257818 400586 258054
rect 400822 257818 436586 258054
rect 436822 257818 472586 258054
rect 472822 257818 508586 258054
rect 508822 257818 544586 258054
rect 544822 257818 580586 258054
rect 580822 257818 587382 258054
rect 587618 257818 588740 258054
rect -4816 257734 588740 257818
rect -4816 257498 -3694 257734
rect -3458 257498 4586 257734
rect 4822 257498 40586 257734
rect 40822 257498 76586 257734
rect 76822 257498 112586 257734
rect 112822 257498 148586 257734
rect 148822 257498 184586 257734
rect 184822 257498 220586 257734
rect 220822 257498 256586 257734
rect 256822 257498 292586 257734
rect 292822 257498 328586 257734
rect 328822 257498 364586 257734
rect 364822 257498 400586 257734
rect 400822 257498 436586 257734
rect 436822 257498 472586 257734
rect 472822 257498 508586 257734
rect 508822 257498 544586 257734
rect 544822 257498 580586 257734
rect 580822 257498 587382 257734
rect 587618 257498 588740 257734
rect -4816 257476 588740 257498
rect -3876 257474 -3276 257476
rect 4404 257474 5004 257476
rect 40404 257474 41004 257476
rect 76404 257474 77004 257476
rect 112404 257474 113004 257476
rect 148404 257474 149004 257476
rect 184404 257474 185004 257476
rect 220404 257474 221004 257476
rect 256404 257474 257004 257476
rect 292404 257474 293004 257476
rect 328404 257474 329004 257476
rect 364404 257474 365004 257476
rect 400404 257474 401004 257476
rect 436404 257474 437004 257476
rect 472404 257474 473004 257476
rect 508404 257474 509004 257476
rect 544404 257474 545004 257476
rect 580404 257474 581004 257476
rect 587200 257474 587800 257476
rect -1996 254476 -1396 254478
rect 804 254476 1404 254478
rect 36804 254476 37404 254478
rect 72804 254476 73404 254478
rect 108804 254476 109404 254478
rect 144804 254476 145404 254478
rect 180804 254476 181404 254478
rect 216804 254476 217404 254478
rect 252804 254476 253404 254478
rect 288804 254476 289404 254478
rect 324804 254476 325404 254478
rect 360804 254476 361404 254478
rect 396804 254476 397404 254478
rect 432804 254476 433404 254478
rect 468804 254476 469404 254478
rect 504804 254476 505404 254478
rect 540804 254476 541404 254478
rect 576804 254476 577404 254478
rect 585320 254476 585920 254478
rect -2936 254454 586860 254476
rect -2936 254218 -1814 254454
rect -1578 254218 986 254454
rect 1222 254218 36986 254454
rect 37222 254218 72986 254454
rect 73222 254218 108986 254454
rect 109222 254218 144986 254454
rect 145222 254218 180986 254454
rect 181222 254218 216986 254454
rect 217222 254218 252986 254454
rect 253222 254218 288986 254454
rect 289222 254218 324986 254454
rect 325222 254218 360986 254454
rect 361222 254218 396986 254454
rect 397222 254218 432986 254454
rect 433222 254218 468986 254454
rect 469222 254218 504986 254454
rect 505222 254218 540986 254454
rect 541222 254218 576986 254454
rect 577222 254218 585502 254454
rect 585738 254218 586860 254454
rect -2936 254134 586860 254218
rect -2936 253898 -1814 254134
rect -1578 253898 986 254134
rect 1222 253898 36986 254134
rect 37222 253898 72986 254134
rect 73222 253898 108986 254134
rect 109222 253898 144986 254134
rect 145222 253898 180986 254134
rect 181222 253898 216986 254134
rect 217222 253898 252986 254134
rect 253222 253898 288986 254134
rect 289222 253898 324986 254134
rect 325222 253898 360986 254134
rect 361222 253898 396986 254134
rect 397222 253898 432986 254134
rect 433222 253898 468986 254134
rect 469222 253898 504986 254134
rect 505222 253898 540986 254134
rect 541222 253898 576986 254134
rect 577222 253898 585502 254134
rect 585738 253898 586860 254134
rect -2936 253876 586860 253898
rect -1996 253874 -1396 253876
rect 804 253874 1404 253876
rect 36804 253874 37404 253876
rect 72804 253874 73404 253876
rect 108804 253874 109404 253876
rect 144804 253874 145404 253876
rect 180804 253874 181404 253876
rect 216804 253874 217404 253876
rect 252804 253874 253404 253876
rect 288804 253874 289404 253876
rect 324804 253874 325404 253876
rect 360804 253874 361404 253876
rect 396804 253874 397404 253876
rect 432804 253874 433404 253876
rect 468804 253874 469404 253876
rect 504804 253874 505404 253876
rect 540804 253874 541404 253876
rect 576804 253874 577404 253876
rect 585320 253874 585920 253876
rect -8576 247276 -7976 247278
rect 29604 247276 30204 247278
rect 65604 247276 66204 247278
rect 101604 247276 102204 247278
rect 137604 247276 138204 247278
rect 173604 247276 174204 247278
rect 209604 247276 210204 247278
rect 245604 247276 246204 247278
rect 281604 247276 282204 247278
rect 317604 247276 318204 247278
rect 353604 247276 354204 247278
rect 389604 247276 390204 247278
rect 425604 247276 426204 247278
rect 461604 247276 462204 247278
rect 497604 247276 498204 247278
rect 533604 247276 534204 247278
rect 569604 247276 570204 247278
rect 591900 247276 592500 247278
rect -8576 247254 592500 247276
rect -8576 247018 -8394 247254
rect -8158 247018 29786 247254
rect 30022 247018 65786 247254
rect 66022 247018 101786 247254
rect 102022 247018 137786 247254
rect 138022 247018 173786 247254
rect 174022 247018 209786 247254
rect 210022 247018 245786 247254
rect 246022 247018 281786 247254
rect 282022 247018 317786 247254
rect 318022 247018 353786 247254
rect 354022 247018 389786 247254
rect 390022 247018 425786 247254
rect 426022 247018 461786 247254
rect 462022 247018 497786 247254
rect 498022 247018 533786 247254
rect 534022 247018 569786 247254
rect 570022 247018 592082 247254
rect 592318 247018 592500 247254
rect -8576 246934 592500 247018
rect -8576 246698 -8394 246934
rect -8158 246698 29786 246934
rect 30022 246698 65786 246934
rect 66022 246698 101786 246934
rect 102022 246698 137786 246934
rect 138022 246698 173786 246934
rect 174022 246698 209786 246934
rect 210022 246698 245786 246934
rect 246022 246698 281786 246934
rect 282022 246698 317786 246934
rect 318022 246698 353786 246934
rect 354022 246698 389786 246934
rect 390022 246698 425786 246934
rect 426022 246698 461786 246934
rect 462022 246698 497786 246934
rect 498022 246698 533786 246934
rect 534022 246698 569786 246934
rect 570022 246698 592082 246934
rect 592318 246698 592500 246934
rect -8576 246676 592500 246698
rect -8576 246674 -7976 246676
rect 29604 246674 30204 246676
rect 65604 246674 66204 246676
rect 101604 246674 102204 246676
rect 137604 246674 138204 246676
rect 173604 246674 174204 246676
rect 209604 246674 210204 246676
rect 245604 246674 246204 246676
rect 281604 246674 282204 246676
rect 317604 246674 318204 246676
rect 353604 246674 354204 246676
rect 389604 246674 390204 246676
rect 425604 246674 426204 246676
rect 461604 246674 462204 246676
rect 497604 246674 498204 246676
rect 533604 246674 534204 246676
rect 569604 246674 570204 246676
rect 591900 246674 592500 246676
rect -6696 243676 -6096 243678
rect 26004 243676 26604 243678
rect 62004 243676 62604 243678
rect 98004 243676 98604 243678
rect 134004 243676 134604 243678
rect 170004 243676 170604 243678
rect 206004 243676 206604 243678
rect 242004 243676 242604 243678
rect 278004 243676 278604 243678
rect 314004 243676 314604 243678
rect 350004 243676 350604 243678
rect 386004 243676 386604 243678
rect 422004 243676 422604 243678
rect 458004 243676 458604 243678
rect 494004 243676 494604 243678
rect 530004 243676 530604 243678
rect 566004 243676 566604 243678
rect 590020 243676 590620 243678
rect -6696 243654 590620 243676
rect -6696 243418 -6514 243654
rect -6278 243418 26186 243654
rect 26422 243418 62186 243654
rect 62422 243418 98186 243654
rect 98422 243418 134186 243654
rect 134422 243418 170186 243654
rect 170422 243418 206186 243654
rect 206422 243418 242186 243654
rect 242422 243418 278186 243654
rect 278422 243418 314186 243654
rect 314422 243418 350186 243654
rect 350422 243418 386186 243654
rect 386422 243418 422186 243654
rect 422422 243418 458186 243654
rect 458422 243418 494186 243654
rect 494422 243418 530186 243654
rect 530422 243418 566186 243654
rect 566422 243418 590202 243654
rect 590438 243418 590620 243654
rect -6696 243334 590620 243418
rect -6696 243098 -6514 243334
rect -6278 243098 26186 243334
rect 26422 243098 62186 243334
rect 62422 243098 98186 243334
rect 98422 243098 134186 243334
rect 134422 243098 170186 243334
rect 170422 243098 206186 243334
rect 206422 243098 242186 243334
rect 242422 243098 278186 243334
rect 278422 243098 314186 243334
rect 314422 243098 350186 243334
rect 350422 243098 386186 243334
rect 386422 243098 422186 243334
rect 422422 243098 458186 243334
rect 458422 243098 494186 243334
rect 494422 243098 530186 243334
rect 530422 243098 566186 243334
rect 566422 243098 590202 243334
rect 590438 243098 590620 243334
rect -6696 243076 590620 243098
rect -6696 243074 -6096 243076
rect 26004 243074 26604 243076
rect 62004 243074 62604 243076
rect 98004 243074 98604 243076
rect 134004 243074 134604 243076
rect 170004 243074 170604 243076
rect 206004 243074 206604 243076
rect 242004 243074 242604 243076
rect 278004 243074 278604 243076
rect 314004 243074 314604 243076
rect 350004 243074 350604 243076
rect 386004 243074 386604 243076
rect 422004 243074 422604 243076
rect 458004 243074 458604 243076
rect 494004 243074 494604 243076
rect 530004 243074 530604 243076
rect 566004 243074 566604 243076
rect 590020 243074 590620 243076
rect -4816 240076 -4216 240078
rect 22404 240076 23004 240078
rect 58404 240076 59004 240078
rect 94404 240076 95004 240078
rect 130404 240076 131004 240078
rect 166404 240076 167004 240078
rect 202404 240076 203004 240078
rect 238404 240076 239004 240078
rect 274404 240076 275004 240078
rect 310404 240076 311004 240078
rect 346404 240076 347004 240078
rect 382404 240076 383004 240078
rect 418404 240076 419004 240078
rect 454404 240076 455004 240078
rect 490404 240076 491004 240078
rect 526404 240076 527004 240078
rect 562404 240076 563004 240078
rect 588140 240076 588740 240078
rect -4816 240054 588740 240076
rect -4816 239818 -4634 240054
rect -4398 239818 22586 240054
rect 22822 239818 58586 240054
rect 58822 239818 94586 240054
rect 94822 239818 130586 240054
rect 130822 239818 166586 240054
rect 166822 239818 202586 240054
rect 202822 239818 238586 240054
rect 238822 239818 274586 240054
rect 274822 239818 310586 240054
rect 310822 239818 346586 240054
rect 346822 239818 382586 240054
rect 382822 239818 418586 240054
rect 418822 239818 454586 240054
rect 454822 239818 490586 240054
rect 490822 239818 526586 240054
rect 526822 239818 562586 240054
rect 562822 239818 588322 240054
rect 588558 239818 588740 240054
rect -4816 239734 588740 239818
rect -4816 239498 -4634 239734
rect -4398 239498 22586 239734
rect 22822 239498 58586 239734
rect 58822 239498 94586 239734
rect 94822 239498 130586 239734
rect 130822 239498 166586 239734
rect 166822 239498 202586 239734
rect 202822 239498 238586 239734
rect 238822 239498 274586 239734
rect 274822 239498 310586 239734
rect 310822 239498 346586 239734
rect 346822 239498 382586 239734
rect 382822 239498 418586 239734
rect 418822 239498 454586 239734
rect 454822 239498 490586 239734
rect 490822 239498 526586 239734
rect 526822 239498 562586 239734
rect 562822 239498 588322 239734
rect 588558 239498 588740 239734
rect -4816 239476 588740 239498
rect -4816 239474 -4216 239476
rect 22404 239474 23004 239476
rect 58404 239474 59004 239476
rect 94404 239474 95004 239476
rect 130404 239474 131004 239476
rect 166404 239474 167004 239476
rect 202404 239474 203004 239476
rect 238404 239474 239004 239476
rect 274404 239474 275004 239476
rect 310404 239474 311004 239476
rect 346404 239474 347004 239476
rect 382404 239474 383004 239476
rect 418404 239474 419004 239476
rect 454404 239474 455004 239476
rect 490404 239474 491004 239476
rect 526404 239474 527004 239476
rect 562404 239474 563004 239476
rect 588140 239474 588740 239476
rect -2936 236476 -2336 236478
rect 18804 236476 19404 236478
rect 54804 236476 55404 236478
rect 90804 236476 91404 236478
rect 126804 236476 127404 236478
rect 162804 236476 163404 236478
rect 198804 236476 199404 236478
rect 234804 236476 235404 236478
rect 270804 236476 271404 236478
rect 306804 236476 307404 236478
rect 342804 236476 343404 236478
rect 378804 236476 379404 236478
rect 414804 236476 415404 236478
rect 450804 236476 451404 236478
rect 486804 236476 487404 236478
rect 522804 236476 523404 236478
rect 558804 236476 559404 236478
rect 586260 236476 586860 236478
rect -2936 236454 586860 236476
rect -2936 236218 -2754 236454
rect -2518 236218 18986 236454
rect 19222 236218 54986 236454
rect 55222 236218 90986 236454
rect 91222 236218 126986 236454
rect 127222 236218 162986 236454
rect 163222 236218 198986 236454
rect 199222 236218 234986 236454
rect 235222 236218 270986 236454
rect 271222 236218 306986 236454
rect 307222 236218 342986 236454
rect 343222 236218 378986 236454
rect 379222 236218 414986 236454
rect 415222 236218 450986 236454
rect 451222 236218 486986 236454
rect 487222 236218 522986 236454
rect 523222 236218 558986 236454
rect 559222 236218 586442 236454
rect 586678 236218 586860 236454
rect -2936 236134 586860 236218
rect -2936 235898 -2754 236134
rect -2518 235898 18986 236134
rect 19222 235898 54986 236134
rect 55222 235898 90986 236134
rect 91222 235898 126986 236134
rect 127222 235898 162986 236134
rect 163222 235898 198986 236134
rect 199222 235898 234986 236134
rect 235222 235898 270986 236134
rect 271222 235898 306986 236134
rect 307222 235898 342986 236134
rect 343222 235898 378986 236134
rect 379222 235898 414986 236134
rect 415222 235898 450986 236134
rect 451222 235898 486986 236134
rect 487222 235898 522986 236134
rect 523222 235898 558986 236134
rect 559222 235898 586442 236134
rect 586678 235898 586860 236134
rect -2936 235876 586860 235898
rect -2936 235874 -2336 235876
rect 18804 235874 19404 235876
rect 54804 235874 55404 235876
rect 90804 235874 91404 235876
rect 126804 235874 127404 235876
rect 162804 235874 163404 235876
rect 198804 235874 199404 235876
rect 234804 235874 235404 235876
rect 270804 235874 271404 235876
rect 306804 235874 307404 235876
rect 342804 235874 343404 235876
rect 378804 235874 379404 235876
rect 414804 235874 415404 235876
rect 450804 235874 451404 235876
rect 486804 235874 487404 235876
rect 522804 235874 523404 235876
rect 558804 235874 559404 235876
rect 586260 235874 586860 235876
rect -7636 229276 -7036 229278
rect 11604 229276 12204 229278
rect 47604 229276 48204 229278
rect 83604 229276 84204 229278
rect 119604 229276 120204 229278
rect 155604 229276 156204 229278
rect 191604 229276 192204 229278
rect 227604 229276 228204 229278
rect 263604 229276 264204 229278
rect 299604 229276 300204 229278
rect 335604 229276 336204 229278
rect 371604 229276 372204 229278
rect 407604 229276 408204 229278
rect 443604 229276 444204 229278
rect 479604 229276 480204 229278
rect 515604 229276 516204 229278
rect 551604 229276 552204 229278
rect 590960 229276 591560 229278
rect -8576 229254 592500 229276
rect -8576 229018 -7454 229254
rect -7218 229018 11786 229254
rect 12022 229018 47786 229254
rect 48022 229018 83786 229254
rect 84022 229018 119786 229254
rect 120022 229018 155786 229254
rect 156022 229018 191786 229254
rect 192022 229018 227786 229254
rect 228022 229018 263786 229254
rect 264022 229018 299786 229254
rect 300022 229018 335786 229254
rect 336022 229018 371786 229254
rect 372022 229018 407786 229254
rect 408022 229018 443786 229254
rect 444022 229018 479786 229254
rect 480022 229018 515786 229254
rect 516022 229018 551786 229254
rect 552022 229018 591142 229254
rect 591378 229018 592500 229254
rect -8576 228934 592500 229018
rect -8576 228698 -7454 228934
rect -7218 228698 11786 228934
rect 12022 228698 47786 228934
rect 48022 228698 83786 228934
rect 84022 228698 119786 228934
rect 120022 228698 155786 228934
rect 156022 228698 191786 228934
rect 192022 228698 227786 228934
rect 228022 228698 263786 228934
rect 264022 228698 299786 228934
rect 300022 228698 335786 228934
rect 336022 228698 371786 228934
rect 372022 228698 407786 228934
rect 408022 228698 443786 228934
rect 444022 228698 479786 228934
rect 480022 228698 515786 228934
rect 516022 228698 551786 228934
rect 552022 228698 591142 228934
rect 591378 228698 592500 228934
rect -8576 228676 592500 228698
rect -7636 228674 -7036 228676
rect 11604 228674 12204 228676
rect 47604 228674 48204 228676
rect 83604 228674 84204 228676
rect 119604 228674 120204 228676
rect 155604 228674 156204 228676
rect 191604 228674 192204 228676
rect 227604 228674 228204 228676
rect 263604 228674 264204 228676
rect 299604 228674 300204 228676
rect 335604 228674 336204 228676
rect 371604 228674 372204 228676
rect 407604 228674 408204 228676
rect 443604 228674 444204 228676
rect 479604 228674 480204 228676
rect 515604 228674 516204 228676
rect 551604 228674 552204 228676
rect 590960 228674 591560 228676
rect -5756 225676 -5156 225678
rect 8004 225676 8604 225678
rect 44004 225676 44604 225678
rect 80004 225676 80604 225678
rect 116004 225676 116604 225678
rect 152004 225676 152604 225678
rect 188004 225676 188604 225678
rect 224004 225676 224604 225678
rect 260004 225676 260604 225678
rect 296004 225676 296604 225678
rect 332004 225676 332604 225678
rect 368004 225676 368604 225678
rect 404004 225676 404604 225678
rect 440004 225676 440604 225678
rect 476004 225676 476604 225678
rect 512004 225676 512604 225678
rect 548004 225676 548604 225678
rect 589080 225676 589680 225678
rect -6696 225654 590620 225676
rect -6696 225418 -5574 225654
rect -5338 225418 8186 225654
rect 8422 225418 44186 225654
rect 44422 225418 80186 225654
rect 80422 225418 116186 225654
rect 116422 225418 152186 225654
rect 152422 225418 188186 225654
rect 188422 225418 224186 225654
rect 224422 225418 260186 225654
rect 260422 225418 296186 225654
rect 296422 225418 332186 225654
rect 332422 225418 368186 225654
rect 368422 225418 404186 225654
rect 404422 225418 440186 225654
rect 440422 225418 476186 225654
rect 476422 225418 512186 225654
rect 512422 225418 548186 225654
rect 548422 225418 589262 225654
rect 589498 225418 590620 225654
rect -6696 225334 590620 225418
rect -6696 225098 -5574 225334
rect -5338 225098 8186 225334
rect 8422 225098 44186 225334
rect 44422 225098 80186 225334
rect 80422 225098 116186 225334
rect 116422 225098 152186 225334
rect 152422 225098 188186 225334
rect 188422 225098 224186 225334
rect 224422 225098 260186 225334
rect 260422 225098 296186 225334
rect 296422 225098 332186 225334
rect 332422 225098 368186 225334
rect 368422 225098 404186 225334
rect 404422 225098 440186 225334
rect 440422 225098 476186 225334
rect 476422 225098 512186 225334
rect 512422 225098 548186 225334
rect 548422 225098 589262 225334
rect 589498 225098 590620 225334
rect -6696 225076 590620 225098
rect -5756 225074 -5156 225076
rect 8004 225074 8604 225076
rect 44004 225074 44604 225076
rect 80004 225074 80604 225076
rect 116004 225074 116604 225076
rect 152004 225074 152604 225076
rect 188004 225074 188604 225076
rect 224004 225074 224604 225076
rect 260004 225074 260604 225076
rect 296004 225074 296604 225076
rect 332004 225074 332604 225076
rect 368004 225074 368604 225076
rect 404004 225074 404604 225076
rect 440004 225074 440604 225076
rect 476004 225074 476604 225076
rect 512004 225074 512604 225076
rect 548004 225074 548604 225076
rect 589080 225074 589680 225076
rect -3876 222076 -3276 222078
rect 4404 222076 5004 222078
rect 40404 222076 41004 222078
rect 76404 222076 77004 222078
rect 112404 222076 113004 222078
rect 148404 222076 149004 222078
rect 184404 222076 185004 222078
rect 220404 222076 221004 222078
rect 256404 222076 257004 222078
rect 292404 222076 293004 222078
rect 328404 222076 329004 222078
rect 364404 222076 365004 222078
rect 400404 222076 401004 222078
rect 436404 222076 437004 222078
rect 472404 222076 473004 222078
rect 508404 222076 509004 222078
rect 544404 222076 545004 222078
rect 580404 222076 581004 222078
rect 587200 222076 587800 222078
rect -4816 222054 588740 222076
rect -4816 221818 -3694 222054
rect -3458 221818 4586 222054
rect 4822 221818 40586 222054
rect 40822 221818 76586 222054
rect 76822 221818 112586 222054
rect 112822 221818 148586 222054
rect 148822 221818 184586 222054
rect 184822 221818 220586 222054
rect 220822 221818 256586 222054
rect 256822 221818 292586 222054
rect 292822 221818 328586 222054
rect 328822 221818 364586 222054
rect 364822 221818 400586 222054
rect 400822 221818 436586 222054
rect 436822 221818 472586 222054
rect 472822 221818 508586 222054
rect 508822 221818 544586 222054
rect 544822 221818 580586 222054
rect 580822 221818 587382 222054
rect 587618 221818 588740 222054
rect -4816 221734 588740 221818
rect -4816 221498 -3694 221734
rect -3458 221498 4586 221734
rect 4822 221498 40586 221734
rect 40822 221498 76586 221734
rect 76822 221498 112586 221734
rect 112822 221498 148586 221734
rect 148822 221498 184586 221734
rect 184822 221498 220586 221734
rect 220822 221498 256586 221734
rect 256822 221498 292586 221734
rect 292822 221498 328586 221734
rect 328822 221498 364586 221734
rect 364822 221498 400586 221734
rect 400822 221498 436586 221734
rect 436822 221498 472586 221734
rect 472822 221498 508586 221734
rect 508822 221498 544586 221734
rect 544822 221498 580586 221734
rect 580822 221498 587382 221734
rect 587618 221498 588740 221734
rect -4816 221476 588740 221498
rect -3876 221474 -3276 221476
rect 4404 221474 5004 221476
rect 40404 221474 41004 221476
rect 76404 221474 77004 221476
rect 112404 221474 113004 221476
rect 148404 221474 149004 221476
rect 184404 221474 185004 221476
rect 220404 221474 221004 221476
rect 256404 221474 257004 221476
rect 292404 221474 293004 221476
rect 328404 221474 329004 221476
rect 364404 221474 365004 221476
rect 400404 221474 401004 221476
rect 436404 221474 437004 221476
rect 472404 221474 473004 221476
rect 508404 221474 509004 221476
rect 544404 221474 545004 221476
rect 580404 221474 581004 221476
rect 587200 221474 587800 221476
rect -1996 218476 -1396 218478
rect 804 218476 1404 218478
rect 36804 218476 37404 218478
rect 72804 218476 73404 218478
rect 108804 218476 109404 218478
rect 144804 218476 145404 218478
rect 180804 218476 181404 218478
rect 216804 218476 217404 218478
rect 252804 218476 253404 218478
rect 288804 218476 289404 218478
rect 324804 218476 325404 218478
rect 360804 218476 361404 218478
rect 396804 218476 397404 218478
rect 432804 218476 433404 218478
rect 468804 218476 469404 218478
rect 504804 218476 505404 218478
rect 540804 218476 541404 218478
rect 576804 218476 577404 218478
rect 585320 218476 585920 218478
rect -2936 218454 586860 218476
rect -2936 218218 -1814 218454
rect -1578 218218 986 218454
rect 1222 218218 36986 218454
rect 37222 218218 72986 218454
rect 73222 218218 108986 218454
rect 109222 218218 144986 218454
rect 145222 218218 180986 218454
rect 181222 218218 216986 218454
rect 217222 218218 252986 218454
rect 253222 218218 288986 218454
rect 289222 218218 324986 218454
rect 325222 218218 360986 218454
rect 361222 218218 396986 218454
rect 397222 218218 432986 218454
rect 433222 218218 468986 218454
rect 469222 218218 504986 218454
rect 505222 218218 540986 218454
rect 541222 218218 576986 218454
rect 577222 218218 585502 218454
rect 585738 218218 586860 218454
rect -2936 218134 586860 218218
rect -2936 217898 -1814 218134
rect -1578 217898 986 218134
rect 1222 217898 36986 218134
rect 37222 217898 72986 218134
rect 73222 217898 108986 218134
rect 109222 217898 144986 218134
rect 145222 217898 180986 218134
rect 181222 217898 216986 218134
rect 217222 217898 252986 218134
rect 253222 217898 288986 218134
rect 289222 217898 324986 218134
rect 325222 217898 360986 218134
rect 361222 217898 396986 218134
rect 397222 217898 432986 218134
rect 433222 217898 468986 218134
rect 469222 217898 504986 218134
rect 505222 217898 540986 218134
rect 541222 217898 576986 218134
rect 577222 217898 585502 218134
rect 585738 217898 586860 218134
rect -2936 217876 586860 217898
rect -1996 217874 -1396 217876
rect 804 217874 1404 217876
rect 36804 217874 37404 217876
rect 72804 217874 73404 217876
rect 108804 217874 109404 217876
rect 144804 217874 145404 217876
rect 180804 217874 181404 217876
rect 216804 217874 217404 217876
rect 252804 217874 253404 217876
rect 288804 217874 289404 217876
rect 324804 217874 325404 217876
rect 360804 217874 361404 217876
rect 396804 217874 397404 217876
rect 432804 217874 433404 217876
rect 468804 217874 469404 217876
rect 504804 217874 505404 217876
rect 540804 217874 541404 217876
rect 576804 217874 577404 217876
rect 585320 217874 585920 217876
rect -8576 211276 -7976 211278
rect 29604 211276 30204 211278
rect 65604 211276 66204 211278
rect 101604 211276 102204 211278
rect 137604 211276 138204 211278
rect 173604 211276 174204 211278
rect 209604 211276 210204 211278
rect 245604 211276 246204 211278
rect 281604 211276 282204 211278
rect 317604 211276 318204 211278
rect 353604 211276 354204 211278
rect 389604 211276 390204 211278
rect 425604 211276 426204 211278
rect 461604 211276 462204 211278
rect 497604 211276 498204 211278
rect 533604 211276 534204 211278
rect 569604 211276 570204 211278
rect 591900 211276 592500 211278
rect -8576 211254 592500 211276
rect -8576 211018 -8394 211254
rect -8158 211018 29786 211254
rect 30022 211018 65786 211254
rect 66022 211018 101786 211254
rect 102022 211018 137786 211254
rect 138022 211018 173786 211254
rect 174022 211018 209786 211254
rect 210022 211018 245786 211254
rect 246022 211018 281786 211254
rect 282022 211018 317786 211254
rect 318022 211018 353786 211254
rect 354022 211018 389786 211254
rect 390022 211018 425786 211254
rect 426022 211018 461786 211254
rect 462022 211018 497786 211254
rect 498022 211018 533786 211254
rect 534022 211018 569786 211254
rect 570022 211018 592082 211254
rect 592318 211018 592500 211254
rect -8576 210934 592500 211018
rect -8576 210698 -8394 210934
rect -8158 210698 29786 210934
rect 30022 210698 65786 210934
rect 66022 210698 101786 210934
rect 102022 210698 137786 210934
rect 138022 210698 173786 210934
rect 174022 210698 209786 210934
rect 210022 210698 245786 210934
rect 246022 210698 281786 210934
rect 282022 210698 317786 210934
rect 318022 210698 353786 210934
rect 354022 210698 389786 210934
rect 390022 210698 425786 210934
rect 426022 210698 461786 210934
rect 462022 210698 497786 210934
rect 498022 210698 533786 210934
rect 534022 210698 569786 210934
rect 570022 210698 592082 210934
rect 592318 210698 592500 210934
rect -8576 210676 592500 210698
rect -8576 210674 -7976 210676
rect 29604 210674 30204 210676
rect 65604 210674 66204 210676
rect 101604 210674 102204 210676
rect 137604 210674 138204 210676
rect 173604 210674 174204 210676
rect 209604 210674 210204 210676
rect 245604 210674 246204 210676
rect 281604 210674 282204 210676
rect 317604 210674 318204 210676
rect 353604 210674 354204 210676
rect 389604 210674 390204 210676
rect 425604 210674 426204 210676
rect 461604 210674 462204 210676
rect 497604 210674 498204 210676
rect 533604 210674 534204 210676
rect 569604 210674 570204 210676
rect 591900 210674 592500 210676
rect -6696 207676 -6096 207678
rect 26004 207676 26604 207678
rect 62004 207676 62604 207678
rect 98004 207676 98604 207678
rect 134004 207676 134604 207678
rect 170004 207676 170604 207678
rect 206004 207676 206604 207678
rect 242004 207676 242604 207678
rect 278004 207676 278604 207678
rect 314004 207676 314604 207678
rect 350004 207676 350604 207678
rect 386004 207676 386604 207678
rect 422004 207676 422604 207678
rect 458004 207676 458604 207678
rect 494004 207676 494604 207678
rect 530004 207676 530604 207678
rect 566004 207676 566604 207678
rect 590020 207676 590620 207678
rect -6696 207654 590620 207676
rect -6696 207418 -6514 207654
rect -6278 207418 26186 207654
rect 26422 207418 62186 207654
rect 62422 207418 98186 207654
rect 98422 207418 134186 207654
rect 134422 207418 170186 207654
rect 170422 207418 206186 207654
rect 206422 207418 242186 207654
rect 242422 207418 278186 207654
rect 278422 207418 314186 207654
rect 314422 207418 350186 207654
rect 350422 207418 386186 207654
rect 386422 207418 422186 207654
rect 422422 207418 458186 207654
rect 458422 207418 494186 207654
rect 494422 207418 530186 207654
rect 530422 207418 566186 207654
rect 566422 207418 590202 207654
rect 590438 207418 590620 207654
rect -6696 207334 590620 207418
rect -6696 207098 -6514 207334
rect -6278 207098 26186 207334
rect 26422 207098 62186 207334
rect 62422 207098 98186 207334
rect 98422 207098 134186 207334
rect 134422 207098 170186 207334
rect 170422 207098 206186 207334
rect 206422 207098 242186 207334
rect 242422 207098 278186 207334
rect 278422 207098 314186 207334
rect 314422 207098 350186 207334
rect 350422 207098 386186 207334
rect 386422 207098 422186 207334
rect 422422 207098 458186 207334
rect 458422 207098 494186 207334
rect 494422 207098 530186 207334
rect 530422 207098 566186 207334
rect 566422 207098 590202 207334
rect 590438 207098 590620 207334
rect -6696 207076 590620 207098
rect -6696 207074 -6096 207076
rect 26004 207074 26604 207076
rect 62004 207074 62604 207076
rect 98004 207074 98604 207076
rect 134004 207074 134604 207076
rect 170004 207074 170604 207076
rect 206004 207074 206604 207076
rect 242004 207074 242604 207076
rect 278004 207074 278604 207076
rect 314004 207074 314604 207076
rect 350004 207074 350604 207076
rect 386004 207074 386604 207076
rect 422004 207074 422604 207076
rect 458004 207074 458604 207076
rect 494004 207074 494604 207076
rect 530004 207074 530604 207076
rect 566004 207074 566604 207076
rect 590020 207074 590620 207076
rect -4816 204076 -4216 204078
rect 22404 204076 23004 204078
rect 58404 204076 59004 204078
rect 94404 204076 95004 204078
rect 130404 204076 131004 204078
rect 166404 204076 167004 204078
rect 202404 204076 203004 204078
rect 238404 204076 239004 204078
rect 274404 204076 275004 204078
rect 310404 204076 311004 204078
rect 346404 204076 347004 204078
rect 382404 204076 383004 204078
rect 418404 204076 419004 204078
rect 454404 204076 455004 204078
rect 490404 204076 491004 204078
rect 526404 204076 527004 204078
rect 562404 204076 563004 204078
rect 588140 204076 588740 204078
rect -4816 204054 588740 204076
rect -4816 203818 -4634 204054
rect -4398 203818 22586 204054
rect 22822 203818 58586 204054
rect 58822 203818 94586 204054
rect 94822 203818 130586 204054
rect 130822 203818 166586 204054
rect 166822 203818 202586 204054
rect 202822 203818 238586 204054
rect 238822 203818 274586 204054
rect 274822 203818 310586 204054
rect 310822 203818 346586 204054
rect 346822 203818 382586 204054
rect 382822 203818 418586 204054
rect 418822 203818 454586 204054
rect 454822 203818 490586 204054
rect 490822 203818 526586 204054
rect 526822 203818 562586 204054
rect 562822 203818 588322 204054
rect 588558 203818 588740 204054
rect -4816 203734 588740 203818
rect -4816 203498 -4634 203734
rect -4398 203498 22586 203734
rect 22822 203498 58586 203734
rect 58822 203498 94586 203734
rect 94822 203498 130586 203734
rect 130822 203498 166586 203734
rect 166822 203498 202586 203734
rect 202822 203498 238586 203734
rect 238822 203498 274586 203734
rect 274822 203498 310586 203734
rect 310822 203498 346586 203734
rect 346822 203498 382586 203734
rect 382822 203498 418586 203734
rect 418822 203498 454586 203734
rect 454822 203498 490586 203734
rect 490822 203498 526586 203734
rect 526822 203498 562586 203734
rect 562822 203498 588322 203734
rect 588558 203498 588740 203734
rect -4816 203476 588740 203498
rect -4816 203474 -4216 203476
rect 22404 203474 23004 203476
rect 58404 203474 59004 203476
rect 94404 203474 95004 203476
rect 130404 203474 131004 203476
rect 166404 203474 167004 203476
rect 202404 203474 203004 203476
rect 238404 203474 239004 203476
rect 274404 203474 275004 203476
rect 310404 203474 311004 203476
rect 346404 203474 347004 203476
rect 382404 203474 383004 203476
rect 418404 203474 419004 203476
rect 454404 203474 455004 203476
rect 490404 203474 491004 203476
rect 526404 203474 527004 203476
rect 562404 203474 563004 203476
rect 588140 203474 588740 203476
rect -2936 200476 -2336 200478
rect 18804 200476 19404 200478
rect 54804 200476 55404 200478
rect 90804 200476 91404 200478
rect 126804 200476 127404 200478
rect 162804 200476 163404 200478
rect 198804 200476 199404 200478
rect 234804 200476 235404 200478
rect 270804 200476 271404 200478
rect 306804 200476 307404 200478
rect 342804 200476 343404 200478
rect 378804 200476 379404 200478
rect 414804 200476 415404 200478
rect 450804 200476 451404 200478
rect 486804 200476 487404 200478
rect 522804 200476 523404 200478
rect 558804 200476 559404 200478
rect 586260 200476 586860 200478
rect -2936 200454 586860 200476
rect -2936 200218 -2754 200454
rect -2518 200218 18986 200454
rect 19222 200218 54986 200454
rect 55222 200218 90986 200454
rect 91222 200218 126986 200454
rect 127222 200218 162986 200454
rect 163222 200218 198986 200454
rect 199222 200218 234986 200454
rect 235222 200218 270986 200454
rect 271222 200218 306986 200454
rect 307222 200218 342986 200454
rect 343222 200218 378986 200454
rect 379222 200218 414986 200454
rect 415222 200218 450986 200454
rect 451222 200218 486986 200454
rect 487222 200218 522986 200454
rect 523222 200218 558986 200454
rect 559222 200218 586442 200454
rect 586678 200218 586860 200454
rect -2936 200134 586860 200218
rect -2936 199898 -2754 200134
rect -2518 199898 18986 200134
rect 19222 199898 54986 200134
rect 55222 199898 90986 200134
rect 91222 199898 126986 200134
rect 127222 199898 162986 200134
rect 163222 199898 198986 200134
rect 199222 199898 234986 200134
rect 235222 199898 270986 200134
rect 271222 199898 306986 200134
rect 307222 199898 342986 200134
rect 343222 199898 378986 200134
rect 379222 199898 414986 200134
rect 415222 199898 450986 200134
rect 451222 199898 486986 200134
rect 487222 199898 522986 200134
rect 523222 199898 558986 200134
rect 559222 199898 586442 200134
rect 586678 199898 586860 200134
rect -2936 199876 586860 199898
rect -2936 199874 -2336 199876
rect 18804 199874 19404 199876
rect 54804 199874 55404 199876
rect 90804 199874 91404 199876
rect 126804 199874 127404 199876
rect 162804 199874 163404 199876
rect 198804 199874 199404 199876
rect 234804 199874 235404 199876
rect 270804 199874 271404 199876
rect 306804 199874 307404 199876
rect 342804 199874 343404 199876
rect 378804 199874 379404 199876
rect 414804 199874 415404 199876
rect 450804 199874 451404 199876
rect 486804 199874 487404 199876
rect 522804 199874 523404 199876
rect 558804 199874 559404 199876
rect 586260 199874 586860 199876
rect -7636 193276 -7036 193278
rect 11604 193276 12204 193278
rect 47604 193276 48204 193278
rect 83604 193276 84204 193278
rect 119604 193276 120204 193278
rect 155604 193276 156204 193278
rect 191604 193276 192204 193278
rect 227604 193276 228204 193278
rect 263604 193276 264204 193278
rect 299604 193276 300204 193278
rect 335604 193276 336204 193278
rect 371604 193276 372204 193278
rect 407604 193276 408204 193278
rect 443604 193276 444204 193278
rect 479604 193276 480204 193278
rect 515604 193276 516204 193278
rect 551604 193276 552204 193278
rect 590960 193276 591560 193278
rect -8576 193254 592500 193276
rect -8576 193018 -7454 193254
rect -7218 193018 11786 193254
rect 12022 193018 47786 193254
rect 48022 193018 83786 193254
rect 84022 193018 119786 193254
rect 120022 193018 155786 193254
rect 156022 193018 191786 193254
rect 192022 193018 227786 193254
rect 228022 193018 263786 193254
rect 264022 193018 299786 193254
rect 300022 193018 335786 193254
rect 336022 193018 371786 193254
rect 372022 193018 407786 193254
rect 408022 193018 443786 193254
rect 444022 193018 479786 193254
rect 480022 193018 515786 193254
rect 516022 193018 551786 193254
rect 552022 193018 591142 193254
rect 591378 193018 592500 193254
rect -8576 192934 592500 193018
rect -8576 192698 -7454 192934
rect -7218 192698 11786 192934
rect 12022 192698 47786 192934
rect 48022 192698 83786 192934
rect 84022 192698 119786 192934
rect 120022 192698 155786 192934
rect 156022 192698 191786 192934
rect 192022 192698 227786 192934
rect 228022 192698 263786 192934
rect 264022 192698 299786 192934
rect 300022 192698 335786 192934
rect 336022 192698 371786 192934
rect 372022 192698 407786 192934
rect 408022 192698 443786 192934
rect 444022 192698 479786 192934
rect 480022 192698 515786 192934
rect 516022 192698 551786 192934
rect 552022 192698 591142 192934
rect 591378 192698 592500 192934
rect -8576 192676 592500 192698
rect -7636 192674 -7036 192676
rect 11604 192674 12204 192676
rect 47604 192674 48204 192676
rect 83604 192674 84204 192676
rect 119604 192674 120204 192676
rect 155604 192674 156204 192676
rect 191604 192674 192204 192676
rect 227604 192674 228204 192676
rect 263604 192674 264204 192676
rect 299604 192674 300204 192676
rect 335604 192674 336204 192676
rect 371604 192674 372204 192676
rect 407604 192674 408204 192676
rect 443604 192674 444204 192676
rect 479604 192674 480204 192676
rect 515604 192674 516204 192676
rect 551604 192674 552204 192676
rect 590960 192674 591560 192676
rect -5756 189676 -5156 189678
rect 8004 189676 8604 189678
rect 44004 189676 44604 189678
rect 80004 189676 80604 189678
rect 116004 189676 116604 189678
rect 152004 189676 152604 189678
rect 188004 189676 188604 189678
rect 224004 189676 224604 189678
rect 260004 189676 260604 189678
rect 296004 189676 296604 189678
rect 332004 189676 332604 189678
rect 368004 189676 368604 189678
rect 404004 189676 404604 189678
rect 440004 189676 440604 189678
rect 476004 189676 476604 189678
rect 512004 189676 512604 189678
rect 548004 189676 548604 189678
rect 589080 189676 589680 189678
rect -6696 189654 590620 189676
rect -6696 189418 -5574 189654
rect -5338 189418 8186 189654
rect 8422 189418 44186 189654
rect 44422 189418 80186 189654
rect 80422 189418 116186 189654
rect 116422 189418 152186 189654
rect 152422 189418 188186 189654
rect 188422 189418 224186 189654
rect 224422 189418 260186 189654
rect 260422 189418 296186 189654
rect 296422 189418 332186 189654
rect 332422 189418 368186 189654
rect 368422 189418 404186 189654
rect 404422 189418 440186 189654
rect 440422 189418 476186 189654
rect 476422 189418 512186 189654
rect 512422 189418 548186 189654
rect 548422 189418 589262 189654
rect 589498 189418 590620 189654
rect -6696 189334 590620 189418
rect -6696 189098 -5574 189334
rect -5338 189098 8186 189334
rect 8422 189098 44186 189334
rect 44422 189098 80186 189334
rect 80422 189098 116186 189334
rect 116422 189098 152186 189334
rect 152422 189098 188186 189334
rect 188422 189098 224186 189334
rect 224422 189098 260186 189334
rect 260422 189098 296186 189334
rect 296422 189098 332186 189334
rect 332422 189098 368186 189334
rect 368422 189098 404186 189334
rect 404422 189098 440186 189334
rect 440422 189098 476186 189334
rect 476422 189098 512186 189334
rect 512422 189098 548186 189334
rect 548422 189098 589262 189334
rect 589498 189098 590620 189334
rect -6696 189076 590620 189098
rect -5756 189074 -5156 189076
rect 8004 189074 8604 189076
rect 44004 189074 44604 189076
rect 80004 189074 80604 189076
rect 116004 189074 116604 189076
rect 152004 189074 152604 189076
rect 188004 189074 188604 189076
rect 224004 189074 224604 189076
rect 260004 189074 260604 189076
rect 296004 189074 296604 189076
rect 332004 189074 332604 189076
rect 368004 189074 368604 189076
rect 404004 189074 404604 189076
rect 440004 189074 440604 189076
rect 476004 189074 476604 189076
rect 512004 189074 512604 189076
rect 548004 189074 548604 189076
rect 589080 189074 589680 189076
rect -3876 186076 -3276 186078
rect 4404 186076 5004 186078
rect 40404 186076 41004 186078
rect 76404 186076 77004 186078
rect 112404 186076 113004 186078
rect 148404 186076 149004 186078
rect 184404 186076 185004 186078
rect 220404 186076 221004 186078
rect 256404 186076 257004 186078
rect 292404 186076 293004 186078
rect 328404 186076 329004 186078
rect 364404 186076 365004 186078
rect 400404 186076 401004 186078
rect 436404 186076 437004 186078
rect 472404 186076 473004 186078
rect 508404 186076 509004 186078
rect 544404 186076 545004 186078
rect 580404 186076 581004 186078
rect 587200 186076 587800 186078
rect -4816 186054 588740 186076
rect -4816 185818 -3694 186054
rect -3458 185818 4586 186054
rect 4822 185818 40586 186054
rect 40822 185818 76586 186054
rect 76822 185818 112586 186054
rect 112822 185818 148586 186054
rect 148822 185818 184586 186054
rect 184822 185818 220586 186054
rect 220822 185818 256586 186054
rect 256822 185818 292586 186054
rect 292822 185818 328586 186054
rect 328822 185818 364586 186054
rect 364822 185818 400586 186054
rect 400822 185818 436586 186054
rect 436822 185818 472586 186054
rect 472822 185818 508586 186054
rect 508822 185818 544586 186054
rect 544822 185818 580586 186054
rect 580822 185818 587382 186054
rect 587618 185818 588740 186054
rect -4816 185734 588740 185818
rect -4816 185498 -3694 185734
rect -3458 185498 4586 185734
rect 4822 185498 40586 185734
rect 40822 185498 76586 185734
rect 76822 185498 112586 185734
rect 112822 185498 148586 185734
rect 148822 185498 184586 185734
rect 184822 185498 220586 185734
rect 220822 185498 256586 185734
rect 256822 185498 292586 185734
rect 292822 185498 328586 185734
rect 328822 185498 364586 185734
rect 364822 185498 400586 185734
rect 400822 185498 436586 185734
rect 436822 185498 472586 185734
rect 472822 185498 508586 185734
rect 508822 185498 544586 185734
rect 544822 185498 580586 185734
rect 580822 185498 587382 185734
rect 587618 185498 588740 185734
rect -4816 185476 588740 185498
rect -3876 185474 -3276 185476
rect 4404 185474 5004 185476
rect 40404 185474 41004 185476
rect 76404 185474 77004 185476
rect 112404 185474 113004 185476
rect 148404 185474 149004 185476
rect 184404 185474 185004 185476
rect 220404 185474 221004 185476
rect 256404 185474 257004 185476
rect 292404 185474 293004 185476
rect 328404 185474 329004 185476
rect 364404 185474 365004 185476
rect 400404 185474 401004 185476
rect 436404 185474 437004 185476
rect 472404 185474 473004 185476
rect 508404 185474 509004 185476
rect 544404 185474 545004 185476
rect 580404 185474 581004 185476
rect 587200 185474 587800 185476
rect -1996 182476 -1396 182478
rect 804 182476 1404 182478
rect 36804 182476 37404 182478
rect 72804 182476 73404 182478
rect 108804 182476 109404 182478
rect 144804 182476 145404 182478
rect 180804 182476 181404 182478
rect 216804 182476 217404 182478
rect 252804 182476 253404 182478
rect 288804 182476 289404 182478
rect 324804 182476 325404 182478
rect 360804 182476 361404 182478
rect 396804 182476 397404 182478
rect 432804 182476 433404 182478
rect 468804 182476 469404 182478
rect 504804 182476 505404 182478
rect 540804 182476 541404 182478
rect 576804 182476 577404 182478
rect 585320 182476 585920 182478
rect -2936 182454 586860 182476
rect -2936 182218 -1814 182454
rect -1578 182218 986 182454
rect 1222 182218 36986 182454
rect 37222 182218 72986 182454
rect 73222 182218 108986 182454
rect 109222 182218 144986 182454
rect 145222 182218 180986 182454
rect 181222 182218 216986 182454
rect 217222 182218 252986 182454
rect 253222 182218 288986 182454
rect 289222 182218 324986 182454
rect 325222 182218 360986 182454
rect 361222 182218 396986 182454
rect 397222 182218 432986 182454
rect 433222 182218 468986 182454
rect 469222 182218 504986 182454
rect 505222 182218 540986 182454
rect 541222 182218 576986 182454
rect 577222 182218 585502 182454
rect 585738 182218 586860 182454
rect -2936 182134 586860 182218
rect -2936 181898 -1814 182134
rect -1578 181898 986 182134
rect 1222 181898 36986 182134
rect 37222 181898 72986 182134
rect 73222 181898 108986 182134
rect 109222 181898 144986 182134
rect 145222 181898 180986 182134
rect 181222 181898 216986 182134
rect 217222 181898 252986 182134
rect 253222 181898 288986 182134
rect 289222 181898 324986 182134
rect 325222 181898 360986 182134
rect 361222 181898 396986 182134
rect 397222 181898 432986 182134
rect 433222 181898 468986 182134
rect 469222 181898 504986 182134
rect 505222 181898 540986 182134
rect 541222 181898 576986 182134
rect 577222 181898 585502 182134
rect 585738 181898 586860 182134
rect -2936 181876 586860 181898
rect -1996 181874 -1396 181876
rect 804 181874 1404 181876
rect 36804 181874 37404 181876
rect 72804 181874 73404 181876
rect 108804 181874 109404 181876
rect 144804 181874 145404 181876
rect 180804 181874 181404 181876
rect 216804 181874 217404 181876
rect 252804 181874 253404 181876
rect 288804 181874 289404 181876
rect 324804 181874 325404 181876
rect 360804 181874 361404 181876
rect 396804 181874 397404 181876
rect 432804 181874 433404 181876
rect 468804 181874 469404 181876
rect 504804 181874 505404 181876
rect 540804 181874 541404 181876
rect 576804 181874 577404 181876
rect 585320 181874 585920 181876
rect -8576 175276 -7976 175278
rect 29604 175276 30204 175278
rect 65604 175276 66204 175278
rect 101604 175276 102204 175278
rect 137604 175276 138204 175278
rect 173604 175276 174204 175278
rect 209604 175276 210204 175278
rect 245604 175276 246204 175278
rect 281604 175276 282204 175278
rect 317604 175276 318204 175278
rect 353604 175276 354204 175278
rect 389604 175276 390204 175278
rect 425604 175276 426204 175278
rect 461604 175276 462204 175278
rect 497604 175276 498204 175278
rect 533604 175276 534204 175278
rect 569604 175276 570204 175278
rect 591900 175276 592500 175278
rect -8576 175254 592500 175276
rect -8576 175018 -8394 175254
rect -8158 175018 29786 175254
rect 30022 175018 65786 175254
rect 66022 175018 101786 175254
rect 102022 175018 137786 175254
rect 138022 175018 173786 175254
rect 174022 175018 209786 175254
rect 210022 175018 245786 175254
rect 246022 175018 281786 175254
rect 282022 175018 317786 175254
rect 318022 175018 353786 175254
rect 354022 175018 389786 175254
rect 390022 175018 425786 175254
rect 426022 175018 461786 175254
rect 462022 175018 497786 175254
rect 498022 175018 533786 175254
rect 534022 175018 569786 175254
rect 570022 175018 592082 175254
rect 592318 175018 592500 175254
rect -8576 174934 592500 175018
rect -8576 174698 -8394 174934
rect -8158 174698 29786 174934
rect 30022 174698 65786 174934
rect 66022 174698 101786 174934
rect 102022 174698 137786 174934
rect 138022 174698 173786 174934
rect 174022 174698 209786 174934
rect 210022 174698 245786 174934
rect 246022 174698 281786 174934
rect 282022 174698 317786 174934
rect 318022 174698 353786 174934
rect 354022 174698 389786 174934
rect 390022 174698 425786 174934
rect 426022 174698 461786 174934
rect 462022 174698 497786 174934
rect 498022 174698 533786 174934
rect 534022 174698 569786 174934
rect 570022 174698 592082 174934
rect 592318 174698 592500 174934
rect -8576 174676 592500 174698
rect -8576 174674 -7976 174676
rect 29604 174674 30204 174676
rect 65604 174674 66204 174676
rect 101604 174674 102204 174676
rect 137604 174674 138204 174676
rect 173604 174674 174204 174676
rect 209604 174674 210204 174676
rect 245604 174674 246204 174676
rect 281604 174674 282204 174676
rect 317604 174674 318204 174676
rect 353604 174674 354204 174676
rect 389604 174674 390204 174676
rect 425604 174674 426204 174676
rect 461604 174674 462204 174676
rect 497604 174674 498204 174676
rect 533604 174674 534204 174676
rect 569604 174674 570204 174676
rect 591900 174674 592500 174676
rect -6696 171676 -6096 171678
rect 26004 171676 26604 171678
rect 62004 171676 62604 171678
rect 98004 171676 98604 171678
rect 134004 171676 134604 171678
rect 170004 171676 170604 171678
rect 206004 171676 206604 171678
rect 242004 171676 242604 171678
rect 278004 171676 278604 171678
rect 314004 171676 314604 171678
rect 350004 171676 350604 171678
rect 386004 171676 386604 171678
rect 422004 171676 422604 171678
rect 458004 171676 458604 171678
rect 494004 171676 494604 171678
rect 530004 171676 530604 171678
rect 566004 171676 566604 171678
rect 590020 171676 590620 171678
rect -6696 171654 590620 171676
rect -6696 171418 -6514 171654
rect -6278 171418 26186 171654
rect 26422 171418 62186 171654
rect 62422 171418 98186 171654
rect 98422 171418 134186 171654
rect 134422 171418 170186 171654
rect 170422 171418 206186 171654
rect 206422 171418 242186 171654
rect 242422 171418 278186 171654
rect 278422 171418 314186 171654
rect 314422 171418 350186 171654
rect 350422 171418 386186 171654
rect 386422 171418 422186 171654
rect 422422 171418 458186 171654
rect 458422 171418 494186 171654
rect 494422 171418 530186 171654
rect 530422 171418 566186 171654
rect 566422 171418 590202 171654
rect 590438 171418 590620 171654
rect -6696 171334 590620 171418
rect -6696 171098 -6514 171334
rect -6278 171098 26186 171334
rect 26422 171098 62186 171334
rect 62422 171098 98186 171334
rect 98422 171098 134186 171334
rect 134422 171098 170186 171334
rect 170422 171098 206186 171334
rect 206422 171098 242186 171334
rect 242422 171098 278186 171334
rect 278422 171098 314186 171334
rect 314422 171098 350186 171334
rect 350422 171098 386186 171334
rect 386422 171098 422186 171334
rect 422422 171098 458186 171334
rect 458422 171098 494186 171334
rect 494422 171098 530186 171334
rect 530422 171098 566186 171334
rect 566422 171098 590202 171334
rect 590438 171098 590620 171334
rect -6696 171076 590620 171098
rect -6696 171074 -6096 171076
rect 26004 171074 26604 171076
rect 62004 171074 62604 171076
rect 98004 171074 98604 171076
rect 134004 171074 134604 171076
rect 170004 171074 170604 171076
rect 206004 171074 206604 171076
rect 242004 171074 242604 171076
rect 278004 171074 278604 171076
rect 314004 171074 314604 171076
rect 350004 171074 350604 171076
rect 386004 171074 386604 171076
rect 422004 171074 422604 171076
rect 458004 171074 458604 171076
rect 494004 171074 494604 171076
rect 530004 171074 530604 171076
rect 566004 171074 566604 171076
rect 590020 171074 590620 171076
rect -4816 168076 -4216 168078
rect 22404 168076 23004 168078
rect 58404 168076 59004 168078
rect 94404 168076 95004 168078
rect 130404 168076 131004 168078
rect 166404 168076 167004 168078
rect 202404 168076 203004 168078
rect 238404 168076 239004 168078
rect 274404 168076 275004 168078
rect 310404 168076 311004 168078
rect 346404 168076 347004 168078
rect 382404 168076 383004 168078
rect 418404 168076 419004 168078
rect 454404 168076 455004 168078
rect 490404 168076 491004 168078
rect 526404 168076 527004 168078
rect 562404 168076 563004 168078
rect 588140 168076 588740 168078
rect -4816 168054 588740 168076
rect -4816 167818 -4634 168054
rect -4398 167818 22586 168054
rect 22822 167818 58586 168054
rect 58822 167818 94586 168054
rect 94822 167818 130586 168054
rect 130822 167818 166586 168054
rect 166822 167818 202586 168054
rect 202822 167818 238586 168054
rect 238822 167818 274586 168054
rect 274822 167818 310586 168054
rect 310822 167818 346586 168054
rect 346822 167818 382586 168054
rect 382822 167818 418586 168054
rect 418822 167818 454586 168054
rect 454822 167818 490586 168054
rect 490822 167818 526586 168054
rect 526822 167818 562586 168054
rect 562822 167818 588322 168054
rect 588558 167818 588740 168054
rect -4816 167734 588740 167818
rect -4816 167498 -4634 167734
rect -4398 167498 22586 167734
rect 22822 167498 58586 167734
rect 58822 167498 94586 167734
rect 94822 167498 130586 167734
rect 130822 167498 166586 167734
rect 166822 167498 202586 167734
rect 202822 167498 238586 167734
rect 238822 167498 274586 167734
rect 274822 167498 310586 167734
rect 310822 167498 346586 167734
rect 346822 167498 382586 167734
rect 382822 167498 418586 167734
rect 418822 167498 454586 167734
rect 454822 167498 490586 167734
rect 490822 167498 526586 167734
rect 526822 167498 562586 167734
rect 562822 167498 588322 167734
rect 588558 167498 588740 167734
rect -4816 167476 588740 167498
rect -4816 167474 -4216 167476
rect 22404 167474 23004 167476
rect 58404 167474 59004 167476
rect 94404 167474 95004 167476
rect 130404 167474 131004 167476
rect 166404 167474 167004 167476
rect 202404 167474 203004 167476
rect 238404 167474 239004 167476
rect 274404 167474 275004 167476
rect 310404 167474 311004 167476
rect 346404 167474 347004 167476
rect 382404 167474 383004 167476
rect 418404 167474 419004 167476
rect 454404 167474 455004 167476
rect 490404 167474 491004 167476
rect 526404 167474 527004 167476
rect 562404 167474 563004 167476
rect 588140 167474 588740 167476
rect -2936 164476 -2336 164478
rect 18804 164476 19404 164478
rect 54804 164476 55404 164478
rect 90804 164476 91404 164478
rect 126804 164476 127404 164478
rect 162804 164476 163404 164478
rect 198804 164476 199404 164478
rect 234804 164476 235404 164478
rect 270804 164476 271404 164478
rect 306804 164476 307404 164478
rect 342804 164476 343404 164478
rect 378804 164476 379404 164478
rect 414804 164476 415404 164478
rect 450804 164476 451404 164478
rect 486804 164476 487404 164478
rect 522804 164476 523404 164478
rect 558804 164476 559404 164478
rect 586260 164476 586860 164478
rect -2936 164454 586860 164476
rect -2936 164218 -2754 164454
rect -2518 164218 18986 164454
rect 19222 164218 54986 164454
rect 55222 164218 90986 164454
rect 91222 164218 126986 164454
rect 127222 164218 162986 164454
rect 163222 164218 198986 164454
rect 199222 164218 234986 164454
rect 235222 164218 270986 164454
rect 271222 164218 306986 164454
rect 307222 164218 342986 164454
rect 343222 164218 378986 164454
rect 379222 164218 414986 164454
rect 415222 164218 450986 164454
rect 451222 164218 486986 164454
rect 487222 164218 522986 164454
rect 523222 164218 558986 164454
rect 559222 164218 586442 164454
rect 586678 164218 586860 164454
rect -2936 164134 586860 164218
rect -2936 163898 -2754 164134
rect -2518 163898 18986 164134
rect 19222 163898 54986 164134
rect 55222 163898 90986 164134
rect 91222 163898 126986 164134
rect 127222 163898 162986 164134
rect 163222 163898 198986 164134
rect 199222 163898 234986 164134
rect 235222 163898 270986 164134
rect 271222 163898 306986 164134
rect 307222 163898 342986 164134
rect 343222 163898 378986 164134
rect 379222 163898 414986 164134
rect 415222 163898 450986 164134
rect 451222 163898 486986 164134
rect 487222 163898 522986 164134
rect 523222 163898 558986 164134
rect 559222 163898 586442 164134
rect 586678 163898 586860 164134
rect -2936 163876 586860 163898
rect -2936 163874 -2336 163876
rect 18804 163874 19404 163876
rect 54804 163874 55404 163876
rect 90804 163874 91404 163876
rect 126804 163874 127404 163876
rect 162804 163874 163404 163876
rect 198804 163874 199404 163876
rect 234804 163874 235404 163876
rect 270804 163874 271404 163876
rect 306804 163874 307404 163876
rect 342804 163874 343404 163876
rect 378804 163874 379404 163876
rect 414804 163874 415404 163876
rect 450804 163874 451404 163876
rect 486804 163874 487404 163876
rect 522804 163874 523404 163876
rect 558804 163874 559404 163876
rect 586260 163874 586860 163876
rect -7636 157276 -7036 157278
rect 11604 157276 12204 157278
rect 47604 157276 48204 157278
rect 83604 157276 84204 157278
rect 119604 157276 120204 157278
rect 155604 157276 156204 157278
rect 191604 157276 192204 157278
rect 227604 157276 228204 157278
rect 263604 157276 264204 157278
rect 299604 157276 300204 157278
rect 335604 157276 336204 157278
rect 371604 157276 372204 157278
rect 407604 157276 408204 157278
rect 443604 157276 444204 157278
rect 479604 157276 480204 157278
rect 515604 157276 516204 157278
rect 551604 157276 552204 157278
rect 590960 157276 591560 157278
rect -8576 157254 592500 157276
rect -8576 157018 -7454 157254
rect -7218 157018 11786 157254
rect 12022 157018 47786 157254
rect 48022 157018 83786 157254
rect 84022 157018 119786 157254
rect 120022 157018 155786 157254
rect 156022 157018 191786 157254
rect 192022 157018 227786 157254
rect 228022 157018 263786 157254
rect 264022 157018 299786 157254
rect 300022 157018 335786 157254
rect 336022 157018 371786 157254
rect 372022 157018 407786 157254
rect 408022 157018 443786 157254
rect 444022 157018 479786 157254
rect 480022 157018 515786 157254
rect 516022 157018 551786 157254
rect 552022 157018 591142 157254
rect 591378 157018 592500 157254
rect -8576 156934 592500 157018
rect -8576 156698 -7454 156934
rect -7218 156698 11786 156934
rect 12022 156698 47786 156934
rect 48022 156698 83786 156934
rect 84022 156698 119786 156934
rect 120022 156698 155786 156934
rect 156022 156698 191786 156934
rect 192022 156698 227786 156934
rect 228022 156698 263786 156934
rect 264022 156698 299786 156934
rect 300022 156698 335786 156934
rect 336022 156698 371786 156934
rect 372022 156698 407786 156934
rect 408022 156698 443786 156934
rect 444022 156698 479786 156934
rect 480022 156698 515786 156934
rect 516022 156698 551786 156934
rect 552022 156698 591142 156934
rect 591378 156698 592500 156934
rect -8576 156676 592500 156698
rect -7636 156674 -7036 156676
rect 11604 156674 12204 156676
rect 47604 156674 48204 156676
rect 83604 156674 84204 156676
rect 119604 156674 120204 156676
rect 155604 156674 156204 156676
rect 191604 156674 192204 156676
rect 227604 156674 228204 156676
rect 263604 156674 264204 156676
rect 299604 156674 300204 156676
rect 335604 156674 336204 156676
rect 371604 156674 372204 156676
rect 407604 156674 408204 156676
rect 443604 156674 444204 156676
rect 479604 156674 480204 156676
rect 515604 156674 516204 156676
rect 551604 156674 552204 156676
rect 590960 156674 591560 156676
rect -5756 153676 -5156 153678
rect 8004 153676 8604 153678
rect 44004 153676 44604 153678
rect 80004 153676 80604 153678
rect 116004 153676 116604 153678
rect 152004 153676 152604 153678
rect 188004 153676 188604 153678
rect 224004 153676 224604 153678
rect 260004 153676 260604 153678
rect 296004 153676 296604 153678
rect 332004 153676 332604 153678
rect 368004 153676 368604 153678
rect 404004 153676 404604 153678
rect 440004 153676 440604 153678
rect 476004 153676 476604 153678
rect 512004 153676 512604 153678
rect 548004 153676 548604 153678
rect 589080 153676 589680 153678
rect -6696 153654 590620 153676
rect -6696 153418 -5574 153654
rect -5338 153418 8186 153654
rect 8422 153418 44186 153654
rect 44422 153418 80186 153654
rect 80422 153418 116186 153654
rect 116422 153418 152186 153654
rect 152422 153418 188186 153654
rect 188422 153418 224186 153654
rect 224422 153418 260186 153654
rect 260422 153418 296186 153654
rect 296422 153418 332186 153654
rect 332422 153418 368186 153654
rect 368422 153418 404186 153654
rect 404422 153418 440186 153654
rect 440422 153418 476186 153654
rect 476422 153418 512186 153654
rect 512422 153418 548186 153654
rect 548422 153418 589262 153654
rect 589498 153418 590620 153654
rect -6696 153334 590620 153418
rect -6696 153098 -5574 153334
rect -5338 153098 8186 153334
rect 8422 153098 44186 153334
rect 44422 153098 80186 153334
rect 80422 153098 116186 153334
rect 116422 153098 152186 153334
rect 152422 153098 188186 153334
rect 188422 153098 224186 153334
rect 224422 153098 260186 153334
rect 260422 153098 296186 153334
rect 296422 153098 332186 153334
rect 332422 153098 368186 153334
rect 368422 153098 404186 153334
rect 404422 153098 440186 153334
rect 440422 153098 476186 153334
rect 476422 153098 512186 153334
rect 512422 153098 548186 153334
rect 548422 153098 589262 153334
rect 589498 153098 590620 153334
rect -6696 153076 590620 153098
rect -5756 153074 -5156 153076
rect 8004 153074 8604 153076
rect 44004 153074 44604 153076
rect 80004 153074 80604 153076
rect 116004 153074 116604 153076
rect 152004 153074 152604 153076
rect 188004 153074 188604 153076
rect 224004 153074 224604 153076
rect 260004 153074 260604 153076
rect 296004 153074 296604 153076
rect 332004 153074 332604 153076
rect 368004 153074 368604 153076
rect 404004 153074 404604 153076
rect 440004 153074 440604 153076
rect 476004 153074 476604 153076
rect 512004 153074 512604 153076
rect 548004 153074 548604 153076
rect 589080 153074 589680 153076
rect -3876 150076 -3276 150078
rect 4404 150076 5004 150078
rect 40404 150076 41004 150078
rect 76404 150076 77004 150078
rect 112404 150076 113004 150078
rect 148404 150076 149004 150078
rect 184404 150076 185004 150078
rect 220404 150076 221004 150078
rect 256404 150076 257004 150078
rect 292404 150076 293004 150078
rect 328404 150076 329004 150078
rect 364404 150076 365004 150078
rect 400404 150076 401004 150078
rect 436404 150076 437004 150078
rect 472404 150076 473004 150078
rect 508404 150076 509004 150078
rect 544404 150076 545004 150078
rect 580404 150076 581004 150078
rect 587200 150076 587800 150078
rect -4816 150054 588740 150076
rect -4816 149818 -3694 150054
rect -3458 149818 4586 150054
rect 4822 149818 40586 150054
rect 40822 149818 76586 150054
rect 76822 149818 112586 150054
rect 112822 149818 148586 150054
rect 148822 149818 184586 150054
rect 184822 149818 220586 150054
rect 220822 149818 256586 150054
rect 256822 149818 292586 150054
rect 292822 149818 328586 150054
rect 328822 149818 364586 150054
rect 364822 149818 400586 150054
rect 400822 149818 436586 150054
rect 436822 149818 472586 150054
rect 472822 149818 508586 150054
rect 508822 149818 544586 150054
rect 544822 149818 580586 150054
rect 580822 149818 587382 150054
rect 587618 149818 588740 150054
rect -4816 149734 588740 149818
rect -4816 149498 -3694 149734
rect -3458 149498 4586 149734
rect 4822 149498 40586 149734
rect 40822 149498 76586 149734
rect 76822 149498 112586 149734
rect 112822 149498 148586 149734
rect 148822 149498 184586 149734
rect 184822 149498 220586 149734
rect 220822 149498 256586 149734
rect 256822 149498 292586 149734
rect 292822 149498 328586 149734
rect 328822 149498 364586 149734
rect 364822 149498 400586 149734
rect 400822 149498 436586 149734
rect 436822 149498 472586 149734
rect 472822 149498 508586 149734
rect 508822 149498 544586 149734
rect 544822 149498 580586 149734
rect 580822 149498 587382 149734
rect 587618 149498 588740 149734
rect -4816 149476 588740 149498
rect -3876 149474 -3276 149476
rect 4404 149474 5004 149476
rect 40404 149474 41004 149476
rect 76404 149474 77004 149476
rect 112404 149474 113004 149476
rect 148404 149474 149004 149476
rect 184404 149474 185004 149476
rect 220404 149474 221004 149476
rect 256404 149474 257004 149476
rect 292404 149474 293004 149476
rect 328404 149474 329004 149476
rect 364404 149474 365004 149476
rect 400404 149474 401004 149476
rect 436404 149474 437004 149476
rect 472404 149474 473004 149476
rect 508404 149474 509004 149476
rect 544404 149474 545004 149476
rect 580404 149474 581004 149476
rect 587200 149474 587800 149476
rect -1996 146476 -1396 146478
rect 804 146476 1404 146478
rect 36804 146476 37404 146478
rect 72804 146476 73404 146478
rect 108804 146476 109404 146478
rect 144804 146476 145404 146478
rect 180804 146476 181404 146478
rect 216804 146476 217404 146478
rect 252804 146476 253404 146478
rect 288804 146476 289404 146478
rect 324804 146476 325404 146478
rect 360804 146476 361404 146478
rect 396804 146476 397404 146478
rect 432804 146476 433404 146478
rect 468804 146476 469404 146478
rect 504804 146476 505404 146478
rect 540804 146476 541404 146478
rect 576804 146476 577404 146478
rect 585320 146476 585920 146478
rect -2936 146454 586860 146476
rect -2936 146218 -1814 146454
rect -1578 146218 986 146454
rect 1222 146218 36986 146454
rect 37222 146218 72986 146454
rect 73222 146218 108986 146454
rect 109222 146218 144986 146454
rect 145222 146218 180986 146454
rect 181222 146218 216986 146454
rect 217222 146218 252986 146454
rect 253222 146218 288986 146454
rect 289222 146218 324986 146454
rect 325222 146218 360986 146454
rect 361222 146218 396986 146454
rect 397222 146218 432986 146454
rect 433222 146218 468986 146454
rect 469222 146218 504986 146454
rect 505222 146218 540986 146454
rect 541222 146218 576986 146454
rect 577222 146218 585502 146454
rect 585738 146218 586860 146454
rect -2936 146134 586860 146218
rect -2936 145898 -1814 146134
rect -1578 145898 986 146134
rect 1222 145898 36986 146134
rect 37222 145898 72986 146134
rect 73222 145898 108986 146134
rect 109222 145898 144986 146134
rect 145222 145898 180986 146134
rect 181222 145898 216986 146134
rect 217222 145898 252986 146134
rect 253222 145898 288986 146134
rect 289222 145898 324986 146134
rect 325222 145898 360986 146134
rect 361222 145898 396986 146134
rect 397222 145898 432986 146134
rect 433222 145898 468986 146134
rect 469222 145898 504986 146134
rect 505222 145898 540986 146134
rect 541222 145898 576986 146134
rect 577222 145898 585502 146134
rect 585738 145898 586860 146134
rect -2936 145876 586860 145898
rect -1996 145874 -1396 145876
rect 804 145874 1404 145876
rect 36804 145874 37404 145876
rect 72804 145874 73404 145876
rect 108804 145874 109404 145876
rect 144804 145874 145404 145876
rect 180804 145874 181404 145876
rect 216804 145874 217404 145876
rect 252804 145874 253404 145876
rect 288804 145874 289404 145876
rect 324804 145874 325404 145876
rect 360804 145874 361404 145876
rect 396804 145874 397404 145876
rect 432804 145874 433404 145876
rect 468804 145874 469404 145876
rect 504804 145874 505404 145876
rect 540804 145874 541404 145876
rect 576804 145874 577404 145876
rect 585320 145874 585920 145876
rect -8576 139276 -7976 139278
rect 29604 139276 30204 139278
rect 65604 139276 66204 139278
rect 101604 139276 102204 139278
rect 137604 139276 138204 139278
rect 173604 139276 174204 139278
rect 209604 139276 210204 139278
rect 245604 139276 246204 139278
rect 281604 139276 282204 139278
rect 317604 139276 318204 139278
rect 353604 139276 354204 139278
rect 389604 139276 390204 139278
rect 425604 139276 426204 139278
rect 461604 139276 462204 139278
rect 497604 139276 498204 139278
rect 533604 139276 534204 139278
rect 569604 139276 570204 139278
rect 591900 139276 592500 139278
rect -8576 139254 592500 139276
rect -8576 139018 -8394 139254
rect -8158 139018 29786 139254
rect 30022 139018 65786 139254
rect 66022 139018 101786 139254
rect 102022 139018 137786 139254
rect 138022 139018 173786 139254
rect 174022 139018 209786 139254
rect 210022 139018 245786 139254
rect 246022 139018 281786 139254
rect 282022 139018 317786 139254
rect 318022 139018 353786 139254
rect 354022 139018 389786 139254
rect 390022 139018 425786 139254
rect 426022 139018 461786 139254
rect 462022 139018 497786 139254
rect 498022 139018 533786 139254
rect 534022 139018 569786 139254
rect 570022 139018 592082 139254
rect 592318 139018 592500 139254
rect -8576 138934 592500 139018
rect -8576 138698 -8394 138934
rect -8158 138698 29786 138934
rect 30022 138698 65786 138934
rect 66022 138698 101786 138934
rect 102022 138698 137786 138934
rect 138022 138698 173786 138934
rect 174022 138698 209786 138934
rect 210022 138698 245786 138934
rect 246022 138698 281786 138934
rect 282022 138698 317786 138934
rect 318022 138698 353786 138934
rect 354022 138698 389786 138934
rect 390022 138698 425786 138934
rect 426022 138698 461786 138934
rect 462022 138698 497786 138934
rect 498022 138698 533786 138934
rect 534022 138698 569786 138934
rect 570022 138698 592082 138934
rect 592318 138698 592500 138934
rect -8576 138676 592500 138698
rect -8576 138674 -7976 138676
rect 29604 138674 30204 138676
rect 65604 138674 66204 138676
rect 101604 138674 102204 138676
rect 137604 138674 138204 138676
rect 173604 138674 174204 138676
rect 209604 138674 210204 138676
rect 245604 138674 246204 138676
rect 281604 138674 282204 138676
rect 317604 138674 318204 138676
rect 353604 138674 354204 138676
rect 389604 138674 390204 138676
rect 425604 138674 426204 138676
rect 461604 138674 462204 138676
rect 497604 138674 498204 138676
rect 533604 138674 534204 138676
rect 569604 138674 570204 138676
rect 591900 138674 592500 138676
rect -6696 135676 -6096 135678
rect 26004 135676 26604 135678
rect 62004 135676 62604 135678
rect 98004 135676 98604 135678
rect 134004 135676 134604 135678
rect 170004 135676 170604 135678
rect 206004 135676 206604 135678
rect 242004 135676 242604 135678
rect 278004 135676 278604 135678
rect 314004 135676 314604 135678
rect 350004 135676 350604 135678
rect 386004 135676 386604 135678
rect 422004 135676 422604 135678
rect 458004 135676 458604 135678
rect 494004 135676 494604 135678
rect 530004 135676 530604 135678
rect 566004 135676 566604 135678
rect 590020 135676 590620 135678
rect -6696 135654 590620 135676
rect -6696 135418 -6514 135654
rect -6278 135418 26186 135654
rect 26422 135418 62186 135654
rect 62422 135418 98186 135654
rect 98422 135418 134186 135654
rect 134422 135418 170186 135654
rect 170422 135418 206186 135654
rect 206422 135418 242186 135654
rect 242422 135418 278186 135654
rect 278422 135418 314186 135654
rect 314422 135418 350186 135654
rect 350422 135418 386186 135654
rect 386422 135418 422186 135654
rect 422422 135418 458186 135654
rect 458422 135418 494186 135654
rect 494422 135418 530186 135654
rect 530422 135418 566186 135654
rect 566422 135418 590202 135654
rect 590438 135418 590620 135654
rect -6696 135334 590620 135418
rect -6696 135098 -6514 135334
rect -6278 135098 26186 135334
rect 26422 135098 62186 135334
rect 62422 135098 98186 135334
rect 98422 135098 134186 135334
rect 134422 135098 170186 135334
rect 170422 135098 206186 135334
rect 206422 135098 242186 135334
rect 242422 135098 278186 135334
rect 278422 135098 314186 135334
rect 314422 135098 350186 135334
rect 350422 135098 386186 135334
rect 386422 135098 422186 135334
rect 422422 135098 458186 135334
rect 458422 135098 494186 135334
rect 494422 135098 530186 135334
rect 530422 135098 566186 135334
rect 566422 135098 590202 135334
rect 590438 135098 590620 135334
rect -6696 135076 590620 135098
rect -6696 135074 -6096 135076
rect 26004 135074 26604 135076
rect 62004 135074 62604 135076
rect 98004 135074 98604 135076
rect 134004 135074 134604 135076
rect 170004 135074 170604 135076
rect 206004 135074 206604 135076
rect 242004 135074 242604 135076
rect 278004 135074 278604 135076
rect 314004 135074 314604 135076
rect 350004 135074 350604 135076
rect 386004 135074 386604 135076
rect 422004 135074 422604 135076
rect 458004 135074 458604 135076
rect 494004 135074 494604 135076
rect 530004 135074 530604 135076
rect 566004 135074 566604 135076
rect 590020 135074 590620 135076
rect -4816 132076 -4216 132078
rect 22404 132076 23004 132078
rect 58404 132076 59004 132078
rect 94404 132076 95004 132078
rect 130404 132076 131004 132078
rect 166404 132076 167004 132078
rect 202404 132076 203004 132078
rect 238404 132076 239004 132078
rect 274404 132076 275004 132078
rect 310404 132076 311004 132078
rect 346404 132076 347004 132078
rect 382404 132076 383004 132078
rect 418404 132076 419004 132078
rect 454404 132076 455004 132078
rect 490404 132076 491004 132078
rect 526404 132076 527004 132078
rect 562404 132076 563004 132078
rect 588140 132076 588740 132078
rect -4816 132054 588740 132076
rect -4816 131818 -4634 132054
rect -4398 131818 22586 132054
rect 22822 131818 58586 132054
rect 58822 131818 94586 132054
rect 94822 131818 130586 132054
rect 130822 131818 166586 132054
rect 166822 131818 202586 132054
rect 202822 131818 238586 132054
rect 238822 131818 274586 132054
rect 274822 131818 310586 132054
rect 310822 131818 346586 132054
rect 346822 131818 382586 132054
rect 382822 131818 418586 132054
rect 418822 131818 454586 132054
rect 454822 131818 490586 132054
rect 490822 131818 526586 132054
rect 526822 131818 562586 132054
rect 562822 131818 588322 132054
rect 588558 131818 588740 132054
rect -4816 131734 588740 131818
rect -4816 131498 -4634 131734
rect -4398 131498 22586 131734
rect 22822 131498 58586 131734
rect 58822 131498 94586 131734
rect 94822 131498 130586 131734
rect 130822 131498 166586 131734
rect 166822 131498 202586 131734
rect 202822 131498 238586 131734
rect 238822 131498 274586 131734
rect 274822 131498 310586 131734
rect 310822 131498 346586 131734
rect 346822 131498 382586 131734
rect 382822 131498 418586 131734
rect 418822 131498 454586 131734
rect 454822 131498 490586 131734
rect 490822 131498 526586 131734
rect 526822 131498 562586 131734
rect 562822 131498 588322 131734
rect 588558 131498 588740 131734
rect -4816 131476 588740 131498
rect -4816 131474 -4216 131476
rect 22404 131474 23004 131476
rect 58404 131474 59004 131476
rect 94404 131474 95004 131476
rect 130404 131474 131004 131476
rect 166404 131474 167004 131476
rect 202404 131474 203004 131476
rect 238404 131474 239004 131476
rect 274404 131474 275004 131476
rect 310404 131474 311004 131476
rect 346404 131474 347004 131476
rect 382404 131474 383004 131476
rect 418404 131474 419004 131476
rect 454404 131474 455004 131476
rect 490404 131474 491004 131476
rect 526404 131474 527004 131476
rect 562404 131474 563004 131476
rect 588140 131474 588740 131476
rect -2936 128476 -2336 128478
rect 18804 128476 19404 128478
rect 54804 128476 55404 128478
rect 90804 128476 91404 128478
rect 126804 128476 127404 128478
rect 162804 128476 163404 128478
rect 198804 128476 199404 128478
rect 234804 128476 235404 128478
rect 270804 128476 271404 128478
rect 306804 128476 307404 128478
rect 342804 128476 343404 128478
rect 378804 128476 379404 128478
rect 414804 128476 415404 128478
rect 450804 128476 451404 128478
rect 486804 128476 487404 128478
rect 522804 128476 523404 128478
rect 558804 128476 559404 128478
rect 586260 128476 586860 128478
rect -2936 128454 586860 128476
rect -2936 128218 -2754 128454
rect -2518 128218 18986 128454
rect 19222 128218 54986 128454
rect 55222 128218 90986 128454
rect 91222 128218 126986 128454
rect 127222 128218 162986 128454
rect 163222 128218 198986 128454
rect 199222 128218 234986 128454
rect 235222 128218 270986 128454
rect 271222 128218 306986 128454
rect 307222 128218 342986 128454
rect 343222 128218 378986 128454
rect 379222 128218 414986 128454
rect 415222 128218 450986 128454
rect 451222 128218 486986 128454
rect 487222 128218 522986 128454
rect 523222 128218 558986 128454
rect 559222 128218 586442 128454
rect 586678 128218 586860 128454
rect -2936 128134 586860 128218
rect -2936 127898 -2754 128134
rect -2518 127898 18986 128134
rect 19222 127898 54986 128134
rect 55222 127898 90986 128134
rect 91222 127898 126986 128134
rect 127222 127898 162986 128134
rect 163222 127898 198986 128134
rect 199222 127898 234986 128134
rect 235222 127898 270986 128134
rect 271222 127898 306986 128134
rect 307222 127898 342986 128134
rect 343222 127898 378986 128134
rect 379222 127898 414986 128134
rect 415222 127898 450986 128134
rect 451222 127898 486986 128134
rect 487222 127898 522986 128134
rect 523222 127898 558986 128134
rect 559222 127898 586442 128134
rect 586678 127898 586860 128134
rect -2936 127876 586860 127898
rect -2936 127874 -2336 127876
rect 18804 127874 19404 127876
rect 54804 127874 55404 127876
rect 90804 127874 91404 127876
rect 126804 127874 127404 127876
rect 162804 127874 163404 127876
rect 198804 127874 199404 127876
rect 234804 127874 235404 127876
rect 270804 127874 271404 127876
rect 306804 127874 307404 127876
rect 342804 127874 343404 127876
rect 378804 127874 379404 127876
rect 414804 127874 415404 127876
rect 450804 127874 451404 127876
rect 486804 127874 487404 127876
rect 522804 127874 523404 127876
rect 558804 127874 559404 127876
rect 586260 127874 586860 127876
rect -7636 121276 -7036 121278
rect 11604 121276 12204 121278
rect 47604 121276 48204 121278
rect 83604 121276 84204 121278
rect 119604 121276 120204 121278
rect 155604 121276 156204 121278
rect 191604 121276 192204 121278
rect 227604 121276 228204 121278
rect 263604 121276 264204 121278
rect 299604 121276 300204 121278
rect 335604 121276 336204 121278
rect 371604 121276 372204 121278
rect 407604 121276 408204 121278
rect 443604 121276 444204 121278
rect 479604 121276 480204 121278
rect 515604 121276 516204 121278
rect 551604 121276 552204 121278
rect 590960 121276 591560 121278
rect -8576 121254 592500 121276
rect -8576 121018 -7454 121254
rect -7218 121018 11786 121254
rect 12022 121018 47786 121254
rect 48022 121018 83786 121254
rect 84022 121018 119786 121254
rect 120022 121018 155786 121254
rect 156022 121018 191786 121254
rect 192022 121018 227786 121254
rect 228022 121018 263786 121254
rect 264022 121018 299786 121254
rect 300022 121018 335786 121254
rect 336022 121018 371786 121254
rect 372022 121018 407786 121254
rect 408022 121018 443786 121254
rect 444022 121018 479786 121254
rect 480022 121018 515786 121254
rect 516022 121018 551786 121254
rect 552022 121018 591142 121254
rect 591378 121018 592500 121254
rect -8576 120934 592500 121018
rect -8576 120698 -7454 120934
rect -7218 120698 11786 120934
rect 12022 120698 47786 120934
rect 48022 120698 83786 120934
rect 84022 120698 119786 120934
rect 120022 120698 155786 120934
rect 156022 120698 191786 120934
rect 192022 120698 227786 120934
rect 228022 120698 263786 120934
rect 264022 120698 299786 120934
rect 300022 120698 335786 120934
rect 336022 120698 371786 120934
rect 372022 120698 407786 120934
rect 408022 120698 443786 120934
rect 444022 120698 479786 120934
rect 480022 120698 515786 120934
rect 516022 120698 551786 120934
rect 552022 120698 591142 120934
rect 591378 120698 592500 120934
rect -8576 120676 592500 120698
rect -7636 120674 -7036 120676
rect 11604 120674 12204 120676
rect 47604 120674 48204 120676
rect 83604 120674 84204 120676
rect 119604 120674 120204 120676
rect 155604 120674 156204 120676
rect 191604 120674 192204 120676
rect 227604 120674 228204 120676
rect 263604 120674 264204 120676
rect 299604 120674 300204 120676
rect 335604 120674 336204 120676
rect 371604 120674 372204 120676
rect 407604 120674 408204 120676
rect 443604 120674 444204 120676
rect 479604 120674 480204 120676
rect 515604 120674 516204 120676
rect 551604 120674 552204 120676
rect 590960 120674 591560 120676
rect -5756 117676 -5156 117678
rect 8004 117676 8604 117678
rect 44004 117676 44604 117678
rect 80004 117676 80604 117678
rect 116004 117676 116604 117678
rect 152004 117676 152604 117678
rect 188004 117676 188604 117678
rect 224004 117676 224604 117678
rect 260004 117676 260604 117678
rect 296004 117676 296604 117678
rect 332004 117676 332604 117678
rect 368004 117676 368604 117678
rect 404004 117676 404604 117678
rect 440004 117676 440604 117678
rect 476004 117676 476604 117678
rect 512004 117676 512604 117678
rect 548004 117676 548604 117678
rect 589080 117676 589680 117678
rect -6696 117654 590620 117676
rect -6696 117418 -5574 117654
rect -5338 117418 8186 117654
rect 8422 117418 44186 117654
rect 44422 117418 80186 117654
rect 80422 117418 116186 117654
rect 116422 117418 152186 117654
rect 152422 117418 188186 117654
rect 188422 117418 224186 117654
rect 224422 117418 260186 117654
rect 260422 117418 296186 117654
rect 296422 117418 332186 117654
rect 332422 117418 368186 117654
rect 368422 117418 404186 117654
rect 404422 117418 440186 117654
rect 440422 117418 476186 117654
rect 476422 117418 512186 117654
rect 512422 117418 548186 117654
rect 548422 117418 589262 117654
rect 589498 117418 590620 117654
rect -6696 117334 590620 117418
rect -6696 117098 -5574 117334
rect -5338 117098 8186 117334
rect 8422 117098 44186 117334
rect 44422 117098 80186 117334
rect 80422 117098 116186 117334
rect 116422 117098 152186 117334
rect 152422 117098 188186 117334
rect 188422 117098 224186 117334
rect 224422 117098 260186 117334
rect 260422 117098 296186 117334
rect 296422 117098 332186 117334
rect 332422 117098 368186 117334
rect 368422 117098 404186 117334
rect 404422 117098 440186 117334
rect 440422 117098 476186 117334
rect 476422 117098 512186 117334
rect 512422 117098 548186 117334
rect 548422 117098 589262 117334
rect 589498 117098 590620 117334
rect -6696 117076 590620 117098
rect -5756 117074 -5156 117076
rect 8004 117074 8604 117076
rect 44004 117074 44604 117076
rect 80004 117074 80604 117076
rect 116004 117074 116604 117076
rect 152004 117074 152604 117076
rect 188004 117074 188604 117076
rect 224004 117074 224604 117076
rect 260004 117074 260604 117076
rect 296004 117074 296604 117076
rect 332004 117074 332604 117076
rect 368004 117074 368604 117076
rect 404004 117074 404604 117076
rect 440004 117074 440604 117076
rect 476004 117074 476604 117076
rect 512004 117074 512604 117076
rect 548004 117074 548604 117076
rect 589080 117074 589680 117076
rect -3876 114076 -3276 114078
rect 4404 114076 5004 114078
rect 40404 114076 41004 114078
rect 76404 114076 77004 114078
rect 112404 114076 113004 114078
rect 148404 114076 149004 114078
rect 184404 114076 185004 114078
rect 220404 114076 221004 114078
rect 256404 114076 257004 114078
rect 292404 114076 293004 114078
rect 328404 114076 329004 114078
rect 364404 114076 365004 114078
rect 400404 114076 401004 114078
rect 436404 114076 437004 114078
rect 472404 114076 473004 114078
rect 508404 114076 509004 114078
rect 544404 114076 545004 114078
rect 580404 114076 581004 114078
rect 587200 114076 587800 114078
rect -4816 114054 588740 114076
rect -4816 113818 -3694 114054
rect -3458 113818 4586 114054
rect 4822 113818 40586 114054
rect 40822 113818 76586 114054
rect 76822 113818 112586 114054
rect 112822 113818 148586 114054
rect 148822 113818 184586 114054
rect 184822 113818 220586 114054
rect 220822 113818 256586 114054
rect 256822 113818 292586 114054
rect 292822 113818 328586 114054
rect 328822 113818 364586 114054
rect 364822 113818 400586 114054
rect 400822 113818 436586 114054
rect 436822 113818 472586 114054
rect 472822 113818 508586 114054
rect 508822 113818 544586 114054
rect 544822 113818 580586 114054
rect 580822 113818 587382 114054
rect 587618 113818 588740 114054
rect -4816 113734 588740 113818
rect -4816 113498 -3694 113734
rect -3458 113498 4586 113734
rect 4822 113498 40586 113734
rect 40822 113498 76586 113734
rect 76822 113498 112586 113734
rect 112822 113498 148586 113734
rect 148822 113498 184586 113734
rect 184822 113498 220586 113734
rect 220822 113498 256586 113734
rect 256822 113498 292586 113734
rect 292822 113498 328586 113734
rect 328822 113498 364586 113734
rect 364822 113498 400586 113734
rect 400822 113498 436586 113734
rect 436822 113498 472586 113734
rect 472822 113498 508586 113734
rect 508822 113498 544586 113734
rect 544822 113498 580586 113734
rect 580822 113498 587382 113734
rect 587618 113498 588740 113734
rect -4816 113476 588740 113498
rect -3876 113474 -3276 113476
rect 4404 113474 5004 113476
rect 40404 113474 41004 113476
rect 76404 113474 77004 113476
rect 112404 113474 113004 113476
rect 148404 113474 149004 113476
rect 184404 113474 185004 113476
rect 220404 113474 221004 113476
rect 256404 113474 257004 113476
rect 292404 113474 293004 113476
rect 328404 113474 329004 113476
rect 364404 113474 365004 113476
rect 400404 113474 401004 113476
rect 436404 113474 437004 113476
rect 472404 113474 473004 113476
rect 508404 113474 509004 113476
rect 544404 113474 545004 113476
rect 580404 113474 581004 113476
rect 587200 113474 587800 113476
rect -1996 110476 -1396 110478
rect 804 110476 1404 110478
rect 36804 110476 37404 110478
rect 72804 110476 73404 110478
rect 108804 110476 109404 110478
rect 144804 110476 145404 110478
rect 180804 110476 181404 110478
rect 216804 110476 217404 110478
rect 252804 110476 253404 110478
rect 288804 110476 289404 110478
rect 324804 110476 325404 110478
rect 360804 110476 361404 110478
rect 396804 110476 397404 110478
rect 432804 110476 433404 110478
rect 468804 110476 469404 110478
rect 504804 110476 505404 110478
rect 540804 110476 541404 110478
rect 576804 110476 577404 110478
rect 585320 110476 585920 110478
rect -2936 110454 586860 110476
rect -2936 110218 -1814 110454
rect -1578 110218 986 110454
rect 1222 110218 36986 110454
rect 37222 110218 72986 110454
rect 73222 110218 108986 110454
rect 109222 110218 144986 110454
rect 145222 110218 180986 110454
rect 181222 110218 216986 110454
rect 217222 110218 252986 110454
rect 253222 110218 288986 110454
rect 289222 110218 324986 110454
rect 325222 110218 360986 110454
rect 361222 110218 396986 110454
rect 397222 110218 432986 110454
rect 433222 110218 468986 110454
rect 469222 110218 504986 110454
rect 505222 110218 540986 110454
rect 541222 110218 576986 110454
rect 577222 110218 585502 110454
rect 585738 110218 586860 110454
rect -2936 110134 586860 110218
rect -2936 109898 -1814 110134
rect -1578 109898 986 110134
rect 1222 109898 36986 110134
rect 37222 109898 72986 110134
rect 73222 109898 108986 110134
rect 109222 109898 144986 110134
rect 145222 109898 180986 110134
rect 181222 109898 216986 110134
rect 217222 109898 252986 110134
rect 253222 109898 288986 110134
rect 289222 109898 324986 110134
rect 325222 109898 360986 110134
rect 361222 109898 396986 110134
rect 397222 109898 432986 110134
rect 433222 109898 468986 110134
rect 469222 109898 504986 110134
rect 505222 109898 540986 110134
rect 541222 109898 576986 110134
rect 577222 109898 585502 110134
rect 585738 109898 586860 110134
rect -2936 109876 586860 109898
rect -1996 109874 -1396 109876
rect 804 109874 1404 109876
rect 36804 109874 37404 109876
rect 72804 109874 73404 109876
rect 108804 109874 109404 109876
rect 144804 109874 145404 109876
rect 180804 109874 181404 109876
rect 216804 109874 217404 109876
rect 252804 109874 253404 109876
rect 288804 109874 289404 109876
rect 324804 109874 325404 109876
rect 360804 109874 361404 109876
rect 396804 109874 397404 109876
rect 432804 109874 433404 109876
rect 468804 109874 469404 109876
rect 504804 109874 505404 109876
rect 540804 109874 541404 109876
rect 576804 109874 577404 109876
rect 585320 109874 585920 109876
rect -8576 103276 -7976 103278
rect 29604 103276 30204 103278
rect 65604 103276 66204 103278
rect 101604 103276 102204 103278
rect 137604 103276 138204 103278
rect 173604 103276 174204 103278
rect 209604 103276 210204 103278
rect 245604 103276 246204 103278
rect 281604 103276 282204 103278
rect 317604 103276 318204 103278
rect 353604 103276 354204 103278
rect 389604 103276 390204 103278
rect 425604 103276 426204 103278
rect 461604 103276 462204 103278
rect 497604 103276 498204 103278
rect 533604 103276 534204 103278
rect 569604 103276 570204 103278
rect 591900 103276 592500 103278
rect -8576 103254 592500 103276
rect -8576 103018 -8394 103254
rect -8158 103018 29786 103254
rect 30022 103018 65786 103254
rect 66022 103018 101786 103254
rect 102022 103018 137786 103254
rect 138022 103018 173786 103254
rect 174022 103018 209786 103254
rect 210022 103018 245786 103254
rect 246022 103018 281786 103254
rect 282022 103018 317786 103254
rect 318022 103018 353786 103254
rect 354022 103018 389786 103254
rect 390022 103018 425786 103254
rect 426022 103018 461786 103254
rect 462022 103018 497786 103254
rect 498022 103018 533786 103254
rect 534022 103018 569786 103254
rect 570022 103018 592082 103254
rect 592318 103018 592500 103254
rect -8576 102934 592500 103018
rect -8576 102698 -8394 102934
rect -8158 102698 29786 102934
rect 30022 102698 65786 102934
rect 66022 102698 101786 102934
rect 102022 102698 137786 102934
rect 138022 102698 173786 102934
rect 174022 102698 209786 102934
rect 210022 102698 245786 102934
rect 246022 102698 281786 102934
rect 282022 102698 317786 102934
rect 318022 102698 353786 102934
rect 354022 102698 389786 102934
rect 390022 102698 425786 102934
rect 426022 102698 461786 102934
rect 462022 102698 497786 102934
rect 498022 102698 533786 102934
rect 534022 102698 569786 102934
rect 570022 102698 592082 102934
rect 592318 102698 592500 102934
rect -8576 102676 592500 102698
rect -8576 102674 -7976 102676
rect 29604 102674 30204 102676
rect 65604 102674 66204 102676
rect 101604 102674 102204 102676
rect 137604 102674 138204 102676
rect 173604 102674 174204 102676
rect 209604 102674 210204 102676
rect 245604 102674 246204 102676
rect 281604 102674 282204 102676
rect 317604 102674 318204 102676
rect 353604 102674 354204 102676
rect 389604 102674 390204 102676
rect 425604 102674 426204 102676
rect 461604 102674 462204 102676
rect 497604 102674 498204 102676
rect 533604 102674 534204 102676
rect 569604 102674 570204 102676
rect 591900 102674 592500 102676
rect -6696 99676 -6096 99678
rect 26004 99676 26604 99678
rect 62004 99676 62604 99678
rect 98004 99676 98604 99678
rect 134004 99676 134604 99678
rect 170004 99676 170604 99678
rect 206004 99676 206604 99678
rect 242004 99676 242604 99678
rect 278004 99676 278604 99678
rect 314004 99676 314604 99678
rect 350004 99676 350604 99678
rect 386004 99676 386604 99678
rect 422004 99676 422604 99678
rect 458004 99676 458604 99678
rect 494004 99676 494604 99678
rect 530004 99676 530604 99678
rect 566004 99676 566604 99678
rect 590020 99676 590620 99678
rect -6696 99654 590620 99676
rect -6696 99418 -6514 99654
rect -6278 99418 26186 99654
rect 26422 99418 62186 99654
rect 62422 99418 98186 99654
rect 98422 99418 134186 99654
rect 134422 99418 170186 99654
rect 170422 99418 206186 99654
rect 206422 99418 242186 99654
rect 242422 99418 278186 99654
rect 278422 99418 314186 99654
rect 314422 99418 350186 99654
rect 350422 99418 386186 99654
rect 386422 99418 422186 99654
rect 422422 99418 458186 99654
rect 458422 99418 494186 99654
rect 494422 99418 530186 99654
rect 530422 99418 566186 99654
rect 566422 99418 590202 99654
rect 590438 99418 590620 99654
rect -6696 99334 590620 99418
rect -6696 99098 -6514 99334
rect -6278 99098 26186 99334
rect 26422 99098 62186 99334
rect 62422 99098 98186 99334
rect 98422 99098 134186 99334
rect 134422 99098 170186 99334
rect 170422 99098 206186 99334
rect 206422 99098 242186 99334
rect 242422 99098 278186 99334
rect 278422 99098 314186 99334
rect 314422 99098 350186 99334
rect 350422 99098 386186 99334
rect 386422 99098 422186 99334
rect 422422 99098 458186 99334
rect 458422 99098 494186 99334
rect 494422 99098 530186 99334
rect 530422 99098 566186 99334
rect 566422 99098 590202 99334
rect 590438 99098 590620 99334
rect -6696 99076 590620 99098
rect -6696 99074 -6096 99076
rect 26004 99074 26604 99076
rect 62004 99074 62604 99076
rect 98004 99074 98604 99076
rect 134004 99074 134604 99076
rect 170004 99074 170604 99076
rect 206004 99074 206604 99076
rect 242004 99074 242604 99076
rect 278004 99074 278604 99076
rect 314004 99074 314604 99076
rect 350004 99074 350604 99076
rect 386004 99074 386604 99076
rect 422004 99074 422604 99076
rect 458004 99074 458604 99076
rect 494004 99074 494604 99076
rect 530004 99074 530604 99076
rect 566004 99074 566604 99076
rect 590020 99074 590620 99076
rect -4816 96076 -4216 96078
rect 22404 96076 23004 96078
rect 58404 96076 59004 96078
rect 94404 96076 95004 96078
rect 130404 96076 131004 96078
rect 166404 96076 167004 96078
rect 202404 96076 203004 96078
rect 238404 96076 239004 96078
rect 274404 96076 275004 96078
rect 310404 96076 311004 96078
rect 346404 96076 347004 96078
rect 382404 96076 383004 96078
rect 418404 96076 419004 96078
rect 454404 96076 455004 96078
rect 490404 96076 491004 96078
rect 526404 96076 527004 96078
rect 562404 96076 563004 96078
rect 588140 96076 588740 96078
rect -4816 96054 588740 96076
rect -4816 95818 -4634 96054
rect -4398 95818 22586 96054
rect 22822 95818 58586 96054
rect 58822 95818 94586 96054
rect 94822 95818 130586 96054
rect 130822 95818 166586 96054
rect 166822 95818 202586 96054
rect 202822 95818 238586 96054
rect 238822 95818 274586 96054
rect 274822 95818 310586 96054
rect 310822 95818 346586 96054
rect 346822 95818 382586 96054
rect 382822 95818 418586 96054
rect 418822 95818 454586 96054
rect 454822 95818 490586 96054
rect 490822 95818 526586 96054
rect 526822 95818 562586 96054
rect 562822 95818 588322 96054
rect 588558 95818 588740 96054
rect -4816 95734 588740 95818
rect -4816 95498 -4634 95734
rect -4398 95498 22586 95734
rect 22822 95498 58586 95734
rect 58822 95498 94586 95734
rect 94822 95498 130586 95734
rect 130822 95498 166586 95734
rect 166822 95498 202586 95734
rect 202822 95498 238586 95734
rect 238822 95498 274586 95734
rect 274822 95498 310586 95734
rect 310822 95498 346586 95734
rect 346822 95498 382586 95734
rect 382822 95498 418586 95734
rect 418822 95498 454586 95734
rect 454822 95498 490586 95734
rect 490822 95498 526586 95734
rect 526822 95498 562586 95734
rect 562822 95498 588322 95734
rect 588558 95498 588740 95734
rect -4816 95476 588740 95498
rect -4816 95474 -4216 95476
rect 22404 95474 23004 95476
rect 58404 95474 59004 95476
rect 94404 95474 95004 95476
rect 130404 95474 131004 95476
rect 166404 95474 167004 95476
rect 202404 95474 203004 95476
rect 238404 95474 239004 95476
rect 274404 95474 275004 95476
rect 310404 95474 311004 95476
rect 346404 95474 347004 95476
rect 382404 95474 383004 95476
rect 418404 95474 419004 95476
rect 454404 95474 455004 95476
rect 490404 95474 491004 95476
rect 526404 95474 527004 95476
rect 562404 95474 563004 95476
rect 588140 95474 588740 95476
rect -2936 92476 -2336 92478
rect 18804 92476 19404 92478
rect 54804 92476 55404 92478
rect 90804 92476 91404 92478
rect 126804 92476 127404 92478
rect 162804 92476 163404 92478
rect 198804 92476 199404 92478
rect 234804 92476 235404 92478
rect 270804 92476 271404 92478
rect 306804 92476 307404 92478
rect 342804 92476 343404 92478
rect 378804 92476 379404 92478
rect 414804 92476 415404 92478
rect 450804 92476 451404 92478
rect 486804 92476 487404 92478
rect 522804 92476 523404 92478
rect 558804 92476 559404 92478
rect 586260 92476 586860 92478
rect -2936 92454 586860 92476
rect -2936 92218 -2754 92454
rect -2518 92218 18986 92454
rect 19222 92218 54986 92454
rect 55222 92218 90986 92454
rect 91222 92218 126986 92454
rect 127222 92218 162986 92454
rect 163222 92218 198986 92454
rect 199222 92218 234986 92454
rect 235222 92218 270986 92454
rect 271222 92218 306986 92454
rect 307222 92218 342986 92454
rect 343222 92218 378986 92454
rect 379222 92218 414986 92454
rect 415222 92218 450986 92454
rect 451222 92218 486986 92454
rect 487222 92218 522986 92454
rect 523222 92218 558986 92454
rect 559222 92218 586442 92454
rect 586678 92218 586860 92454
rect -2936 92134 586860 92218
rect -2936 91898 -2754 92134
rect -2518 91898 18986 92134
rect 19222 91898 54986 92134
rect 55222 91898 90986 92134
rect 91222 91898 126986 92134
rect 127222 91898 162986 92134
rect 163222 91898 198986 92134
rect 199222 91898 234986 92134
rect 235222 91898 270986 92134
rect 271222 91898 306986 92134
rect 307222 91898 342986 92134
rect 343222 91898 378986 92134
rect 379222 91898 414986 92134
rect 415222 91898 450986 92134
rect 451222 91898 486986 92134
rect 487222 91898 522986 92134
rect 523222 91898 558986 92134
rect 559222 91898 586442 92134
rect 586678 91898 586860 92134
rect -2936 91876 586860 91898
rect -2936 91874 -2336 91876
rect 18804 91874 19404 91876
rect 54804 91874 55404 91876
rect 90804 91874 91404 91876
rect 126804 91874 127404 91876
rect 162804 91874 163404 91876
rect 198804 91874 199404 91876
rect 234804 91874 235404 91876
rect 270804 91874 271404 91876
rect 306804 91874 307404 91876
rect 342804 91874 343404 91876
rect 378804 91874 379404 91876
rect 414804 91874 415404 91876
rect 450804 91874 451404 91876
rect 486804 91874 487404 91876
rect 522804 91874 523404 91876
rect 558804 91874 559404 91876
rect 586260 91874 586860 91876
rect -7636 85276 -7036 85278
rect 11604 85276 12204 85278
rect 47604 85276 48204 85278
rect 83604 85276 84204 85278
rect 119604 85276 120204 85278
rect 155604 85276 156204 85278
rect 191604 85276 192204 85278
rect 227604 85276 228204 85278
rect 263604 85276 264204 85278
rect 299604 85276 300204 85278
rect 335604 85276 336204 85278
rect 371604 85276 372204 85278
rect 407604 85276 408204 85278
rect 443604 85276 444204 85278
rect 479604 85276 480204 85278
rect 515604 85276 516204 85278
rect 551604 85276 552204 85278
rect 590960 85276 591560 85278
rect -8576 85254 592500 85276
rect -8576 85018 -7454 85254
rect -7218 85018 11786 85254
rect 12022 85018 47786 85254
rect 48022 85018 83786 85254
rect 84022 85018 119786 85254
rect 120022 85018 155786 85254
rect 156022 85018 191786 85254
rect 192022 85018 227786 85254
rect 228022 85018 263786 85254
rect 264022 85018 299786 85254
rect 300022 85018 335786 85254
rect 336022 85018 371786 85254
rect 372022 85018 407786 85254
rect 408022 85018 443786 85254
rect 444022 85018 479786 85254
rect 480022 85018 515786 85254
rect 516022 85018 551786 85254
rect 552022 85018 591142 85254
rect 591378 85018 592500 85254
rect -8576 84934 592500 85018
rect -8576 84698 -7454 84934
rect -7218 84698 11786 84934
rect 12022 84698 47786 84934
rect 48022 84698 83786 84934
rect 84022 84698 119786 84934
rect 120022 84698 155786 84934
rect 156022 84698 191786 84934
rect 192022 84698 227786 84934
rect 228022 84698 263786 84934
rect 264022 84698 299786 84934
rect 300022 84698 335786 84934
rect 336022 84698 371786 84934
rect 372022 84698 407786 84934
rect 408022 84698 443786 84934
rect 444022 84698 479786 84934
rect 480022 84698 515786 84934
rect 516022 84698 551786 84934
rect 552022 84698 591142 84934
rect 591378 84698 592500 84934
rect -8576 84676 592500 84698
rect -7636 84674 -7036 84676
rect 11604 84674 12204 84676
rect 47604 84674 48204 84676
rect 83604 84674 84204 84676
rect 119604 84674 120204 84676
rect 155604 84674 156204 84676
rect 191604 84674 192204 84676
rect 227604 84674 228204 84676
rect 263604 84674 264204 84676
rect 299604 84674 300204 84676
rect 335604 84674 336204 84676
rect 371604 84674 372204 84676
rect 407604 84674 408204 84676
rect 443604 84674 444204 84676
rect 479604 84674 480204 84676
rect 515604 84674 516204 84676
rect 551604 84674 552204 84676
rect 590960 84674 591560 84676
rect -5756 81676 -5156 81678
rect 8004 81676 8604 81678
rect 44004 81676 44604 81678
rect 80004 81676 80604 81678
rect 116004 81676 116604 81678
rect 152004 81676 152604 81678
rect 188004 81676 188604 81678
rect 224004 81676 224604 81678
rect 260004 81676 260604 81678
rect 296004 81676 296604 81678
rect 332004 81676 332604 81678
rect 368004 81676 368604 81678
rect 404004 81676 404604 81678
rect 440004 81676 440604 81678
rect 476004 81676 476604 81678
rect 512004 81676 512604 81678
rect 548004 81676 548604 81678
rect 589080 81676 589680 81678
rect -6696 81654 590620 81676
rect -6696 81418 -5574 81654
rect -5338 81418 8186 81654
rect 8422 81418 44186 81654
rect 44422 81418 80186 81654
rect 80422 81418 116186 81654
rect 116422 81418 152186 81654
rect 152422 81418 188186 81654
rect 188422 81418 224186 81654
rect 224422 81418 260186 81654
rect 260422 81418 296186 81654
rect 296422 81418 332186 81654
rect 332422 81418 368186 81654
rect 368422 81418 404186 81654
rect 404422 81418 440186 81654
rect 440422 81418 476186 81654
rect 476422 81418 512186 81654
rect 512422 81418 548186 81654
rect 548422 81418 589262 81654
rect 589498 81418 590620 81654
rect -6696 81334 590620 81418
rect -6696 81098 -5574 81334
rect -5338 81098 8186 81334
rect 8422 81098 44186 81334
rect 44422 81098 80186 81334
rect 80422 81098 116186 81334
rect 116422 81098 152186 81334
rect 152422 81098 188186 81334
rect 188422 81098 224186 81334
rect 224422 81098 260186 81334
rect 260422 81098 296186 81334
rect 296422 81098 332186 81334
rect 332422 81098 368186 81334
rect 368422 81098 404186 81334
rect 404422 81098 440186 81334
rect 440422 81098 476186 81334
rect 476422 81098 512186 81334
rect 512422 81098 548186 81334
rect 548422 81098 589262 81334
rect 589498 81098 590620 81334
rect -6696 81076 590620 81098
rect -5756 81074 -5156 81076
rect 8004 81074 8604 81076
rect 44004 81074 44604 81076
rect 80004 81074 80604 81076
rect 116004 81074 116604 81076
rect 152004 81074 152604 81076
rect 188004 81074 188604 81076
rect 224004 81074 224604 81076
rect 260004 81074 260604 81076
rect 296004 81074 296604 81076
rect 332004 81074 332604 81076
rect 368004 81074 368604 81076
rect 404004 81074 404604 81076
rect 440004 81074 440604 81076
rect 476004 81074 476604 81076
rect 512004 81074 512604 81076
rect 548004 81074 548604 81076
rect 589080 81074 589680 81076
rect -3876 78076 -3276 78078
rect 4404 78076 5004 78078
rect 40404 78076 41004 78078
rect 76404 78076 77004 78078
rect 112404 78076 113004 78078
rect 148404 78076 149004 78078
rect 184404 78076 185004 78078
rect 220404 78076 221004 78078
rect 256404 78076 257004 78078
rect 292404 78076 293004 78078
rect 328404 78076 329004 78078
rect 364404 78076 365004 78078
rect 400404 78076 401004 78078
rect 436404 78076 437004 78078
rect 472404 78076 473004 78078
rect 508404 78076 509004 78078
rect 544404 78076 545004 78078
rect 580404 78076 581004 78078
rect 587200 78076 587800 78078
rect -4816 78054 588740 78076
rect -4816 77818 -3694 78054
rect -3458 77818 4586 78054
rect 4822 77818 40586 78054
rect 40822 77818 76586 78054
rect 76822 77818 112586 78054
rect 112822 77818 148586 78054
rect 148822 77818 184586 78054
rect 184822 77818 220586 78054
rect 220822 77818 256586 78054
rect 256822 77818 292586 78054
rect 292822 77818 328586 78054
rect 328822 77818 364586 78054
rect 364822 77818 400586 78054
rect 400822 77818 436586 78054
rect 436822 77818 472586 78054
rect 472822 77818 508586 78054
rect 508822 77818 544586 78054
rect 544822 77818 580586 78054
rect 580822 77818 587382 78054
rect 587618 77818 588740 78054
rect -4816 77734 588740 77818
rect -4816 77498 -3694 77734
rect -3458 77498 4586 77734
rect 4822 77498 40586 77734
rect 40822 77498 76586 77734
rect 76822 77498 112586 77734
rect 112822 77498 148586 77734
rect 148822 77498 184586 77734
rect 184822 77498 220586 77734
rect 220822 77498 256586 77734
rect 256822 77498 292586 77734
rect 292822 77498 328586 77734
rect 328822 77498 364586 77734
rect 364822 77498 400586 77734
rect 400822 77498 436586 77734
rect 436822 77498 472586 77734
rect 472822 77498 508586 77734
rect 508822 77498 544586 77734
rect 544822 77498 580586 77734
rect 580822 77498 587382 77734
rect 587618 77498 588740 77734
rect -4816 77476 588740 77498
rect -3876 77474 -3276 77476
rect 4404 77474 5004 77476
rect 40404 77474 41004 77476
rect 76404 77474 77004 77476
rect 112404 77474 113004 77476
rect 148404 77474 149004 77476
rect 184404 77474 185004 77476
rect 220404 77474 221004 77476
rect 256404 77474 257004 77476
rect 292404 77474 293004 77476
rect 328404 77474 329004 77476
rect 364404 77474 365004 77476
rect 400404 77474 401004 77476
rect 436404 77474 437004 77476
rect 472404 77474 473004 77476
rect 508404 77474 509004 77476
rect 544404 77474 545004 77476
rect 580404 77474 581004 77476
rect 587200 77474 587800 77476
rect -1996 74476 -1396 74478
rect 804 74476 1404 74478
rect 36804 74476 37404 74478
rect 72804 74476 73404 74478
rect 108804 74476 109404 74478
rect 144804 74476 145404 74478
rect 180804 74476 181404 74478
rect 216804 74476 217404 74478
rect 252804 74476 253404 74478
rect 288804 74476 289404 74478
rect 324804 74476 325404 74478
rect 360804 74476 361404 74478
rect 396804 74476 397404 74478
rect 432804 74476 433404 74478
rect 468804 74476 469404 74478
rect 504804 74476 505404 74478
rect 540804 74476 541404 74478
rect 576804 74476 577404 74478
rect 585320 74476 585920 74478
rect -2936 74454 586860 74476
rect -2936 74218 -1814 74454
rect -1578 74218 986 74454
rect 1222 74218 36986 74454
rect 37222 74218 72986 74454
rect 73222 74218 108986 74454
rect 109222 74218 144986 74454
rect 145222 74218 180986 74454
rect 181222 74218 216986 74454
rect 217222 74218 252986 74454
rect 253222 74218 288986 74454
rect 289222 74218 324986 74454
rect 325222 74218 360986 74454
rect 361222 74218 396986 74454
rect 397222 74218 432986 74454
rect 433222 74218 468986 74454
rect 469222 74218 504986 74454
rect 505222 74218 540986 74454
rect 541222 74218 576986 74454
rect 577222 74218 585502 74454
rect 585738 74218 586860 74454
rect -2936 74134 586860 74218
rect -2936 73898 -1814 74134
rect -1578 73898 986 74134
rect 1222 73898 36986 74134
rect 37222 73898 72986 74134
rect 73222 73898 108986 74134
rect 109222 73898 144986 74134
rect 145222 73898 180986 74134
rect 181222 73898 216986 74134
rect 217222 73898 252986 74134
rect 253222 73898 288986 74134
rect 289222 73898 324986 74134
rect 325222 73898 360986 74134
rect 361222 73898 396986 74134
rect 397222 73898 432986 74134
rect 433222 73898 468986 74134
rect 469222 73898 504986 74134
rect 505222 73898 540986 74134
rect 541222 73898 576986 74134
rect 577222 73898 585502 74134
rect 585738 73898 586860 74134
rect -2936 73876 586860 73898
rect -1996 73874 -1396 73876
rect 804 73874 1404 73876
rect 36804 73874 37404 73876
rect 72804 73874 73404 73876
rect 108804 73874 109404 73876
rect 144804 73874 145404 73876
rect 180804 73874 181404 73876
rect 216804 73874 217404 73876
rect 252804 73874 253404 73876
rect 288804 73874 289404 73876
rect 324804 73874 325404 73876
rect 360804 73874 361404 73876
rect 396804 73874 397404 73876
rect 432804 73874 433404 73876
rect 468804 73874 469404 73876
rect 504804 73874 505404 73876
rect 540804 73874 541404 73876
rect 576804 73874 577404 73876
rect 585320 73874 585920 73876
rect -8576 67276 -7976 67278
rect 29604 67276 30204 67278
rect 65604 67276 66204 67278
rect 101604 67276 102204 67278
rect 137604 67276 138204 67278
rect 173604 67276 174204 67278
rect 209604 67276 210204 67278
rect 245604 67276 246204 67278
rect 281604 67276 282204 67278
rect 317604 67276 318204 67278
rect 353604 67276 354204 67278
rect 389604 67276 390204 67278
rect 425604 67276 426204 67278
rect 461604 67276 462204 67278
rect 497604 67276 498204 67278
rect 533604 67276 534204 67278
rect 569604 67276 570204 67278
rect 591900 67276 592500 67278
rect -8576 67254 592500 67276
rect -8576 67018 -8394 67254
rect -8158 67018 29786 67254
rect 30022 67018 65786 67254
rect 66022 67018 101786 67254
rect 102022 67018 137786 67254
rect 138022 67018 173786 67254
rect 174022 67018 209786 67254
rect 210022 67018 245786 67254
rect 246022 67018 281786 67254
rect 282022 67018 317786 67254
rect 318022 67018 353786 67254
rect 354022 67018 389786 67254
rect 390022 67018 425786 67254
rect 426022 67018 461786 67254
rect 462022 67018 497786 67254
rect 498022 67018 533786 67254
rect 534022 67018 569786 67254
rect 570022 67018 592082 67254
rect 592318 67018 592500 67254
rect -8576 66934 592500 67018
rect -8576 66698 -8394 66934
rect -8158 66698 29786 66934
rect 30022 66698 65786 66934
rect 66022 66698 101786 66934
rect 102022 66698 137786 66934
rect 138022 66698 173786 66934
rect 174022 66698 209786 66934
rect 210022 66698 245786 66934
rect 246022 66698 281786 66934
rect 282022 66698 317786 66934
rect 318022 66698 353786 66934
rect 354022 66698 389786 66934
rect 390022 66698 425786 66934
rect 426022 66698 461786 66934
rect 462022 66698 497786 66934
rect 498022 66698 533786 66934
rect 534022 66698 569786 66934
rect 570022 66698 592082 66934
rect 592318 66698 592500 66934
rect -8576 66676 592500 66698
rect -8576 66674 -7976 66676
rect 29604 66674 30204 66676
rect 65604 66674 66204 66676
rect 101604 66674 102204 66676
rect 137604 66674 138204 66676
rect 173604 66674 174204 66676
rect 209604 66674 210204 66676
rect 245604 66674 246204 66676
rect 281604 66674 282204 66676
rect 317604 66674 318204 66676
rect 353604 66674 354204 66676
rect 389604 66674 390204 66676
rect 425604 66674 426204 66676
rect 461604 66674 462204 66676
rect 497604 66674 498204 66676
rect 533604 66674 534204 66676
rect 569604 66674 570204 66676
rect 591900 66674 592500 66676
rect -6696 63676 -6096 63678
rect 26004 63676 26604 63678
rect 62004 63676 62604 63678
rect 98004 63676 98604 63678
rect 134004 63676 134604 63678
rect 170004 63676 170604 63678
rect 206004 63676 206604 63678
rect 242004 63676 242604 63678
rect 278004 63676 278604 63678
rect 314004 63676 314604 63678
rect 350004 63676 350604 63678
rect 386004 63676 386604 63678
rect 422004 63676 422604 63678
rect 458004 63676 458604 63678
rect 494004 63676 494604 63678
rect 530004 63676 530604 63678
rect 566004 63676 566604 63678
rect 590020 63676 590620 63678
rect -6696 63654 590620 63676
rect -6696 63418 -6514 63654
rect -6278 63418 26186 63654
rect 26422 63418 62186 63654
rect 62422 63418 98186 63654
rect 98422 63418 134186 63654
rect 134422 63418 170186 63654
rect 170422 63418 206186 63654
rect 206422 63418 242186 63654
rect 242422 63418 278186 63654
rect 278422 63418 314186 63654
rect 314422 63418 350186 63654
rect 350422 63418 386186 63654
rect 386422 63418 422186 63654
rect 422422 63418 458186 63654
rect 458422 63418 494186 63654
rect 494422 63418 530186 63654
rect 530422 63418 566186 63654
rect 566422 63418 590202 63654
rect 590438 63418 590620 63654
rect -6696 63334 590620 63418
rect -6696 63098 -6514 63334
rect -6278 63098 26186 63334
rect 26422 63098 62186 63334
rect 62422 63098 98186 63334
rect 98422 63098 134186 63334
rect 134422 63098 170186 63334
rect 170422 63098 206186 63334
rect 206422 63098 242186 63334
rect 242422 63098 278186 63334
rect 278422 63098 314186 63334
rect 314422 63098 350186 63334
rect 350422 63098 386186 63334
rect 386422 63098 422186 63334
rect 422422 63098 458186 63334
rect 458422 63098 494186 63334
rect 494422 63098 530186 63334
rect 530422 63098 566186 63334
rect 566422 63098 590202 63334
rect 590438 63098 590620 63334
rect -6696 63076 590620 63098
rect -6696 63074 -6096 63076
rect 26004 63074 26604 63076
rect 62004 63074 62604 63076
rect 98004 63074 98604 63076
rect 134004 63074 134604 63076
rect 170004 63074 170604 63076
rect 206004 63074 206604 63076
rect 242004 63074 242604 63076
rect 278004 63074 278604 63076
rect 314004 63074 314604 63076
rect 350004 63074 350604 63076
rect 386004 63074 386604 63076
rect 422004 63074 422604 63076
rect 458004 63074 458604 63076
rect 494004 63074 494604 63076
rect 530004 63074 530604 63076
rect 566004 63074 566604 63076
rect 590020 63074 590620 63076
rect -4816 60076 -4216 60078
rect 22404 60076 23004 60078
rect 58404 60076 59004 60078
rect 94404 60076 95004 60078
rect 130404 60076 131004 60078
rect 166404 60076 167004 60078
rect 202404 60076 203004 60078
rect 238404 60076 239004 60078
rect 274404 60076 275004 60078
rect 310404 60076 311004 60078
rect 346404 60076 347004 60078
rect 382404 60076 383004 60078
rect 418404 60076 419004 60078
rect 454404 60076 455004 60078
rect 490404 60076 491004 60078
rect 526404 60076 527004 60078
rect 562404 60076 563004 60078
rect 588140 60076 588740 60078
rect -4816 60054 588740 60076
rect -4816 59818 -4634 60054
rect -4398 59818 22586 60054
rect 22822 59818 58586 60054
rect 58822 59818 94586 60054
rect 94822 59818 130586 60054
rect 130822 59818 166586 60054
rect 166822 59818 202586 60054
rect 202822 59818 238586 60054
rect 238822 59818 274586 60054
rect 274822 59818 310586 60054
rect 310822 59818 346586 60054
rect 346822 59818 382586 60054
rect 382822 59818 418586 60054
rect 418822 59818 454586 60054
rect 454822 59818 490586 60054
rect 490822 59818 526586 60054
rect 526822 59818 562586 60054
rect 562822 59818 588322 60054
rect 588558 59818 588740 60054
rect -4816 59734 588740 59818
rect -4816 59498 -4634 59734
rect -4398 59498 22586 59734
rect 22822 59498 58586 59734
rect 58822 59498 94586 59734
rect 94822 59498 130586 59734
rect 130822 59498 166586 59734
rect 166822 59498 202586 59734
rect 202822 59498 238586 59734
rect 238822 59498 274586 59734
rect 274822 59498 310586 59734
rect 310822 59498 346586 59734
rect 346822 59498 382586 59734
rect 382822 59498 418586 59734
rect 418822 59498 454586 59734
rect 454822 59498 490586 59734
rect 490822 59498 526586 59734
rect 526822 59498 562586 59734
rect 562822 59498 588322 59734
rect 588558 59498 588740 59734
rect -4816 59476 588740 59498
rect -4816 59474 -4216 59476
rect 22404 59474 23004 59476
rect 58404 59474 59004 59476
rect 94404 59474 95004 59476
rect 130404 59474 131004 59476
rect 166404 59474 167004 59476
rect 202404 59474 203004 59476
rect 238404 59474 239004 59476
rect 274404 59474 275004 59476
rect 310404 59474 311004 59476
rect 346404 59474 347004 59476
rect 382404 59474 383004 59476
rect 418404 59474 419004 59476
rect 454404 59474 455004 59476
rect 490404 59474 491004 59476
rect 526404 59474 527004 59476
rect 562404 59474 563004 59476
rect 588140 59474 588740 59476
rect -2936 56476 -2336 56478
rect 18804 56476 19404 56478
rect 54804 56476 55404 56478
rect 90804 56476 91404 56478
rect 126804 56476 127404 56478
rect 162804 56476 163404 56478
rect 198804 56476 199404 56478
rect 234804 56476 235404 56478
rect 270804 56476 271404 56478
rect 306804 56476 307404 56478
rect 342804 56476 343404 56478
rect 378804 56476 379404 56478
rect 414804 56476 415404 56478
rect 450804 56476 451404 56478
rect 486804 56476 487404 56478
rect 522804 56476 523404 56478
rect 558804 56476 559404 56478
rect 586260 56476 586860 56478
rect -2936 56454 586860 56476
rect -2936 56218 -2754 56454
rect -2518 56218 18986 56454
rect 19222 56218 54986 56454
rect 55222 56218 90986 56454
rect 91222 56218 126986 56454
rect 127222 56218 162986 56454
rect 163222 56218 198986 56454
rect 199222 56218 234986 56454
rect 235222 56218 270986 56454
rect 271222 56218 306986 56454
rect 307222 56218 342986 56454
rect 343222 56218 378986 56454
rect 379222 56218 414986 56454
rect 415222 56218 450986 56454
rect 451222 56218 486986 56454
rect 487222 56218 522986 56454
rect 523222 56218 558986 56454
rect 559222 56218 586442 56454
rect 586678 56218 586860 56454
rect -2936 56134 586860 56218
rect -2936 55898 -2754 56134
rect -2518 55898 18986 56134
rect 19222 55898 54986 56134
rect 55222 55898 90986 56134
rect 91222 55898 126986 56134
rect 127222 55898 162986 56134
rect 163222 55898 198986 56134
rect 199222 55898 234986 56134
rect 235222 55898 270986 56134
rect 271222 55898 306986 56134
rect 307222 55898 342986 56134
rect 343222 55898 378986 56134
rect 379222 55898 414986 56134
rect 415222 55898 450986 56134
rect 451222 55898 486986 56134
rect 487222 55898 522986 56134
rect 523222 55898 558986 56134
rect 559222 55898 586442 56134
rect 586678 55898 586860 56134
rect -2936 55876 586860 55898
rect -2936 55874 -2336 55876
rect 18804 55874 19404 55876
rect 54804 55874 55404 55876
rect 90804 55874 91404 55876
rect 126804 55874 127404 55876
rect 162804 55874 163404 55876
rect 198804 55874 199404 55876
rect 234804 55874 235404 55876
rect 270804 55874 271404 55876
rect 306804 55874 307404 55876
rect 342804 55874 343404 55876
rect 378804 55874 379404 55876
rect 414804 55874 415404 55876
rect 450804 55874 451404 55876
rect 486804 55874 487404 55876
rect 522804 55874 523404 55876
rect 558804 55874 559404 55876
rect 586260 55874 586860 55876
rect -7636 49276 -7036 49278
rect 11604 49276 12204 49278
rect 47604 49276 48204 49278
rect 83604 49276 84204 49278
rect 119604 49276 120204 49278
rect 155604 49276 156204 49278
rect 191604 49276 192204 49278
rect 227604 49276 228204 49278
rect 263604 49276 264204 49278
rect 299604 49276 300204 49278
rect 335604 49276 336204 49278
rect 371604 49276 372204 49278
rect 407604 49276 408204 49278
rect 443604 49276 444204 49278
rect 479604 49276 480204 49278
rect 515604 49276 516204 49278
rect 551604 49276 552204 49278
rect 590960 49276 591560 49278
rect -8576 49254 592500 49276
rect -8576 49018 -7454 49254
rect -7218 49018 11786 49254
rect 12022 49018 47786 49254
rect 48022 49018 83786 49254
rect 84022 49018 119786 49254
rect 120022 49018 155786 49254
rect 156022 49018 191786 49254
rect 192022 49018 227786 49254
rect 228022 49018 263786 49254
rect 264022 49018 299786 49254
rect 300022 49018 335786 49254
rect 336022 49018 371786 49254
rect 372022 49018 407786 49254
rect 408022 49018 443786 49254
rect 444022 49018 479786 49254
rect 480022 49018 515786 49254
rect 516022 49018 551786 49254
rect 552022 49018 591142 49254
rect 591378 49018 592500 49254
rect -8576 48934 592500 49018
rect -8576 48698 -7454 48934
rect -7218 48698 11786 48934
rect 12022 48698 47786 48934
rect 48022 48698 83786 48934
rect 84022 48698 119786 48934
rect 120022 48698 155786 48934
rect 156022 48698 191786 48934
rect 192022 48698 227786 48934
rect 228022 48698 263786 48934
rect 264022 48698 299786 48934
rect 300022 48698 335786 48934
rect 336022 48698 371786 48934
rect 372022 48698 407786 48934
rect 408022 48698 443786 48934
rect 444022 48698 479786 48934
rect 480022 48698 515786 48934
rect 516022 48698 551786 48934
rect 552022 48698 591142 48934
rect 591378 48698 592500 48934
rect -8576 48676 592500 48698
rect -7636 48674 -7036 48676
rect 11604 48674 12204 48676
rect 47604 48674 48204 48676
rect 83604 48674 84204 48676
rect 119604 48674 120204 48676
rect 155604 48674 156204 48676
rect 191604 48674 192204 48676
rect 227604 48674 228204 48676
rect 263604 48674 264204 48676
rect 299604 48674 300204 48676
rect 335604 48674 336204 48676
rect 371604 48674 372204 48676
rect 407604 48674 408204 48676
rect 443604 48674 444204 48676
rect 479604 48674 480204 48676
rect 515604 48674 516204 48676
rect 551604 48674 552204 48676
rect 590960 48674 591560 48676
rect -5756 45676 -5156 45678
rect 8004 45676 8604 45678
rect 44004 45676 44604 45678
rect 80004 45676 80604 45678
rect 116004 45676 116604 45678
rect 152004 45676 152604 45678
rect 188004 45676 188604 45678
rect 224004 45676 224604 45678
rect 260004 45676 260604 45678
rect 296004 45676 296604 45678
rect 332004 45676 332604 45678
rect 368004 45676 368604 45678
rect 404004 45676 404604 45678
rect 440004 45676 440604 45678
rect 476004 45676 476604 45678
rect 512004 45676 512604 45678
rect 548004 45676 548604 45678
rect 589080 45676 589680 45678
rect -6696 45654 590620 45676
rect -6696 45418 -5574 45654
rect -5338 45418 8186 45654
rect 8422 45418 44186 45654
rect 44422 45418 80186 45654
rect 80422 45418 116186 45654
rect 116422 45418 152186 45654
rect 152422 45418 188186 45654
rect 188422 45418 224186 45654
rect 224422 45418 260186 45654
rect 260422 45418 296186 45654
rect 296422 45418 332186 45654
rect 332422 45418 368186 45654
rect 368422 45418 404186 45654
rect 404422 45418 440186 45654
rect 440422 45418 476186 45654
rect 476422 45418 512186 45654
rect 512422 45418 548186 45654
rect 548422 45418 589262 45654
rect 589498 45418 590620 45654
rect -6696 45334 590620 45418
rect -6696 45098 -5574 45334
rect -5338 45098 8186 45334
rect 8422 45098 44186 45334
rect 44422 45098 80186 45334
rect 80422 45098 116186 45334
rect 116422 45098 152186 45334
rect 152422 45098 188186 45334
rect 188422 45098 224186 45334
rect 224422 45098 260186 45334
rect 260422 45098 296186 45334
rect 296422 45098 332186 45334
rect 332422 45098 368186 45334
rect 368422 45098 404186 45334
rect 404422 45098 440186 45334
rect 440422 45098 476186 45334
rect 476422 45098 512186 45334
rect 512422 45098 548186 45334
rect 548422 45098 589262 45334
rect 589498 45098 590620 45334
rect -6696 45076 590620 45098
rect -5756 45074 -5156 45076
rect 8004 45074 8604 45076
rect 44004 45074 44604 45076
rect 80004 45074 80604 45076
rect 116004 45074 116604 45076
rect 152004 45074 152604 45076
rect 188004 45074 188604 45076
rect 224004 45074 224604 45076
rect 260004 45074 260604 45076
rect 296004 45074 296604 45076
rect 332004 45074 332604 45076
rect 368004 45074 368604 45076
rect 404004 45074 404604 45076
rect 440004 45074 440604 45076
rect 476004 45074 476604 45076
rect 512004 45074 512604 45076
rect 548004 45074 548604 45076
rect 589080 45074 589680 45076
rect -3876 42076 -3276 42078
rect 4404 42076 5004 42078
rect 40404 42076 41004 42078
rect 76404 42076 77004 42078
rect 112404 42076 113004 42078
rect 148404 42076 149004 42078
rect 184404 42076 185004 42078
rect 220404 42076 221004 42078
rect 256404 42076 257004 42078
rect 292404 42076 293004 42078
rect 328404 42076 329004 42078
rect 364404 42076 365004 42078
rect 400404 42076 401004 42078
rect 436404 42076 437004 42078
rect 472404 42076 473004 42078
rect 508404 42076 509004 42078
rect 544404 42076 545004 42078
rect 580404 42076 581004 42078
rect 587200 42076 587800 42078
rect -4816 42054 588740 42076
rect -4816 41818 -3694 42054
rect -3458 41818 4586 42054
rect 4822 41818 40586 42054
rect 40822 41818 76586 42054
rect 76822 41818 112586 42054
rect 112822 41818 148586 42054
rect 148822 41818 184586 42054
rect 184822 41818 220586 42054
rect 220822 41818 256586 42054
rect 256822 41818 292586 42054
rect 292822 41818 328586 42054
rect 328822 41818 364586 42054
rect 364822 41818 400586 42054
rect 400822 41818 436586 42054
rect 436822 41818 472586 42054
rect 472822 41818 508586 42054
rect 508822 41818 544586 42054
rect 544822 41818 580586 42054
rect 580822 41818 587382 42054
rect 587618 41818 588740 42054
rect -4816 41734 588740 41818
rect -4816 41498 -3694 41734
rect -3458 41498 4586 41734
rect 4822 41498 40586 41734
rect 40822 41498 76586 41734
rect 76822 41498 112586 41734
rect 112822 41498 148586 41734
rect 148822 41498 184586 41734
rect 184822 41498 220586 41734
rect 220822 41498 256586 41734
rect 256822 41498 292586 41734
rect 292822 41498 328586 41734
rect 328822 41498 364586 41734
rect 364822 41498 400586 41734
rect 400822 41498 436586 41734
rect 436822 41498 472586 41734
rect 472822 41498 508586 41734
rect 508822 41498 544586 41734
rect 544822 41498 580586 41734
rect 580822 41498 587382 41734
rect 587618 41498 588740 41734
rect -4816 41476 588740 41498
rect -3876 41474 -3276 41476
rect 4404 41474 5004 41476
rect 40404 41474 41004 41476
rect 76404 41474 77004 41476
rect 112404 41474 113004 41476
rect 148404 41474 149004 41476
rect 184404 41474 185004 41476
rect 220404 41474 221004 41476
rect 256404 41474 257004 41476
rect 292404 41474 293004 41476
rect 328404 41474 329004 41476
rect 364404 41474 365004 41476
rect 400404 41474 401004 41476
rect 436404 41474 437004 41476
rect 472404 41474 473004 41476
rect 508404 41474 509004 41476
rect 544404 41474 545004 41476
rect 580404 41474 581004 41476
rect 587200 41474 587800 41476
rect -1996 38476 -1396 38478
rect 804 38476 1404 38478
rect 36804 38476 37404 38478
rect 72804 38476 73404 38478
rect 108804 38476 109404 38478
rect 144804 38476 145404 38478
rect 180804 38476 181404 38478
rect 216804 38476 217404 38478
rect 252804 38476 253404 38478
rect 288804 38476 289404 38478
rect 324804 38476 325404 38478
rect 360804 38476 361404 38478
rect 396804 38476 397404 38478
rect 432804 38476 433404 38478
rect 468804 38476 469404 38478
rect 504804 38476 505404 38478
rect 540804 38476 541404 38478
rect 576804 38476 577404 38478
rect 585320 38476 585920 38478
rect -2936 38454 586860 38476
rect -2936 38218 -1814 38454
rect -1578 38218 986 38454
rect 1222 38218 36986 38454
rect 37222 38218 72986 38454
rect 73222 38218 108986 38454
rect 109222 38218 144986 38454
rect 145222 38218 180986 38454
rect 181222 38218 216986 38454
rect 217222 38218 252986 38454
rect 253222 38218 288986 38454
rect 289222 38218 324986 38454
rect 325222 38218 360986 38454
rect 361222 38218 396986 38454
rect 397222 38218 432986 38454
rect 433222 38218 468986 38454
rect 469222 38218 504986 38454
rect 505222 38218 540986 38454
rect 541222 38218 576986 38454
rect 577222 38218 585502 38454
rect 585738 38218 586860 38454
rect -2936 38134 586860 38218
rect -2936 37898 -1814 38134
rect -1578 37898 986 38134
rect 1222 37898 36986 38134
rect 37222 37898 72986 38134
rect 73222 37898 108986 38134
rect 109222 37898 144986 38134
rect 145222 37898 180986 38134
rect 181222 37898 216986 38134
rect 217222 37898 252986 38134
rect 253222 37898 288986 38134
rect 289222 37898 324986 38134
rect 325222 37898 360986 38134
rect 361222 37898 396986 38134
rect 397222 37898 432986 38134
rect 433222 37898 468986 38134
rect 469222 37898 504986 38134
rect 505222 37898 540986 38134
rect 541222 37898 576986 38134
rect 577222 37898 585502 38134
rect 585738 37898 586860 38134
rect -2936 37876 586860 37898
rect -1996 37874 -1396 37876
rect 804 37874 1404 37876
rect 36804 37874 37404 37876
rect 72804 37874 73404 37876
rect 108804 37874 109404 37876
rect 144804 37874 145404 37876
rect 180804 37874 181404 37876
rect 216804 37874 217404 37876
rect 252804 37874 253404 37876
rect 288804 37874 289404 37876
rect 324804 37874 325404 37876
rect 360804 37874 361404 37876
rect 396804 37874 397404 37876
rect 432804 37874 433404 37876
rect 468804 37874 469404 37876
rect 504804 37874 505404 37876
rect 540804 37874 541404 37876
rect 576804 37874 577404 37876
rect 585320 37874 585920 37876
rect -8576 31276 -7976 31278
rect 29604 31276 30204 31278
rect 65604 31276 66204 31278
rect 101604 31276 102204 31278
rect 137604 31276 138204 31278
rect 173604 31276 174204 31278
rect 209604 31276 210204 31278
rect 245604 31276 246204 31278
rect 281604 31276 282204 31278
rect 317604 31276 318204 31278
rect 353604 31276 354204 31278
rect 389604 31276 390204 31278
rect 425604 31276 426204 31278
rect 461604 31276 462204 31278
rect 497604 31276 498204 31278
rect 533604 31276 534204 31278
rect 569604 31276 570204 31278
rect 591900 31276 592500 31278
rect -8576 31254 592500 31276
rect -8576 31018 -8394 31254
rect -8158 31018 29786 31254
rect 30022 31018 65786 31254
rect 66022 31018 101786 31254
rect 102022 31018 137786 31254
rect 138022 31018 173786 31254
rect 174022 31018 209786 31254
rect 210022 31018 245786 31254
rect 246022 31018 281786 31254
rect 282022 31018 317786 31254
rect 318022 31018 353786 31254
rect 354022 31018 389786 31254
rect 390022 31018 425786 31254
rect 426022 31018 461786 31254
rect 462022 31018 497786 31254
rect 498022 31018 533786 31254
rect 534022 31018 569786 31254
rect 570022 31018 592082 31254
rect 592318 31018 592500 31254
rect -8576 30934 592500 31018
rect -8576 30698 -8394 30934
rect -8158 30698 29786 30934
rect 30022 30698 65786 30934
rect 66022 30698 101786 30934
rect 102022 30698 137786 30934
rect 138022 30698 173786 30934
rect 174022 30698 209786 30934
rect 210022 30698 245786 30934
rect 246022 30698 281786 30934
rect 282022 30698 317786 30934
rect 318022 30698 353786 30934
rect 354022 30698 389786 30934
rect 390022 30698 425786 30934
rect 426022 30698 461786 30934
rect 462022 30698 497786 30934
rect 498022 30698 533786 30934
rect 534022 30698 569786 30934
rect 570022 30698 592082 30934
rect 592318 30698 592500 30934
rect -8576 30676 592500 30698
rect -8576 30674 -7976 30676
rect 29604 30674 30204 30676
rect 65604 30674 66204 30676
rect 101604 30674 102204 30676
rect 137604 30674 138204 30676
rect 173604 30674 174204 30676
rect 209604 30674 210204 30676
rect 245604 30674 246204 30676
rect 281604 30674 282204 30676
rect 317604 30674 318204 30676
rect 353604 30674 354204 30676
rect 389604 30674 390204 30676
rect 425604 30674 426204 30676
rect 461604 30674 462204 30676
rect 497604 30674 498204 30676
rect 533604 30674 534204 30676
rect 569604 30674 570204 30676
rect 591900 30674 592500 30676
rect -6696 27676 -6096 27678
rect 26004 27676 26604 27678
rect 62004 27676 62604 27678
rect 98004 27676 98604 27678
rect 134004 27676 134604 27678
rect 170004 27676 170604 27678
rect 206004 27676 206604 27678
rect 242004 27676 242604 27678
rect 278004 27676 278604 27678
rect 314004 27676 314604 27678
rect 350004 27676 350604 27678
rect 386004 27676 386604 27678
rect 422004 27676 422604 27678
rect 458004 27676 458604 27678
rect 494004 27676 494604 27678
rect 530004 27676 530604 27678
rect 566004 27676 566604 27678
rect 590020 27676 590620 27678
rect -6696 27654 590620 27676
rect -6696 27418 -6514 27654
rect -6278 27418 26186 27654
rect 26422 27418 62186 27654
rect 62422 27418 98186 27654
rect 98422 27418 134186 27654
rect 134422 27418 170186 27654
rect 170422 27418 206186 27654
rect 206422 27418 242186 27654
rect 242422 27418 278186 27654
rect 278422 27418 314186 27654
rect 314422 27418 350186 27654
rect 350422 27418 386186 27654
rect 386422 27418 422186 27654
rect 422422 27418 458186 27654
rect 458422 27418 494186 27654
rect 494422 27418 530186 27654
rect 530422 27418 566186 27654
rect 566422 27418 590202 27654
rect 590438 27418 590620 27654
rect -6696 27334 590620 27418
rect -6696 27098 -6514 27334
rect -6278 27098 26186 27334
rect 26422 27098 62186 27334
rect 62422 27098 98186 27334
rect 98422 27098 134186 27334
rect 134422 27098 170186 27334
rect 170422 27098 206186 27334
rect 206422 27098 242186 27334
rect 242422 27098 278186 27334
rect 278422 27098 314186 27334
rect 314422 27098 350186 27334
rect 350422 27098 386186 27334
rect 386422 27098 422186 27334
rect 422422 27098 458186 27334
rect 458422 27098 494186 27334
rect 494422 27098 530186 27334
rect 530422 27098 566186 27334
rect 566422 27098 590202 27334
rect 590438 27098 590620 27334
rect -6696 27076 590620 27098
rect -6696 27074 -6096 27076
rect 26004 27074 26604 27076
rect 62004 27074 62604 27076
rect 98004 27074 98604 27076
rect 134004 27074 134604 27076
rect 170004 27074 170604 27076
rect 206004 27074 206604 27076
rect 242004 27074 242604 27076
rect 278004 27074 278604 27076
rect 314004 27074 314604 27076
rect 350004 27074 350604 27076
rect 386004 27074 386604 27076
rect 422004 27074 422604 27076
rect 458004 27074 458604 27076
rect 494004 27074 494604 27076
rect 530004 27074 530604 27076
rect 566004 27074 566604 27076
rect 590020 27074 590620 27076
rect -4816 24076 -4216 24078
rect 22404 24076 23004 24078
rect 58404 24076 59004 24078
rect 94404 24076 95004 24078
rect 130404 24076 131004 24078
rect 166404 24076 167004 24078
rect 202404 24076 203004 24078
rect 238404 24076 239004 24078
rect 274404 24076 275004 24078
rect 310404 24076 311004 24078
rect 346404 24076 347004 24078
rect 382404 24076 383004 24078
rect 418404 24076 419004 24078
rect 454404 24076 455004 24078
rect 490404 24076 491004 24078
rect 526404 24076 527004 24078
rect 562404 24076 563004 24078
rect 588140 24076 588740 24078
rect -4816 24054 588740 24076
rect -4816 23818 -4634 24054
rect -4398 23818 22586 24054
rect 22822 23818 58586 24054
rect 58822 23818 94586 24054
rect 94822 23818 130586 24054
rect 130822 23818 166586 24054
rect 166822 23818 202586 24054
rect 202822 23818 238586 24054
rect 238822 23818 274586 24054
rect 274822 23818 310586 24054
rect 310822 23818 346586 24054
rect 346822 23818 382586 24054
rect 382822 23818 418586 24054
rect 418822 23818 454586 24054
rect 454822 23818 490586 24054
rect 490822 23818 526586 24054
rect 526822 23818 562586 24054
rect 562822 23818 588322 24054
rect 588558 23818 588740 24054
rect -4816 23734 588740 23818
rect -4816 23498 -4634 23734
rect -4398 23498 22586 23734
rect 22822 23498 58586 23734
rect 58822 23498 94586 23734
rect 94822 23498 130586 23734
rect 130822 23498 166586 23734
rect 166822 23498 202586 23734
rect 202822 23498 238586 23734
rect 238822 23498 274586 23734
rect 274822 23498 310586 23734
rect 310822 23498 346586 23734
rect 346822 23498 382586 23734
rect 382822 23498 418586 23734
rect 418822 23498 454586 23734
rect 454822 23498 490586 23734
rect 490822 23498 526586 23734
rect 526822 23498 562586 23734
rect 562822 23498 588322 23734
rect 588558 23498 588740 23734
rect -4816 23476 588740 23498
rect -4816 23474 -4216 23476
rect 22404 23474 23004 23476
rect 58404 23474 59004 23476
rect 94404 23474 95004 23476
rect 130404 23474 131004 23476
rect 166404 23474 167004 23476
rect 202404 23474 203004 23476
rect 238404 23474 239004 23476
rect 274404 23474 275004 23476
rect 310404 23474 311004 23476
rect 346404 23474 347004 23476
rect 382404 23474 383004 23476
rect 418404 23474 419004 23476
rect 454404 23474 455004 23476
rect 490404 23474 491004 23476
rect 526404 23474 527004 23476
rect 562404 23474 563004 23476
rect 588140 23474 588740 23476
rect -2936 20476 -2336 20478
rect 18804 20476 19404 20478
rect 54804 20476 55404 20478
rect 90804 20476 91404 20478
rect 126804 20476 127404 20478
rect 162804 20476 163404 20478
rect 198804 20476 199404 20478
rect 234804 20476 235404 20478
rect 270804 20476 271404 20478
rect 306804 20476 307404 20478
rect 342804 20476 343404 20478
rect 378804 20476 379404 20478
rect 414804 20476 415404 20478
rect 450804 20476 451404 20478
rect 486804 20476 487404 20478
rect 522804 20476 523404 20478
rect 558804 20476 559404 20478
rect 586260 20476 586860 20478
rect -2936 20454 586860 20476
rect -2936 20218 -2754 20454
rect -2518 20218 18986 20454
rect 19222 20218 54986 20454
rect 55222 20218 90986 20454
rect 91222 20218 126986 20454
rect 127222 20218 162986 20454
rect 163222 20218 198986 20454
rect 199222 20218 234986 20454
rect 235222 20218 270986 20454
rect 271222 20218 306986 20454
rect 307222 20218 342986 20454
rect 343222 20218 378986 20454
rect 379222 20218 414986 20454
rect 415222 20218 450986 20454
rect 451222 20218 486986 20454
rect 487222 20218 522986 20454
rect 523222 20218 558986 20454
rect 559222 20218 586442 20454
rect 586678 20218 586860 20454
rect -2936 20134 586860 20218
rect -2936 19898 -2754 20134
rect -2518 19898 18986 20134
rect 19222 19898 54986 20134
rect 55222 19898 90986 20134
rect 91222 19898 126986 20134
rect 127222 19898 162986 20134
rect 163222 19898 198986 20134
rect 199222 19898 234986 20134
rect 235222 19898 270986 20134
rect 271222 19898 306986 20134
rect 307222 19898 342986 20134
rect 343222 19898 378986 20134
rect 379222 19898 414986 20134
rect 415222 19898 450986 20134
rect 451222 19898 486986 20134
rect 487222 19898 522986 20134
rect 523222 19898 558986 20134
rect 559222 19898 586442 20134
rect 586678 19898 586860 20134
rect -2936 19876 586860 19898
rect -2936 19874 -2336 19876
rect 18804 19874 19404 19876
rect 54804 19874 55404 19876
rect 90804 19874 91404 19876
rect 126804 19874 127404 19876
rect 162804 19874 163404 19876
rect 198804 19874 199404 19876
rect 234804 19874 235404 19876
rect 270804 19874 271404 19876
rect 306804 19874 307404 19876
rect 342804 19874 343404 19876
rect 378804 19874 379404 19876
rect 414804 19874 415404 19876
rect 450804 19874 451404 19876
rect 486804 19874 487404 19876
rect 522804 19874 523404 19876
rect 558804 19874 559404 19876
rect 586260 19874 586860 19876
rect -7636 13276 -7036 13278
rect 11604 13276 12204 13278
rect 47604 13276 48204 13278
rect 83604 13276 84204 13278
rect 119604 13276 120204 13278
rect 155604 13276 156204 13278
rect 191604 13276 192204 13278
rect 227604 13276 228204 13278
rect 263604 13276 264204 13278
rect 299604 13276 300204 13278
rect 335604 13276 336204 13278
rect 371604 13276 372204 13278
rect 407604 13276 408204 13278
rect 443604 13276 444204 13278
rect 479604 13276 480204 13278
rect 515604 13276 516204 13278
rect 551604 13276 552204 13278
rect 590960 13276 591560 13278
rect -8576 13254 592500 13276
rect -8576 13018 -7454 13254
rect -7218 13018 11786 13254
rect 12022 13018 47786 13254
rect 48022 13018 83786 13254
rect 84022 13018 119786 13254
rect 120022 13018 155786 13254
rect 156022 13018 191786 13254
rect 192022 13018 227786 13254
rect 228022 13018 263786 13254
rect 264022 13018 299786 13254
rect 300022 13018 335786 13254
rect 336022 13018 371786 13254
rect 372022 13018 407786 13254
rect 408022 13018 443786 13254
rect 444022 13018 479786 13254
rect 480022 13018 515786 13254
rect 516022 13018 551786 13254
rect 552022 13018 591142 13254
rect 591378 13018 592500 13254
rect -8576 12934 592500 13018
rect -8576 12698 -7454 12934
rect -7218 12698 11786 12934
rect 12022 12698 47786 12934
rect 48022 12698 83786 12934
rect 84022 12698 119786 12934
rect 120022 12698 155786 12934
rect 156022 12698 191786 12934
rect 192022 12698 227786 12934
rect 228022 12698 263786 12934
rect 264022 12698 299786 12934
rect 300022 12698 335786 12934
rect 336022 12698 371786 12934
rect 372022 12698 407786 12934
rect 408022 12698 443786 12934
rect 444022 12698 479786 12934
rect 480022 12698 515786 12934
rect 516022 12698 551786 12934
rect 552022 12698 591142 12934
rect 591378 12698 592500 12934
rect -8576 12676 592500 12698
rect -7636 12674 -7036 12676
rect 11604 12674 12204 12676
rect 47604 12674 48204 12676
rect 83604 12674 84204 12676
rect 119604 12674 120204 12676
rect 155604 12674 156204 12676
rect 191604 12674 192204 12676
rect 227604 12674 228204 12676
rect 263604 12674 264204 12676
rect 299604 12674 300204 12676
rect 335604 12674 336204 12676
rect 371604 12674 372204 12676
rect 407604 12674 408204 12676
rect 443604 12674 444204 12676
rect 479604 12674 480204 12676
rect 515604 12674 516204 12676
rect 551604 12674 552204 12676
rect 590960 12674 591560 12676
rect -5756 9676 -5156 9678
rect 8004 9676 8604 9678
rect 44004 9676 44604 9678
rect 80004 9676 80604 9678
rect 116004 9676 116604 9678
rect 152004 9676 152604 9678
rect 188004 9676 188604 9678
rect 224004 9676 224604 9678
rect 260004 9676 260604 9678
rect 296004 9676 296604 9678
rect 332004 9676 332604 9678
rect 368004 9676 368604 9678
rect 404004 9676 404604 9678
rect 440004 9676 440604 9678
rect 476004 9676 476604 9678
rect 512004 9676 512604 9678
rect 548004 9676 548604 9678
rect 589080 9676 589680 9678
rect -6696 9654 590620 9676
rect -6696 9418 -5574 9654
rect -5338 9418 8186 9654
rect 8422 9418 44186 9654
rect 44422 9418 80186 9654
rect 80422 9418 116186 9654
rect 116422 9418 152186 9654
rect 152422 9418 188186 9654
rect 188422 9418 224186 9654
rect 224422 9418 260186 9654
rect 260422 9418 296186 9654
rect 296422 9418 332186 9654
rect 332422 9418 368186 9654
rect 368422 9418 404186 9654
rect 404422 9418 440186 9654
rect 440422 9418 476186 9654
rect 476422 9418 512186 9654
rect 512422 9418 548186 9654
rect 548422 9418 589262 9654
rect 589498 9418 590620 9654
rect -6696 9334 590620 9418
rect -6696 9098 -5574 9334
rect -5338 9098 8186 9334
rect 8422 9098 44186 9334
rect 44422 9098 80186 9334
rect 80422 9098 116186 9334
rect 116422 9098 152186 9334
rect 152422 9098 188186 9334
rect 188422 9098 224186 9334
rect 224422 9098 260186 9334
rect 260422 9098 296186 9334
rect 296422 9098 332186 9334
rect 332422 9098 368186 9334
rect 368422 9098 404186 9334
rect 404422 9098 440186 9334
rect 440422 9098 476186 9334
rect 476422 9098 512186 9334
rect 512422 9098 548186 9334
rect 548422 9098 589262 9334
rect 589498 9098 590620 9334
rect -6696 9076 590620 9098
rect -5756 9074 -5156 9076
rect 8004 9074 8604 9076
rect 44004 9074 44604 9076
rect 80004 9074 80604 9076
rect 116004 9074 116604 9076
rect 152004 9074 152604 9076
rect 188004 9074 188604 9076
rect 224004 9074 224604 9076
rect 260004 9074 260604 9076
rect 296004 9074 296604 9076
rect 332004 9074 332604 9076
rect 368004 9074 368604 9076
rect 404004 9074 404604 9076
rect 440004 9074 440604 9076
rect 476004 9074 476604 9076
rect 512004 9074 512604 9076
rect 548004 9074 548604 9076
rect 589080 9074 589680 9076
rect -3876 6076 -3276 6078
rect 4404 6076 5004 6078
rect 40404 6076 41004 6078
rect 76404 6076 77004 6078
rect 112404 6076 113004 6078
rect 148404 6076 149004 6078
rect 184404 6076 185004 6078
rect 220404 6076 221004 6078
rect 256404 6076 257004 6078
rect 292404 6076 293004 6078
rect 328404 6076 329004 6078
rect 364404 6076 365004 6078
rect 400404 6076 401004 6078
rect 436404 6076 437004 6078
rect 472404 6076 473004 6078
rect 508404 6076 509004 6078
rect 544404 6076 545004 6078
rect 580404 6076 581004 6078
rect 587200 6076 587800 6078
rect -4816 6054 588740 6076
rect -4816 5818 -3694 6054
rect -3458 5818 4586 6054
rect 4822 5818 40586 6054
rect 40822 5818 76586 6054
rect 76822 5818 112586 6054
rect 112822 5818 148586 6054
rect 148822 5818 184586 6054
rect 184822 5818 220586 6054
rect 220822 5818 256586 6054
rect 256822 5818 292586 6054
rect 292822 5818 328586 6054
rect 328822 5818 364586 6054
rect 364822 5818 400586 6054
rect 400822 5818 436586 6054
rect 436822 5818 472586 6054
rect 472822 5818 508586 6054
rect 508822 5818 544586 6054
rect 544822 5818 580586 6054
rect 580822 5818 587382 6054
rect 587618 5818 588740 6054
rect -4816 5734 588740 5818
rect -4816 5498 -3694 5734
rect -3458 5498 4586 5734
rect 4822 5498 40586 5734
rect 40822 5498 76586 5734
rect 76822 5498 112586 5734
rect 112822 5498 148586 5734
rect 148822 5498 184586 5734
rect 184822 5498 220586 5734
rect 220822 5498 256586 5734
rect 256822 5498 292586 5734
rect 292822 5498 328586 5734
rect 328822 5498 364586 5734
rect 364822 5498 400586 5734
rect 400822 5498 436586 5734
rect 436822 5498 472586 5734
rect 472822 5498 508586 5734
rect 508822 5498 544586 5734
rect 544822 5498 580586 5734
rect 580822 5498 587382 5734
rect 587618 5498 588740 5734
rect -4816 5476 588740 5498
rect -3876 5474 -3276 5476
rect 4404 5474 5004 5476
rect 40404 5474 41004 5476
rect 76404 5474 77004 5476
rect 112404 5474 113004 5476
rect 148404 5474 149004 5476
rect 184404 5474 185004 5476
rect 220404 5474 221004 5476
rect 256404 5474 257004 5476
rect 292404 5474 293004 5476
rect 328404 5474 329004 5476
rect 364404 5474 365004 5476
rect 400404 5474 401004 5476
rect 436404 5474 437004 5476
rect 472404 5474 473004 5476
rect 508404 5474 509004 5476
rect 544404 5474 545004 5476
rect 580404 5474 581004 5476
rect 587200 5474 587800 5476
rect -1996 2476 -1396 2478
rect 804 2476 1404 2478
rect 36804 2476 37404 2478
rect 72804 2476 73404 2478
rect 108804 2476 109404 2478
rect 144804 2476 145404 2478
rect 180804 2476 181404 2478
rect 216804 2476 217404 2478
rect 252804 2476 253404 2478
rect 288804 2476 289404 2478
rect 324804 2476 325404 2478
rect 360804 2476 361404 2478
rect 396804 2476 397404 2478
rect 432804 2476 433404 2478
rect 468804 2476 469404 2478
rect 504804 2476 505404 2478
rect 540804 2476 541404 2478
rect 576804 2476 577404 2478
rect 585320 2476 585920 2478
rect -2936 2454 586860 2476
rect -2936 2218 -1814 2454
rect -1578 2218 986 2454
rect 1222 2218 36986 2454
rect 37222 2218 72986 2454
rect 73222 2218 108986 2454
rect 109222 2218 144986 2454
rect 145222 2218 180986 2454
rect 181222 2218 216986 2454
rect 217222 2218 252986 2454
rect 253222 2218 288986 2454
rect 289222 2218 324986 2454
rect 325222 2218 360986 2454
rect 361222 2218 396986 2454
rect 397222 2218 432986 2454
rect 433222 2218 468986 2454
rect 469222 2218 504986 2454
rect 505222 2218 540986 2454
rect 541222 2218 576986 2454
rect 577222 2218 585502 2454
rect 585738 2218 586860 2454
rect -2936 2134 586860 2218
rect -2936 1898 -1814 2134
rect -1578 1898 986 2134
rect 1222 1898 36986 2134
rect 37222 1898 72986 2134
rect 73222 1898 108986 2134
rect 109222 1898 144986 2134
rect 145222 1898 180986 2134
rect 181222 1898 216986 2134
rect 217222 1898 252986 2134
rect 253222 1898 288986 2134
rect 289222 1898 324986 2134
rect 325222 1898 360986 2134
rect 361222 1898 396986 2134
rect 397222 1898 432986 2134
rect 433222 1898 468986 2134
rect 469222 1898 504986 2134
rect 505222 1898 540986 2134
rect 541222 1898 576986 2134
rect 577222 1898 585502 2134
rect 585738 1898 586860 2134
rect -2936 1876 586860 1898
rect -1996 1874 -1396 1876
rect 804 1874 1404 1876
rect 36804 1874 37404 1876
rect 72804 1874 73404 1876
rect 108804 1874 109404 1876
rect 144804 1874 145404 1876
rect 180804 1874 181404 1876
rect 216804 1874 217404 1876
rect 252804 1874 253404 1876
rect 288804 1874 289404 1876
rect 324804 1874 325404 1876
rect 360804 1874 361404 1876
rect 396804 1874 397404 1876
rect 432804 1874 433404 1876
rect 468804 1874 469404 1876
rect 504804 1874 505404 1876
rect 540804 1874 541404 1876
rect 576804 1874 577404 1876
rect 585320 1874 585920 1876
rect -1996 -324 -1396 -322
rect 804 -324 1404 -322
rect 36804 -324 37404 -322
rect 72804 -324 73404 -322
rect 108804 -324 109404 -322
rect 144804 -324 145404 -322
rect 180804 -324 181404 -322
rect 216804 -324 217404 -322
rect 252804 -324 253404 -322
rect 288804 -324 289404 -322
rect 324804 -324 325404 -322
rect 360804 -324 361404 -322
rect 396804 -324 397404 -322
rect 432804 -324 433404 -322
rect 468804 -324 469404 -322
rect 504804 -324 505404 -322
rect 540804 -324 541404 -322
rect 576804 -324 577404 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 986 -346
rect 1222 -582 36986 -346
rect 37222 -582 72986 -346
rect 73222 -582 108986 -346
rect 109222 -582 144986 -346
rect 145222 -582 180986 -346
rect 181222 -582 216986 -346
rect 217222 -582 252986 -346
rect 253222 -582 288986 -346
rect 289222 -582 324986 -346
rect 325222 -582 360986 -346
rect 361222 -582 396986 -346
rect 397222 -582 432986 -346
rect 433222 -582 468986 -346
rect 469222 -582 504986 -346
rect 505222 -582 540986 -346
rect 541222 -582 576986 -346
rect 577222 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 986 -666
rect 1222 -902 36986 -666
rect 37222 -902 72986 -666
rect 73222 -902 108986 -666
rect 109222 -902 144986 -666
rect 145222 -902 180986 -666
rect 181222 -902 216986 -666
rect 217222 -902 252986 -666
rect 253222 -902 288986 -666
rect 289222 -902 324986 -666
rect 325222 -902 360986 -666
rect 361222 -902 396986 -666
rect 397222 -902 432986 -666
rect 433222 -902 468986 -666
rect 469222 -902 504986 -666
rect 505222 -902 540986 -666
rect 541222 -902 576986 -666
rect 577222 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 108804 -926 109404 -924
rect 144804 -926 145404 -924
rect 180804 -926 181404 -924
rect 216804 -926 217404 -924
rect 252804 -926 253404 -924
rect 288804 -926 289404 -924
rect 324804 -926 325404 -924
rect 360804 -926 361404 -924
rect 396804 -926 397404 -924
rect 432804 -926 433404 -924
rect 468804 -926 469404 -924
rect 504804 -926 505404 -924
rect 540804 -926 541404 -924
rect 576804 -926 577404 -924
rect 585320 -926 585920 -924
rect -2936 -1264 -2336 -1262
rect 18804 -1264 19404 -1262
rect 54804 -1264 55404 -1262
rect 90804 -1264 91404 -1262
rect 126804 -1264 127404 -1262
rect 162804 -1264 163404 -1262
rect 198804 -1264 199404 -1262
rect 234804 -1264 235404 -1262
rect 270804 -1264 271404 -1262
rect 306804 -1264 307404 -1262
rect 342804 -1264 343404 -1262
rect 378804 -1264 379404 -1262
rect 414804 -1264 415404 -1262
rect 450804 -1264 451404 -1262
rect 486804 -1264 487404 -1262
rect 522804 -1264 523404 -1262
rect 558804 -1264 559404 -1262
rect 586260 -1264 586860 -1262
rect -2936 -1286 586860 -1264
rect -2936 -1522 -2754 -1286
rect -2518 -1522 18986 -1286
rect 19222 -1522 54986 -1286
rect 55222 -1522 90986 -1286
rect 91222 -1522 126986 -1286
rect 127222 -1522 162986 -1286
rect 163222 -1522 198986 -1286
rect 199222 -1522 234986 -1286
rect 235222 -1522 270986 -1286
rect 271222 -1522 306986 -1286
rect 307222 -1522 342986 -1286
rect 343222 -1522 378986 -1286
rect 379222 -1522 414986 -1286
rect 415222 -1522 450986 -1286
rect 451222 -1522 486986 -1286
rect 487222 -1522 522986 -1286
rect 523222 -1522 558986 -1286
rect 559222 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect -2936 -1606 586860 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 18986 -1606
rect 19222 -1842 54986 -1606
rect 55222 -1842 90986 -1606
rect 91222 -1842 126986 -1606
rect 127222 -1842 162986 -1606
rect 163222 -1842 198986 -1606
rect 199222 -1842 234986 -1606
rect 235222 -1842 270986 -1606
rect 271222 -1842 306986 -1606
rect 307222 -1842 342986 -1606
rect 343222 -1842 378986 -1606
rect 379222 -1842 414986 -1606
rect 415222 -1842 450986 -1606
rect 451222 -1842 486986 -1606
rect 487222 -1842 522986 -1606
rect 523222 -1842 558986 -1606
rect 559222 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect -2936 -1864 586860 -1842
rect -2936 -1866 -2336 -1864
rect 18804 -1866 19404 -1864
rect 54804 -1866 55404 -1864
rect 90804 -1866 91404 -1864
rect 126804 -1866 127404 -1864
rect 162804 -1866 163404 -1864
rect 198804 -1866 199404 -1864
rect 234804 -1866 235404 -1864
rect 270804 -1866 271404 -1864
rect 306804 -1866 307404 -1864
rect 342804 -1866 343404 -1864
rect 378804 -1866 379404 -1864
rect 414804 -1866 415404 -1864
rect 450804 -1866 451404 -1864
rect 486804 -1866 487404 -1864
rect 522804 -1866 523404 -1864
rect 558804 -1866 559404 -1864
rect 586260 -1866 586860 -1864
rect -3876 -2204 -3276 -2202
rect 4404 -2204 5004 -2202
rect 40404 -2204 41004 -2202
rect 76404 -2204 77004 -2202
rect 112404 -2204 113004 -2202
rect 148404 -2204 149004 -2202
rect 184404 -2204 185004 -2202
rect 220404 -2204 221004 -2202
rect 256404 -2204 257004 -2202
rect 292404 -2204 293004 -2202
rect 328404 -2204 329004 -2202
rect 364404 -2204 365004 -2202
rect 400404 -2204 401004 -2202
rect 436404 -2204 437004 -2202
rect 472404 -2204 473004 -2202
rect 508404 -2204 509004 -2202
rect 544404 -2204 545004 -2202
rect 580404 -2204 581004 -2202
rect 587200 -2204 587800 -2202
rect -3876 -2226 587800 -2204
rect -3876 -2462 -3694 -2226
rect -3458 -2462 4586 -2226
rect 4822 -2462 40586 -2226
rect 40822 -2462 76586 -2226
rect 76822 -2462 112586 -2226
rect 112822 -2462 148586 -2226
rect 148822 -2462 184586 -2226
rect 184822 -2462 220586 -2226
rect 220822 -2462 256586 -2226
rect 256822 -2462 292586 -2226
rect 292822 -2462 328586 -2226
rect 328822 -2462 364586 -2226
rect 364822 -2462 400586 -2226
rect 400822 -2462 436586 -2226
rect 436822 -2462 472586 -2226
rect 472822 -2462 508586 -2226
rect 508822 -2462 544586 -2226
rect 544822 -2462 580586 -2226
rect 580822 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect -3876 -2546 587800 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 4586 -2546
rect 4822 -2782 40586 -2546
rect 40822 -2782 76586 -2546
rect 76822 -2782 112586 -2546
rect 112822 -2782 148586 -2546
rect 148822 -2782 184586 -2546
rect 184822 -2782 220586 -2546
rect 220822 -2782 256586 -2546
rect 256822 -2782 292586 -2546
rect 292822 -2782 328586 -2546
rect 328822 -2782 364586 -2546
rect 364822 -2782 400586 -2546
rect 400822 -2782 436586 -2546
rect 436822 -2782 472586 -2546
rect 472822 -2782 508586 -2546
rect 508822 -2782 544586 -2546
rect 544822 -2782 580586 -2546
rect 580822 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect -3876 -2804 587800 -2782
rect -3876 -2806 -3276 -2804
rect 4404 -2806 5004 -2804
rect 40404 -2806 41004 -2804
rect 76404 -2806 77004 -2804
rect 112404 -2806 113004 -2804
rect 148404 -2806 149004 -2804
rect 184404 -2806 185004 -2804
rect 220404 -2806 221004 -2804
rect 256404 -2806 257004 -2804
rect 292404 -2806 293004 -2804
rect 328404 -2806 329004 -2804
rect 364404 -2806 365004 -2804
rect 400404 -2806 401004 -2804
rect 436404 -2806 437004 -2804
rect 472404 -2806 473004 -2804
rect 508404 -2806 509004 -2804
rect 544404 -2806 545004 -2804
rect 580404 -2806 581004 -2804
rect 587200 -2806 587800 -2804
rect -4816 -3144 -4216 -3142
rect 22404 -3144 23004 -3142
rect 58404 -3144 59004 -3142
rect 94404 -3144 95004 -3142
rect 130404 -3144 131004 -3142
rect 166404 -3144 167004 -3142
rect 202404 -3144 203004 -3142
rect 238404 -3144 239004 -3142
rect 274404 -3144 275004 -3142
rect 310404 -3144 311004 -3142
rect 346404 -3144 347004 -3142
rect 382404 -3144 383004 -3142
rect 418404 -3144 419004 -3142
rect 454404 -3144 455004 -3142
rect 490404 -3144 491004 -3142
rect 526404 -3144 527004 -3142
rect 562404 -3144 563004 -3142
rect 588140 -3144 588740 -3142
rect -4816 -3166 588740 -3144
rect -4816 -3402 -4634 -3166
rect -4398 -3402 22586 -3166
rect 22822 -3402 58586 -3166
rect 58822 -3402 94586 -3166
rect 94822 -3402 130586 -3166
rect 130822 -3402 166586 -3166
rect 166822 -3402 202586 -3166
rect 202822 -3402 238586 -3166
rect 238822 -3402 274586 -3166
rect 274822 -3402 310586 -3166
rect 310822 -3402 346586 -3166
rect 346822 -3402 382586 -3166
rect 382822 -3402 418586 -3166
rect 418822 -3402 454586 -3166
rect 454822 -3402 490586 -3166
rect 490822 -3402 526586 -3166
rect 526822 -3402 562586 -3166
rect 562822 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect -4816 -3486 588740 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 22586 -3486
rect 22822 -3722 58586 -3486
rect 58822 -3722 94586 -3486
rect 94822 -3722 130586 -3486
rect 130822 -3722 166586 -3486
rect 166822 -3722 202586 -3486
rect 202822 -3722 238586 -3486
rect 238822 -3722 274586 -3486
rect 274822 -3722 310586 -3486
rect 310822 -3722 346586 -3486
rect 346822 -3722 382586 -3486
rect 382822 -3722 418586 -3486
rect 418822 -3722 454586 -3486
rect 454822 -3722 490586 -3486
rect 490822 -3722 526586 -3486
rect 526822 -3722 562586 -3486
rect 562822 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect -4816 -3744 588740 -3722
rect -4816 -3746 -4216 -3744
rect 22404 -3746 23004 -3744
rect 58404 -3746 59004 -3744
rect 94404 -3746 95004 -3744
rect 130404 -3746 131004 -3744
rect 166404 -3746 167004 -3744
rect 202404 -3746 203004 -3744
rect 238404 -3746 239004 -3744
rect 274404 -3746 275004 -3744
rect 310404 -3746 311004 -3744
rect 346404 -3746 347004 -3744
rect 382404 -3746 383004 -3744
rect 418404 -3746 419004 -3744
rect 454404 -3746 455004 -3744
rect 490404 -3746 491004 -3744
rect 526404 -3746 527004 -3744
rect 562404 -3746 563004 -3744
rect 588140 -3746 588740 -3744
rect -5756 -4084 -5156 -4082
rect 8004 -4084 8604 -4082
rect 44004 -4084 44604 -4082
rect 80004 -4084 80604 -4082
rect 116004 -4084 116604 -4082
rect 152004 -4084 152604 -4082
rect 188004 -4084 188604 -4082
rect 224004 -4084 224604 -4082
rect 260004 -4084 260604 -4082
rect 296004 -4084 296604 -4082
rect 332004 -4084 332604 -4082
rect 368004 -4084 368604 -4082
rect 404004 -4084 404604 -4082
rect 440004 -4084 440604 -4082
rect 476004 -4084 476604 -4082
rect 512004 -4084 512604 -4082
rect 548004 -4084 548604 -4082
rect 589080 -4084 589680 -4082
rect -5756 -4106 589680 -4084
rect -5756 -4342 -5574 -4106
rect -5338 -4342 8186 -4106
rect 8422 -4342 44186 -4106
rect 44422 -4342 80186 -4106
rect 80422 -4342 116186 -4106
rect 116422 -4342 152186 -4106
rect 152422 -4342 188186 -4106
rect 188422 -4342 224186 -4106
rect 224422 -4342 260186 -4106
rect 260422 -4342 296186 -4106
rect 296422 -4342 332186 -4106
rect 332422 -4342 368186 -4106
rect 368422 -4342 404186 -4106
rect 404422 -4342 440186 -4106
rect 440422 -4342 476186 -4106
rect 476422 -4342 512186 -4106
rect 512422 -4342 548186 -4106
rect 548422 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect -5756 -4426 589680 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 8186 -4426
rect 8422 -4662 44186 -4426
rect 44422 -4662 80186 -4426
rect 80422 -4662 116186 -4426
rect 116422 -4662 152186 -4426
rect 152422 -4662 188186 -4426
rect 188422 -4662 224186 -4426
rect 224422 -4662 260186 -4426
rect 260422 -4662 296186 -4426
rect 296422 -4662 332186 -4426
rect 332422 -4662 368186 -4426
rect 368422 -4662 404186 -4426
rect 404422 -4662 440186 -4426
rect 440422 -4662 476186 -4426
rect 476422 -4662 512186 -4426
rect 512422 -4662 548186 -4426
rect 548422 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect -5756 -4684 589680 -4662
rect -5756 -4686 -5156 -4684
rect 8004 -4686 8604 -4684
rect 44004 -4686 44604 -4684
rect 80004 -4686 80604 -4684
rect 116004 -4686 116604 -4684
rect 152004 -4686 152604 -4684
rect 188004 -4686 188604 -4684
rect 224004 -4686 224604 -4684
rect 260004 -4686 260604 -4684
rect 296004 -4686 296604 -4684
rect 332004 -4686 332604 -4684
rect 368004 -4686 368604 -4684
rect 404004 -4686 404604 -4684
rect 440004 -4686 440604 -4684
rect 476004 -4686 476604 -4684
rect 512004 -4686 512604 -4684
rect 548004 -4686 548604 -4684
rect 589080 -4686 589680 -4684
rect -6696 -5024 -6096 -5022
rect 26004 -5024 26604 -5022
rect 62004 -5024 62604 -5022
rect 98004 -5024 98604 -5022
rect 134004 -5024 134604 -5022
rect 170004 -5024 170604 -5022
rect 206004 -5024 206604 -5022
rect 242004 -5024 242604 -5022
rect 278004 -5024 278604 -5022
rect 314004 -5024 314604 -5022
rect 350004 -5024 350604 -5022
rect 386004 -5024 386604 -5022
rect 422004 -5024 422604 -5022
rect 458004 -5024 458604 -5022
rect 494004 -5024 494604 -5022
rect 530004 -5024 530604 -5022
rect 566004 -5024 566604 -5022
rect 590020 -5024 590620 -5022
rect -6696 -5046 590620 -5024
rect -6696 -5282 -6514 -5046
rect -6278 -5282 26186 -5046
rect 26422 -5282 62186 -5046
rect 62422 -5282 98186 -5046
rect 98422 -5282 134186 -5046
rect 134422 -5282 170186 -5046
rect 170422 -5282 206186 -5046
rect 206422 -5282 242186 -5046
rect 242422 -5282 278186 -5046
rect 278422 -5282 314186 -5046
rect 314422 -5282 350186 -5046
rect 350422 -5282 386186 -5046
rect 386422 -5282 422186 -5046
rect 422422 -5282 458186 -5046
rect 458422 -5282 494186 -5046
rect 494422 -5282 530186 -5046
rect 530422 -5282 566186 -5046
rect 566422 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect -6696 -5366 590620 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 26186 -5366
rect 26422 -5602 62186 -5366
rect 62422 -5602 98186 -5366
rect 98422 -5602 134186 -5366
rect 134422 -5602 170186 -5366
rect 170422 -5602 206186 -5366
rect 206422 -5602 242186 -5366
rect 242422 -5602 278186 -5366
rect 278422 -5602 314186 -5366
rect 314422 -5602 350186 -5366
rect 350422 -5602 386186 -5366
rect 386422 -5602 422186 -5366
rect 422422 -5602 458186 -5366
rect 458422 -5602 494186 -5366
rect 494422 -5602 530186 -5366
rect 530422 -5602 566186 -5366
rect 566422 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect -6696 -5624 590620 -5602
rect -6696 -5626 -6096 -5624
rect 26004 -5626 26604 -5624
rect 62004 -5626 62604 -5624
rect 98004 -5626 98604 -5624
rect 134004 -5626 134604 -5624
rect 170004 -5626 170604 -5624
rect 206004 -5626 206604 -5624
rect 242004 -5626 242604 -5624
rect 278004 -5626 278604 -5624
rect 314004 -5626 314604 -5624
rect 350004 -5626 350604 -5624
rect 386004 -5626 386604 -5624
rect 422004 -5626 422604 -5624
rect 458004 -5626 458604 -5624
rect 494004 -5626 494604 -5624
rect 530004 -5626 530604 -5624
rect 566004 -5626 566604 -5624
rect 590020 -5626 590620 -5624
rect -7636 -5964 -7036 -5962
rect 11604 -5964 12204 -5962
rect 47604 -5964 48204 -5962
rect 83604 -5964 84204 -5962
rect 119604 -5964 120204 -5962
rect 155604 -5964 156204 -5962
rect 191604 -5964 192204 -5962
rect 227604 -5964 228204 -5962
rect 263604 -5964 264204 -5962
rect 299604 -5964 300204 -5962
rect 335604 -5964 336204 -5962
rect 371604 -5964 372204 -5962
rect 407604 -5964 408204 -5962
rect 443604 -5964 444204 -5962
rect 479604 -5964 480204 -5962
rect 515604 -5964 516204 -5962
rect 551604 -5964 552204 -5962
rect 590960 -5964 591560 -5962
rect -7636 -5986 591560 -5964
rect -7636 -6222 -7454 -5986
rect -7218 -6222 11786 -5986
rect 12022 -6222 47786 -5986
rect 48022 -6222 83786 -5986
rect 84022 -6222 119786 -5986
rect 120022 -6222 155786 -5986
rect 156022 -6222 191786 -5986
rect 192022 -6222 227786 -5986
rect 228022 -6222 263786 -5986
rect 264022 -6222 299786 -5986
rect 300022 -6222 335786 -5986
rect 336022 -6222 371786 -5986
rect 372022 -6222 407786 -5986
rect 408022 -6222 443786 -5986
rect 444022 -6222 479786 -5986
rect 480022 -6222 515786 -5986
rect 516022 -6222 551786 -5986
rect 552022 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect -7636 -6306 591560 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 11786 -6306
rect 12022 -6542 47786 -6306
rect 48022 -6542 83786 -6306
rect 84022 -6542 119786 -6306
rect 120022 -6542 155786 -6306
rect 156022 -6542 191786 -6306
rect 192022 -6542 227786 -6306
rect 228022 -6542 263786 -6306
rect 264022 -6542 299786 -6306
rect 300022 -6542 335786 -6306
rect 336022 -6542 371786 -6306
rect 372022 -6542 407786 -6306
rect 408022 -6542 443786 -6306
rect 444022 -6542 479786 -6306
rect 480022 -6542 515786 -6306
rect 516022 -6542 551786 -6306
rect 552022 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect -7636 -6564 591560 -6542
rect -7636 -6566 -7036 -6564
rect 11604 -6566 12204 -6564
rect 47604 -6566 48204 -6564
rect 83604 -6566 84204 -6564
rect 119604 -6566 120204 -6564
rect 155604 -6566 156204 -6564
rect 191604 -6566 192204 -6564
rect 227604 -6566 228204 -6564
rect 263604 -6566 264204 -6564
rect 299604 -6566 300204 -6564
rect 335604 -6566 336204 -6564
rect 371604 -6566 372204 -6564
rect 407604 -6566 408204 -6564
rect 443604 -6566 444204 -6564
rect 479604 -6566 480204 -6564
rect 515604 -6566 516204 -6564
rect 551604 -6566 552204 -6564
rect 590960 -6566 591560 -6564
rect -8576 -6904 -7976 -6902
rect 29604 -6904 30204 -6902
rect 65604 -6904 66204 -6902
rect 101604 -6904 102204 -6902
rect 137604 -6904 138204 -6902
rect 173604 -6904 174204 -6902
rect 209604 -6904 210204 -6902
rect 245604 -6904 246204 -6902
rect 281604 -6904 282204 -6902
rect 317604 -6904 318204 -6902
rect 353604 -6904 354204 -6902
rect 389604 -6904 390204 -6902
rect 425604 -6904 426204 -6902
rect 461604 -6904 462204 -6902
rect 497604 -6904 498204 -6902
rect 533604 -6904 534204 -6902
rect 569604 -6904 570204 -6902
rect 591900 -6904 592500 -6902
rect -8576 -6926 592500 -6904
rect -8576 -7162 -8394 -6926
rect -8158 -7162 29786 -6926
rect 30022 -7162 65786 -6926
rect 66022 -7162 101786 -6926
rect 102022 -7162 137786 -6926
rect 138022 -7162 173786 -6926
rect 174022 -7162 209786 -6926
rect 210022 -7162 245786 -6926
rect 246022 -7162 281786 -6926
rect 282022 -7162 317786 -6926
rect 318022 -7162 353786 -6926
rect 354022 -7162 389786 -6926
rect 390022 -7162 425786 -6926
rect 426022 -7162 461786 -6926
rect 462022 -7162 497786 -6926
rect 498022 -7162 533786 -6926
rect 534022 -7162 569786 -6926
rect 570022 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect -8576 -7246 592500 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 29786 -7246
rect 30022 -7482 65786 -7246
rect 66022 -7482 101786 -7246
rect 102022 -7482 137786 -7246
rect 138022 -7482 173786 -7246
rect 174022 -7482 209786 -7246
rect 210022 -7482 245786 -7246
rect 246022 -7482 281786 -7246
rect 282022 -7482 317786 -7246
rect 318022 -7482 353786 -7246
rect 354022 -7482 389786 -7246
rect 390022 -7482 425786 -7246
rect 426022 -7482 461786 -7246
rect 462022 -7482 497786 -7246
rect 498022 -7482 533786 -7246
rect 534022 -7482 569786 -7246
rect 570022 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect -8576 -7504 592500 -7482
rect -8576 -7506 -7976 -7504
rect 29604 -7506 30204 -7504
rect 65604 -7506 66204 -7504
rect 101604 -7506 102204 -7504
rect 137604 -7506 138204 -7504
rect 173604 -7506 174204 -7504
rect 209604 -7506 210204 -7504
rect 245604 -7506 246204 -7504
rect 281604 -7506 282204 -7504
rect 317604 -7506 318204 -7504
rect 353604 -7506 354204 -7504
rect 389604 -7506 390204 -7504
rect 425604 -7506 426204 -7504
rect 461604 -7506 462204 -7504
rect 497604 -7506 498204 -7504
rect 533604 -7506 534204 -7504
rect 569604 -7506 570204 -7504
rect 591900 -7506 592500 -7504
use sram_1rw1r_32_256_8_sky130  sram3
timestamp 1608446478
transform -1 0 417296 0 -1 411247
box 0 0 77296 91247
use sram_1rw1r_32_256_8_sky130  sram2
timestamp 1608446478
transform 1 0 310000 0 1 560000
box 0 0 77296 91247
use sram_1rw1r_32_256_8_sky130  sram1
timestamp 1608446478
transform 1 0 190000 0 1 560000
box 0 0 77296 91247
use sram_1rw1r_32_256_8_sky130  sram0
timestamp 1608446478
transform 1 0 60000 0 1 560000
box 0 0 77296 91247
use hs32_core1  core1
timestamp 1608446478
transform 1 0 60000 0 1 320000
box 0 0 220000 220000
<< labels >>
rlabel metal3 s 583520 5796 584960 6036 6 analog_io[0]
port 0 nsew default bidirectional
rlabel metal3 s 583520 474996 584960 475236 6 analog_io[10]
port 1 nsew default bidirectional
rlabel metal3 s 583520 521916 584960 522156 6 analog_io[11]
port 2 nsew default bidirectional
rlabel metal3 s 583520 568836 584960 569076 6 analog_io[12]
port 3 nsew default bidirectional
rlabel metal3 s 583520 615756 584960 615996 6 analog_io[13]
port 4 nsew default bidirectional
rlabel metal3 s 583520 662676 584960 662916 6 analog_io[14]
port 5 nsew default bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[15]
port 6 nsew default bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[16]
port 7 nsew default bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[17]
port 8 nsew default bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[18]
port 9 nsew default bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[19]
port 10 nsew default bidirectional
rlabel metal3 s 583520 52716 584960 52956 6 analog_io[1]
port 11 nsew default bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[20]
port 12 nsew default bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[21]
port 13 nsew default bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[22]
port 14 nsew default bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[23]
port 15 nsew default bidirectional
rlabel metal3 s -960 696540 480 696780 4 analog_io[24]
port 16 nsew default bidirectional
rlabel metal3 s -960 639012 480 639252 4 analog_io[25]
port 17 nsew default bidirectional
rlabel metal3 s -960 581620 480 581860 4 analog_io[26]
port 18 nsew default bidirectional
rlabel metal3 s -960 524092 480 524332 4 analog_io[27]
port 19 nsew default bidirectional
rlabel metal3 s -960 466700 480 466940 4 analog_io[28]
port 20 nsew default bidirectional
rlabel metal3 s -960 409172 480 409412 4 analog_io[29]
port 21 nsew default bidirectional
rlabel metal3 s 583520 99636 584960 99876 6 analog_io[2]
port 22 nsew default bidirectional
rlabel metal3 s -960 351780 480 352020 4 analog_io[30]
port 23 nsew default bidirectional
rlabel metal3 s 583520 146556 584960 146796 6 analog_io[3]
port 24 nsew default bidirectional
rlabel metal3 s 583520 193476 584960 193716 6 analog_io[4]
port 25 nsew default bidirectional
rlabel metal3 s 583520 240396 584960 240636 6 analog_io[5]
port 26 nsew default bidirectional
rlabel metal3 s 583520 287316 584960 287556 6 analog_io[6]
port 27 nsew default bidirectional
rlabel metal3 s 583520 334236 584960 334476 6 analog_io[7]
port 28 nsew default bidirectional
rlabel metal3 s 583520 381156 584960 381396 6 analog_io[8]
port 29 nsew default bidirectional
rlabel metal3 s 583520 428076 584960 428316 6 analog_io[9]
port 30 nsew default bidirectional
rlabel metal3 s 583520 17492 584960 17732 6 io_in[0]
port 31 nsew default input
rlabel metal3 s 583520 486692 584960 486932 6 io_in[10]
port 32 nsew default input
rlabel metal3 s 583520 533748 584960 533988 6 io_in[11]
port 33 nsew default input
rlabel metal3 s 583520 580668 584960 580908 6 io_in[12]
port 34 nsew default input
rlabel metal3 s 583520 627588 584960 627828 6 io_in[13]
port 35 nsew default input
rlabel metal3 s 583520 674508 584960 674748 6 io_in[14]
port 36 nsew default input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 37 nsew default input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 38 nsew default input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 39 nsew default input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 40 nsew default input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 41 nsew default input
rlabel metal3 s 583520 64412 584960 64652 6 io_in[1]
port 42 nsew default input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 43 nsew default input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 44 nsew default input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 45 nsew default input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 46 nsew default input
rlabel metal3 s -960 682124 480 682364 4 io_in[24]
port 47 nsew default input
rlabel metal3 s -960 624732 480 624972 4 io_in[25]
port 48 nsew default input
rlabel metal3 s -960 567204 480 567444 4 io_in[26]
port 49 nsew default input
rlabel metal3 s -960 509812 480 510052 4 io_in[27]
port 50 nsew default input
rlabel metal3 s -960 452284 480 452524 4 io_in[28]
port 51 nsew default input
rlabel metal3 s -960 394892 480 395132 4 io_in[29]
port 52 nsew default input
rlabel metal3 s 583520 111332 584960 111572 6 io_in[2]
port 53 nsew default input
rlabel metal3 s -960 337364 480 337604 4 io_in[30]
port 54 nsew default input
rlabel metal3 s -960 294252 480 294492 4 io_in[31]
port 55 nsew default input
rlabel metal3 s -960 251140 480 251380 4 io_in[32]
port 56 nsew default input
rlabel metal3 s -960 208028 480 208268 4 io_in[33]
port 57 nsew default input
rlabel metal3 s -960 164916 480 165156 4 io_in[34]
port 58 nsew default input
rlabel metal3 s -960 121940 480 122180 4 io_in[35]
port 59 nsew default input
rlabel metal3 s -960 78828 480 79068 4 io_in[36]
port 60 nsew default input
rlabel metal3 s -960 35716 480 35956 4 io_in[37]
port 61 nsew default input
rlabel metal3 s 583520 158252 584960 158492 6 io_in[3]
port 62 nsew default input
rlabel metal3 s 583520 205172 584960 205412 6 io_in[4]
port 63 nsew default input
rlabel metal3 s 583520 252092 584960 252332 6 io_in[5]
port 64 nsew default input
rlabel metal3 s 583520 299012 584960 299252 6 io_in[6]
port 65 nsew default input
rlabel metal3 s 583520 345932 584960 346172 6 io_in[7]
port 66 nsew default input
rlabel metal3 s 583520 392852 584960 393092 6 io_in[8]
port 67 nsew default input
rlabel metal3 s 583520 439772 584960 440012 6 io_in[9]
port 68 nsew default input
rlabel metal3 s 583520 40884 584960 41124 6 io_oeb[0]
port 69 nsew default tristate
rlabel metal3 s 583520 510220 584960 510460 6 io_oeb[10]
port 70 nsew default tristate
rlabel metal3 s 583520 557140 584960 557380 6 io_oeb[11]
port 71 nsew default tristate
rlabel metal3 s 583520 604060 584960 604300 6 io_oeb[12]
port 72 nsew default tristate
rlabel metal3 s 583520 650980 584960 651220 6 io_oeb[13]
port 73 nsew default tristate
rlabel metal3 s 583520 697900 584960 698140 6 io_oeb[14]
port 74 nsew default tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 75 nsew default tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 76 nsew default tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 77 nsew default tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 78 nsew default tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 79 nsew default tristate
rlabel metal3 s 583520 87804 584960 88044 6 io_oeb[1]
port 80 nsew default tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 81 nsew default tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 82 nsew default tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 83 nsew default tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 84 nsew default tristate
rlabel metal3 s -960 653428 480 653668 4 io_oeb[24]
port 85 nsew default tristate
rlabel metal3 s -960 595900 480 596140 4 io_oeb[25]
port 86 nsew default tristate
rlabel metal3 s -960 538508 480 538748 4 io_oeb[26]
port 87 nsew default tristate
rlabel metal3 s -960 480980 480 481220 4 io_oeb[27]
port 88 nsew default tristate
rlabel metal3 s -960 423588 480 423828 4 io_oeb[28]
port 89 nsew default tristate
rlabel metal3 s -960 366060 480 366300 4 io_oeb[29]
port 90 nsew default tristate
rlabel metal3 s 583520 134724 584960 134964 6 io_oeb[2]
port 91 nsew default tristate
rlabel metal3 s -960 308668 480 308908 4 io_oeb[30]
port 92 nsew default tristate
rlabel metal3 s -960 265556 480 265796 4 io_oeb[31]
port 93 nsew default tristate
rlabel metal3 s -960 222444 480 222684 4 io_oeb[32]
port 94 nsew default tristate
rlabel metal3 s -960 179332 480 179572 4 io_oeb[33]
port 95 nsew default tristate
rlabel metal3 s -960 136220 480 136460 4 io_oeb[34]
port 96 nsew default tristate
rlabel metal3 s -960 93108 480 93348 4 io_oeb[35]
port 97 nsew default tristate
rlabel metal3 s -960 49996 480 50236 4 io_oeb[36]
port 98 nsew default tristate
rlabel metal3 s -960 7020 480 7260 4 io_oeb[37]
port 99 nsew default tristate
rlabel metal3 s 583520 181780 584960 182020 6 io_oeb[3]
port 100 nsew default tristate
rlabel metal3 s 583520 228700 584960 228940 6 io_oeb[4]
port 101 nsew default tristate
rlabel metal3 s 583520 275620 584960 275860 6 io_oeb[5]
port 102 nsew default tristate
rlabel metal3 s 583520 322540 584960 322780 6 io_oeb[6]
port 103 nsew default tristate
rlabel metal3 s 583520 369460 584960 369700 6 io_oeb[7]
port 104 nsew default tristate
rlabel metal3 s 583520 416380 584960 416620 6 io_oeb[8]
port 105 nsew default tristate
rlabel metal3 s 583520 463300 584960 463540 6 io_oeb[9]
port 106 nsew default tristate
rlabel metal3 s 583520 29188 584960 29428 6 io_out[0]
port 107 nsew default tristate
rlabel metal3 s 583520 498524 584960 498764 6 io_out[10]
port 108 nsew default tristate
rlabel metal3 s 583520 545444 584960 545684 6 io_out[11]
port 109 nsew default tristate
rlabel metal3 s 583520 592364 584960 592604 6 io_out[12]
port 110 nsew default tristate
rlabel metal3 s 583520 639284 584960 639524 6 io_out[13]
port 111 nsew default tristate
rlabel metal3 s 583520 686204 584960 686444 6 io_out[14]
port 112 nsew default tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 113 nsew default tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 114 nsew default tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 115 nsew default tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 116 nsew default tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 117 nsew default tristate
rlabel metal3 s 583520 76108 584960 76348 6 io_out[1]
port 118 nsew default tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 119 nsew default tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 120 nsew default tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 121 nsew default tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 122 nsew default tristate
rlabel metal3 s -960 667844 480 668084 4 io_out[24]
port 123 nsew default tristate
rlabel metal3 s -960 610316 480 610556 4 io_out[25]
port 124 nsew default tristate
rlabel metal3 s -960 552924 480 553164 4 io_out[26]
port 125 nsew default tristate
rlabel metal3 s -960 495396 480 495636 4 io_out[27]
port 126 nsew default tristate
rlabel metal3 s -960 437868 480 438108 4 io_out[28]
port 127 nsew default tristate
rlabel metal3 s -960 380476 480 380716 4 io_out[29]
port 128 nsew default tristate
rlabel metal3 s 583520 123028 584960 123268 6 io_out[2]
port 129 nsew default tristate
rlabel metal3 s -960 322948 480 323188 4 io_out[30]
port 130 nsew default tristate
rlabel metal3 s -960 279972 480 280212 4 io_out[31]
port 131 nsew default tristate
rlabel metal3 s -960 236860 480 237100 4 io_out[32]
port 132 nsew default tristate
rlabel metal3 s -960 193748 480 193988 4 io_out[33]
port 133 nsew default tristate
rlabel metal3 s -960 150636 480 150876 4 io_out[34]
port 134 nsew default tristate
rlabel metal3 s -960 107524 480 107764 4 io_out[35]
port 135 nsew default tristate
rlabel metal3 s -960 64412 480 64652 4 io_out[36]
port 136 nsew default tristate
rlabel metal3 s -960 21300 480 21540 4 io_out[37]
port 137 nsew default tristate
rlabel metal3 s 583520 169948 584960 170188 6 io_out[3]
port 138 nsew default tristate
rlabel metal3 s 583520 216868 584960 217108 6 io_out[4]
port 139 nsew default tristate
rlabel metal3 s 583520 263788 584960 264028 6 io_out[5]
port 140 nsew default tristate
rlabel metal3 s 583520 310708 584960 310948 6 io_out[6]
port 141 nsew default tristate
rlabel metal3 s 583520 357764 584960 358004 6 io_out[7]
port 142 nsew default tristate
rlabel metal3 s 583520 404684 584960 404924 6 io_out[8]
port 143 nsew default tristate
rlabel metal3 s 583520 451604 584960 451844 6 io_out[9]
port 144 nsew default tristate
rlabel metal2 s 126582 -960 126694 480 8 la_data_in[0]
port 145 nsew default input
rlabel metal2 s 483450 -960 483562 480 8 la_data_in[100]
port 146 nsew default input
rlabel metal2 s 486946 -960 487058 480 8 la_data_in[101]
port 147 nsew default input
rlabel metal2 s 490534 -960 490646 480 8 la_data_in[102]
port 148 nsew default input
rlabel metal2 s 494122 -960 494234 480 8 la_data_in[103]
port 149 nsew default input
rlabel metal2 s 497710 -960 497822 480 8 la_data_in[104]
port 150 nsew default input
rlabel metal2 s 501206 -960 501318 480 8 la_data_in[105]
port 151 nsew default input
rlabel metal2 s 504794 -960 504906 480 8 la_data_in[106]
port 152 nsew default input
rlabel metal2 s 508382 -960 508494 480 8 la_data_in[107]
port 153 nsew default input
rlabel metal2 s 511970 -960 512082 480 8 la_data_in[108]
port 154 nsew default input
rlabel metal2 s 515558 -960 515670 480 8 la_data_in[109]
port 155 nsew default input
rlabel metal2 s 162278 -960 162390 480 8 la_data_in[10]
port 156 nsew default input
rlabel metal2 s 519054 -960 519166 480 8 la_data_in[110]
port 157 nsew default input
rlabel metal2 s 522642 -960 522754 480 8 la_data_in[111]
port 158 nsew default input
rlabel metal2 s 526230 -960 526342 480 8 la_data_in[112]
port 159 nsew default input
rlabel metal2 s 529818 -960 529930 480 8 la_data_in[113]
port 160 nsew default input
rlabel metal2 s 533406 -960 533518 480 8 la_data_in[114]
port 161 nsew default input
rlabel metal2 s 536902 -960 537014 480 8 la_data_in[115]
port 162 nsew default input
rlabel metal2 s 540490 -960 540602 480 8 la_data_in[116]
port 163 nsew default input
rlabel metal2 s 544078 -960 544190 480 8 la_data_in[117]
port 164 nsew default input
rlabel metal2 s 547666 -960 547778 480 8 la_data_in[118]
port 165 nsew default input
rlabel metal2 s 551162 -960 551274 480 8 la_data_in[119]
port 166 nsew default input
rlabel metal2 s 165866 -960 165978 480 8 la_data_in[11]
port 167 nsew default input
rlabel metal2 s 554750 -960 554862 480 8 la_data_in[120]
port 168 nsew default input
rlabel metal2 s 558338 -960 558450 480 8 la_data_in[121]
port 169 nsew default input
rlabel metal2 s 561926 -960 562038 480 8 la_data_in[122]
port 170 nsew default input
rlabel metal2 s 565514 -960 565626 480 8 la_data_in[123]
port 171 nsew default input
rlabel metal2 s 569010 -960 569122 480 8 la_data_in[124]
port 172 nsew default input
rlabel metal2 s 572598 -960 572710 480 8 la_data_in[125]
port 173 nsew default input
rlabel metal2 s 576186 -960 576298 480 8 la_data_in[126]
port 174 nsew default input
rlabel metal2 s 579774 -960 579886 480 8 la_data_in[127]
port 175 nsew default input
rlabel metal2 s 169362 -960 169474 480 8 la_data_in[12]
port 176 nsew default input
rlabel metal2 s 172950 -960 173062 480 8 la_data_in[13]
port 177 nsew default input
rlabel metal2 s 176538 -960 176650 480 8 la_data_in[14]
port 178 nsew default input
rlabel metal2 s 180126 -960 180238 480 8 la_data_in[15]
port 179 nsew default input
rlabel metal2 s 183714 -960 183826 480 8 la_data_in[16]
port 180 nsew default input
rlabel metal2 s 187210 -960 187322 480 8 la_data_in[17]
port 181 nsew default input
rlabel metal2 s 190798 -960 190910 480 8 la_data_in[18]
port 182 nsew default input
rlabel metal2 s 194386 -960 194498 480 8 la_data_in[19]
port 183 nsew default input
rlabel metal2 s 130170 -960 130282 480 8 la_data_in[1]
port 184 nsew default input
rlabel metal2 s 197974 -960 198086 480 8 la_data_in[20]
port 185 nsew default input
rlabel metal2 s 201470 -960 201582 480 8 la_data_in[21]
port 186 nsew default input
rlabel metal2 s 205058 -960 205170 480 8 la_data_in[22]
port 187 nsew default input
rlabel metal2 s 208646 -960 208758 480 8 la_data_in[23]
port 188 nsew default input
rlabel metal2 s 212234 -960 212346 480 8 la_data_in[24]
port 189 nsew default input
rlabel metal2 s 215822 -960 215934 480 8 la_data_in[25]
port 190 nsew default input
rlabel metal2 s 219318 -960 219430 480 8 la_data_in[26]
port 191 nsew default input
rlabel metal2 s 222906 -960 223018 480 8 la_data_in[27]
port 192 nsew default input
rlabel metal2 s 226494 -960 226606 480 8 la_data_in[28]
port 193 nsew default input
rlabel metal2 s 230082 -960 230194 480 8 la_data_in[29]
port 194 nsew default input
rlabel metal2 s 133758 -960 133870 480 8 la_data_in[2]
port 195 nsew default input
rlabel metal2 s 233670 -960 233782 480 8 la_data_in[30]
port 196 nsew default input
rlabel metal2 s 237166 -960 237278 480 8 la_data_in[31]
port 197 nsew default input
rlabel metal2 s 240754 -960 240866 480 8 la_data_in[32]
port 198 nsew default input
rlabel metal2 s 244342 -960 244454 480 8 la_data_in[33]
port 199 nsew default input
rlabel metal2 s 247930 -960 248042 480 8 la_data_in[34]
port 200 nsew default input
rlabel metal2 s 251426 -960 251538 480 8 la_data_in[35]
port 201 nsew default input
rlabel metal2 s 255014 -960 255126 480 8 la_data_in[36]
port 202 nsew default input
rlabel metal2 s 258602 -960 258714 480 8 la_data_in[37]
port 203 nsew default input
rlabel metal2 s 262190 -960 262302 480 8 la_data_in[38]
port 204 nsew default input
rlabel metal2 s 265778 -960 265890 480 8 la_data_in[39]
port 205 nsew default input
rlabel metal2 s 137254 -960 137366 480 8 la_data_in[3]
port 206 nsew default input
rlabel metal2 s 269274 -960 269386 480 8 la_data_in[40]
port 207 nsew default input
rlabel metal2 s 272862 -960 272974 480 8 la_data_in[41]
port 208 nsew default input
rlabel metal2 s 276450 -960 276562 480 8 la_data_in[42]
port 209 nsew default input
rlabel metal2 s 280038 -960 280150 480 8 la_data_in[43]
port 210 nsew default input
rlabel metal2 s 283626 -960 283738 480 8 la_data_in[44]
port 211 nsew default input
rlabel metal2 s 287122 -960 287234 480 8 la_data_in[45]
port 212 nsew default input
rlabel metal2 s 290710 -960 290822 480 8 la_data_in[46]
port 213 nsew default input
rlabel metal2 s 294298 -960 294410 480 8 la_data_in[47]
port 214 nsew default input
rlabel metal2 s 297886 -960 297998 480 8 la_data_in[48]
port 215 nsew default input
rlabel metal2 s 301382 -960 301494 480 8 la_data_in[49]
port 216 nsew default input
rlabel metal2 s 140842 -960 140954 480 8 la_data_in[4]
port 217 nsew default input
rlabel metal2 s 304970 -960 305082 480 8 la_data_in[50]
port 218 nsew default input
rlabel metal2 s 308558 -960 308670 480 8 la_data_in[51]
port 219 nsew default input
rlabel metal2 s 312146 -960 312258 480 8 la_data_in[52]
port 220 nsew default input
rlabel metal2 s 315734 -960 315846 480 8 la_data_in[53]
port 221 nsew default input
rlabel metal2 s 319230 -960 319342 480 8 la_data_in[54]
port 222 nsew default input
rlabel metal2 s 322818 -960 322930 480 8 la_data_in[55]
port 223 nsew default input
rlabel metal2 s 326406 -960 326518 480 8 la_data_in[56]
port 224 nsew default input
rlabel metal2 s 329994 -960 330106 480 8 la_data_in[57]
port 225 nsew default input
rlabel metal2 s 333582 -960 333694 480 8 la_data_in[58]
port 226 nsew default input
rlabel metal2 s 337078 -960 337190 480 8 la_data_in[59]
port 227 nsew default input
rlabel metal2 s 144430 -960 144542 480 8 la_data_in[5]
port 228 nsew default input
rlabel metal2 s 340666 -960 340778 480 8 la_data_in[60]
port 229 nsew default input
rlabel metal2 s 344254 -960 344366 480 8 la_data_in[61]
port 230 nsew default input
rlabel metal2 s 347842 -960 347954 480 8 la_data_in[62]
port 231 nsew default input
rlabel metal2 s 351338 -960 351450 480 8 la_data_in[63]
port 232 nsew default input
rlabel metal2 s 354926 -960 355038 480 8 la_data_in[64]
port 233 nsew default input
rlabel metal2 s 358514 -960 358626 480 8 la_data_in[65]
port 234 nsew default input
rlabel metal2 s 362102 -960 362214 480 8 la_data_in[66]
port 235 nsew default input
rlabel metal2 s 365690 -960 365802 480 8 la_data_in[67]
port 236 nsew default input
rlabel metal2 s 369186 -960 369298 480 8 la_data_in[68]
port 237 nsew default input
rlabel metal2 s 372774 -960 372886 480 8 la_data_in[69]
port 238 nsew default input
rlabel metal2 s 148018 -960 148130 480 8 la_data_in[6]
port 239 nsew default input
rlabel metal2 s 376362 -960 376474 480 8 la_data_in[70]
port 240 nsew default input
rlabel metal2 s 379950 -960 380062 480 8 la_data_in[71]
port 241 nsew default input
rlabel metal2 s 383538 -960 383650 480 8 la_data_in[72]
port 242 nsew default input
rlabel metal2 s 387034 -960 387146 480 8 la_data_in[73]
port 243 nsew default input
rlabel metal2 s 390622 -960 390734 480 8 la_data_in[74]
port 244 nsew default input
rlabel metal2 s 394210 -960 394322 480 8 la_data_in[75]
port 245 nsew default input
rlabel metal2 s 397798 -960 397910 480 8 la_data_in[76]
port 246 nsew default input
rlabel metal2 s 401294 -960 401406 480 8 la_data_in[77]
port 247 nsew default input
rlabel metal2 s 404882 -960 404994 480 8 la_data_in[78]
port 248 nsew default input
rlabel metal2 s 408470 -960 408582 480 8 la_data_in[79]
port 249 nsew default input
rlabel metal2 s 151514 -960 151626 480 8 la_data_in[7]
port 250 nsew default input
rlabel metal2 s 412058 -960 412170 480 8 la_data_in[80]
port 251 nsew default input
rlabel metal2 s 415646 -960 415758 480 8 la_data_in[81]
port 252 nsew default input
rlabel metal2 s 419142 -960 419254 480 8 la_data_in[82]
port 253 nsew default input
rlabel metal2 s 422730 -960 422842 480 8 la_data_in[83]
port 254 nsew default input
rlabel metal2 s 426318 -960 426430 480 8 la_data_in[84]
port 255 nsew default input
rlabel metal2 s 429906 -960 430018 480 8 la_data_in[85]
port 256 nsew default input
rlabel metal2 s 433494 -960 433606 480 8 la_data_in[86]
port 257 nsew default input
rlabel metal2 s 436990 -960 437102 480 8 la_data_in[87]
port 258 nsew default input
rlabel metal2 s 440578 -960 440690 480 8 la_data_in[88]
port 259 nsew default input
rlabel metal2 s 444166 -960 444278 480 8 la_data_in[89]
port 260 nsew default input
rlabel metal2 s 155102 -960 155214 480 8 la_data_in[8]
port 261 nsew default input
rlabel metal2 s 447754 -960 447866 480 8 la_data_in[90]
port 262 nsew default input
rlabel metal2 s 451250 -960 451362 480 8 la_data_in[91]
port 263 nsew default input
rlabel metal2 s 454838 -960 454950 480 8 la_data_in[92]
port 264 nsew default input
rlabel metal2 s 458426 -960 458538 480 8 la_data_in[93]
port 265 nsew default input
rlabel metal2 s 462014 -960 462126 480 8 la_data_in[94]
port 266 nsew default input
rlabel metal2 s 465602 -960 465714 480 8 la_data_in[95]
port 267 nsew default input
rlabel metal2 s 469098 -960 469210 480 8 la_data_in[96]
port 268 nsew default input
rlabel metal2 s 472686 -960 472798 480 8 la_data_in[97]
port 269 nsew default input
rlabel metal2 s 476274 -960 476386 480 8 la_data_in[98]
port 270 nsew default input
rlabel metal2 s 479862 -960 479974 480 8 la_data_in[99]
port 271 nsew default input
rlabel metal2 s 158690 -960 158802 480 8 la_data_in[9]
port 272 nsew default input
rlabel metal2 s 127778 -960 127890 480 8 la_data_out[0]
port 273 nsew default tristate
rlabel metal2 s 484554 -960 484666 480 8 la_data_out[100]
port 274 nsew default tristate
rlabel metal2 s 488142 -960 488254 480 8 la_data_out[101]
port 275 nsew default tristate
rlabel metal2 s 491730 -960 491842 480 8 la_data_out[102]
port 276 nsew default tristate
rlabel metal2 s 495318 -960 495430 480 8 la_data_out[103]
port 277 nsew default tristate
rlabel metal2 s 498906 -960 499018 480 8 la_data_out[104]
port 278 nsew default tristate
rlabel metal2 s 502402 -960 502514 480 8 la_data_out[105]
port 279 nsew default tristate
rlabel metal2 s 505990 -960 506102 480 8 la_data_out[106]
port 280 nsew default tristate
rlabel metal2 s 509578 -960 509690 480 8 la_data_out[107]
port 281 nsew default tristate
rlabel metal2 s 513166 -960 513278 480 8 la_data_out[108]
port 282 nsew default tristate
rlabel metal2 s 516754 -960 516866 480 8 la_data_out[109]
port 283 nsew default tristate
rlabel metal2 s 163474 -960 163586 480 8 la_data_out[10]
port 284 nsew default tristate
rlabel metal2 s 520250 -960 520362 480 8 la_data_out[110]
port 285 nsew default tristate
rlabel metal2 s 523838 -960 523950 480 8 la_data_out[111]
port 286 nsew default tristate
rlabel metal2 s 527426 -960 527538 480 8 la_data_out[112]
port 287 nsew default tristate
rlabel metal2 s 531014 -960 531126 480 8 la_data_out[113]
port 288 nsew default tristate
rlabel metal2 s 534510 -960 534622 480 8 la_data_out[114]
port 289 nsew default tristate
rlabel metal2 s 538098 -960 538210 480 8 la_data_out[115]
port 290 nsew default tristate
rlabel metal2 s 541686 -960 541798 480 8 la_data_out[116]
port 291 nsew default tristate
rlabel metal2 s 545274 -960 545386 480 8 la_data_out[117]
port 292 nsew default tristate
rlabel metal2 s 548862 -960 548974 480 8 la_data_out[118]
port 293 nsew default tristate
rlabel metal2 s 552358 -960 552470 480 8 la_data_out[119]
port 294 nsew default tristate
rlabel metal2 s 167062 -960 167174 480 8 la_data_out[11]
port 295 nsew default tristate
rlabel metal2 s 555946 -960 556058 480 8 la_data_out[120]
port 296 nsew default tristate
rlabel metal2 s 559534 -960 559646 480 8 la_data_out[121]
port 297 nsew default tristate
rlabel metal2 s 563122 -960 563234 480 8 la_data_out[122]
port 298 nsew default tristate
rlabel metal2 s 566710 -960 566822 480 8 la_data_out[123]
port 299 nsew default tristate
rlabel metal2 s 570206 -960 570318 480 8 la_data_out[124]
port 300 nsew default tristate
rlabel metal2 s 573794 -960 573906 480 8 la_data_out[125]
port 301 nsew default tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[126]
port 302 nsew default tristate
rlabel metal2 s 580970 -960 581082 480 8 la_data_out[127]
port 303 nsew default tristate
rlabel metal2 s 170558 -960 170670 480 8 la_data_out[12]
port 304 nsew default tristate
rlabel metal2 s 174146 -960 174258 480 8 la_data_out[13]
port 305 nsew default tristate
rlabel metal2 s 177734 -960 177846 480 8 la_data_out[14]
port 306 nsew default tristate
rlabel metal2 s 181322 -960 181434 480 8 la_data_out[15]
port 307 nsew default tristate
rlabel metal2 s 184818 -960 184930 480 8 la_data_out[16]
port 308 nsew default tristate
rlabel metal2 s 188406 -960 188518 480 8 la_data_out[17]
port 309 nsew default tristate
rlabel metal2 s 191994 -960 192106 480 8 la_data_out[18]
port 310 nsew default tristate
rlabel metal2 s 195582 -960 195694 480 8 la_data_out[19]
port 311 nsew default tristate
rlabel metal2 s 131366 -960 131478 480 8 la_data_out[1]
port 312 nsew default tristate
rlabel metal2 s 199170 -960 199282 480 8 la_data_out[20]
port 313 nsew default tristate
rlabel metal2 s 202666 -960 202778 480 8 la_data_out[21]
port 314 nsew default tristate
rlabel metal2 s 206254 -960 206366 480 8 la_data_out[22]
port 315 nsew default tristate
rlabel metal2 s 209842 -960 209954 480 8 la_data_out[23]
port 316 nsew default tristate
rlabel metal2 s 213430 -960 213542 480 8 la_data_out[24]
port 317 nsew default tristate
rlabel metal2 s 217018 -960 217130 480 8 la_data_out[25]
port 318 nsew default tristate
rlabel metal2 s 220514 -960 220626 480 8 la_data_out[26]
port 319 nsew default tristate
rlabel metal2 s 224102 -960 224214 480 8 la_data_out[27]
port 320 nsew default tristate
rlabel metal2 s 227690 -960 227802 480 8 la_data_out[28]
port 321 nsew default tristate
rlabel metal2 s 231278 -960 231390 480 8 la_data_out[29]
port 322 nsew default tristate
rlabel metal2 s 134862 -960 134974 480 8 la_data_out[2]
port 323 nsew default tristate
rlabel metal2 s 234774 -960 234886 480 8 la_data_out[30]
port 324 nsew default tristate
rlabel metal2 s 238362 -960 238474 480 8 la_data_out[31]
port 325 nsew default tristate
rlabel metal2 s 241950 -960 242062 480 8 la_data_out[32]
port 326 nsew default tristate
rlabel metal2 s 245538 -960 245650 480 8 la_data_out[33]
port 327 nsew default tristate
rlabel metal2 s 249126 -960 249238 480 8 la_data_out[34]
port 328 nsew default tristate
rlabel metal2 s 252622 -960 252734 480 8 la_data_out[35]
port 329 nsew default tristate
rlabel metal2 s 256210 -960 256322 480 8 la_data_out[36]
port 330 nsew default tristate
rlabel metal2 s 259798 -960 259910 480 8 la_data_out[37]
port 331 nsew default tristate
rlabel metal2 s 263386 -960 263498 480 8 la_data_out[38]
port 332 nsew default tristate
rlabel metal2 s 266974 -960 267086 480 8 la_data_out[39]
port 333 nsew default tristate
rlabel metal2 s 138450 -960 138562 480 8 la_data_out[3]
port 334 nsew default tristate
rlabel metal2 s 270470 -960 270582 480 8 la_data_out[40]
port 335 nsew default tristate
rlabel metal2 s 274058 -960 274170 480 8 la_data_out[41]
port 336 nsew default tristate
rlabel metal2 s 277646 -960 277758 480 8 la_data_out[42]
port 337 nsew default tristate
rlabel metal2 s 281234 -960 281346 480 8 la_data_out[43]
port 338 nsew default tristate
rlabel metal2 s 284730 -960 284842 480 8 la_data_out[44]
port 339 nsew default tristate
rlabel metal2 s 288318 -960 288430 480 8 la_data_out[45]
port 340 nsew default tristate
rlabel metal2 s 291906 -960 292018 480 8 la_data_out[46]
port 341 nsew default tristate
rlabel metal2 s 295494 -960 295606 480 8 la_data_out[47]
port 342 nsew default tristate
rlabel metal2 s 299082 -960 299194 480 8 la_data_out[48]
port 343 nsew default tristate
rlabel metal2 s 302578 -960 302690 480 8 la_data_out[49]
port 344 nsew default tristate
rlabel metal2 s 142038 -960 142150 480 8 la_data_out[4]
port 345 nsew default tristate
rlabel metal2 s 306166 -960 306278 480 8 la_data_out[50]
port 346 nsew default tristate
rlabel metal2 s 309754 -960 309866 480 8 la_data_out[51]
port 347 nsew default tristate
rlabel metal2 s 313342 -960 313454 480 8 la_data_out[52]
port 348 nsew default tristate
rlabel metal2 s 316930 -960 317042 480 8 la_data_out[53]
port 349 nsew default tristate
rlabel metal2 s 320426 -960 320538 480 8 la_data_out[54]
port 350 nsew default tristate
rlabel metal2 s 324014 -960 324126 480 8 la_data_out[55]
port 351 nsew default tristate
rlabel metal2 s 327602 -960 327714 480 8 la_data_out[56]
port 352 nsew default tristate
rlabel metal2 s 331190 -960 331302 480 8 la_data_out[57]
port 353 nsew default tristate
rlabel metal2 s 334686 -960 334798 480 8 la_data_out[58]
port 354 nsew default tristate
rlabel metal2 s 338274 -960 338386 480 8 la_data_out[59]
port 355 nsew default tristate
rlabel metal2 s 145626 -960 145738 480 8 la_data_out[5]
port 356 nsew default tristate
rlabel metal2 s 341862 -960 341974 480 8 la_data_out[60]
port 357 nsew default tristate
rlabel metal2 s 345450 -960 345562 480 8 la_data_out[61]
port 358 nsew default tristate
rlabel metal2 s 349038 -960 349150 480 8 la_data_out[62]
port 359 nsew default tristate
rlabel metal2 s 352534 -960 352646 480 8 la_data_out[63]
port 360 nsew default tristate
rlabel metal2 s 356122 -960 356234 480 8 la_data_out[64]
port 361 nsew default tristate
rlabel metal2 s 359710 -960 359822 480 8 la_data_out[65]
port 362 nsew default tristate
rlabel metal2 s 363298 -960 363410 480 8 la_data_out[66]
port 363 nsew default tristate
rlabel metal2 s 366886 -960 366998 480 8 la_data_out[67]
port 364 nsew default tristate
rlabel metal2 s 370382 -960 370494 480 8 la_data_out[68]
port 365 nsew default tristate
rlabel metal2 s 373970 -960 374082 480 8 la_data_out[69]
port 366 nsew default tristate
rlabel metal2 s 149214 -960 149326 480 8 la_data_out[6]
port 367 nsew default tristate
rlabel metal2 s 377558 -960 377670 480 8 la_data_out[70]
port 368 nsew default tristate
rlabel metal2 s 381146 -960 381258 480 8 la_data_out[71]
port 369 nsew default tristate
rlabel metal2 s 384642 -960 384754 480 8 la_data_out[72]
port 370 nsew default tristate
rlabel metal2 s 388230 -960 388342 480 8 la_data_out[73]
port 371 nsew default tristate
rlabel metal2 s 391818 -960 391930 480 8 la_data_out[74]
port 372 nsew default tristate
rlabel metal2 s 395406 -960 395518 480 8 la_data_out[75]
port 373 nsew default tristate
rlabel metal2 s 398994 -960 399106 480 8 la_data_out[76]
port 374 nsew default tristate
rlabel metal2 s 402490 -960 402602 480 8 la_data_out[77]
port 375 nsew default tristate
rlabel metal2 s 406078 -960 406190 480 8 la_data_out[78]
port 376 nsew default tristate
rlabel metal2 s 409666 -960 409778 480 8 la_data_out[79]
port 377 nsew default tristate
rlabel metal2 s 152710 -960 152822 480 8 la_data_out[7]
port 378 nsew default tristate
rlabel metal2 s 413254 -960 413366 480 8 la_data_out[80]
port 379 nsew default tristate
rlabel metal2 s 416842 -960 416954 480 8 la_data_out[81]
port 380 nsew default tristate
rlabel metal2 s 420338 -960 420450 480 8 la_data_out[82]
port 381 nsew default tristate
rlabel metal2 s 423926 -960 424038 480 8 la_data_out[83]
port 382 nsew default tristate
rlabel metal2 s 427514 -960 427626 480 8 la_data_out[84]
port 383 nsew default tristate
rlabel metal2 s 431102 -960 431214 480 8 la_data_out[85]
port 384 nsew default tristate
rlabel metal2 s 434598 -960 434710 480 8 la_data_out[86]
port 385 nsew default tristate
rlabel metal2 s 438186 -960 438298 480 8 la_data_out[87]
port 386 nsew default tristate
rlabel metal2 s 441774 -960 441886 480 8 la_data_out[88]
port 387 nsew default tristate
rlabel metal2 s 445362 -960 445474 480 8 la_data_out[89]
port 388 nsew default tristate
rlabel metal2 s 156298 -960 156410 480 8 la_data_out[8]
port 389 nsew default tristate
rlabel metal2 s 448950 -960 449062 480 8 la_data_out[90]
port 390 nsew default tristate
rlabel metal2 s 452446 -960 452558 480 8 la_data_out[91]
port 391 nsew default tristate
rlabel metal2 s 456034 -960 456146 480 8 la_data_out[92]
port 392 nsew default tristate
rlabel metal2 s 459622 -960 459734 480 8 la_data_out[93]
port 393 nsew default tristate
rlabel metal2 s 463210 -960 463322 480 8 la_data_out[94]
port 394 nsew default tristate
rlabel metal2 s 466798 -960 466910 480 8 la_data_out[95]
port 395 nsew default tristate
rlabel metal2 s 470294 -960 470406 480 8 la_data_out[96]
port 396 nsew default tristate
rlabel metal2 s 473882 -960 473994 480 8 la_data_out[97]
port 397 nsew default tristate
rlabel metal2 s 477470 -960 477582 480 8 la_data_out[98]
port 398 nsew default tristate
rlabel metal2 s 481058 -960 481170 480 8 la_data_out[99]
port 399 nsew default tristate
rlabel metal2 s 159886 -960 159998 480 8 la_data_out[9]
port 400 nsew default tristate
rlabel metal2 s 128974 -960 129086 480 8 la_oen[0]
port 401 nsew default input
rlabel metal2 s 485750 -960 485862 480 8 la_oen[100]
port 402 nsew default input
rlabel metal2 s 489338 -960 489450 480 8 la_oen[101]
port 403 nsew default input
rlabel metal2 s 492926 -960 493038 480 8 la_oen[102]
port 404 nsew default input
rlabel metal2 s 496514 -960 496626 480 8 la_oen[103]
port 405 nsew default input
rlabel metal2 s 500102 -960 500214 480 8 la_oen[104]
port 406 nsew default input
rlabel metal2 s 503598 -960 503710 480 8 la_oen[105]
port 407 nsew default input
rlabel metal2 s 507186 -960 507298 480 8 la_oen[106]
port 408 nsew default input
rlabel metal2 s 510774 -960 510886 480 8 la_oen[107]
port 409 nsew default input
rlabel metal2 s 514362 -960 514474 480 8 la_oen[108]
port 410 nsew default input
rlabel metal2 s 517858 -960 517970 480 8 la_oen[109]
port 411 nsew default input
rlabel metal2 s 164670 -960 164782 480 8 la_oen[10]
port 412 nsew default input
rlabel metal2 s 521446 -960 521558 480 8 la_oen[110]
port 413 nsew default input
rlabel metal2 s 525034 -960 525146 480 8 la_oen[111]
port 414 nsew default input
rlabel metal2 s 528622 -960 528734 480 8 la_oen[112]
port 415 nsew default input
rlabel metal2 s 532210 -960 532322 480 8 la_oen[113]
port 416 nsew default input
rlabel metal2 s 535706 -960 535818 480 8 la_oen[114]
port 417 nsew default input
rlabel metal2 s 539294 -960 539406 480 8 la_oen[115]
port 418 nsew default input
rlabel metal2 s 542882 -960 542994 480 8 la_oen[116]
port 419 nsew default input
rlabel metal2 s 546470 -960 546582 480 8 la_oen[117]
port 420 nsew default input
rlabel metal2 s 550058 -960 550170 480 8 la_oen[118]
port 421 nsew default input
rlabel metal2 s 553554 -960 553666 480 8 la_oen[119]
port 422 nsew default input
rlabel metal2 s 168166 -960 168278 480 8 la_oen[11]
port 423 nsew default input
rlabel metal2 s 557142 -960 557254 480 8 la_oen[120]
port 424 nsew default input
rlabel metal2 s 560730 -960 560842 480 8 la_oen[121]
port 425 nsew default input
rlabel metal2 s 564318 -960 564430 480 8 la_oen[122]
port 426 nsew default input
rlabel metal2 s 567814 -960 567926 480 8 la_oen[123]
port 427 nsew default input
rlabel metal2 s 571402 -960 571514 480 8 la_oen[124]
port 428 nsew default input
rlabel metal2 s 574990 -960 575102 480 8 la_oen[125]
port 429 nsew default input
rlabel metal2 s 578578 -960 578690 480 8 la_oen[126]
port 430 nsew default input
rlabel metal2 s 582166 -960 582278 480 8 la_oen[127]
port 431 nsew default input
rlabel metal2 s 171754 -960 171866 480 8 la_oen[12]
port 432 nsew default input
rlabel metal2 s 175342 -960 175454 480 8 la_oen[13]
port 433 nsew default input
rlabel metal2 s 178930 -960 179042 480 8 la_oen[14]
port 434 nsew default input
rlabel metal2 s 182518 -960 182630 480 8 la_oen[15]
port 435 nsew default input
rlabel metal2 s 186014 -960 186126 480 8 la_oen[16]
port 436 nsew default input
rlabel metal2 s 189602 -960 189714 480 8 la_oen[17]
port 437 nsew default input
rlabel metal2 s 193190 -960 193302 480 8 la_oen[18]
port 438 nsew default input
rlabel metal2 s 196778 -960 196890 480 8 la_oen[19]
port 439 nsew default input
rlabel metal2 s 132562 -960 132674 480 8 la_oen[1]
port 440 nsew default input
rlabel metal2 s 200366 -960 200478 480 8 la_oen[20]
port 441 nsew default input
rlabel metal2 s 203862 -960 203974 480 8 la_oen[21]
port 442 nsew default input
rlabel metal2 s 207450 -960 207562 480 8 la_oen[22]
port 443 nsew default input
rlabel metal2 s 211038 -960 211150 480 8 la_oen[23]
port 444 nsew default input
rlabel metal2 s 214626 -960 214738 480 8 la_oen[24]
port 445 nsew default input
rlabel metal2 s 218122 -960 218234 480 8 la_oen[25]
port 446 nsew default input
rlabel metal2 s 221710 -960 221822 480 8 la_oen[26]
port 447 nsew default input
rlabel metal2 s 225298 -960 225410 480 8 la_oen[27]
port 448 nsew default input
rlabel metal2 s 228886 -960 228998 480 8 la_oen[28]
port 449 nsew default input
rlabel metal2 s 232474 -960 232586 480 8 la_oen[29]
port 450 nsew default input
rlabel metal2 s 136058 -960 136170 480 8 la_oen[2]
port 451 nsew default input
rlabel metal2 s 235970 -960 236082 480 8 la_oen[30]
port 452 nsew default input
rlabel metal2 s 239558 -960 239670 480 8 la_oen[31]
port 453 nsew default input
rlabel metal2 s 243146 -960 243258 480 8 la_oen[32]
port 454 nsew default input
rlabel metal2 s 246734 -960 246846 480 8 la_oen[33]
port 455 nsew default input
rlabel metal2 s 250322 -960 250434 480 8 la_oen[34]
port 456 nsew default input
rlabel metal2 s 253818 -960 253930 480 8 la_oen[35]
port 457 nsew default input
rlabel metal2 s 257406 -960 257518 480 8 la_oen[36]
port 458 nsew default input
rlabel metal2 s 260994 -960 261106 480 8 la_oen[37]
port 459 nsew default input
rlabel metal2 s 264582 -960 264694 480 8 la_oen[38]
port 460 nsew default input
rlabel metal2 s 268078 -960 268190 480 8 la_oen[39]
port 461 nsew default input
rlabel metal2 s 139646 -960 139758 480 8 la_oen[3]
port 462 nsew default input
rlabel metal2 s 271666 -960 271778 480 8 la_oen[40]
port 463 nsew default input
rlabel metal2 s 275254 -960 275366 480 8 la_oen[41]
port 464 nsew default input
rlabel metal2 s 278842 -960 278954 480 8 la_oen[42]
port 465 nsew default input
rlabel metal2 s 282430 -960 282542 480 8 la_oen[43]
port 466 nsew default input
rlabel metal2 s 285926 -960 286038 480 8 la_oen[44]
port 467 nsew default input
rlabel metal2 s 289514 -960 289626 480 8 la_oen[45]
port 468 nsew default input
rlabel metal2 s 293102 -960 293214 480 8 la_oen[46]
port 469 nsew default input
rlabel metal2 s 296690 -960 296802 480 8 la_oen[47]
port 470 nsew default input
rlabel metal2 s 300278 -960 300390 480 8 la_oen[48]
port 471 nsew default input
rlabel metal2 s 303774 -960 303886 480 8 la_oen[49]
port 472 nsew default input
rlabel metal2 s 143234 -960 143346 480 8 la_oen[4]
port 473 nsew default input
rlabel metal2 s 307362 -960 307474 480 8 la_oen[50]
port 474 nsew default input
rlabel metal2 s 310950 -960 311062 480 8 la_oen[51]
port 475 nsew default input
rlabel metal2 s 314538 -960 314650 480 8 la_oen[52]
port 476 nsew default input
rlabel metal2 s 318034 -960 318146 480 8 la_oen[53]
port 477 nsew default input
rlabel metal2 s 321622 -960 321734 480 8 la_oen[54]
port 478 nsew default input
rlabel metal2 s 325210 -960 325322 480 8 la_oen[55]
port 479 nsew default input
rlabel metal2 s 328798 -960 328910 480 8 la_oen[56]
port 480 nsew default input
rlabel metal2 s 332386 -960 332498 480 8 la_oen[57]
port 481 nsew default input
rlabel metal2 s 335882 -960 335994 480 8 la_oen[58]
port 482 nsew default input
rlabel metal2 s 339470 -960 339582 480 8 la_oen[59]
port 483 nsew default input
rlabel metal2 s 146822 -960 146934 480 8 la_oen[5]
port 484 nsew default input
rlabel metal2 s 343058 -960 343170 480 8 la_oen[60]
port 485 nsew default input
rlabel metal2 s 346646 -960 346758 480 8 la_oen[61]
port 486 nsew default input
rlabel metal2 s 350234 -960 350346 480 8 la_oen[62]
port 487 nsew default input
rlabel metal2 s 353730 -960 353842 480 8 la_oen[63]
port 488 nsew default input
rlabel metal2 s 357318 -960 357430 480 8 la_oen[64]
port 489 nsew default input
rlabel metal2 s 360906 -960 361018 480 8 la_oen[65]
port 490 nsew default input
rlabel metal2 s 364494 -960 364606 480 8 la_oen[66]
port 491 nsew default input
rlabel metal2 s 367990 -960 368102 480 8 la_oen[67]
port 492 nsew default input
rlabel metal2 s 371578 -960 371690 480 8 la_oen[68]
port 493 nsew default input
rlabel metal2 s 375166 -960 375278 480 8 la_oen[69]
port 494 nsew default input
rlabel metal2 s 150410 -960 150522 480 8 la_oen[6]
port 495 nsew default input
rlabel metal2 s 378754 -960 378866 480 8 la_oen[70]
port 496 nsew default input
rlabel metal2 s 382342 -960 382454 480 8 la_oen[71]
port 497 nsew default input
rlabel metal2 s 385838 -960 385950 480 8 la_oen[72]
port 498 nsew default input
rlabel metal2 s 389426 -960 389538 480 8 la_oen[73]
port 499 nsew default input
rlabel metal2 s 393014 -960 393126 480 8 la_oen[74]
port 500 nsew default input
rlabel metal2 s 396602 -960 396714 480 8 la_oen[75]
port 501 nsew default input
rlabel metal2 s 400190 -960 400302 480 8 la_oen[76]
port 502 nsew default input
rlabel metal2 s 403686 -960 403798 480 8 la_oen[77]
port 503 nsew default input
rlabel metal2 s 407274 -960 407386 480 8 la_oen[78]
port 504 nsew default input
rlabel metal2 s 410862 -960 410974 480 8 la_oen[79]
port 505 nsew default input
rlabel metal2 s 153906 -960 154018 480 8 la_oen[7]
port 506 nsew default input
rlabel metal2 s 414450 -960 414562 480 8 la_oen[80]
port 507 nsew default input
rlabel metal2 s 417946 -960 418058 480 8 la_oen[81]
port 508 nsew default input
rlabel metal2 s 421534 -960 421646 480 8 la_oen[82]
port 509 nsew default input
rlabel metal2 s 425122 -960 425234 480 8 la_oen[83]
port 510 nsew default input
rlabel metal2 s 428710 -960 428822 480 8 la_oen[84]
port 511 nsew default input
rlabel metal2 s 432298 -960 432410 480 8 la_oen[85]
port 512 nsew default input
rlabel metal2 s 435794 -960 435906 480 8 la_oen[86]
port 513 nsew default input
rlabel metal2 s 439382 -960 439494 480 8 la_oen[87]
port 514 nsew default input
rlabel metal2 s 442970 -960 443082 480 8 la_oen[88]
port 515 nsew default input
rlabel metal2 s 446558 -960 446670 480 8 la_oen[89]
port 516 nsew default input
rlabel metal2 s 157494 -960 157606 480 8 la_oen[8]
port 517 nsew default input
rlabel metal2 s 450146 -960 450258 480 8 la_oen[90]
port 518 nsew default input
rlabel metal2 s 453642 -960 453754 480 8 la_oen[91]
port 519 nsew default input
rlabel metal2 s 457230 -960 457342 480 8 la_oen[92]
port 520 nsew default input
rlabel metal2 s 460818 -960 460930 480 8 la_oen[93]
port 521 nsew default input
rlabel metal2 s 464406 -960 464518 480 8 la_oen[94]
port 522 nsew default input
rlabel metal2 s 467902 -960 468014 480 8 la_oen[95]
port 523 nsew default input
rlabel metal2 s 471490 -960 471602 480 8 la_oen[96]
port 524 nsew default input
rlabel metal2 s 475078 -960 475190 480 8 la_oen[97]
port 525 nsew default input
rlabel metal2 s 478666 -960 478778 480 8 la_oen[98]
port 526 nsew default input
rlabel metal2 s 482254 -960 482366 480 8 la_oen[99]
port 527 nsew default input
rlabel metal2 s 161082 -960 161194 480 8 la_oen[9]
port 528 nsew default input
rlabel metal2 s 583362 -960 583474 480 8 user_clock2
port 529 nsew default input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 530 nsew default input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 531 nsew default input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 532 nsew default tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 533 nsew default input
rlabel metal2 s 48106 -960 48218 480 8 wbs_adr_i[10]
port 534 nsew default input
rlabel metal2 s 51602 -960 51714 480 8 wbs_adr_i[11]
port 535 nsew default input
rlabel metal2 s 55190 -960 55302 480 8 wbs_adr_i[12]
port 536 nsew default input
rlabel metal2 s 58778 -960 58890 480 8 wbs_adr_i[13]
port 537 nsew default input
rlabel metal2 s 62366 -960 62478 480 8 wbs_adr_i[14]
port 538 nsew default input
rlabel metal2 s 65954 -960 66066 480 8 wbs_adr_i[15]
port 539 nsew default input
rlabel metal2 s 69450 -960 69562 480 8 wbs_adr_i[16]
port 540 nsew default input
rlabel metal2 s 73038 -960 73150 480 8 wbs_adr_i[17]
port 541 nsew default input
rlabel metal2 s 76626 -960 76738 480 8 wbs_adr_i[18]
port 542 nsew default input
rlabel metal2 s 80214 -960 80326 480 8 wbs_adr_i[19]
port 543 nsew default input
rlabel metal2 s 12410 -960 12522 480 8 wbs_adr_i[1]
port 544 nsew default input
rlabel metal2 s 83802 -960 83914 480 8 wbs_adr_i[20]
port 545 nsew default input
rlabel metal2 s 87298 -960 87410 480 8 wbs_adr_i[21]
port 546 nsew default input
rlabel metal2 s 90886 -960 90998 480 8 wbs_adr_i[22]
port 547 nsew default input
rlabel metal2 s 94474 -960 94586 480 8 wbs_adr_i[23]
port 548 nsew default input
rlabel metal2 s 98062 -960 98174 480 8 wbs_adr_i[24]
port 549 nsew default input
rlabel metal2 s 101558 -960 101670 480 8 wbs_adr_i[25]
port 550 nsew default input
rlabel metal2 s 105146 -960 105258 480 8 wbs_adr_i[26]
port 551 nsew default input
rlabel metal2 s 108734 -960 108846 480 8 wbs_adr_i[27]
port 552 nsew default input
rlabel metal2 s 112322 -960 112434 480 8 wbs_adr_i[28]
port 553 nsew default input
rlabel metal2 s 115910 -960 116022 480 8 wbs_adr_i[29]
port 554 nsew default input
rlabel metal2 s 17194 -960 17306 480 8 wbs_adr_i[2]
port 555 nsew default input
rlabel metal2 s 119406 -960 119518 480 8 wbs_adr_i[30]
port 556 nsew default input
rlabel metal2 s 122994 -960 123106 480 8 wbs_adr_i[31]
port 557 nsew default input
rlabel metal2 s 21886 -960 21998 480 8 wbs_adr_i[3]
port 558 nsew default input
rlabel metal2 s 26670 -960 26782 480 8 wbs_adr_i[4]
port 559 nsew default input
rlabel metal2 s 30258 -960 30370 480 8 wbs_adr_i[5]
port 560 nsew default input
rlabel metal2 s 33846 -960 33958 480 8 wbs_adr_i[6]
port 561 nsew default input
rlabel metal2 s 37342 -960 37454 480 8 wbs_adr_i[7]
port 562 nsew default input
rlabel metal2 s 40930 -960 41042 480 8 wbs_adr_i[8]
port 563 nsew default input
rlabel metal2 s 44518 -960 44630 480 8 wbs_adr_i[9]
port 564 nsew default input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 565 nsew default input
rlabel metal2 s 8822 -960 8934 480 8 wbs_dat_i[0]
port 566 nsew default input
rlabel metal2 s 49302 -960 49414 480 8 wbs_dat_i[10]
port 567 nsew default input
rlabel metal2 s 52798 -960 52910 480 8 wbs_dat_i[11]
port 568 nsew default input
rlabel metal2 s 56386 -960 56498 480 8 wbs_dat_i[12]
port 569 nsew default input
rlabel metal2 s 59974 -960 60086 480 8 wbs_dat_i[13]
port 570 nsew default input
rlabel metal2 s 63562 -960 63674 480 8 wbs_dat_i[14]
port 571 nsew default input
rlabel metal2 s 67150 -960 67262 480 8 wbs_dat_i[15]
port 572 nsew default input
rlabel metal2 s 70646 -960 70758 480 8 wbs_dat_i[16]
port 573 nsew default input
rlabel metal2 s 74234 -960 74346 480 8 wbs_dat_i[17]
port 574 nsew default input
rlabel metal2 s 77822 -960 77934 480 8 wbs_dat_i[18]
port 575 nsew default input
rlabel metal2 s 81410 -960 81522 480 8 wbs_dat_i[19]
port 576 nsew default input
rlabel metal2 s 13606 -960 13718 480 8 wbs_dat_i[1]
port 577 nsew default input
rlabel metal2 s 84906 -960 85018 480 8 wbs_dat_i[20]
port 578 nsew default input
rlabel metal2 s 88494 -960 88606 480 8 wbs_dat_i[21]
port 579 nsew default input
rlabel metal2 s 92082 -960 92194 480 8 wbs_dat_i[22]
port 580 nsew default input
rlabel metal2 s 95670 -960 95782 480 8 wbs_dat_i[23]
port 581 nsew default input
rlabel metal2 s 99258 -960 99370 480 8 wbs_dat_i[24]
port 582 nsew default input
rlabel metal2 s 102754 -960 102866 480 8 wbs_dat_i[25]
port 583 nsew default input
rlabel metal2 s 106342 -960 106454 480 8 wbs_dat_i[26]
port 584 nsew default input
rlabel metal2 s 109930 -960 110042 480 8 wbs_dat_i[27]
port 585 nsew default input
rlabel metal2 s 113518 -960 113630 480 8 wbs_dat_i[28]
port 586 nsew default input
rlabel metal2 s 117106 -960 117218 480 8 wbs_dat_i[29]
port 587 nsew default input
rlabel metal2 s 18298 -960 18410 480 8 wbs_dat_i[2]
port 588 nsew default input
rlabel metal2 s 120602 -960 120714 480 8 wbs_dat_i[30]
port 589 nsew default input
rlabel metal2 s 124190 -960 124302 480 8 wbs_dat_i[31]
port 590 nsew default input
rlabel metal2 s 23082 -960 23194 480 8 wbs_dat_i[3]
port 591 nsew default input
rlabel metal2 s 27866 -960 27978 480 8 wbs_dat_i[4]
port 592 nsew default input
rlabel metal2 s 31454 -960 31566 480 8 wbs_dat_i[5]
port 593 nsew default input
rlabel metal2 s 34950 -960 35062 480 8 wbs_dat_i[6]
port 594 nsew default input
rlabel metal2 s 38538 -960 38650 480 8 wbs_dat_i[7]
port 595 nsew default input
rlabel metal2 s 42126 -960 42238 480 8 wbs_dat_i[8]
port 596 nsew default input
rlabel metal2 s 45714 -960 45826 480 8 wbs_dat_i[9]
port 597 nsew default input
rlabel metal2 s 10018 -960 10130 480 8 wbs_dat_o[0]
port 598 nsew default tristate
rlabel metal2 s 50498 -960 50610 480 8 wbs_dat_o[10]
port 599 nsew default tristate
rlabel metal2 s 53994 -960 54106 480 8 wbs_dat_o[11]
port 600 nsew default tristate
rlabel metal2 s 57582 -960 57694 480 8 wbs_dat_o[12]
port 601 nsew default tristate
rlabel metal2 s 61170 -960 61282 480 8 wbs_dat_o[13]
port 602 nsew default tristate
rlabel metal2 s 64758 -960 64870 480 8 wbs_dat_o[14]
port 603 nsew default tristate
rlabel metal2 s 68254 -960 68366 480 8 wbs_dat_o[15]
port 604 nsew default tristate
rlabel metal2 s 71842 -960 71954 480 8 wbs_dat_o[16]
port 605 nsew default tristate
rlabel metal2 s 75430 -960 75542 480 8 wbs_dat_o[17]
port 606 nsew default tristate
rlabel metal2 s 79018 -960 79130 480 8 wbs_dat_o[18]
port 607 nsew default tristate
rlabel metal2 s 82606 -960 82718 480 8 wbs_dat_o[19]
port 608 nsew default tristate
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[1]
port 609 nsew default tristate
rlabel metal2 s 86102 -960 86214 480 8 wbs_dat_o[20]
port 610 nsew default tristate
rlabel metal2 s 89690 -960 89802 480 8 wbs_dat_o[21]
port 611 nsew default tristate
rlabel metal2 s 93278 -960 93390 480 8 wbs_dat_o[22]
port 612 nsew default tristate
rlabel metal2 s 96866 -960 96978 480 8 wbs_dat_o[23]
port 613 nsew default tristate
rlabel metal2 s 100454 -960 100566 480 8 wbs_dat_o[24]
port 614 nsew default tristate
rlabel metal2 s 103950 -960 104062 480 8 wbs_dat_o[25]
port 615 nsew default tristate
rlabel metal2 s 107538 -960 107650 480 8 wbs_dat_o[26]
port 616 nsew default tristate
rlabel metal2 s 111126 -960 111238 480 8 wbs_dat_o[27]
port 617 nsew default tristate
rlabel metal2 s 114714 -960 114826 480 8 wbs_dat_o[28]
port 618 nsew default tristate
rlabel metal2 s 118210 -960 118322 480 8 wbs_dat_o[29]
port 619 nsew default tristate
rlabel metal2 s 19494 -960 19606 480 8 wbs_dat_o[2]
port 620 nsew default tristate
rlabel metal2 s 121798 -960 121910 480 8 wbs_dat_o[30]
port 621 nsew default tristate
rlabel metal2 s 125386 -960 125498 480 8 wbs_dat_o[31]
port 622 nsew default tristate
rlabel metal2 s 24278 -960 24390 480 8 wbs_dat_o[3]
port 623 nsew default tristate
rlabel metal2 s 29062 -960 29174 480 8 wbs_dat_o[4]
port 624 nsew default tristate
rlabel metal2 s 32650 -960 32762 480 8 wbs_dat_o[5]
port 625 nsew default tristate
rlabel metal2 s 36146 -960 36258 480 8 wbs_dat_o[6]
port 626 nsew default tristate
rlabel metal2 s 39734 -960 39846 480 8 wbs_dat_o[7]
port 627 nsew default tristate
rlabel metal2 s 43322 -960 43434 480 8 wbs_dat_o[8]
port 628 nsew default tristate
rlabel metal2 s 46910 -960 47022 480 8 wbs_dat_o[9]
port 629 nsew default tristate
rlabel metal2 s 11214 -960 11326 480 8 wbs_sel_i[0]
port 630 nsew default input
rlabel metal2 s 15998 -960 16110 480 8 wbs_sel_i[1]
port 631 nsew default input
rlabel metal2 s 20690 -960 20802 480 8 wbs_sel_i[2]
port 632 nsew default input
rlabel metal2 s 25474 -960 25586 480 8 wbs_sel_i[3]
port 633 nsew default input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 634 nsew default input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 635 nsew default input
rlabel metal5 s -1996 -924 585920 -324 8 vccd1
port 636 nsew default input
rlabel metal5 s -2936 -1864 586860 -1264 8 vssd1
port 637 nsew default input
rlabel metal5 s -3876 -2804 587800 -2204 8 vccd2
port 638 nsew default input
rlabel metal5 s -4816 -3744 588740 -3144 8 vssd2
port 639 nsew default input
rlabel metal5 s -5756 -4684 589680 -4084 8 vdda1
port 640 nsew default input
rlabel metal5 s -6696 -5624 590620 -5024 8 vssa1
port 641 nsew default input
rlabel metal5 s -7636 -6564 591560 -5964 8 vdda2
port 642 nsew default input
rlabel metal5 s -8576 -7504 592500 -6904 8 vssa2
port 643 nsew default input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
