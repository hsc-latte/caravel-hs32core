magic
tech sky130A
magscale 1 2
timestamp 1612306080
<< metal1 >>
rect 478506 700884 478512 700936
rect 478564 700924 478570 700936
rect 539594 700924 539600 700936
rect 478564 700896 539600 700924
rect 478564 700884 478570 700896
rect 539594 700884 539600 700896
rect 539652 700884 539658 700936
rect 413646 700816 413652 700868
rect 413704 700856 413710 700868
rect 539686 700856 539692 700868
rect 413704 700828 539692 700856
rect 413704 700816 413710 700828
rect 539686 700816 539692 700828
rect 539744 700816 539750 700868
rect 348786 700748 348792 700800
rect 348844 700788 348850 700800
rect 539778 700788 539784 700800
rect 348844 700760 539784 700788
rect 348844 700748 348850 700760
rect 539778 700748 539784 700760
rect 539836 700748 539842 700800
rect 332502 700680 332508 700732
rect 332560 700720 332566 700732
rect 539134 700720 539140 700732
rect 332560 700692 539140 700720
rect 332560 700680 332566 700692
rect 539134 700680 539140 700692
rect 539192 700680 539198 700732
rect 235166 700612 235172 700664
rect 235224 700652 235230 700664
rect 235902 700652 235908 700664
rect 235224 700624 235908 700652
rect 235224 700612 235230 700624
rect 235902 700612 235908 700624
rect 235960 700612 235966 700664
rect 283834 700612 283840 700664
rect 283892 700652 283898 700664
rect 539226 700652 539232 700664
rect 283892 700624 539232 700652
rect 283892 700612 283898 700624
rect 539226 700612 539232 700624
rect 539284 700612 539290 700664
rect 218974 700544 218980 700596
rect 219032 700584 219038 700596
rect 539962 700584 539968 700596
rect 219032 700556 539968 700584
rect 219032 700544 219038 700556
rect 539962 700544 539968 700556
rect 540020 700544 540026 700596
rect 202782 700476 202788 700528
rect 202840 700516 202846 700528
rect 539870 700516 539876 700528
rect 202840 700488 539876 700516
rect 202840 700476 202846 700488
rect 539870 700476 539876 700488
rect 539928 700476 539934 700528
rect 154114 700408 154120 700460
rect 154172 700448 154178 700460
rect 540054 700448 540060 700460
rect 154172 700420 540060 700448
rect 154172 700408 154178 700420
rect 540054 700408 540060 700420
rect 540112 700408 540118 700460
rect 72970 700340 72976 700392
rect 73028 700380 73034 700392
rect 540146 700380 540152 700392
rect 73028 700352 540152 700380
rect 73028 700340 73034 700352
rect 540146 700340 540152 700352
rect 540204 700340 540210 700392
rect 40494 700272 40500 700324
rect 40552 700312 40558 700324
rect 541066 700312 541072 700324
rect 40552 700284 541072 700312
rect 40552 700272 40558 700284
rect 541066 700272 541072 700284
rect 541124 700272 541130 700324
rect 549898 700272 549904 700324
rect 549956 700312 549962 700324
rect 559650 700312 559656 700324
rect 549956 700284 559656 700312
rect 549956 700272 549962 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 397454 699932 397460 699984
rect 397512 699972 397518 699984
rect 398742 699972 398748 699984
rect 397512 699944 398748 699972
rect 397512 699932 397518 699944
rect 398742 699932 398748 699944
rect 398800 699932 398806 699984
rect 494790 699796 494796 699848
rect 494848 699836 494854 699848
rect 495342 699836 495348 699848
rect 494848 699808 495348 699836
rect 494848 699796 494854 699808
rect 495342 699796 495348 699808
rect 495400 699796 495406 699848
rect 105446 699660 105452 699712
rect 105504 699700 105510 699712
rect 106182 699700 106188 699712
rect 105504 699672 106188 699700
rect 105504 699660 105510 699672
rect 106182 699660 106188 699672
rect 106240 699660 106246 699712
rect 170306 699660 170312 699712
rect 170364 699700 170370 699712
rect 171042 699700 171048 699712
rect 170364 699672 171048 699700
rect 170364 699660 170370 699672
rect 171042 699660 171048 699672
rect 171100 699660 171106 699712
rect 300118 699660 300124 699712
rect 300176 699700 300182 699712
rect 300762 699700 300768 699712
rect 300176 699672 300768 699700
rect 300176 699660 300182 699672
rect 300762 699660 300768 699672
rect 300820 699660 300826 699712
rect 364978 699660 364984 699712
rect 365036 699700 365042 699712
rect 365622 699700 365628 699712
rect 365036 699672 365628 699700
rect 365036 699660 365042 699672
rect 365622 699660 365628 699672
rect 365680 699660 365686 699712
rect 429838 699660 429844 699712
rect 429896 699700 429902 699712
rect 430482 699700 430488 699712
rect 429896 699672 430488 699700
rect 429896 699660 429902 699672
rect 430482 699660 430488 699672
rect 430540 699660 430546 699712
rect 462314 699660 462320 699712
rect 462372 699700 462378 699712
rect 463602 699700 463608 699712
rect 462372 699672 463608 699700
rect 462372 699660 462378 699672
rect 463602 699660 463608 699672
rect 463660 699660 463666 699712
rect 527174 699660 527180 699712
rect 527232 699700 527238 699712
rect 528462 699700 528468 699712
rect 527232 699672 528468 699700
rect 527232 699660 527238 699672
rect 528462 699660 528468 699672
rect 528520 699660 528526 699712
rect 563698 696940 563704 696992
rect 563756 696980 563762 696992
rect 580166 696980 580172 696992
rect 563756 696952 580172 696980
rect 563756 696940 563762 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 554038 685856 554044 685908
rect 554096 685896 554102 685908
rect 580166 685896 580172 685908
rect 554096 685868 580172 685896
rect 554096 685856 554102 685868
rect 580166 685856 580172 685868
rect 580224 685856 580230 685908
rect 3510 681708 3516 681760
rect 3568 681748 3574 681760
rect 541158 681748 541164 681760
rect 3568 681720 541164 681748
rect 3568 681708 3574 681720
rect 541158 681708 541164 681720
rect 541216 681708 541222 681760
rect 543274 676132 543280 676184
rect 543332 676172 543338 676184
rect 543550 676172 543556 676184
rect 543332 676144 543556 676172
rect 543332 676132 543338 676144
rect 543550 676132 543556 676144
rect 543608 676132 543614 676184
rect 547138 673480 547144 673532
rect 547196 673520 547202 673532
rect 580166 673520 580172 673532
rect 547196 673492 580172 673520
rect 547196 673480 547202 673492
rect 580166 673480 580172 673492
rect 580224 673480 580230 673532
rect 3418 667904 3424 667956
rect 3476 667944 3482 667956
rect 541250 667944 541256 667956
rect 3476 667916 541256 667944
rect 3476 667904 3482 667916
rect 541250 667904 541256 667916
rect 541308 667904 541314 667956
rect 3050 652740 3056 652792
rect 3108 652780 3114 652792
rect 540238 652780 540244 652792
rect 3108 652752 540244 652780
rect 3108 652740 3114 652752
rect 540238 652740 540244 652752
rect 540296 652740 540302 652792
rect 560938 650020 560944 650072
rect 560996 650060 561002 650072
rect 580166 650060 580172 650072
rect 560996 650032 580172 650060
rect 560996 650020 561002 650032
rect 580166 650020 580172 650032
rect 580224 650020 580230 650072
rect 543458 647232 543464 647284
rect 543516 647272 543522 647284
rect 543550 647272 543556 647284
rect 543516 647244 543556 647272
rect 543516 647232 543522 647244
rect 543550 647232 543556 647244
rect 543608 647232 543614 647284
rect 543458 640364 543464 640416
rect 543516 640404 543522 640416
rect 543550 640404 543556 640416
rect 543516 640376 543556 640404
rect 543516 640364 543522 640376
rect 543550 640364 543556 640376
rect 543608 640364 543614 640416
rect 565078 638936 565084 638988
rect 565136 638976 565142 638988
rect 580166 638976 580172 638988
rect 565136 638948 580172 638976
rect 565136 638936 565142 638948
rect 580166 638936 580172 638948
rect 580224 638936 580230 638988
rect 543366 630640 543372 630692
rect 543424 630680 543430 630692
rect 543550 630680 543556 630692
rect 543424 630652 543556 630680
rect 543424 630640 543430 630652
rect 543550 630640 543556 630652
rect 543608 630640 543614 630692
rect 545758 626560 545764 626612
rect 545816 626600 545822 626612
rect 580166 626600 580172 626612
rect 545816 626572 580172 626600
rect 545816 626560 545822 626572
rect 580166 626560 580172 626572
rect 580224 626560 580230 626612
rect 267642 620236 267648 620288
rect 267700 620276 267706 620288
rect 540330 620276 540336 620288
rect 267700 620248 540336 620276
rect 267700 620236 267706 620248
rect 540330 620236 540336 620248
rect 540388 620236 540394 620288
rect 488534 613368 488540 613420
rect 488592 613408 488598 613420
rect 493962 613408 493968 613420
rect 488592 613380 493968 613408
rect 488592 613368 488598 613380
rect 493962 613368 493968 613380
rect 494020 613368 494026 613420
rect 373626 612756 373632 612808
rect 373684 612796 373690 612808
rect 379606 612796 379612 612808
rect 373684 612768 379612 612796
rect 373684 612756 373690 612768
rect 379606 612756 379612 612768
rect 379664 612796 379670 612808
rect 488534 612796 488540 612808
rect 379664 612768 488540 612796
rect 379664 612756 379670 612768
rect 488534 612756 488540 612768
rect 488592 612756 488598 612808
rect 493962 612756 493968 612808
rect 494020 612796 494026 612808
rect 499574 612796 499580 612808
rect 494020 612768 499580 612796
rect 494020 612756 494026 612768
rect 499574 612756 499580 612768
rect 499632 612756 499638 612808
rect 543366 611328 543372 611380
rect 543424 611368 543430 611380
rect 543550 611368 543556 611380
rect 543424 611340 543556 611368
rect 543424 611328 543430 611340
rect 543550 611328 543556 611340
rect 543608 611328 543614 611380
rect 495342 610784 495348 610836
rect 495400 610824 495406 610836
rect 541342 610824 541348 610836
rect 495400 610796 541348 610824
rect 495400 610784 495406 610796
rect 541342 610784 541348 610796
rect 541400 610784 541406 610836
rect 463602 610716 463608 610768
rect 463660 610756 463666 610768
rect 539318 610756 539324 610768
rect 463660 610728 539324 610756
rect 463660 610716 463666 610728
rect 539318 610716 539324 610728
rect 539376 610716 539382 610768
rect 430482 610648 430488 610700
rect 430540 610688 430546 610700
rect 541434 610688 541440 610700
rect 430540 610660 541440 610688
rect 430540 610648 430546 610660
rect 541434 610648 541440 610660
rect 541492 610648 541498 610700
rect 365622 610580 365628 610632
rect 365680 610620 365686 610632
rect 541526 610620 541532 610632
rect 365680 610592 541532 610620
rect 365680 610580 365686 610592
rect 541526 610580 541532 610592
rect 541584 610580 541590 610632
rect 379974 610376 379980 610428
rect 380032 610416 380038 610428
rect 496446 610416 496452 610428
rect 380032 610388 496452 610416
rect 380032 610376 380038 610388
rect 496446 610376 496452 610388
rect 496504 610376 496510 610428
rect 3418 610308 3424 610360
rect 3476 610348 3482 610360
rect 541710 610348 541716 610360
rect 3476 610320 541716 610348
rect 3476 610308 3482 610320
rect 541710 610308 541716 610320
rect 541768 610308 541774 610360
rect 387702 605820 387708 605872
rect 387760 605860 387766 605872
rect 416774 605860 416780 605872
rect 387760 605832 416780 605860
rect 387760 605820 387766 605832
rect 416774 605820 416780 605832
rect 416832 605820 416838 605872
rect 384942 604460 384948 604512
rect 385000 604500 385006 604512
rect 416774 604500 416780 604512
rect 385000 604472 416780 604500
rect 385000 604460 385006 604472
rect 416774 604460 416780 604472
rect 416832 604460 416838 604512
rect 382182 603100 382188 603152
rect 382240 603140 382246 603152
rect 416774 603140 416780 603152
rect 382240 603112 416780 603140
rect 382240 603100 382246 603112
rect 416774 603100 416780 603112
rect 416832 603100 416838 603152
rect 558178 603100 558184 603152
rect 558236 603140 558242 603152
rect 580166 603140 580172 603152
rect 558236 603112 580172 603140
rect 558236 603100 558242 603112
rect 580166 603100 580172 603112
rect 580224 603100 580230 603152
rect 379422 601672 379428 601724
rect 379480 601712 379486 601724
rect 416774 601712 416780 601724
rect 379480 601684 416780 601712
rect 379480 601672 379486 601684
rect 416774 601672 416780 601684
rect 416832 601672 416838 601724
rect 378042 600312 378048 600364
rect 378100 600352 378106 600364
rect 416774 600352 416780 600364
rect 378100 600324 416780 600352
rect 378100 600312 378106 600324
rect 416774 600312 416780 600324
rect 416832 600312 416838 600364
rect 543366 592016 543372 592068
rect 543424 592056 543430 592068
rect 543550 592056 543556 592068
rect 543424 592028 543556 592056
rect 543424 592016 543430 592028
rect 543550 592016 543556 592028
rect 543608 592016 543614 592068
rect 574738 592016 574744 592068
rect 574796 592056 574802 592068
rect 580166 592056 580172 592068
rect 574796 592028 580172 592056
rect 574796 592016 574802 592028
rect 580166 592016 580172 592028
rect 580224 592016 580230 592068
rect 544378 579640 544384 579692
rect 544436 579680 544442 579692
rect 580166 579680 580172 579692
rect 544436 579652 580172 579680
rect 544436 579640 544442 579652
rect 580166 579640 580172 579652
rect 580224 579640 580230 579692
rect 543366 572704 543372 572756
rect 543424 572744 543430 572756
rect 543550 572744 543556 572756
rect 543424 572716 543556 572744
rect 543424 572704 543430 572716
rect 543550 572704 543556 572716
rect 543608 572704 543614 572756
rect 556798 556180 556804 556232
rect 556856 556220 556862 556232
rect 580166 556220 580172 556232
rect 556856 556192 580172 556220
rect 556856 556180 556862 556192
rect 580166 556180 580172 556192
rect 580224 556180 580230 556232
rect 543366 553392 543372 553444
rect 543424 553432 543430 553444
rect 543550 553432 543556 553444
rect 543424 553404 543556 553432
rect 543424 553392 543430 553404
rect 543550 553392 543556 553404
rect 543608 553392 543614 553444
rect 573358 545096 573364 545148
rect 573416 545136 573422 545148
rect 580166 545136 580172 545148
rect 573416 545108 580172 545136
rect 573416 545096 573422 545108
rect 580166 545096 580172 545108
rect 580224 545096 580230 545148
rect 413922 539588 413928 539640
rect 413980 539628 413986 539640
rect 416958 539628 416964 539640
rect 413980 539600 416964 539628
rect 413980 539588 413986 539600
rect 416958 539588 416964 539600
rect 417016 539588 417022 539640
rect 379514 538228 379520 538280
rect 379572 538268 379578 538280
rect 379790 538268 379796 538280
rect 379572 538240 379796 538268
rect 379572 538228 379578 538240
rect 379790 538228 379796 538240
rect 379848 538228 379854 538280
rect 410518 538228 410524 538280
rect 410576 538268 410582 538280
rect 416774 538268 416780 538280
rect 410576 538240 416780 538268
rect 410576 538228 410582 538240
rect 416774 538228 416780 538240
rect 416832 538228 416838 538280
rect 379514 536052 379520 536104
rect 379572 536092 379578 536104
rect 379790 536092 379796 536104
rect 379572 536064 379796 536092
rect 379572 536052 379578 536064
rect 379790 536052 379796 536064
rect 379848 536052 379854 536104
rect 543366 534080 543372 534132
rect 543424 534120 543430 534132
rect 543550 534120 543556 534132
rect 543424 534092 543556 534120
rect 543424 534080 543430 534092
rect 543550 534080 543556 534092
rect 543608 534080 543614 534132
rect 544470 532720 544476 532772
rect 544528 532760 544534 532772
rect 580166 532760 580172 532772
rect 544528 532732 580172 532760
rect 544528 532720 544534 532732
rect 580166 532720 580172 532732
rect 580224 532720 580230 532772
rect 409874 521568 409880 521620
rect 409932 521608 409938 521620
rect 410518 521608 410524 521620
rect 409932 521580 410524 521608
rect 409932 521568 409938 521580
rect 410518 521568 410524 521580
rect 410576 521568 410582 521620
rect 297266 520888 297272 520940
rect 297324 520928 297330 520940
rect 409874 520928 409880 520940
rect 297324 520900 409880 520928
rect 297324 520888 297330 520900
rect 409874 520888 409880 520900
rect 409932 520888 409938 520940
rect 379606 518916 379612 518968
rect 379664 518956 379670 518968
rect 379790 518956 379796 518968
rect 379664 518928 379796 518956
rect 379664 518916 379670 518928
rect 379790 518916 379796 518928
rect 379848 518916 379854 518968
rect 320082 518848 320088 518900
rect 320140 518888 320146 518900
rect 328914 518888 328920 518900
rect 320140 518860 328920 518888
rect 320140 518848 320146 518860
rect 328914 518848 328920 518860
rect 328972 518888 328978 518900
rect 329650 518888 329656 518900
rect 328972 518860 329656 518888
rect 328972 518848 328978 518860
rect 329650 518848 329656 518860
rect 329708 518848 329714 518900
rect 348970 518848 348976 518900
rect 349028 518888 349034 518900
rect 455414 518888 455420 518900
rect 349028 518860 455420 518888
rect 349028 518848 349034 518860
rect 455414 518848 455420 518860
rect 455472 518848 455478 518900
rect 289722 518780 289728 518832
rect 289780 518820 289786 518832
rect 322934 518820 322940 518832
rect 289780 518792 322940 518820
rect 289780 518780 289786 518792
rect 322934 518780 322940 518792
rect 322992 518780 322998 518832
rect 327350 518780 327356 518832
rect 327408 518820 327414 518832
rect 336918 518820 336924 518832
rect 327408 518792 336924 518820
rect 327408 518780 327414 518792
rect 336918 518780 336924 518792
rect 336976 518780 336982 518832
rect 345290 518780 345296 518832
rect 345348 518820 345354 518832
rect 448514 518820 448520 518832
rect 345348 518792 448520 518820
rect 345348 518780 345354 518792
rect 448514 518780 448520 518792
rect 448572 518780 448578 518832
rect 448698 518780 448704 518832
rect 448756 518820 448762 518832
rect 458358 518820 458364 518832
rect 448756 518792 458364 518820
rect 448756 518780 448762 518792
rect 458358 518780 458364 518792
rect 458416 518780 458422 518832
rect 307662 518712 307668 518764
rect 307720 518752 307726 518764
rect 331306 518752 331312 518764
rect 307720 518724 331312 518752
rect 307720 518712 307726 518724
rect 331306 518712 331312 518724
rect 331364 518712 331370 518764
rect 331398 518712 331404 518764
rect 331456 518752 331462 518764
rect 340598 518752 340604 518764
rect 331456 518724 340604 518752
rect 331456 518712 331462 518724
rect 340598 518712 340604 518724
rect 340656 518712 340662 518764
rect 346578 518712 346584 518764
rect 346636 518752 346642 518764
rect 449894 518752 449900 518764
rect 346636 518724 449900 518752
rect 346636 518712 346642 518724
rect 449894 518712 449900 518724
rect 449952 518712 449958 518764
rect 451274 518712 451280 518764
rect 451332 518752 451338 518764
rect 459554 518752 459560 518764
rect 451332 518724 459560 518752
rect 451332 518712 451338 518724
rect 459554 518712 459560 518724
rect 459612 518712 459618 518764
rect 314562 518644 314568 518696
rect 314620 518684 314626 518696
rect 323118 518684 323124 518696
rect 314620 518656 323124 518684
rect 314620 518644 314626 518656
rect 323118 518644 323124 518656
rect 323176 518684 323182 518696
rect 332410 518684 332416 518696
rect 323176 518656 332416 518684
rect 323176 518644 323182 518656
rect 332410 518644 332416 518656
rect 332468 518684 332474 518696
rect 341518 518684 341524 518696
rect 332468 518656 341524 518684
rect 332468 518644 332474 518656
rect 341518 518644 341524 518656
rect 341576 518644 341582 518696
rect 443178 518644 443184 518696
rect 443236 518684 443242 518696
rect 452562 518684 452568 518696
rect 443236 518656 452568 518684
rect 443236 518644 443242 518656
rect 452562 518644 452568 518656
rect 452620 518684 452626 518696
rect 452620 518656 452792 518684
rect 452620 518644 452626 518656
rect 318702 518576 318708 518628
rect 318760 518616 318766 518628
rect 327350 518616 327356 518628
rect 318760 518588 327356 518616
rect 318760 518576 318766 518588
rect 327350 518576 327356 518588
rect 327408 518576 327414 518628
rect 329650 518576 329656 518628
rect 329708 518616 329714 518628
rect 338114 518616 338120 518628
rect 329708 518588 338120 518616
rect 329708 518576 329714 518588
rect 338114 518576 338120 518588
rect 338172 518616 338178 518628
rect 347682 518616 347688 518628
rect 338172 518588 347688 518616
rect 338172 518576 338178 518588
rect 347682 518576 347688 518588
rect 347740 518616 347746 518628
rect 452654 518616 452660 518628
rect 347740 518588 452660 518616
rect 347740 518576 347746 518588
rect 452654 518576 452660 518588
rect 452712 518576 452718 518628
rect 321094 518508 321100 518560
rect 321152 518548 321158 518560
rect 330110 518548 330116 518560
rect 321152 518520 330116 518548
rect 321152 518508 321158 518520
rect 330110 518508 330116 518520
rect 330168 518548 330174 518560
rect 339494 518548 339500 518560
rect 330168 518520 339500 518548
rect 330168 518508 330174 518520
rect 339494 518508 339500 518520
rect 339552 518548 339558 518560
rect 348970 518548 348976 518560
rect 339552 518520 348976 518548
rect 339552 518508 339558 518520
rect 348970 518508 348976 518520
rect 349028 518508 349034 518560
rect 442534 518508 442540 518560
rect 442592 518548 442598 518560
rect 451274 518548 451280 518560
rect 442592 518520 451280 518548
rect 442592 518508 442598 518520
rect 451274 518508 451280 518520
rect 451332 518508 451338 518560
rect 452764 518548 452792 518656
rect 457070 518644 457076 518696
rect 457128 518684 457134 518696
rect 466454 518684 466460 518696
rect 457128 518656 466460 518684
rect 457128 518644 457134 518656
rect 466454 518644 466460 518656
rect 466512 518644 466518 518696
rect 461026 518548 461032 518560
rect 452764 518520 461032 518548
rect 461026 518508 461032 518520
rect 461084 518508 461090 518560
rect 274542 518440 274548 518492
rect 274600 518480 274606 518492
rect 316034 518480 316040 518492
rect 274600 518452 316040 518480
rect 274600 518440 274606 518452
rect 316034 518440 316040 518452
rect 316092 518440 316098 518492
rect 317322 518440 317328 518492
rect 317380 518480 317386 518492
rect 326430 518480 326436 518492
rect 317380 518452 326436 518480
rect 317380 518440 317386 518452
rect 326430 518440 326436 518452
rect 326488 518480 326494 518492
rect 335814 518480 335820 518492
rect 326488 518452 335820 518480
rect 326488 518440 326494 518452
rect 335814 518440 335820 518452
rect 335872 518480 335878 518492
rect 345290 518480 345296 518492
rect 335872 518452 345296 518480
rect 335872 518440 335878 518452
rect 345290 518440 345296 518452
rect 345348 518440 345354 518492
rect 447962 518440 447968 518492
rect 448020 518480 448026 518492
rect 457070 518480 457076 518492
rect 448020 518452 457076 518480
rect 448020 518440 448026 518452
rect 457070 518440 457076 518452
rect 457128 518440 457134 518492
rect 458358 518440 458364 518492
rect 458416 518480 458422 518492
rect 466454 518480 466460 518492
rect 458416 518452 466460 518480
rect 458416 518440 458422 518452
rect 466454 518440 466460 518452
rect 466512 518440 466518 518492
rect 313182 518372 313188 518424
rect 313240 518412 313246 518424
rect 313240 518384 317092 518412
rect 313240 518372 313246 518384
rect 271782 518304 271788 518356
rect 271840 518344 271846 518356
rect 314654 518344 314660 518356
rect 271840 518316 314660 518344
rect 271840 518304 271846 518316
rect 314654 518304 314660 518316
rect 314712 518304 314718 518356
rect 317064 518344 317092 518384
rect 317230 518372 317236 518424
rect 317288 518412 317294 518424
rect 325418 518412 325424 518424
rect 317288 518384 325424 518412
rect 317288 518372 317294 518384
rect 325418 518372 325424 518384
rect 325476 518372 325482 518424
rect 325510 518372 325516 518424
rect 325568 518412 325574 518424
rect 331398 518412 331404 518424
rect 325568 518384 331404 518412
rect 325568 518372 325574 518384
rect 331398 518372 331404 518384
rect 331456 518372 331462 518424
rect 333790 518372 333796 518424
rect 333848 518412 333854 518424
rect 342990 518412 342996 518424
rect 333848 518384 342996 518412
rect 333848 518372 333854 518384
rect 342990 518372 342996 518384
rect 343048 518372 343054 518424
rect 369762 518372 369768 518424
rect 369820 518412 369826 518424
rect 426434 518412 426440 518424
rect 369820 518384 426440 518412
rect 369820 518372 369826 518384
rect 426434 518372 426440 518384
rect 426492 518372 426498 518424
rect 444282 518372 444288 518424
rect 444340 518412 444346 518424
rect 453758 518412 453764 518424
rect 444340 518384 453764 518412
rect 444340 518372 444346 518384
rect 453758 518372 453764 518384
rect 453816 518412 453822 518424
rect 462314 518412 462320 518424
rect 453816 518384 462320 518412
rect 453816 518372 453822 518384
rect 462314 518372 462320 518384
rect 462372 518372 462378 518424
rect 318794 518344 318800 518356
rect 317064 518316 318800 518344
rect 318794 518304 318800 518316
rect 318852 518304 318858 518356
rect 336918 518304 336924 518356
rect 336976 518344 336982 518356
rect 346578 518344 346584 518356
rect 336976 518316 346584 518344
rect 336976 518304 336982 518316
rect 346578 518304 346584 518316
rect 346636 518304 346642 518356
rect 357342 518304 357348 518356
rect 357400 518344 357406 518356
rect 430574 518344 430580 518356
rect 357400 518316 430580 518344
rect 357400 518304 357406 518316
rect 430574 518304 430580 518316
rect 430632 518304 430638 518356
rect 435910 518304 435916 518356
rect 435968 518344 435974 518356
rect 444300 518344 444328 518372
rect 435968 518316 444328 518344
rect 435968 518304 435974 518316
rect 445386 518304 445392 518356
rect 445444 518344 445450 518356
rect 455322 518344 455328 518356
rect 445444 518316 455328 518344
rect 445444 518304 445450 518316
rect 455322 518304 455328 518316
rect 455380 518344 455386 518356
rect 463694 518344 463700 518356
rect 455380 518316 463700 518344
rect 455380 518304 455386 518316
rect 463694 518304 463700 518316
rect 463752 518304 463758 518356
rect 269022 518236 269028 518288
rect 269080 518276 269086 518288
rect 313274 518276 313280 518288
rect 269080 518248 313280 518276
rect 269080 518236 269086 518248
rect 313274 518236 313280 518248
rect 313332 518236 313338 518288
rect 315850 518236 315856 518288
rect 315908 518276 315914 518288
rect 320174 518276 320180 518288
rect 315908 518248 320180 518276
rect 315908 518236 315914 518248
rect 320174 518236 320180 518248
rect 320232 518236 320238 518288
rect 325418 518236 325424 518288
rect 325476 518276 325482 518288
rect 334710 518276 334716 518288
rect 325476 518248 334716 518276
rect 325476 518236 325482 518248
rect 334710 518236 334716 518248
rect 334768 518276 334774 518288
rect 343726 518276 343732 518288
rect 334768 518248 343732 518276
rect 334768 518236 334774 518248
rect 343726 518236 343732 518248
rect 343784 518276 343790 518288
rect 344370 518276 344376 518288
rect 343784 518248 344376 518276
rect 343784 518236 343790 518248
rect 344370 518236 344376 518248
rect 344428 518236 344434 518288
rect 354582 518236 354588 518288
rect 354640 518276 354646 518288
rect 429286 518276 429292 518288
rect 354640 518248 429292 518276
rect 354640 518236 354646 518248
rect 429286 518236 429292 518248
rect 429344 518236 429350 518288
rect 303614 518168 303620 518220
rect 303672 518208 303678 518220
rect 423674 518208 423680 518220
rect 303672 518180 423680 518208
rect 303672 518168 303678 518180
rect 423674 518168 423680 518180
rect 423732 518168 423738 518220
rect 436922 518168 436928 518220
rect 436980 518208 436986 518220
rect 445404 518208 445432 518304
rect 446398 518236 446404 518288
rect 446456 518276 446462 518288
rect 456058 518276 456064 518288
rect 446456 518248 456064 518276
rect 446456 518236 446462 518248
rect 456058 518236 456064 518248
rect 456116 518276 456122 518288
rect 465074 518276 465080 518288
rect 456116 518248 465080 518276
rect 456116 518236 456122 518248
rect 465074 518236 465080 518248
rect 465132 518236 465138 518288
rect 450170 518208 450176 518220
rect 436980 518180 445432 518208
rect 447796 518180 450176 518208
rect 436980 518168 436986 518180
rect 286962 518100 286968 518152
rect 287020 518140 287026 518152
rect 321738 518140 321744 518152
rect 287020 518112 321744 518140
rect 287020 518100 287026 518112
rect 321738 518100 321744 518112
rect 321796 518100 321802 518152
rect 331122 518100 331128 518152
rect 331180 518140 331186 518152
rect 340874 518140 340880 518152
rect 331180 518112 340880 518140
rect 331180 518100 331186 518112
rect 340874 518100 340880 518112
rect 340932 518100 340938 518152
rect 351822 518100 351828 518152
rect 351880 518140 351886 518152
rect 429194 518140 429200 518152
rect 351880 518112 429200 518140
rect 351880 518100 351886 518112
rect 429194 518100 429200 518112
rect 429252 518100 429258 518152
rect 440878 518100 440884 518152
rect 440936 518140 440942 518152
rect 447796 518140 447824 518180
rect 450170 518168 450176 518180
rect 450228 518208 450234 518220
rect 459554 518208 459560 518220
rect 450228 518180 459560 518208
rect 450228 518168 450234 518180
rect 459554 518168 459560 518180
rect 459612 518208 459618 518220
rect 467834 518208 467840 518220
rect 459612 518180 467840 518208
rect 459612 518168 459618 518180
rect 467834 518168 467840 518180
rect 467892 518168 467898 518220
rect 440936 518112 447824 518140
rect 440936 518100 440942 518112
rect 285582 518032 285588 518084
rect 285640 518072 285646 518084
rect 315850 518072 315856 518084
rect 285640 518044 315856 518072
rect 285640 518032 285646 518044
rect 315850 518032 315856 518044
rect 315908 518032 315914 518084
rect 315942 518032 315948 518084
rect 316000 518072 316006 518084
rect 324314 518072 324320 518084
rect 316000 518044 324320 518072
rect 316000 518032 316006 518044
rect 324314 518032 324320 518044
rect 324372 518072 324378 518084
rect 325510 518072 325516 518084
rect 324372 518044 325516 518072
rect 324372 518032 324378 518044
rect 325510 518032 325516 518044
rect 325568 518032 325574 518084
rect 325602 518032 325608 518084
rect 325660 518072 325666 518084
rect 339494 518072 339500 518084
rect 325660 518044 339500 518072
rect 325660 518032 325666 518044
rect 339494 518032 339500 518044
rect 339552 518032 339558 518084
rect 349062 518032 349068 518084
rect 349120 518072 349126 518084
rect 425330 518072 425336 518084
rect 349120 518044 425336 518072
rect 349120 518032 349126 518044
rect 425330 518032 425336 518044
rect 425388 518032 425394 518084
rect 432598 518032 432604 518084
rect 432656 518072 432662 518084
rect 442534 518072 442540 518084
rect 432656 518044 442540 518072
rect 432656 518032 432662 518044
rect 442534 518032 442540 518044
rect 442592 518032 442598 518084
rect 282822 517964 282828 518016
rect 282880 518004 282886 518016
rect 318794 518004 318800 518016
rect 282880 517976 318800 518004
rect 282880 517964 282886 517976
rect 318794 517964 318800 517976
rect 318852 517964 318858 518016
rect 328362 517964 328368 518016
rect 328420 518004 328426 518016
rect 339586 518004 339592 518016
rect 328420 517976 339592 518004
rect 328420 517964 328426 517976
rect 339586 517964 339592 517976
rect 339644 517964 339650 518016
rect 340598 517964 340604 518016
rect 340656 518004 340662 518016
rect 437474 518004 437480 518016
rect 340656 517976 437480 518004
rect 340656 517964 340662 517976
rect 437474 517964 437480 517976
rect 437532 517964 437538 518016
rect 439498 517964 439504 518016
rect 439556 518004 439562 518016
rect 448698 518004 448704 518016
rect 439556 517976 448704 518004
rect 439556 517964 439562 517976
rect 448698 517964 448704 517976
rect 448756 517964 448762 518016
rect 280062 517896 280068 517948
rect 280120 517936 280126 517948
rect 317506 517936 317512 517948
rect 280120 517908 317512 517936
rect 280120 517896 280126 517908
rect 317506 517896 317512 517908
rect 317564 517896 317570 517948
rect 322842 517896 322848 517948
rect 322900 517936 322906 517948
rect 338114 517936 338120 517948
rect 322900 517908 338120 517936
rect 322900 517896 322906 517908
rect 338114 517896 338120 517908
rect 338172 517896 338178 517948
rect 341518 517896 341524 517948
rect 341576 517936 341582 517948
rect 440234 517936 440240 517948
rect 341576 517908 440240 517936
rect 341576 517896 341582 517908
rect 440234 517896 440240 517908
rect 440292 517896 440298 517948
rect 444098 517896 444104 517948
rect 444156 517936 444162 517948
rect 469858 517936 469864 517948
rect 444156 517908 469864 517936
rect 444156 517896 444162 517908
rect 469858 517896 469864 517908
rect 469916 517896 469922 517948
rect 277302 517828 277308 517880
rect 277360 517868 277366 517880
rect 317414 517868 317420 517880
rect 277360 517840 317420 517868
rect 277360 517828 277366 517840
rect 317414 517828 317420 517840
rect 317472 517828 317478 517880
rect 321462 517828 321468 517880
rect 321520 517868 321526 517880
rect 336734 517868 336740 517880
rect 321520 517840 336740 517868
rect 321520 517828 321526 517840
rect 336734 517828 336740 517840
rect 336792 517828 336798 517880
rect 342990 517828 342996 517880
rect 343048 517868 343054 517880
rect 442994 517868 443000 517880
rect 343048 517840 443000 517868
rect 343048 517828 343054 517840
rect 442994 517828 443000 517840
rect 443052 517828 443058 517880
rect 445570 517828 445576 517880
rect 445628 517868 445634 517880
rect 476758 517868 476764 517880
rect 445628 517840 476764 517868
rect 445628 517828 445634 517840
rect 476758 517828 476764 517840
rect 476816 517828 476822 517880
rect 315942 517760 315948 517812
rect 316000 517800 316006 517812
rect 333974 517800 333980 517812
rect 316000 517772 333980 517800
rect 316000 517760 316006 517772
rect 333974 517760 333980 517772
rect 334032 517760 334038 517812
rect 344370 517760 344376 517812
rect 344428 517800 344434 517812
rect 445754 517800 445760 517812
rect 344428 517772 445760 517800
rect 344428 517760 344434 517772
rect 445754 517760 445760 517772
rect 445812 517760 445818 517812
rect 313182 517692 313188 517744
rect 313240 517732 313246 517744
rect 332686 517732 332692 517744
rect 313240 517704 332692 517732
rect 313240 517692 313246 517704
rect 332686 517692 332692 517704
rect 332744 517692 332750 517744
rect 333882 517692 333888 517744
rect 333940 517732 333946 517744
rect 342254 517732 342260 517744
rect 333940 517704 342260 517732
rect 333940 517692 333946 517704
rect 342254 517692 342260 517704
rect 342312 517692 342318 517744
rect 344278 517692 344284 517744
rect 344336 517732 344342 517744
rect 347866 517732 347872 517744
rect 344336 517704 347872 517732
rect 344336 517692 344342 517704
rect 347866 517692 347872 517704
rect 347924 517692 347930 517744
rect 447042 517692 447048 517744
rect 447100 517732 447106 517744
rect 473998 517732 474004 517744
rect 447100 517704 474004 517732
rect 447100 517692 447106 517704
rect 473998 517692 474004 517704
rect 474056 517692 474062 517744
rect 261110 517624 261116 517676
rect 261168 517664 261174 517676
rect 303614 517664 303620 517676
rect 261168 517636 303620 517664
rect 261168 517624 261174 517636
rect 303614 517624 303620 517636
rect 303672 517624 303678 517676
rect 304902 517624 304908 517676
rect 304960 517664 304966 517676
rect 329834 517664 329840 517676
rect 304960 517636 329840 517664
rect 304960 517624 304966 517636
rect 329834 517624 329840 517636
rect 329892 517624 329898 517676
rect 337378 517624 337384 517676
rect 337436 517664 337442 517676
rect 343634 517664 343640 517676
rect 337436 517636 343640 517664
rect 337436 517624 337442 517636
rect 343634 517624 343640 517636
rect 343692 517624 343698 517676
rect 438118 517624 438124 517676
rect 438176 517664 438182 517676
rect 447134 517664 447140 517676
rect 438176 517636 447140 517664
rect 438176 517624 438182 517636
rect 447134 517624 447140 517636
rect 447192 517624 447198 517676
rect 448330 517624 448336 517676
rect 448388 517664 448394 517676
rect 471238 517664 471244 517676
rect 448388 517636 471244 517664
rect 448388 517624 448394 517636
rect 471238 517624 471244 517636
rect 471296 517624 471302 517676
rect 310422 517556 310428 517608
rect 310480 517596 310486 517608
rect 332594 517596 332600 517608
rect 310480 517568 332600 517596
rect 310480 517556 310486 517568
rect 332594 517556 332600 517568
rect 332652 517556 332658 517608
rect 340782 517556 340788 517608
rect 340840 517596 340846 517608
rect 346394 517596 346400 517608
rect 340840 517568 346400 517596
rect 340840 517556 340846 517568
rect 346394 517556 346400 517568
rect 346452 517556 346458 517608
rect 436738 517556 436744 517608
rect 436796 517596 436802 517608
rect 437290 517596 437296 517608
rect 436796 517568 437296 517596
rect 436796 517556 436802 517568
rect 437290 517556 437296 517568
rect 437348 517596 437354 517608
rect 446398 517596 446404 517608
rect 437348 517568 446404 517596
rect 437348 517556 437354 517568
rect 446398 517556 446404 517568
rect 446456 517556 446462 517608
rect 266262 517488 266268 517540
rect 266320 517528 266326 517540
rect 312170 517528 312176 517540
rect 266320 517500 312176 517528
rect 266320 517488 266326 517500
rect 312170 517488 312176 517500
rect 312228 517488 312234 517540
rect 325510 517488 325516 517540
rect 325568 517528 325574 517540
rect 333790 517528 333796 517540
rect 325568 517500 333796 517528
rect 325568 517488 325574 517500
rect 333790 517488 333796 517500
rect 333848 517488 333854 517540
rect 339402 517488 339408 517540
rect 339460 517528 339466 517540
rect 345198 517528 345204 517540
rect 339460 517500 345204 517528
rect 339460 517488 339466 517500
rect 345198 517488 345204 517500
rect 345256 517488 345262 517540
rect 346302 517488 346308 517540
rect 346360 517528 346366 517540
rect 347774 517528 347780 517540
rect 346360 517500 347780 517528
rect 346360 517488 346366 517500
rect 347774 517488 347780 517500
rect 347832 517488 347838 517540
rect 434162 517488 434168 517540
rect 434220 517528 434226 517540
rect 443178 517528 443184 517540
rect 434220 517500 443184 517528
rect 434220 517488 434226 517500
rect 443178 517488 443184 517500
rect 443236 517488 443242 517540
rect 445478 517488 445484 517540
rect 445536 517528 445542 517540
rect 479518 517528 479524 517540
rect 445536 517500 479524 517528
rect 445536 517488 445542 517500
rect 479518 517488 479524 517500
rect 479576 517488 479582 517540
rect 543366 514768 543372 514820
rect 543424 514808 543430 514820
rect 543550 514808 543556 514820
rect 543424 514780 543556 514808
rect 543424 514768 543430 514780
rect 543550 514768 543556 514780
rect 543608 514768 543614 514820
rect 379606 514020 379612 514072
rect 379664 514060 379670 514072
rect 379790 514060 379796 514072
rect 379664 514032 379796 514060
rect 379664 514020 379670 514032
rect 379790 514020 379796 514032
rect 379848 514020 379854 514072
rect 434070 511980 434076 512032
rect 434128 512020 434134 512032
rect 434162 512020 434168 512032
rect 434128 511992 434168 512020
rect 434128 511980 434134 511992
rect 434162 511980 434168 511992
rect 434220 511980 434226 512032
rect 3234 509260 3240 509312
rect 3292 509300 3298 509312
rect 539502 509300 539508 509312
rect 3292 509272 539508 509300
rect 3292 509260 3298 509272
rect 539502 509260 539508 509272
rect 539560 509260 539566 509312
rect 555418 509260 555424 509312
rect 555476 509300 555482 509312
rect 580166 509300 580172 509312
rect 555476 509272 580172 509300
rect 555476 509260 555482 509272
rect 580166 509260 580172 509272
rect 580224 509260 580230 509312
rect 543274 502324 543280 502376
rect 543332 502364 543338 502376
rect 543550 502364 543556 502376
rect 543332 502336 543556 502364
rect 543332 502324 543338 502336
rect 543550 502324 543556 502336
rect 543608 502324 543614 502376
rect 379606 499536 379612 499588
rect 379664 499576 379670 499588
rect 379790 499576 379796 499588
rect 379664 499548 379796 499576
rect 379664 499536 379670 499548
rect 379790 499536 379796 499548
rect 379848 499536 379854 499588
rect 571978 498176 571984 498228
rect 572036 498216 572042 498228
rect 580166 498216 580172 498228
rect 572036 498188 580172 498216
rect 572036 498176 572042 498188
rect 580166 498176 580172 498188
rect 580224 498176 580230 498228
rect 3326 495456 3332 495508
rect 3384 495496 3390 495508
rect 540974 495496 540980 495508
rect 3384 495468 540980 495496
rect 3384 495456 3390 495468
rect 540974 495456 540980 495468
rect 541032 495456 541038 495508
rect 379606 494708 379612 494760
rect 379664 494748 379670 494760
rect 379790 494748 379796 494760
rect 379664 494720 379796 494748
rect 379664 494708 379670 494720
rect 379790 494708 379796 494720
rect 379848 494708 379854 494760
rect 433610 492600 433616 492652
rect 433668 492640 433674 492652
rect 433886 492640 433892 492652
rect 433668 492612 433892 492640
rect 433668 492600 433674 492612
rect 433886 492600 433892 492612
rect 433944 492600 433950 492652
rect 543274 492600 543280 492652
rect 543332 492640 543338 492652
rect 543550 492640 543556 492652
rect 543332 492612 543556 492640
rect 543332 492600 543338 492612
rect 543550 492600 543556 492612
rect 543608 492600 543614 492652
rect 398742 487772 398748 487824
rect 398800 487812 398806 487824
rect 539410 487812 539416 487824
rect 398800 487784 539416 487812
rect 398800 487772 398806 487784
rect 539410 487772 539416 487784
rect 539468 487772 539474 487824
rect 544562 485800 544568 485852
rect 544620 485840 544626 485852
rect 580166 485840 580172 485852
rect 544620 485812 580172 485840
rect 544620 485800 544626 485812
rect 580166 485800 580172 485812
rect 580224 485800 580230 485852
rect 281718 482944 281724 482996
rect 281776 482984 281782 482996
rect 282822 482984 282828 482996
rect 281776 482956 282828 482984
rect 281776 482944 281782 482956
rect 282822 482944 282828 482956
rect 282880 482944 282886 482996
rect 311802 482944 311808 482996
rect 311860 482984 311866 482996
rect 366450 482984 366456 482996
rect 311860 482956 366456 482984
rect 311860 482944 311866 482956
rect 366450 482944 366456 482956
rect 366508 482944 366514 482996
rect 371602 482944 371608 482996
rect 371660 482984 371666 482996
rect 417510 482984 417516 482996
rect 371660 482956 417516 482984
rect 371660 482944 371666 482956
rect 417510 482944 417516 482956
rect 417568 482944 417574 482996
rect 433150 482944 433156 482996
rect 433208 482984 433214 482996
rect 439498 482984 439504 482996
rect 433208 482956 439504 482984
rect 433208 482944 433214 482956
rect 439498 482944 439504 482956
rect 439556 482944 439562 482996
rect 455322 482944 455328 482996
rect 455380 482984 455386 482996
rect 507762 482984 507768 482996
rect 455380 482956 507768 482984
rect 455380 482944 455386 482956
rect 507762 482944 507768 482956
rect 507820 482944 507826 482996
rect 307570 482876 307576 482928
rect 307628 482916 307634 482928
rect 307628 482888 386644 482916
rect 307628 482876 307634 482888
rect 297450 482808 297456 482860
rect 297508 482848 297514 482860
rect 386506 482848 386512 482860
rect 297508 482820 386512 482848
rect 297508 482808 297514 482820
rect 386506 482808 386512 482820
rect 386564 482808 386570 482860
rect 386616 482848 386644 482888
rect 386966 482876 386972 482928
rect 387024 482916 387030 482928
rect 387702 482916 387708 482928
rect 387024 482888 387708 482916
rect 387024 482876 387030 482888
rect 387702 482876 387708 482888
rect 387760 482876 387766 482928
rect 453942 482876 453948 482928
rect 454000 482916 454006 482928
rect 505186 482916 505192 482928
rect 454000 482888 505192 482916
rect 454000 482876 454006 482888
rect 505186 482876 505192 482888
rect 505244 482876 505250 482928
rect 389542 482848 389548 482860
rect 386616 482820 389548 482848
rect 389542 482808 389548 482820
rect 389600 482808 389606 482860
rect 456702 482808 456708 482860
rect 456760 482848 456766 482860
rect 510246 482848 510252 482860
rect 456760 482820 510252 482848
rect 456760 482808 456766 482820
rect 510246 482808 510252 482820
rect 510304 482808 510310 482860
rect 297542 482740 297548 482792
rect 297600 482780 297606 482792
rect 394694 482780 394700 482792
rect 297600 482752 394700 482780
rect 297600 482740 297606 482752
rect 394694 482740 394700 482752
rect 394752 482740 394758 482792
rect 430666 482740 430672 482792
rect 430724 482780 430730 482792
rect 438118 482780 438124 482792
rect 430724 482752 438124 482780
rect 430724 482740 430730 482752
rect 438118 482740 438124 482752
rect 438176 482740 438182 482792
rect 458082 482740 458088 482792
rect 458140 482780 458146 482792
rect 512822 482780 512828 482792
rect 458140 482752 512828 482780
rect 458140 482740 458146 482752
rect 512822 482740 512828 482752
rect 512880 482740 512886 482792
rect 284294 482672 284300 482724
rect 284352 482712 284358 482724
rect 285582 482712 285588 482724
rect 284352 482684 285588 482712
rect 284352 482672 284358 482684
rect 285582 482672 285588 482684
rect 285640 482672 285646 482724
rect 297634 482672 297640 482724
rect 297692 482712 297698 482724
rect 397270 482712 397276 482724
rect 297692 482684 397276 482712
rect 297692 482672 297698 482684
rect 397270 482672 397276 482684
rect 397328 482672 397334 482724
rect 428090 482672 428096 482724
rect 428148 482712 428154 482724
rect 436738 482712 436744 482724
rect 428148 482684 436744 482712
rect 428148 482672 428154 482684
rect 436738 482672 436744 482684
rect 436796 482672 436802 482724
rect 459462 482672 459468 482724
rect 459520 482712 459526 482724
rect 515398 482712 515404 482724
rect 459520 482684 515404 482712
rect 459520 482672 459526 482684
rect 515398 482672 515404 482684
rect 515456 482672 515462 482724
rect 297726 482604 297732 482656
rect 297784 482644 297790 482656
rect 399846 482644 399852 482656
rect 297784 482616 399852 482644
rect 297784 482604 297790 482616
rect 399846 482604 399852 482616
rect 399904 482604 399910 482656
rect 425514 482604 425520 482656
rect 425572 482644 425578 482656
rect 436922 482644 436928 482656
rect 425572 482616 436928 482644
rect 425572 482604 425578 482616
rect 436922 482604 436928 482616
rect 436980 482604 436986 482656
rect 460842 482604 460848 482656
rect 460900 482644 460906 482656
rect 517974 482644 517980 482656
rect 460900 482616 517980 482644
rect 460900 482604 460906 482616
rect 517974 482604 517980 482616
rect 518032 482604 518038 482656
rect 279142 482536 279148 482588
rect 279200 482576 279206 482588
rect 280062 482576 280068 482588
rect 279200 482548 280068 482576
rect 279200 482536 279206 482548
rect 280062 482536 280068 482548
rect 280120 482536 280126 482588
rect 297818 482536 297824 482588
rect 297876 482576 297882 482588
rect 402422 482576 402428 482588
rect 297876 482548 402428 482576
rect 297876 482536 297882 482548
rect 402422 482536 402428 482548
rect 402480 482536 402486 482588
rect 412726 482536 412732 482588
rect 412784 482576 412790 482588
rect 413922 482576 413928 482588
rect 412784 482548 413928 482576
rect 412784 482536 412790 482548
rect 413922 482536 413928 482548
rect 413980 482536 413986 482588
rect 422938 482536 422944 482588
rect 422996 482576 423002 482588
rect 435358 482576 435364 482588
rect 422996 482548 435364 482576
rect 422996 482536 423002 482548
rect 435358 482536 435364 482548
rect 435416 482536 435422 482588
rect 460750 482536 460756 482588
rect 460808 482576 460814 482588
rect 520550 482576 520556 482588
rect 460808 482548 520556 482576
rect 460808 482536 460814 482548
rect 520550 482536 520556 482548
rect 520608 482536 520614 482588
rect 297910 482468 297916 482520
rect 297968 482508 297974 482520
rect 404998 482508 405004 482520
rect 297968 482480 405004 482508
rect 297968 482468 297974 482480
rect 404998 482468 405004 482480
rect 405056 482468 405062 482520
rect 433242 482468 433248 482520
rect 433300 482508 433306 482520
rect 458910 482508 458916 482520
rect 433300 482480 458916 482508
rect 433300 482468 433306 482480
rect 458910 482468 458916 482480
rect 458968 482468 458974 482520
rect 463602 482468 463608 482520
rect 463660 482508 463666 482520
rect 525702 482508 525708 482520
rect 463660 482480 525708 482508
rect 463660 482468 463666 482480
rect 525702 482468 525708 482480
rect 525760 482468 525766 482520
rect 298002 482400 298008 482452
rect 298060 482440 298066 482452
rect 407574 482440 407580 482452
rect 298060 482412 407580 482440
rect 298060 482400 298066 482412
rect 407574 482400 407580 482412
rect 407632 482400 407638 482452
rect 434622 482400 434628 482452
rect 434680 482440 434686 482452
rect 461486 482440 461492 482452
rect 434680 482412 461492 482440
rect 434680 482400 434686 482412
rect 461486 482400 461492 482412
rect 461544 482400 461550 482452
rect 462222 482400 462228 482452
rect 462280 482440 462286 482452
rect 523126 482440 523132 482452
rect 462280 482412 523132 482440
rect 462280 482400 462286 482412
rect 523126 482400 523132 482412
rect 523184 482400 523190 482452
rect 297358 482332 297364 482384
rect 297416 482372 297422 482384
rect 415302 482372 415308 482384
rect 297416 482344 415308 482372
rect 297416 482332 297422 482344
rect 415302 482332 415308 482344
rect 415360 482332 415366 482384
rect 420362 482332 420368 482384
rect 420420 482372 420426 482384
rect 433794 482372 433800 482384
rect 420420 482344 433800 482372
rect 420420 482332 420426 482344
rect 433794 482332 433800 482344
rect 433852 482332 433858 482384
rect 436002 482332 436008 482384
rect 436060 482372 436066 482384
rect 464062 482372 464068 482384
rect 436060 482344 464068 482372
rect 436060 482332 436066 482344
rect 464062 482332 464068 482344
rect 464120 482332 464126 482384
rect 464982 482332 464988 482384
rect 465040 482372 465046 482384
rect 528278 482372 528284 482384
rect 465040 482344 528284 482372
rect 465040 482332 465046 482344
rect 528278 482332 528284 482344
rect 528336 482332 528342 482384
rect 261202 482264 261208 482316
rect 261260 482304 261266 482316
rect 261260 482276 374132 482304
rect 261260 482264 261266 482276
rect 310330 482196 310336 482248
rect 310388 482236 310394 482248
rect 363874 482236 363880 482248
rect 310388 482208 363880 482236
rect 310388 482196 310394 482208
rect 363874 482196 363880 482208
rect 363932 482196 363938 482248
rect 310238 482128 310244 482180
rect 310296 482168 310302 482180
rect 361298 482168 361304 482180
rect 310296 482140 361304 482168
rect 310296 482128 310302 482140
rect 361298 482128 361304 482140
rect 361356 482128 361362 482180
rect 309042 482060 309048 482112
rect 309100 482100 309106 482112
rect 358722 482100 358728 482112
rect 309100 482072 358728 482100
rect 309100 482060 309106 482072
rect 358722 482060 358728 482072
rect 358780 482060 358786 482112
rect 374104 482100 374132 482276
rect 376754 482264 376760 482316
rect 376812 482304 376818 482316
rect 378042 482304 378048 482316
rect 376812 482276 378048 482304
rect 376812 482264 376818 482276
rect 378042 482264 378048 482276
rect 378100 482264 378106 482316
rect 386506 482264 386512 482316
rect 386564 482304 386570 482316
rect 392118 482304 392124 482316
rect 386564 482276 392124 482304
rect 386564 482264 386570 482276
rect 392118 482264 392124 482276
rect 392176 482264 392182 482316
rect 417786 482264 417792 482316
rect 417844 482304 417850 482316
rect 432598 482304 432604 482316
rect 417844 482276 432604 482304
rect 417844 482264 417850 482276
rect 432598 482264 432604 482276
rect 432656 482264 432662 482316
rect 437382 482264 437388 482316
rect 437440 482304 437446 482316
rect 466638 482304 466644 482316
rect 437440 482276 466644 482304
rect 437440 482264 437446 482276
rect 466638 482264 466644 482276
rect 466696 482264 466702 482316
rect 467742 482264 467748 482316
rect 467800 482304 467806 482316
rect 533430 482304 533436 482316
rect 467800 482276 533436 482304
rect 467800 482264 467806 482276
rect 533430 482264 533436 482276
rect 533488 482264 533494 482316
rect 374178 482196 374184 482248
rect 374236 482236 374242 482248
rect 417418 482236 417424 482248
rect 374236 482208 417424 482236
rect 374236 482196 374242 482208
rect 417418 482196 417424 482208
rect 417476 482196 417482 482248
rect 453850 482196 453856 482248
rect 453908 482236 453914 482248
rect 502610 482236 502616 482248
rect 453908 482208 502616 482236
rect 453908 482196 453914 482208
rect 502610 482196 502616 482208
rect 502668 482196 502674 482248
rect 435818 482128 435824 482180
rect 435876 482168 435882 482180
rect 440878 482168 440884 482180
rect 435876 482140 440884 482168
rect 435876 482128 435882 482140
rect 440878 482128 440884 482140
rect 440936 482128 440942 482180
rect 452562 482128 452568 482180
rect 452620 482168 452626 482180
rect 500034 482168 500040 482180
rect 452620 482140 500040 482168
rect 452620 482128 452626 482140
rect 500034 482128 500040 482140
rect 500092 482128 500098 482180
rect 379790 482100 379796 482112
rect 374104 482072 379796 482100
rect 379790 482060 379796 482072
rect 379848 482060 379854 482112
rect 451182 482060 451188 482112
rect 451240 482100 451246 482112
rect 497458 482100 497464 482112
rect 451240 482072 497464 482100
rect 451240 482060 451246 482072
rect 497458 482060 497464 482072
rect 497516 482060 497522 482112
rect 276566 481992 276572 482044
rect 276624 482032 276630 482044
rect 277302 482032 277308 482044
rect 276624 482004 277308 482032
rect 276624 481992 276630 482004
rect 277302 481992 277308 482004
rect 277360 481992 277366 482044
rect 292022 481992 292028 482044
rect 292080 482032 292086 482044
rect 320174 482032 320180 482044
rect 292080 482004 320180 482032
rect 292080 481992 292086 482004
rect 320174 481992 320180 482004
rect 320232 481992 320238 482044
rect 320266 481992 320272 482044
rect 320324 482032 320330 482044
rect 321462 482032 321468 482044
rect 320324 482004 321468 482032
rect 320324 481992 320330 482004
rect 321462 481992 321468 482004
rect 321520 481992 321526 482044
rect 321554 481992 321560 482044
rect 321612 482032 321618 482044
rect 324498 482032 324504 482044
rect 321612 482004 324504 482032
rect 321612 481992 321618 482004
rect 324498 481992 324504 482004
rect 324556 481992 324562 482044
rect 333054 481992 333060 482044
rect 333112 482032 333118 482044
rect 333882 482032 333888 482044
rect 333112 482004 333888 482032
rect 333112 481992 333118 482004
rect 333882 481992 333888 482004
rect 333940 481992 333946 482044
rect 338206 481992 338212 482044
rect 338264 482032 338270 482044
rect 339402 482032 339408 482044
rect 338264 482004 339408 482032
rect 338264 481992 338270 482004
rect 339402 481992 339408 482004
rect 339460 481992 339466 482044
rect 343358 481992 343364 482044
rect 343416 482032 343422 482044
rect 344278 482032 344284 482044
rect 343416 482004 344284 482032
rect 343416 481992 343422 482004
rect 344278 481992 344284 482004
rect 344336 481992 344342 482044
rect 351086 481992 351092 482044
rect 351144 482032 351150 482044
rect 351822 482032 351828 482044
rect 351144 482004 351828 482032
rect 351144 481992 351150 482004
rect 351822 481992 351828 482004
rect 351880 481992 351886 482044
rect 353662 481992 353668 482044
rect 353720 482032 353726 482044
rect 354582 482032 354588 482044
rect 353720 482004 354588 482032
rect 353720 481992 353726 482004
rect 354582 481992 354588 482004
rect 354640 481992 354646 482044
rect 449802 481992 449808 482044
rect 449860 482032 449866 482044
rect 494882 482032 494888 482044
rect 449860 482004 494888 482032
rect 449860 481992 449866 482004
rect 494882 481992 494888 482004
rect 494940 481992 494946 482044
rect 294506 481924 294512 481976
rect 294564 481964 294570 481976
rect 324406 481964 324412 481976
rect 294564 481936 324412 481964
rect 294564 481924 294570 481936
rect 324406 481924 324412 481936
rect 324464 481924 324470 481976
rect 325786 481924 325792 481976
rect 325844 481964 325850 481976
rect 325844 481936 330524 481964
rect 325844 481924 325850 481936
rect 297082 481856 297088 481908
rect 297140 481896 297146 481908
rect 325694 481896 325700 481908
rect 297140 481868 325700 481896
rect 297140 481856 297146 481868
rect 325694 481856 325700 481868
rect 325752 481856 325758 481908
rect 299658 481788 299664 481840
rect 299716 481828 299722 481840
rect 327166 481828 327172 481840
rect 299716 481800 327172 481828
rect 299716 481788 299722 481800
rect 327166 481788 327172 481800
rect 327224 481788 327230 481840
rect 302234 481720 302240 481772
rect 302292 481760 302298 481772
rect 328454 481760 328460 481772
rect 302292 481732 328460 481760
rect 302292 481720 302298 481732
rect 328454 481720 328460 481732
rect 328512 481720 328518 481772
rect 330496 481760 330524 481936
rect 442902 481924 442908 481976
rect 442960 481964 442966 481976
rect 479426 481964 479432 481976
rect 442960 481936 479432 481964
rect 442960 481924 442966 481936
rect 479426 481924 479432 481936
rect 479484 481924 479490 481976
rect 479518 481924 479524 481976
rect 479576 481964 479582 481976
rect 484578 481964 484584 481976
rect 479576 481936 484584 481964
rect 479576 481924 479582 481936
rect 484578 481924 484584 481936
rect 484636 481924 484642 481976
rect 356146 481856 356152 481908
rect 356204 481896 356210 481908
rect 357342 481896 357348 481908
rect 356204 481868 357348 481896
rect 356204 481856 356210 481868
rect 357342 481856 357348 481868
rect 357400 481856 357406 481908
rect 441522 481856 441528 481908
rect 441580 481896 441586 481908
rect 476942 481896 476948 481908
rect 441580 481868 476948 481896
rect 441580 481856 441586 481868
rect 476942 481856 476948 481868
rect 477000 481856 477006 481908
rect 487154 481896 487160 481908
rect 477052 481868 487160 481896
rect 440142 481788 440148 481840
rect 440200 481828 440206 481840
rect 474366 481828 474372 481840
rect 440200 481800 474372 481828
rect 440200 481788 440206 481800
rect 474366 481788 474372 481800
rect 474424 481788 474430 481840
rect 476758 481788 476764 481840
rect 476816 481828 476822 481840
rect 477052 481828 477080 481868
rect 487154 481856 487160 481868
rect 487212 481856 487218 481908
rect 489730 481828 489736 481840
rect 476816 481800 477080 481828
rect 477144 481800 489736 481828
rect 476816 481788 476822 481800
rect 335354 481760 335360 481772
rect 330496 481732 335360 481760
rect 335354 481720 335360 481732
rect 335412 481720 335418 481772
rect 335630 481720 335636 481772
rect 335688 481760 335694 481772
rect 337378 481760 337384 481772
rect 335688 481732 337384 481760
rect 335688 481720 335694 481732
rect 337378 481720 337384 481732
rect 337436 481720 337442 481772
rect 438762 481720 438768 481772
rect 438820 481760 438826 481772
rect 471790 481760 471796 481772
rect 438820 481732 471796 481760
rect 438820 481720 438826 481732
rect 471790 481720 471796 481732
rect 471848 481720 471854 481772
rect 473998 481720 474004 481772
rect 474056 481760 474062 481772
rect 477144 481760 477172 481800
rect 489730 481788 489736 481800
rect 489788 481788 489794 481840
rect 474056 481732 477172 481760
rect 474056 481720 474062 481732
rect 477218 481720 477224 481772
rect 477276 481760 477282 481772
rect 492306 481760 492312 481772
rect 477276 481732 492312 481760
rect 477276 481720 477282 481732
rect 492306 481720 492312 481732
rect 492364 481720 492370 481772
rect 315114 481652 315120 481704
rect 315172 481692 315178 481704
rect 315942 481692 315948 481704
rect 315172 481664 315948 481692
rect 315172 481652 315178 481664
rect 315942 481652 315948 481664
rect 316000 481652 316006 481704
rect 317690 481652 317696 481704
rect 317748 481692 317754 481704
rect 325694 481692 325700 481704
rect 317748 481664 325700 481692
rect 317748 481652 317754 481664
rect 325694 481652 325700 481664
rect 325752 481652 325758 481704
rect 438670 481652 438676 481704
rect 438728 481692 438734 481704
rect 469214 481692 469220 481704
rect 438728 481664 469220 481692
rect 438728 481652 438734 481664
rect 469214 481652 469220 481664
rect 469272 481652 469278 481704
rect 469858 481652 469864 481704
rect 469916 481692 469922 481704
rect 477126 481692 477132 481704
rect 469916 481664 473860 481692
rect 469916 481652 469922 481664
rect 473832 481556 473860 481664
rect 474016 481664 477132 481692
rect 474016 481556 474044 481664
rect 477126 481652 477132 481664
rect 477184 481652 477190 481704
rect 477310 481652 477316 481704
rect 477368 481692 477374 481704
rect 482002 481692 482008 481704
rect 477368 481664 482008 481692
rect 477368 481652 477374 481664
rect 482002 481652 482008 481664
rect 482060 481652 482066 481704
rect 473832 481528 474044 481556
rect 3142 480224 3148 480276
rect 3200 480264 3206 480276
rect 540606 480264 540612 480276
rect 3200 480236 540612 480264
rect 3200 480224 3206 480236
rect 540606 480224 540612 480236
rect 540664 480224 540670 480276
rect 528462 479816 528468 479868
rect 528520 479856 528526 479868
rect 541802 479856 541808 479868
rect 528520 479828 541808 479856
rect 528520 479816 528526 479828
rect 541802 479816 541808 479828
rect 541860 479816 541866 479868
rect 300762 479748 300768 479800
rect 300820 479788 300826 479800
rect 541894 479788 541900 479800
rect 300820 479760 541900 479788
rect 300820 479748 300826 479760
rect 541894 479748 541900 479760
rect 541952 479748 541958 479800
rect 235902 479680 235908 479732
rect 235960 479720 235966 479732
rect 541986 479720 541992 479732
rect 235960 479692 541992 479720
rect 235960 479680 235966 479692
rect 541986 479680 541992 479692
rect 542044 479680 542050 479732
rect 171042 479612 171048 479664
rect 171100 479652 171106 479664
rect 542078 479652 542084 479664
rect 171100 479624 542084 479652
rect 171100 479612 171106 479624
rect 542078 479612 542084 479624
rect 542136 479612 542142 479664
rect 106182 479544 106188 479596
rect 106240 479584 106246 479596
rect 542170 479584 542176 479596
rect 106240 479556 542176 479584
rect 106240 479544 106246 479556
rect 542170 479544 542176 479556
rect 542228 479544 542234 479596
rect 3510 479476 3516 479528
rect 3568 479516 3574 479528
rect 540514 479516 540520 479528
rect 3568 479488 540520 479516
rect 3568 479476 3574 479488
rect 540514 479476 540520 479488
rect 540572 479476 540578 479528
rect 260650 479136 260656 479188
rect 260708 479176 260714 479188
rect 540882 479176 540888 479188
rect 260708 479148 540888 479176
rect 260708 479136 260714 479148
rect 540882 479136 540888 479148
rect 540940 479136 540946 479188
rect 260558 479068 260564 479120
rect 260616 479108 260622 479120
rect 540790 479108 540796 479120
rect 260616 479080 540796 479108
rect 260616 479068 260622 479080
rect 540790 479068 540796 479080
rect 540848 479068 540854 479120
rect 260374 479000 260380 479052
rect 260432 479040 260438 479052
rect 543458 479040 543464 479052
rect 260432 479012 543464 479040
rect 260432 479000 260438 479012
rect 543458 479000 543464 479012
rect 543516 479000 543522 479052
rect 260098 478932 260104 478984
rect 260156 478972 260162 478984
rect 542446 478972 542452 478984
rect 260156 478944 542452 478972
rect 260156 478932 260162 478944
rect 542446 478932 542452 478944
rect 542504 478932 542510 478984
rect 135162 478864 135168 478916
rect 135220 478904 135226 478916
rect 256694 478904 256700 478916
rect 135220 478876 256700 478904
rect 135220 478864 135226 478876
rect 256694 478864 256700 478876
rect 256752 478864 256758 478916
rect 259914 478864 259920 478916
rect 259972 478904 259978 478916
rect 543182 478904 543188 478916
rect 259972 478876 543188 478904
rect 259972 478864 259978 478876
rect 543182 478864 543188 478876
rect 543240 478864 543246 478916
rect 259822 478524 259828 478576
rect 259880 478564 259886 478576
rect 540698 478564 540704 478576
rect 259880 478536 540704 478564
rect 259880 478524 259886 478536
rect 540698 478524 540704 478536
rect 540756 478524 540762 478576
rect 260742 478456 260748 478508
rect 260800 478496 260806 478508
rect 542722 478496 542728 478508
rect 260800 478468 542728 478496
rect 260800 478456 260806 478468
rect 542722 478456 542728 478468
rect 542780 478456 542786 478508
rect 260466 478388 260472 478440
rect 260524 478428 260530 478440
rect 542630 478428 542636 478440
rect 260524 478400 542636 478428
rect 260524 478388 260530 478400
rect 542630 478388 542636 478400
rect 542688 478388 542694 478440
rect 260282 478320 260288 478372
rect 260340 478360 260346 478372
rect 543550 478360 543556 478372
rect 260340 478332 543556 478360
rect 260340 478320 260346 478332
rect 543550 478320 543556 478332
rect 543608 478320 543614 478372
rect 3694 478252 3700 478304
rect 3752 478292 3758 478304
rect 542906 478292 542912 478304
rect 3752 478264 542912 478292
rect 3752 478252 3758 478264
rect 542906 478252 542912 478264
rect 542964 478252 542970 478304
rect 3418 478184 3424 478236
rect 3476 478224 3482 478236
rect 542814 478224 542820 478236
rect 3476 478196 542820 478224
rect 3476 478184 3482 478196
rect 542814 478184 542820 478196
rect 542872 478184 542878 478236
rect 3602 478116 3608 478168
rect 3660 478156 3666 478168
rect 542998 478156 543004 478168
rect 3660 478128 543004 478156
rect 3660 478116 3666 478128
rect 542998 478116 543004 478128
rect 543056 478116 543062 478168
rect 260006 478048 260012 478100
rect 260064 478088 260070 478100
rect 543090 478088 543096 478100
rect 260064 478060 543096 478088
rect 260064 478048 260070 478060
rect 543090 478048 543096 478060
rect 543148 478048 543154 478100
rect 260190 477980 260196 478032
rect 260248 478020 260254 478032
rect 543274 478020 543280 478032
rect 260248 477992 543280 478020
rect 260248 477980 260254 477992
rect 543274 477980 543280 477992
rect 543332 477980 543338 478032
rect 133782 476076 133788 476128
rect 133840 476116 133846 476128
rect 256694 476116 256700 476128
rect 133840 476088 256700 476116
rect 133840 476076 133846 476088
rect 256694 476076 256700 476088
rect 256752 476076 256758 476128
rect 543366 476076 543372 476128
rect 543424 476116 543430 476128
rect 543642 476116 543648 476128
rect 543424 476088 543648 476116
rect 543424 476076 543430 476088
rect 543642 476076 543648 476088
rect 543700 476076 543706 476128
rect 132402 473356 132408 473408
rect 132460 473396 132466 473408
rect 256694 473396 256700 473408
rect 132460 473368 256700 473396
rect 132460 473356 132466 473368
rect 256694 473356 256700 473368
rect 256752 473356 256758 473408
rect 131022 471996 131028 472048
rect 131080 472036 131086 472048
rect 256694 472036 256700 472048
rect 131080 472008 256700 472036
rect 131080 471996 131086 472008
rect 256694 471996 256700 472008
rect 256752 471996 256758 472048
rect 129642 469208 129648 469260
rect 129700 469248 129706 469260
rect 256694 469248 256700 469260
rect 129700 469220 256700 469248
rect 129700 469208 129706 469220
rect 256694 469208 256700 469220
rect 256752 469208 256758 469260
rect 128262 467848 128268 467900
rect 128320 467888 128326 467900
rect 256694 467888 256700 467900
rect 128320 467860 256700 467888
rect 128320 467848 128326 467860
rect 256694 467848 256700 467860
rect 256752 467848 256758 467900
rect 126882 465060 126888 465112
rect 126940 465100 126946 465112
rect 256694 465100 256700 465112
rect 126940 465072 256700 465100
rect 126940 465060 126946 465072
rect 256694 465060 256700 465072
rect 256752 465060 256758 465112
rect 125502 463700 125508 463752
rect 125560 463740 125566 463752
rect 256694 463740 256700 463752
rect 125560 463712 256700 463740
rect 125560 463700 125566 463712
rect 256694 463700 256700 463712
rect 256752 463700 256758 463752
rect 567838 462340 567844 462392
rect 567896 462380 567902 462392
rect 580166 462380 580172 462392
rect 567896 462352 580172 462380
rect 567896 462340 567902 462352
rect 580166 462340 580172 462352
rect 580224 462340 580230 462392
rect 125410 460912 125416 460964
rect 125468 460952 125474 460964
rect 256694 460952 256700 460964
rect 125468 460924 256700 460952
rect 125468 460912 125474 460924
rect 256694 460912 256700 460924
rect 256752 460912 256758 460964
rect 543366 460912 543372 460964
rect 543424 460952 543430 460964
rect 543642 460952 543648 460964
rect 543424 460924 543648 460952
rect 543424 460912 543430 460924
rect 543642 460912 543648 460924
rect 543700 460912 543706 460964
rect 124122 459552 124128 459604
rect 124180 459592 124186 459604
rect 256694 459592 256700 459604
rect 124180 459564 256700 459592
rect 124180 459552 124186 459564
rect 256694 459552 256700 459564
rect 256752 459552 256758 459604
rect 122742 456764 122748 456816
rect 122800 456804 122806 456816
rect 256694 456804 256700 456816
rect 122800 456776 256700 456804
rect 122800 456764 122806 456776
rect 256694 456764 256700 456776
rect 256752 456764 256758 456816
rect 121362 455404 121368 455456
rect 121420 455444 121426 455456
rect 256694 455444 256700 455456
rect 121420 455416 256700 455444
rect 121420 455404 121426 455416
rect 256694 455404 256700 455416
rect 256752 455404 256758 455456
rect 119982 452616 119988 452668
rect 120040 452656 120046 452668
rect 256694 452656 256700 452668
rect 120040 452628 256700 452656
rect 120040 452616 120046 452628
rect 256694 452616 256700 452628
rect 256752 452616 256758 452668
rect 3418 452548 3424 452600
rect 3476 452588 3482 452600
rect 259822 452588 259828 452600
rect 3476 452560 259828 452588
rect 3476 452548 3482 452560
rect 259822 452548 259828 452560
rect 259880 452548 259886 452600
rect 542354 451936 542360 451988
rect 542412 451976 542418 451988
rect 543366 451976 543372 451988
rect 542412 451948 543372 451976
rect 542412 451936 542418 451948
rect 543366 451936 543372 451948
rect 543424 451936 543430 451988
rect 118602 451256 118608 451308
rect 118660 451296 118666 451308
rect 256694 451296 256700 451308
rect 118660 451268 256700 451296
rect 118660 451256 118666 451268
rect 256694 451256 256700 451268
rect 256752 451256 256758 451308
rect 563790 451256 563796 451308
rect 563848 451296 563854 451308
rect 580166 451296 580172 451308
rect 563848 451268 580172 451296
rect 563848 451256 563854 451268
rect 580166 451256 580172 451268
rect 580224 451256 580230 451308
rect 117222 448536 117228 448588
rect 117280 448576 117286 448588
rect 256694 448576 256700 448588
rect 117280 448548 256700 448576
rect 117280 448536 117286 448548
rect 256694 448536 256700 448548
rect 256752 448536 256758 448588
rect 117130 445748 117136 445800
rect 117188 445788 117194 445800
rect 256694 445788 256700 445800
rect 117188 445760 256700 445788
rect 117188 445748 117194 445760
rect 256694 445748 256700 445760
rect 256752 445748 256758 445800
rect 542354 445272 542360 445324
rect 542412 445312 542418 445324
rect 543734 445312 543740 445324
rect 542412 445284 543740 445312
rect 542412 445272 542418 445284
rect 543734 445272 543740 445284
rect 543792 445272 543798 445324
rect 115842 444388 115848 444440
rect 115900 444428 115906 444440
rect 256694 444428 256700 444440
rect 115900 444400 256700 444428
rect 115900 444388 115906 444400
rect 256694 444388 256700 444400
rect 256752 444388 256758 444440
rect 114462 441600 114468 441652
rect 114520 441640 114526 441652
rect 256694 441640 256700 441652
rect 114520 441612 256700 441640
rect 114520 441600 114526 441612
rect 256694 441600 256700 441612
rect 256752 441600 256758 441652
rect 543366 441600 543372 441652
rect 543424 441640 543430 441652
rect 543734 441640 543740 441652
rect 543424 441612 543740 441640
rect 543424 441600 543430 441612
rect 543734 441600 543740 441612
rect 543792 441600 543798 441652
rect 113082 440240 113088 440292
rect 113140 440280 113146 440292
rect 256694 440280 256700 440292
rect 113140 440252 256700 440280
rect 113140 440240 113146 440252
rect 256694 440240 256700 440252
rect 256752 440240 256758 440292
rect 554130 438880 554136 438932
rect 554188 438920 554194 438932
rect 580166 438920 580172 438932
rect 554188 438892 580172 438920
rect 554188 438880 554194 438892
rect 580166 438880 580172 438892
rect 580224 438880 580230 438932
rect 3142 438812 3148 438864
rect 3200 438852 3206 438864
rect 259914 438852 259920 438864
rect 3200 438824 259920 438852
rect 3200 438812 3206 438824
rect 259914 438812 259920 438824
rect 259972 438812 259978 438864
rect 111702 437452 111708 437504
rect 111760 437492 111766 437504
rect 256694 437492 256700 437504
rect 111760 437464 256700 437492
rect 111760 437452 111766 437464
rect 256694 437452 256700 437464
rect 256752 437452 256758 437504
rect 543366 437384 543372 437436
rect 543424 437384 543430 437436
rect 543274 436636 543280 436688
rect 543332 436676 543338 436688
rect 543384 436676 543412 437384
rect 543332 436648 543412 436676
rect 543332 436636 543338 436648
rect 110322 436092 110328 436144
rect 110380 436132 110386 436144
rect 256694 436132 256700 436144
rect 110380 436104 256700 436132
rect 110380 436092 110386 436104
rect 256694 436092 256700 436104
rect 256752 436092 256758 436144
rect 108942 433304 108948 433356
rect 109000 433344 109006 433356
rect 256694 433344 256700 433356
rect 109000 433316 256700 433344
rect 109000 433304 109006 433316
rect 256694 433304 256700 433316
rect 256752 433304 256758 433356
rect 107562 431944 107568 431996
rect 107620 431984 107626 431996
rect 256694 431984 256700 431996
rect 107620 431956 256700 431984
rect 107620 431944 107626 431956
rect 256694 431944 256700 431956
rect 256752 431944 256758 431996
rect 107470 429156 107476 429208
rect 107528 429196 107534 429208
rect 256694 429196 256700 429208
rect 107528 429168 256700 429196
rect 107528 429156 107534 429168
rect 256694 429156 256700 429168
rect 256752 429156 256758 429208
rect 106182 427796 106188 427848
rect 106240 427836 106246 427848
rect 256694 427836 256700 427848
rect 106240 427808 256700 427836
rect 106240 427796 106246 427808
rect 256694 427796 256700 427808
rect 256752 427796 256758 427848
rect 543274 427796 543280 427848
rect 543332 427796 543338 427848
rect 543292 427768 543320 427796
rect 543366 427768 543372 427780
rect 543292 427740 543372 427768
rect 543366 427728 543372 427740
rect 543424 427728 543430 427780
rect 104802 425076 104808 425128
rect 104860 425116 104866 425128
rect 256694 425116 256700 425128
rect 104860 425088 256700 425116
rect 104860 425076 104866 425088
rect 256694 425076 256700 425088
rect 256752 425076 256758 425128
rect 3234 425008 3240 425060
rect 3292 425048 3298 425060
rect 260006 425048 260012 425060
rect 3292 425020 260012 425048
rect 3292 425008 3298 425020
rect 260006 425008 260012 425020
rect 260064 425008 260070 425060
rect 103422 423648 103428 423700
rect 103480 423688 103486 423700
rect 256694 423688 256700 423700
rect 103480 423660 256700 423688
rect 103480 423648 103486 423660
rect 256694 423648 256700 423660
rect 256752 423648 256758 423700
rect 102042 420928 102048 420980
rect 102100 420968 102106 420980
rect 256694 420968 256700 420980
rect 102100 420940 256700 420968
rect 102100 420928 102106 420940
rect 256694 420928 256700 420940
rect 256752 420928 256758 420980
rect 100662 418140 100668 418192
rect 100720 418180 100726 418192
rect 256694 418180 256700 418192
rect 100720 418152 256700 418180
rect 100720 418140 100726 418152
rect 256694 418140 256700 418152
rect 256752 418140 256758 418192
rect 543366 418140 543372 418192
rect 543424 418140 543430 418192
rect 543384 418044 543412 418140
rect 543458 418044 543464 418056
rect 543384 418016 543464 418044
rect 543458 418004 543464 418016
rect 543516 418004 543522 418056
rect 99282 416780 99288 416832
rect 99340 416820 99346 416832
rect 256694 416820 256700 416832
rect 99340 416792 256700 416820
rect 99340 416780 99346 416792
rect 256694 416780 256700 416792
rect 256752 416780 256758 416832
rect 565170 415420 565176 415472
rect 565228 415460 565234 415472
rect 580166 415460 580172 415472
rect 565228 415432 580172 415460
rect 565228 415420 565234 415432
rect 580166 415420 580172 415432
rect 580224 415420 580230 415472
rect 99190 413992 99196 414044
rect 99248 414032 99254 414044
rect 256694 414032 256700 414044
rect 99248 414004 256700 414032
rect 99248 413992 99254 414004
rect 256694 413992 256700 414004
rect 256752 413992 256758 414044
rect 540606 413516 540612 413568
rect 540664 413556 540670 413568
rect 540790 413556 540796 413568
rect 540664 413528 540796 413556
rect 540664 413516 540670 413528
rect 540790 413516 540796 413528
rect 540848 413516 540854 413568
rect 97902 412632 97908 412684
rect 97960 412672 97966 412684
rect 256694 412672 256700 412684
rect 97960 412644 256700 412672
rect 97960 412632 97966 412644
rect 256694 412632 256700 412644
rect 256752 412632 256758 412684
rect 96522 409844 96528 409896
rect 96580 409884 96586 409896
rect 256694 409884 256700 409896
rect 96580 409856 256700 409884
rect 96580 409844 96586 409856
rect 256694 409844 256700 409856
rect 256752 409844 256758 409896
rect 95142 408484 95148 408536
rect 95200 408524 95206 408536
rect 256694 408524 256700 408536
rect 95200 408496 256700 408524
rect 95200 408484 95206 408496
rect 256694 408484 256700 408496
rect 256752 408484 256758 408536
rect 93762 405696 93768 405748
rect 93820 405736 93826 405748
rect 256694 405736 256700 405748
rect 93820 405708 256700 405736
rect 93820 405696 93826 405708
rect 256694 405696 256700 405708
rect 256752 405696 256758 405748
rect 543458 404472 543464 404524
rect 543516 404472 543522 404524
rect 543476 404388 543504 404472
rect 92382 404336 92388 404388
rect 92440 404376 92446 404388
rect 256694 404376 256700 404388
rect 92440 404348 256700 404376
rect 92440 404336 92446 404348
rect 256694 404336 256700 404348
rect 256752 404336 256758 404388
rect 543458 404336 543464 404388
rect 543516 404336 543522 404388
rect 549990 404336 549996 404388
rect 550048 404376 550054 404388
rect 580166 404376 580172 404388
rect 550048 404348 580172 404376
rect 550048 404336 550054 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 91002 401616 91008 401668
rect 91060 401656 91066 401668
rect 256694 401656 256700 401668
rect 91060 401628 256700 401656
rect 91060 401616 91066 401628
rect 256694 401616 256700 401628
rect 256752 401616 256758 401668
rect 90910 400188 90916 400240
rect 90968 400228 90974 400240
rect 256694 400228 256700 400240
rect 90968 400200 256700 400228
rect 90968 400188 90974 400200
rect 256694 400188 256700 400200
rect 256752 400188 256758 400240
rect 89622 397468 89628 397520
rect 89680 397508 89686 397520
rect 256694 397508 256700 397520
rect 89680 397480 256700 397508
rect 89680 397468 89686 397480
rect 256694 397468 256700 397480
rect 256752 397468 256758 397520
rect 88242 396040 88248 396092
rect 88300 396080 88306 396092
rect 256694 396080 256700 396092
rect 88300 396052 256700 396080
rect 88300 396040 88306 396052
rect 256694 396040 256700 396052
rect 256752 396040 256758 396092
rect 3142 395972 3148 396024
rect 3200 396012 3206 396024
rect 260742 396012 260748 396024
rect 3200 395984 260748 396012
rect 3200 395972 3206 395984
rect 260742 395972 260748 395984
rect 260800 395972 260806 396024
rect 86862 393320 86868 393372
rect 86920 393360 86926 393372
rect 256694 393360 256700 393372
rect 86920 393332 256700 393360
rect 86920 393320 86926 393332
rect 256694 393320 256700 393332
rect 256752 393320 256758 393372
rect 544654 391960 544660 392012
rect 544712 392000 544718 392012
rect 580166 392000 580172 392012
rect 544712 391972 580172 392000
rect 544712 391960 544718 391972
rect 580166 391960 580172 391972
rect 580224 391960 580230 392012
rect 85482 390532 85488 390584
rect 85540 390572 85546 390584
rect 256694 390572 256700 390584
rect 85540 390544 256700 390572
rect 85540 390532 85546 390544
rect 256694 390532 256700 390544
rect 256752 390532 256758 390584
rect 84102 389172 84108 389224
rect 84160 389212 84166 389224
rect 256694 389212 256700 389224
rect 84160 389184 256700 389212
rect 84160 389172 84166 389184
rect 256694 389172 256700 389184
rect 256752 389172 256758 389224
rect 82722 386384 82728 386436
rect 82780 386424 82786 386436
rect 256694 386424 256700 386436
rect 82780 386396 256700 386424
rect 82780 386384 82786 386396
rect 256694 386384 256700 386396
rect 256752 386384 256758 386436
rect 543182 386316 543188 386368
rect 543240 386356 543246 386368
rect 543458 386356 543464 386368
rect 543240 386328 543464 386356
rect 543240 386316 543246 386328
rect 543458 386316 543464 386328
rect 543516 386316 543522 386368
rect 82630 385024 82636 385076
rect 82688 385064 82694 385076
rect 256694 385064 256700 385076
rect 82688 385036 256700 385064
rect 82688 385024 82694 385036
rect 256694 385024 256700 385036
rect 256752 385024 256758 385076
rect 81342 382236 81348 382288
rect 81400 382276 81406 382288
rect 256694 382276 256700 382288
rect 81400 382248 256700 382276
rect 81400 382236 81406 382248
rect 256694 382236 256700 382248
rect 256752 382236 256758 382288
rect 79962 380876 79968 380928
rect 80020 380916 80026 380928
rect 256694 380916 256700 380928
rect 80020 380888 256700 380916
rect 80020 380876 80026 380888
rect 256694 380876 256700 380888
rect 256752 380876 256758 380928
rect 3234 380808 3240 380860
rect 3292 380848 3298 380860
rect 260650 380848 260656 380860
rect 3292 380820 260656 380848
rect 3292 380808 3298 380820
rect 260650 380808 260656 380820
rect 260708 380808 260714 380860
rect 78582 378156 78588 378208
rect 78640 378196 78646 378208
rect 256694 378196 256700 378208
rect 78640 378168 256700 378196
rect 78640 378156 78646 378168
rect 256694 378156 256700 378168
rect 256752 378156 256758 378208
rect 77202 376728 77208 376780
rect 77260 376768 77266 376780
rect 256694 376768 256700 376780
rect 77260 376740 256700 376768
rect 77260 376728 77266 376740
rect 256694 376728 256700 376740
rect 256752 376728 256758 376780
rect 543182 376728 543188 376780
rect 543240 376768 543246 376780
rect 543366 376768 543372 376780
rect 543240 376740 543372 376768
rect 543240 376728 543246 376740
rect 543366 376728 543372 376740
rect 543424 376728 543430 376780
rect 75822 374008 75828 374060
rect 75880 374048 75886 374060
rect 256694 374048 256700 374060
rect 75880 374020 256700 374048
rect 75880 374008 75886 374020
rect 256694 374008 256700 374020
rect 256752 374008 256758 374060
rect 74442 372580 74448 372632
rect 74500 372620 74506 372632
rect 256694 372620 256700 372632
rect 74500 372592 256700 372620
rect 74500 372580 74506 372592
rect 256694 372580 256700 372592
rect 256752 372580 256758 372632
rect 73062 369860 73068 369912
rect 73120 369900 73126 369912
rect 256694 369900 256700 369912
rect 73120 369872 256700 369900
rect 73120 369860 73126 369872
rect 256694 369860 256700 369872
rect 256752 369860 256758 369912
rect 72970 368500 72976 368552
rect 73028 368540 73034 368552
rect 256694 368540 256700 368552
rect 73028 368512 256700 368540
rect 73028 368500 73034 368512
rect 256694 368500 256700 368512
rect 256752 368500 256758 368552
rect 3142 367004 3148 367056
rect 3200 367044 3206 367056
rect 260558 367044 260564 367056
rect 3200 367016 260564 367044
rect 3200 367004 3206 367016
rect 260558 367004 260564 367016
rect 260616 367004 260622 367056
rect 543182 367004 543188 367056
rect 543240 367044 543246 367056
rect 543458 367044 543464 367056
rect 543240 367016 543464 367044
rect 543240 367004 543246 367016
rect 543458 367004 543464 367016
rect 543516 367004 543522 367056
rect 71682 365712 71688 365764
rect 71740 365752 71746 365764
rect 256694 365752 256700 365764
rect 71740 365724 256700 365752
rect 71740 365712 71746 365724
rect 256694 365712 256700 365724
rect 256752 365712 256758 365764
rect 539226 365644 539232 365696
rect 539284 365684 539290 365696
rect 539502 365684 539508 365696
rect 539284 365656 539508 365684
rect 539284 365644 539290 365656
rect 539502 365644 539508 365656
rect 539560 365644 539566 365696
rect 70302 362924 70308 362976
rect 70360 362964 70366 362976
rect 256694 362964 256700 362976
rect 70360 362936 256700 362964
rect 70360 362924 70366 362936
rect 256694 362924 256700 362936
rect 256752 362924 256758 362976
rect 68922 361564 68928 361616
rect 68980 361604 68986 361616
rect 256694 361604 256700 361616
rect 68980 361576 256700 361604
rect 68980 361564 68986 361576
rect 256694 361564 256700 361576
rect 256752 361564 256758 361616
rect 67542 358776 67548 358828
rect 67600 358816 67606 358828
rect 256694 358816 256700 358828
rect 67600 358788 256700 358816
rect 67600 358776 67606 358788
rect 256694 358776 256700 358788
rect 256752 358776 256758 358828
rect 66162 357416 66168 357468
rect 66220 357456 66226 357468
rect 256694 357456 256700 357468
rect 66220 357428 256700 357456
rect 66220 357416 66226 357428
rect 256694 357416 256700 357428
rect 256752 357416 256758 357468
rect 539318 357416 539324 357468
rect 539376 357416 539382 357468
rect 543182 357416 543188 357468
rect 543240 357456 543246 357468
rect 543366 357456 543372 357468
rect 543240 357428 543372 357456
rect 543240 357416 543246 357428
rect 543366 357416 543372 357428
rect 543424 357416 543430 357468
rect 539336 357264 539364 357416
rect 539318 357212 539324 357264
rect 539376 357212 539382 357264
rect 64782 354696 64788 354748
rect 64840 354736 64846 354748
rect 256694 354736 256700 354748
rect 64840 354708 256700 354736
rect 64840 354696 64846 354708
rect 256694 354696 256700 354708
rect 256752 354696 256758 354748
rect 64690 353268 64696 353320
rect 64748 353308 64754 353320
rect 256694 353308 256700 353320
rect 64748 353280 256700 353308
rect 64748 353268 64754 353280
rect 256694 353268 256700 353280
rect 256752 353268 256758 353320
rect 63402 350548 63408 350600
rect 63460 350588 63466 350600
rect 256694 350588 256700 350600
rect 63460 350560 256700 350588
rect 63460 350548 63466 350560
rect 256694 350548 256700 350560
rect 256752 350548 256758 350600
rect 62022 349120 62028 349172
rect 62080 349160 62086 349172
rect 256694 349160 256700 349172
rect 62080 349132 256700 349160
rect 62080 349120 62086 349132
rect 256694 349120 256700 349132
rect 256752 349120 256758 349172
rect 60642 346400 60648 346452
rect 60700 346440 60706 346452
rect 256694 346440 256700 346452
rect 60700 346412 256700 346440
rect 60700 346400 60706 346412
rect 256694 346400 256700 346412
rect 256752 346400 256758 346452
rect 59262 345040 59268 345092
rect 59320 345080 59326 345092
rect 256694 345080 256700 345092
rect 59320 345052 256700 345080
rect 59320 345040 59326 345052
rect 256694 345040 256700 345052
rect 256752 345040 256758 345092
rect 57882 342252 57888 342304
rect 57940 342292 57946 342304
rect 256694 342292 256700 342304
rect 57940 342264 256700 342292
rect 57940 342252 57946 342264
rect 256694 342252 256700 342264
rect 256752 342252 256758 342304
rect 56502 340892 56508 340944
rect 56560 340932 56566 340944
rect 256694 340932 256700 340944
rect 56560 340904 256700 340932
rect 56560 340892 56566 340904
rect 256694 340892 256700 340904
rect 256752 340892 256758 340944
rect 539778 339464 539784 339516
rect 539836 339504 539842 339516
rect 539962 339504 539968 339516
rect 539836 339476 539968 339504
rect 539836 339464 539842 339476
rect 539962 339464 539968 339476
rect 540020 339464 540026 339516
rect 56410 338104 56416 338156
rect 56468 338144 56474 338156
rect 256694 338144 256700 338156
rect 56468 338116 256700 338144
rect 56468 338104 56474 338116
rect 256694 338104 256700 338116
rect 256752 338104 256758 338156
rect 3418 338036 3424 338088
rect 3476 338076 3482 338088
rect 260466 338076 260472 338088
rect 3476 338048 260472 338076
rect 3476 338036 3482 338048
rect 260466 338036 260472 338048
rect 260524 338036 260530 338088
rect 542630 336200 542636 336252
rect 542688 336240 542694 336252
rect 549898 336240 549904 336252
rect 542688 336212 549904 336240
rect 542688 336200 542694 336212
rect 549898 336200 549904 336212
rect 549956 336200 549962 336252
rect 55122 335316 55128 335368
rect 55180 335356 55186 335368
rect 256694 335356 256700 335368
rect 55180 335328 256700 335356
rect 55180 335316 55186 335328
rect 256694 335316 256700 335328
rect 256752 335316 256758 335368
rect 53742 333956 53748 334008
rect 53800 333996 53806 334008
rect 256694 333996 256700 334008
rect 53800 333968 256700 333996
rect 53800 333956 53806 333968
rect 256694 333956 256700 333968
rect 256752 333956 256758 334008
rect 542630 333888 542636 333940
rect 542688 333928 542694 333940
rect 554038 333928 554044 333940
rect 542688 333900 554044 333928
rect 542688 333888 542694 333900
rect 554038 333888 554044 333900
rect 554096 333888 554102 333940
rect 542630 332528 542636 332580
rect 542688 332568 542694 332580
rect 563698 332568 563704 332580
rect 542688 332540 563704 332568
rect 542688 332528 542694 332540
rect 563698 332528 563704 332540
rect 563756 332528 563762 332580
rect 52362 331236 52368 331288
rect 52420 331276 52426 331288
rect 256694 331276 256700 331288
rect 52420 331248 256700 331276
rect 52420 331236 52426 331248
rect 256694 331236 256700 331248
rect 256752 331236 256758 331288
rect 50982 329808 50988 329860
rect 51040 329848 51046 329860
rect 256694 329848 256700 329860
rect 51040 329820 256700 329848
rect 51040 329808 51046 329820
rect 256694 329808 256700 329820
rect 256752 329808 256758 329860
rect 542630 328856 542636 328908
rect 542688 328896 542694 328908
rect 547138 328896 547144 328908
rect 542688 328868 547144 328896
rect 542688 328856 542694 328868
rect 547138 328856 547144 328868
rect 547196 328856 547202 328908
rect 542630 328380 542636 328432
rect 542688 328420 542694 328432
rect 565078 328420 565084 328432
rect 542688 328392 565084 328420
rect 542688 328380 542694 328392
rect 565078 328380 565084 328392
rect 565136 328380 565142 328432
rect 49602 327088 49608 327140
rect 49660 327128 49666 327140
rect 256694 327128 256700 327140
rect 49660 327100 256700 327128
rect 49660 327088 49666 327100
rect 256694 327088 256700 327100
rect 256752 327088 256758 327140
rect 48222 325660 48228 325712
rect 48280 325700 48286 325712
rect 256694 325700 256700 325712
rect 48280 325672 256700 325700
rect 48280 325660 48286 325672
rect 256694 325660 256700 325672
rect 256752 325660 256758 325712
rect 542630 325592 542636 325644
rect 542688 325632 542694 325644
rect 560938 325632 560944 325644
rect 542688 325604 560944 325632
rect 542688 325592 542694 325604
rect 560938 325592 560944 325604
rect 560996 325592 561002 325644
rect 3234 324232 3240 324284
rect 3292 324272 3298 324284
rect 260374 324272 260380 324284
rect 3292 324244 260380 324272
rect 3292 324232 3298 324244
rect 260374 324232 260380 324244
rect 260432 324232 260438 324284
rect 542630 324164 542636 324216
rect 542688 324204 542694 324216
rect 545758 324204 545764 324216
rect 542688 324176 545764 324204
rect 542688 324164 542694 324176
rect 545758 324164 545764 324176
rect 545816 324164 545822 324216
rect 48130 322940 48136 322992
rect 48188 322980 48194 322992
rect 256694 322980 256700 322992
rect 48188 322952 256700 322980
rect 48188 322940 48194 322952
rect 256694 322940 256700 322952
rect 256752 322940 256758 322992
rect 46842 321580 46848 321632
rect 46900 321620 46906 321632
rect 256694 321620 256700 321632
rect 46900 321592 256700 321620
rect 46900 321580 46906 321592
rect 256694 321580 256700 321592
rect 256752 321580 256758 321632
rect 542630 321512 542636 321564
rect 542688 321552 542694 321564
rect 574738 321552 574744 321564
rect 542688 321524 574744 321552
rect 542688 321512 542694 321524
rect 574738 321512 574744 321524
rect 574796 321512 574802 321564
rect 542630 320084 542636 320136
rect 542688 320124 542694 320136
rect 558178 320124 558184 320136
rect 542688 320096 558184 320124
rect 542688 320084 542694 320096
rect 558178 320084 558184 320096
rect 558236 320084 558242 320136
rect 45462 318792 45468 318844
rect 45520 318832 45526 318844
rect 256694 318832 256700 318844
rect 45520 318804 256700 318832
rect 45520 318792 45526 318804
rect 256694 318792 256700 318804
rect 256752 318792 256758 318844
rect 44082 317432 44088 317484
rect 44140 317472 44146 317484
rect 256694 317472 256700 317484
rect 44140 317444 256700 317472
rect 44140 317432 44146 317444
rect 256694 317432 256700 317444
rect 256752 317432 256758 317484
rect 542630 316888 542636 316940
rect 542688 316928 542694 316940
rect 544378 316928 544384 316940
rect 542688 316900 544384 316928
rect 542688 316888 542694 316900
rect 544378 316888 544384 316900
rect 544436 316888 544442 316940
rect 42702 314644 42708 314696
rect 42760 314684 42766 314696
rect 256694 314684 256700 314696
rect 42760 314656 256700 314684
rect 42760 314644 42766 314656
rect 256694 314644 256700 314656
rect 256752 314644 256758 314696
rect 542630 314576 542636 314628
rect 542688 314616 542694 314628
rect 573358 314616 573364 314628
rect 542688 314588 573364 314616
rect 542688 314576 542694 314588
rect 573358 314576 573364 314588
rect 573416 314576 573422 314628
rect 41322 313284 41328 313336
rect 41380 313324 41386 313336
rect 256694 313324 256700 313336
rect 41380 313296 256700 313324
rect 41380 313284 41386 313296
rect 256694 313284 256700 313296
rect 256752 313284 256758 313336
rect 542630 313216 542636 313268
rect 542688 313256 542694 313268
rect 556798 313256 556804 313268
rect 542688 313228 556804 313256
rect 542688 313216 542694 313228
rect 556798 313216 556804 313228
rect 556856 313216 556862 313268
rect 39942 310496 39948 310548
rect 40000 310536 40006 310548
rect 256694 310536 256700 310548
rect 40000 310508 256700 310536
rect 40000 310496 40006 310508
rect 256694 310496 256700 310508
rect 256752 310496 256758 310548
rect 542630 309952 542636 310004
rect 542688 309992 542694 310004
rect 544470 309992 544476 310004
rect 542688 309964 544476 309992
rect 542688 309952 542694 309964
rect 544470 309952 544476 309964
rect 544528 309952 544534 310004
rect 3326 309068 3332 309120
rect 3384 309108 3390 309120
rect 260282 309108 260288 309120
rect 3384 309080 260288 309108
rect 3384 309068 3390 309080
rect 260282 309068 260288 309080
rect 260340 309068 260346 309120
rect 542630 309068 542636 309120
rect 542688 309108 542694 309120
rect 571978 309108 571984 309120
rect 542688 309080 571984 309108
rect 542688 309068 542694 309080
rect 571978 309068 571984 309080
rect 572036 309068 572042 309120
rect 38562 307776 38568 307828
rect 38620 307816 38626 307828
rect 256694 307816 256700 307828
rect 38620 307788 256700 307816
rect 38620 307776 38626 307788
rect 256694 307776 256700 307788
rect 256752 307776 256758 307828
rect 38470 306348 38476 306400
rect 38528 306388 38534 306400
rect 256694 306388 256700 306400
rect 38528 306360 256700 306388
rect 38528 306348 38534 306360
rect 256694 306348 256700 306360
rect 256752 306348 256758 306400
rect 542630 306280 542636 306332
rect 542688 306320 542694 306332
rect 555418 306320 555424 306332
rect 542688 306292 555424 306320
rect 542688 306280 542694 306292
rect 555418 306280 555424 306292
rect 555476 306280 555482 306332
rect 542630 304852 542636 304904
rect 542688 304892 542694 304904
rect 544562 304892 544568 304904
rect 542688 304864 544568 304892
rect 542688 304852 542694 304864
rect 544562 304852 544568 304864
rect 544620 304852 544626 304904
rect 37182 303628 37188 303680
rect 37240 303668 37246 303680
rect 256694 303668 256700 303680
rect 37240 303640 256700 303668
rect 37240 303628 37246 303640
rect 256694 303628 256700 303640
rect 256752 303628 256758 303680
rect 35802 302200 35808 302252
rect 35860 302240 35866 302252
rect 256694 302240 256700 302252
rect 35860 302212 256700 302240
rect 35860 302200 35866 302212
rect 256694 302200 256700 302212
rect 256752 302200 256758 302252
rect 542630 302132 542636 302184
rect 542688 302172 542694 302184
rect 563790 302172 563796 302184
rect 542688 302144 563796 302172
rect 542688 302132 542694 302144
rect 563790 302132 563796 302144
rect 563848 302132 563854 302184
rect 542630 300772 542636 300824
rect 542688 300812 542694 300824
rect 567838 300812 567844 300824
rect 542688 300784 567844 300812
rect 542688 300772 542694 300784
rect 567838 300772 567844 300784
rect 567896 300772 567902 300824
rect 34422 299480 34428 299532
rect 34480 299520 34486 299532
rect 256694 299520 256700 299532
rect 34480 299492 256700 299520
rect 34480 299480 34486 299492
rect 256694 299480 256700 299492
rect 256752 299480 256758 299532
rect 33042 298120 33048 298172
rect 33100 298160 33106 298172
rect 256694 298160 256700 298172
rect 33100 298132 256700 298160
rect 33100 298120 33106 298132
rect 256694 298120 256700 298132
rect 256752 298120 256758 298172
rect 542630 298052 542636 298104
rect 542688 298092 542694 298104
rect 554130 298092 554136 298104
rect 542688 298064 554136 298092
rect 542688 298052 542694 298064
rect 554130 298052 554136 298064
rect 554188 298052 554194 298104
rect 542630 296624 542636 296676
rect 542688 296664 542694 296676
rect 549990 296664 549996 296676
rect 542688 296636 549996 296664
rect 542688 296624 542694 296636
rect 549990 296624 549996 296636
rect 550048 296624 550054 296676
rect 31662 295332 31668 295384
rect 31720 295372 31726 295384
rect 256694 295372 256700 295384
rect 31720 295344 256700 295372
rect 31720 295332 31726 295344
rect 256694 295332 256700 295344
rect 256752 295332 256758 295384
rect 3418 295264 3424 295316
rect 3476 295304 3482 295316
rect 260190 295304 260196 295316
rect 3476 295276 260196 295304
rect 3476 295264 3482 295276
rect 260190 295264 260196 295276
rect 260248 295264 260254 295316
rect 30282 293972 30288 294024
rect 30340 294012 30346 294024
rect 256694 294012 256700 294024
rect 30340 293984 256700 294012
rect 30340 293972 30346 293984
rect 256694 293972 256700 293984
rect 256752 293972 256758 294024
rect 542630 293904 542636 293956
rect 542688 293944 542694 293956
rect 565170 293944 565176 293956
rect 542688 293916 565176 293944
rect 542688 293904 542694 293916
rect 565170 293904 565176 293916
rect 565228 293904 565234 293956
rect 542630 291252 542636 291304
rect 542688 291292 542694 291304
rect 544654 291292 544660 291304
rect 542688 291264 544660 291292
rect 542688 291252 542694 291264
rect 544654 291252 544660 291264
rect 544712 291252 544718 291304
rect 30190 291184 30196 291236
rect 30248 291224 30254 291236
rect 256694 291224 256700 291236
rect 30248 291196 256700 291224
rect 30248 291184 30254 291196
rect 256694 291184 256700 291196
rect 256752 291184 256758 291236
rect 28902 289824 28908 289876
rect 28960 289864 28966 289876
rect 256694 289864 256700 289876
rect 28960 289836 256700 289864
rect 28960 289824 28966 289836
rect 256694 289824 256700 289836
rect 256752 289824 256758 289876
rect 542630 289756 542636 289808
rect 542688 289796 542694 289808
rect 580350 289796 580356 289808
rect 542688 289768 580356 289796
rect 542688 289756 542694 289768
rect 580350 289756 580356 289768
rect 580408 289756 580414 289808
rect 542630 288328 542636 288380
rect 542688 288368 542694 288380
rect 580258 288368 580264 288380
rect 542688 288340 580264 288368
rect 542688 288328 542694 288340
rect 580258 288328 580264 288340
rect 580316 288328 580322 288380
rect 27522 287036 27528 287088
rect 27580 287076 27586 287088
rect 256694 287076 256700 287088
rect 27580 287048 256700 287076
rect 27580 287036 27586 287048
rect 256694 287036 256700 287048
rect 256752 287036 256758 287088
rect 26142 285676 26148 285728
rect 26200 285716 26206 285728
rect 256694 285716 256700 285728
rect 26200 285688 256700 285716
rect 26200 285676 26206 285688
rect 256694 285676 256700 285688
rect 256752 285676 256758 285728
rect 542630 285608 542636 285660
rect 542688 285648 542694 285660
rect 580442 285648 580448 285660
rect 542688 285620 580448 285648
rect 542688 285608 542694 285620
rect 580442 285608 580448 285620
rect 580500 285608 580506 285660
rect 542630 284248 542636 284300
rect 542688 284288 542694 284300
rect 580626 284288 580632 284300
rect 542688 284260 580632 284288
rect 542688 284248 542694 284260
rect 580626 284248 580632 284260
rect 580684 284248 580690 284300
rect 24762 282888 24768 282940
rect 24820 282928 24826 282940
rect 256694 282928 256700 282940
rect 24820 282900 256700 282928
rect 24820 282888 24826 282900
rect 256694 282888 256700 282900
rect 256752 282888 256758 282940
rect 542630 281460 542636 281512
rect 542688 281500 542694 281512
rect 580534 281500 580540 281512
rect 542688 281472 580540 281500
rect 542688 281460 542694 281472
rect 580534 281460 580540 281472
rect 580592 281460 580598 281512
rect 23382 280168 23388 280220
rect 23440 280208 23446 280220
rect 256694 280208 256700 280220
rect 23440 280180 256700 280208
rect 23440 280168 23446 280180
rect 256694 280168 256700 280180
rect 256752 280168 256758 280220
rect 3418 280100 3424 280152
rect 3476 280140 3482 280152
rect 260098 280140 260104 280152
rect 3476 280112 260104 280140
rect 3476 280100 3482 280112
rect 260098 280100 260104 280112
rect 260156 280100 260162 280152
rect 541158 280100 541164 280152
rect 541216 280140 541222 280152
rect 580718 280140 580724 280152
rect 541216 280112 580724 280140
rect 541216 280100 541222 280112
rect 580718 280100 580724 280112
rect 580776 280100 580782 280152
rect 22002 278740 22008 278792
rect 22060 278780 22066 278792
rect 256694 278780 256700 278792
rect 22060 278752 256700 278780
rect 22060 278740 22066 278752
rect 256694 278740 256700 278752
rect 256752 278740 256758 278792
rect 21910 276020 21916 276072
rect 21968 276060 21974 276072
rect 256694 276060 256700 276072
rect 21968 276032 256700 276060
rect 21968 276020 21974 276032
rect 256694 276020 256700 276032
rect 256752 276020 256758 276072
rect 542630 275272 542636 275324
rect 542688 275312 542694 275324
rect 580166 275312 580172 275324
rect 542688 275284 580172 275312
rect 542688 275272 542694 275284
rect 580166 275272 580172 275284
rect 580224 275272 580230 275324
rect 20622 274660 20628 274712
rect 20680 274700 20686 274712
rect 256694 274700 256700 274712
rect 20680 274672 256700 274700
rect 20680 274660 20686 274672
rect 256694 274660 256700 274672
rect 256752 274660 256758 274712
rect 19242 271872 19248 271924
rect 19300 271912 19306 271924
rect 256694 271912 256700 271924
rect 19300 271884 256700 271912
rect 19300 271872 19306 271884
rect 256694 271872 256700 271884
rect 256752 271872 256758 271924
rect 17862 270512 17868 270564
rect 17920 270552 17926 270564
rect 256694 270552 256700 270564
rect 17920 270524 256700 270552
rect 17920 270512 17926 270524
rect 256694 270512 256700 270524
rect 256752 270512 256758 270564
rect 16482 267724 16488 267776
rect 16540 267764 16546 267776
rect 256694 267764 256700 267776
rect 16540 267736 256700 267764
rect 16540 267724 16546 267736
rect 256694 267724 256700 267736
rect 256752 267724 256758 267776
rect 15102 266364 15108 266416
rect 15160 266404 15166 266416
rect 256694 266404 256700 266416
rect 15160 266376 256700 266404
rect 15160 266364 15166 266376
rect 256694 266364 256700 266376
rect 256752 266364 256758 266416
rect 543090 264868 543096 264920
rect 543148 264908 543154 264920
rect 580166 264908 580172 264920
rect 543148 264880 580172 264908
rect 543148 264868 543154 264880
rect 580166 264868 580172 264880
rect 580224 264868 580230 264920
rect 13722 263576 13728 263628
rect 13780 263616 13786 263628
rect 256694 263616 256700 263628
rect 13780 263588 256700 263616
rect 13780 263576 13786 263588
rect 256694 263576 256700 263588
rect 256752 263576 256758 263628
rect 13630 262216 13636 262268
rect 13688 262256 13694 262268
rect 256694 262256 256700 262268
rect 13688 262228 256700 262256
rect 13688 262216 13694 262228
rect 256694 262216 256700 262228
rect 256752 262216 256758 262268
rect 12342 259428 12348 259480
rect 12400 259468 12406 259480
rect 256694 259468 256700 259480
rect 12400 259440 256700 259468
rect 12400 259428 12406 259440
rect 256694 259428 256700 259440
rect 256752 259428 256758 259480
rect 10962 256708 10968 256760
rect 11020 256748 11026 256760
rect 256694 256748 256700 256760
rect 11020 256720 256700 256748
rect 11020 256708 11026 256720
rect 256694 256708 256700 256720
rect 256752 256708 256758 256760
rect 542630 256708 542636 256760
rect 542688 256748 542694 256760
rect 558178 256748 558184 256760
rect 542688 256720 558184 256748
rect 542688 256708 542694 256720
rect 558178 256708 558184 256720
rect 558236 256708 558242 256760
rect 9582 255280 9588 255332
rect 9640 255320 9646 255332
rect 256694 255320 256700 255332
rect 9640 255292 256700 255320
rect 9640 255280 9646 255292
rect 256694 255280 256700 255292
rect 256752 255280 256758 255332
rect 542630 255280 542636 255332
rect 542688 255320 542694 255332
rect 556798 255320 556804 255332
rect 542688 255292 556804 255320
rect 542688 255280 542694 255292
rect 556798 255280 556804 255292
rect 556856 255280 556862 255332
rect 8202 252560 8208 252612
rect 8260 252600 8266 252612
rect 256694 252600 256700 252612
rect 8260 252572 256700 252600
rect 8260 252560 8266 252572
rect 256694 252560 256700 252572
rect 256752 252560 256758 252612
rect 542630 252560 542636 252612
rect 542688 252600 542694 252612
rect 549898 252600 549904 252612
rect 542688 252572 549904 252600
rect 542688 252560 542694 252572
rect 549898 252560 549904 252572
rect 549956 252560 549962 252612
rect 542998 252492 543004 252544
rect 543056 252532 543062 252544
rect 579798 252532 579804 252544
rect 543056 252504 579804 252532
rect 543056 252492 543062 252504
rect 579798 252492 579804 252504
rect 579856 252492 579862 252544
rect 6822 251200 6828 251252
rect 6880 251240 6886 251252
rect 256694 251240 256700 251252
rect 6880 251212 256700 251240
rect 6880 251200 6886 251212
rect 256694 251200 256700 251212
rect 256752 251200 256758 251252
rect 5442 248412 5448 248464
rect 5500 248452 5506 248464
rect 256694 248452 256700 248464
rect 5500 248424 256700 248452
rect 5500 248412 5506 248424
rect 256694 248412 256700 248424
rect 256752 248412 256758 248464
rect 542630 248412 542636 248464
rect 542688 248452 542694 248464
rect 555418 248452 555424 248464
rect 542688 248424 555424 248452
rect 542688 248412 542694 248424
rect 555418 248412 555424 248424
rect 555476 248412 555482 248464
rect 542630 247052 542636 247104
rect 542688 247092 542694 247104
rect 547138 247092 547144 247104
rect 542688 247064 547144 247092
rect 542688 247052 542694 247064
rect 547138 247052 547144 247064
rect 547196 247052 547202 247104
rect 542446 243176 542452 243228
rect 542504 243216 542510 243228
rect 542722 243216 542728 243228
rect 542504 243188 542728 243216
rect 542504 243176 542510 243188
rect 542722 243176 542728 243188
rect 542780 243176 542786 243228
rect 2682 242904 2688 242956
rect 2740 242944 2746 242956
rect 256970 242944 256976 242956
rect 2740 242916 256976 242944
rect 2740 242904 2746 242916
rect 256970 242904 256976 242916
rect 257028 242904 257034 242956
rect 542446 242904 542452 242956
rect 542504 242944 542510 242956
rect 554038 242944 554044 242956
rect 542504 242916 554044 242944
rect 542504 242904 542510 242916
rect 554038 242904 554044 242916
rect 554096 242904 554102 242956
rect 3418 241068 3424 241120
rect 3476 241108 3482 241120
rect 542722 241108 542728 241120
rect 3476 241080 542728 241108
rect 3476 241068 3482 241080
rect 542722 241068 542728 241080
rect 542780 241068 542786 241120
rect 282840 240944 289860 240972
rect 282840 240700 282868 240944
rect 289832 240712 289860 240944
rect 311728 240876 318840 240904
rect 311728 240836 311756 240876
rect 299400 240808 311756 240836
rect 299400 240712 299428 240808
rect 318812 240712 318840 240876
rect 328380 240808 331260 240836
rect 328380 240712 328408 240808
rect 331232 240768 331260 240808
rect 331232 240740 331444 240768
rect 280080 240672 282868 240700
rect 270402 240592 270408 240644
rect 270460 240632 270466 240644
rect 273254 240632 273260 240644
rect 270460 240604 273260 240632
rect 270460 240592 270466 240604
rect 273254 240592 273260 240604
rect 273312 240592 273318 240644
rect 273346 240592 273352 240644
rect 273404 240632 273410 240644
rect 280080 240632 280108 240672
rect 289814 240660 289820 240712
rect 289872 240660 289878 240712
rect 299382 240660 299388 240712
rect 299440 240660 299446 240712
rect 318794 240660 318800 240712
rect 318852 240660 318858 240712
rect 328362 240660 328368 240712
rect 328420 240660 328426 240712
rect 331416 240700 331444 240740
rect 347792 240740 357480 240768
rect 347792 240700 347820 240740
rect 357452 240712 357480 240740
rect 331416 240672 347820 240700
rect 357434 240660 357440 240712
rect 357492 240660 357498 240712
rect 367002 240660 367008 240712
rect 367060 240700 367066 240712
rect 368014 240700 368020 240712
rect 367060 240672 368020 240700
rect 367060 240660 367066 240672
rect 368014 240660 368020 240672
rect 368072 240660 368078 240712
rect 273404 240604 280108 240632
rect 273404 240592 273410 240604
rect 257982 240524 257988 240576
rect 258040 240564 258046 240576
rect 260834 240564 260840 240576
rect 258040 240536 260840 240564
rect 258040 240524 258046 240536
rect 260834 240524 260840 240536
rect 260892 240524 260898 240576
rect 289814 240524 289820 240576
rect 289872 240564 289878 240576
rect 299382 240564 299388 240576
rect 289872 240536 299388 240564
rect 289872 240524 289878 240536
rect 299382 240524 299388 240536
rect 299440 240524 299446 240576
rect 318794 240524 318800 240576
rect 318852 240564 318858 240576
rect 328362 240564 328368 240576
rect 318852 240536 328368 240564
rect 318852 240524 318858 240536
rect 328362 240524 328368 240536
rect 328420 240524 328426 240576
rect 260834 240388 260840 240440
rect 260892 240428 260898 240440
rect 261110 240428 261116 240440
rect 260892 240400 261116 240428
rect 260892 240388 260898 240400
rect 261110 240388 261116 240400
rect 261168 240428 261174 240440
rect 270402 240428 270408 240440
rect 261168 240400 270408 240428
rect 261168 240388 261174 240400
rect 270402 240388 270408 240400
rect 270460 240388 270466 240440
rect 1302 240116 1308 240168
rect 1360 240156 1366 240168
rect 257982 240156 257988 240168
rect 1360 240128 257988 240156
rect 1360 240116 1366 240128
rect 257982 240116 257988 240128
rect 258040 240116 258046 240168
rect 542446 240116 542452 240168
rect 542504 240156 542510 240168
rect 545758 240156 545764 240168
rect 542504 240128 545764 240156
rect 542504 240116 542510 240128
rect 545758 240116 545764 240128
rect 545816 240116 545822 240168
rect 368014 240048 368020 240100
rect 368072 240088 368078 240100
rect 373258 240088 373264 240100
rect 368072 240060 373264 240088
rect 368072 240048 368078 240060
rect 373258 240048 373264 240060
rect 373316 240048 373322 240100
rect 331122 238688 331128 238740
rect 331180 238728 331186 238740
rect 340782 238728 340788 238740
rect 331180 238700 340788 238728
rect 331180 238688 331186 238700
rect 340782 238688 340788 238700
rect 340840 238688 340846 238740
rect 433242 238688 433248 238740
rect 433300 238728 433306 238740
rect 449158 238728 449164 238740
rect 433300 238700 449164 238728
rect 433300 238688 433306 238700
rect 449158 238688 449164 238700
rect 449216 238688 449222 238740
rect 464062 238688 464068 238740
rect 464120 238728 464126 238740
rect 477034 238728 477040 238740
rect 464120 238700 477040 238728
rect 464120 238688 464126 238700
rect 477034 238688 477040 238700
rect 477092 238688 477098 238740
rect 477218 238688 477224 238740
rect 477276 238728 477282 238740
rect 497458 238728 497464 238740
rect 477276 238700 497464 238728
rect 477276 238688 477282 238700
rect 497458 238688 497464 238700
rect 497516 238688 497522 238740
rect 325326 238620 325332 238672
rect 325384 238660 325390 238672
rect 336734 238660 336740 238672
rect 325384 238632 336740 238660
rect 325384 238620 325390 238632
rect 336734 238620 336740 238632
rect 336792 238620 336798 238672
rect 391198 238620 391204 238672
rect 391256 238660 391262 238672
rect 404998 238660 405004 238672
rect 391256 238632 405004 238660
rect 391256 238620 391262 238632
rect 404998 238620 405004 238632
rect 405056 238620 405062 238672
rect 430666 238620 430672 238672
rect 430724 238660 430730 238672
rect 450538 238660 450544 238672
rect 430724 238632 450544 238660
rect 430724 238620 430730 238632
rect 450538 238620 450544 238632
rect 450596 238620 450602 238672
rect 458910 238620 458916 238672
rect 458968 238660 458974 238672
rect 479518 238660 479524 238672
rect 458968 238632 479524 238660
rect 458968 238620 458974 238632
rect 479518 238620 479524 238632
rect 479576 238620 479582 238672
rect 263686 238552 263692 238604
rect 263744 238592 263750 238604
rect 297818 238592 297824 238604
rect 263744 238564 297824 238592
rect 263744 238552 263750 238564
rect 297818 238552 297824 238564
rect 297876 238552 297882 238604
rect 329742 238552 329748 238604
rect 329800 238592 329806 238604
rect 343358 238592 343364 238604
rect 329800 238564 343364 238592
rect 329800 238552 329806 238564
rect 343358 238552 343364 238564
rect 343416 238552 343422 238604
rect 388438 238552 388444 238604
rect 388496 238592 388502 238604
rect 402422 238592 402428 238604
rect 388496 238564 402428 238592
rect 388496 238552 388502 238564
rect 402422 238552 402428 238564
rect 402480 238552 402486 238604
rect 428090 238552 428096 238604
rect 428148 238592 428154 238604
rect 451918 238592 451924 238604
rect 428148 238564 451924 238592
rect 428148 238552 428154 238564
rect 451918 238552 451924 238564
rect 451976 238552 451982 238604
rect 463602 238552 463608 238604
rect 463660 238592 463666 238604
rect 505186 238592 505192 238604
rect 463660 238564 505192 238592
rect 463660 238552 463666 238564
rect 505186 238552 505192 238564
rect 505244 238552 505250 238604
rect 261202 238484 261208 238536
rect 261260 238524 261266 238536
rect 297358 238524 297364 238536
rect 261260 238496 297364 238524
rect 261260 238484 261266 238496
rect 297358 238484 297364 238496
rect 297416 238484 297422 238536
rect 328362 238484 328368 238536
rect 328420 238524 328426 238536
rect 345934 238524 345940 238536
rect 328420 238496 345940 238524
rect 328420 238484 328426 238496
rect 345934 238484 345940 238496
rect 345992 238484 345998 238536
rect 380342 238484 380348 238536
rect 380400 238524 380406 238536
rect 394694 238524 394700 238536
rect 380400 238496 394700 238524
rect 380400 238484 380406 238496
rect 394694 238484 394700 238496
rect 394752 238484 394758 238536
rect 420362 238484 420368 238536
rect 420420 238524 420426 238536
rect 456242 238524 456248 238536
rect 420420 238496 456248 238524
rect 420420 238484 420426 238496
rect 456242 238484 456248 238496
rect 456300 238484 456306 238536
rect 460842 238484 460848 238536
rect 460900 238524 460906 238536
rect 512822 238524 512828 238536
rect 460900 238496 512828 238524
rect 460900 238484 460906 238496
rect 512822 238484 512828 238496
rect 512880 238484 512886 238536
rect 297082 238416 297088 238468
rect 297140 238456 297146 238468
rect 347038 238456 347044 238468
rect 297140 238428 347044 238456
rect 297140 238416 297146 238428
rect 347038 238416 347044 238428
rect 347096 238416 347102 238468
rect 380250 238416 380256 238468
rect 380308 238456 380314 238468
rect 397270 238456 397276 238468
rect 380308 238428 397276 238456
rect 380308 238416 380314 238428
rect 397270 238416 397276 238428
rect 397328 238416 397334 238468
rect 417786 238416 417792 238468
rect 417844 238456 417850 238468
rect 456058 238456 456064 238468
rect 417844 238428 456064 238456
rect 417844 238416 417850 238428
rect 456058 238416 456064 238428
rect 456116 238416 456122 238468
rect 458082 238416 458088 238468
rect 458140 238456 458146 238468
rect 517974 238456 517980 238468
rect 458140 238428 517980 238456
rect 458140 238416 458146 238428
rect 517974 238416 517980 238428
rect 518032 238416 518038 238468
rect 294506 238348 294512 238400
rect 294564 238388 294570 238400
rect 344278 238388 344284 238400
rect 294564 238360 344284 238388
rect 294564 238348 294570 238360
rect 344278 238348 344284 238360
rect 344336 238348 344342 238400
rect 371142 238348 371148 238400
rect 371200 238388 371206 238400
rect 389542 238388 389548 238400
rect 371200 238360 389548 238388
rect 371200 238348 371206 238360
rect 389542 238348 389548 238360
rect 389600 238348 389606 238400
rect 393958 238348 393964 238400
rect 394016 238388 394022 238400
rect 407574 238388 407580 238400
rect 394016 238360 407580 238388
rect 394016 238348 394022 238360
rect 407574 238348 407580 238360
rect 407632 238348 407638 238400
rect 422938 238348 422944 238400
rect 422996 238388 423002 238400
rect 454678 238388 454684 238400
rect 422996 238360 454684 238388
rect 422996 238348 423002 238360
rect 454678 238348 454684 238360
rect 454736 238348 454742 238400
rect 455230 238348 455236 238400
rect 455288 238388 455294 238400
rect 523126 238388 523132 238400
rect 455288 238360 523132 238388
rect 455288 238348 455294 238360
rect 523126 238348 523132 238360
rect 523184 238348 523190 238400
rect 289446 238280 289452 238332
rect 289504 238320 289510 238332
rect 341518 238320 341524 238332
rect 289504 238292 341524 238320
rect 289504 238280 289510 238292
rect 341518 238280 341524 238292
rect 341576 238280 341582 238332
rect 380434 238280 380440 238332
rect 380492 238320 380498 238332
rect 415302 238320 415308 238332
rect 380492 238292 415308 238320
rect 380492 238280 380498 238292
rect 415302 238280 415308 238292
rect 415360 238280 415366 238332
rect 425514 238280 425520 238332
rect 425572 238320 425578 238332
rect 453298 238320 453304 238332
rect 425572 238292 453304 238320
rect 425572 238280 425578 238292
rect 453298 238280 453304 238292
rect 453356 238280 453362 238332
rect 453942 238280 453948 238332
rect 454000 238320 454006 238332
rect 528278 238320 528284 238332
rect 454000 238292 528284 238320
rect 454000 238280 454006 238292
rect 528278 238280 528284 238292
rect 528336 238280 528342 238332
rect 284294 238212 284300 238264
rect 284352 238252 284358 238264
rect 338758 238252 338764 238264
rect 284352 238224 338764 238252
rect 284352 238212 284358 238224
rect 338758 238212 338764 238224
rect 338816 238212 338822 238264
rect 384482 238212 384488 238264
rect 384540 238252 384546 238264
rect 447778 238252 447784 238264
rect 384540 238224 447784 238252
rect 384540 238212 384546 238224
rect 447778 238212 447784 238224
rect 447836 238212 447842 238264
rect 451182 238212 451188 238264
rect 451240 238252 451246 238264
rect 533430 238252 533436 238264
rect 451240 238224 533436 238252
rect 451240 238212 451246 238224
rect 533430 238212 533436 238224
rect 533488 238212 533494 238264
rect 286870 238144 286876 238196
rect 286928 238184 286934 238196
rect 340138 238184 340144 238196
rect 286928 238156 340144 238184
rect 286928 238144 286934 238156
rect 340138 238144 340144 238156
rect 340196 238144 340202 238196
rect 380158 238144 380164 238196
rect 380216 238184 380222 238196
rect 399846 238184 399852 238196
rect 380216 238156 399852 238184
rect 380216 238144 380222 238156
rect 399846 238144 399852 238156
rect 399904 238144 399910 238196
rect 412726 238144 412732 238196
rect 412784 238184 412790 238196
rect 496354 238184 496360 238196
rect 412784 238156 496360 238184
rect 412784 238144 412790 238156
rect 496354 238144 496360 238156
rect 496412 238144 496418 238196
rect 292022 238076 292028 238128
rect 292080 238116 292086 238128
rect 345750 238116 345756 238128
rect 292080 238088 345756 238116
rect 292080 238076 292086 238088
rect 345750 238076 345756 238088
rect 345808 238076 345814 238128
rect 356146 238076 356152 238128
rect 356204 238116 356210 238128
rect 478230 238116 478236 238128
rect 356204 238088 478236 238116
rect 356204 238076 356210 238088
rect 478230 238076 478236 238088
rect 478288 238076 478294 238128
rect 266262 238008 266268 238060
rect 266320 238048 266326 238060
rect 345658 238048 345664 238060
rect 266320 238020 345664 238048
rect 266320 238008 266326 238020
rect 345658 238008 345664 238020
rect 345716 238008 345722 238060
rect 353662 238008 353668 238060
rect 353720 238048 353726 238060
rect 477126 238048 477132 238060
rect 353720 238020 477132 238048
rect 353720 238008 353726 238020
rect 477126 238008 477132 238020
rect 477184 238008 477190 238060
rect 478322 238008 478328 238060
rect 478380 238048 478386 238060
rect 500034 238048 500040 238060
rect 478380 238020 500040 238048
rect 478380 238008 478386 238020
rect 500034 238008 500040 238020
rect 500092 238008 500098 238060
rect 435818 237940 435824 237992
rect 435876 237980 435882 237992
rect 447870 237980 447876 237992
rect 435876 237952 447876 237980
rect 435876 237940 435882 237952
rect 447870 237940 447876 237952
rect 447928 237940 447934 237992
rect 471882 237940 471888 237992
rect 471940 237980 471946 237992
rect 487154 237980 487160 237992
rect 471940 237952 487160 237980
rect 471940 237940 471946 237952
rect 487154 237940 487160 237952
rect 487212 237940 487218 237992
rect 473262 237872 473268 237924
rect 473320 237912 473326 237924
rect 484578 237912 484584 237924
rect 473320 237884 484584 237912
rect 473320 237872 473326 237884
rect 484578 237872 484584 237884
rect 484636 237872 484642 237924
rect 466638 237804 466644 237856
rect 466696 237844 466702 237856
rect 476758 237844 476764 237856
rect 466696 237816 476764 237844
rect 466696 237804 466702 237816
rect 476758 237804 476764 237816
rect 476816 237804 476822 237856
rect 469214 237736 469220 237788
rect 469272 237776 469278 237788
rect 478138 237776 478144 237788
rect 469272 237748 478144 237776
rect 469272 237736 469278 237748
rect 478138 237736 478144 237748
rect 478196 237736 478202 237788
rect 471790 237600 471796 237652
rect 471848 237640 471854 237652
rect 477586 237640 477592 237652
rect 471848 237612 477592 237640
rect 471848 237600 471854 237612
rect 477586 237600 477592 237612
rect 477644 237600 477650 237652
rect 332502 237532 332508 237584
rect 332560 237572 332566 237584
rect 338206 237572 338212 237584
rect 332560 237544 338212 237572
rect 332560 237532 332566 237544
rect 338206 237532 338212 237544
rect 338264 237532 338270 237584
rect 476022 237532 476028 237584
rect 476080 237572 476086 237584
rect 479426 237572 479432 237584
rect 476080 237544 479432 237572
rect 476080 237532 476086 237544
rect 479426 237532 479432 237544
rect 479484 237532 479490 237584
rect 333882 237464 333888 237516
rect 333940 237504 333946 237516
rect 335630 237504 335636 237516
rect 333940 237476 335636 237504
rect 333940 237464 333946 237476
rect 335630 237464 335636 237476
rect 335688 237464 335694 237516
rect 476942 237464 476948 237516
rect 477000 237504 477006 237516
rect 482002 237504 482008 237516
rect 477000 237476 482008 237504
rect 477000 237464 477006 237476
rect 482002 237464 482008 237476
rect 482060 237464 482066 237516
rect 276566 237396 276572 237448
rect 276624 237436 276630 237448
rect 277302 237436 277308 237448
rect 276624 237408 277308 237436
rect 276624 237396 276630 237408
rect 277302 237396 277308 237408
rect 277360 237396 277366 237448
rect 279142 237396 279148 237448
rect 279200 237436 279206 237448
rect 280062 237436 280068 237448
rect 279200 237408 280068 237436
rect 279200 237396 279206 237408
rect 280062 237396 280068 237408
rect 280120 237396 280126 237448
rect 281718 237396 281724 237448
rect 281776 237436 281782 237448
rect 282822 237436 282828 237448
rect 281776 237408 282828 237436
rect 281776 237396 281782 237408
rect 282822 237396 282828 237408
rect 282880 237396 282886 237448
rect 299658 237396 299664 237448
rect 299716 237436 299722 237448
rect 300762 237436 300768 237448
rect 299716 237408 300768 237436
rect 299716 237396 299722 237408
rect 300762 237396 300768 237408
rect 300820 237396 300826 237448
rect 302234 237396 302240 237448
rect 302292 237436 302298 237448
rect 303522 237436 303528 237448
rect 302292 237408 303528 237436
rect 302292 237396 302298 237408
rect 303522 237396 303528 237408
rect 303580 237396 303586 237448
rect 315114 237396 315120 237448
rect 315172 237436 315178 237448
rect 315942 237436 315948 237448
rect 315172 237408 315948 237436
rect 315172 237396 315178 237408
rect 315942 237396 315948 237408
rect 316000 237396 316006 237448
rect 317690 237396 317696 237448
rect 317748 237436 317754 237448
rect 318702 237436 318708 237448
rect 317748 237408 318708 237436
rect 317748 237396 317754 237408
rect 318702 237396 318708 237408
rect 318760 237396 318766 237448
rect 320266 237396 320272 237448
rect 320324 237436 320330 237448
rect 321462 237436 321468 237448
rect 320324 237408 321468 237436
rect 320324 237396 320330 237408
rect 321462 237396 321468 237408
rect 321520 237396 321526 237448
rect 333054 237396 333060 237448
rect 333112 237436 333118 237448
rect 333974 237436 333980 237448
rect 333112 237408 333980 237436
rect 333112 237396 333118 237408
rect 333974 237396 333980 237408
rect 334032 237396 334038 237448
rect 351086 237396 351092 237448
rect 351144 237436 351150 237448
rect 351822 237436 351828 237448
rect 351144 237408 351828 237436
rect 351144 237396 351150 237408
rect 351822 237396 351828 237408
rect 351880 237396 351886 237448
rect 361298 237396 361304 237448
rect 361356 237436 361362 237448
rect 362218 237436 362224 237448
rect 361356 237408 362224 237436
rect 361356 237396 361362 237408
rect 362218 237396 362224 237408
rect 362276 237396 362282 237448
rect 371602 237396 371608 237448
rect 371660 237436 371666 237448
rect 372522 237436 372528 237448
rect 371660 237408 372528 237436
rect 371660 237396 371666 237408
rect 372522 237396 372528 237408
rect 372580 237396 372586 237448
rect 374178 237396 374184 237448
rect 374236 237436 374242 237448
rect 375282 237436 375288 237448
rect 374236 237408 375288 237436
rect 374236 237396 374242 237408
rect 375282 237396 375288 237408
rect 375340 237396 375346 237448
rect 376754 237396 376760 237448
rect 376812 237436 376818 237448
rect 378042 237436 378048 237448
rect 376812 237408 378048 237436
rect 376812 237396 376818 237408
rect 378042 237396 378048 237408
rect 378100 237396 378106 237448
rect 386966 237396 386972 237448
rect 387024 237436 387030 237448
rect 387702 237436 387708 237448
rect 387024 237408 387708 237436
rect 387024 237396 387030 237408
rect 387702 237396 387708 237408
rect 387760 237396 387766 237448
rect 461486 237396 461492 237448
rect 461544 237436 461550 237448
rect 462222 237436 462228 237448
rect 461544 237408 462228 237436
rect 461544 237396 461550 237408
rect 462222 237396 462228 237408
rect 462280 237396 462286 237448
rect 474366 237396 474372 237448
rect 474424 237436 474430 237448
rect 477494 237436 477500 237448
rect 474424 237408 477500 237436
rect 474424 237396 474430 237408
rect 477494 237396 477500 237408
rect 477552 237396 477558 237448
rect 3418 237328 3424 237380
rect 3476 237368 3482 237380
rect 540422 237368 540428 237380
rect 3476 237340 540428 237368
rect 3476 237328 3482 237340
rect 540422 237328 540428 237340
rect 540480 237328 540486 237380
rect 542170 234608 542176 234660
rect 542228 234648 542234 234660
rect 542814 234648 542820 234660
rect 542228 234620 542820 234648
rect 542228 234608 542234 234620
rect 542814 234608 542820 234620
rect 542872 234608 542878 234660
rect 542630 231752 542636 231804
rect 542688 231792 542694 231804
rect 542814 231792 542820 231804
rect 542688 231764 542820 231792
rect 542688 231752 542694 231764
rect 542814 231752 542820 231764
rect 542872 231752 542878 231804
rect 543550 229032 543556 229084
rect 543608 229072 543614 229084
rect 580166 229072 580172 229084
rect 543608 229044 580172 229072
rect 543608 229032 543614 229044
rect 580166 229032 580172 229044
rect 580224 229032 580230 229084
rect 3142 223524 3148 223576
rect 3200 223564 3206 223576
rect 542354 223564 542360 223576
rect 3200 223536 542360 223564
rect 3200 223524 3206 223536
rect 542354 223524 542360 223536
rect 542412 223524 542418 223576
rect 542630 222164 542636 222216
rect 542688 222204 542694 222216
rect 542906 222204 542912 222216
rect 542688 222176 542912 222204
rect 542688 222164 542694 222176
rect 542906 222164 542912 222176
rect 542964 222164 542970 222216
rect 543458 217948 543464 218000
rect 543516 217988 543522 218000
rect 580166 217988 580172 218000
rect 543516 217960 580172 217988
rect 543516 217948 543522 217960
rect 580166 217948 580172 217960
rect 580224 217948 580230 218000
rect 542906 215404 542912 215416
rect 542832 215376 542912 215404
rect 542832 215280 542860 215376
rect 542906 215364 542912 215376
rect 542964 215364 542970 215416
rect 542814 215228 542820 215280
rect 542872 215228 542878 215280
rect 542722 212440 542728 212492
rect 542780 212480 542786 212492
rect 542814 212480 542820 212492
rect 542780 212452 542820 212480
rect 542780 212440 542786 212452
rect 542814 212440 542820 212452
rect 542872 212440 542878 212492
rect 3418 208292 3424 208344
rect 3476 208332 3482 208344
rect 541618 208332 541624 208344
rect 3476 208304 541624 208332
rect 3476 208292 3482 208304
rect 541618 208292 541624 208304
rect 541676 208292 541682 208344
rect 543366 205572 543372 205624
rect 543424 205612 543430 205624
rect 579798 205612 579804 205624
rect 543424 205584 579804 205612
rect 543424 205572 543430 205584
rect 579798 205572 579804 205584
rect 579856 205572 579862 205624
rect 470502 205164 470508 205216
rect 470560 205204 470566 205216
rect 488534 205204 488540 205216
rect 470560 205176 488540 205204
rect 470560 205164 470566 205176
rect 488534 205164 488540 205176
rect 488592 205164 488598 205216
rect 470410 205028 470416 205080
rect 470468 205068 470474 205080
rect 491294 205068 491300 205080
rect 470468 205040 491300 205068
rect 470468 205028 470474 205040
rect 491294 205028 491300 205040
rect 491352 205028 491358 205080
rect 469122 204960 469128 205012
rect 469180 205000 469186 205012
rect 494054 205000 494060 205012
rect 469180 204972 494060 205000
rect 469180 204960 469186 204972
rect 494054 204960 494060 204972
rect 494112 204960 494118 205012
rect 369762 204892 369768 204944
rect 369820 204932 369826 204944
rect 490190 204932 490196 204944
rect 369820 204904 490196 204932
rect 369820 204892 369826 204904
rect 490190 204892 490196 204904
rect 490248 204892 490254 204944
rect 473814 204416 473820 204468
rect 473872 204456 473878 204468
rect 477218 204456 477224 204468
rect 473872 204428 477224 204456
rect 473872 204416 473878 204428
rect 477218 204416 477224 204428
rect 477276 204416 477282 204468
rect 345382 204320 345388 204332
rect 342916 204292 345388 204320
rect 331030 204212 331036 204264
rect 331088 204252 331094 204264
rect 334066 204252 334072 204264
rect 331088 204224 334072 204252
rect 331088 204212 331094 204224
rect 334066 204212 334072 204224
rect 334124 204212 334130 204264
rect 336366 204212 336372 204264
rect 336424 204252 336430 204264
rect 342162 204252 342168 204264
rect 336424 204224 342168 204252
rect 336424 204212 336430 204224
rect 342162 204212 342168 204224
rect 342220 204212 342226 204264
rect 282822 204144 282828 204196
rect 282880 204184 282886 204196
rect 342916 204184 342944 204292
rect 345382 204280 345388 204292
rect 345440 204280 345446 204332
rect 345290 204212 345296 204264
rect 345348 204252 345354 204264
rect 349154 204252 349160 204264
rect 345348 204224 349160 204252
rect 345348 204212 345354 204224
rect 349154 204212 349160 204224
rect 349212 204212 349218 204264
rect 364242 204212 364248 204264
rect 364300 204252 364306 204264
rect 365714 204252 365720 204264
rect 364300 204224 365720 204252
rect 364300 204212 364306 204224
rect 365714 204212 365720 204224
rect 365772 204212 365778 204264
rect 456058 204212 456064 204264
rect 456116 204252 456122 204264
rect 456610 204252 456616 204264
rect 456116 204224 456616 204252
rect 456116 204212 456122 204224
rect 456610 204212 456616 204224
rect 456668 204252 456674 204264
rect 465074 204252 465080 204264
rect 456668 204224 465080 204252
rect 456668 204212 456674 204224
rect 465074 204212 465080 204224
rect 465132 204212 465138 204264
rect 477034 204212 477040 204264
rect 477092 204252 477098 204264
rect 481634 204252 481640 204264
rect 477092 204224 481640 204252
rect 477092 204212 477098 204224
rect 481634 204212 481640 204224
rect 481692 204212 481698 204264
rect 282880 204156 342944 204184
rect 282880 204144 282886 204156
rect 345382 204144 345388 204196
rect 345440 204184 345446 204196
rect 357434 204184 357440 204196
rect 345440 204156 357440 204184
rect 345440 204144 345446 204156
rect 357434 204144 357440 204156
rect 357492 204144 357498 204196
rect 362218 204144 362224 204196
rect 362276 204184 362282 204196
rect 367094 204184 367100 204196
rect 362276 204156 367100 204184
rect 362276 204144 362282 204156
rect 367094 204144 367100 204156
rect 367152 204144 367158 204196
rect 467742 204144 467748 204196
rect 467800 204184 467806 204196
rect 473814 204184 473820 204196
rect 467800 204156 473820 204184
rect 467800 204144 467806 204156
rect 473814 204144 473820 204156
rect 473872 204144 473878 204196
rect 478230 204144 478236 204196
rect 478288 204184 478294 204196
rect 485774 204184 485780 204196
rect 478288 204156 485780 204184
rect 478288 204144 478294 204156
rect 485774 204144 485780 204156
rect 485832 204144 485838 204196
rect 300762 204076 300768 204128
rect 300820 204116 300826 204128
rect 345290 204116 345296 204128
rect 300820 204088 345296 204116
rect 300820 204076 300826 204088
rect 345290 204076 345296 204088
rect 345348 204076 345354 204128
rect 345750 204076 345756 204128
rect 345808 204116 345814 204128
rect 351914 204116 351920 204128
rect 345808 204088 351920 204116
rect 345808 204076 345814 204088
rect 351914 204076 351920 204088
rect 351972 204076 351978 204128
rect 449802 204076 449808 204128
rect 449860 204116 449866 204128
rect 535454 204116 535460 204128
rect 449860 204088 535460 204116
rect 449860 204076 449866 204088
rect 535454 204076 535460 204088
rect 535512 204076 535518 204128
rect 303522 204008 303528 204060
rect 303580 204048 303586 204060
rect 343818 204048 343824 204060
rect 303580 204020 343824 204048
rect 303580 204008 303586 204020
rect 343818 204008 343824 204020
rect 343876 204008 343882 204060
rect 346394 204048 346400 204060
rect 343928 204020 346400 204048
rect 304902 203940 304908 203992
rect 304960 203980 304966 203992
rect 343928 203980 343956 204020
rect 346394 204008 346400 204020
rect 346452 204008 346458 204060
rect 349246 204008 349252 204060
rect 349304 204048 349310 204060
rect 357526 204048 357532 204060
rect 349304 204020 357532 204048
rect 349304 204008 349310 204020
rect 357526 204008 357532 204020
rect 357584 204008 357590 204060
rect 360010 204008 360016 204060
rect 360068 204048 360074 204060
rect 448514 204048 448520 204060
rect 360068 204020 448520 204048
rect 360068 204008 360074 204020
rect 448514 204008 448520 204020
rect 448572 204008 448578 204060
rect 449158 204008 449164 204060
rect 449216 204048 449222 204060
rect 459002 204048 459008 204060
rect 449216 204020 459008 204048
rect 449216 204008 449222 204020
rect 459002 204008 459008 204020
rect 459060 204048 459066 204060
rect 465166 204048 465172 204060
rect 459060 204020 465172 204048
rect 459060 204008 459066 204020
rect 465166 204008 465172 204020
rect 465224 204008 465230 204060
rect 466546 204008 466552 204060
rect 466604 204048 466610 204060
rect 474182 204048 474188 204060
rect 466604 204020 474188 204048
rect 466604 204008 466610 204020
rect 474182 204008 474188 204020
rect 474240 204048 474246 204060
rect 476666 204048 476672 204060
rect 474240 204020 476672 204048
rect 474240 204008 474246 204020
rect 476666 204008 476672 204020
rect 476724 204008 476730 204060
rect 476758 204008 476764 204060
rect 476816 204048 476822 204060
rect 480438 204048 480444 204060
rect 476816 204020 480444 204048
rect 476816 204008 476822 204020
rect 480438 204008 480444 204020
rect 480496 204008 480502 204060
rect 304960 203952 343956 203980
rect 304960 203940 304966 203952
rect 344278 203940 344284 203992
rect 344336 203980 344342 203992
rect 351086 203980 351092 203992
rect 344336 203952 351092 203980
rect 344336 203940 344342 203952
rect 351086 203940 351092 203952
rect 351144 203940 351150 203992
rect 351730 203940 351736 203992
rect 351788 203980 351794 203992
rect 361298 203980 361304 203992
rect 351788 203952 361304 203980
rect 351788 203940 351794 203952
rect 361298 203940 361304 203952
rect 361356 203980 361362 203992
rect 445754 203980 445760 203992
rect 361356 203952 445760 203980
rect 361356 203940 361362 203952
rect 445754 203940 445760 203952
rect 445812 203940 445818 203992
rect 459462 203940 459468 203992
rect 459520 203980 459526 203992
rect 514754 203980 514760 203992
rect 459520 203952 514760 203980
rect 459520 203940 459526 203952
rect 514754 203940 514760 203952
rect 514812 203940 514818 203992
rect 307662 203872 307668 203924
rect 307720 203912 307726 203924
rect 345014 203912 345020 203924
rect 307720 203884 345020 203912
rect 307720 203872 307726 203884
rect 345014 203872 345020 203884
rect 345072 203872 345078 203924
rect 345658 203872 345664 203924
rect 345716 203912 345722 203924
rect 364334 203912 364340 203924
rect 345716 203884 364340 203912
rect 345716 203872 345722 203884
rect 364334 203872 364340 203884
rect 364392 203872 364398 203924
rect 450538 203872 450544 203924
rect 450596 203912 450602 203924
rect 460566 203912 460572 203924
rect 450596 203884 460572 203912
rect 450596 203872 450602 203884
rect 460566 203872 460572 203884
rect 460624 203872 460630 203924
rect 462130 203872 462136 203924
rect 462188 203912 462194 203924
rect 509234 203912 509240 203924
rect 462188 203884 509240 203912
rect 462188 203872 462194 203884
rect 509234 203872 509240 203884
rect 509292 203872 509298 203924
rect 310422 203804 310428 203856
rect 310480 203844 310486 203856
rect 343634 203844 343640 203856
rect 310480 203816 343640 203844
rect 310480 203804 310486 203816
rect 343634 203804 343640 203816
rect 343692 203804 343698 203856
rect 343818 203804 343824 203856
rect 343876 203844 343882 203856
rect 347774 203844 347780 203856
rect 343876 203816 347780 203844
rect 343876 203804 343882 203816
rect 347774 203804 347780 203816
rect 347832 203804 347838 203856
rect 363506 203844 363512 203856
rect 354968 203816 363512 203844
rect 313182 203736 313188 203788
rect 313240 203776 313246 203788
rect 332318 203776 332324 203788
rect 313240 203748 332324 203776
rect 313240 203736 313246 203748
rect 332318 203736 332324 203748
rect 332376 203736 332382 203788
rect 332410 203736 332416 203788
rect 332468 203776 332474 203788
rect 336366 203776 336372 203788
rect 332468 203748 336372 203776
rect 332468 203736 332474 203748
rect 336366 203736 336372 203748
rect 336424 203736 336430 203788
rect 336458 203736 336464 203788
rect 336516 203776 336522 203788
rect 340046 203776 340052 203788
rect 336516 203748 340052 203776
rect 336516 203736 336522 203748
rect 340046 203736 340052 203748
rect 340104 203736 340110 203788
rect 340138 203736 340144 203788
rect 340196 203776 340202 203788
rect 354674 203776 354680 203788
rect 340196 203748 354680 203776
rect 340196 203736 340202 203748
rect 354674 203736 354680 203748
rect 354732 203736 354738 203788
rect 340782 203668 340788 203720
rect 340840 203708 340846 203720
rect 342254 203708 342260 203720
rect 340840 203680 342260 203708
rect 340840 203668 340846 203680
rect 342254 203668 342260 203680
rect 342312 203668 342318 203720
rect 344922 203668 344928 203720
rect 344980 203708 344986 203720
rect 354306 203708 354312 203720
rect 344980 203680 354312 203708
rect 344980 203668 344986 203680
rect 354306 203668 354312 203680
rect 354364 203708 354370 203720
rect 354968 203708 354996 203816
rect 363506 203804 363512 203816
rect 363564 203844 363570 203856
rect 440234 203844 440240 203856
rect 363564 203816 440240 203844
rect 363564 203804 363570 203816
rect 440234 203804 440240 203816
rect 440292 203804 440298 203856
rect 451918 203804 451924 203856
rect 451976 203844 451982 203856
rect 461394 203844 461400 203856
rect 451976 203816 461400 203844
rect 451976 203804 451982 203816
rect 461394 203804 461400 203816
rect 461452 203804 461458 203856
rect 463510 203804 463516 203856
rect 463568 203844 463574 203856
rect 506474 203844 506480 203856
rect 463568 203816 506480 203844
rect 463568 203804 463574 203816
rect 506474 203804 506480 203816
rect 506532 203804 506538 203856
rect 355594 203736 355600 203788
rect 355652 203776 355658 203788
rect 364702 203776 364708 203788
rect 355652 203748 364708 203776
rect 355652 203736 355658 203748
rect 364702 203736 364708 203748
rect 364760 203776 364766 203788
rect 437474 203776 437480 203788
rect 364760 203748 437480 203776
rect 364760 203736 364766 203748
rect 437474 203736 437480 203748
rect 437532 203736 437538 203788
rect 447870 203736 447876 203788
rect 447928 203776 447934 203788
rect 448422 203776 448428 203788
rect 447928 203748 448428 203776
rect 447928 203736 447934 203748
rect 448422 203736 448428 203748
rect 448480 203776 448486 203788
rect 457990 203776 457996 203788
rect 448480 203748 457996 203776
rect 448480 203736 448486 203748
rect 457990 203736 457996 203748
rect 458048 203736 458054 203788
rect 464982 203736 464988 203788
rect 465040 203776 465046 203788
rect 502334 203776 502340 203788
rect 465040 203748 502340 203776
rect 465040 203736 465046 203748
rect 502334 203736 502340 203748
rect 502392 203736 502398 203788
rect 354364 203680 354996 203708
rect 354364 203668 354370 203680
rect 462222 203668 462228 203720
rect 462280 203708 462286 203720
rect 483014 203708 483020 203720
rect 462280 203680 483020 203708
rect 462280 203668 462286 203680
rect 483014 203668 483020 203680
rect 483072 203668 483078 203720
rect 318702 203600 318708 203652
rect 318760 203640 318766 203652
rect 340874 203640 340880 203652
rect 318760 203612 340880 203640
rect 318760 203600 318766 203612
rect 340874 203600 340880 203612
rect 340932 203600 340938 203652
rect 349246 203640 349252 203652
rect 346872 203612 349252 203640
rect 321462 203532 321468 203584
rect 321520 203572 321526 203584
rect 339402 203572 339408 203584
rect 321520 203544 339408 203572
rect 321520 203532 321526 203544
rect 339402 203532 339408 203544
rect 339460 203532 339466 203584
rect 346762 203572 346768 203584
rect 339512 203544 346768 203572
rect 322842 203464 322848 203516
rect 322900 203504 322906 203516
rect 338114 203504 338120 203516
rect 322900 203476 338120 203504
rect 322900 203464 322906 203476
rect 338114 203464 338120 203476
rect 338172 203464 338178 203516
rect 338206 203464 338212 203516
rect 338264 203504 338270 203516
rect 339218 203504 339224 203516
rect 338264 203476 339224 203504
rect 338264 203464 338270 203476
rect 339218 203464 339224 203476
rect 339276 203504 339282 203516
rect 339512 203504 339540 203544
rect 346762 203532 346768 203544
rect 346820 203532 346826 203584
rect 339276 203476 339540 203504
rect 339276 203464 339282 203476
rect 339586 203464 339592 203516
rect 339644 203504 339650 203516
rect 346872 203504 346900 203612
rect 349246 203600 349252 203612
rect 349304 203600 349310 203652
rect 349338 203600 349344 203652
rect 349396 203640 349402 203652
rect 350994 203640 351000 203652
rect 349396 203612 351000 203640
rect 349396 203600 349402 203612
rect 350994 203600 351000 203612
rect 351052 203600 351058 203652
rect 353202 203600 353208 203652
rect 353260 203640 353266 203652
rect 362494 203640 362500 203652
rect 353260 203612 362500 203640
rect 353260 203600 353266 203612
rect 362494 203600 362500 203612
rect 362552 203640 362558 203652
rect 442994 203640 443000 203652
rect 362552 203612 443000 203640
rect 362552 203600 362558 203612
rect 442994 203600 443000 203612
rect 443052 203600 443058 203652
rect 466454 203600 466460 203652
rect 466512 203640 466518 203652
rect 478322 203640 478328 203652
rect 466512 203612 478328 203640
rect 466512 203600 466518 203612
rect 478322 203600 478328 203612
rect 478380 203600 478386 203652
rect 479518 203600 479524 203652
rect 479576 203640 479582 203652
rect 484394 203640 484400 203652
rect 479576 203612 484400 203640
rect 479576 203600 479582 203612
rect 484394 203600 484400 203612
rect 484452 203600 484458 203652
rect 346946 203532 346952 203584
rect 347004 203572 347010 203584
rect 348326 203572 348332 203584
rect 347004 203544 348332 203572
rect 347004 203532 347010 203544
rect 348326 203532 348332 203544
rect 348384 203572 348390 203584
rect 357802 203572 357808 203584
rect 348384 203544 357808 203572
rect 348384 203532 348390 203544
rect 357802 203532 357808 203544
rect 357860 203572 357866 203584
rect 452654 203572 452660 203584
rect 357860 203544 452660 203572
rect 357860 203532 357866 203544
rect 452654 203532 452660 203544
rect 452712 203532 452718 203584
rect 461394 203532 461400 203584
rect 461452 203572 461458 203584
rect 470686 203572 470692 203584
rect 461452 203544 470692 203572
rect 461452 203532 461458 203544
rect 470686 203532 470692 203544
rect 470744 203532 470750 203584
rect 347130 203504 347136 203516
rect 339644 203476 346900 203504
rect 346964 203476 347136 203504
rect 339644 203464 339650 203476
rect 328362 203396 328368 203448
rect 328420 203436 328426 203448
rect 337930 203436 337936 203448
rect 328420 203408 337936 203436
rect 328420 203396 328426 203408
rect 337930 203396 337936 203408
rect 337988 203436 337994 203448
rect 346964 203436 346992 203476
rect 347130 203464 347136 203476
rect 347188 203504 347194 203516
rect 469398 203504 469404 203516
rect 347188 203476 349292 203504
rect 347188 203464 347194 203476
rect 337988 203408 346992 203436
rect 337988 203396 337994 203408
rect 347038 203396 347044 203448
rect 347096 203436 347102 203448
rect 349154 203436 349160 203448
rect 347096 203408 349160 203436
rect 347096 203396 347102 203408
rect 349154 203396 349160 203408
rect 349212 203396 349218 203448
rect 349264 203436 349292 203476
rect 465092 203476 469404 203504
rect 356422 203436 356428 203448
rect 349264 203408 356428 203436
rect 356422 203396 356428 203408
rect 356480 203436 356486 203448
rect 455414 203436 455420 203448
rect 356480 203408 455420 203436
rect 356480 203396 356486 203408
rect 455414 203396 455420 203408
rect 455472 203396 455478 203448
rect 456150 203396 456156 203448
rect 456208 203436 456214 203448
rect 456208 203408 457944 203436
rect 456208 203396 456214 203408
rect 328270 203328 328276 203380
rect 328328 203368 328334 203380
rect 335354 203368 335360 203380
rect 328328 203340 335360 203368
rect 328328 203328 328334 203340
rect 335354 203328 335360 203340
rect 335412 203328 335418 203380
rect 336642 203328 336648 203380
rect 336700 203368 336706 203380
rect 345934 203368 345940 203380
rect 336700 203340 345940 203368
rect 336700 203328 336706 203340
rect 345934 203328 345940 203340
rect 345992 203368 345998 203380
rect 355594 203368 355600 203380
rect 345992 203340 355600 203368
rect 345992 203328 345998 203340
rect 355594 203328 355600 203340
rect 355652 203328 355658 203380
rect 358722 203328 358728 203380
rect 358780 203368 358786 203380
rect 368474 203368 368480 203380
rect 358780 203340 368480 203368
rect 358780 203328 358786 203340
rect 368474 203328 368480 203340
rect 368532 203328 368538 203380
rect 331122 203260 331128 203312
rect 331180 203300 331186 203312
rect 331180 203272 333836 203300
rect 331180 203260 331186 203272
rect 329742 203192 329748 203244
rect 329800 203232 329806 203244
rect 333808 203232 333836 203272
rect 333882 203260 333888 203312
rect 333940 203300 333946 203312
rect 342438 203300 342444 203312
rect 333940 203272 342444 203300
rect 333940 203260 333946 203272
rect 342438 203260 342444 203272
rect 342496 203300 342502 203312
rect 351730 203300 351736 203312
rect 342496 203272 351736 203300
rect 342496 203260 342502 203272
rect 351730 203260 351736 203272
rect 351788 203260 351794 203312
rect 357526 203260 357532 203312
rect 357584 203300 357590 203312
rect 358630 203300 358636 203312
rect 357584 203272 358636 203300
rect 357584 203260 357590 203272
rect 358630 203260 358636 203272
rect 358688 203300 358694 203312
rect 449894 203300 449900 203312
rect 358688 203272 449900 203300
rect 358688 203260 358694 203272
rect 449894 203260 449900 203272
rect 449952 203260 449958 203312
rect 457916 203300 457944 203408
rect 460566 203396 460572 203448
rect 460624 203436 460630 203448
rect 465092 203436 465120 203476
rect 469398 203464 469404 203476
rect 469456 203504 469462 203516
rect 477586 203504 477592 203516
rect 469456 203476 477592 203504
rect 469456 203464 469462 203476
rect 477586 203464 477592 203476
rect 477644 203464 477650 203516
rect 460624 203408 465120 203436
rect 460624 203396 460630 203408
rect 465166 203396 465172 203448
rect 465224 203436 465230 203448
rect 468478 203436 468484 203448
rect 465224 203408 468484 203436
rect 465224 203396 465230 203408
rect 468478 203396 468484 203408
rect 468536 203436 468542 203448
rect 468536 203408 476252 203436
rect 468536 203396 468542 203408
rect 457990 203328 457996 203380
rect 458048 203368 458054 203380
rect 467282 203368 467288 203380
rect 458048 203340 467288 203368
rect 458048 203328 458054 203340
rect 467282 203328 467288 203340
rect 467340 203368 467346 203380
rect 476114 203368 476120 203380
rect 467340 203340 476120 203368
rect 467340 203328 467346 203340
rect 476114 203328 476120 203340
rect 476172 203328 476178 203380
rect 476224 203368 476252 203408
rect 477126 203396 477132 203448
rect 477184 203436 477190 203448
rect 485774 203436 485780 203448
rect 477184 203408 485780 203436
rect 477184 203396 477190 203408
rect 485774 203396 485780 203408
rect 485832 203396 485838 203448
rect 477494 203368 477500 203380
rect 476224 203340 477500 203368
rect 477494 203328 477500 203340
rect 477552 203328 477558 203380
rect 477678 203328 477684 203380
rect 477736 203368 477742 203380
rect 477736 203340 479288 203368
rect 477736 203328 477742 203340
rect 464614 203300 464620 203312
rect 457916 203272 464620 203300
rect 464614 203260 464620 203272
rect 464672 203300 464678 203312
rect 466454 203300 466460 203312
rect 464672 203272 466460 203300
rect 464672 203260 464678 203272
rect 466454 203260 466460 203272
rect 466512 203260 466518 203312
rect 466546 203260 466552 203312
rect 466604 203300 466610 203312
rect 475562 203300 475568 203312
rect 466604 203272 475568 203300
rect 466604 203260 466610 203272
rect 475562 203260 475568 203272
rect 475620 203300 475626 203312
rect 479260 203300 479288 203340
rect 483014 203300 483020 203312
rect 475620 203272 479196 203300
rect 479260 203272 483020 203300
rect 475620 203260 475626 203272
rect 335170 203232 335176 203244
rect 329800 203204 333744 203232
rect 333808 203204 335176 203232
rect 329800 203192 329806 203204
rect 333716 203164 333744 203204
rect 335170 203192 335176 203204
rect 335228 203192 335234 203244
rect 335262 203192 335268 203244
rect 335320 203232 335326 203244
rect 343634 203232 343640 203244
rect 335320 203204 343640 203232
rect 335320 203192 335326 203204
rect 343634 203192 343640 203204
rect 343692 203232 343698 203244
rect 353202 203232 353208 203244
rect 343692 203204 353208 203232
rect 343692 203192 343698 203204
rect 353202 203192 353208 203204
rect 353260 203192 353266 203244
rect 472894 203232 472900 203244
rect 471716 203204 472900 203232
rect 338206 203164 338212 203176
rect 333716 203136 338212 203164
rect 338206 203124 338212 203136
rect 338264 203124 338270 203176
rect 338758 203124 338764 203176
rect 338816 203164 338822 203176
rect 356054 203164 356060 203176
rect 338816 203136 356060 203164
rect 338816 203124 338822 203136
rect 356054 203124 356060 203136
rect 356112 203124 356118 203176
rect 455046 203124 455052 203176
rect 455104 203164 455110 203176
rect 463602 203164 463608 203176
rect 455104 203136 463608 203164
rect 455104 203124 455110 203136
rect 463602 203124 463608 203136
rect 463660 203164 463666 203176
rect 471716 203164 471744 203204
rect 472894 203192 472900 203204
rect 472952 203232 472958 203244
rect 479168 203232 479196 203272
rect 483014 203260 483020 203272
rect 483072 203260 483078 203312
rect 484394 203232 484400 203244
rect 472952 203204 479104 203232
rect 479168 203204 484400 203232
rect 472952 203192 472958 203204
rect 479076 203164 479104 203204
rect 484394 203192 484400 203204
rect 484452 203192 484458 203244
rect 481634 203164 481640 203176
rect 463660 203136 471744 203164
rect 471808 203136 479012 203164
rect 479076 203136 481640 203164
rect 463660 203124 463666 203136
rect 471808 203108 471836 203136
rect 332318 203056 332324 203108
rect 332376 203096 332382 203108
rect 336458 203096 336464 203108
rect 332376 203068 336464 203096
rect 332376 203056 332382 203068
rect 336458 203056 336464 203068
rect 336516 203056 336522 203108
rect 336642 203056 336648 203108
rect 336700 203096 336706 203108
rect 344922 203096 344928 203108
rect 336700 203068 344928 203096
rect 336700 203056 336706 203068
rect 344922 203056 344928 203068
rect 344980 203056 344986 203108
rect 350994 203056 351000 203108
rect 351052 203096 351058 203108
rect 360010 203096 360016 203108
rect 351052 203068 360016 203096
rect 351052 203056 351058 203068
rect 360010 203056 360016 203068
rect 360068 203056 360074 203108
rect 453298 203056 453304 203108
rect 453356 203096 453362 203108
rect 462406 203096 462412 203108
rect 453356 203068 462412 203096
rect 453356 203056 453362 203068
rect 462406 203056 462412 203068
rect 462464 203096 462470 203108
rect 471790 203096 471796 203108
rect 462464 203068 471796 203096
rect 462464 203056 462470 203068
rect 471790 203056 471796 203068
rect 471848 203056 471854 203108
rect 471882 203056 471888 203108
rect 471940 203096 471946 203108
rect 478874 203096 478880 203108
rect 471940 203068 478880 203096
rect 471940 203056 471946 203068
rect 478874 203056 478880 203068
rect 478932 203056 478938 203108
rect 478984 203096 479012 203136
rect 481634 203124 481640 203136
rect 481692 203124 481698 203176
rect 480622 203096 480628 203108
rect 478984 203068 480628 203096
rect 480622 203056 480628 203068
rect 480680 203056 480686 203108
rect 341518 202988 341524 203040
rect 341576 203028 341582 203040
rect 353294 203028 353300 203040
rect 341576 203000 353300 203028
rect 341576 202988 341582 203000
rect 353294 202988 353300 203000
rect 353352 202988 353358 203040
rect 455322 202988 455328 203040
rect 455380 203028 455386 203040
rect 524414 203028 524420 203040
rect 455380 203000 524420 203028
rect 455380 202988 455386 203000
rect 524414 202988 524420 203000
rect 524472 202988 524478 203040
rect 280062 202920 280068 202972
rect 280120 202960 280126 202972
rect 357434 202960 357440 202972
rect 280120 202932 357440 202960
rect 280120 202920 280126 202932
rect 357434 202920 357440 202932
rect 357492 202920 357498 202972
rect 452562 202920 452568 202972
rect 452620 202960 452626 202972
rect 529934 202960 529940 202972
rect 452620 202932 529940 202960
rect 452620 202920 452626 202932
rect 529934 202920 529940 202932
rect 529992 202920 529998 202972
rect 315942 202852 315948 202904
rect 316000 202892 316006 202904
rect 342254 202892 342260 202904
rect 316000 202864 342260 202892
rect 316000 202852 316006 202864
rect 342254 202852 342260 202864
rect 342312 202852 342318 202904
rect 349338 202892 349344 202904
rect 342364 202864 349344 202892
rect 297358 202784 297364 202836
rect 297416 202824 297422 202836
rect 297910 202824 297916 202836
rect 297416 202796 297916 202824
rect 297416 202784 297422 202796
rect 297910 202784 297916 202796
rect 297968 202784 297974 202836
rect 342162 202784 342168 202836
rect 342220 202824 342226 202836
rect 342364 202824 342392 202864
rect 349338 202852 349344 202864
rect 349396 202852 349402 202904
rect 456610 202852 456616 202904
rect 456668 202892 456674 202904
rect 520274 202892 520280 202904
rect 456668 202864 520280 202892
rect 456668 202852 456674 202864
rect 520274 202852 520280 202864
rect 520332 202852 520338 202904
rect 542722 202852 542728 202904
rect 542780 202892 542786 202904
rect 542906 202892 542912 202904
rect 542780 202864 542912 202892
rect 542780 202852 542786 202864
rect 542906 202852 542912 202864
rect 542964 202852 542970 202904
rect 342220 202796 342392 202824
rect 342220 202784 342226 202796
rect 409874 202784 409880 202836
rect 409932 202824 409938 202836
rect 410518 202824 410524 202836
rect 409932 202796 410524 202824
rect 409932 202784 409938 202796
rect 410518 202784 410524 202796
rect 410576 202784 410582 202836
rect 387702 202172 387708 202224
rect 387760 202212 387766 202224
rect 500218 202212 500224 202224
rect 387760 202184 500224 202212
rect 387760 202172 387766 202184
rect 500218 202172 500224 202184
rect 500276 202172 500282 202224
rect 382182 202104 382188 202156
rect 382240 202144 382246 202156
rect 499758 202144 499764 202156
rect 382240 202116 499764 202144
rect 382240 202104 382246 202116
rect 499758 202104 499764 202116
rect 499816 202104 499822 202156
rect 410518 201560 410524 201612
rect 410576 201600 410582 201612
rect 500310 201600 500316 201612
rect 410576 201572 500316 201600
rect 410576 201560 410582 201572
rect 500310 201560 500316 201572
rect 500368 201560 500374 201612
rect 297910 201492 297916 201544
rect 297968 201532 297974 201544
rect 417418 201532 417424 201544
rect 297968 201504 417424 201532
rect 297968 201492 297974 201504
rect 417418 201492 417424 201504
rect 417476 201492 417482 201544
rect 447778 201152 447784 201204
rect 447836 201192 447842 201204
rect 499666 201192 499672 201204
rect 447836 201164 499672 201192
rect 447836 201152 447842 201164
rect 499666 201152 499672 201164
rect 499724 201152 499730 201204
rect 379422 201084 379428 201136
rect 379480 201124 379486 201136
rect 499850 201124 499856 201136
rect 379480 201096 499856 201124
rect 379480 201084 379486 201096
rect 499850 201084 499856 201096
rect 499908 201084 499914 201136
rect 378042 201016 378048 201068
rect 378100 201056 378106 201068
rect 499942 201056 499948 201068
rect 378100 201028 499948 201056
rect 378100 201016 378106 201028
rect 499942 201016 499948 201028
rect 500000 201016 500006 201068
rect 375282 200948 375288 201000
rect 375340 200988 375346 201000
rect 500034 200988 500040 201000
rect 375340 200960 500040 200988
rect 375340 200948 375346 200960
rect 500034 200948 500040 200960
rect 500092 200948 500098 201000
rect 372522 200880 372528 200932
rect 372580 200920 372586 200932
rect 500126 200920 500132 200932
rect 372580 200892 500132 200920
rect 372580 200880 372586 200892
rect 500126 200880 500132 200892
rect 500184 200880 500190 200932
rect 4062 200812 4068 200864
rect 4120 200852 4126 200864
rect 543642 200852 543648 200864
rect 4120 200824 543648 200852
rect 4120 200812 4126 200824
rect 543642 200812 543648 200824
rect 543700 200812 543706 200864
rect 3510 200744 3516 200796
rect 3568 200784 3574 200796
rect 542538 200784 542544 200796
rect 3568 200756 542544 200784
rect 3568 200744 3574 200756
rect 542538 200744 542544 200756
rect 542596 200744 542602 200796
rect 542906 196092 542912 196104
rect 542832 196064 542912 196092
rect 542832 195968 542860 196064
rect 542906 196052 542912 196064
rect 542964 196052 542970 196104
rect 542814 195916 542820 195968
rect 542872 195916 542878 195968
rect 379790 183472 379796 183524
rect 379848 183512 379854 183524
rect 410518 183512 410524 183524
rect 379848 183484 410524 183512
rect 379848 183472 379854 183484
rect 410518 183472 410524 183484
rect 410576 183472 410582 183524
rect 543274 182112 543280 182164
rect 543332 182152 543338 182164
rect 580166 182152 580172 182164
rect 543332 182124 580172 182152
rect 543332 182112 543338 182124
rect 580166 182112 580172 182124
rect 580224 182112 580230 182164
rect 542814 173884 542820 173936
rect 542872 173924 542878 173936
rect 542998 173924 543004 173936
rect 542872 173896 543004 173924
rect 542872 173884 542878 173896
rect 542998 173884 543004 173896
rect 543056 173884 543062 173936
rect 544378 171028 544384 171080
rect 544436 171068 544442 171080
rect 580166 171068 580172 171080
rect 544436 171040 580172 171068
rect 544436 171028 544442 171040
rect 580166 171028 580172 171040
rect 580224 171028 580230 171080
rect 542814 162800 542820 162852
rect 542872 162840 542878 162852
rect 542998 162840 543004 162852
rect 542872 162812 543004 162840
rect 542872 162800 542878 162812
rect 542998 162800 543004 162812
rect 543056 162800 543062 162852
rect 543182 158652 543188 158704
rect 543240 158692 543246 158704
rect 579798 158692 579804 158704
rect 543240 158664 579804 158692
rect 543240 158652 543246 158664
rect 579798 158652 579804 158664
rect 579856 158652 579862 158704
rect 542814 153212 542820 153264
rect 542872 153252 542878 153264
rect 542998 153252 543004 153264
rect 542872 153224 543004 153252
rect 542872 153212 542878 153224
rect 542998 153212 543004 153224
rect 543056 153212 543062 153264
rect 542998 143488 543004 143540
rect 543056 143528 543062 143540
rect 543182 143528 543188 143540
rect 543056 143500 543188 143528
rect 543056 143488 543062 143500
rect 543182 143488 543188 143500
rect 543240 143488 543246 143540
rect 380066 137912 380072 137964
rect 380124 137952 380130 137964
rect 380158 137952 380164 137964
rect 380124 137924 380164 137952
rect 380124 137912 380130 137924
rect 380158 137912 380164 137924
rect 380216 137912 380222 137964
rect 379790 135192 379796 135244
rect 379848 135232 379854 135244
rect 380066 135232 380072 135244
rect 379848 135204 380072 135232
rect 379848 135192 379854 135204
rect 380066 135192 380072 135204
rect 380124 135192 380130 135244
rect 556798 135192 556804 135244
rect 556856 135232 556862 135244
rect 580166 135232 580172 135244
rect 556856 135204 580172 135232
rect 556856 135192 556862 135204
rect 580166 135192 580172 135204
rect 580224 135192 580230 135244
rect 542998 133900 543004 133952
rect 543056 133940 543062 133952
rect 543182 133940 543188 133952
rect 543056 133912 543188 133940
rect 543056 133900 543062 133912
rect 543182 133900 543188 133912
rect 543240 133900 543246 133952
rect 380802 124108 380808 124160
rect 380860 124148 380866 124160
rect 391934 124148 391940 124160
rect 380860 124120 391940 124148
rect 380860 124108 380866 124120
rect 391934 124108 391940 124120
rect 391992 124108 391998 124160
rect 542998 124108 543004 124160
rect 543056 124148 543062 124160
rect 543366 124148 543372 124160
rect 543056 124120 543372 124148
rect 543056 124108 543062 124120
rect 543366 124108 543372 124120
rect 543424 124108 543430 124160
rect 558178 124108 558184 124160
rect 558236 124148 558242 124160
rect 580166 124148 580172 124160
rect 558236 124120 580172 124148
rect 558236 124108 558242 124120
rect 580166 124108 580172 124120
rect 580224 124108 580230 124160
rect 380802 118396 380808 118448
rect 380860 118436 380866 118448
rect 388438 118436 388444 118448
rect 380860 118408 388444 118436
rect 380860 118396 380866 118408
rect 388438 118396 388444 118408
rect 388496 118396 388502 118448
rect 380710 115880 380716 115932
rect 380768 115920 380774 115932
rect 393958 115920 393964 115932
rect 380768 115892 393964 115920
rect 380768 115880 380774 115892
rect 393958 115880 393964 115892
rect 394016 115880 394022 115932
rect 380802 115812 380808 115864
rect 380860 115852 380866 115864
rect 391198 115852 391204 115864
rect 380860 115824 391204 115852
rect 380860 115812 380866 115824
rect 391198 115812 391204 115824
rect 391256 115812 391262 115864
rect 549898 111732 549904 111784
rect 549956 111772 549962 111784
rect 579798 111772 579804 111784
rect 549956 111744 579804 111772
rect 549956 111732 549962 111744
rect 579798 111732 579804 111744
rect 579856 111732 579862 111784
rect 300762 110916 300768 110968
rect 300820 110956 300826 110968
rect 416774 110956 416780 110968
rect 300820 110928 416780 110956
rect 300820 110916 300826 110928
rect 416774 110916 416780 110928
rect 416832 110916 416838 110968
rect 543090 109080 543096 109132
rect 543148 109080 543154 109132
rect 543108 108996 543136 109080
rect 3234 108944 3240 108996
rect 3292 108984 3298 108996
rect 542262 108984 542268 108996
rect 3292 108956 542268 108984
rect 3292 108944 3298 108956
rect 542262 108944 542268 108956
rect 542320 108944 542326 108996
rect 543090 108944 543096 108996
rect 543148 108944 543154 108996
rect 297910 108876 297916 108928
rect 297968 108916 297974 108928
rect 303614 108916 303620 108928
rect 297968 108888 303620 108916
rect 297968 108876 297974 108888
rect 303614 108876 303620 108888
rect 303672 108916 303678 108928
rect 305638 108916 305644 108928
rect 303672 108888 305644 108916
rect 303672 108876 303678 108888
rect 305638 108876 305644 108888
rect 305696 108916 305702 108928
rect 307754 108916 307760 108928
rect 305696 108888 307760 108916
rect 305696 108876 305702 108888
rect 307754 108876 307760 108888
rect 307812 108876 307818 108928
rect 418062 108876 418068 108928
rect 418120 108916 418126 108928
rect 424226 108916 424232 108928
rect 418120 108888 424232 108916
rect 418120 108876 418126 108888
rect 424226 108876 424232 108888
rect 424284 108916 424290 108928
rect 427814 108916 427820 108928
rect 424284 108888 427820 108916
rect 424284 108876 424290 108888
rect 427814 108876 427820 108888
rect 427872 108876 427878 108928
rect 542998 99356 543004 99408
rect 543056 99396 543062 99408
rect 543182 99396 543188 99408
rect 543056 99368 543188 99396
rect 543056 99356 543062 99368
rect 543182 99356 543188 99368
rect 543240 99356 543246 99408
rect 542814 96568 542820 96620
rect 542872 96608 542878 96620
rect 542906 96608 542912 96620
rect 542872 96580 542912 96608
rect 542872 96568 542878 96580
rect 542906 96568 542912 96580
rect 542964 96568 542970 96620
rect 48222 93712 48228 93764
rect 48280 93712 48286 93764
rect 48240 93560 48268 93712
rect 144914 93644 144920 93696
rect 144972 93684 144978 93696
rect 154482 93684 154488 93696
rect 144972 93656 154488 93684
rect 144972 93644 144978 93656
rect 154482 93644 154488 93656
rect 154540 93644 154546 93696
rect 38654 93508 38660 93560
rect 38712 93548 38718 93560
rect 48130 93548 48136 93560
rect 38712 93520 48136 93548
rect 38712 93508 38718 93520
rect 48130 93508 48136 93520
rect 48188 93508 48194 93560
rect 48222 93508 48228 93560
rect 48280 93508 48286 93560
rect 9582 93440 9588 93492
rect 9640 93440 9646 93492
rect 9600 93356 9628 93440
rect 9582 93304 9588 93356
rect 9640 93304 9646 93356
rect 542814 89700 542820 89752
rect 542872 89700 542878 89752
rect 542832 89672 542860 89700
rect 542906 89672 542912 89684
rect 542832 89644 542912 89672
rect 542906 89632 542912 89644
rect 542964 89632 542970 89684
rect 555418 88272 555424 88324
rect 555476 88312 555482 88324
rect 580166 88312 580172 88324
rect 555476 88284 580172 88312
rect 555476 88272 555482 88284
rect 580166 88272 580172 88284
rect 580224 88272 580230 88324
rect 542814 86912 542820 86964
rect 542872 86952 542878 86964
rect 543274 86952 543280 86964
rect 542872 86924 543280 86952
rect 542872 86912 542878 86924
rect 543274 86912 543280 86924
rect 543332 86912 543338 86964
rect 580166 77228 580172 77240
rect 543108 77200 580172 77228
rect 543108 77172 543136 77200
rect 580166 77188 580172 77200
rect 580224 77188 580230 77240
rect 543090 77120 543096 77172
rect 543148 77120 543154 77172
rect 542906 67600 542912 67652
rect 542964 67640 542970 67652
rect 543090 67640 543096 67652
rect 542964 67612 543096 67640
rect 542964 67600 542970 67612
rect 543090 67600 543096 67612
rect 543148 67600 543154 67652
rect 547138 64812 547144 64864
rect 547196 64852 547202 64864
rect 579798 64852 579804 64864
rect 547196 64824 579804 64852
rect 547196 64812 547202 64824
rect 579798 64812 579804 64824
rect 579856 64812 579862 64864
rect 543090 60772 543096 60784
rect 542832 60744 543096 60772
rect 542832 60716 542860 60744
rect 543090 60732 543096 60744
rect 543148 60732 543154 60784
rect 542814 60664 542820 60716
rect 542872 60664 542878 60716
rect 542814 51008 542820 51060
rect 542872 51048 542878 51060
rect 542998 51048 543004 51060
rect 542872 51020 543004 51048
rect 542872 51008 542878 51020
rect 542998 51008 543004 51020
rect 543056 51008 543062 51060
rect 542998 48220 543004 48272
rect 543056 48260 543062 48272
rect 543274 48260 543280 48272
rect 543056 48232 543280 48260
rect 543056 48220 543062 48232
rect 543274 48220 543280 48232
rect 543332 48220 543338 48272
rect 554038 41352 554044 41404
rect 554096 41392 554102 41404
rect 580166 41392 580172 41404
rect 554096 41364 580172 41392
rect 554096 41352 554102 41364
rect 580166 41352 580172 41364
rect 580224 41352 580230 41404
rect 543090 38632 543096 38684
rect 543148 38672 543154 38684
rect 543274 38672 543280 38684
rect 543148 38644 543280 38672
rect 543148 38632 543154 38644
rect 543274 38632 543280 38644
rect 543332 38632 543338 38684
rect 543090 30268 543096 30320
rect 543148 30308 543154 30320
rect 580166 30308 580172 30320
rect 543148 30280 580172 30308
rect 543148 30268 543154 30280
rect 580166 30268 580172 30280
rect 580224 30268 580230 30320
rect 545758 17892 545764 17944
rect 545816 17932 545822 17944
rect 579798 17932 579804 17944
rect 545816 17904 579804 17932
rect 545816 17892 545822 17904
rect 579798 17892 579804 17904
rect 579856 17892 579862 17944
rect 7650 3544 7656 3596
rect 7708 3584 7714 3596
rect 8202 3584 8208 3596
rect 7708 3556 8208 3584
rect 7708 3544 7714 3556
rect 8202 3544 8208 3556
rect 8260 3544 8266 3596
rect 8846 3544 8852 3596
rect 8904 3584 8910 3596
rect 9582 3584 9588 3596
rect 8904 3556 9588 3584
rect 8904 3544 8910 3556
rect 9582 3544 9588 3556
rect 9640 3544 9646 3596
rect 10042 3544 10048 3596
rect 10100 3584 10106 3596
rect 10962 3584 10968 3596
rect 10100 3556 10968 3584
rect 10100 3544 10106 3556
rect 10962 3544 10968 3556
rect 11020 3544 11026 3596
rect 11238 3544 11244 3596
rect 11296 3584 11302 3596
rect 12342 3584 12348 3596
rect 11296 3556 12348 3584
rect 11296 3544 11302 3556
rect 12342 3544 12348 3556
rect 12400 3544 12406 3596
rect 12434 3544 12440 3596
rect 12492 3584 12498 3596
rect 13630 3584 13636 3596
rect 12492 3556 13636 3584
rect 12492 3544 12498 3556
rect 13630 3544 13636 3556
rect 13688 3544 13694 3596
rect 16022 3544 16028 3596
rect 16080 3584 16086 3596
rect 16482 3584 16488 3596
rect 16080 3556 16488 3584
rect 16080 3544 16086 3556
rect 16482 3544 16488 3556
rect 16540 3544 16546 3596
rect 17218 3544 17224 3596
rect 17276 3584 17282 3596
rect 17862 3584 17868 3596
rect 17276 3556 17868 3584
rect 17276 3544 17282 3556
rect 17862 3544 17868 3556
rect 17920 3544 17926 3596
rect 18322 3544 18328 3596
rect 18380 3584 18386 3596
rect 19242 3584 19248 3596
rect 18380 3556 19248 3584
rect 18380 3544 18386 3556
rect 19242 3544 19248 3556
rect 19300 3544 19306 3596
rect 19518 3544 19524 3596
rect 19576 3584 19582 3596
rect 20622 3584 20628 3596
rect 19576 3556 20628 3584
rect 19576 3544 19582 3556
rect 20622 3544 20628 3556
rect 20680 3544 20686 3596
rect 20714 3544 20720 3596
rect 20772 3584 20778 3596
rect 21910 3584 21916 3596
rect 20772 3556 21916 3584
rect 20772 3544 20778 3556
rect 21910 3544 21916 3556
rect 21968 3544 21974 3596
rect 24302 3544 24308 3596
rect 24360 3584 24366 3596
rect 24762 3584 24768 3596
rect 24360 3556 24768 3584
rect 24360 3544 24366 3556
rect 24762 3544 24768 3556
rect 24820 3544 24826 3596
rect 25498 3544 25504 3596
rect 25556 3584 25562 3596
rect 26142 3584 26148 3596
rect 25556 3556 26148 3584
rect 25556 3544 25562 3556
rect 26142 3544 26148 3556
rect 26200 3544 26206 3596
rect 26694 3544 26700 3596
rect 26752 3584 26758 3596
rect 27522 3584 27528 3596
rect 26752 3556 27528 3584
rect 26752 3544 26758 3556
rect 27522 3544 27528 3556
rect 27580 3544 27586 3596
rect 27890 3544 27896 3596
rect 27948 3584 27954 3596
rect 28902 3584 28908 3596
rect 27948 3556 28908 3584
rect 27948 3544 27954 3556
rect 28902 3544 28908 3556
rect 28960 3544 28966 3596
rect 29086 3544 29092 3596
rect 29144 3584 29150 3596
rect 30190 3584 30196 3596
rect 29144 3556 30196 3584
rect 29144 3544 29150 3556
rect 30190 3544 30196 3556
rect 30248 3544 30254 3596
rect 33870 3544 33876 3596
rect 33928 3584 33934 3596
rect 34422 3584 34428 3596
rect 33928 3556 34428 3584
rect 33928 3544 33934 3556
rect 34422 3544 34428 3556
rect 34480 3544 34486 3596
rect 34974 3544 34980 3596
rect 35032 3584 35038 3596
rect 35802 3584 35808 3596
rect 35032 3556 35808 3584
rect 35032 3544 35038 3556
rect 35802 3544 35808 3556
rect 35860 3544 35866 3596
rect 36170 3544 36176 3596
rect 36228 3584 36234 3596
rect 37182 3584 37188 3596
rect 36228 3556 37188 3584
rect 36228 3544 36234 3556
rect 37182 3544 37188 3556
rect 37240 3544 37246 3596
rect 37366 3544 37372 3596
rect 37424 3584 37430 3596
rect 38470 3584 38476 3596
rect 37424 3556 38476 3584
rect 37424 3544 37430 3556
rect 38470 3544 38476 3556
rect 38528 3544 38534 3596
rect 42150 3544 42156 3596
rect 42208 3584 42214 3596
rect 42702 3584 42708 3596
rect 42208 3556 42708 3584
rect 42208 3544 42214 3556
rect 42702 3544 42708 3556
rect 42760 3544 42766 3596
rect 43346 3544 43352 3596
rect 43404 3584 43410 3596
rect 44082 3584 44088 3596
rect 43404 3556 44088 3584
rect 43404 3544 43410 3556
rect 44082 3544 44088 3556
rect 44140 3544 44146 3596
rect 44542 3544 44548 3596
rect 44600 3584 44606 3596
rect 45462 3584 45468 3596
rect 44600 3556 45468 3584
rect 44600 3544 44606 3556
rect 45462 3544 45468 3556
rect 45520 3544 45526 3596
rect 45738 3544 45744 3596
rect 45796 3584 45802 3596
rect 46842 3584 46848 3596
rect 45796 3556 46848 3584
rect 45796 3544 45802 3556
rect 46842 3544 46848 3556
rect 46900 3544 46906 3596
rect 46934 3544 46940 3596
rect 46992 3584 46998 3596
rect 48130 3584 48136 3596
rect 46992 3556 48136 3584
rect 46992 3544 46998 3556
rect 48130 3544 48136 3556
rect 48188 3544 48194 3596
rect 50522 3544 50528 3596
rect 50580 3584 50586 3596
rect 50982 3584 50988 3596
rect 50580 3556 50988 3584
rect 50580 3544 50586 3556
rect 50982 3544 50988 3556
rect 51040 3544 51046 3596
rect 51626 3544 51632 3596
rect 51684 3584 51690 3596
rect 52362 3584 52368 3596
rect 51684 3556 52368 3584
rect 51684 3544 51690 3556
rect 52362 3544 52368 3556
rect 52420 3544 52426 3596
rect 52822 3544 52828 3596
rect 52880 3584 52886 3596
rect 53742 3584 53748 3596
rect 52880 3556 53748 3584
rect 52880 3544 52886 3556
rect 53742 3544 53748 3556
rect 53800 3544 53806 3596
rect 54018 3544 54024 3596
rect 54076 3584 54082 3596
rect 55122 3584 55128 3596
rect 54076 3556 55128 3584
rect 54076 3544 54082 3556
rect 55122 3544 55128 3556
rect 55180 3544 55186 3596
rect 55214 3544 55220 3596
rect 55272 3584 55278 3596
rect 56410 3584 56416 3596
rect 55272 3556 56416 3584
rect 55272 3544 55278 3556
rect 56410 3544 56416 3556
rect 56468 3544 56474 3596
rect 58802 3544 58808 3596
rect 58860 3584 58866 3596
rect 59262 3584 59268 3596
rect 58860 3556 59268 3584
rect 58860 3544 58866 3556
rect 59262 3544 59268 3556
rect 59320 3544 59326 3596
rect 59998 3544 60004 3596
rect 60056 3584 60062 3596
rect 60642 3584 60648 3596
rect 60056 3556 60648 3584
rect 60056 3544 60062 3556
rect 60642 3544 60648 3556
rect 60700 3544 60706 3596
rect 61194 3544 61200 3596
rect 61252 3584 61258 3596
rect 62022 3584 62028 3596
rect 61252 3556 62028 3584
rect 61252 3544 61258 3556
rect 62022 3544 62028 3556
rect 62080 3544 62086 3596
rect 63586 3544 63592 3596
rect 63644 3584 63650 3596
rect 64690 3584 64696 3596
rect 63644 3556 64696 3584
rect 63644 3544 63650 3556
rect 64690 3544 64696 3556
rect 64748 3544 64754 3596
rect 68278 3544 68284 3596
rect 68336 3584 68342 3596
rect 68922 3584 68928 3596
rect 68336 3556 68928 3584
rect 68336 3544 68342 3556
rect 68922 3544 68928 3556
rect 68980 3544 68986 3596
rect 69474 3544 69480 3596
rect 69532 3584 69538 3596
rect 70302 3584 70308 3596
rect 69532 3556 70308 3584
rect 69532 3544 69538 3556
rect 70302 3544 70308 3556
rect 70360 3544 70366 3596
rect 70670 3544 70676 3596
rect 70728 3584 70734 3596
rect 71682 3584 71688 3596
rect 70728 3556 71688 3584
rect 70728 3544 70734 3556
rect 71682 3544 71688 3556
rect 71740 3544 71746 3596
rect 71866 3544 71872 3596
rect 71924 3584 71930 3596
rect 72970 3584 72976 3596
rect 71924 3556 72976 3584
rect 71924 3544 71930 3556
rect 72970 3544 72976 3556
rect 73028 3544 73034 3596
rect 76650 3544 76656 3596
rect 76708 3584 76714 3596
rect 77202 3584 77208 3596
rect 76708 3556 77208 3584
rect 76708 3544 76714 3556
rect 77202 3544 77208 3556
rect 77260 3544 77266 3596
rect 77846 3544 77852 3596
rect 77904 3584 77910 3596
rect 78582 3584 78588 3596
rect 77904 3556 78588 3584
rect 77904 3544 77910 3556
rect 78582 3544 78588 3556
rect 78640 3544 78646 3596
rect 79042 3544 79048 3596
rect 79100 3584 79106 3596
rect 79962 3584 79968 3596
rect 79100 3556 79968 3584
rect 79100 3544 79106 3556
rect 79962 3544 79968 3556
rect 80020 3544 80026 3596
rect 80238 3544 80244 3596
rect 80296 3584 80302 3596
rect 81342 3584 81348 3596
rect 80296 3556 81348 3584
rect 80296 3544 80302 3556
rect 81342 3544 81348 3556
rect 81400 3544 81406 3596
rect 81434 3544 81440 3596
rect 81492 3584 81498 3596
rect 82630 3584 82636 3596
rect 81492 3556 82636 3584
rect 81492 3544 81498 3556
rect 82630 3544 82636 3556
rect 82688 3544 82694 3596
rect 84930 3544 84936 3596
rect 84988 3584 84994 3596
rect 85482 3584 85488 3596
rect 84988 3556 85488 3584
rect 84988 3544 84994 3556
rect 85482 3544 85488 3556
rect 85540 3544 85546 3596
rect 86126 3544 86132 3596
rect 86184 3584 86190 3596
rect 86862 3584 86868 3596
rect 86184 3556 86868 3584
rect 86184 3544 86190 3556
rect 86862 3544 86868 3556
rect 86920 3544 86926 3596
rect 87322 3544 87328 3596
rect 87380 3584 87386 3596
rect 88242 3584 88248 3596
rect 87380 3556 88248 3584
rect 87380 3544 87386 3556
rect 88242 3544 88248 3556
rect 88300 3544 88306 3596
rect 88518 3544 88524 3596
rect 88576 3584 88582 3596
rect 89622 3584 89628 3596
rect 88576 3556 89628 3584
rect 88576 3544 88582 3556
rect 89622 3544 89628 3556
rect 89680 3544 89686 3596
rect 89714 3544 89720 3596
rect 89772 3584 89778 3596
rect 90910 3584 90916 3596
rect 89772 3556 90916 3584
rect 89772 3544 89778 3556
rect 90910 3544 90916 3556
rect 90968 3544 90974 3596
rect 93302 3544 93308 3596
rect 93360 3584 93366 3596
rect 93762 3584 93768 3596
rect 93360 3556 93768 3584
rect 93360 3544 93366 3556
rect 93762 3544 93768 3556
rect 93820 3544 93826 3596
rect 94498 3544 94504 3596
rect 94556 3584 94562 3596
rect 95142 3584 95148 3596
rect 94556 3556 95148 3584
rect 94556 3544 94562 3556
rect 95142 3544 95148 3556
rect 95200 3544 95206 3596
rect 95694 3544 95700 3596
rect 95752 3584 95758 3596
rect 96522 3584 96528 3596
rect 95752 3556 96528 3584
rect 95752 3544 95758 3556
rect 96522 3544 96528 3556
rect 96580 3544 96586 3596
rect 96890 3544 96896 3596
rect 96948 3584 96954 3596
rect 97902 3584 97908 3596
rect 96948 3556 97908 3584
rect 96948 3544 96954 3556
rect 97902 3544 97908 3556
rect 97960 3544 97966 3596
rect 98086 3544 98092 3596
rect 98144 3584 98150 3596
rect 99190 3584 99196 3596
rect 98144 3556 99196 3584
rect 98144 3544 98150 3556
rect 99190 3544 99196 3556
rect 99248 3544 99254 3596
rect 102778 3544 102784 3596
rect 102836 3584 102842 3596
rect 103422 3584 103428 3596
rect 102836 3556 103428 3584
rect 102836 3544 102842 3556
rect 103422 3544 103428 3556
rect 103480 3544 103486 3596
rect 103974 3544 103980 3596
rect 104032 3584 104038 3596
rect 104802 3584 104808 3596
rect 104032 3556 104808 3584
rect 104032 3544 104038 3556
rect 104802 3544 104808 3556
rect 104860 3544 104866 3596
rect 105170 3544 105176 3596
rect 105228 3584 105234 3596
rect 106182 3584 106188 3596
rect 105228 3556 106188 3584
rect 105228 3544 105234 3556
rect 106182 3544 106188 3556
rect 106240 3544 106246 3596
rect 106366 3544 106372 3596
rect 106424 3584 106430 3596
rect 107470 3584 107476 3596
rect 106424 3556 107476 3584
rect 106424 3544 106430 3556
rect 107470 3544 107476 3556
rect 107528 3544 107534 3596
rect 111150 3544 111156 3596
rect 111208 3584 111214 3596
rect 111702 3584 111708 3596
rect 111208 3556 111708 3584
rect 111208 3544 111214 3556
rect 111702 3544 111708 3556
rect 111760 3544 111766 3596
rect 112346 3544 112352 3596
rect 112404 3584 112410 3596
rect 113082 3584 113088 3596
rect 112404 3556 113088 3584
rect 112404 3544 112410 3556
rect 113082 3544 113088 3556
rect 113140 3544 113146 3596
rect 113542 3544 113548 3596
rect 113600 3584 113606 3596
rect 114462 3584 114468 3596
rect 113600 3556 114468 3584
rect 113600 3544 113606 3556
rect 114462 3544 114468 3556
rect 114520 3544 114526 3596
rect 114738 3544 114744 3596
rect 114796 3584 114802 3596
rect 115842 3584 115848 3596
rect 114796 3556 115848 3584
rect 114796 3544 114802 3556
rect 115842 3544 115848 3556
rect 115900 3544 115906 3596
rect 115934 3544 115940 3596
rect 115992 3584 115998 3596
rect 117130 3584 117136 3596
rect 115992 3556 117136 3584
rect 115992 3544 115998 3556
rect 117130 3544 117136 3556
rect 117188 3544 117194 3596
rect 119430 3544 119436 3596
rect 119488 3584 119494 3596
rect 119982 3584 119988 3596
rect 119488 3556 119988 3584
rect 119488 3544 119494 3556
rect 119982 3544 119988 3556
rect 120040 3544 120046 3596
rect 120626 3544 120632 3596
rect 120684 3584 120690 3596
rect 121362 3584 121368 3596
rect 120684 3556 121368 3584
rect 120684 3544 120690 3556
rect 121362 3544 121368 3556
rect 121420 3544 121426 3596
rect 121822 3544 121828 3596
rect 121880 3584 121886 3596
rect 122742 3584 122748 3596
rect 121880 3556 122748 3584
rect 121880 3544 121886 3556
rect 122742 3544 122748 3556
rect 122800 3544 122806 3596
rect 123018 3544 123024 3596
rect 123076 3584 123082 3596
rect 124122 3584 124128 3596
rect 123076 3556 124128 3584
rect 123076 3544 123082 3556
rect 124122 3544 124128 3556
rect 124180 3544 124186 3596
rect 124214 3544 124220 3596
rect 124272 3584 124278 3596
rect 125410 3584 125416 3596
rect 124272 3556 125416 3584
rect 124272 3544 124278 3556
rect 125410 3544 125416 3556
rect 125468 3544 125474 3596
rect 127802 3544 127808 3596
rect 127860 3584 127866 3596
rect 128262 3584 128268 3596
rect 127860 3556 128268 3584
rect 127860 3544 127866 3556
rect 128262 3544 128268 3556
rect 128320 3544 128326 3596
rect 128998 3544 129004 3596
rect 129056 3584 129062 3596
rect 129642 3584 129648 3596
rect 129056 3556 129648 3584
rect 129056 3544 129062 3556
rect 129642 3544 129648 3556
rect 129700 3544 129706 3596
rect 130194 3544 130200 3596
rect 130252 3584 130258 3596
rect 131022 3584 131028 3596
rect 130252 3556 131028 3584
rect 130252 3544 130258 3556
rect 131022 3544 131028 3556
rect 131080 3544 131086 3596
rect 131390 3544 131396 3596
rect 131448 3584 131454 3596
rect 132402 3584 132408 3596
rect 131448 3556 132408 3584
rect 131448 3544 131454 3556
rect 132402 3544 132408 3556
rect 132460 3544 132466 3596
rect 132586 3544 132592 3596
rect 132644 3584 132650 3596
rect 133782 3584 133788 3596
rect 132644 3556 133788 3584
rect 132644 3544 132650 3556
rect 133782 3544 133788 3556
rect 133840 3544 133846 3596
rect 566 3476 572 3528
rect 624 3516 630 3528
rect 1302 3516 1308 3528
rect 624 3488 1308 3516
rect 624 3476 630 3488
rect 1302 3476 1308 3488
rect 1360 3476 1366 3528
rect 1670 3476 1676 3528
rect 1728 3516 1734 3528
rect 2682 3516 2688 3528
rect 1728 3488 2688 3516
rect 1728 3476 1734 3488
rect 2682 3476 2688 3488
rect 2740 3476 2746 3528
rect 2866 3476 2872 3528
rect 2924 3516 2930 3528
rect 257430 3516 257436 3528
rect 2924 3488 257436 3516
rect 2924 3476 2930 3488
rect 257430 3476 257436 3488
rect 257488 3476 257494 3528
rect 4062 3408 4068 3460
rect 4120 3448 4126 3460
rect 257338 3448 257344 3460
rect 4120 3420 257344 3448
rect 4120 3408 4126 3420
rect 257338 3408 257344 3420
rect 257396 3408 257402 3460
rect 101582 3272 101588 3324
rect 101640 3312 101646 3324
rect 102042 3312 102048 3324
rect 101640 3284 102048 3312
rect 101640 3272 101646 3284
rect 102042 3272 102048 3284
rect 102100 3272 102106 3324
rect 62390 3136 62396 3188
rect 62448 3176 62454 3188
rect 63402 3176 63408 3188
rect 62448 3148 63408 3176
rect 62448 3136 62454 3148
rect 63402 3136 63408 3148
rect 63460 3136 63466 3188
rect 142062 2796 142068 2848
rect 142120 2836 142126 2848
rect 145650 2836 145656 2848
rect 142120 2808 145656 2836
rect 142120 2796 142126 2808
rect 145650 2796 145656 2808
rect 145708 2836 145714 2848
rect 149238 2836 149244 2848
rect 145708 2808 149244 2836
rect 145708 2796 145714 2808
rect 149238 2796 149244 2808
rect 149296 2836 149302 2848
rect 152734 2836 152740 2848
rect 149296 2808 152740 2836
rect 149296 2796 149302 2808
rect 152734 2796 152740 2808
rect 152792 2836 152798 2848
rect 156322 2836 156328 2848
rect 152792 2808 156328 2836
rect 152792 2796 152798 2808
rect 156322 2796 156328 2808
rect 156380 2836 156386 2848
rect 159910 2836 159916 2848
rect 156380 2808 159916 2836
rect 156380 2796 156386 2808
rect 159910 2796 159916 2808
rect 159968 2836 159974 2848
rect 163498 2836 163504 2848
rect 159968 2808 163504 2836
rect 159968 2796 159974 2808
rect 163498 2796 163504 2808
rect 163556 2836 163562 2848
rect 167086 2836 167092 2848
rect 163556 2808 167092 2836
rect 163556 2796 163562 2808
rect 167086 2796 167092 2808
rect 167144 2836 167150 2848
rect 170582 2836 170588 2848
rect 167144 2808 170588 2836
rect 167144 2796 167150 2808
rect 170582 2796 170588 2808
rect 170640 2836 170646 2848
rect 174170 2836 174176 2848
rect 170640 2808 174176 2836
rect 170640 2796 170646 2808
rect 174170 2796 174176 2808
rect 174228 2836 174234 2848
rect 177758 2836 177764 2848
rect 174228 2808 177764 2836
rect 174228 2796 174234 2808
rect 177758 2796 177764 2808
rect 177816 2836 177822 2848
rect 181346 2836 181352 2848
rect 177816 2808 181352 2836
rect 177816 2796 177822 2808
rect 181346 2796 181352 2808
rect 181404 2836 181410 2848
rect 184842 2836 184848 2848
rect 181404 2808 184848 2836
rect 181404 2796 181410 2808
rect 184842 2796 184848 2808
rect 184900 2836 184906 2848
rect 188430 2836 188436 2848
rect 184900 2808 188436 2836
rect 184900 2796 184906 2808
rect 188430 2796 188436 2808
rect 188488 2836 188494 2848
rect 192018 2836 192024 2848
rect 188488 2808 192024 2836
rect 188488 2796 188494 2808
rect 192018 2796 192024 2808
rect 192076 2836 192082 2848
rect 195606 2836 195612 2848
rect 192076 2808 195612 2836
rect 192076 2796 192082 2808
rect 195606 2796 195612 2808
rect 195664 2836 195670 2848
rect 199194 2836 199200 2848
rect 195664 2808 199200 2836
rect 195664 2796 195670 2808
rect 199194 2796 199200 2808
rect 199252 2836 199258 2848
rect 202690 2836 202696 2848
rect 199252 2808 202696 2836
rect 199252 2796 199258 2808
rect 202690 2796 202696 2808
rect 202748 2836 202754 2848
rect 206278 2836 206284 2848
rect 202748 2808 206284 2836
rect 202748 2796 202754 2808
rect 206278 2796 206284 2808
rect 206336 2836 206342 2848
rect 209866 2836 209872 2848
rect 206336 2808 209872 2836
rect 206336 2796 206342 2808
rect 209866 2796 209872 2808
rect 209924 2836 209930 2848
rect 213454 2836 213460 2848
rect 209924 2808 213460 2836
rect 209924 2796 209930 2808
rect 213454 2796 213460 2808
rect 213512 2836 213518 2848
rect 217042 2836 217048 2848
rect 213512 2808 217048 2836
rect 213512 2796 213518 2808
rect 217042 2796 217048 2808
rect 217100 2836 217106 2848
rect 220538 2836 220544 2848
rect 217100 2808 220544 2836
rect 217100 2796 217106 2808
rect 220538 2796 220544 2808
rect 220596 2836 220602 2848
rect 224126 2836 224132 2848
rect 220596 2808 224132 2836
rect 220596 2796 220602 2808
rect 224126 2796 224132 2808
rect 224184 2836 224190 2848
rect 227714 2836 227720 2848
rect 224184 2808 227720 2836
rect 224184 2796 224190 2808
rect 227714 2796 227720 2808
rect 227772 2836 227778 2848
rect 231302 2836 231308 2848
rect 227772 2808 231308 2836
rect 227772 2796 227778 2808
rect 231302 2796 231308 2808
rect 231360 2836 231366 2848
rect 234798 2836 234804 2848
rect 231360 2808 234804 2836
rect 231360 2796 231366 2808
rect 234798 2796 234804 2808
rect 234856 2836 234862 2848
rect 238386 2836 238392 2848
rect 234856 2808 238392 2836
rect 234856 2796 234862 2808
rect 238386 2796 238392 2808
rect 238444 2836 238450 2848
rect 241974 2836 241980 2848
rect 238444 2808 241980 2836
rect 238444 2796 238450 2808
rect 241974 2796 241980 2808
rect 242032 2836 242038 2848
rect 245562 2836 245568 2848
rect 242032 2808 245568 2836
rect 242032 2796 242038 2808
rect 245562 2796 245568 2808
rect 245620 2836 245626 2848
rect 249150 2836 249156 2848
rect 245620 2808 249156 2836
rect 245620 2796 245626 2808
rect 249150 2796 249156 2808
rect 249208 2836 249214 2848
rect 252646 2836 252652 2848
rect 249208 2808 252652 2836
rect 249208 2796 249214 2808
rect 252646 2796 252652 2808
rect 252704 2836 252710 2848
rect 256234 2836 256240 2848
rect 252704 2808 256240 2836
rect 252704 2796 252710 2808
rect 256234 2796 256240 2808
rect 256292 2836 256298 2848
rect 259822 2836 259828 2848
rect 256292 2808 259828 2836
rect 256292 2796 256298 2808
rect 259822 2796 259828 2808
rect 259880 2836 259886 2848
rect 263410 2836 263416 2848
rect 259880 2808 263416 2836
rect 259880 2796 259886 2808
rect 263410 2796 263416 2808
rect 263468 2836 263474 2848
rect 266998 2836 267004 2848
rect 263468 2808 267004 2836
rect 263468 2796 263474 2808
rect 266998 2796 267004 2808
rect 267056 2836 267062 2848
rect 270494 2836 270500 2848
rect 267056 2808 270500 2836
rect 267056 2796 267062 2808
rect 270494 2796 270500 2808
rect 270552 2836 270558 2848
rect 274082 2836 274088 2848
rect 270552 2808 274088 2836
rect 270552 2796 270558 2808
rect 274082 2796 274088 2808
rect 274140 2836 274146 2848
rect 277670 2836 277676 2848
rect 274140 2808 277676 2836
rect 274140 2796 274146 2808
rect 277670 2796 277676 2808
rect 277728 2836 277734 2848
rect 281258 2836 281264 2848
rect 277728 2808 281264 2836
rect 277728 2796 277734 2808
rect 281258 2796 281264 2808
rect 281316 2836 281322 2848
rect 284754 2836 284760 2848
rect 281316 2808 284760 2836
rect 281316 2796 281322 2808
rect 284754 2796 284760 2808
rect 284812 2836 284818 2848
rect 288342 2836 288348 2848
rect 284812 2808 288348 2836
rect 284812 2796 284818 2808
rect 288342 2796 288348 2808
rect 288400 2836 288406 2848
rect 291930 2836 291936 2848
rect 288400 2808 291936 2836
rect 288400 2796 288406 2808
rect 291930 2796 291936 2808
rect 291988 2836 291994 2848
rect 295518 2836 295524 2848
rect 291988 2808 295524 2836
rect 291988 2796 291994 2808
rect 295518 2796 295524 2808
rect 295576 2836 295582 2848
rect 299106 2836 299112 2848
rect 295576 2808 299112 2836
rect 295576 2796 295582 2808
rect 299106 2796 299112 2808
rect 299164 2836 299170 2848
rect 302602 2836 302608 2848
rect 299164 2808 302608 2836
rect 299164 2796 299170 2808
rect 302602 2796 302608 2808
rect 302660 2836 302666 2848
rect 305638 2836 305644 2848
rect 302660 2808 305644 2836
rect 302660 2796 302666 2808
rect 305638 2796 305644 2808
rect 305696 2836 305702 2848
rect 306190 2836 306196 2848
rect 305696 2808 306196 2836
rect 305696 2796 305702 2808
rect 306190 2796 306196 2808
rect 306248 2836 306254 2848
rect 309778 2836 309784 2848
rect 306248 2808 309784 2836
rect 306248 2796 306254 2808
rect 309778 2796 309784 2808
rect 309836 2836 309842 2848
rect 313366 2836 313372 2848
rect 309836 2808 313372 2836
rect 309836 2796 309842 2808
rect 313366 2796 313372 2808
rect 313424 2836 313430 2848
rect 316954 2836 316960 2848
rect 313424 2808 316960 2836
rect 313424 2796 313430 2808
rect 316954 2796 316960 2808
rect 317012 2836 317018 2848
rect 320450 2836 320456 2848
rect 317012 2808 320456 2836
rect 317012 2796 317018 2808
rect 320450 2796 320456 2808
rect 320508 2836 320514 2848
rect 324038 2836 324044 2848
rect 320508 2808 324044 2836
rect 320508 2796 320514 2808
rect 324038 2796 324044 2808
rect 324096 2836 324102 2848
rect 327626 2836 327632 2848
rect 324096 2808 327632 2836
rect 324096 2796 324102 2808
rect 327626 2796 327632 2808
rect 327684 2836 327690 2848
rect 331214 2836 331220 2848
rect 327684 2808 331220 2836
rect 327684 2796 327690 2808
rect 331214 2796 331220 2808
rect 331272 2836 331278 2848
rect 334710 2836 334716 2848
rect 331272 2808 334716 2836
rect 331272 2796 331278 2808
rect 334710 2796 334716 2808
rect 334768 2836 334774 2848
rect 338298 2836 338304 2848
rect 334768 2808 338304 2836
rect 334768 2796 334774 2808
rect 338298 2796 338304 2808
rect 338356 2836 338362 2848
rect 341886 2836 341892 2848
rect 338356 2808 341892 2836
rect 338356 2796 338362 2808
rect 341886 2796 341892 2808
rect 341944 2836 341950 2848
rect 345474 2836 345480 2848
rect 341944 2808 345480 2836
rect 341944 2796 341950 2808
rect 345474 2796 345480 2808
rect 345532 2836 345538 2848
rect 349062 2836 349068 2848
rect 345532 2808 349068 2836
rect 345532 2796 345538 2808
rect 349062 2796 349068 2808
rect 349120 2836 349126 2848
rect 352558 2836 352564 2848
rect 349120 2808 352564 2836
rect 349120 2796 349126 2808
rect 352558 2796 352564 2808
rect 352616 2836 352622 2848
rect 356146 2836 356152 2848
rect 352616 2808 356152 2836
rect 352616 2796 352622 2808
rect 356146 2796 356152 2808
rect 356204 2836 356210 2848
rect 359734 2836 359740 2848
rect 356204 2808 359740 2836
rect 356204 2796 356210 2808
rect 359734 2796 359740 2808
rect 359792 2836 359798 2848
rect 363322 2836 363328 2848
rect 359792 2808 363328 2836
rect 359792 2796 359798 2808
rect 363322 2796 363328 2808
rect 363380 2836 363386 2848
rect 366910 2836 366916 2848
rect 363380 2808 366916 2836
rect 363380 2796 363386 2808
rect 366910 2796 366916 2808
rect 366968 2836 366974 2848
rect 370406 2836 370412 2848
rect 366968 2808 370412 2836
rect 366968 2796 366974 2808
rect 370406 2796 370412 2808
rect 370464 2836 370470 2848
rect 373994 2836 374000 2848
rect 370464 2808 374000 2836
rect 370464 2796 370470 2808
rect 373994 2796 374000 2808
rect 374052 2836 374058 2848
rect 377582 2836 377588 2848
rect 374052 2808 377588 2836
rect 374052 2796 374058 2808
rect 377582 2796 377588 2808
rect 377640 2836 377646 2848
rect 381170 2836 381176 2848
rect 377640 2808 381176 2836
rect 377640 2796 377646 2808
rect 381170 2796 381176 2808
rect 381228 2836 381234 2848
rect 384666 2836 384672 2848
rect 381228 2808 384672 2836
rect 381228 2796 381234 2808
rect 384666 2796 384672 2808
rect 384724 2836 384730 2848
rect 388254 2836 388260 2848
rect 384724 2808 388260 2836
rect 384724 2796 384730 2808
rect 388254 2796 388260 2808
rect 388312 2836 388318 2848
rect 391842 2836 391848 2848
rect 388312 2808 391848 2836
rect 388312 2796 388318 2808
rect 391842 2796 391848 2808
rect 391900 2836 391906 2848
rect 395430 2836 395436 2848
rect 391900 2808 395436 2836
rect 391900 2796 391906 2808
rect 395430 2796 395436 2808
rect 395488 2836 395494 2848
rect 399018 2836 399024 2848
rect 395488 2808 399024 2836
rect 395488 2796 395494 2808
rect 399018 2796 399024 2808
rect 399076 2836 399082 2848
rect 402514 2836 402520 2848
rect 399076 2808 402520 2836
rect 399076 2796 399082 2808
rect 402514 2796 402520 2808
rect 402572 2836 402578 2848
rect 406102 2836 406108 2848
rect 402572 2808 406108 2836
rect 402572 2796 402578 2808
rect 406102 2796 406108 2808
rect 406160 2836 406166 2848
rect 409690 2836 409696 2848
rect 406160 2808 409696 2836
rect 406160 2796 406166 2808
rect 409690 2796 409696 2808
rect 409748 2836 409754 2848
rect 413278 2836 413284 2848
rect 409748 2808 413284 2836
rect 409748 2796 409754 2808
rect 413278 2796 413284 2808
rect 413336 2836 413342 2848
rect 416866 2836 416872 2848
rect 413336 2808 416872 2836
rect 413336 2796 413342 2808
rect 416866 2796 416872 2808
rect 416924 2836 416930 2848
rect 420362 2836 420368 2848
rect 416924 2808 420368 2836
rect 416924 2796 416930 2808
rect 420362 2796 420368 2808
rect 420420 2836 420426 2848
rect 423950 2836 423956 2848
rect 420420 2808 423956 2836
rect 420420 2796 420426 2808
rect 423950 2796 423956 2808
rect 424008 2836 424014 2848
rect 427538 2836 427544 2848
rect 424008 2808 427544 2836
rect 424008 2796 424014 2808
rect 427538 2796 427544 2808
rect 427596 2836 427602 2848
rect 431126 2836 431132 2848
rect 427596 2808 431132 2836
rect 427596 2796 427602 2808
rect 431126 2796 431132 2808
rect 431184 2836 431190 2848
rect 434622 2836 434628 2848
rect 431184 2808 434628 2836
rect 431184 2796 431190 2808
rect 434622 2796 434628 2808
rect 434680 2836 434686 2848
rect 438210 2836 438216 2848
rect 434680 2808 438216 2836
rect 434680 2796 434686 2808
rect 438210 2796 438216 2808
rect 438268 2836 438274 2848
rect 441798 2836 441804 2848
rect 438268 2808 441804 2836
rect 438268 2796 438274 2808
rect 441798 2796 441804 2808
rect 441856 2836 441862 2848
rect 445386 2836 445392 2848
rect 441856 2808 445392 2836
rect 441856 2796 441862 2808
rect 445386 2796 445392 2808
rect 445444 2836 445450 2848
rect 448974 2836 448980 2848
rect 445444 2808 448980 2836
rect 445444 2796 445450 2808
rect 448974 2796 448980 2808
rect 449032 2836 449038 2848
rect 452470 2836 452476 2848
rect 449032 2808 452476 2836
rect 449032 2796 449038 2808
rect 452470 2796 452476 2808
rect 452528 2836 452534 2848
rect 456058 2836 456064 2848
rect 452528 2808 456064 2836
rect 452528 2796 452534 2808
rect 456058 2796 456064 2808
rect 456116 2836 456122 2848
rect 459646 2836 459652 2848
rect 456116 2808 459652 2836
rect 456116 2796 456122 2808
rect 459646 2796 459652 2808
rect 459704 2836 459710 2848
rect 463234 2836 463240 2848
rect 459704 2808 463240 2836
rect 459704 2796 459710 2808
rect 463234 2796 463240 2808
rect 463292 2836 463298 2848
rect 466822 2836 466828 2848
rect 463292 2808 466828 2836
rect 463292 2796 463298 2808
rect 466822 2796 466828 2808
rect 466880 2836 466886 2848
rect 470318 2836 470324 2848
rect 466880 2808 470324 2836
rect 466880 2796 466886 2808
rect 470318 2796 470324 2808
rect 470376 2836 470382 2848
rect 473906 2836 473912 2848
rect 470376 2808 473912 2836
rect 470376 2796 470382 2808
rect 473906 2796 473912 2808
rect 473964 2836 473970 2848
rect 477494 2836 477500 2848
rect 473964 2808 477500 2836
rect 473964 2796 473970 2808
rect 477494 2796 477500 2808
rect 477552 2836 477558 2848
rect 481082 2836 481088 2848
rect 477552 2808 481088 2836
rect 477552 2796 477558 2808
rect 481082 2796 481088 2808
rect 481140 2836 481146 2848
rect 484578 2836 484584 2848
rect 481140 2808 484584 2836
rect 481140 2796 481146 2808
rect 484578 2796 484584 2808
rect 484636 2836 484642 2848
rect 488166 2836 488172 2848
rect 484636 2808 488172 2836
rect 484636 2796 484642 2808
rect 488166 2796 488172 2808
rect 488224 2836 488230 2848
rect 491754 2836 491760 2848
rect 488224 2808 491760 2836
rect 488224 2796 488230 2808
rect 491754 2796 491760 2808
rect 491812 2836 491818 2848
rect 495342 2836 495348 2848
rect 491812 2808 495348 2836
rect 491812 2796 491818 2808
rect 495342 2796 495348 2808
rect 495400 2836 495406 2848
rect 498930 2836 498936 2848
rect 495400 2808 498936 2836
rect 495400 2796 495406 2808
rect 498930 2796 498936 2808
rect 498988 2836 498994 2848
rect 502426 2836 502432 2848
rect 498988 2808 502432 2836
rect 498988 2796 498994 2808
rect 502426 2796 502432 2808
rect 502484 2836 502490 2848
rect 506014 2836 506020 2848
rect 502484 2808 506020 2836
rect 502484 2796 502490 2808
rect 506014 2796 506020 2808
rect 506072 2836 506078 2848
rect 509602 2836 509608 2848
rect 506072 2808 509608 2836
rect 506072 2796 506078 2808
rect 509602 2796 509608 2808
rect 509660 2836 509666 2848
rect 513190 2836 513196 2848
rect 509660 2808 513196 2836
rect 509660 2796 509666 2808
rect 513190 2796 513196 2808
rect 513248 2836 513254 2848
rect 516778 2836 516784 2848
rect 513248 2808 516784 2836
rect 513248 2796 513254 2808
rect 516778 2796 516784 2808
rect 516836 2836 516842 2848
rect 520274 2836 520280 2848
rect 516836 2808 520280 2836
rect 516836 2796 516842 2808
rect 520274 2796 520280 2808
rect 520332 2836 520338 2848
rect 523862 2836 523868 2848
rect 520332 2808 523868 2836
rect 520332 2796 520338 2808
rect 523862 2796 523868 2808
rect 523920 2836 523926 2848
rect 527450 2836 527456 2848
rect 523920 2808 527456 2836
rect 523920 2796 523926 2808
rect 527450 2796 527456 2808
rect 527508 2836 527514 2848
rect 531038 2836 531044 2848
rect 527508 2808 531044 2836
rect 527508 2796 527514 2808
rect 531038 2796 531044 2808
rect 531096 2836 531102 2848
rect 534534 2836 534540 2848
rect 531096 2808 534540 2836
rect 531096 2796 531102 2808
rect 534534 2796 534540 2808
rect 534592 2836 534598 2848
rect 538122 2836 538128 2848
rect 534592 2808 538128 2836
rect 534592 2796 534598 2808
rect 538122 2796 538128 2808
rect 538180 2836 538186 2848
rect 541710 2836 541716 2848
rect 538180 2808 541716 2836
rect 538180 2796 538186 2808
rect 541710 2796 541716 2808
rect 541768 2836 541774 2848
rect 545298 2836 545304 2848
rect 541768 2808 545304 2836
rect 541768 2796 541774 2808
rect 545298 2796 545304 2808
rect 545356 2836 545362 2848
rect 548886 2836 548892 2848
rect 545356 2808 548892 2836
rect 545356 2796 545362 2808
rect 548886 2796 548892 2808
rect 548944 2836 548950 2848
rect 552382 2836 552388 2848
rect 548944 2808 552388 2836
rect 548944 2796 548950 2808
rect 552382 2796 552388 2808
rect 552440 2836 552446 2848
rect 555970 2836 555976 2848
rect 552440 2808 555976 2836
rect 552440 2796 552446 2808
rect 555970 2796 555976 2808
rect 556028 2836 556034 2848
rect 559558 2836 559564 2848
rect 556028 2808 559564 2836
rect 556028 2796 556034 2808
rect 559558 2796 559564 2808
rect 559616 2836 559622 2848
rect 563146 2836 563152 2848
rect 559616 2808 563152 2836
rect 559616 2796 559622 2808
rect 563146 2796 563152 2808
rect 563204 2836 563210 2848
rect 566734 2836 566740 2848
rect 563204 2808 566740 2836
rect 563204 2796 563210 2808
rect 566734 2796 566740 2808
rect 566792 2836 566798 2848
rect 570230 2836 570236 2848
rect 566792 2808 570236 2836
rect 566792 2796 566798 2808
rect 570230 2796 570236 2808
rect 570288 2836 570294 2848
rect 573818 2836 573824 2848
rect 570288 2808 573824 2836
rect 570288 2796 570294 2808
rect 573818 2796 573824 2808
rect 573876 2836 573882 2848
rect 577406 2836 577412 2848
rect 573876 2808 577412 2836
rect 573876 2796 573882 2808
rect 577406 2796 577412 2808
rect 577464 2836 577470 2848
rect 580994 2836 581000 2848
rect 577464 2808 581000 2836
rect 577464 2796 577470 2808
rect 580994 2796 581000 2808
rect 581052 2796 581058 2848
rect 5258 552 5264 604
rect 5316 592 5322 604
rect 5442 592 5448 604
rect 5316 564 5448 592
rect 5316 552 5322 564
rect 5442 552 5448 564
rect 5500 552 5506 604
rect 138474 552 138480 604
rect 138532 592 138538 604
rect 142062 592 142068 604
rect 138532 564 142068 592
rect 138532 552 138538 564
rect 142062 552 142068 564
rect 142120 552 142126 604
<< via1 >>
rect 478512 700884 478564 700936
rect 539600 700884 539652 700936
rect 413652 700816 413704 700868
rect 539692 700816 539744 700868
rect 348792 700748 348844 700800
rect 539784 700748 539836 700800
rect 332508 700680 332560 700732
rect 539140 700680 539192 700732
rect 235172 700612 235224 700664
rect 235908 700612 235960 700664
rect 283840 700612 283892 700664
rect 539232 700612 539284 700664
rect 218980 700544 219032 700596
rect 539968 700544 540020 700596
rect 202788 700476 202840 700528
rect 539876 700476 539928 700528
rect 154120 700408 154172 700460
rect 540060 700408 540112 700460
rect 72976 700340 73028 700392
rect 540152 700340 540204 700392
rect 40500 700272 40552 700324
rect 541072 700272 541124 700324
rect 549904 700272 549956 700324
rect 559656 700272 559708 700324
rect 397460 699932 397512 699984
rect 398748 699932 398800 699984
rect 494796 699796 494848 699848
rect 495348 699796 495400 699848
rect 105452 699660 105504 699712
rect 106188 699660 106240 699712
rect 170312 699660 170364 699712
rect 171048 699660 171100 699712
rect 300124 699660 300176 699712
rect 300768 699660 300820 699712
rect 364984 699660 365036 699712
rect 365628 699660 365680 699712
rect 429844 699660 429896 699712
rect 430488 699660 430540 699712
rect 462320 699660 462372 699712
rect 463608 699660 463660 699712
rect 527180 699660 527232 699712
rect 528468 699660 528520 699712
rect 563704 696940 563756 696992
rect 580172 696940 580224 696992
rect 554044 685856 554096 685908
rect 580172 685856 580224 685908
rect 3516 681708 3568 681760
rect 541164 681708 541216 681760
rect 543280 676132 543332 676184
rect 543556 676132 543608 676184
rect 547144 673480 547196 673532
rect 580172 673480 580224 673532
rect 3424 667904 3476 667956
rect 541256 667904 541308 667956
rect 3056 652740 3108 652792
rect 540244 652740 540296 652792
rect 560944 650020 560996 650072
rect 580172 650020 580224 650072
rect 543464 647232 543516 647284
rect 543556 647232 543608 647284
rect 543464 640364 543516 640416
rect 543556 640364 543608 640416
rect 565084 638936 565136 638988
rect 580172 638936 580224 638988
rect 543372 630640 543424 630692
rect 543556 630640 543608 630692
rect 545764 626560 545816 626612
rect 580172 626560 580224 626612
rect 267648 620236 267700 620288
rect 540336 620236 540388 620288
rect 488540 613368 488592 613420
rect 493968 613368 494020 613420
rect 373632 612756 373684 612808
rect 379612 612756 379664 612808
rect 488540 612756 488592 612808
rect 493968 612756 494020 612808
rect 499580 612756 499632 612808
rect 543372 611328 543424 611380
rect 543556 611328 543608 611380
rect 495348 610784 495400 610836
rect 541348 610784 541400 610836
rect 463608 610716 463660 610768
rect 539324 610716 539376 610768
rect 430488 610648 430540 610700
rect 541440 610648 541492 610700
rect 365628 610580 365680 610632
rect 541532 610580 541584 610632
rect 379980 610376 380032 610428
rect 496452 610376 496504 610428
rect 3424 610308 3476 610360
rect 541716 610308 541768 610360
rect 387708 605820 387760 605872
rect 416780 605820 416832 605872
rect 384948 604460 385000 604512
rect 416780 604460 416832 604512
rect 382188 603100 382240 603152
rect 416780 603100 416832 603152
rect 558184 603100 558236 603152
rect 580172 603100 580224 603152
rect 379428 601672 379480 601724
rect 416780 601672 416832 601724
rect 378048 600312 378100 600364
rect 416780 600312 416832 600364
rect 543372 592016 543424 592068
rect 543556 592016 543608 592068
rect 574744 592016 574796 592068
rect 580172 592016 580224 592068
rect 544384 579640 544436 579692
rect 580172 579640 580224 579692
rect 543372 572704 543424 572756
rect 543556 572704 543608 572756
rect 556804 556180 556856 556232
rect 580172 556180 580224 556232
rect 543372 553392 543424 553444
rect 543556 553392 543608 553444
rect 573364 545096 573416 545148
rect 580172 545096 580224 545148
rect 413928 539588 413980 539640
rect 416964 539588 417016 539640
rect 379520 538228 379572 538280
rect 379796 538228 379848 538280
rect 410524 538228 410576 538280
rect 416780 538228 416832 538280
rect 379520 536052 379572 536104
rect 379796 536052 379848 536104
rect 543372 534080 543424 534132
rect 543556 534080 543608 534132
rect 544476 532720 544528 532772
rect 580172 532720 580224 532772
rect 409880 521568 409932 521620
rect 410524 521568 410576 521620
rect 297272 520888 297324 520940
rect 409880 520888 409932 520940
rect 379612 518916 379664 518968
rect 379796 518916 379848 518968
rect 320088 518848 320140 518900
rect 328920 518848 328972 518900
rect 329656 518848 329708 518900
rect 348976 518848 349028 518900
rect 455420 518848 455472 518900
rect 289728 518780 289780 518832
rect 322940 518780 322992 518832
rect 327356 518780 327408 518832
rect 336924 518780 336976 518832
rect 345296 518780 345348 518832
rect 448520 518780 448572 518832
rect 448704 518780 448756 518832
rect 458364 518780 458416 518832
rect 307668 518712 307720 518764
rect 331312 518712 331364 518764
rect 331404 518712 331456 518764
rect 340604 518712 340656 518764
rect 346584 518712 346636 518764
rect 449900 518712 449952 518764
rect 451280 518712 451332 518764
rect 459560 518712 459612 518764
rect 314568 518644 314620 518696
rect 323124 518644 323176 518696
rect 332416 518644 332468 518696
rect 341524 518644 341576 518696
rect 443184 518644 443236 518696
rect 452568 518644 452620 518696
rect 318708 518576 318760 518628
rect 327356 518576 327408 518628
rect 329656 518576 329708 518628
rect 338120 518576 338172 518628
rect 347688 518576 347740 518628
rect 452660 518576 452712 518628
rect 321100 518508 321152 518560
rect 330116 518508 330168 518560
rect 339500 518508 339552 518560
rect 348976 518508 349028 518560
rect 442540 518508 442592 518560
rect 451280 518508 451332 518560
rect 457076 518644 457128 518696
rect 466460 518644 466512 518696
rect 461032 518508 461084 518560
rect 274548 518440 274600 518492
rect 316040 518440 316092 518492
rect 317328 518440 317380 518492
rect 326436 518440 326488 518492
rect 335820 518440 335872 518492
rect 345296 518440 345348 518492
rect 447968 518440 448020 518492
rect 457076 518440 457128 518492
rect 458364 518440 458416 518492
rect 466460 518440 466512 518492
rect 313188 518372 313240 518424
rect 271788 518304 271840 518356
rect 314660 518304 314712 518356
rect 317236 518372 317288 518424
rect 325424 518372 325476 518424
rect 325516 518372 325568 518424
rect 331404 518372 331456 518424
rect 333796 518372 333848 518424
rect 342996 518372 343048 518424
rect 369768 518372 369820 518424
rect 426440 518372 426492 518424
rect 444288 518372 444340 518424
rect 453764 518372 453816 518424
rect 462320 518372 462372 518424
rect 318800 518304 318852 518356
rect 336924 518304 336976 518356
rect 346584 518304 346636 518356
rect 357348 518304 357400 518356
rect 430580 518304 430632 518356
rect 435916 518304 435968 518356
rect 445392 518304 445444 518356
rect 455328 518304 455380 518356
rect 463700 518304 463752 518356
rect 269028 518236 269080 518288
rect 313280 518236 313332 518288
rect 315856 518236 315908 518288
rect 320180 518236 320232 518288
rect 325424 518236 325476 518288
rect 334716 518236 334768 518288
rect 343732 518236 343784 518288
rect 344376 518236 344428 518288
rect 354588 518236 354640 518288
rect 429292 518236 429344 518288
rect 303620 518168 303672 518220
rect 423680 518168 423732 518220
rect 436928 518168 436980 518220
rect 446404 518236 446456 518288
rect 456064 518236 456116 518288
rect 465080 518236 465132 518288
rect 286968 518100 287020 518152
rect 321744 518100 321796 518152
rect 331128 518100 331180 518152
rect 340880 518100 340932 518152
rect 351828 518100 351880 518152
rect 429200 518100 429252 518152
rect 440884 518100 440936 518152
rect 450176 518168 450228 518220
rect 459560 518168 459612 518220
rect 467840 518168 467892 518220
rect 285588 518032 285640 518084
rect 315856 518032 315908 518084
rect 315948 518032 316000 518084
rect 324320 518032 324372 518084
rect 325516 518032 325568 518084
rect 325608 518032 325660 518084
rect 339500 518032 339552 518084
rect 349068 518032 349120 518084
rect 425336 518032 425388 518084
rect 432604 518032 432656 518084
rect 442540 518032 442592 518084
rect 282828 517964 282880 518016
rect 318800 517964 318852 518016
rect 328368 517964 328420 518016
rect 339592 517964 339644 518016
rect 340604 517964 340656 518016
rect 437480 517964 437532 518016
rect 439504 517964 439556 518016
rect 448704 517964 448756 518016
rect 280068 517896 280120 517948
rect 317512 517896 317564 517948
rect 322848 517896 322900 517948
rect 338120 517896 338172 517948
rect 341524 517896 341576 517948
rect 440240 517896 440292 517948
rect 444104 517896 444156 517948
rect 469864 517896 469916 517948
rect 277308 517828 277360 517880
rect 317420 517828 317472 517880
rect 321468 517828 321520 517880
rect 336740 517828 336792 517880
rect 342996 517828 343048 517880
rect 443000 517828 443052 517880
rect 445576 517828 445628 517880
rect 476764 517828 476816 517880
rect 315948 517760 316000 517812
rect 333980 517760 334032 517812
rect 344376 517760 344428 517812
rect 445760 517760 445812 517812
rect 313188 517692 313240 517744
rect 332692 517692 332744 517744
rect 333888 517692 333940 517744
rect 342260 517692 342312 517744
rect 344284 517692 344336 517744
rect 347872 517692 347924 517744
rect 447048 517692 447100 517744
rect 474004 517692 474056 517744
rect 261116 517624 261168 517676
rect 303620 517624 303672 517676
rect 304908 517624 304960 517676
rect 329840 517624 329892 517676
rect 337384 517624 337436 517676
rect 343640 517624 343692 517676
rect 438124 517624 438176 517676
rect 447140 517624 447192 517676
rect 448336 517624 448388 517676
rect 471244 517624 471296 517676
rect 310428 517556 310480 517608
rect 332600 517556 332652 517608
rect 340788 517556 340840 517608
rect 346400 517556 346452 517608
rect 436744 517556 436796 517608
rect 437296 517556 437348 517608
rect 446404 517556 446456 517608
rect 266268 517488 266320 517540
rect 312176 517488 312228 517540
rect 325516 517488 325568 517540
rect 333796 517488 333848 517540
rect 339408 517488 339460 517540
rect 345204 517488 345256 517540
rect 346308 517488 346360 517540
rect 347780 517488 347832 517540
rect 434168 517488 434220 517540
rect 443184 517488 443236 517540
rect 445484 517488 445536 517540
rect 479524 517488 479576 517540
rect 543372 514768 543424 514820
rect 543556 514768 543608 514820
rect 379612 514020 379664 514072
rect 379796 514020 379848 514072
rect 434076 511980 434128 512032
rect 434168 511980 434220 512032
rect 3240 509260 3292 509312
rect 539508 509260 539560 509312
rect 555424 509260 555476 509312
rect 580172 509260 580224 509312
rect 543280 502324 543332 502376
rect 543556 502324 543608 502376
rect 379612 499536 379664 499588
rect 379796 499536 379848 499588
rect 571984 498176 572036 498228
rect 580172 498176 580224 498228
rect 3332 495456 3384 495508
rect 540980 495456 541032 495508
rect 379612 494708 379664 494760
rect 379796 494708 379848 494760
rect 433616 492600 433668 492652
rect 433892 492600 433944 492652
rect 543280 492600 543332 492652
rect 543556 492600 543608 492652
rect 398748 487772 398800 487824
rect 539416 487772 539468 487824
rect 544568 485800 544620 485852
rect 580172 485800 580224 485852
rect 281724 482944 281776 482996
rect 282828 482944 282880 482996
rect 311808 482944 311860 482996
rect 366456 482944 366508 482996
rect 371608 482944 371660 482996
rect 417516 482944 417568 482996
rect 433156 482944 433208 482996
rect 439504 482944 439556 482996
rect 455328 482944 455380 482996
rect 507768 482944 507820 482996
rect 307576 482876 307628 482928
rect 297456 482808 297508 482860
rect 386512 482808 386564 482860
rect 386972 482876 387024 482928
rect 387708 482876 387760 482928
rect 453948 482876 454000 482928
rect 505192 482876 505244 482928
rect 389548 482808 389600 482860
rect 456708 482808 456760 482860
rect 510252 482808 510304 482860
rect 297548 482740 297600 482792
rect 394700 482740 394752 482792
rect 430672 482740 430724 482792
rect 438124 482740 438176 482792
rect 458088 482740 458140 482792
rect 512828 482740 512880 482792
rect 284300 482672 284352 482724
rect 285588 482672 285640 482724
rect 297640 482672 297692 482724
rect 397276 482672 397328 482724
rect 428096 482672 428148 482724
rect 436744 482672 436796 482724
rect 459468 482672 459520 482724
rect 515404 482672 515456 482724
rect 297732 482604 297784 482656
rect 399852 482604 399904 482656
rect 425520 482604 425572 482656
rect 436928 482604 436980 482656
rect 460848 482604 460900 482656
rect 517980 482604 518032 482656
rect 279148 482536 279200 482588
rect 280068 482536 280120 482588
rect 297824 482536 297876 482588
rect 402428 482536 402480 482588
rect 412732 482536 412784 482588
rect 413928 482536 413980 482588
rect 422944 482536 422996 482588
rect 435364 482536 435416 482588
rect 460756 482536 460808 482588
rect 520556 482536 520608 482588
rect 297916 482468 297968 482520
rect 405004 482468 405056 482520
rect 433248 482468 433300 482520
rect 458916 482468 458968 482520
rect 463608 482468 463660 482520
rect 525708 482468 525760 482520
rect 298008 482400 298060 482452
rect 407580 482400 407632 482452
rect 434628 482400 434680 482452
rect 461492 482400 461544 482452
rect 462228 482400 462280 482452
rect 523132 482400 523184 482452
rect 297364 482332 297416 482384
rect 415308 482332 415360 482384
rect 420368 482332 420420 482384
rect 433800 482332 433852 482384
rect 436008 482332 436060 482384
rect 464068 482332 464120 482384
rect 464988 482332 465040 482384
rect 528284 482332 528336 482384
rect 261208 482264 261260 482316
rect 310336 482196 310388 482248
rect 363880 482196 363932 482248
rect 310244 482128 310296 482180
rect 361304 482128 361356 482180
rect 309048 482060 309100 482112
rect 358728 482060 358780 482112
rect 376760 482264 376812 482316
rect 378048 482264 378100 482316
rect 386512 482264 386564 482316
rect 392124 482264 392176 482316
rect 417792 482264 417844 482316
rect 432604 482264 432656 482316
rect 437388 482264 437440 482316
rect 466644 482264 466696 482316
rect 467748 482264 467800 482316
rect 533436 482264 533488 482316
rect 374184 482196 374236 482248
rect 417424 482196 417476 482248
rect 453856 482196 453908 482248
rect 502616 482196 502668 482248
rect 435824 482128 435876 482180
rect 440884 482128 440936 482180
rect 452568 482128 452620 482180
rect 500040 482128 500092 482180
rect 379796 482060 379848 482112
rect 451188 482060 451240 482112
rect 497464 482060 497516 482112
rect 276572 481992 276624 482044
rect 277308 481992 277360 482044
rect 292028 481992 292080 482044
rect 320180 481992 320232 482044
rect 320272 481992 320324 482044
rect 321468 481992 321520 482044
rect 321560 481992 321612 482044
rect 324504 481992 324556 482044
rect 333060 481992 333112 482044
rect 333888 481992 333940 482044
rect 338212 481992 338264 482044
rect 339408 481992 339460 482044
rect 343364 481992 343416 482044
rect 344284 481992 344336 482044
rect 351092 481992 351144 482044
rect 351828 481992 351880 482044
rect 353668 481992 353720 482044
rect 354588 481992 354640 482044
rect 449808 481992 449860 482044
rect 494888 481992 494940 482044
rect 294512 481924 294564 481976
rect 324412 481924 324464 481976
rect 325792 481924 325844 481976
rect 297088 481856 297140 481908
rect 325700 481856 325752 481908
rect 299664 481788 299716 481840
rect 327172 481788 327224 481840
rect 302240 481720 302292 481772
rect 328460 481720 328512 481772
rect 442908 481924 442960 481976
rect 479432 481924 479484 481976
rect 479524 481924 479576 481976
rect 484584 481924 484636 481976
rect 356152 481856 356204 481908
rect 357348 481856 357400 481908
rect 441528 481856 441580 481908
rect 476948 481856 477000 481908
rect 440148 481788 440200 481840
rect 474372 481788 474424 481840
rect 476764 481788 476816 481840
rect 487160 481856 487212 481908
rect 335360 481720 335412 481772
rect 335636 481720 335688 481772
rect 337384 481720 337436 481772
rect 438768 481720 438820 481772
rect 471796 481720 471848 481772
rect 474004 481720 474056 481772
rect 489736 481788 489788 481840
rect 477224 481720 477276 481772
rect 492312 481720 492364 481772
rect 315120 481652 315172 481704
rect 315948 481652 316000 481704
rect 317696 481652 317748 481704
rect 325700 481652 325752 481704
rect 438676 481652 438728 481704
rect 469220 481652 469272 481704
rect 469864 481652 469916 481704
rect 477132 481652 477184 481704
rect 477316 481652 477368 481704
rect 482008 481652 482060 481704
rect 3148 480224 3200 480276
rect 540612 480224 540664 480276
rect 528468 479816 528520 479868
rect 541808 479816 541860 479868
rect 300768 479748 300820 479800
rect 541900 479748 541952 479800
rect 235908 479680 235960 479732
rect 541992 479680 542044 479732
rect 171048 479612 171100 479664
rect 542084 479612 542136 479664
rect 106188 479544 106240 479596
rect 542176 479544 542228 479596
rect 3516 479476 3568 479528
rect 540520 479476 540572 479528
rect 260656 479136 260708 479188
rect 540888 479136 540940 479188
rect 260564 479068 260616 479120
rect 540796 479068 540848 479120
rect 260380 479000 260432 479052
rect 543464 479000 543516 479052
rect 260104 478932 260156 478984
rect 542452 478932 542504 478984
rect 135168 478864 135220 478916
rect 256700 478864 256752 478916
rect 259920 478864 259972 478916
rect 543188 478864 543240 478916
rect 259828 478524 259880 478576
rect 540704 478524 540756 478576
rect 260748 478456 260800 478508
rect 542728 478456 542780 478508
rect 260472 478388 260524 478440
rect 542636 478388 542688 478440
rect 260288 478320 260340 478372
rect 543556 478320 543608 478372
rect 3700 478252 3752 478304
rect 542912 478252 542964 478304
rect 3424 478184 3476 478236
rect 542820 478184 542872 478236
rect 3608 478116 3660 478168
rect 543004 478116 543056 478168
rect 260012 478048 260064 478100
rect 543096 478048 543148 478100
rect 260196 477980 260248 478032
rect 543280 477980 543332 478032
rect 133788 476076 133840 476128
rect 256700 476076 256752 476128
rect 543372 476076 543424 476128
rect 543648 476076 543700 476128
rect 132408 473356 132460 473408
rect 256700 473356 256752 473408
rect 131028 471996 131080 472048
rect 256700 471996 256752 472048
rect 129648 469208 129700 469260
rect 256700 469208 256752 469260
rect 128268 467848 128320 467900
rect 256700 467848 256752 467900
rect 126888 465060 126940 465112
rect 256700 465060 256752 465112
rect 125508 463700 125560 463752
rect 256700 463700 256752 463752
rect 567844 462340 567896 462392
rect 580172 462340 580224 462392
rect 125416 460912 125468 460964
rect 256700 460912 256752 460964
rect 543372 460912 543424 460964
rect 543648 460912 543700 460964
rect 124128 459552 124180 459604
rect 256700 459552 256752 459604
rect 122748 456764 122800 456816
rect 256700 456764 256752 456816
rect 121368 455404 121420 455456
rect 256700 455404 256752 455456
rect 119988 452616 120040 452668
rect 256700 452616 256752 452668
rect 3424 452548 3476 452600
rect 259828 452548 259880 452600
rect 542360 451936 542412 451988
rect 543372 451936 543424 451988
rect 118608 451256 118660 451308
rect 256700 451256 256752 451308
rect 563796 451256 563848 451308
rect 580172 451256 580224 451308
rect 117228 448536 117280 448588
rect 256700 448536 256752 448588
rect 117136 445748 117188 445800
rect 256700 445748 256752 445800
rect 542360 445272 542412 445324
rect 543740 445272 543792 445324
rect 115848 444388 115900 444440
rect 256700 444388 256752 444440
rect 114468 441600 114520 441652
rect 256700 441600 256752 441652
rect 543372 441600 543424 441652
rect 543740 441600 543792 441652
rect 113088 440240 113140 440292
rect 256700 440240 256752 440292
rect 554136 438880 554188 438932
rect 580172 438880 580224 438932
rect 3148 438812 3200 438864
rect 259920 438812 259972 438864
rect 111708 437452 111760 437504
rect 256700 437452 256752 437504
rect 543372 437384 543424 437436
rect 543280 436636 543332 436688
rect 110328 436092 110380 436144
rect 256700 436092 256752 436144
rect 108948 433304 109000 433356
rect 256700 433304 256752 433356
rect 107568 431944 107620 431996
rect 256700 431944 256752 431996
rect 107476 429156 107528 429208
rect 256700 429156 256752 429208
rect 106188 427796 106240 427848
rect 256700 427796 256752 427848
rect 543280 427796 543332 427848
rect 543372 427728 543424 427780
rect 104808 425076 104860 425128
rect 256700 425076 256752 425128
rect 3240 425008 3292 425060
rect 260012 425008 260064 425060
rect 103428 423648 103480 423700
rect 256700 423648 256752 423700
rect 102048 420928 102100 420980
rect 256700 420928 256752 420980
rect 100668 418140 100720 418192
rect 256700 418140 256752 418192
rect 543372 418140 543424 418192
rect 543464 418004 543516 418056
rect 99288 416780 99340 416832
rect 256700 416780 256752 416832
rect 565176 415420 565228 415472
rect 580172 415420 580224 415472
rect 99196 413992 99248 414044
rect 256700 413992 256752 414044
rect 540612 413516 540664 413568
rect 540796 413516 540848 413568
rect 97908 412632 97960 412684
rect 256700 412632 256752 412684
rect 96528 409844 96580 409896
rect 256700 409844 256752 409896
rect 95148 408484 95200 408536
rect 256700 408484 256752 408536
rect 93768 405696 93820 405748
rect 256700 405696 256752 405748
rect 543464 404472 543516 404524
rect 92388 404336 92440 404388
rect 256700 404336 256752 404388
rect 543464 404336 543516 404388
rect 549996 404336 550048 404388
rect 580172 404336 580224 404388
rect 91008 401616 91060 401668
rect 256700 401616 256752 401668
rect 90916 400188 90968 400240
rect 256700 400188 256752 400240
rect 89628 397468 89680 397520
rect 256700 397468 256752 397520
rect 88248 396040 88300 396092
rect 256700 396040 256752 396092
rect 3148 395972 3200 396024
rect 260748 395972 260800 396024
rect 86868 393320 86920 393372
rect 256700 393320 256752 393372
rect 544660 391960 544712 392012
rect 580172 391960 580224 392012
rect 85488 390532 85540 390584
rect 256700 390532 256752 390584
rect 84108 389172 84160 389224
rect 256700 389172 256752 389224
rect 82728 386384 82780 386436
rect 256700 386384 256752 386436
rect 543188 386316 543240 386368
rect 543464 386316 543516 386368
rect 82636 385024 82688 385076
rect 256700 385024 256752 385076
rect 81348 382236 81400 382288
rect 256700 382236 256752 382288
rect 79968 380876 80020 380928
rect 256700 380876 256752 380928
rect 3240 380808 3292 380860
rect 260656 380808 260708 380860
rect 78588 378156 78640 378208
rect 256700 378156 256752 378208
rect 77208 376728 77260 376780
rect 256700 376728 256752 376780
rect 543188 376728 543240 376780
rect 543372 376728 543424 376780
rect 75828 374008 75880 374060
rect 256700 374008 256752 374060
rect 74448 372580 74500 372632
rect 256700 372580 256752 372632
rect 73068 369860 73120 369912
rect 256700 369860 256752 369912
rect 72976 368500 73028 368552
rect 256700 368500 256752 368552
rect 3148 367004 3200 367056
rect 260564 367004 260616 367056
rect 543188 367004 543240 367056
rect 543464 367004 543516 367056
rect 71688 365712 71740 365764
rect 256700 365712 256752 365764
rect 539232 365644 539284 365696
rect 539508 365644 539560 365696
rect 70308 362924 70360 362976
rect 256700 362924 256752 362976
rect 68928 361564 68980 361616
rect 256700 361564 256752 361616
rect 67548 358776 67600 358828
rect 256700 358776 256752 358828
rect 66168 357416 66220 357468
rect 256700 357416 256752 357468
rect 539324 357416 539376 357468
rect 543188 357416 543240 357468
rect 543372 357416 543424 357468
rect 539324 357212 539376 357264
rect 64788 354696 64840 354748
rect 256700 354696 256752 354748
rect 64696 353268 64748 353320
rect 256700 353268 256752 353320
rect 63408 350548 63460 350600
rect 256700 350548 256752 350600
rect 62028 349120 62080 349172
rect 256700 349120 256752 349172
rect 60648 346400 60700 346452
rect 256700 346400 256752 346452
rect 59268 345040 59320 345092
rect 256700 345040 256752 345092
rect 57888 342252 57940 342304
rect 256700 342252 256752 342304
rect 56508 340892 56560 340944
rect 256700 340892 256752 340944
rect 539784 339464 539836 339516
rect 539968 339464 540020 339516
rect 56416 338104 56468 338156
rect 256700 338104 256752 338156
rect 3424 338036 3476 338088
rect 260472 338036 260524 338088
rect 542636 336200 542688 336252
rect 549904 336200 549956 336252
rect 55128 335316 55180 335368
rect 256700 335316 256752 335368
rect 53748 333956 53800 334008
rect 256700 333956 256752 334008
rect 542636 333888 542688 333940
rect 554044 333888 554096 333940
rect 542636 332528 542688 332580
rect 563704 332528 563756 332580
rect 52368 331236 52420 331288
rect 256700 331236 256752 331288
rect 50988 329808 51040 329860
rect 256700 329808 256752 329860
rect 542636 328856 542688 328908
rect 547144 328856 547196 328908
rect 542636 328380 542688 328432
rect 565084 328380 565136 328432
rect 49608 327088 49660 327140
rect 256700 327088 256752 327140
rect 48228 325660 48280 325712
rect 256700 325660 256752 325712
rect 542636 325592 542688 325644
rect 560944 325592 560996 325644
rect 3240 324232 3292 324284
rect 260380 324232 260432 324284
rect 542636 324164 542688 324216
rect 545764 324164 545816 324216
rect 48136 322940 48188 322992
rect 256700 322940 256752 322992
rect 46848 321580 46900 321632
rect 256700 321580 256752 321632
rect 542636 321512 542688 321564
rect 574744 321512 574796 321564
rect 542636 320084 542688 320136
rect 558184 320084 558236 320136
rect 45468 318792 45520 318844
rect 256700 318792 256752 318844
rect 44088 317432 44140 317484
rect 256700 317432 256752 317484
rect 542636 316888 542688 316940
rect 544384 316888 544436 316940
rect 42708 314644 42760 314696
rect 256700 314644 256752 314696
rect 542636 314576 542688 314628
rect 573364 314576 573416 314628
rect 41328 313284 41380 313336
rect 256700 313284 256752 313336
rect 542636 313216 542688 313268
rect 556804 313216 556856 313268
rect 39948 310496 40000 310548
rect 256700 310496 256752 310548
rect 542636 309952 542688 310004
rect 544476 309952 544528 310004
rect 3332 309068 3384 309120
rect 260288 309068 260340 309120
rect 542636 309068 542688 309120
rect 571984 309068 572036 309120
rect 38568 307776 38620 307828
rect 256700 307776 256752 307828
rect 38476 306348 38528 306400
rect 256700 306348 256752 306400
rect 542636 306280 542688 306332
rect 555424 306280 555476 306332
rect 542636 304852 542688 304904
rect 544568 304852 544620 304904
rect 37188 303628 37240 303680
rect 256700 303628 256752 303680
rect 35808 302200 35860 302252
rect 256700 302200 256752 302252
rect 542636 302132 542688 302184
rect 563796 302132 563848 302184
rect 542636 300772 542688 300824
rect 567844 300772 567896 300824
rect 34428 299480 34480 299532
rect 256700 299480 256752 299532
rect 33048 298120 33100 298172
rect 256700 298120 256752 298172
rect 542636 298052 542688 298104
rect 554136 298052 554188 298104
rect 542636 296624 542688 296676
rect 549996 296624 550048 296676
rect 31668 295332 31720 295384
rect 256700 295332 256752 295384
rect 3424 295264 3476 295316
rect 260196 295264 260248 295316
rect 30288 293972 30340 294024
rect 256700 293972 256752 294024
rect 542636 293904 542688 293956
rect 565176 293904 565228 293956
rect 542636 291252 542688 291304
rect 544660 291252 544712 291304
rect 30196 291184 30248 291236
rect 256700 291184 256752 291236
rect 28908 289824 28960 289876
rect 256700 289824 256752 289876
rect 542636 289756 542688 289808
rect 580356 289756 580408 289808
rect 542636 288328 542688 288380
rect 580264 288328 580316 288380
rect 27528 287036 27580 287088
rect 256700 287036 256752 287088
rect 26148 285676 26200 285728
rect 256700 285676 256752 285728
rect 542636 285608 542688 285660
rect 580448 285608 580500 285660
rect 542636 284248 542688 284300
rect 580632 284248 580684 284300
rect 24768 282888 24820 282940
rect 256700 282888 256752 282940
rect 542636 281460 542688 281512
rect 580540 281460 580592 281512
rect 23388 280168 23440 280220
rect 256700 280168 256752 280220
rect 3424 280100 3476 280152
rect 260104 280100 260156 280152
rect 541164 280100 541216 280152
rect 580724 280100 580776 280152
rect 22008 278740 22060 278792
rect 256700 278740 256752 278792
rect 21916 276020 21968 276072
rect 256700 276020 256752 276072
rect 542636 275272 542688 275324
rect 580172 275272 580224 275324
rect 20628 274660 20680 274712
rect 256700 274660 256752 274712
rect 19248 271872 19300 271924
rect 256700 271872 256752 271924
rect 17868 270512 17920 270564
rect 256700 270512 256752 270564
rect 16488 267724 16540 267776
rect 256700 267724 256752 267776
rect 15108 266364 15160 266416
rect 256700 266364 256752 266416
rect 543096 264868 543148 264920
rect 580172 264868 580224 264920
rect 13728 263576 13780 263628
rect 256700 263576 256752 263628
rect 13636 262216 13688 262268
rect 256700 262216 256752 262268
rect 12348 259428 12400 259480
rect 256700 259428 256752 259480
rect 10968 256708 11020 256760
rect 256700 256708 256752 256760
rect 542636 256708 542688 256760
rect 558184 256708 558236 256760
rect 9588 255280 9640 255332
rect 256700 255280 256752 255332
rect 542636 255280 542688 255332
rect 556804 255280 556856 255332
rect 8208 252560 8260 252612
rect 256700 252560 256752 252612
rect 542636 252560 542688 252612
rect 549904 252560 549956 252612
rect 543004 252492 543056 252544
rect 579804 252492 579856 252544
rect 6828 251200 6880 251252
rect 256700 251200 256752 251252
rect 5448 248412 5500 248464
rect 256700 248412 256752 248464
rect 542636 248412 542688 248464
rect 555424 248412 555476 248464
rect 542636 247052 542688 247104
rect 547144 247052 547196 247104
rect 542452 243176 542504 243228
rect 542728 243176 542780 243228
rect 2688 242904 2740 242956
rect 256976 242904 257028 242956
rect 542452 242904 542504 242956
rect 554044 242904 554096 242956
rect 3424 241068 3476 241120
rect 542728 241068 542780 241120
rect 270408 240592 270460 240644
rect 273260 240592 273312 240644
rect 273352 240592 273404 240644
rect 289820 240660 289872 240712
rect 299388 240660 299440 240712
rect 318800 240660 318852 240712
rect 328368 240660 328420 240712
rect 357440 240660 357492 240712
rect 367008 240660 367060 240712
rect 368020 240660 368072 240712
rect 257988 240524 258040 240576
rect 260840 240524 260892 240576
rect 289820 240524 289872 240576
rect 299388 240524 299440 240576
rect 318800 240524 318852 240576
rect 328368 240524 328420 240576
rect 260840 240388 260892 240440
rect 261116 240388 261168 240440
rect 270408 240388 270460 240440
rect 1308 240116 1360 240168
rect 257988 240116 258040 240168
rect 542452 240116 542504 240168
rect 545764 240116 545816 240168
rect 368020 240048 368072 240100
rect 373264 240048 373316 240100
rect 331128 238688 331180 238740
rect 340788 238688 340840 238740
rect 433248 238688 433300 238740
rect 449164 238688 449216 238740
rect 464068 238688 464120 238740
rect 477040 238688 477092 238740
rect 477224 238688 477276 238740
rect 497464 238688 497516 238740
rect 325332 238620 325384 238672
rect 336740 238620 336792 238672
rect 391204 238620 391256 238672
rect 405004 238620 405056 238672
rect 430672 238620 430724 238672
rect 450544 238620 450596 238672
rect 458916 238620 458968 238672
rect 479524 238620 479576 238672
rect 263692 238552 263744 238604
rect 297824 238552 297876 238604
rect 329748 238552 329800 238604
rect 343364 238552 343416 238604
rect 388444 238552 388496 238604
rect 402428 238552 402480 238604
rect 428096 238552 428148 238604
rect 451924 238552 451976 238604
rect 463608 238552 463660 238604
rect 505192 238552 505244 238604
rect 261208 238484 261260 238536
rect 297364 238484 297416 238536
rect 328368 238484 328420 238536
rect 345940 238484 345992 238536
rect 380348 238484 380400 238536
rect 394700 238484 394752 238536
rect 420368 238484 420420 238536
rect 456248 238484 456300 238536
rect 460848 238484 460900 238536
rect 512828 238484 512880 238536
rect 297088 238416 297140 238468
rect 347044 238416 347096 238468
rect 380256 238416 380308 238468
rect 397276 238416 397328 238468
rect 417792 238416 417844 238468
rect 456064 238416 456116 238468
rect 458088 238416 458140 238468
rect 517980 238416 518032 238468
rect 294512 238348 294564 238400
rect 344284 238348 344336 238400
rect 371148 238348 371200 238400
rect 389548 238348 389600 238400
rect 393964 238348 394016 238400
rect 407580 238348 407632 238400
rect 422944 238348 422996 238400
rect 454684 238348 454736 238400
rect 455236 238348 455288 238400
rect 523132 238348 523184 238400
rect 289452 238280 289504 238332
rect 341524 238280 341576 238332
rect 380440 238280 380492 238332
rect 415308 238280 415360 238332
rect 425520 238280 425572 238332
rect 453304 238280 453356 238332
rect 453948 238280 454000 238332
rect 528284 238280 528336 238332
rect 284300 238212 284352 238264
rect 338764 238212 338816 238264
rect 384488 238212 384540 238264
rect 447784 238212 447836 238264
rect 451188 238212 451240 238264
rect 533436 238212 533488 238264
rect 286876 238144 286928 238196
rect 340144 238144 340196 238196
rect 380164 238144 380216 238196
rect 399852 238144 399904 238196
rect 412732 238144 412784 238196
rect 496360 238144 496412 238196
rect 292028 238076 292080 238128
rect 345756 238076 345808 238128
rect 356152 238076 356204 238128
rect 478236 238076 478288 238128
rect 266268 238008 266320 238060
rect 345664 238008 345716 238060
rect 353668 238008 353720 238060
rect 477132 238008 477184 238060
rect 478328 238008 478380 238060
rect 500040 238008 500092 238060
rect 435824 237940 435876 237992
rect 447876 237940 447928 237992
rect 471888 237940 471940 237992
rect 487160 237940 487212 237992
rect 473268 237872 473320 237924
rect 484584 237872 484636 237924
rect 466644 237804 466696 237856
rect 476764 237804 476816 237856
rect 469220 237736 469272 237788
rect 478144 237736 478196 237788
rect 471796 237600 471848 237652
rect 477592 237600 477644 237652
rect 332508 237532 332560 237584
rect 338212 237532 338264 237584
rect 476028 237532 476080 237584
rect 479432 237532 479484 237584
rect 333888 237464 333940 237516
rect 335636 237464 335688 237516
rect 476948 237464 477000 237516
rect 482008 237464 482060 237516
rect 276572 237396 276624 237448
rect 277308 237396 277360 237448
rect 279148 237396 279200 237448
rect 280068 237396 280120 237448
rect 281724 237396 281776 237448
rect 282828 237396 282880 237448
rect 299664 237396 299716 237448
rect 300768 237396 300820 237448
rect 302240 237396 302292 237448
rect 303528 237396 303580 237448
rect 315120 237396 315172 237448
rect 315948 237396 316000 237448
rect 317696 237396 317748 237448
rect 318708 237396 318760 237448
rect 320272 237396 320324 237448
rect 321468 237396 321520 237448
rect 333060 237396 333112 237448
rect 333980 237396 334032 237448
rect 351092 237396 351144 237448
rect 351828 237396 351880 237448
rect 361304 237396 361356 237448
rect 362224 237396 362276 237448
rect 371608 237396 371660 237448
rect 372528 237396 372580 237448
rect 374184 237396 374236 237448
rect 375288 237396 375340 237448
rect 376760 237396 376812 237448
rect 378048 237396 378100 237448
rect 386972 237396 387024 237448
rect 387708 237396 387760 237448
rect 461492 237396 461544 237448
rect 462228 237396 462280 237448
rect 474372 237396 474424 237448
rect 477500 237396 477552 237448
rect 3424 237328 3476 237380
rect 540428 237328 540480 237380
rect 542176 234608 542228 234660
rect 542820 234608 542872 234660
rect 542636 231752 542688 231804
rect 542820 231752 542872 231804
rect 543556 229032 543608 229084
rect 580172 229032 580224 229084
rect 3148 223524 3200 223576
rect 542360 223524 542412 223576
rect 542636 222164 542688 222216
rect 542912 222164 542964 222216
rect 543464 217948 543516 218000
rect 580172 217948 580224 218000
rect 542912 215364 542964 215416
rect 542820 215228 542872 215280
rect 542728 212440 542780 212492
rect 542820 212440 542872 212492
rect 3424 208292 3476 208344
rect 541624 208292 541676 208344
rect 543372 205572 543424 205624
rect 579804 205572 579856 205624
rect 470508 205164 470560 205216
rect 488540 205164 488592 205216
rect 470416 205028 470468 205080
rect 491300 205028 491352 205080
rect 469128 204960 469180 205012
rect 494060 204960 494112 205012
rect 369768 204892 369820 204944
rect 490196 204892 490248 204944
rect 473820 204416 473872 204468
rect 477224 204416 477276 204468
rect 331036 204212 331088 204264
rect 334072 204212 334124 204264
rect 336372 204212 336424 204264
rect 342168 204212 342220 204264
rect 282828 204144 282880 204196
rect 345388 204280 345440 204332
rect 345296 204212 345348 204264
rect 349160 204212 349212 204264
rect 364248 204212 364300 204264
rect 365720 204212 365772 204264
rect 456064 204212 456116 204264
rect 456616 204212 456668 204264
rect 465080 204212 465132 204264
rect 477040 204212 477092 204264
rect 481640 204212 481692 204264
rect 345388 204144 345440 204196
rect 357440 204144 357492 204196
rect 362224 204144 362276 204196
rect 367100 204144 367152 204196
rect 467748 204144 467800 204196
rect 473820 204144 473872 204196
rect 478236 204144 478288 204196
rect 485780 204144 485832 204196
rect 300768 204076 300820 204128
rect 345296 204076 345348 204128
rect 345756 204076 345808 204128
rect 351920 204076 351972 204128
rect 449808 204076 449860 204128
rect 535460 204076 535512 204128
rect 303528 204008 303580 204060
rect 343824 204008 343876 204060
rect 304908 203940 304960 203992
rect 346400 204008 346452 204060
rect 349252 204008 349304 204060
rect 357532 204008 357584 204060
rect 360016 204008 360068 204060
rect 448520 204008 448572 204060
rect 449164 204008 449216 204060
rect 459008 204008 459060 204060
rect 465172 204008 465224 204060
rect 466552 204008 466604 204060
rect 474188 204008 474240 204060
rect 476672 204008 476724 204060
rect 476764 204008 476816 204060
rect 480444 204008 480496 204060
rect 344284 203940 344336 203992
rect 351092 203940 351144 203992
rect 351736 203940 351788 203992
rect 361304 203940 361356 203992
rect 445760 203940 445812 203992
rect 459468 203940 459520 203992
rect 514760 203940 514812 203992
rect 307668 203872 307720 203924
rect 345020 203872 345072 203924
rect 345664 203872 345716 203924
rect 364340 203872 364392 203924
rect 450544 203872 450596 203924
rect 460572 203872 460624 203924
rect 462136 203872 462188 203924
rect 509240 203872 509292 203924
rect 310428 203804 310480 203856
rect 343640 203804 343692 203856
rect 343824 203804 343876 203856
rect 347780 203804 347832 203856
rect 313188 203736 313240 203788
rect 332324 203736 332376 203788
rect 332416 203736 332468 203788
rect 336372 203736 336424 203788
rect 336464 203736 336516 203788
rect 340052 203736 340104 203788
rect 340144 203736 340196 203788
rect 354680 203736 354732 203788
rect 340788 203668 340840 203720
rect 342260 203668 342312 203720
rect 344928 203668 344980 203720
rect 354312 203668 354364 203720
rect 363512 203804 363564 203856
rect 440240 203804 440292 203856
rect 451924 203804 451976 203856
rect 461400 203804 461452 203856
rect 463516 203804 463568 203856
rect 506480 203804 506532 203856
rect 355600 203736 355652 203788
rect 364708 203736 364760 203788
rect 437480 203736 437532 203788
rect 447876 203736 447928 203788
rect 448428 203736 448480 203788
rect 457996 203736 458048 203788
rect 464988 203736 465040 203788
rect 502340 203736 502392 203788
rect 462228 203668 462280 203720
rect 483020 203668 483072 203720
rect 318708 203600 318760 203652
rect 340880 203600 340932 203652
rect 321468 203532 321520 203584
rect 339408 203532 339460 203584
rect 322848 203464 322900 203516
rect 338120 203464 338172 203516
rect 338212 203464 338264 203516
rect 339224 203464 339276 203516
rect 346768 203532 346820 203584
rect 339592 203464 339644 203516
rect 349252 203600 349304 203652
rect 349344 203600 349396 203652
rect 351000 203600 351052 203652
rect 353208 203600 353260 203652
rect 362500 203600 362552 203652
rect 443000 203600 443052 203652
rect 466460 203600 466512 203652
rect 478328 203600 478380 203652
rect 479524 203600 479576 203652
rect 484400 203600 484452 203652
rect 346952 203532 347004 203584
rect 348332 203532 348384 203584
rect 357808 203532 357860 203584
rect 452660 203532 452712 203584
rect 461400 203532 461452 203584
rect 470692 203532 470744 203584
rect 328368 203396 328420 203448
rect 337936 203396 337988 203448
rect 347136 203464 347188 203516
rect 347044 203396 347096 203448
rect 349160 203396 349212 203448
rect 356428 203396 356480 203448
rect 455420 203396 455472 203448
rect 456156 203396 456208 203448
rect 328276 203328 328328 203380
rect 335360 203328 335412 203380
rect 336648 203328 336700 203380
rect 345940 203328 345992 203380
rect 355600 203328 355652 203380
rect 358728 203328 358780 203380
rect 368480 203328 368532 203380
rect 331128 203260 331180 203312
rect 329748 203192 329800 203244
rect 333888 203260 333940 203312
rect 342444 203260 342496 203312
rect 351736 203260 351788 203312
rect 357532 203260 357584 203312
rect 358636 203260 358688 203312
rect 449900 203260 449952 203312
rect 460572 203396 460624 203448
rect 469404 203464 469456 203516
rect 477592 203464 477644 203516
rect 465172 203396 465224 203448
rect 468484 203396 468536 203448
rect 457996 203328 458048 203380
rect 467288 203328 467340 203380
rect 476120 203328 476172 203380
rect 477132 203396 477184 203448
rect 485780 203396 485832 203448
rect 477500 203328 477552 203380
rect 477684 203328 477736 203380
rect 464620 203260 464672 203312
rect 466460 203260 466512 203312
rect 466552 203260 466604 203312
rect 475568 203260 475620 203312
rect 335176 203192 335228 203244
rect 335268 203192 335320 203244
rect 343640 203192 343692 203244
rect 353208 203192 353260 203244
rect 338212 203124 338264 203176
rect 338764 203124 338816 203176
rect 356060 203124 356112 203176
rect 455052 203124 455104 203176
rect 463608 203124 463660 203176
rect 472900 203192 472952 203244
rect 483020 203260 483072 203312
rect 484400 203192 484452 203244
rect 332324 203056 332376 203108
rect 336464 203056 336516 203108
rect 336648 203056 336700 203108
rect 344928 203056 344980 203108
rect 351000 203056 351052 203108
rect 360016 203056 360068 203108
rect 453304 203056 453356 203108
rect 462412 203056 462464 203108
rect 471796 203056 471848 203108
rect 471888 203056 471940 203108
rect 478880 203056 478932 203108
rect 481640 203124 481692 203176
rect 480628 203056 480680 203108
rect 341524 202988 341576 203040
rect 353300 202988 353352 203040
rect 455328 202988 455380 203040
rect 524420 202988 524472 203040
rect 280068 202920 280120 202972
rect 357440 202920 357492 202972
rect 452568 202920 452620 202972
rect 529940 202920 529992 202972
rect 315948 202852 316000 202904
rect 342260 202852 342312 202904
rect 297364 202784 297416 202836
rect 297916 202784 297968 202836
rect 342168 202784 342220 202836
rect 349344 202852 349396 202904
rect 456616 202852 456668 202904
rect 520280 202852 520332 202904
rect 542728 202852 542780 202904
rect 542912 202852 542964 202904
rect 409880 202784 409932 202836
rect 410524 202784 410576 202836
rect 387708 202172 387760 202224
rect 500224 202172 500276 202224
rect 382188 202104 382240 202156
rect 499764 202104 499816 202156
rect 410524 201560 410576 201612
rect 500316 201560 500368 201612
rect 297916 201492 297968 201544
rect 417424 201492 417476 201544
rect 447784 201152 447836 201204
rect 499672 201152 499724 201204
rect 379428 201084 379480 201136
rect 499856 201084 499908 201136
rect 378048 201016 378100 201068
rect 499948 201016 500000 201068
rect 375288 200948 375340 201000
rect 500040 200948 500092 201000
rect 372528 200880 372580 200932
rect 500132 200880 500184 200932
rect 4068 200812 4120 200864
rect 543648 200812 543700 200864
rect 3516 200744 3568 200796
rect 542544 200744 542596 200796
rect 542912 196052 542964 196104
rect 542820 195916 542872 195968
rect 379796 183472 379848 183524
rect 410524 183472 410576 183524
rect 543280 182112 543332 182164
rect 580172 182112 580224 182164
rect 542820 173884 542872 173936
rect 543004 173884 543056 173936
rect 544384 171028 544436 171080
rect 580172 171028 580224 171080
rect 542820 162800 542872 162852
rect 543004 162800 543056 162852
rect 543188 158652 543240 158704
rect 579804 158652 579856 158704
rect 542820 153212 542872 153264
rect 543004 153212 543056 153264
rect 543004 143488 543056 143540
rect 543188 143488 543240 143540
rect 380072 137912 380124 137964
rect 380164 137912 380216 137964
rect 379796 135192 379848 135244
rect 380072 135192 380124 135244
rect 556804 135192 556856 135244
rect 580172 135192 580224 135244
rect 543004 133900 543056 133952
rect 543188 133900 543240 133952
rect 380808 124108 380860 124160
rect 391940 124108 391992 124160
rect 543004 124108 543056 124160
rect 543372 124108 543424 124160
rect 558184 124108 558236 124160
rect 580172 124108 580224 124160
rect 380808 118396 380860 118448
rect 388444 118396 388496 118448
rect 380716 115880 380768 115932
rect 393964 115880 394016 115932
rect 380808 115812 380860 115864
rect 391204 115812 391256 115864
rect 549904 111732 549956 111784
rect 579804 111732 579856 111784
rect 300768 110916 300820 110968
rect 416780 110916 416832 110968
rect 543096 109080 543148 109132
rect 3240 108944 3292 108996
rect 542268 108944 542320 108996
rect 543096 108944 543148 108996
rect 297916 108876 297968 108928
rect 303620 108876 303672 108928
rect 305644 108876 305696 108928
rect 307760 108876 307812 108928
rect 418068 108876 418120 108928
rect 424232 108876 424284 108928
rect 427820 108876 427872 108928
rect 543004 99356 543056 99408
rect 543188 99356 543240 99408
rect 542820 96568 542872 96620
rect 542912 96568 542964 96620
rect 48228 93712 48280 93764
rect 144920 93644 144972 93696
rect 154488 93644 154540 93696
rect 38660 93508 38712 93560
rect 48136 93508 48188 93560
rect 48228 93508 48280 93560
rect 9588 93440 9640 93492
rect 9588 93304 9640 93356
rect 542820 89700 542872 89752
rect 542912 89632 542964 89684
rect 555424 88272 555476 88324
rect 580172 88272 580224 88324
rect 542820 86912 542872 86964
rect 543280 86912 543332 86964
rect 580172 77188 580224 77240
rect 543096 77120 543148 77172
rect 542912 67600 542964 67652
rect 543096 67600 543148 67652
rect 547144 64812 547196 64864
rect 579804 64812 579856 64864
rect 543096 60732 543148 60784
rect 542820 60664 542872 60716
rect 542820 51008 542872 51060
rect 543004 51008 543056 51060
rect 543004 48220 543056 48272
rect 543280 48220 543332 48272
rect 554044 41352 554096 41404
rect 580172 41352 580224 41404
rect 543096 38632 543148 38684
rect 543280 38632 543332 38684
rect 543096 30268 543148 30320
rect 580172 30268 580224 30320
rect 545764 17892 545816 17944
rect 579804 17892 579856 17944
rect 7656 3544 7708 3596
rect 8208 3544 8260 3596
rect 8852 3544 8904 3596
rect 9588 3544 9640 3596
rect 10048 3544 10100 3596
rect 10968 3544 11020 3596
rect 11244 3544 11296 3596
rect 12348 3544 12400 3596
rect 12440 3544 12492 3596
rect 13636 3544 13688 3596
rect 16028 3544 16080 3596
rect 16488 3544 16540 3596
rect 17224 3544 17276 3596
rect 17868 3544 17920 3596
rect 18328 3544 18380 3596
rect 19248 3544 19300 3596
rect 19524 3544 19576 3596
rect 20628 3544 20680 3596
rect 20720 3544 20772 3596
rect 21916 3544 21968 3596
rect 24308 3544 24360 3596
rect 24768 3544 24820 3596
rect 25504 3544 25556 3596
rect 26148 3544 26200 3596
rect 26700 3544 26752 3596
rect 27528 3544 27580 3596
rect 27896 3544 27948 3596
rect 28908 3544 28960 3596
rect 29092 3544 29144 3596
rect 30196 3544 30248 3596
rect 33876 3544 33928 3596
rect 34428 3544 34480 3596
rect 34980 3544 35032 3596
rect 35808 3544 35860 3596
rect 36176 3544 36228 3596
rect 37188 3544 37240 3596
rect 37372 3544 37424 3596
rect 38476 3544 38528 3596
rect 42156 3544 42208 3596
rect 42708 3544 42760 3596
rect 43352 3544 43404 3596
rect 44088 3544 44140 3596
rect 44548 3544 44600 3596
rect 45468 3544 45520 3596
rect 45744 3544 45796 3596
rect 46848 3544 46900 3596
rect 46940 3544 46992 3596
rect 48136 3544 48188 3596
rect 50528 3544 50580 3596
rect 50988 3544 51040 3596
rect 51632 3544 51684 3596
rect 52368 3544 52420 3596
rect 52828 3544 52880 3596
rect 53748 3544 53800 3596
rect 54024 3544 54076 3596
rect 55128 3544 55180 3596
rect 55220 3544 55272 3596
rect 56416 3544 56468 3596
rect 58808 3544 58860 3596
rect 59268 3544 59320 3596
rect 60004 3544 60056 3596
rect 60648 3544 60700 3596
rect 61200 3544 61252 3596
rect 62028 3544 62080 3596
rect 63592 3544 63644 3596
rect 64696 3544 64748 3596
rect 68284 3544 68336 3596
rect 68928 3544 68980 3596
rect 69480 3544 69532 3596
rect 70308 3544 70360 3596
rect 70676 3544 70728 3596
rect 71688 3544 71740 3596
rect 71872 3544 71924 3596
rect 72976 3544 73028 3596
rect 76656 3544 76708 3596
rect 77208 3544 77260 3596
rect 77852 3544 77904 3596
rect 78588 3544 78640 3596
rect 79048 3544 79100 3596
rect 79968 3544 80020 3596
rect 80244 3544 80296 3596
rect 81348 3544 81400 3596
rect 81440 3544 81492 3596
rect 82636 3544 82688 3596
rect 84936 3544 84988 3596
rect 85488 3544 85540 3596
rect 86132 3544 86184 3596
rect 86868 3544 86920 3596
rect 87328 3544 87380 3596
rect 88248 3544 88300 3596
rect 88524 3544 88576 3596
rect 89628 3544 89680 3596
rect 89720 3544 89772 3596
rect 90916 3544 90968 3596
rect 93308 3544 93360 3596
rect 93768 3544 93820 3596
rect 94504 3544 94556 3596
rect 95148 3544 95200 3596
rect 95700 3544 95752 3596
rect 96528 3544 96580 3596
rect 96896 3544 96948 3596
rect 97908 3544 97960 3596
rect 98092 3544 98144 3596
rect 99196 3544 99248 3596
rect 102784 3544 102836 3596
rect 103428 3544 103480 3596
rect 103980 3544 104032 3596
rect 104808 3544 104860 3596
rect 105176 3544 105228 3596
rect 106188 3544 106240 3596
rect 106372 3544 106424 3596
rect 107476 3544 107528 3596
rect 111156 3544 111208 3596
rect 111708 3544 111760 3596
rect 112352 3544 112404 3596
rect 113088 3544 113140 3596
rect 113548 3544 113600 3596
rect 114468 3544 114520 3596
rect 114744 3544 114796 3596
rect 115848 3544 115900 3596
rect 115940 3544 115992 3596
rect 117136 3544 117188 3596
rect 119436 3544 119488 3596
rect 119988 3544 120040 3596
rect 120632 3544 120684 3596
rect 121368 3544 121420 3596
rect 121828 3544 121880 3596
rect 122748 3544 122800 3596
rect 123024 3544 123076 3596
rect 124128 3544 124180 3596
rect 124220 3544 124272 3596
rect 125416 3544 125468 3596
rect 127808 3544 127860 3596
rect 128268 3544 128320 3596
rect 129004 3544 129056 3596
rect 129648 3544 129700 3596
rect 130200 3544 130252 3596
rect 131028 3544 131080 3596
rect 131396 3544 131448 3596
rect 132408 3544 132460 3596
rect 132592 3544 132644 3596
rect 133788 3544 133840 3596
rect 572 3476 624 3528
rect 1308 3476 1360 3528
rect 1676 3476 1728 3528
rect 2688 3476 2740 3528
rect 2872 3476 2924 3528
rect 257436 3476 257488 3528
rect 4068 3408 4120 3460
rect 257344 3408 257396 3460
rect 101588 3272 101640 3324
rect 102048 3272 102100 3324
rect 62396 3136 62448 3188
rect 63408 3136 63460 3188
rect 142068 2796 142120 2848
rect 145656 2796 145708 2848
rect 149244 2796 149296 2848
rect 152740 2796 152792 2848
rect 156328 2796 156380 2848
rect 159916 2796 159968 2848
rect 163504 2796 163556 2848
rect 167092 2796 167144 2848
rect 170588 2796 170640 2848
rect 174176 2796 174228 2848
rect 177764 2796 177816 2848
rect 181352 2796 181404 2848
rect 184848 2796 184900 2848
rect 188436 2796 188488 2848
rect 192024 2796 192076 2848
rect 195612 2796 195664 2848
rect 199200 2796 199252 2848
rect 202696 2796 202748 2848
rect 206284 2796 206336 2848
rect 209872 2796 209924 2848
rect 213460 2796 213512 2848
rect 217048 2796 217100 2848
rect 220544 2796 220596 2848
rect 224132 2796 224184 2848
rect 227720 2796 227772 2848
rect 231308 2796 231360 2848
rect 234804 2796 234856 2848
rect 238392 2796 238444 2848
rect 241980 2796 242032 2848
rect 245568 2796 245620 2848
rect 249156 2796 249208 2848
rect 252652 2796 252704 2848
rect 256240 2796 256292 2848
rect 259828 2796 259880 2848
rect 263416 2796 263468 2848
rect 267004 2796 267056 2848
rect 270500 2796 270552 2848
rect 274088 2796 274140 2848
rect 277676 2796 277728 2848
rect 281264 2796 281316 2848
rect 284760 2796 284812 2848
rect 288348 2796 288400 2848
rect 291936 2796 291988 2848
rect 295524 2796 295576 2848
rect 299112 2796 299164 2848
rect 302608 2796 302660 2848
rect 305644 2796 305696 2848
rect 306196 2796 306248 2848
rect 309784 2796 309836 2848
rect 313372 2796 313424 2848
rect 316960 2796 317012 2848
rect 320456 2796 320508 2848
rect 324044 2796 324096 2848
rect 327632 2796 327684 2848
rect 331220 2796 331272 2848
rect 334716 2796 334768 2848
rect 338304 2796 338356 2848
rect 341892 2796 341944 2848
rect 345480 2796 345532 2848
rect 349068 2796 349120 2848
rect 352564 2796 352616 2848
rect 356152 2796 356204 2848
rect 359740 2796 359792 2848
rect 363328 2796 363380 2848
rect 366916 2796 366968 2848
rect 370412 2796 370464 2848
rect 374000 2796 374052 2848
rect 377588 2796 377640 2848
rect 381176 2796 381228 2848
rect 384672 2796 384724 2848
rect 388260 2796 388312 2848
rect 391848 2796 391900 2848
rect 395436 2796 395488 2848
rect 399024 2796 399076 2848
rect 402520 2796 402572 2848
rect 406108 2796 406160 2848
rect 409696 2796 409748 2848
rect 413284 2796 413336 2848
rect 416872 2796 416924 2848
rect 420368 2796 420420 2848
rect 423956 2796 424008 2848
rect 427544 2796 427596 2848
rect 431132 2796 431184 2848
rect 434628 2796 434680 2848
rect 438216 2796 438268 2848
rect 441804 2796 441856 2848
rect 445392 2796 445444 2848
rect 448980 2796 449032 2848
rect 452476 2796 452528 2848
rect 456064 2796 456116 2848
rect 459652 2796 459704 2848
rect 463240 2796 463292 2848
rect 466828 2796 466880 2848
rect 470324 2796 470376 2848
rect 473912 2796 473964 2848
rect 477500 2796 477552 2848
rect 481088 2796 481140 2848
rect 484584 2796 484636 2848
rect 488172 2796 488224 2848
rect 491760 2796 491812 2848
rect 495348 2796 495400 2848
rect 498936 2796 498988 2848
rect 502432 2796 502484 2848
rect 506020 2796 506072 2848
rect 509608 2796 509660 2848
rect 513196 2796 513248 2848
rect 516784 2796 516836 2848
rect 520280 2796 520332 2848
rect 523868 2796 523920 2848
rect 527456 2796 527508 2848
rect 531044 2796 531096 2848
rect 534540 2796 534592 2848
rect 538128 2796 538180 2848
rect 541716 2796 541768 2848
rect 545304 2796 545356 2848
rect 548892 2796 548944 2848
rect 552388 2796 552440 2848
rect 555976 2796 556028 2848
rect 559564 2796 559616 2848
rect 563152 2796 563204 2848
rect 566740 2796 566792 2848
rect 570236 2796 570288 2848
rect 573824 2796 573876 2848
rect 577412 2796 577464 2848
rect 581000 2796 581052 2848
rect 5264 552 5316 604
rect 5448 552 5500 604
rect 138480 552 138532 604
rect 142068 552 142120 604
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 700369 8156 703520
rect 24320 700505 24348 703520
rect 24306 700496 24362 700505
rect 24306 700431 24362 700440
rect 8114 700360 8170 700369
rect 40512 700330 40540 703520
rect 72988 700398 73016 703520
rect 89180 700641 89208 703520
rect 89166 700632 89222 700641
rect 89166 700567 89222 700576
rect 72976 700392 73028 700398
rect 72976 700334 73028 700340
rect 8114 700295 8170 700304
rect 40500 700324 40552 700330
rect 40500 700266 40552 700272
rect 105464 699718 105492 703520
rect 137848 700777 137876 703520
rect 137834 700768 137890 700777
rect 137834 700703 137890 700712
rect 154132 700466 154160 703520
rect 154120 700460 154172 700466
rect 154120 700402 154172 700408
rect 170324 699718 170352 703520
rect 202800 700534 202828 703520
rect 218992 700602 219020 703520
rect 235184 700670 235212 703520
rect 235172 700664 235224 700670
rect 235172 700606 235224 700612
rect 235908 700664 235960 700670
rect 235908 700606 235960 700612
rect 218980 700596 219032 700602
rect 218980 700538 219032 700544
rect 202788 700528 202840 700534
rect 202788 700470 202840 700476
rect 105452 699712 105504 699718
rect 105452 699654 105504 699660
rect 106188 699712 106240 699718
rect 106188 699654 106240 699660
rect 170312 699712 170364 699718
rect 170312 699654 170364 699660
rect 171048 699712 171100 699718
rect 171048 699654 171100 699660
rect 3514 682272 3570 682281
rect 3514 682207 3570 682216
rect 3528 681766 3556 682207
rect 3516 681760 3568 681766
rect 3516 681702 3568 681708
rect 3422 667992 3478 668001
rect 3422 667927 3424 667936
rect 3476 667927 3478 667936
rect 3424 667898 3476 667904
rect 3054 653576 3110 653585
rect 3054 653511 3110 653520
rect 3068 652798 3096 653511
rect 3056 652792 3108 652798
rect 3056 652734 3108 652740
rect 3422 624880 3478 624889
rect 3422 624815 3478 624824
rect 3436 623801 3464 624815
rect 3422 623792 3478 623801
rect 3422 623727 3478 623736
rect 3422 610464 3478 610473
rect 3422 610399 3478 610408
rect 3436 610366 3464 610399
rect 3424 610360 3476 610366
rect 3424 610302 3476 610308
rect 3422 596048 3478 596057
rect 3422 595983 3478 595992
rect 3238 509960 3294 509969
rect 3238 509895 3294 509904
rect 3252 509318 3280 509895
rect 3240 509312 3292 509318
rect 3240 509254 3292 509260
rect 3330 495544 3386 495553
rect 3330 495479 3332 495488
rect 3384 495479 3386 495488
rect 3332 495450 3384 495456
rect 3146 481128 3202 481137
rect 3146 481063 3202 481072
rect 3160 480282 3188 481063
rect 3148 480276 3200 480282
rect 3148 480218 3200 480224
rect 3436 478242 3464 595983
rect 3514 567352 3570 567361
rect 3514 567287 3570 567296
rect 3528 479534 3556 567287
rect 3606 553072 3662 553081
rect 3606 553007 3662 553016
rect 3516 479528 3568 479534
rect 3516 479470 3568 479476
rect 3424 478236 3476 478242
rect 3424 478178 3476 478184
rect 3620 478174 3648 553007
rect 3698 538656 3754 538665
rect 3698 538591 3754 538600
rect 3712 478310 3740 538591
rect 106200 479602 106228 699654
rect 171060 479670 171088 699654
rect 235920 479738 235948 700606
rect 267660 620294 267688 703520
rect 283852 700670 283880 703520
rect 283840 700664 283892 700670
rect 283840 700606 283892 700612
rect 300136 699718 300164 703520
rect 332520 700738 332548 703520
rect 348804 700806 348832 703520
rect 348792 700800 348844 700806
rect 348792 700742 348844 700748
rect 332508 700732 332560 700738
rect 332508 700674 332560 700680
rect 364996 699718 365024 703520
rect 397472 699990 397500 703520
rect 413664 700874 413692 703520
rect 413652 700868 413704 700874
rect 413652 700810 413704 700816
rect 397460 699984 397512 699990
rect 397460 699926 397512 699932
rect 398748 699984 398800 699990
rect 398748 699926 398800 699932
rect 300124 699712 300176 699718
rect 300124 699654 300176 699660
rect 300768 699712 300820 699718
rect 300768 699654 300820 699660
rect 364984 699712 365036 699718
rect 364984 699654 365036 699660
rect 365628 699712 365680 699718
rect 365628 699654 365680 699660
rect 267648 620288 267700 620294
rect 267648 620230 267700 620236
rect 298006 606656 298062 606665
rect 298006 606591 298062 606600
rect 297914 605432 297970 605441
rect 297914 605367 297970 605376
rect 297822 603800 297878 603809
rect 297822 603735 297878 603744
rect 297730 602576 297786 602585
rect 297730 602511 297786 602520
rect 297638 600944 297694 600953
rect 297638 600879 297694 600888
rect 297546 599856 297602 599865
rect 297546 599791 297602 599800
rect 297454 598088 297510 598097
rect 297454 598023 297510 598032
rect 297362 540288 297418 540297
rect 297362 540223 297418 540232
rect 297270 538520 297326 538529
rect 297270 538455 297326 538464
rect 297284 520946 297312 538455
rect 297272 520940 297324 520946
rect 297272 520882 297324 520888
rect 289728 518832 289780 518838
rect 289728 518774 289780 518780
rect 274548 518492 274600 518498
rect 274548 518434 274600 518440
rect 271788 518356 271840 518362
rect 271788 518298 271840 518304
rect 269028 518288 269080 518294
rect 269028 518230 269080 518236
rect 261116 517676 261168 517682
rect 261116 517618 261168 517624
rect 235908 479732 235960 479738
rect 235908 479674 235960 479680
rect 171048 479664 171100 479670
rect 171048 479606 171100 479612
rect 106188 479596 106240 479602
rect 106188 479538 106240 479544
rect 260656 479188 260708 479194
rect 260656 479130 260708 479136
rect 260564 479120 260616 479126
rect 260564 479062 260616 479068
rect 260380 479052 260432 479058
rect 260380 478994 260432 479000
rect 260104 478984 260156 478990
rect 256698 478952 256754 478961
rect 135168 478916 135220 478922
rect 260104 478926 260156 478932
rect 256698 478887 256700 478896
rect 135168 478858 135220 478864
rect 256752 478887 256754 478896
rect 259920 478916 259972 478922
rect 256700 478858 256752 478864
rect 259920 478858 259972 478864
rect 3700 478304 3752 478310
rect 3700 478246 3752 478252
rect 3608 478168 3660 478174
rect 3608 478110 3660 478116
rect 133788 476128 133840 476134
rect 133788 476070 133840 476076
rect 132408 473408 132460 473414
rect 132408 473350 132460 473356
rect 131028 472048 131080 472054
rect 131028 471990 131080 471996
rect 129648 469260 129700 469266
rect 129648 469202 129700 469208
rect 128268 467900 128320 467906
rect 128268 467842 128320 467848
rect 126888 465112 126940 465118
rect 126888 465054 126940 465060
rect 125508 463752 125560 463758
rect 125508 463694 125560 463700
rect 125416 460964 125468 460970
rect 125416 460906 125468 460912
rect 124128 459604 124180 459610
rect 124128 459546 124180 459552
rect 122748 456816 122800 456822
rect 122748 456758 122800 456764
rect 121368 455456 121420 455462
rect 121368 455398 121420 455404
rect 119988 452668 120040 452674
rect 119988 452610 120040 452616
rect 3424 452600 3476 452606
rect 3424 452542 3476 452548
rect 3436 452441 3464 452542
rect 3422 452432 3478 452441
rect 3422 452367 3478 452376
rect 118608 451308 118660 451314
rect 118608 451250 118660 451256
rect 117228 448588 117280 448594
rect 117228 448530 117280 448536
rect 117136 445800 117188 445806
rect 117136 445742 117188 445748
rect 115848 444440 115900 444446
rect 115848 444382 115900 444388
rect 114468 441652 114520 441658
rect 114468 441594 114520 441600
rect 113088 440292 113140 440298
rect 113088 440234 113140 440240
rect 3148 438864 3200 438870
rect 3148 438806 3200 438812
rect 3160 438025 3188 438806
rect 3146 438016 3202 438025
rect 3146 437951 3202 437960
rect 111708 437504 111760 437510
rect 111708 437446 111760 437452
rect 110328 436144 110380 436150
rect 110328 436086 110380 436092
rect 108948 433356 109000 433362
rect 108948 433298 109000 433304
rect 107568 431996 107620 432002
rect 107568 431938 107620 431944
rect 107476 429208 107528 429214
rect 107476 429150 107528 429156
rect 106188 427848 106240 427854
rect 106188 427790 106240 427796
rect 104808 425128 104860 425134
rect 104808 425070 104860 425076
rect 3240 425060 3292 425066
rect 3240 425002 3292 425008
rect 3252 423745 3280 425002
rect 3238 423736 3294 423745
rect 3238 423671 3294 423680
rect 103428 423700 103480 423706
rect 103428 423642 103480 423648
rect 102048 420980 102100 420986
rect 102048 420922 102100 420928
rect 100668 418192 100720 418198
rect 100668 418134 100720 418140
rect 99288 416832 99340 416838
rect 99288 416774 99340 416780
rect 99196 414044 99248 414050
rect 99196 413986 99248 413992
rect 97908 412684 97960 412690
rect 97908 412626 97960 412632
rect 96528 409896 96580 409902
rect 96528 409838 96580 409844
rect 95148 408536 95200 408542
rect 95148 408478 95200 408484
rect 93768 405748 93820 405754
rect 93768 405690 93820 405696
rect 92388 404388 92440 404394
rect 92388 404330 92440 404336
rect 91008 401668 91060 401674
rect 91008 401610 91060 401616
rect 90916 400240 90968 400246
rect 90916 400182 90968 400188
rect 89628 397520 89680 397526
rect 89628 397462 89680 397468
rect 88248 396092 88300 396098
rect 88248 396034 88300 396040
rect 3148 396024 3200 396030
rect 3148 395966 3200 395972
rect 3160 395049 3188 395966
rect 3146 395040 3202 395049
rect 3146 394975 3202 394984
rect 86868 393372 86920 393378
rect 86868 393314 86920 393320
rect 85488 390584 85540 390590
rect 85488 390526 85540 390532
rect 84108 389224 84160 389230
rect 84108 389166 84160 389172
rect 82728 386436 82780 386442
rect 82728 386378 82780 386384
rect 82636 385076 82688 385082
rect 82636 385018 82688 385024
rect 81348 382288 81400 382294
rect 81348 382230 81400 382236
rect 79968 380928 80020 380934
rect 79968 380870 80020 380876
rect 3240 380860 3292 380866
rect 3240 380802 3292 380808
rect 3252 380633 3280 380802
rect 3238 380624 3294 380633
rect 3238 380559 3294 380568
rect 78588 378208 78640 378214
rect 78588 378150 78640 378156
rect 77208 376780 77260 376786
rect 77208 376722 77260 376728
rect 75828 374060 75880 374066
rect 75828 374002 75880 374008
rect 74448 372632 74500 372638
rect 74448 372574 74500 372580
rect 73068 369912 73120 369918
rect 73068 369854 73120 369860
rect 72976 368552 73028 368558
rect 72976 368494 73028 368500
rect 3148 367056 3200 367062
rect 3148 366998 3200 367004
rect 3160 366217 3188 366998
rect 3146 366208 3202 366217
rect 3146 366143 3202 366152
rect 71688 365764 71740 365770
rect 71688 365706 71740 365712
rect 70308 362976 70360 362982
rect 70308 362918 70360 362924
rect 68928 361616 68980 361622
rect 68928 361558 68980 361564
rect 67548 358828 67600 358834
rect 67548 358770 67600 358776
rect 66168 357468 66220 357474
rect 66168 357410 66220 357416
rect 64788 354748 64840 354754
rect 64788 354690 64840 354696
rect 64696 353320 64748 353326
rect 64696 353262 64748 353268
rect 63408 350600 63460 350606
rect 63408 350542 63460 350548
rect 62028 349172 62080 349178
rect 62028 349114 62080 349120
rect 60648 346452 60700 346458
rect 60648 346394 60700 346400
rect 59268 345092 59320 345098
rect 59268 345034 59320 345040
rect 57888 342304 57940 342310
rect 57888 342246 57940 342252
rect 56508 340944 56560 340950
rect 56508 340886 56560 340892
rect 56416 338156 56468 338162
rect 56416 338098 56468 338104
rect 3424 338088 3476 338094
rect 3424 338030 3476 338036
rect 3436 337521 3464 338030
rect 3422 337512 3478 337521
rect 3422 337447 3478 337456
rect 55128 335368 55180 335374
rect 55128 335310 55180 335316
rect 53748 334008 53800 334014
rect 53748 333950 53800 333956
rect 52368 331288 52420 331294
rect 52368 331230 52420 331236
rect 50988 329860 51040 329866
rect 50988 329802 51040 329808
rect 49608 327140 49660 327146
rect 49608 327082 49660 327088
rect 48228 325712 48280 325718
rect 48228 325654 48280 325660
rect 3240 324284 3292 324290
rect 3240 324226 3292 324232
rect 3252 323105 3280 324226
rect 3238 323096 3294 323105
rect 3238 323031 3294 323040
rect 48136 322992 48188 322998
rect 48136 322934 48188 322940
rect 46848 321632 46900 321638
rect 46848 321574 46900 321580
rect 45468 318844 45520 318850
rect 45468 318786 45520 318792
rect 44088 317484 44140 317490
rect 44088 317426 44140 317432
rect 42708 314696 42760 314702
rect 42708 314638 42760 314644
rect 41328 313336 41380 313342
rect 41328 313278 41380 313284
rect 39948 310548 40000 310554
rect 39948 310490 40000 310496
rect 3332 309120 3384 309126
rect 3332 309062 3384 309068
rect 3344 308825 3372 309062
rect 3330 308816 3386 308825
rect 3330 308751 3386 308760
rect 38568 307828 38620 307834
rect 38568 307770 38620 307776
rect 38476 306400 38528 306406
rect 38476 306342 38528 306348
rect 37188 303680 37240 303686
rect 37188 303622 37240 303628
rect 35808 302252 35860 302258
rect 35808 302194 35860 302200
rect 34428 299532 34480 299538
rect 34428 299474 34480 299480
rect 33048 298172 33100 298178
rect 33048 298114 33100 298120
rect 31668 295384 31720 295390
rect 31668 295326 31720 295332
rect 3424 295316 3476 295322
rect 3424 295258 3476 295264
rect 3436 294409 3464 295258
rect 3422 294400 3478 294409
rect 3422 294335 3478 294344
rect 30288 294024 30340 294030
rect 30288 293966 30340 293972
rect 30196 291236 30248 291242
rect 30196 291178 30248 291184
rect 28908 289876 28960 289882
rect 28908 289818 28960 289824
rect 27528 287088 27580 287094
rect 27528 287030 27580 287036
rect 26148 285728 26200 285734
rect 26148 285670 26200 285676
rect 24768 282940 24820 282946
rect 24768 282882 24820 282888
rect 23388 280220 23440 280226
rect 23388 280162 23440 280168
rect 3424 280152 3476 280158
rect 3422 280120 3424 280129
rect 3476 280120 3478 280129
rect 3422 280055 3478 280064
rect 22008 278792 22060 278798
rect 22008 278734 22060 278740
rect 21916 276072 21968 276078
rect 21916 276014 21968 276020
rect 20628 274712 20680 274718
rect 20628 274654 20680 274660
rect 19248 271924 19300 271930
rect 19248 271866 19300 271872
rect 17868 270564 17920 270570
rect 17868 270506 17920 270512
rect 16488 267776 16540 267782
rect 16488 267718 16540 267724
rect 15108 266416 15160 266422
rect 15108 266358 15160 266364
rect 3422 265704 3478 265713
rect 3422 265639 3478 265648
rect 2688 242956 2740 242962
rect 2688 242898 2740 242904
rect 1308 240168 1360 240174
rect 1308 240110 1360 240116
rect 1320 3534 1348 240110
rect 2700 3534 2728 242898
rect 3436 241126 3464 265639
rect 13728 263628 13780 263634
rect 13728 263570 13780 263576
rect 13636 262268 13688 262274
rect 13636 262210 13688 262216
rect 12348 259480 12400 259486
rect 12348 259422 12400 259428
rect 10968 256760 11020 256766
rect 10968 256702 11020 256708
rect 9588 255332 9640 255338
rect 9588 255274 9640 255280
rect 8208 252612 8260 252618
rect 8208 252554 8260 252560
rect 3514 251288 3570 251297
rect 3514 251223 3570 251232
rect 6828 251252 6880 251258
rect 3424 241120 3476 241126
rect 3424 241062 3476 241068
rect 3528 240825 3556 251223
rect 6828 251194 6880 251200
rect 5448 248464 5500 248470
rect 5448 248406 5500 248412
rect 3514 240816 3570 240825
rect 3514 240751 3570 240760
rect 3424 237380 3476 237386
rect 3424 237322 3476 237328
rect 3436 237017 3464 237322
rect 3422 237008 3478 237017
rect 3422 236943 3478 236952
rect 3148 223576 3200 223582
rect 3148 223518 3200 223524
rect 3160 222601 3188 223518
rect 3146 222592 3202 222601
rect 3146 222527 3202 222536
rect 3424 208344 3476 208350
rect 3424 208286 3476 208292
rect 3436 208185 3464 208286
rect 3422 208176 3478 208185
rect 3422 208111 3478 208120
rect 3974 201104 4030 201113
rect 3974 201039 4030 201048
rect 3422 200968 3478 200977
rect 3422 200903 3478 200912
rect 3436 122097 3464 200903
rect 3790 200832 3846 200841
rect 3516 200796 3568 200802
rect 3790 200767 3846 200776
rect 3516 200738 3568 200744
rect 3528 179489 3556 200738
rect 3606 200696 3662 200705
rect 3606 200631 3662 200640
rect 3514 179480 3570 179489
rect 3514 179415 3570 179424
rect 3620 136377 3648 200631
rect 3804 150793 3832 200767
rect 3988 165073 4016 201039
rect 4068 200864 4120 200870
rect 4068 200806 4120 200812
rect 4080 193905 4108 200806
rect 4066 193896 4122 193905
rect 4066 193831 4122 193840
rect 3974 165064 4030 165073
rect 3974 164999 4030 165008
rect 3790 150784 3846 150793
rect 3790 150719 3846 150728
rect 3606 136368 3662 136377
rect 3606 136303 3662 136312
rect 3422 122088 3478 122097
rect 3422 122023 3478 122032
rect 3240 108996 3292 109002
rect 3240 108938 3292 108944
rect 3252 107681 3280 108938
rect 3238 107672 3294 107681
rect 3238 107607 3294 107616
rect 3422 80064 3478 80073
rect 3422 79999 3478 80008
rect 3436 78985 3464 79999
rect 3422 78976 3478 78985
rect 3422 78911 3478 78920
rect 3330 50960 3386 50969
rect 3330 50895 3386 50904
rect 3344 50153 3372 50895
rect 3330 50144 3386 50153
rect 3330 50079 3386 50088
rect 3422 8256 3478 8265
rect 3422 8191 3478 8200
rect 3436 7177 3464 8191
rect 3422 7168 3478 7177
rect 3422 7103 3478 7112
rect 572 3528 624 3534
rect 572 3470 624 3476
rect 1308 3528 1360 3534
rect 1308 3470 1360 3476
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 2688 3528 2740 3534
rect 2688 3470 2740 3476
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 584 480 612 3470
rect 1688 480 1716 3470
rect 2884 480 2912 3470
rect 4068 3460 4120 3466
rect 4068 3402 4120 3408
rect 4080 480 4108 3402
rect 5460 610 5488 248406
rect 6840 626 6868 251194
rect 8220 3602 8248 252554
rect 9600 93498 9628 255274
rect 9588 93492 9640 93498
rect 9588 93434 9640 93440
rect 9588 93356 9640 93362
rect 9588 93298 9640 93304
rect 9600 3602 9628 93298
rect 10980 3602 11008 256702
rect 12360 3602 12388 259422
rect 13648 3602 13676 262210
rect 7656 3596 7708 3602
rect 7656 3538 7708 3544
rect 8208 3596 8260 3602
rect 8208 3538 8260 3544
rect 8852 3596 8904 3602
rect 8852 3538 8904 3544
rect 9588 3596 9640 3602
rect 9588 3538 9640 3544
rect 10048 3596 10100 3602
rect 10048 3538 10100 3544
rect 10968 3596 11020 3602
rect 10968 3538 11020 3544
rect 11244 3596 11296 3602
rect 11244 3538 11296 3544
rect 12348 3596 12400 3602
rect 12348 3538 12400 3544
rect 12440 3596 12492 3602
rect 12440 3538 12492 3544
rect 13636 3596 13688 3602
rect 13636 3538 13688 3544
rect 5264 604 5316 610
rect 5264 546 5316 552
rect 5448 604 5500 610
rect 5448 546 5500 552
rect 6472 598 6868 626
rect 5276 480 5304 546
rect 6472 480 6500 598
rect 7668 480 7696 3538
rect 8864 480 8892 3538
rect 10060 480 10088 3538
rect 11256 480 11284 3538
rect 12452 480 12480 3538
rect 13740 3482 13768 263570
rect 15120 3482 15148 266358
rect 16500 3602 16528 267718
rect 17880 3602 17908 270506
rect 19260 3602 19288 271866
rect 20640 3602 20668 274654
rect 21928 3602 21956 276014
rect 16028 3596 16080 3602
rect 16028 3538 16080 3544
rect 16488 3596 16540 3602
rect 16488 3538 16540 3544
rect 17224 3596 17276 3602
rect 17224 3538 17276 3544
rect 17868 3596 17920 3602
rect 17868 3538 17920 3544
rect 18328 3596 18380 3602
rect 18328 3538 18380 3544
rect 19248 3596 19300 3602
rect 19248 3538 19300 3544
rect 19524 3596 19576 3602
rect 19524 3538 19576 3544
rect 20628 3596 20680 3602
rect 20628 3538 20680 3544
rect 20720 3596 20772 3602
rect 20720 3538 20772 3544
rect 21916 3596 21968 3602
rect 21916 3538 21968 3544
rect 13648 3454 13768 3482
rect 14844 3454 15148 3482
rect 13648 480 13676 3454
rect 14844 480 14872 3454
rect 16040 480 16068 3538
rect 17236 480 17264 3538
rect 18340 480 18368 3538
rect 19536 480 19564 3538
rect 20732 480 20760 3538
rect 22020 3482 22048 278734
rect 23400 3482 23428 280162
rect 24780 3602 24808 282882
rect 26160 3602 26188 285670
rect 27540 3602 27568 287030
rect 28920 3602 28948 289818
rect 30208 3602 30236 291178
rect 24308 3596 24360 3602
rect 24308 3538 24360 3544
rect 24768 3596 24820 3602
rect 24768 3538 24820 3544
rect 25504 3596 25556 3602
rect 25504 3538 25556 3544
rect 26148 3596 26200 3602
rect 26148 3538 26200 3544
rect 26700 3596 26752 3602
rect 26700 3538 26752 3544
rect 27528 3596 27580 3602
rect 27528 3538 27580 3544
rect 27896 3596 27948 3602
rect 27896 3538 27948 3544
rect 28908 3596 28960 3602
rect 28908 3538 28960 3544
rect 29092 3596 29144 3602
rect 29092 3538 29144 3544
rect 30196 3596 30248 3602
rect 30196 3538 30248 3544
rect 21928 3454 22048 3482
rect 23124 3454 23428 3482
rect 21928 480 21956 3454
rect 23124 480 23152 3454
rect 24320 480 24348 3538
rect 25516 480 25544 3538
rect 26712 480 26740 3538
rect 27908 480 27936 3538
rect 29104 480 29132 3538
rect 30300 480 30328 293966
rect 31680 3482 31708 295326
rect 33060 3482 33088 298114
rect 34440 3602 34468 299474
rect 35820 3602 35848 302194
rect 37200 3602 37228 303622
rect 38488 3602 38516 306342
rect 33876 3596 33928 3602
rect 33876 3538 33928 3544
rect 34428 3596 34480 3602
rect 34428 3538 34480 3544
rect 34980 3596 35032 3602
rect 34980 3538 35032 3544
rect 35808 3596 35860 3602
rect 35808 3538 35860 3544
rect 36176 3596 36228 3602
rect 36176 3538 36228 3544
rect 37188 3596 37240 3602
rect 37188 3538 37240 3544
rect 37372 3596 37424 3602
rect 37372 3538 37424 3544
rect 38476 3596 38528 3602
rect 38476 3538 38528 3544
rect 31496 3454 31708 3482
rect 32692 3454 33088 3482
rect 31496 480 31524 3454
rect 32692 480 32720 3454
rect 33888 480 33916 3538
rect 34992 480 35020 3538
rect 36188 480 36216 3538
rect 37384 480 37412 3538
rect 38580 480 38608 307770
rect 38660 93560 38712 93566
rect 38658 93528 38660 93537
rect 38712 93528 38714 93537
rect 38658 93463 38714 93472
rect 39960 3482 39988 310490
rect 41340 3482 41368 313278
rect 42720 3602 42748 314638
rect 44100 3602 44128 317426
rect 45480 3602 45508 318786
rect 46860 3602 46888 321574
rect 48148 93786 48176 322934
rect 48056 93758 48176 93786
rect 48240 93770 48268 325654
rect 48228 93764 48280 93770
rect 48056 86986 48084 93758
rect 48228 93706 48280 93712
rect 48134 93664 48190 93673
rect 48134 93599 48190 93608
rect 48148 93566 48176 93599
rect 48136 93560 48188 93566
rect 48136 93502 48188 93508
rect 48228 93560 48280 93566
rect 48228 93502 48280 93508
rect 48056 86958 48176 86986
rect 48148 3602 48176 86958
rect 42156 3596 42208 3602
rect 42156 3538 42208 3544
rect 42708 3596 42760 3602
rect 42708 3538 42760 3544
rect 43352 3596 43404 3602
rect 43352 3538 43404 3544
rect 44088 3596 44140 3602
rect 44088 3538 44140 3544
rect 44548 3596 44600 3602
rect 44548 3538 44600 3544
rect 45468 3596 45520 3602
rect 45468 3538 45520 3544
rect 45744 3596 45796 3602
rect 45744 3538 45796 3544
rect 46848 3596 46900 3602
rect 46848 3538 46900 3544
rect 46940 3596 46992 3602
rect 46940 3538 46992 3544
rect 48136 3596 48188 3602
rect 48136 3538 48188 3544
rect 39776 3454 39988 3482
rect 40972 3454 41368 3482
rect 39776 480 39804 3454
rect 40972 480 41000 3454
rect 42168 480 42196 3538
rect 43364 480 43392 3538
rect 44560 480 44588 3538
rect 45756 480 45784 3538
rect 46952 480 46980 3538
rect 48240 3482 48268 93502
rect 49620 3482 49648 327082
rect 51000 3602 51028 329802
rect 52380 3602 52408 331230
rect 53760 3602 53788 333950
rect 55140 3602 55168 335310
rect 56428 3602 56456 338098
rect 50528 3596 50580 3602
rect 50528 3538 50580 3544
rect 50988 3596 51040 3602
rect 50988 3538 51040 3544
rect 51632 3596 51684 3602
rect 51632 3538 51684 3544
rect 52368 3596 52420 3602
rect 52368 3538 52420 3544
rect 52828 3596 52880 3602
rect 52828 3538 52880 3544
rect 53748 3596 53800 3602
rect 53748 3538 53800 3544
rect 54024 3596 54076 3602
rect 54024 3538 54076 3544
rect 55128 3596 55180 3602
rect 55128 3538 55180 3544
rect 55220 3596 55272 3602
rect 55220 3538 55272 3544
rect 56416 3596 56468 3602
rect 56416 3538 56468 3544
rect 48148 3454 48268 3482
rect 49344 3454 49648 3482
rect 48148 480 48176 3454
rect 49344 480 49372 3454
rect 50540 480 50568 3538
rect 51644 480 51672 3538
rect 52840 480 52868 3538
rect 54036 480 54064 3538
rect 55232 480 55260 3538
rect 56520 3482 56548 340886
rect 57900 3482 57928 342246
rect 59280 3602 59308 345034
rect 60660 3602 60688 346394
rect 62040 3602 62068 349114
rect 58808 3596 58860 3602
rect 58808 3538 58860 3544
rect 59268 3596 59320 3602
rect 59268 3538 59320 3544
rect 60004 3596 60056 3602
rect 60004 3538 60056 3544
rect 60648 3596 60700 3602
rect 60648 3538 60700 3544
rect 61200 3596 61252 3602
rect 61200 3538 61252 3544
rect 62028 3596 62080 3602
rect 62028 3538 62080 3544
rect 56428 3454 56548 3482
rect 57624 3454 57928 3482
rect 56428 480 56456 3454
rect 57624 480 57652 3454
rect 58820 480 58848 3538
rect 60016 480 60044 3538
rect 61212 480 61240 3538
rect 63420 3194 63448 350542
rect 64708 3602 64736 353262
rect 63592 3596 63644 3602
rect 63592 3538 63644 3544
rect 64696 3596 64748 3602
rect 64696 3538 64748 3544
rect 62396 3188 62448 3194
rect 62396 3130 62448 3136
rect 63408 3188 63460 3194
rect 63408 3130 63460 3136
rect 62408 480 62436 3130
rect 63604 480 63632 3538
rect 64800 480 64828 354690
rect 66180 3482 66208 357410
rect 67560 3482 67588 358770
rect 68940 3602 68968 361558
rect 70320 3602 70348 362918
rect 71700 3602 71728 365706
rect 72422 93936 72478 93945
rect 72422 93871 72478 93880
rect 72436 93673 72464 93871
rect 72422 93664 72478 93673
rect 72422 93599 72478 93608
rect 72988 3602 73016 368494
rect 68284 3596 68336 3602
rect 68284 3538 68336 3544
rect 68928 3596 68980 3602
rect 68928 3538 68980 3544
rect 69480 3596 69532 3602
rect 69480 3538 69532 3544
rect 70308 3596 70360 3602
rect 70308 3538 70360 3544
rect 70676 3596 70728 3602
rect 70676 3538 70728 3544
rect 71688 3596 71740 3602
rect 71688 3538 71740 3544
rect 71872 3596 71924 3602
rect 71872 3538 71924 3544
rect 72976 3596 73028 3602
rect 72976 3538 73028 3544
rect 65996 3454 66208 3482
rect 67192 3454 67588 3482
rect 65996 480 66024 3454
rect 67192 480 67220 3454
rect 68296 480 68324 3538
rect 69492 480 69520 3538
rect 70688 480 70716 3538
rect 71884 480 71912 3538
rect 73080 480 73108 369854
rect 74460 3482 74488 372574
rect 75840 3482 75868 374002
rect 77220 3602 77248 376722
rect 78600 3602 78628 378150
rect 79980 3602 80008 380870
rect 81360 3602 81388 382230
rect 82648 3602 82676 385018
rect 76656 3596 76708 3602
rect 76656 3538 76708 3544
rect 77208 3596 77260 3602
rect 77208 3538 77260 3544
rect 77852 3596 77904 3602
rect 77852 3538 77904 3544
rect 78588 3596 78640 3602
rect 78588 3538 78640 3544
rect 79048 3596 79100 3602
rect 79048 3538 79100 3544
rect 79968 3596 80020 3602
rect 79968 3538 80020 3544
rect 80244 3596 80296 3602
rect 80244 3538 80296 3544
rect 81348 3596 81400 3602
rect 81348 3538 81400 3544
rect 81440 3596 81492 3602
rect 81440 3538 81492 3544
rect 82636 3596 82688 3602
rect 82636 3538 82688 3544
rect 74276 3454 74488 3482
rect 75472 3454 75868 3482
rect 74276 480 74304 3454
rect 75472 480 75500 3454
rect 76668 480 76696 3538
rect 77864 480 77892 3538
rect 79060 480 79088 3538
rect 80256 480 80284 3538
rect 81452 480 81480 3538
rect 82740 3482 82768 386378
rect 84120 3482 84148 389166
rect 85500 3602 85528 390526
rect 86880 3602 86908 393314
rect 88260 3602 88288 396034
rect 89640 3602 89668 397462
rect 90928 3602 90956 400182
rect 84936 3596 84988 3602
rect 84936 3538 84988 3544
rect 85488 3596 85540 3602
rect 85488 3538 85540 3544
rect 86132 3596 86184 3602
rect 86132 3538 86184 3544
rect 86868 3596 86920 3602
rect 86868 3538 86920 3544
rect 87328 3596 87380 3602
rect 87328 3538 87380 3544
rect 88248 3596 88300 3602
rect 88248 3538 88300 3544
rect 88524 3596 88576 3602
rect 88524 3538 88576 3544
rect 89628 3596 89680 3602
rect 89628 3538 89680 3544
rect 89720 3596 89772 3602
rect 89720 3538 89772 3544
rect 90916 3596 90968 3602
rect 90916 3538 90968 3544
rect 82648 3454 82768 3482
rect 83844 3454 84148 3482
rect 82648 480 82676 3454
rect 83844 480 83872 3454
rect 84948 480 84976 3538
rect 86144 480 86172 3538
rect 87340 480 87368 3538
rect 88536 480 88564 3538
rect 89732 480 89760 3538
rect 91020 3482 91048 401610
rect 91742 93936 91798 93945
rect 91742 93871 91798 93880
rect 91756 93673 91784 93871
rect 91742 93664 91798 93673
rect 91742 93599 91798 93608
rect 92400 3482 92428 404330
rect 93780 3602 93808 405690
rect 95160 3602 95188 408478
rect 96540 3602 96568 409838
rect 97920 3602 97948 412626
rect 99208 3602 99236 413986
rect 93308 3596 93360 3602
rect 93308 3538 93360 3544
rect 93768 3596 93820 3602
rect 93768 3538 93820 3544
rect 94504 3596 94556 3602
rect 94504 3538 94556 3544
rect 95148 3596 95200 3602
rect 95148 3538 95200 3544
rect 95700 3596 95752 3602
rect 95700 3538 95752 3544
rect 96528 3596 96580 3602
rect 96528 3538 96580 3544
rect 96896 3596 96948 3602
rect 96896 3538 96948 3544
rect 97908 3596 97960 3602
rect 97908 3538 97960 3544
rect 98092 3596 98144 3602
rect 98092 3538 98144 3544
rect 99196 3596 99248 3602
rect 99196 3538 99248 3544
rect 90928 3454 91048 3482
rect 92124 3454 92428 3482
rect 90928 480 90956 3454
rect 92124 480 92152 3454
rect 93320 480 93348 3538
rect 94516 480 94544 3538
rect 95712 480 95740 3538
rect 96908 480 96936 3538
rect 98104 480 98132 3538
rect 99300 480 99328 416774
rect 100680 3482 100708 418134
rect 100496 3454 100708 3482
rect 100496 480 100524 3454
rect 102060 3330 102088 420922
rect 103440 3602 103468 423642
rect 104820 3602 104848 425070
rect 106200 3602 106228 427790
rect 107488 3602 107516 429150
rect 102784 3596 102836 3602
rect 102784 3538 102836 3544
rect 103428 3596 103480 3602
rect 103428 3538 103480 3544
rect 103980 3596 104032 3602
rect 103980 3538 104032 3544
rect 104808 3596 104860 3602
rect 104808 3538 104860 3544
rect 105176 3596 105228 3602
rect 105176 3538 105228 3544
rect 106188 3596 106240 3602
rect 106188 3538 106240 3544
rect 106372 3596 106424 3602
rect 106372 3538 106424 3544
rect 107476 3596 107528 3602
rect 107476 3538 107528 3544
rect 101588 3324 101640 3330
rect 101588 3266 101640 3272
rect 102048 3324 102100 3330
rect 102048 3266 102100 3272
rect 101600 480 101628 3266
rect 102796 480 102824 3538
rect 103992 480 104020 3538
rect 105188 480 105216 3538
rect 106384 480 106412 3538
rect 107580 480 107608 431938
rect 108960 3482 108988 433298
rect 110340 3482 110368 436086
rect 111062 93936 111118 93945
rect 111062 93871 111118 93880
rect 111076 93673 111104 93871
rect 111062 93664 111118 93673
rect 111062 93599 111118 93608
rect 111720 3602 111748 437446
rect 113100 3602 113128 440234
rect 114480 3602 114508 441594
rect 115860 3602 115888 444382
rect 117148 3602 117176 445742
rect 111156 3596 111208 3602
rect 111156 3538 111208 3544
rect 111708 3596 111760 3602
rect 111708 3538 111760 3544
rect 112352 3596 112404 3602
rect 112352 3538 112404 3544
rect 113088 3596 113140 3602
rect 113088 3538 113140 3544
rect 113548 3596 113600 3602
rect 113548 3538 113600 3544
rect 114468 3596 114520 3602
rect 114468 3538 114520 3544
rect 114744 3596 114796 3602
rect 114744 3538 114796 3544
rect 115848 3596 115900 3602
rect 115848 3538 115900 3544
rect 115940 3596 115992 3602
rect 115940 3538 115992 3544
rect 117136 3596 117188 3602
rect 117136 3538 117188 3544
rect 108776 3454 108988 3482
rect 109972 3454 110368 3482
rect 108776 480 108804 3454
rect 109972 480 110000 3454
rect 111168 480 111196 3538
rect 112364 480 112392 3538
rect 113560 480 113588 3538
rect 114756 480 114784 3538
rect 115952 480 115980 3538
rect 117240 3482 117268 448530
rect 118620 3482 118648 451250
rect 120000 3602 120028 452610
rect 121380 3602 121408 455398
rect 122760 3602 122788 456758
rect 124140 3602 124168 459546
rect 125428 3602 125456 460906
rect 119436 3596 119488 3602
rect 119436 3538 119488 3544
rect 119988 3596 120040 3602
rect 119988 3538 120040 3544
rect 120632 3596 120684 3602
rect 120632 3538 120684 3544
rect 121368 3596 121420 3602
rect 121368 3538 121420 3544
rect 121828 3596 121880 3602
rect 121828 3538 121880 3544
rect 122748 3596 122800 3602
rect 122748 3538 122800 3544
rect 123024 3596 123076 3602
rect 123024 3538 123076 3544
rect 124128 3596 124180 3602
rect 124128 3538 124180 3544
rect 124220 3596 124272 3602
rect 124220 3538 124272 3544
rect 125416 3596 125468 3602
rect 125416 3538 125468 3544
rect 117148 3454 117268 3482
rect 118252 3454 118648 3482
rect 117148 480 117176 3454
rect 118252 480 118280 3454
rect 119448 480 119476 3538
rect 120644 480 120672 3538
rect 121840 480 121868 3538
rect 123036 480 123064 3538
rect 124232 480 124260 3538
rect 125520 3482 125548 463694
rect 126900 3482 126928 465054
rect 128280 3602 128308 467842
rect 129660 3602 129688 469202
rect 130382 93936 130438 93945
rect 130382 93871 130438 93880
rect 130396 93673 130424 93871
rect 130382 93664 130438 93673
rect 130382 93599 130438 93608
rect 131040 3602 131068 471990
rect 132420 3602 132448 473350
rect 133800 3602 133828 476070
rect 127808 3596 127860 3602
rect 127808 3538 127860 3544
rect 128268 3596 128320 3602
rect 128268 3538 128320 3544
rect 129004 3596 129056 3602
rect 129004 3538 129056 3544
rect 129648 3596 129700 3602
rect 129648 3538 129700 3544
rect 130200 3596 130252 3602
rect 130200 3538 130252 3544
rect 131028 3596 131080 3602
rect 131028 3538 131080 3544
rect 131396 3596 131448 3602
rect 131396 3538 131448 3544
rect 132408 3596 132460 3602
rect 132408 3538 132460 3544
rect 132592 3596 132644 3602
rect 132592 3538 132644 3544
rect 133788 3596 133840 3602
rect 133788 3538 133840 3544
rect 125428 3454 125548 3482
rect 126624 3454 126928 3482
rect 125428 480 125456 3454
rect 126624 480 126652 3454
rect 127820 480 127848 3538
rect 129016 480 129044 3538
rect 130212 480 130240 3538
rect 131408 480 131436 3538
rect 132604 480 132632 3538
rect 135180 626 135208 478858
rect 259828 478576 259880 478582
rect 259828 478518 259880 478524
rect 256698 476776 256754 476785
rect 256698 476711 256754 476720
rect 256712 476134 256740 476711
rect 256700 476128 256752 476134
rect 256700 476070 256752 476076
rect 256698 474736 256754 474745
rect 256698 474671 256754 474680
rect 256712 473414 256740 474671
rect 256700 473408 256752 473414
rect 256700 473350 256752 473356
rect 256698 472560 256754 472569
rect 256698 472495 256754 472504
rect 256712 472054 256740 472495
rect 256700 472048 256752 472054
rect 256700 471990 256752 471996
rect 256698 470384 256754 470393
rect 256698 470319 256754 470328
rect 256712 469266 256740 470319
rect 256700 469260 256752 469266
rect 256700 469202 256752 469208
rect 256698 468344 256754 468353
rect 256698 468279 256754 468288
rect 256712 467906 256740 468279
rect 256700 467900 256752 467906
rect 256700 467842 256752 467848
rect 256698 466168 256754 466177
rect 256698 466103 256754 466112
rect 256712 465118 256740 466103
rect 256700 465112 256752 465118
rect 256700 465054 256752 465060
rect 256698 464128 256754 464137
rect 256698 464063 256754 464072
rect 256712 463758 256740 464063
rect 256700 463752 256752 463758
rect 256700 463694 256752 463700
rect 256698 461952 256754 461961
rect 256698 461887 256754 461896
rect 256712 460970 256740 461887
rect 256700 460964 256752 460970
rect 256700 460906 256752 460912
rect 256698 459776 256754 459785
rect 256698 459711 256754 459720
rect 256712 459610 256740 459711
rect 256700 459604 256752 459610
rect 256700 459546 256752 459552
rect 256698 457736 256754 457745
rect 256698 457671 256754 457680
rect 256712 456822 256740 457671
rect 256700 456816 256752 456822
rect 256700 456758 256752 456764
rect 256698 455560 256754 455569
rect 256698 455495 256754 455504
rect 256712 455462 256740 455495
rect 256700 455456 256752 455462
rect 256700 455398 256752 455404
rect 256698 453384 256754 453393
rect 256698 453319 256754 453328
rect 256712 452674 256740 453319
rect 256700 452668 256752 452674
rect 256700 452610 256752 452616
rect 259840 452606 259868 478518
rect 259828 452600 259880 452606
rect 259828 452542 259880 452548
rect 256698 451344 256754 451353
rect 256698 451279 256700 451288
rect 256752 451279 256754 451288
rect 256700 451250 256752 451256
rect 256698 449168 256754 449177
rect 256698 449103 256754 449112
rect 256712 448594 256740 449103
rect 256700 448588 256752 448594
rect 256700 448530 256752 448536
rect 256698 447128 256754 447137
rect 256698 447063 256754 447072
rect 256712 445806 256740 447063
rect 256700 445800 256752 445806
rect 256700 445742 256752 445748
rect 256698 444952 256754 444961
rect 256698 444887 256754 444896
rect 256712 444446 256740 444887
rect 256700 444440 256752 444446
rect 256700 444382 256752 444388
rect 256698 442776 256754 442785
rect 256698 442711 256754 442720
rect 256712 441658 256740 442711
rect 256700 441652 256752 441658
rect 256700 441594 256752 441600
rect 256698 440736 256754 440745
rect 256698 440671 256754 440680
rect 256712 440298 256740 440671
rect 256700 440292 256752 440298
rect 256700 440234 256752 440240
rect 259932 438870 259960 478858
rect 260012 478100 260064 478106
rect 260012 478042 260064 478048
rect 259920 438864 259972 438870
rect 259920 438806 259972 438812
rect 256698 438560 256754 438569
rect 256698 438495 256754 438504
rect 256712 437510 256740 438495
rect 256700 437504 256752 437510
rect 256700 437446 256752 437452
rect 256698 436384 256754 436393
rect 256698 436319 256754 436328
rect 256712 436150 256740 436319
rect 256700 436144 256752 436150
rect 256700 436086 256752 436092
rect 256698 434344 256754 434353
rect 256698 434279 256754 434288
rect 256712 433362 256740 434279
rect 256700 433356 256752 433362
rect 256700 433298 256752 433304
rect 256698 432168 256754 432177
rect 256698 432103 256754 432112
rect 256712 432002 256740 432103
rect 256700 431996 256752 432002
rect 256700 431938 256752 431944
rect 256698 430128 256754 430137
rect 256698 430063 256754 430072
rect 256712 429214 256740 430063
rect 256700 429208 256752 429214
rect 256700 429150 256752 429156
rect 256698 427952 256754 427961
rect 256698 427887 256754 427896
rect 256712 427854 256740 427887
rect 256700 427848 256752 427854
rect 256700 427790 256752 427796
rect 256698 425776 256754 425785
rect 256698 425711 256754 425720
rect 256712 425134 256740 425711
rect 256700 425128 256752 425134
rect 256700 425070 256752 425076
rect 260024 425066 260052 478042
rect 260012 425060 260064 425066
rect 260012 425002 260064 425008
rect 256698 423736 256754 423745
rect 256698 423671 256700 423680
rect 256752 423671 256754 423680
rect 256700 423642 256752 423648
rect 256698 421560 256754 421569
rect 256698 421495 256754 421504
rect 256712 420986 256740 421495
rect 256700 420980 256752 420986
rect 256700 420922 256752 420928
rect 256698 419520 256754 419529
rect 256698 419455 256754 419464
rect 256712 418198 256740 419455
rect 256700 418192 256752 418198
rect 256700 418134 256752 418140
rect 256698 417344 256754 417353
rect 256698 417279 256754 417288
rect 256712 416838 256740 417279
rect 256700 416832 256752 416838
rect 256700 416774 256752 416780
rect 256698 415168 256754 415177
rect 256698 415103 256754 415112
rect 256712 414050 256740 415103
rect 256700 414044 256752 414050
rect 256700 413986 256752 413992
rect 256698 413128 256754 413137
rect 256698 413063 256754 413072
rect 256712 412690 256740 413063
rect 256700 412684 256752 412690
rect 256700 412626 256752 412632
rect 256698 410952 256754 410961
rect 256698 410887 256754 410896
rect 256712 409902 256740 410887
rect 256700 409896 256752 409902
rect 256700 409838 256752 409844
rect 256698 408776 256754 408785
rect 256698 408711 256754 408720
rect 256712 408542 256740 408711
rect 256700 408536 256752 408542
rect 256700 408478 256752 408484
rect 256698 406736 256754 406745
rect 256698 406671 256754 406680
rect 256712 405754 256740 406671
rect 256700 405748 256752 405754
rect 256700 405690 256752 405696
rect 256698 404560 256754 404569
rect 256698 404495 256754 404504
rect 256712 404394 256740 404495
rect 256700 404388 256752 404394
rect 256700 404330 256752 404336
rect 256698 402520 256754 402529
rect 256698 402455 256754 402464
rect 256712 401674 256740 402455
rect 256700 401668 256752 401674
rect 256700 401610 256752 401616
rect 256698 400344 256754 400353
rect 256698 400279 256754 400288
rect 256712 400246 256740 400279
rect 256700 400240 256752 400246
rect 256700 400182 256752 400188
rect 256698 398168 256754 398177
rect 256698 398103 256754 398112
rect 256712 397526 256740 398103
rect 256700 397520 256752 397526
rect 256700 397462 256752 397468
rect 256698 396128 256754 396137
rect 256698 396063 256700 396072
rect 256752 396063 256754 396072
rect 256700 396034 256752 396040
rect 256698 393952 256754 393961
rect 256698 393887 256754 393896
rect 256712 393378 256740 393887
rect 256700 393372 256752 393378
rect 256700 393314 256752 393320
rect 256698 391776 256754 391785
rect 256698 391711 256754 391720
rect 256712 390590 256740 391711
rect 256700 390584 256752 390590
rect 256700 390526 256752 390532
rect 256698 389736 256754 389745
rect 256698 389671 256754 389680
rect 256712 389230 256740 389671
rect 256700 389224 256752 389230
rect 256700 389166 256752 389172
rect 256698 387560 256754 387569
rect 256698 387495 256754 387504
rect 256712 386442 256740 387495
rect 256700 386436 256752 386442
rect 256700 386378 256752 386384
rect 256698 385520 256754 385529
rect 256698 385455 256754 385464
rect 256712 385082 256740 385455
rect 256700 385076 256752 385082
rect 256700 385018 256752 385024
rect 256698 383344 256754 383353
rect 256698 383279 256754 383288
rect 256712 382294 256740 383279
rect 256700 382288 256752 382294
rect 256700 382230 256752 382236
rect 256698 381168 256754 381177
rect 256698 381103 256754 381112
rect 256712 380934 256740 381103
rect 256700 380928 256752 380934
rect 256700 380870 256752 380876
rect 256698 379128 256754 379137
rect 256698 379063 256754 379072
rect 256712 378214 256740 379063
rect 256700 378208 256752 378214
rect 256700 378150 256752 378156
rect 256698 376952 256754 376961
rect 256698 376887 256754 376896
rect 256712 376786 256740 376887
rect 256700 376780 256752 376786
rect 256700 376722 256752 376728
rect 256698 374912 256754 374921
rect 256698 374847 256754 374856
rect 256712 374066 256740 374847
rect 256700 374060 256752 374066
rect 256700 374002 256752 374008
rect 256698 372736 256754 372745
rect 256698 372671 256754 372680
rect 256712 372638 256740 372671
rect 256700 372632 256752 372638
rect 256700 372574 256752 372580
rect 256698 370560 256754 370569
rect 256698 370495 256754 370504
rect 256712 369918 256740 370495
rect 256700 369912 256752 369918
rect 256700 369854 256752 369860
rect 256700 368552 256752 368558
rect 256698 368520 256700 368529
rect 256752 368520 256754 368529
rect 256698 368455 256754 368464
rect 256698 366344 256754 366353
rect 256698 366279 256754 366288
rect 256712 365770 256740 366279
rect 256700 365764 256752 365770
rect 256700 365706 256752 365712
rect 256698 364168 256754 364177
rect 256698 364103 256754 364112
rect 256712 362982 256740 364103
rect 256700 362976 256752 362982
rect 256700 362918 256752 362924
rect 256698 362128 256754 362137
rect 256698 362063 256754 362072
rect 256712 361622 256740 362063
rect 256700 361616 256752 361622
rect 256700 361558 256752 361564
rect 256698 359952 256754 359961
rect 256698 359887 256754 359896
rect 256712 358834 256740 359887
rect 256700 358828 256752 358834
rect 256700 358770 256752 358776
rect 256698 357912 256754 357921
rect 256698 357847 256754 357856
rect 256712 357474 256740 357847
rect 256700 357468 256752 357474
rect 256700 357410 256752 357416
rect 256698 355736 256754 355745
rect 256698 355671 256754 355680
rect 256712 354754 256740 355671
rect 256700 354748 256752 354754
rect 256700 354690 256752 354696
rect 256698 353560 256754 353569
rect 256698 353495 256754 353504
rect 256712 353326 256740 353495
rect 256700 353320 256752 353326
rect 256700 353262 256752 353268
rect 256698 351520 256754 351529
rect 256698 351455 256754 351464
rect 256712 350606 256740 351455
rect 256700 350600 256752 350606
rect 256700 350542 256752 350548
rect 256698 349344 256754 349353
rect 256698 349279 256754 349288
rect 256712 349178 256740 349279
rect 256700 349172 256752 349178
rect 256700 349114 256752 349120
rect 256698 347168 256754 347177
rect 256698 347103 256754 347112
rect 256712 346458 256740 347103
rect 256700 346452 256752 346458
rect 256700 346394 256752 346400
rect 256698 345128 256754 345137
rect 256698 345063 256700 345072
rect 256752 345063 256754 345072
rect 256700 345034 256752 345040
rect 256698 342952 256754 342961
rect 256698 342887 256754 342896
rect 256712 342310 256740 342887
rect 256700 342304 256752 342310
rect 256700 342246 256752 342252
rect 256700 340944 256752 340950
rect 256698 340912 256700 340921
rect 256752 340912 256754 340921
rect 256698 340847 256754 340856
rect 256698 338736 256754 338745
rect 256698 338671 256754 338680
rect 256712 338162 256740 338671
rect 256700 338156 256752 338162
rect 256700 338098 256752 338104
rect 256698 336560 256754 336569
rect 256698 336495 256754 336504
rect 256712 335374 256740 336495
rect 256700 335368 256752 335374
rect 256700 335310 256752 335316
rect 256698 334520 256754 334529
rect 256698 334455 256754 334464
rect 256712 334014 256740 334455
rect 256700 334008 256752 334014
rect 256700 333950 256752 333956
rect 256698 332344 256754 332353
rect 256698 332279 256754 332288
rect 256712 331294 256740 332279
rect 256700 331288 256752 331294
rect 256700 331230 256752 331236
rect 256698 330304 256754 330313
rect 256698 330239 256754 330248
rect 256712 329866 256740 330239
rect 256700 329860 256752 329866
rect 256700 329802 256752 329808
rect 256698 328128 256754 328137
rect 256698 328063 256754 328072
rect 256712 327146 256740 328063
rect 256700 327140 256752 327146
rect 256700 327082 256752 327088
rect 256698 325952 256754 325961
rect 256698 325887 256754 325896
rect 256712 325718 256740 325887
rect 256700 325712 256752 325718
rect 256700 325654 256752 325660
rect 256698 323912 256754 323921
rect 256698 323847 256754 323856
rect 256712 322998 256740 323847
rect 256700 322992 256752 322998
rect 256700 322934 256752 322940
rect 256698 321736 256754 321745
rect 256698 321671 256754 321680
rect 256712 321638 256740 321671
rect 256700 321632 256752 321638
rect 256700 321574 256752 321580
rect 256698 319560 256754 319569
rect 256698 319495 256754 319504
rect 256712 318850 256740 319495
rect 256700 318844 256752 318850
rect 256700 318786 256752 318792
rect 256698 317520 256754 317529
rect 256698 317455 256700 317464
rect 256752 317455 256754 317464
rect 256700 317426 256752 317432
rect 256698 315344 256754 315353
rect 256698 315279 256754 315288
rect 256712 314702 256740 315279
rect 256700 314696 256752 314702
rect 256700 314638 256752 314644
rect 256700 313336 256752 313342
rect 256698 313304 256700 313313
rect 256752 313304 256754 313313
rect 256698 313239 256754 313248
rect 256698 311128 256754 311137
rect 256698 311063 256754 311072
rect 256712 310554 256740 311063
rect 256700 310548 256752 310554
rect 256700 310490 256752 310496
rect 256698 308952 256754 308961
rect 256698 308887 256754 308896
rect 256712 307834 256740 308887
rect 256700 307828 256752 307834
rect 256700 307770 256752 307776
rect 256698 306912 256754 306921
rect 256698 306847 256754 306856
rect 256712 306406 256740 306847
rect 256700 306400 256752 306406
rect 256700 306342 256752 306348
rect 256698 304736 256754 304745
rect 256698 304671 256754 304680
rect 256712 303686 256740 304671
rect 256700 303680 256752 303686
rect 256700 303622 256752 303628
rect 256698 302560 256754 302569
rect 256698 302495 256754 302504
rect 256712 302258 256740 302495
rect 256700 302252 256752 302258
rect 256700 302194 256752 302200
rect 256698 300520 256754 300529
rect 256698 300455 256754 300464
rect 256712 299538 256740 300455
rect 256700 299532 256752 299538
rect 256700 299474 256752 299480
rect 256698 298344 256754 298353
rect 256698 298279 256754 298288
rect 256712 298178 256740 298279
rect 256700 298172 256752 298178
rect 256700 298114 256752 298120
rect 256698 296304 256754 296313
rect 256698 296239 256754 296248
rect 256712 295390 256740 296239
rect 256700 295384 256752 295390
rect 256700 295326 256752 295332
rect 256698 294128 256754 294137
rect 256698 294063 256754 294072
rect 256712 294030 256740 294063
rect 256700 294024 256752 294030
rect 256700 293966 256752 293972
rect 256698 291952 256754 291961
rect 256698 291887 256754 291896
rect 256712 291242 256740 291887
rect 256700 291236 256752 291242
rect 256700 291178 256752 291184
rect 256698 289912 256754 289921
rect 256698 289847 256700 289856
rect 256752 289847 256754 289856
rect 256700 289818 256752 289824
rect 256698 287736 256754 287745
rect 256698 287671 256754 287680
rect 256712 287094 256740 287671
rect 256700 287088 256752 287094
rect 256700 287030 256752 287036
rect 256700 285728 256752 285734
rect 256698 285696 256700 285705
rect 256752 285696 256754 285705
rect 256698 285631 256754 285640
rect 256698 283520 256754 283529
rect 256698 283455 256754 283464
rect 256712 282946 256740 283455
rect 256700 282940 256752 282946
rect 256700 282882 256752 282888
rect 256698 281344 256754 281353
rect 256698 281279 256754 281288
rect 256712 280226 256740 281279
rect 256700 280220 256752 280226
rect 256700 280162 256752 280168
rect 260116 280158 260144 478926
rect 260288 478372 260340 478378
rect 260288 478314 260340 478320
rect 260196 478032 260248 478038
rect 260196 477974 260248 477980
rect 260208 295322 260236 477974
rect 260300 309126 260328 478314
rect 260392 324290 260420 478994
rect 260472 478440 260524 478446
rect 260472 478382 260524 478388
rect 260484 338094 260512 478382
rect 260576 367062 260604 479062
rect 260668 380866 260696 479130
rect 260748 478508 260800 478514
rect 260748 478450 260800 478456
rect 260760 396030 260788 478450
rect 260748 396024 260800 396030
rect 260748 395966 260800 395972
rect 260656 380860 260708 380866
rect 260656 380802 260708 380808
rect 260564 367056 260616 367062
rect 260564 366998 260616 367004
rect 260472 338088 260524 338094
rect 260472 338030 260524 338036
rect 260380 324284 260432 324290
rect 260380 324226 260432 324232
rect 260288 309120 260340 309126
rect 260288 309062 260340 309068
rect 260196 295316 260248 295322
rect 260196 295258 260248 295264
rect 260104 280152 260156 280158
rect 260104 280094 260156 280100
rect 256698 279304 256754 279313
rect 256698 279239 256754 279248
rect 256712 278798 256740 279239
rect 256700 278792 256752 278798
rect 256700 278734 256752 278740
rect 256698 277128 256754 277137
rect 256698 277063 256754 277072
rect 256712 276078 256740 277063
rect 256700 276072 256752 276078
rect 256700 276014 256752 276020
rect 256698 274952 256754 274961
rect 256698 274887 256754 274896
rect 256712 274718 256740 274887
rect 256700 274712 256752 274718
rect 256700 274654 256752 274660
rect 256698 272912 256754 272921
rect 256698 272847 256754 272856
rect 256712 271930 256740 272847
rect 256700 271924 256752 271930
rect 256700 271866 256752 271872
rect 256698 270736 256754 270745
rect 256698 270671 256754 270680
rect 256712 270570 256740 270671
rect 256700 270564 256752 270570
rect 256700 270506 256752 270512
rect 256698 268696 256754 268705
rect 256698 268631 256754 268640
rect 256712 267782 256740 268631
rect 256700 267776 256752 267782
rect 256700 267718 256752 267724
rect 256698 266520 256754 266529
rect 256698 266455 256754 266464
rect 256712 266422 256740 266455
rect 256700 266416 256752 266422
rect 256700 266358 256752 266364
rect 256698 264344 256754 264353
rect 256698 264279 256754 264288
rect 256712 263634 256740 264279
rect 256700 263628 256752 263634
rect 256700 263570 256752 263576
rect 256698 262304 256754 262313
rect 256698 262239 256700 262248
rect 256752 262239 256754 262248
rect 256700 262210 256752 262216
rect 256698 260128 256754 260137
rect 256698 260063 256754 260072
rect 256712 259486 256740 260063
rect 256700 259480 256752 259486
rect 256700 259422 256752 259428
rect 256698 257952 256754 257961
rect 256698 257887 256754 257896
rect 256712 256766 256740 257887
rect 256700 256760 256752 256766
rect 256700 256702 256752 256708
rect 256698 255912 256754 255921
rect 256698 255847 256754 255856
rect 256712 255338 256740 255847
rect 256700 255332 256752 255338
rect 256700 255274 256752 255280
rect 256698 253736 256754 253745
rect 256698 253671 256754 253680
rect 256712 252618 256740 253671
rect 256700 252612 256752 252618
rect 256700 252554 256752 252560
rect 256698 251696 256754 251705
rect 256698 251631 256754 251640
rect 256712 251258 256740 251631
rect 256700 251252 256752 251258
rect 256700 251194 256752 251200
rect 256698 249520 256754 249529
rect 256698 249455 256754 249464
rect 256712 248470 256740 249455
rect 256700 248464 256752 248470
rect 256700 248406 256752 248412
rect 257342 247344 257398 247353
rect 257342 247279 257398 247288
rect 256974 243128 257030 243137
rect 256974 243063 257030 243072
rect 256988 242962 257016 243063
rect 256976 242956 257028 242962
rect 256976 242898 257028 242904
rect 154486 93800 154542 93809
rect 154486 93735 154542 93744
rect 154500 93702 154528 93735
rect 144920 93696 144972 93702
rect 140042 93664 140098 93673
rect 140042 93599 140098 93608
rect 144918 93664 144920 93673
rect 154488 93696 154540 93702
rect 144972 93664 144974 93673
rect 154488 93638 154540 93644
rect 144918 93599 144974 93608
rect 140056 93265 140084 93599
rect 140042 93256 140098 93265
rect 140042 93191 140098 93200
rect 257356 3466 257384 247279
rect 257434 245304 257490 245313
rect 257434 245239 257490 245248
rect 257448 3534 257476 245239
rect 257986 241088 258042 241097
rect 257986 241023 258042 241032
rect 258000 240582 258028 241023
rect 257988 240576 258040 240582
rect 257988 240518 258040 240524
rect 260840 240576 260892 240582
rect 260840 240518 260892 240524
rect 258000 240174 258028 240518
rect 260852 240446 260880 240518
rect 261128 240446 261156 517618
rect 266268 517540 266320 517546
rect 266268 517482 266320 517488
rect 261208 482316 261260 482322
rect 261208 482258 261260 482264
rect 261220 479876 261248 482258
rect 263690 482216 263746 482225
rect 263690 482151 263746 482160
rect 263704 479876 263732 482151
rect 266280 479876 266308 517482
rect 269040 479890 269068 518230
rect 271800 479890 271828 518298
rect 268870 479862 269068 479890
rect 271446 479862 271828 479890
rect 274560 479754 274588 518434
rect 286968 518152 287020 518158
rect 286968 518094 287020 518100
rect 285588 518084 285640 518090
rect 285588 518026 285640 518032
rect 282828 518016 282880 518022
rect 282828 517958 282880 517964
rect 280068 517948 280120 517954
rect 280068 517890 280120 517896
rect 277308 517880 277360 517886
rect 277308 517822 277360 517828
rect 277320 482050 277348 517822
rect 280080 482594 280108 517890
rect 282840 483002 282868 517958
rect 281724 482996 281776 483002
rect 281724 482938 281776 482944
rect 282828 482996 282880 483002
rect 282828 482938 282880 482944
rect 279148 482588 279200 482594
rect 279148 482530 279200 482536
rect 280068 482588 280120 482594
rect 280068 482530 280120 482536
rect 276572 482044 276624 482050
rect 276572 481986 276624 481992
rect 277308 482044 277360 482050
rect 277308 481986 277360 481992
rect 276584 479876 276612 481986
rect 279160 479876 279188 482530
rect 281736 479876 281764 482938
rect 285600 482730 285628 518026
rect 284300 482724 284352 482730
rect 284300 482666 284352 482672
rect 285588 482724 285640 482730
rect 285588 482666 285640 482672
rect 284312 479876 284340 482666
rect 286980 479890 287008 518094
rect 289740 479890 289768 518774
rect 297376 482390 297404 540223
rect 297468 482866 297496 598023
rect 297456 482860 297508 482866
rect 297456 482802 297508 482808
rect 297560 482798 297588 599791
rect 297548 482792 297600 482798
rect 297548 482734 297600 482740
rect 297652 482730 297680 600879
rect 297640 482724 297692 482730
rect 297640 482666 297692 482672
rect 297744 482662 297772 602511
rect 297732 482656 297784 482662
rect 297732 482598 297784 482604
rect 297836 482594 297864 603735
rect 297824 482588 297876 482594
rect 297824 482530 297876 482536
rect 297928 482526 297956 605367
rect 297916 482520 297968 482526
rect 297916 482462 297968 482468
rect 298020 482458 298048 606591
rect 298008 482452 298060 482458
rect 298008 482394 298060 482400
rect 297364 482384 297416 482390
rect 297364 482326 297416 482332
rect 292028 482044 292080 482050
rect 292028 481986 292080 481992
rect 286902 479862 287008 479890
rect 289478 479862 289768 479890
rect 292040 479876 292068 481986
rect 294512 481976 294564 481982
rect 294512 481918 294564 481924
rect 294524 479876 294552 481918
rect 297088 481908 297140 481914
rect 297088 481850 297140 481856
rect 297100 479876 297128 481850
rect 299664 481840 299716 481846
rect 299664 481782 299716 481788
rect 299676 479876 299704 481782
rect 300780 479806 300808 699654
rect 365640 610638 365668 699654
rect 373632 612808 373684 612814
rect 373630 612776 373632 612785
rect 379612 612808 379664 612814
rect 373684 612776 373686 612785
rect 379612 612750 379664 612756
rect 373630 612711 373686 612720
rect 365628 610632 365680 610638
rect 365628 610574 365680 610580
rect 379428 601724 379480 601730
rect 379428 601666 379480 601672
rect 378048 600364 378100 600370
rect 378048 600306 378100 600312
rect 320088 518900 320140 518906
rect 328920 518900 328972 518906
rect 320088 518842 320140 518848
rect 320100 518809 320128 518842
rect 327368 518838 327396 518869
rect 328920 518842 328972 518848
rect 329656 518900 329708 518906
rect 329656 518842 329708 518848
rect 348976 518900 349028 518906
rect 348976 518842 349028 518848
rect 322940 518832 322992 518838
rect 314566 518800 314622 518809
rect 307668 518764 307720 518770
rect 314566 518735 314622 518744
rect 320086 518800 320142 518809
rect 320086 518735 320142 518744
rect 322938 518800 322940 518809
rect 327356 518832 327408 518838
rect 322992 518800 322994 518809
rect 322938 518735 322994 518744
rect 324318 518800 324374 518809
rect 324318 518735 324374 518744
rect 325422 518800 325478 518809
rect 325422 518735 325478 518744
rect 326434 518800 326490 518809
rect 326434 518735 326490 518744
rect 327354 518800 327356 518809
rect 328932 518809 328960 518842
rect 327408 518800 327410 518809
rect 327354 518735 327410 518744
rect 328918 518800 328974 518809
rect 328918 518735 328974 518744
rect 307668 518706 307720 518712
rect 303618 518256 303674 518265
rect 303618 518191 303620 518200
rect 303672 518191 303674 518200
rect 303620 518162 303672 518168
rect 303632 517682 303660 518162
rect 303620 517676 303672 517682
rect 303620 517618 303672 517624
rect 304908 517676 304960 517682
rect 304908 517618 304960 517624
rect 302240 481772 302292 481778
rect 302240 481714 302292 481720
rect 302252 479876 302280 481714
rect 304920 479890 304948 517618
rect 307574 517576 307630 517585
rect 307574 517511 307630 517520
rect 307588 482934 307616 517511
rect 307576 482928 307628 482934
rect 307576 482870 307628 482876
rect 307680 479890 307708 518706
rect 314580 518702 314608 518735
rect 314568 518696 314620 518702
rect 313186 518664 313242 518673
rect 323124 518696 323176 518702
rect 314568 518638 314620 518644
rect 317234 518664 317290 518673
rect 313186 518599 313242 518608
rect 317234 518599 317290 518608
rect 318706 518664 318762 518673
rect 318706 518599 318708 518608
rect 313200 518430 313228 518599
rect 314658 518528 314714 518537
rect 314658 518463 314714 518472
rect 316038 518528 316094 518537
rect 316038 518463 316040 518472
rect 313188 518424 313240 518430
rect 313188 518366 313240 518372
rect 313278 518392 313334 518401
rect 314672 518362 314700 518463
rect 316092 518463 316094 518472
rect 316040 518434 316092 518440
rect 317248 518430 317276 518599
rect 318760 518599 318762 518608
rect 321098 518664 321154 518673
rect 321098 518599 321154 518608
rect 323122 518664 323124 518673
rect 323176 518664 323178 518673
rect 323122 518599 323178 518608
rect 318708 518570 318760 518576
rect 321112 518566 321140 518599
rect 321100 518560 321152 518566
rect 317326 518528 317382 518537
rect 317326 518463 317328 518472
rect 317380 518463 317382 518472
rect 317510 518528 317566 518537
rect 321100 518502 321152 518508
rect 317510 518463 317566 518472
rect 317328 518434 317380 518440
rect 317236 518424 317288 518430
rect 317236 518366 317288 518372
rect 313278 518327 313334 518336
rect 314660 518356 314712 518362
rect 313292 518294 313320 518327
rect 314660 518298 314712 518304
rect 313280 518288 313332 518294
rect 313280 518230 313332 518236
rect 315856 518288 315908 518294
rect 315856 518230 315908 518236
rect 315868 518090 315896 518230
rect 315946 518120 316002 518129
rect 315856 518084 315908 518090
rect 315946 518055 315948 518064
rect 315856 518026 315908 518032
rect 316000 518055 316002 518064
rect 315948 518026 316000 518032
rect 317418 517984 317474 517993
rect 317524 517954 317552 518463
rect 318798 518392 318854 518401
rect 318798 518327 318800 518336
rect 318852 518327 318854 518336
rect 320178 518392 320234 518401
rect 320178 518327 320234 518336
rect 318800 518298 318852 518304
rect 320192 518294 320220 518327
rect 320180 518288 320232 518294
rect 320180 518230 320232 518236
rect 321742 518256 321798 518265
rect 321742 518191 321798 518200
rect 321756 518158 321784 518191
rect 321744 518152 321796 518158
rect 318798 518120 318854 518129
rect 321744 518094 321796 518100
rect 324332 518090 324360 518735
rect 325436 518430 325464 518735
rect 325514 518528 325570 518537
rect 326448 518498 326476 518735
rect 327368 518634 327396 518735
rect 329668 518634 329696 518842
rect 336924 518832 336976 518838
rect 330114 518800 330170 518809
rect 330114 518735 330170 518744
rect 331310 518800 331366 518809
rect 332414 518800 332470 518809
rect 331310 518735 331312 518744
rect 327356 518628 327408 518634
rect 327356 518570 327408 518576
rect 329656 518628 329708 518634
rect 329656 518570 329708 518576
rect 330128 518566 330156 518735
rect 331364 518735 331366 518744
rect 331404 518764 331456 518770
rect 331312 518706 331364 518712
rect 332414 518735 332470 518744
rect 333794 518800 333850 518809
rect 333794 518735 333850 518744
rect 334714 518800 334770 518809
rect 334714 518735 334770 518744
rect 335818 518800 335874 518809
rect 335818 518735 335874 518744
rect 336922 518800 336924 518809
rect 345296 518832 345348 518838
rect 336976 518800 336978 518809
rect 336922 518735 336978 518744
rect 338118 518800 338174 518809
rect 338118 518735 338174 518744
rect 339498 518800 339554 518809
rect 339498 518735 339554 518744
rect 340602 518800 340658 518809
rect 340602 518735 340604 518744
rect 331404 518706 331456 518712
rect 331416 518673 331444 518706
rect 332428 518702 332456 518735
rect 332416 518696 332468 518702
rect 331402 518664 331458 518673
rect 332416 518638 332468 518644
rect 331402 518599 331458 518608
rect 330116 518560 330168 518566
rect 329838 518528 329894 518537
rect 325514 518463 325570 518472
rect 326436 518492 326488 518498
rect 325528 518430 325556 518463
rect 330116 518502 330168 518508
rect 329838 518463 329894 518472
rect 326436 518434 326488 518440
rect 325424 518424 325476 518430
rect 325424 518366 325476 518372
rect 325516 518424 325568 518430
rect 325516 518366 325568 518372
rect 325436 518294 325464 518366
rect 325424 518288 325476 518294
rect 325424 518230 325476 518236
rect 318798 518055 318854 518064
rect 324320 518084 324372 518090
rect 318812 518022 318840 518055
rect 324320 518026 324372 518032
rect 325516 518084 325568 518090
rect 325516 518026 325568 518032
rect 325608 518084 325660 518090
rect 325608 518026 325660 518032
rect 318800 518016 318852 518022
rect 318800 517958 318852 517964
rect 317418 517919 317474 517928
rect 317512 517948 317564 517954
rect 317432 517886 317460 517919
rect 317512 517890 317564 517896
rect 322848 517948 322900 517954
rect 322848 517890 322900 517896
rect 317420 517880 317472 517886
rect 312174 517848 312230 517857
rect 317420 517822 317472 517828
rect 321468 517880 321520 517886
rect 321468 517822 321520 517828
rect 312174 517783 312230 517792
rect 315948 517812 316000 517818
rect 310242 517712 310298 517721
rect 310242 517647 310298 517656
rect 309046 517576 309102 517585
rect 309046 517511 309102 517520
rect 309060 482118 309088 517511
rect 310256 482186 310284 517647
rect 310428 517608 310480 517614
rect 310334 517576 310390 517585
rect 310428 517550 310480 517556
rect 311806 517576 311862 517585
rect 310334 517511 310390 517520
rect 310348 482254 310376 517511
rect 310336 482248 310388 482254
rect 310336 482190 310388 482196
rect 310244 482180 310296 482186
rect 310244 482122 310296 482128
rect 309048 482112 309100 482118
rect 309048 482054 309100 482060
rect 310440 479890 310468 517550
rect 312188 517546 312216 517783
rect 315948 517754 316000 517760
rect 313188 517744 313240 517750
rect 313188 517686 313240 517692
rect 311806 517511 311862 517520
rect 312176 517540 312228 517546
rect 311820 483002 311848 517511
rect 312176 517482 312228 517488
rect 311808 482996 311860 483002
rect 311808 482938 311860 482944
rect 304842 479862 304948 479890
rect 307418 479862 307708 479890
rect 309994 479862 310468 479890
rect 274022 479726 274588 479754
rect 300768 479800 300820 479806
rect 313200 479754 313228 517686
rect 315960 481710 315988 517754
rect 320178 482080 320234 482089
rect 321480 482050 321508 517822
rect 321558 482080 321614 482089
rect 320178 482015 320180 482024
rect 320232 482015 320234 482024
rect 320272 482044 320324 482050
rect 320180 481986 320232 481992
rect 320272 481986 320324 481992
rect 321468 482044 321520 482050
rect 321558 482015 321560 482024
rect 321468 481986 321520 481992
rect 321612 482015 321614 482024
rect 321560 481986 321612 481992
rect 315120 481704 315172 481710
rect 315120 481646 315172 481652
rect 315948 481704 316000 481710
rect 315948 481646 316000 481652
rect 317696 481704 317748 481710
rect 317696 481646 317748 481652
rect 315132 479876 315160 481646
rect 317708 479876 317736 481646
rect 320284 479876 320312 481986
rect 322860 479876 322888 517890
rect 324502 517712 324558 517721
rect 324502 517647 324558 517656
rect 324410 517576 324466 517585
rect 324410 517511 324466 517520
rect 324424 481982 324452 517511
rect 324516 482050 324544 517647
rect 325528 517546 325556 518026
rect 325516 517540 325568 517546
rect 325516 517482 325568 517488
rect 324504 482044 324556 482050
rect 324504 481986 324556 481992
rect 324412 481976 324464 481982
rect 324412 481918 324464 481924
rect 325620 479890 325648 518026
rect 328368 518016 328420 518022
rect 328368 517958 328420 517964
rect 325698 517712 325754 517721
rect 325698 517647 325754 517656
rect 327170 517712 327226 517721
rect 327170 517647 327226 517656
rect 325712 481914 325740 517647
rect 325792 481976 325844 481982
rect 325792 481918 325844 481924
rect 325700 481908 325752 481914
rect 325700 481850 325752 481856
rect 325700 481704 325752 481710
rect 325804 481692 325832 481918
rect 327184 481846 327212 517647
rect 327172 481840 327224 481846
rect 327172 481782 327224 481788
rect 325752 481664 325832 481692
rect 325700 481646 325752 481652
rect 325358 479862 325648 479890
rect 328380 479754 328408 517958
rect 328458 517712 328514 517721
rect 329852 517682 329880 518463
rect 331416 518430 331444 518599
rect 333808 518430 333836 518735
rect 331404 518424 331456 518430
rect 331404 518366 331456 518372
rect 333796 518424 333848 518430
rect 333796 518366 333848 518372
rect 332690 518256 332746 518265
rect 332690 518191 332746 518200
rect 331128 518152 331180 518158
rect 331128 518094 331180 518100
rect 328458 517647 328514 517656
rect 329840 517676 329892 517682
rect 328472 481778 328500 517647
rect 329840 517618 329892 517624
rect 328460 481772 328512 481778
rect 328460 481714 328512 481720
rect 331140 479754 331168 518094
rect 332704 517750 332732 518191
rect 332692 517744 332744 517750
rect 332598 517712 332654 517721
rect 332692 517686 332744 517692
rect 332598 517647 332654 517656
rect 332612 517614 332640 517647
rect 332600 517608 332652 517614
rect 332600 517550 332652 517556
rect 333808 517546 333836 518366
rect 334728 518294 334756 518735
rect 335832 518498 335860 518735
rect 335820 518492 335872 518498
rect 335820 518434 335872 518440
rect 336738 518392 336794 518401
rect 336936 518362 336964 518735
rect 338132 518634 338160 518735
rect 338120 518628 338172 518634
rect 338120 518570 338172 518576
rect 339512 518566 339540 518735
rect 340656 518735 340658 518744
rect 341522 518800 341578 518809
rect 341522 518735 341578 518744
rect 345294 518800 345296 518809
rect 348988 518809 349016 518842
rect 345348 518800 345350 518809
rect 345294 518735 345350 518744
rect 346582 518800 346638 518809
rect 346582 518735 346584 518744
rect 340604 518706 340656 518712
rect 339590 518664 339646 518673
rect 339590 518599 339646 518608
rect 339500 518560 339552 518566
rect 339500 518502 339552 518508
rect 338118 518392 338174 518401
rect 336738 518327 336794 518336
rect 336924 518356 336976 518362
rect 334716 518288 334768 518294
rect 334716 518230 334768 518236
rect 336752 517886 336780 518327
rect 338118 518327 338174 518336
rect 339498 518392 339554 518401
rect 339498 518327 339554 518336
rect 336924 518298 336976 518304
rect 338132 517954 338160 518327
rect 339512 518090 339540 518327
rect 339500 518084 339552 518090
rect 339500 518026 339552 518032
rect 339604 518022 339632 518599
rect 340616 518022 340644 518706
rect 341536 518702 341564 518735
rect 341524 518696 341576 518702
rect 341524 518638 341576 518644
rect 340878 518256 340934 518265
rect 340878 518191 340934 518200
rect 340892 518158 340920 518191
rect 340880 518152 340932 518158
rect 340880 518094 340932 518100
rect 339592 518016 339644 518022
rect 339592 517958 339644 517964
rect 340604 518016 340656 518022
rect 340604 517958 340656 517964
rect 341536 517954 341564 518638
rect 342994 518528 343050 518537
rect 345308 518498 345336 518735
rect 346636 518735 346638 518744
rect 348974 518800 349030 518809
rect 348974 518735 349030 518744
rect 346584 518706 346636 518712
rect 342994 518463 343050 518472
rect 345296 518492 345348 518498
rect 343008 518430 343036 518463
rect 345296 518434 345348 518440
rect 342996 518424 343048 518430
rect 342996 518366 343048 518372
rect 343730 518392 343786 518401
rect 338120 517948 338172 517954
rect 338120 517890 338172 517896
rect 341524 517948 341576 517954
rect 341524 517890 341576 517896
rect 343008 517886 343036 518366
rect 346596 518362 346624 518706
rect 347686 518664 347742 518673
rect 347686 518599 347688 518608
rect 347740 518599 347742 518608
rect 347688 518570 347740 518576
rect 348988 518566 349016 518735
rect 348976 518560 349028 518566
rect 347778 518528 347834 518537
rect 348976 518502 349028 518508
rect 347778 518463 347834 518472
rect 343730 518327 343786 518336
rect 346584 518356 346636 518362
rect 343744 518294 343772 518327
rect 346584 518298 346636 518304
rect 343732 518288 343784 518294
rect 343732 518230 343784 518236
rect 344376 518288 344428 518294
rect 344376 518230 344428 518236
rect 336740 517880 336792 517886
rect 333978 517848 334034 517857
rect 342996 517880 343048 517886
rect 336740 517822 336792 517828
rect 342258 517848 342314 517857
rect 333978 517783 333980 517792
rect 334032 517783 334034 517792
rect 342996 517822 343048 517828
rect 344388 517818 344416 518230
rect 342258 517783 342314 517792
rect 344376 517812 344428 517818
rect 333980 517754 334032 517760
rect 342272 517750 342300 517783
rect 344376 517754 344428 517760
rect 333888 517744 333940 517750
rect 342260 517744 342312 517750
rect 333888 517686 333940 517692
rect 335358 517712 335414 517721
rect 333796 517540 333848 517546
rect 333796 517482 333848 517488
rect 333900 482050 333928 517686
rect 344284 517744 344336 517750
rect 342260 517686 342312 517692
rect 343638 517712 343694 517721
rect 335358 517647 335414 517656
rect 337384 517676 337436 517682
rect 333060 482044 333112 482050
rect 333060 481986 333112 481992
rect 333888 482044 333940 482050
rect 333888 481986 333940 481992
rect 333072 479876 333100 481986
rect 335372 481778 335400 517647
rect 344284 517686 344336 517692
rect 345202 517712 345258 517721
rect 343638 517647 343640 517656
rect 337384 517618 337436 517624
rect 343692 517647 343694 517656
rect 343640 517618 343692 517624
rect 337396 481778 337424 517618
rect 340788 517608 340840 517614
rect 340788 517550 340840 517556
rect 339408 517540 339460 517546
rect 339408 517482 339460 517488
rect 339420 482050 339448 517482
rect 338212 482044 338264 482050
rect 338212 481986 338264 481992
rect 339408 482044 339460 482050
rect 339408 481986 339460 481992
rect 335360 481772 335412 481778
rect 335360 481714 335412 481720
rect 335636 481772 335688 481778
rect 335636 481714 335688 481720
rect 337384 481772 337436 481778
rect 337384 481714 337436 481720
rect 335648 479876 335676 481714
rect 338224 479876 338252 481986
rect 340800 479876 340828 517550
rect 344296 482050 344324 517686
rect 345202 517647 345258 517656
rect 346398 517712 346454 517721
rect 346398 517647 346454 517656
rect 345216 517546 345244 517647
rect 346412 517614 346440 517647
rect 346400 517608 346452 517614
rect 346400 517550 346452 517556
rect 347792 517546 347820 518463
rect 369768 518424 369820 518430
rect 369768 518366 369820 518372
rect 357348 518356 357400 518362
rect 357348 518298 357400 518304
rect 354588 518288 354640 518294
rect 354588 518230 354640 518236
rect 351828 518152 351880 518158
rect 351828 518094 351880 518100
rect 349068 518084 349120 518090
rect 349068 518026 349120 518032
rect 347870 517848 347926 517857
rect 347870 517783 347926 517792
rect 347884 517750 347912 517783
rect 347872 517744 347924 517750
rect 347872 517686 347924 517692
rect 345204 517540 345256 517546
rect 345204 517482 345256 517488
rect 346308 517540 346360 517546
rect 346308 517482 346360 517488
rect 347780 517540 347832 517546
rect 347780 517482 347832 517488
rect 343364 482044 343416 482050
rect 343364 481986 343416 481992
rect 344284 482044 344336 482050
rect 344284 481986 344336 481992
rect 343376 479876 343404 481986
rect 346320 479890 346348 517482
rect 345966 479862 346348 479890
rect 349080 479754 349108 518026
rect 351840 482050 351868 518094
rect 354600 482050 354628 518230
rect 351092 482044 351144 482050
rect 351092 481986 351144 481992
rect 351828 482044 351880 482050
rect 351828 481986 351880 481992
rect 353668 482044 353720 482050
rect 353668 481986 353720 481992
rect 354588 482044 354640 482050
rect 354588 481986 354640 481992
rect 351104 479876 351132 481986
rect 353680 479876 353708 481986
rect 357360 481914 357388 518298
rect 366456 482996 366508 483002
rect 366456 482938 366508 482944
rect 363880 482248 363932 482254
rect 363880 482190 363932 482196
rect 361304 482180 361356 482186
rect 361304 482122 361356 482128
rect 358728 482112 358780 482118
rect 358728 482054 358780 482060
rect 356152 481908 356204 481914
rect 356152 481850 356204 481856
rect 357348 481908 357400 481914
rect 357348 481850 357400 481856
rect 356164 479876 356192 481850
rect 358740 479876 358768 482054
rect 361316 479876 361344 482122
rect 363892 479876 363920 482190
rect 366468 479876 366496 482938
rect 369780 479754 369808 518366
rect 371608 482996 371660 483002
rect 371608 482938 371660 482944
rect 371620 479876 371648 482938
rect 378060 482322 378088 600306
rect 376760 482316 376812 482322
rect 376760 482258 376812 482264
rect 378048 482316 378100 482322
rect 378048 482258 378100 482264
rect 374184 482248 374236 482254
rect 374184 482190 374236 482196
rect 374196 479876 374224 482190
rect 376772 479876 376800 482258
rect 379440 479890 379468 601666
rect 379624 549409 379652 612750
rect 379980 610428 380032 610434
rect 379980 610370 380032 610376
rect 379992 609657 380020 610370
rect 379702 609648 379758 609657
rect 379702 609583 379758 609592
rect 379978 609648 380034 609657
rect 379978 609583 380034 609592
rect 379610 549400 379666 549409
rect 379610 549335 379666 549344
rect 379520 538280 379572 538286
rect 379520 538222 379572 538228
rect 379532 536110 379560 538222
rect 379520 536104 379572 536110
rect 379520 536046 379572 536052
rect 379612 518968 379664 518974
rect 379612 518910 379664 518916
rect 379624 514078 379652 518910
rect 379612 514072 379664 514078
rect 379612 514014 379664 514020
rect 379612 499588 379664 499594
rect 379612 499530 379664 499536
rect 379624 494766 379652 499530
rect 379612 494760 379664 494766
rect 379612 494702 379664 494708
rect 379716 482225 379744 609583
rect 387708 605872 387760 605878
rect 387708 605814 387760 605820
rect 384948 604512 385000 604518
rect 384948 604454 385000 604460
rect 382188 603152 382240 603158
rect 382188 603094 382240 603100
rect 379794 540968 379850 540977
rect 379794 540903 379850 540912
rect 379808 538286 379836 540903
rect 379796 538280 379848 538286
rect 379796 538222 379848 538228
rect 379796 536104 379848 536110
rect 379796 536046 379848 536052
rect 379808 518974 379836 536046
rect 379796 518968 379848 518974
rect 379796 518910 379848 518916
rect 379796 514072 379848 514078
rect 379796 514014 379848 514020
rect 379808 499594 379836 514014
rect 379796 499588 379848 499594
rect 379796 499530 379848 499536
rect 379796 494760 379848 494766
rect 379796 494702 379848 494708
rect 379702 482216 379758 482225
rect 379702 482151 379758 482160
rect 379808 482118 379836 494702
rect 379796 482112 379848 482118
rect 379796 482054 379848 482060
rect 382200 479890 382228 603094
rect 384960 479890 384988 604454
rect 387720 482934 387748 605814
rect 398760 487830 398788 699926
rect 429856 699718 429884 703520
rect 462332 699718 462360 703520
rect 478524 700942 478552 703520
rect 478512 700936 478564 700942
rect 478512 700878 478564 700884
rect 494808 699854 494836 703520
rect 494796 699848 494848 699854
rect 494796 699790 494848 699796
rect 495348 699848 495400 699854
rect 495348 699790 495400 699796
rect 429844 699712 429896 699718
rect 429844 699654 429896 699660
rect 430488 699712 430540 699718
rect 430488 699654 430540 699660
rect 462320 699712 462372 699718
rect 462320 699654 462372 699660
rect 463608 699712 463660 699718
rect 463608 699654 463660 699660
rect 430500 610706 430528 699654
rect 463620 610774 463648 699654
rect 488540 613420 488592 613426
rect 488540 613362 488592 613368
rect 493968 613420 494020 613426
rect 493968 613362 494020 613368
rect 488552 612814 488580 613362
rect 493980 612814 494008 613362
rect 488540 612808 488592 612814
rect 488538 612776 488540 612785
rect 493968 612808 494020 612814
rect 488592 612776 488594 612785
rect 488538 612711 488594 612720
rect 493966 612776 493968 612785
rect 494020 612776 494022 612785
rect 493966 612711 494022 612720
rect 495360 610842 495388 699790
rect 527192 699718 527220 703520
rect 539600 700936 539652 700942
rect 539600 700878 539652 700884
rect 539140 700732 539192 700738
rect 539140 700674 539192 700680
rect 527180 699712 527232 699718
rect 527180 699654 527232 699660
rect 528468 699712 528520 699718
rect 528468 699654 528520 699660
rect 499580 612808 499632 612814
rect 499580 612750 499632 612756
rect 495348 610836 495400 610842
rect 495348 610778 495400 610784
rect 463608 610768 463660 610774
rect 463608 610710 463660 610716
rect 430488 610700 430540 610706
rect 430488 610642 430540 610648
rect 496452 610428 496504 610434
rect 496452 610370 496504 610376
rect 496464 609929 496492 610370
rect 496450 609920 496506 609929
rect 496450 609855 496506 609864
rect 416778 606112 416834 606121
rect 416778 606047 416834 606056
rect 416792 605878 416820 606047
rect 416780 605872 416832 605878
rect 416780 605814 416832 605820
rect 416778 604888 416834 604897
rect 416778 604823 416834 604832
rect 416792 604518 416820 604823
rect 416780 604512 416832 604518
rect 416780 604454 416832 604460
rect 416778 603256 416834 603265
rect 416778 603191 416834 603200
rect 416792 603158 416820 603191
rect 416780 603152 416832 603158
rect 416780 603094 416832 603100
rect 416778 602032 416834 602041
rect 416778 601967 416834 601976
rect 416792 601730 416820 601967
rect 416780 601724 416832 601730
rect 416780 601666 416832 601672
rect 416778 600536 416834 600545
rect 416778 600471 416834 600480
rect 416792 600370 416820 600471
rect 416780 600364 416832 600370
rect 416780 600306 416832 600312
rect 417422 599312 417478 599321
rect 417422 599247 417478 599256
rect 416962 539744 417018 539753
rect 416962 539679 417018 539688
rect 416976 539646 417004 539679
rect 413928 539640 413980 539646
rect 413928 539582 413980 539588
rect 416964 539640 417016 539646
rect 416964 539582 417016 539588
rect 410524 538280 410576 538286
rect 410524 538222 410576 538228
rect 410536 521626 410564 538222
rect 409880 521620 409932 521626
rect 409880 521562 409932 521568
rect 410524 521620 410576 521626
rect 410524 521562 410576 521568
rect 409892 520946 409920 521562
rect 409880 520940 409932 520946
rect 409880 520882 409932 520888
rect 398748 487824 398800 487830
rect 398748 487766 398800 487772
rect 386972 482928 387024 482934
rect 386972 482870 387024 482876
rect 387708 482928 387760 482934
rect 387708 482870 387760 482876
rect 386512 482860 386564 482866
rect 386512 482802 386564 482808
rect 386524 482322 386552 482802
rect 386512 482316 386564 482322
rect 386512 482258 386564 482264
rect 379362 479862 379468 479890
rect 381938 479862 382228 479890
rect 384514 479862 384988 479890
rect 386984 479876 387012 482870
rect 389548 482860 389600 482866
rect 389548 482802 389600 482808
rect 389560 479876 389588 482802
rect 394700 482792 394752 482798
rect 394700 482734 394752 482740
rect 392124 482316 392176 482322
rect 392124 482258 392176 482264
rect 392136 479876 392164 482258
rect 394712 479876 394740 482734
rect 397276 482724 397328 482730
rect 397276 482666 397328 482672
rect 397288 479876 397316 482666
rect 399852 482656 399904 482662
rect 399852 482598 399904 482604
rect 399864 479876 399892 482598
rect 402428 482588 402480 482594
rect 402428 482530 402480 482536
rect 402440 479876 402468 482530
rect 405004 482520 405056 482526
rect 405004 482462 405056 482468
rect 405016 479876 405044 482462
rect 407580 482452 407632 482458
rect 407580 482394 407632 482400
rect 407592 479876 407620 482394
rect 409892 479890 409920 520882
rect 413940 482594 413968 539582
rect 416778 538384 416834 538393
rect 416778 538319 416834 538328
rect 416792 538286 416820 538319
rect 416780 538280 416832 538286
rect 416780 538222 416832 538228
rect 412732 482588 412784 482594
rect 412732 482530 412784 482536
rect 413928 482588 413980 482594
rect 413928 482530 413980 482536
rect 409892 479862 410182 479890
rect 412744 479876 412772 482530
rect 415308 482384 415360 482390
rect 415308 482326 415360 482332
rect 415320 479876 415348 482326
rect 417436 482254 417464 599247
rect 417514 597680 417570 597689
rect 417514 597615 417570 597624
rect 417528 483002 417556 597615
rect 499592 549545 499620 612750
rect 499578 549536 499634 549545
rect 499578 549471 499634 549480
rect 499578 542056 499634 542065
rect 499578 541991 499634 542000
rect 499592 540977 499620 541991
rect 499578 540968 499634 540977
rect 499578 540903 499634 540912
rect 425334 519752 425390 519761
rect 425334 519687 425390 519696
rect 434166 519752 434222 519761
rect 434166 519687 434222 519696
rect 423678 518256 423734 518265
rect 423678 518191 423680 518200
rect 423732 518191 423734 518200
rect 423680 518162 423732 518168
rect 425348 518090 425376 519687
rect 429290 518664 429346 518673
rect 429290 518599 429346 518608
rect 426438 518528 426494 518537
rect 426438 518463 426494 518472
rect 426452 518430 426480 518463
rect 426440 518424 426492 518430
rect 426440 518366 426492 518372
rect 429304 518294 429332 518599
rect 430578 518392 430634 518401
rect 430578 518327 430580 518336
rect 430632 518327 430634 518336
rect 430580 518298 430632 518304
rect 429292 518288 429344 518294
rect 429198 518256 429254 518265
rect 429292 518230 429344 518236
rect 429198 518191 429254 518200
rect 429212 518158 429240 518191
rect 429200 518152 429252 518158
rect 429200 518094 429252 518100
rect 425336 518084 425388 518090
rect 425336 518026 425388 518032
rect 432604 518084 432656 518090
rect 432604 518026 432656 518032
rect 432616 517857 432644 518026
rect 432602 517848 432658 517857
rect 432602 517783 432658 517792
rect 417516 482996 417568 483002
rect 417516 482938 417568 482944
rect 430672 482792 430724 482798
rect 430672 482734 430724 482740
rect 428096 482724 428148 482730
rect 428096 482666 428148 482672
rect 425520 482656 425572 482662
rect 425520 482598 425572 482604
rect 422944 482588 422996 482594
rect 422944 482530 422996 482536
rect 420368 482384 420420 482390
rect 420368 482326 420420 482332
rect 417792 482316 417844 482322
rect 417792 482258 417844 482264
rect 417424 482248 417476 482254
rect 417424 482190 417476 482196
rect 417804 479876 417832 482258
rect 420380 479876 420408 482326
rect 422956 479876 422984 482530
rect 425532 479876 425560 482598
rect 428108 479876 428136 482666
rect 430684 479876 430712 482734
rect 432616 482322 432644 517783
rect 433246 517712 433302 517721
rect 433246 517647 433302 517656
rect 433156 482996 433208 483002
rect 433156 482938 433208 482944
rect 432604 482316 432656 482322
rect 432604 482258 432656 482264
rect 433168 479890 433196 482938
rect 433260 482526 433288 517647
rect 434180 517546 434208 519687
rect 455420 518900 455472 518906
rect 455420 518842 455472 518848
rect 448520 518832 448572 518838
rect 443182 518800 443238 518809
rect 448520 518774 448572 518780
rect 448704 518832 448756 518838
rect 448704 518774 448756 518780
rect 451278 518800 451334 518809
rect 443182 518735 443238 518744
rect 443196 518702 443224 518735
rect 443184 518696 443236 518702
rect 442538 518664 442594 518673
rect 443184 518638 443236 518644
rect 444286 518664 444342 518673
rect 442538 518599 442594 518608
rect 442552 518566 442580 518599
rect 442540 518560 442592 518566
rect 442540 518502 442592 518508
rect 435362 518392 435418 518401
rect 435362 518327 435418 518336
rect 435914 518392 435970 518401
rect 435914 518327 435916 518336
rect 434626 517712 434682 517721
rect 434626 517647 434682 517656
rect 434168 517540 434220 517546
rect 434168 517482 434220 517488
rect 434180 512038 434208 517482
rect 434076 512032 434128 512038
rect 434076 511974 434128 511980
rect 434168 512032 434220 512038
rect 434168 511974 434220 511980
rect 434088 495553 434116 511974
rect 434074 495544 434130 495553
rect 434074 495479 434130 495488
rect 433890 492688 433946 492697
rect 433616 492652 433668 492658
rect 433890 492623 433892 492632
rect 433616 492594 433668 492600
rect 433944 492623 433946 492632
rect 433892 492594 433944 492600
rect 433628 483041 433656 492594
rect 433614 483032 433670 483041
rect 433614 482967 433670 482976
rect 433798 483032 433854 483041
rect 433798 482967 433854 482976
rect 433248 482520 433300 482526
rect 433248 482462 433300 482468
rect 433812 482390 433840 482967
rect 434640 482458 434668 517647
rect 435376 482594 435404 518327
rect 435968 518327 435970 518336
rect 435916 518298 435968 518304
rect 436926 518256 436982 518265
rect 436926 518191 436928 518200
rect 436980 518191 436982 518200
rect 440882 518256 440938 518265
rect 440882 518191 440938 518200
rect 436928 518162 436980 518168
rect 436006 517712 436062 517721
rect 436006 517647 436062 517656
rect 435364 482588 435416 482594
rect 435364 482530 435416 482536
rect 434628 482452 434680 482458
rect 434628 482394 434680 482400
rect 436020 482390 436048 517647
rect 436744 517608 436796 517614
rect 436744 517550 436796 517556
rect 436756 482730 436784 517550
rect 436744 482724 436796 482730
rect 436744 482666 436796 482672
rect 436940 482662 436968 518162
rect 440896 518158 440924 518191
rect 440884 518152 440936 518158
rect 440884 518094 440936 518100
rect 437480 518016 437532 518022
rect 437480 517958 437532 517964
rect 439504 518016 439556 518022
rect 439504 517958 439556 517964
rect 437294 517848 437350 517857
rect 437294 517783 437350 517792
rect 437308 517614 437336 517783
rect 437386 517712 437442 517721
rect 437386 517647 437442 517656
rect 437296 517608 437348 517614
rect 437296 517550 437348 517556
rect 436928 482656 436980 482662
rect 436928 482598 436980 482604
rect 433800 482384 433852 482390
rect 433800 482326 433852 482332
rect 436008 482384 436060 482390
rect 436008 482326 436060 482332
rect 437400 482322 437428 517647
rect 437388 482316 437440 482322
rect 437388 482258 437440 482264
rect 435824 482180 435876 482186
rect 435824 482122 435876 482128
rect 433168 479862 433274 479890
rect 435836 479876 435864 482122
rect 437492 480026 437520 517958
rect 438674 517712 438730 517721
rect 438124 517676 438176 517682
rect 438674 517647 438730 517656
rect 438124 517618 438176 517624
rect 438136 517585 438164 517618
rect 438122 517576 438178 517585
rect 438122 517511 438178 517520
rect 438136 482798 438164 517511
rect 438124 482792 438176 482798
rect 438124 482734 438176 482740
rect 438688 481710 438716 517647
rect 439516 517585 439544 517958
rect 440240 517948 440292 517954
rect 440240 517890 440292 517896
rect 438766 517576 438822 517585
rect 438766 517511 438822 517520
rect 439502 517576 439558 517585
rect 439502 517511 439558 517520
rect 440146 517576 440202 517585
rect 440146 517511 440202 517520
rect 438780 481778 438808 517511
rect 439516 483002 439544 517511
rect 439504 482996 439556 483002
rect 439504 482938 439556 482944
rect 440160 481846 440188 517511
rect 440148 481840 440200 481846
rect 440148 481782 440200 481788
rect 438768 481772 438820 481778
rect 438768 481714 438820 481720
rect 438676 481704 438728 481710
rect 438676 481646 438728 481652
rect 437492 479998 437980 480026
rect 300768 479742 300820 479748
rect 312570 479726 313228 479754
rect 327934 479726 328408 479754
rect 330510 479726 331168 479754
rect 348542 479726 349108 479754
rect 369058 479726 369808 479754
rect 437952 479754 437980 479998
rect 440252 479890 440280 517890
rect 440896 482186 440924 518094
rect 442552 518090 442580 518502
rect 442540 518084 442592 518090
rect 442540 518026 442592 518032
rect 443000 517880 443052 517886
rect 443000 517822 443052 517828
rect 441526 517576 441582 517585
rect 441526 517511 441582 517520
rect 442906 517576 442962 517585
rect 442906 517511 442962 517520
rect 440884 482180 440936 482186
rect 440884 482122 440936 482128
rect 441540 481914 441568 517511
rect 442920 481982 442948 517511
rect 442908 481976 442960 481982
rect 442908 481918 442960 481924
rect 441528 481908 441580 481914
rect 441528 481850 441580 481856
rect 440252 479862 440556 479890
rect 440528 479754 440556 479862
rect 443012 479754 443040 517822
rect 443196 517546 443224 518638
rect 444286 518599 444342 518608
rect 445390 518664 445446 518673
rect 445390 518599 445446 518608
rect 446402 518664 446458 518673
rect 446402 518599 446458 518608
rect 444102 518528 444158 518537
rect 444102 518463 444158 518472
rect 444116 517954 444144 518463
rect 444300 518430 444328 518599
rect 444288 518424 444340 518430
rect 444288 518366 444340 518372
rect 445404 518362 445432 518599
rect 445482 518528 445538 518537
rect 445482 518463 445538 518472
rect 445392 518356 445444 518362
rect 445392 518298 445444 518304
rect 444104 517948 444156 517954
rect 444104 517890 444156 517896
rect 445496 517546 445524 518463
rect 445574 518392 445630 518401
rect 445574 518327 445630 518336
rect 445588 517886 445616 518327
rect 446416 518294 446444 518599
rect 447138 518528 447194 518537
rect 447138 518463 447194 518472
rect 447966 518528 448022 518537
rect 447966 518463 447968 518472
rect 447046 518392 447102 518401
rect 447046 518327 447102 518336
rect 446404 518288 446456 518294
rect 446404 518230 446456 518236
rect 445576 517880 445628 517886
rect 445576 517822 445628 517828
rect 445760 517812 445812 517818
rect 445760 517754 445812 517760
rect 443184 517540 443236 517546
rect 443184 517482 443236 517488
rect 445484 517540 445536 517546
rect 445484 517482 445536 517488
rect 445772 479890 445800 517754
rect 446416 517614 446444 518230
rect 447060 517750 447088 518327
rect 447048 517744 447100 517750
rect 447048 517686 447100 517692
rect 447152 517682 447180 518463
rect 448020 518463 448022 518472
rect 447968 518434 448020 518440
rect 448334 518256 448390 518265
rect 448334 518191 448390 518200
rect 448348 517682 448376 518191
rect 447140 517676 447192 517682
rect 447140 517618 447192 517624
rect 448336 517676 448388 517682
rect 448336 517618 448388 517624
rect 446404 517608 446456 517614
rect 446404 517550 446456 517556
rect 448532 479890 448560 518774
rect 448716 518537 448744 518774
rect 449900 518764 449952 518770
rect 451278 518735 451280 518744
rect 449900 518706 449952 518712
rect 451332 518735 451334 518744
rect 452566 518800 452622 518809
rect 452566 518735 452622 518744
rect 451280 518706 451332 518712
rect 448702 518528 448758 518537
rect 448702 518463 448758 518472
rect 448716 518022 448744 518463
rect 448704 518016 448756 518022
rect 448704 517958 448756 517964
rect 449806 517576 449862 517585
rect 449806 517511 449862 517520
rect 449820 482050 449848 517511
rect 449808 482044 449860 482050
rect 449808 481986 449860 481992
rect 449912 480026 449940 518706
rect 451292 518566 451320 518706
rect 452580 518702 452608 518735
rect 452568 518696 452620 518702
rect 452568 518638 452620 518644
rect 452660 518628 452712 518634
rect 452660 518570 452712 518576
rect 451280 518560 451332 518566
rect 451280 518502 451332 518508
rect 450174 518392 450230 518401
rect 450174 518327 450230 518336
rect 450188 518226 450216 518327
rect 450176 518220 450228 518226
rect 450176 518162 450228 518168
rect 451186 517576 451242 517585
rect 451186 517511 451242 517520
rect 452566 517576 452622 517585
rect 452566 517511 452622 517520
rect 451200 482118 451228 517511
rect 452580 482186 452608 517511
rect 452568 482180 452620 482186
rect 452568 482122 452620 482128
rect 451188 482112 451240 482118
rect 451188 482054 451240 482060
rect 452672 480026 452700 518570
rect 453762 518528 453818 518537
rect 453762 518463 453818 518472
rect 455326 518528 455382 518537
rect 455326 518463 455382 518472
rect 453776 518430 453804 518463
rect 453764 518424 453816 518430
rect 453764 518366 453816 518372
rect 455340 518362 455368 518463
rect 455328 518356 455380 518362
rect 455328 518298 455380 518304
rect 453854 517712 453910 517721
rect 453854 517647 453910 517656
rect 453868 482254 453896 517647
rect 453946 517576 454002 517585
rect 453946 517511 454002 517520
rect 455326 517576 455382 517585
rect 455326 517511 455382 517520
rect 453960 482934 453988 517511
rect 455340 483002 455368 517511
rect 455328 482996 455380 483002
rect 455328 482938 455380 482944
rect 453948 482928 454000 482934
rect 453948 482870 454000 482876
rect 453856 482248 453908 482254
rect 453856 482190 453908 482196
rect 455432 480026 455460 518842
rect 458364 518832 458416 518838
rect 458362 518800 458364 518809
rect 458416 518800 458418 518809
rect 458362 518735 458418 518744
rect 459558 518800 459614 518809
rect 459558 518735 459560 518744
rect 457088 518702 457116 518733
rect 457076 518696 457128 518702
rect 457074 518664 457076 518673
rect 457128 518664 457130 518673
rect 457074 518599 457130 518608
rect 456062 518528 456118 518537
rect 457088 518498 457116 518599
rect 458376 518498 458404 518735
rect 459612 518735 459614 518744
rect 466458 518800 466514 518809
rect 466458 518735 466514 518744
rect 459560 518706 459612 518712
rect 466472 518702 466500 518735
rect 466460 518696 466512 518702
rect 461030 518664 461086 518673
rect 466460 518638 466512 518644
rect 461030 518599 461086 518608
rect 461044 518566 461072 518599
rect 461032 518560 461084 518566
rect 461032 518502 461084 518508
rect 462318 518528 462374 518537
rect 456062 518463 456118 518472
rect 457076 518492 457128 518498
rect 456076 518294 456104 518463
rect 457076 518434 457128 518440
rect 458364 518492 458416 518498
rect 462318 518463 462374 518472
rect 463698 518528 463754 518537
rect 463698 518463 463754 518472
rect 466458 518528 466514 518537
rect 466458 518463 466460 518472
rect 458364 518434 458416 518440
rect 462332 518430 462360 518463
rect 462320 518424 462372 518430
rect 459558 518392 459614 518401
rect 462320 518366 462372 518372
rect 463712 518362 463740 518463
rect 466512 518463 466514 518472
rect 466460 518434 466512 518440
rect 465078 518392 465134 518401
rect 459558 518327 459614 518336
rect 463700 518356 463752 518362
rect 456064 518288 456116 518294
rect 456064 518230 456116 518236
rect 459572 518226 459600 518327
rect 465078 518327 465134 518336
rect 463700 518298 463752 518304
rect 465092 518294 465120 518327
rect 465080 518288 465132 518294
rect 465080 518230 465132 518236
rect 467838 518256 467894 518265
rect 459560 518220 459612 518226
rect 467838 518191 467840 518200
rect 459560 518162 459612 518168
rect 467892 518191 467894 518200
rect 467840 518162 467892 518168
rect 469864 517948 469916 517954
rect 469864 517890 469916 517896
rect 460846 517712 460902 517721
rect 460846 517647 460902 517656
rect 469034 517712 469090 517721
rect 469034 517647 469090 517656
rect 456706 517576 456762 517585
rect 456706 517511 456762 517520
rect 458086 517576 458142 517585
rect 458086 517511 458142 517520
rect 459466 517576 459522 517585
rect 459466 517511 459522 517520
rect 460754 517576 460810 517585
rect 460754 517511 460810 517520
rect 456720 482866 456748 517511
rect 456708 482860 456760 482866
rect 456708 482802 456760 482808
rect 458100 482798 458128 517511
rect 458088 482792 458140 482798
rect 458088 482734 458140 482740
rect 459480 482730 459508 517511
rect 459468 482724 459520 482730
rect 459468 482666 459520 482672
rect 460768 482594 460796 517511
rect 460860 482662 460888 517647
rect 462226 517576 462282 517585
rect 462226 517511 462282 517520
rect 463606 517576 463662 517585
rect 463606 517511 463662 517520
rect 464986 517576 465042 517585
rect 464986 517511 465042 517520
rect 466366 517576 466422 517585
rect 466366 517511 466422 517520
rect 467746 517576 467802 517585
rect 467746 517511 467802 517520
rect 460848 482656 460900 482662
rect 460848 482598 460900 482604
rect 460756 482588 460808 482594
rect 460756 482530 460808 482536
rect 458916 482520 458968 482526
rect 458916 482462 458968 482468
rect 449912 479998 450676 480026
rect 452672 479998 453252 480026
rect 455432 479998 455828 480026
rect 445772 479862 446154 479890
rect 448532 479862 448638 479890
rect 450648 479754 450676 479998
rect 453224 479754 453252 479998
rect 455800 479754 455828 479998
rect 458928 479876 458956 482462
rect 462240 482458 462268 517511
rect 463620 482526 463648 517511
rect 463608 482520 463660 482526
rect 463608 482462 463660 482468
rect 461492 482452 461544 482458
rect 461492 482394 461544 482400
rect 462228 482452 462280 482458
rect 462228 482394 462280 482400
rect 461504 479876 461532 482394
rect 465000 482390 465028 517511
rect 466380 482497 466408 517511
rect 466366 482488 466422 482497
rect 466366 482423 466422 482432
rect 464068 482384 464120 482390
rect 464068 482326 464120 482332
rect 464988 482384 465040 482390
rect 464988 482326 465040 482332
rect 464080 479876 464108 482326
rect 467760 482322 467788 517511
rect 469048 482361 469076 517647
rect 469126 517576 469182 517585
rect 469126 517511 469182 517520
rect 469034 482352 469090 482361
rect 466644 482316 466696 482322
rect 466644 482258 466696 482264
rect 467748 482316 467800 482322
rect 469034 482287 469090 482296
rect 467748 482258 467800 482264
rect 466656 479876 466684 482258
rect 469140 482225 469168 517511
rect 469126 482216 469182 482225
rect 469126 482151 469182 482160
rect 469876 481710 469904 517890
rect 476764 517880 476816 517886
rect 476764 517822 476816 517828
rect 474004 517744 474056 517750
rect 474004 517686 474056 517692
rect 471244 517676 471296 517682
rect 471244 517618 471296 517624
rect 471256 481817 471284 517618
rect 471242 481808 471298 481817
rect 474016 481778 474044 517686
rect 476776 481846 476804 517822
rect 479524 517540 479576 517546
rect 479524 517482 479576 517488
rect 479536 481982 479564 517482
rect 507768 482996 507820 483002
rect 507768 482938 507820 482944
rect 505192 482928 505244 482934
rect 505192 482870 505244 482876
rect 502616 482248 502668 482254
rect 502616 482190 502668 482196
rect 500040 482180 500092 482186
rect 500040 482122 500092 482128
rect 497464 482112 497516 482118
rect 497464 482054 497516 482060
rect 494888 482044 494940 482050
rect 494888 481986 494940 481992
rect 479432 481976 479484 481982
rect 479432 481918 479484 481924
rect 479524 481976 479576 481982
rect 479524 481918 479576 481924
rect 484584 481976 484636 481982
rect 484584 481918 484636 481924
rect 476948 481908 477000 481914
rect 476948 481850 477000 481856
rect 474372 481840 474424 481846
rect 474372 481782 474424 481788
rect 476764 481840 476816 481846
rect 476764 481782 476816 481788
rect 471242 481743 471298 481752
rect 471796 481772 471848 481778
rect 471796 481714 471848 481720
rect 474004 481772 474056 481778
rect 474004 481714 474056 481720
rect 469220 481704 469272 481710
rect 469220 481646 469272 481652
rect 469864 481704 469916 481710
rect 469864 481646 469916 481652
rect 469232 479876 469260 481646
rect 471808 479876 471836 481714
rect 474384 479876 474412 481782
rect 476960 479876 476988 481850
rect 477222 481808 477278 481817
rect 477222 481743 477224 481752
rect 477276 481743 477278 481752
rect 477224 481714 477276 481720
rect 477132 481704 477184 481710
rect 477316 481704 477368 481710
rect 477184 481652 477316 481658
rect 477132 481646 477368 481652
rect 477144 481630 477356 481646
rect 479444 479876 479472 481918
rect 482008 481704 482060 481710
rect 482008 481646 482060 481652
rect 482020 479876 482048 481646
rect 484596 479876 484624 481918
rect 487160 481908 487212 481914
rect 487160 481850 487212 481856
rect 487172 479876 487200 481850
rect 489736 481840 489788 481846
rect 489736 481782 489788 481788
rect 489748 479876 489776 481782
rect 492312 481772 492364 481778
rect 492312 481714 492364 481720
rect 492324 479876 492352 481714
rect 494900 479876 494928 481986
rect 497476 479876 497504 482054
rect 500052 479876 500080 482122
rect 502628 479876 502656 482190
rect 505204 479876 505232 482870
rect 507780 479876 507808 482938
rect 510252 482860 510304 482866
rect 510252 482802 510304 482808
rect 510264 479876 510292 482802
rect 512828 482792 512880 482798
rect 512828 482734 512880 482740
rect 512840 479876 512868 482734
rect 515404 482724 515456 482730
rect 515404 482666 515456 482672
rect 515416 479876 515444 482666
rect 517980 482656 518032 482662
rect 517980 482598 518032 482604
rect 517992 479876 518020 482598
rect 520556 482588 520608 482594
rect 520556 482530 520608 482536
rect 520568 479876 520596 482530
rect 525708 482520 525760 482526
rect 525708 482462 525760 482468
rect 523132 482452 523184 482458
rect 523132 482394 523184 482400
rect 523144 479876 523172 482394
rect 525720 479876 525748 482462
rect 528284 482384 528336 482390
rect 528284 482326 528336 482332
rect 528296 479876 528324 482326
rect 528480 479874 528508 699654
rect 530858 482488 530914 482497
rect 530858 482423 530914 482432
rect 530872 479876 530900 482423
rect 536010 482352 536066 482361
rect 533436 482316 533488 482322
rect 536010 482287 536066 482296
rect 533436 482258 533488 482264
rect 533448 479876 533476 482258
rect 536024 479876 536052 482287
rect 538586 482216 538642 482225
rect 538586 482151 538642 482160
rect 538600 479876 538628 482151
rect 528468 479868 528520 479874
rect 528468 479810 528520 479816
rect 437952 479726 438426 479754
rect 440528 479726 441002 479754
rect 443012 479726 443578 479754
rect 450648 479726 451214 479754
rect 453224 479726 453790 479754
rect 455800 479726 456366 479754
rect 539152 357354 539180 700674
rect 539232 700664 539284 700670
rect 539232 700606 539284 700612
rect 539244 365702 539272 700606
rect 539324 610768 539376 610774
rect 539324 610710 539376 610716
rect 539232 365696 539284 365702
rect 539232 365638 539284 365644
rect 539336 357474 539364 610710
rect 539508 509312 539560 509318
rect 539508 509254 539560 509260
rect 539416 487824 539468 487830
rect 539416 487766 539468 487772
rect 539324 357468 539376 357474
rect 539324 357410 539376 357416
rect 539322 357368 539378 357377
rect 539152 357326 539322 357354
rect 539322 357303 539378 357312
rect 539324 357264 539376 357270
rect 539324 357206 539376 357212
rect 539336 344321 539364 357206
rect 539428 350713 539456 487766
rect 539520 412185 539548 509254
rect 539506 412176 539562 412185
rect 539506 412111 539562 412120
rect 539506 406464 539562 406473
rect 539506 406399 539562 406408
rect 539520 405793 539548 406399
rect 539506 405784 539562 405793
rect 539506 405719 539562 405728
rect 539506 402248 539562 402257
rect 539506 402183 539562 402192
rect 539520 391377 539548 402183
rect 539506 391368 539562 391377
rect 539506 391303 539562 391312
rect 539506 388648 539562 388657
rect 539506 388583 539562 388592
rect 539520 373289 539548 388583
rect 539506 373280 539562 373289
rect 539506 373215 539562 373224
rect 539508 365696 539560 365702
rect 539506 365664 539508 365673
rect 539560 365664 539562 365673
rect 539506 365599 539562 365608
rect 539414 350704 539470 350713
rect 539414 350639 539470 350648
rect 539612 346497 539640 700878
rect 539692 700868 539744 700874
rect 539692 700810 539744 700816
rect 539704 353161 539732 700810
rect 539784 700800 539836 700806
rect 539784 700742 539836 700748
rect 539796 359553 539824 700742
rect 539968 700596 540020 700602
rect 539968 700538 540020 700544
rect 539876 700528 539928 700534
rect 539876 700470 539928 700476
rect 539888 369617 539916 700470
rect 539980 372065 540008 700538
rect 540060 700460 540112 700466
rect 540060 700402 540112 700408
rect 540072 378049 540100 700402
rect 540152 700392 540204 700398
rect 540152 700334 540204 700340
rect 540164 382129 540192 700334
rect 541072 700324 541124 700330
rect 541072 700266 541124 700272
rect 540244 652792 540296 652798
rect 540244 652734 540296 652740
rect 540256 394777 540284 652734
rect 540336 620288 540388 620294
rect 540336 620230 540388 620236
rect 540242 394768 540298 394777
rect 540242 394703 540298 394712
rect 540150 382120 540206 382129
rect 540150 382055 540206 382064
rect 540058 378040 540114 378049
rect 540058 377975 540114 377984
rect 539966 372056 540022 372065
rect 539966 371991 540022 372000
rect 539874 369608 539930 369617
rect 539874 369543 539930 369552
rect 540348 363089 540376 620230
rect 540980 495508 541032 495514
rect 540980 495450 541032 495456
rect 540612 480276 540664 480282
rect 540612 480218 540664 480224
rect 540520 479528 540572 479534
rect 540520 479470 540572 479476
rect 540426 447400 540482 447409
rect 540426 447335 540482 447344
rect 540334 363080 540390 363089
rect 540334 363015 540390 363024
rect 539782 359544 539838 359553
rect 539782 359479 539838 359488
rect 539690 353152 539746 353161
rect 539690 353087 539746 353096
rect 539966 348936 540022 348945
rect 539966 348871 540022 348880
rect 539598 346488 539654 346497
rect 539598 346423 539654 346432
rect 539322 344312 539378 344321
rect 539322 344247 539378 344256
rect 539980 339522 540008 348871
rect 539784 339516 539836 339522
rect 539784 339458 539836 339464
rect 539968 339516 540020 339522
rect 539968 339458 540020 339464
rect 539796 331265 539824 339458
rect 539782 331256 539838 331265
rect 539782 331191 539838 331200
rect 539322 292768 539378 292777
rect 539322 292703 539378 292712
rect 539336 292097 539364 292703
rect 539322 292088 539378 292097
rect 539322 292023 539378 292032
rect 539874 291952 539930 291961
rect 539874 291887 539930 291896
rect 539322 286648 539378 286657
rect 539322 286583 539378 286592
rect 539336 265033 539364 286583
rect 539888 279177 539916 291887
rect 539874 279168 539930 279177
rect 539874 279103 539930 279112
rect 539782 273456 539838 273465
rect 539782 273391 539838 273400
rect 539796 265033 539824 273391
rect 539322 265024 539378 265033
rect 539322 264959 539378 264968
rect 539782 265024 539838 265033
rect 539782 264959 539838 264968
rect 289820 240712 289872 240718
rect 273272 240650 273392 240666
rect 289820 240654 289872 240660
rect 299388 240712 299440 240718
rect 299388 240654 299440 240660
rect 318800 240712 318852 240718
rect 318800 240654 318852 240660
rect 328368 240712 328420 240718
rect 357440 240712 357492 240718
rect 328368 240654 328420 240660
rect 357438 240680 357440 240689
rect 367008 240712 367060 240718
rect 357492 240680 357494 240689
rect 270408 240644 270460 240650
rect 270408 240586 270460 240592
rect 273260 240644 273404 240650
rect 273312 240638 273352 240644
rect 273260 240586 273312 240592
rect 273352 240586 273404 240592
rect 270420 240446 270448 240586
rect 289832 240582 289860 240654
rect 299400 240582 299428 240654
rect 318812 240582 318840 240654
rect 328380 240582 328408 240654
rect 357438 240615 357494 240624
rect 366914 240680 366970 240689
rect 366970 240660 367008 240666
rect 366970 240654 367060 240660
rect 368020 240712 368072 240718
rect 368020 240654 368072 240660
rect 366970 240638 367048 240654
rect 366914 240615 366970 240624
rect 289820 240576 289872 240582
rect 289820 240518 289872 240524
rect 299388 240576 299440 240582
rect 299388 240518 299440 240524
rect 318800 240576 318852 240582
rect 318800 240518 318852 240524
rect 328368 240576 328420 240582
rect 328368 240518 328420 240524
rect 260840 240440 260892 240446
rect 260840 240382 260892 240388
rect 261116 240440 261168 240446
rect 261116 240382 261168 240388
rect 270408 240440 270460 240446
rect 270408 240382 270460 240388
rect 257988 240168 258040 240174
rect 257988 240110 258040 240116
rect 261220 238542 261248 240108
rect 263704 238610 263732 240108
rect 263692 238604 263744 238610
rect 263692 238546 263744 238552
rect 261208 238536 261260 238542
rect 261208 238478 261260 238484
rect 266280 238066 266308 240108
rect 268870 240094 269068 240122
rect 271446 240094 271828 240122
rect 274022 240094 274588 240122
rect 266268 238060 266320 238066
rect 266268 238002 266320 238008
rect 269040 203833 269068 240094
rect 271800 203969 271828 240094
rect 274560 204105 274588 240094
rect 276584 237454 276612 240108
rect 279160 237454 279188 240108
rect 281736 237454 281764 240108
rect 284312 238270 284340 240108
rect 284300 238264 284352 238270
rect 284300 238206 284352 238212
rect 286888 238202 286916 240108
rect 289464 238338 289492 240108
rect 289452 238332 289504 238338
rect 289452 238274 289504 238280
rect 286876 238196 286928 238202
rect 286876 238138 286928 238144
rect 292040 238134 292068 240108
rect 294524 238406 294552 240108
rect 297100 238474 297128 240108
rect 297824 238604 297876 238610
rect 297824 238546 297876 238552
rect 297364 238536 297416 238542
rect 297364 238478 297416 238484
rect 297088 238468 297140 238474
rect 297088 238410 297140 238416
rect 294512 238400 294564 238406
rect 294512 238342 294564 238348
rect 292028 238128 292080 238134
rect 292028 238070 292080 238076
rect 276572 237448 276624 237454
rect 276572 237390 276624 237396
rect 277308 237448 277360 237454
rect 277308 237390 277360 237396
rect 279148 237448 279200 237454
rect 279148 237390 279200 237396
rect 280068 237448 280120 237454
rect 280068 237390 280120 237396
rect 281724 237448 281776 237454
rect 281724 237390 281776 237396
rect 282828 237448 282880 237454
rect 282828 237390 282880 237396
rect 277320 204241 277348 237390
rect 277306 204232 277362 204241
rect 277306 204167 277362 204176
rect 274546 204096 274602 204105
rect 274546 204031 274602 204040
rect 271786 203960 271842 203969
rect 271786 203895 271842 203904
rect 269026 203824 269082 203833
rect 269026 203759 269082 203768
rect 280080 202978 280108 237390
rect 282840 204202 282868 237390
rect 282828 204196 282880 204202
rect 282828 204138 282880 204144
rect 280068 202972 280120 202978
rect 280068 202914 280120 202920
rect 297376 202842 297404 238478
rect 297364 202836 297416 202842
rect 297364 202778 297416 202784
rect 297836 111761 297864 238546
rect 299676 237454 299704 240108
rect 302252 237454 302280 240108
rect 304842 240094 304948 240122
rect 307418 240094 307708 240122
rect 309994 240094 310468 240122
rect 312570 240094 313228 240122
rect 299664 237448 299716 237454
rect 299664 237390 299716 237396
rect 300768 237448 300820 237454
rect 300768 237390 300820 237396
rect 302240 237448 302292 237454
rect 302240 237390 302292 237396
rect 303528 237448 303580 237454
rect 303528 237390 303580 237396
rect 300780 204134 300808 237390
rect 300768 204128 300820 204134
rect 300768 204070 300820 204076
rect 303540 204066 303568 237390
rect 303528 204060 303580 204066
rect 303528 204002 303580 204008
rect 304920 203998 304948 240094
rect 304908 203992 304960 203998
rect 304908 203934 304960 203940
rect 307680 203930 307708 240094
rect 307668 203924 307720 203930
rect 307668 203866 307720 203872
rect 310440 203862 310468 240094
rect 310428 203856 310480 203862
rect 310428 203798 310480 203804
rect 313200 203794 313228 240094
rect 315132 237454 315160 240108
rect 317708 237454 317736 240108
rect 320284 237454 320312 240108
rect 315120 237448 315172 237454
rect 315120 237390 315172 237396
rect 315948 237448 316000 237454
rect 315948 237390 316000 237396
rect 317696 237448 317748 237454
rect 317696 237390 317748 237396
rect 318708 237448 318760 237454
rect 318708 237390 318760 237396
rect 320272 237448 320324 237454
rect 320272 237390 320324 237396
rect 321468 237448 321520 237454
rect 321468 237390 321520 237396
rect 313188 203788 313240 203794
rect 313188 203730 313240 203736
rect 315960 202910 315988 237390
rect 318720 203658 318748 237390
rect 318708 203652 318760 203658
rect 318708 203594 318760 203600
rect 321480 203590 321508 237390
rect 321468 203584 321520 203590
rect 321468 203526 321520 203532
rect 322860 203522 322888 240108
rect 325344 238678 325372 240108
rect 327934 240094 328316 240122
rect 330510 240094 331076 240122
rect 325332 238672 325384 238678
rect 325332 238614 325384 238620
rect 322848 203516 322900 203522
rect 322848 203458 322900 203464
rect 328288 203386 328316 240094
rect 329748 238604 329800 238610
rect 329748 238546 329800 238552
rect 328368 238536 328420 238542
rect 328368 238478 328420 238484
rect 328380 203697 328408 238478
rect 329760 203697 329788 238546
rect 331048 204270 331076 240094
rect 331128 238740 331180 238746
rect 331128 238682 331180 238688
rect 331036 204264 331088 204270
rect 331036 204206 331088 204212
rect 331140 203697 331168 238682
rect 332508 237584 332560 237590
rect 332508 237526 332560 237532
rect 332324 203788 332376 203794
rect 332324 203730 332376 203736
rect 332416 203788 332468 203794
rect 332416 203730 332468 203736
rect 328366 203688 328422 203697
rect 328366 203623 328422 203632
rect 329746 203688 329802 203697
rect 329746 203623 329802 203632
rect 331126 203688 331182 203697
rect 331126 203623 331182 203632
rect 328368 203448 328420 203454
rect 328366 203416 328368 203425
rect 328420 203416 328422 203425
rect 328276 203380 328328 203386
rect 328366 203351 328422 203360
rect 328276 203322 328328 203328
rect 331128 203312 331180 203318
rect 331126 203280 331128 203289
rect 331180 203280 331182 203289
rect 329748 203244 329800 203250
rect 331126 203215 331182 203224
rect 329748 203186 329800 203192
rect 329760 203153 329788 203186
rect 329746 203144 329802 203153
rect 332336 203114 332364 203730
rect 332428 203425 332456 203730
rect 332414 203416 332470 203425
rect 332414 203351 332470 203360
rect 332520 203289 332548 237526
rect 333072 237454 333100 240108
rect 335648 237522 335676 240108
rect 336740 238672 336792 238678
rect 336740 238614 336792 238620
rect 333888 237516 333940 237522
rect 333888 237458 333940 237464
rect 335636 237516 335688 237522
rect 335636 237458 335688 237464
rect 333060 237448 333112 237454
rect 333060 237390 333112 237396
rect 333900 203425 333928 237458
rect 333980 237448 334032 237454
rect 333980 237390 334032 237396
rect 333886 203416 333942 203425
rect 333886 203351 333942 203360
rect 333888 203312 333940 203318
rect 332506 203280 332562 203289
rect 333992 203289 334020 237390
rect 334072 204264 334124 204270
rect 334072 204206 334124 204212
rect 336372 204264 336424 204270
rect 336372 204206 336424 204212
rect 334084 203697 334112 204206
rect 336384 203794 336412 204206
rect 336372 203788 336424 203794
rect 336372 203730 336424 203736
rect 336464 203788 336516 203794
rect 336464 203730 336516 203736
rect 334070 203688 334126 203697
rect 334070 203623 334126 203632
rect 335174 203552 335230 203561
rect 335174 203487 335230 203496
rect 333888 203254 333940 203260
rect 333978 203280 334034 203289
rect 332506 203215 332562 203224
rect 333900 203153 333928 203254
rect 335188 203250 335216 203487
rect 335360 203380 335412 203386
rect 335360 203322 335412 203328
rect 335372 203289 335400 203322
rect 335358 203280 335414 203289
rect 333978 203215 334034 203224
rect 335176 203244 335228 203250
rect 335176 203186 335228 203192
rect 335268 203244 335320 203250
rect 335358 203215 335414 203224
rect 335268 203186 335320 203192
rect 335280 203153 335308 203186
rect 333886 203144 333942 203153
rect 329746 203079 329802 203088
rect 332324 203108 332376 203114
rect 333886 203079 333942 203088
rect 335266 203144 335322 203153
rect 336476 203114 336504 203730
rect 336646 203416 336702 203425
rect 336646 203351 336648 203360
rect 336700 203351 336702 203360
rect 336648 203322 336700 203328
rect 336752 203289 336780 238614
rect 338224 237590 338252 240108
rect 340800 238746 340828 240108
rect 340788 238740 340840 238746
rect 340788 238682 340840 238688
rect 343376 238610 343404 240108
rect 343364 238604 343416 238610
rect 343364 238546 343416 238552
rect 345952 238542 345980 240108
rect 348542 240094 349108 240122
rect 345940 238536 345992 238542
rect 345940 238478 345992 238484
rect 347044 238468 347096 238474
rect 347044 238410 347096 238416
rect 344284 238400 344336 238406
rect 344284 238342 344336 238348
rect 341524 238332 341576 238338
rect 341524 238274 341576 238280
rect 338764 238264 338816 238270
rect 338764 238206 338816 238212
rect 338212 237584 338264 237590
rect 338212 237526 338264 237532
rect 338120 203516 338172 203522
rect 338120 203458 338172 203464
rect 338212 203516 338264 203522
rect 338212 203458 338264 203464
rect 337936 203448 337988 203454
rect 338132 203425 338160 203458
rect 337936 203390 337988 203396
rect 338118 203416 338174 203425
rect 336738 203280 336794 203289
rect 336738 203215 336794 203224
rect 335266 203079 335322 203088
rect 336464 203108 336516 203114
rect 332324 203050 332376 203056
rect 336464 203050 336516 203056
rect 336648 203108 336700 203114
rect 336648 203050 336700 203056
rect 336660 203017 336688 203050
rect 337948 203017 337976 203390
rect 338118 203351 338174 203360
rect 338224 203182 338252 203458
rect 338776 203182 338804 238206
rect 340144 238196 340196 238202
rect 340144 238138 340196 238144
rect 340156 203794 340184 238138
rect 340052 203788 340104 203794
rect 340052 203730 340104 203736
rect 340144 203788 340196 203794
rect 340144 203730 340196 203736
rect 340064 203674 340092 203730
rect 340788 203720 340840 203726
rect 340064 203668 340788 203674
rect 340064 203662 340840 203668
rect 340064 203646 340828 203662
rect 340880 203652 340932 203658
rect 340880 203594 340932 203600
rect 339408 203584 339460 203590
rect 340892 203561 340920 203594
rect 339590 203552 339646 203561
rect 339460 203532 339540 203538
rect 339408 203526 339540 203532
rect 339224 203516 339276 203522
rect 339420 203510 339540 203526
rect 339224 203458 339276 203464
rect 338212 203176 338264 203182
rect 338212 203118 338264 203124
rect 338764 203176 338816 203182
rect 338764 203118 338816 203124
rect 339236 203017 339264 203458
rect 339512 203289 339540 203510
rect 339590 203487 339592 203496
rect 339644 203487 339646 203496
rect 340878 203552 340934 203561
rect 340878 203487 340934 203496
rect 339592 203458 339644 203464
rect 339498 203280 339554 203289
rect 339498 203215 339554 203224
rect 341536 203046 341564 238274
rect 342168 204264 342220 204270
rect 342168 204206 342220 204212
rect 342180 203153 342208 204206
rect 343824 204060 343876 204066
rect 343824 204002 343876 204008
rect 343836 203862 343864 204002
rect 344296 203998 344324 238342
rect 345756 238128 345808 238134
rect 345756 238070 345808 238076
rect 345664 238060 345716 238066
rect 345664 238002 345716 238008
rect 345388 204332 345440 204338
rect 345388 204274 345440 204280
rect 345296 204264 345348 204270
rect 345296 204206 345348 204212
rect 345308 204134 345336 204206
rect 345400 204202 345428 204274
rect 345388 204196 345440 204202
rect 345388 204138 345440 204144
rect 345296 204128 345348 204134
rect 345296 204070 345348 204076
rect 344284 203992 344336 203998
rect 344284 203934 344336 203940
rect 345676 203930 345704 238002
rect 345768 204134 345796 238070
rect 345756 204128 345808 204134
rect 345756 204070 345808 204076
rect 346400 204060 346452 204066
rect 346400 204002 346452 204008
rect 345020 203924 345072 203930
rect 345020 203866 345072 203872
rect 345664 203924 345716 203930
rect 345664 203866 345716 203872
rect 343640 203856 343692 203862
rect 343640 203798 343692 203804
rect 343824 203856 343876 203862
rect 343824 203798 343876 203804
rect 342260 203720 342312 203726
rect 342258 203688 342260 203697
rect 343652 203697 343680 203798
rect 344928 203720 344980 203726
rect 342312 203688 342314 203697
rect 342258 203623 342314 203632
rect 343638 203688 343694 203697
rect 344928 203662 344980 203668
rect 343638 203623 343694 203632
rect 342444 203312 342496 203318
rect 342444 203254 342496 203260
rect 342166 203144 342222 203153
rect 342166 203079 342222 203088
rect 341524 203040 341576 203046
rect 336646 203008 336702 203017
rect 336646 202943 336702 202952
rect 337934 203008 337990 203017
rect 337934 202943 337990 202952
rect 339222 203008 339278 203017
rect 341524 202982 341576 202988
rect 339222 202943 339278 202952
rect 315948 202904 316000 202910
rect 315948 202846 316000 202852
rect 342180 202842 342208 203079
rect 342456 203017 342484 203254
rect 343640 203244 343692 203250
rect 343640 203186 343692 203192
rect 343652 203017 343680 203186
rect 344940 203114 344968 203662
rect 345032 203289 345060 203866
rect 345940 203380 345992 203386
rect 345940 203322 345992 203328
rect 345018 203280 345074 203289
rect 345018 203215 345074 203224
rect 344928 203108 344980 203114
rect 344928 203050 344980 203056
rect 344940 203017 344968 203050
rect 345952 203017 345980 203322
rect 346412 203153 346440 204002
rect 346768 203584 346820 203590
rect 346952 203584 347004 203590
rect 346820 203532 346952 203538
rect 346768 203526 347004 203532
rect 346780 203510 346992 203526
rect 347056 203454 347084 238410
rect 347780 203856 347832 203862
rect 347780 203798 347832 203804
rect 347136 203516 347188 203522
rect 347136 203458 347188 203464
rect 347044 203448 347096 203454
rect 347044 203390 347096 203396
rect 346398 203144 346454 203153
rect 346398 203079 346454 203088
rect 347148 203017 347176 203458
rect 347792 203153 347820 203798
rect 348332 203584 348384 203590
rect 349080 203561 349108 240094
rect 351104 237454 351132 240108
rect 353680 238066 353708 240108
rect 356164 238134 356192 240108
rect 356152 238128 356204 238134
rect 356152 238070 356204 238076
rect 353668 238060 353720 238066
rect 353668 238002 353720 238008
rect 351092 237448 351144 237454
rect 351092 237390 351144 237396
rect 351828 237448 351880 237454
rect 351828 237390 351880 237396
rect 349160 204264 349212 204270
rect 349160 204206 349212 204212
rect 349172 203697 349200 204206
rect 349252 204060 349304 204066
rect 349252 204002 349304 204008
rect 349158 203688 349214 203697
rect 349264 203658 349292 204002
rect 351092 203992 351144 203998
rect 351092 203934 351144 203940
rect 351736 203992 351788 203998
rect 351736 203934 351788 203940
rect 351104 203697 351132 203934
rect 351090 203688 351146 203697
rect 349158 203623 349214 203632
rect 349252 203652 349304 203658
rect 349252 203594 349304 203600
rect 349344 203652 349396 203658
rect 349344 203594 349396 203600
rect 351000 203652 351052 203658
rect 351090 203623 351146 203632
rect 351000 203594 351052 203600
rect 348332 203526 348384 203532
rect 349066 203552 349122 203561
rect 347778 203144 347834 203153
rect 347778 203079 347834 203088
rect 348344 203017 348372 203526
rect 349066 203487 349122 203496
rect 349160 203448 349212 203454
rect 349160 203390 349212 203396
rect 349172 203289 349200 203390
rect 349158 203280 349214 203289
rect 349158 203215 349214 203224
rect 349264 203017 349292 203594
rect 342258 203008 342314 203017
rect 342258 202943 342314 202952
rect 342442 203008 342498 203017
rect 342442 202943 342498 202952
rect 343638 203008 343694 203017
rect 343638 202943 343694 202952
rect 344926 203008 344982 203017
rect 344926 202943 344982 202952
rect 345938 203008 345994 203017
rect 345938 202943 345994 202952
rect 347134 203008 347190 203017
rect 347134 202943 347190 202952
rect 348330 203008 348386 203017
rect 348330 202943 348386 202952
rect 349250 203008 349306 203017
rect 349250 202943 349306 202952
rect 342272 202910 342300 202943
rect 349356 202910 349384 203594
rect 351012 203114 351040 203594
rect 351748 203318 351776 203934
rect 351840 203697 351868 237390
rect 357440 204196 357492 204202
rect 357440 204138 357492 204144
rect 351920 204128 351972 204134
rect 351920 204070 351972 204076
rect 351826 203688 351882 203697
rect 351826 203623 351882 203632
rect 351736 203312 351788 203318
rect 351736 203254 351788 203260
rect 351000 203108 351052 203114
rect 351000 203050 351052 203056
rect 351012 203017 351040 203050
rect 351748 203017 351776 203254
rect 351932 203153 351960 204070
rect 354680 203788 354732 203794
rect 354680 203730 354732 203736
rect 355600 203788 355652 203794
rect 355600 203730 355652 203736
rect 354312 203720 354364 203726
rect 354312 203662 354364 203668
rect 353208 203652 353260 203658
rect 353208 203594 353260 203600
rect 353220 203250 353248 203594
rect 353208 203244 353260 203250
rect 353208 203186 353260 203192
rect 353220 203153 353248 203186
rect 351918 203144 351974 203153
rect 351918 203079 351974 203088
rect 353206 203144 353262 203153
rect 353206 203079 353262 203088
rect 353300 203040 353352 203046
rect 350998 203008 351054 203017
rect 350998 202943 351054 202952
rect 351734 203008 351790 203017
rect 351734 202943 351790 202952
rect 353298 203008 353300 203017
rect 354324 203017 354352 203662
rect 354692 203153 354720 203730
rect 355612 203386 355640 203730
rect 356428 203448 356480 203454
rect 357452 203425 357480 204138
rect 357532 204060 357584 204066
rect 357532 204002 357584 204008
rect 356428 203390 356480 203396
rect 357438 203416 357494 203425
rect 355600 203380 355652 203386
rect 355600 203322 355652 203328
rect 354678 203144 354734 203153
rect 354678 203079 354734 203088
rect 355612 203017 355640 203322
rect 356060 203176 356112 203182
rect 356058 203144 356060 203153
rect 356112 203144 356114 203153
rect 356058 203079 356114 203088
rect 356440 203017 356468 203390
rect 357438 203351 357494 203360
rect 357544 203318 357572 204002
rect 357808 203584 357860 203590
rect 357808 203526 357860 203532
rect 357532 203312 357584 203318
rect 357532 203254 357584 203260
rect 357820 203153 357848 203526
rect 358740 203386 358768 240108
rect 361316 237454 361344 240108
rect 363906 240094 364288 240122
rect 361304 237448 361356 237454
rect 361304 237390 361356 237396
rect 362224 237448 362276 237454
rect 362224 237390 362276 237396
rect 362236 204202 362264 237390
rect 364260 204270 364288 240094
rect 366376 240094 366482 240122
rect 368032 240106 368060 240654
rect 368020 240100 368072 240106
rect 364248 204264 364300 204270
rect 364248 204206 364300 204212
rect 365720 204264 365772 204270
rect 366376 204241 366404 240094
rect 369058 240094 369808 240122
rect 368020 240042 368072 240048
rect 369780 204950 369808 240094
rect 371148 238400 371200 238406
rect 371148 238342 371200 238348
rect 369768 204944 369820 204950
rect 369768 204886 369820 204892
rect 371160 204241 371188 238342
rect 371620 237454 371648 240108
rect 373264 240100 373316 240106
rect 373264 240042 373316 240048
rect 371608 237448 371660 237454
rect 371608 237390 371660 237396
rect 372528 237448 372580 237454
rect 372528 237390 372580 237396
rect 365720 204206 365772 204212
rect 366362 204232 366418 204241
rect 362224 204196 362276 204202
rect 362224 204138 362276 204144
rect 360016 204060 360068 204066
rect 360016 204002 360068 204008
rect 358728 203380 358780 203386
rect 358728 203322 358780 203328
rect 358636 203312 358688 203318
rect 358636 203254 358688 203260
rect 357806 203144 357862 203153
rect 357806 203079 357862 203088
rect 358648 203017 358676 203254
rect 360028 203114 360056 204002
rect 361304 203992 361356 203998
rect 365732 203969 365760 204206
rect 371146 204232 371202 204241
rect 366362 204167 366418 204176
rect 367100 204196 367152 204202
rect 371146 204167 371202 204176
rect 367100 204138 367152 204144
rect 367112 204105 367140 204138
rect 367098 204096 367154 204105
rect 367098 204031 367154 204040
rect 361304 203934 361356 203940
rect 365718 203960 365774 203969
rect 360016 203108 360068 203114
rect 360016 203050 360068 203056
rect 360028 203017 360056 203050
rect 361316 203017 361344 203934
rect 364340 203924 364392 203930
rect 365718 203895 365774 203904
rect 364340 203866 364392 203872
rect 363512 203856 363564 203862
rect 364352 203833 364380 203866
rect 363512 203798 363564 203804
rect 364338 203824 364394 203833
rect 362500 203652 362552 203658
rect 362500 203594 362552 203600
rect 362512 203017 362540 203594
rect 363524 203017 363552 203798
rect 364338 203759 364394 203768
rect 364708 203788 364760 203794
rect 364708 203730 364760 203736
rect 364720 203017 364748 203730
rect 368480 203380 368532 203386
rect 368480 203322 368532 203328
rect 368492 203289 368520 203322
rect 368478 203280 368534 203289
rect 368478 203215 368534 203224
rect 353352 203008 353354 203017
rect 353298 202943 353354 202952
rect 354310 203008 354366 203017
rect 354310 202943 354366 202952
rect 355598 203008 355654 203017
rect 355598 202943 355654 202952
rect 356426 203008 356482 203017
rect 356426 202943 356482 202952
rect 357438 203008 357494 203017
rect 357438 202943 357440 202952
rect 357492 202943 357494 202952
rect 358634 203008 358690 203017
rect 358634 202943 358690 202952
rect 360014 203008 360070 203017
rect 360014 202943 360070 202952
rect 361302 203008 361358 203017
rect 361302 202943 361358 202952
rect 362498 203008 362554 203017
rect 362498 202943 362554 202952
rect 363510 203008 363566 203017
rect 363510 202943 363566 202952
rect 364706 203008 364762 203017
rect 364706 202943 364762 202952
rect 357440 202914 357492 202920
rect 342260 202904 342312 202910
rect 342260 202846 342312 202852
rect 349344 202904 349396 202910
rect 349344 202846 349396 202852
rect 297916 202836 297968 202842
rect 297916 202778 297968 202784
rect 342168 202836 342220 202842
rect 342168 202778 342220 202784
rect 297928 201550 297956 202778
rect 297916 201544 297968 201550
rect 297916 201486 297968 201492
rect 297928 180305 297956 201486
rect 372540 200938 372568 237390
rect 373276 203153 373304 240042
rect 374196 237454 374224 240108
rect 376772 237454 376800 240108
rect 379362 240094 379468 240122
rect 381938 240094 382228 240122
rect 374184 237448 374236 237454
rect 374184 237390 374236 237396
rect 375288 237448 375340 237454
rect 375288 237390 375340 237396
rect 376760 237448 376812 237454
rect 376760 237390 376812 237396
rect 378048 237448 378100 237454
rect 378048 237390 378100 237396
rect 373262 203144 373318 203153
rect 373262 203079 373318 203088
rect 375300 201006 375328 237390
rect 378060 201074 378088 237390
rect 379440 201142 379468 240094
rect 380348 238536 380400 238542
rect 380348 238478 380400 238484
rect 380256 238468 380308 238474
rect 380256 238410 380308 238416
rect 380164 238196 380216 238202
rect 380164 238138 380216 238144
rect 379428 201136 379480 201142
rect 379428 201078 379480 201084
rect 378048 201068 378100 201074
rect 378048 201010 378100 201016
rect 375288 201000 375340 201006
rect 375288 200942 375340 200948
rect 372528 200932 372580 200938
rect 372528 200874 372580 200880
rect 379796 183524 379848 183530
rect 379796 183466 379848 183472
rect 379808 182753 379836 183466
rect 379794 182744 379850 182753
rect 379794 182679 379850 182688
rect 297914 180296 297970 180305
rect 297914 180231 297970 180240
rect 297914 171864 297970 171873
rect 297914 171799 297970 171808
rect 297822 111752 297878 111761
rect 297822 111687 297878 111696
rect 297928 108934 297956 171799
rect 380176 137970 380204 238138
rect 380072 137964 380124 137970
rect 380072 137906 380124 137912
rect 380164 137964 380216 137970
rect 380164 137906 380216 137912
rect 380084 135250 380112 137906
rect 379796 135244 379848 135250
rect 379796 135186 379848 135192
rect 380072 135244 380124 135250
rect 380072 135186 380124 135192
rect 379808 125633 379836 135186
rect 379794 125624 379850 125633
rect 379794 125559 379850 125568
rect 379978 125624 380034 125633
rect 379978 125559 380034 125568
rect 379992 119241 380020 125559
rect 380268 120329 380296 238410
rect 380360 122097 380388 238478
rect 380440 238332 380492 238338
rect 380440 238274 380492 238280
rect 380452 180985 380480 238274
rect 382200 202162 382228 240094
rect 384500 238270 384528 240108
rect 384488 238264 384540 238270
rect 384488 238206 384540 238212
rect 386984 237454 387012 240108
rect 388444 238604 388496 238610
rect 388444 238546 388496 238552
rect 386972 237448 387024 237454
rect 386972 237390 387024 237396
rect 387708 237448 387760 237454
rect 387708 237390 387760 237396
rect 387720 202230 387748 237390
rect 387708 202224 387760 202230
rect 387708 202166 387760 202172
rect 382188 202156 382240 202162
rect 382188 202098 382240 202104
rect 380438 180976 380494 180985
rect 380438 180911 380494 180920
rect 380808 124160 380860 124166
rect 380808 124102 380860 124108
rect 380820 123185 380848 124102
rect 380806 123176 380862 123185
rect 380806 123111 380862 123120
rect 380346 122088 380402 122097
rect 380346 122023 380402 122032
rect 380254 120320 380310 120329
rect 380254 120255 380310 120264
rect 379978 119232 380034 119241
rect 379978 119167 380034 119176
rect 388456 118454 388484 238546
rect 389560 238406 389588 240108
rect 391952 240094 392150 240122
rect 391204 238672 391256 238678
rect 391204 238614 391256 238620
rect 389548 238400 389600 238406
rect 389548 238342 389600 238348
rect 380808 118448 380860 118454
rect 380808 118390 380860 118396
rect 388444 118448 388496 118454
rect 388444 118390 388496 118396
rect 380820 118153 380848 118390
rect 380806 118144 380862 118153
rect 380806 118079 380862 118088
rect 380716 115932 380768 115938
rect 380716 115874 380768 115880
rect 380728 114753 380756 115874
rect 391216 115870 391244 238614
rect 391952 124166 391980 240094
rect 394712 238542 394740 240108
rect 394700 238536 394752 238542
rect 394700 238478 394752 238484
rect 397288 238474 397316 240108
rect 397276 238468 397328 238474
rect 397276 238410 397328 238416
rect 393964 238400 394016 238406
rect 393964 238342 394016 238348
rect 391940 124160 391992 124166
rect 391940 124102 391992 124108
rect 393976 115938 394004 238342
rect 399864 238202 399892 240108
rect 402440 238610 402468 240108
rect 405016 238678 405044 240108
rect 405004 238672 405056 238678
rect 405004 238614 405056 238620
rect 402428 238604 402480 238610
rect 402428 238546 402480 238552
rect 407592 238406 407620 240108
rect 409892 240094 410182 240122
rect 407580 238400 407632 238406
rect 407580 238342 407632 238348
rect 399852 238196 399904 238202
rect 399852 238138 399904 238144
rect 409892 202842 409920 240094
rect 412744 238202 412772 240108
rect 415320 238338 415348 240108
rect 417804 238474 417832 240108
rect 420380 238542 420408 240108
rect 420368 238536 420420 238542
rect 420368 238478 420420 238484
rect 417792 238468 417844 238474
rect 417792 238410 417844 238416
rect 422956 238406 422984 240108
rect 422944 238400 422996 238406
rect 422944 238342 422996 238348
rect 425532 238338 425560 240108
rect 428108 238610 428136 240108
rect 430684 238678 430712 240108
rect 433260 238746 433288 240108
rect 433248 238740 433300 238746
rect 433248 238682 433300 238688
rect 430672 238672 430724 238678
rect 430672 238614 430724 238620
rect 428096 238604 428148 238610
rect 428096 238546 428148 238552
rect 415308 238332 415360 238338
rect 415308 238274 415360 238280
rect 425520 238332 425572 238338
rect 425520 238274 425572 238280
rect 412732 238196 412784 238202
rect 412732 238138 412784 238144
rect 435836 237998 435864 240108
rect 437492 240094 438426 240122
rect 440252 240094 441002 240122
rect 443012 240094 443578 240122
rect 445772 240094 446154 240122
rect 448532 240094 448638 240122
rect 449912 240094 451214 240122
rect 452672 240094 453790 240122
rect 455432 240094 456366 240122
rect 435824 237992 435876 237998
rect 435824 237934 435876 237940
rect 437492 203794 437520 240094
rect 440252 203862 440280 240094
rect 440240 203856 440292 203862
rect 440240 203798 440292 203804
rect 437480 203788 437532 203794
rect 437480 203730 437532 203736
rect 443012 203658 443040 240094
rect 445772 203998 445800 240094
rect 447784 238264 447836 238270
rect 447784 238206 447836 238212
rect 445760 203992 445812 203998
rect 445760 203934 445812 203940
rect 443000 203652 443052 203658
rect 443000 203594 443052 203600
rect 409880 202836 409932 202842
rect 409880 202778 409932 202784
rect 410524 202836 410576 202842
rect 410524 202778 410576 202784
rect 410536 201618 410564 202778
rect 410524 201612 410576 201618
rect 410524 201554 410576 201560
rect 410536 183530 410564 201554
rect 417424 201544 417476 201550
rect 417424 201486 417476 201492
rect 410524 183524 410576 183530
rect 410524 183466 410576 183472
rect 417436 180577 417464 201486
rect 447796 201210 447824 238206
rect 447876 237992 447928 237998
rect 447876 237934 447928 237940
rect 447888 203794 447916 237934
rect 448532 204066 448560 240094
rect 449164 238740 449216 238746
rect 449164 238682 449216 238688
rect 449176 204066 449204 238682
rect 449808 204128 449860 204134
rect 449806 204096 449808 204105
rect 449860 204096 449862 204105
rect 448520 204060 448572 204066
rect 448520 204002 448572 204008
rect 449164 204060 449216 204066
rect 449806 204031 449862 204040
rect 449164 204002 449216 204008
rect 447876 203788 447928 203794
rect 447876 203730 447928 203736
rect 448428 203788 448480 203794
rect 448428 203730 448480 203736
rect 448440 201521 448468 203730
rect 449176 203425 449204 204002
rect 449162 203416 449218 203425
rect 449162 203351 449218 203360
rect 449912 203318 449940 240094
rect 450544 238672 450596 238678
rect 450544 238614 450596 238620
rect 450556 203930 450584 238614
rect 451924 238604 451976 238610
rect 451924 238546 451976 238552
rect 451188 238264 451240 238270
rect 451188 238206 451240 238212
rect 450544 203924 450596 203930
rect 450544 203866 450596 203872
rect 450556 203425 450584 203866
rect 450542 203416 450598 203425
rect 450542 203351 450598 203360
rect 449900 203312 449952 203318
rect 451200 203289 451228 238206
rect 451936 203862 451964 238546
rect 451924 203856 451976 203862
rect 451924 203798 451976 203804
rect 451936 203425 451964 203798
rect 452672 203590 452700 240094
rect 454684 238400 454736 238406
rect 454684 238342 454736 238348
rect 455236 238400 455288 238406
rect 455236 238342 455288 238348
rect 453304 238332 453356 238338
rect 453304 238274 453356 238280
rect 453948 238332 454000 238338
rect 453948 238274 454000 238280
rect 452660 203584 452712 203590
rect 452660 203526 452712 203532
rect 453316 203425 453344 238274
rect 451922 203416 451978 203425
rect 451922 203351 451978 203360
rect 453302 203416 453358 203425
rect 453302 203351 453358 203360
rect 449900 203254 449952 203260
rect 451186 203280 451242 203289
rect 451186 203215 451242 203224
rect 453316 203114 453344 203351
rect 453960 203289 453988 238274
rect 454696 203289 454724 238342
rect 455248 203289 455276 238342
rect 455432 203454 455460 240094
rect 458928 238678 458956 240108
rect 458916 238672 458968 238678
rect 458916 238614 458968 238620
rect 456248 238536 456300 238542
rect 456248 238478 456300 238484
rect 460848 238536 460900 238542
rect 460848 238478 460900 238484
rect 456064 238468 456116 238474
rect 456064 238410 456116 238416
rect 456076 204270 456104 238410
rect 456064 204264 456116 204270
rect 456064 204206 456116 204212
rect 456260 203538 456288 238478
rect 458088 238468 458140 238474
rect 458088 238410 458140 238416
rect 456616 204264 456668 204270
rect 456614 204232 456616 204241
rect 456668 204232 456670 204241
rect 456614 204167 456670 204176
rect 457996 203788 458048 203794
rect 457996 203730 458048 203736
rect 456168 203510 456288 203538
rect 456168 203454 456196 203510
rect 455420 203448 455472 203454
rect 456156 203448 456208 203454
rect 455420 203390 455472 203396
rect 456154 203416 456156 203425
rect 456208 203416 456210 203425
rect 458008 203386 458036 203730
rect 456154 203351 456210 203360
rect 457996 203380 458048 203386
rect 457996 203322 458048 203328
rect 453946 203280 454002 203289
rect 453946 203215 454002 203224
rect 454682 203280 454738 203289
rect 454682 203215 454738 203224
rect 455050 203280 455106 203289
rect 455050 203215 455106 203224
rect 455234 203280 455290 203289
rect 455234 203215 455290 203224
rect 455064 203182 455092 203215
rect 455052 203176 455104 203182
rect 455052 203118 455104 203124
rect 453304 203108 453356 203114
rect 453304 203050 453356 203056
rect 455328 203040 455380 203046
rect 452566 203008 452622 203017
rect 452566 202943 452568 202952
rect 452620 202943 452622 202952
rect 455326 203008 455328 203017
rect 458008 203017 458036 203322
rect 458100 203289 458128 238410
rect 459008 204060 459060 204066
rect 459008 204002 459060 204008
rect 458086 203280 458142 203289
rect 458086 203215 458142 203224
rect 459020 203017 459048 204002
rect 459468 203992 459520 203998
rect 459468 203934 459520 203940
rect 459480 203425 459508 203934
rect 460572 203924 460624 203930
rect 460572 203866 460624 203872
rect 460584 203454 460612 203866
rect 460572 203448 460624 203454
rect 459466 203416 459522 203425
rect 460572 203390 460624 203396
rect 459466 203351 459522 203360
rect 460584 203017 460612 203390
rect 460860 203289 460888 238478
rect 461504 237454 461532 240108
rect 464080 238746 464108 240108
rect 464068 238740 464120 238746
rect 464068 238682 464120 238688
rect 463608 238604 463660 238610
rect 463608 238546 463660 238552
rect 461492 237448 461544 237454
rect 461492 237390 461544 237396
rect 462228 237448 462280 237454
rect 462228 237390 462280 237396
rect 462136 203924 462188 203930
rect 462136 203866 462188 203872
rect 461400 203856 461452 203862
rect 461400 203798 461452 203804
rect 461412 203590 461440 203798
rect 461400 203584 461452 203590
rect 461400 203526 461452 203532
rect 460846 203280 460902 203289
rect 460846 203215 460902 203224
rect 461412 203017 461440 203526
rect 462148 203425 462176 203866
rect 462240 203726 462268 237390
rect 463516 203856 463568 203862
rect 463516 203798 463568 203804
rect 462228 203720 462280 203726
rect 462228 203662 462280 203668
rect 463528 203425 463556 203798
rect 462134 203416 462190 203425
rect 462134 203351 462190 203360
rect 463514 203416 463570 203425
rect 463514 203351 463570 203360
rect 463620 203289 463648 238546
rect 466656 237862 466684 240108
rect 466644 237856 466696 237862
rect 466644 237798 466696 237804
rect 469232 237794 469260 240108
rect 469220 237788 469272 237794
rect 469220 237730 469272 237736
rect 471808 237658 471836 240108
rect 471888 237992 471940 237998
rect 471888 237934 471940 237940
rect 471796 237652 471848 237658
rect 471796 237594 471848 237600
rect 470508 205216 470560 205222
rect 470508 205158 470560 205164
rect 470416 205080 470468 205086
rect 470416 205022 470468 205028
rect 469128 205012 469180 205018
rect 469128 204954 469180 204960
rect 465080 204264 465132 204270
rect 469140 204241 469168 204954
rect 465080 204206 465132 204212
rect 469126 204232 469182 204241
rect 464988 203788 465040 203794
rect 464988 203730 465040 203736
rect 464620 203312 464672 203318
rect 463606 203280 463662 203289
rect 463606 203215 463662 203224
rect 464618 203280 464620 203289
rect 464672 203280 464674 203289
rect 464618 203215 464674 203224
rect 463608 203176 463660 203182
rect 463608 203118 463660 203124
rect 462412 203108 462464 203114
rect 462412 203050 462464 203056
rect 462424 203017 462452 203050
rect 463620 203017 463648 203118
rect 465000 203017 465028 203730
rect 465092 203289 465120 204206
rect 467748 204196 467800 204202
rect 469126 204167 469182 204176
rect 467748 204138 467800 204144
rect 467760 204105 467788 204138
rect 470428 204105 470456 205022
rect 470520 204241 470548 205158
rect 470506 204232 470562 204241
rect 470506 204167 470562 204176
rect 467746 204096 467802 204105
rect 465172 204060 465224 204066
rect 465172 204002 465224 204008
rect 466552 204060 466604 204066
rect 467746 204031 467802 204040
rect 470414 204096 470470 204105
rect 470414 204031 470470 204040
rect 466552 204002 466604 204008
rect 465184 203454 465212 204002
rect 466380 203658 466500 203674
rect 466380 203652 466512 203658
rect 466380 203646 466460 203652
rect 465172 203448 465224 203454
rect 465172 203390 465224 203396
rect 465078 203280 465134 203289
rect 465078 203215 465134 203224
rect 466380 203017 466408 203646
rect 466460 203594 466512 203600
rect 466564 203538 466592 204002
rect 466472 203510 466592 203538
rect 470692 203584 470744 203590
rect 470692 203526 470744 203532
rect 469404 203516 469456 203522
rect 466472 203318 466500 203510
rect 469404 203458 469456 203464
rect 468484 203448 468536 203454
rect 468484 203390 468536 203396
rect 467288 203380 467340 203386
rect 467288 203322 467340 203328
rect 466460 203312 466512 203318
rect 466552 203312 466604 203318
rect 466460 203254 466512 203260
rect 466550 203280 466552 203289
rect 466604 203280 466606 203289
rect 466550 203215 466606 203224
rect 467300 203017 467328 203322
rect 468496 203017 468524 203390
rect 469416 203017 469444 203458
rect 470704 203017 470732 203526
rect 471900 203289 471928 237934
rect 473268 237924 473320 237930
rect 473268 237866 473320 237872
rect 473280 203289 473308 237866
rect 474384 237454 474412 240108
rect 476868 240094 476974 240122
rect 476764 237856 476816 237862
rect 476764 237798 476816 237804
rect 476028 237584 476080 237590
rect 476028 237526 476080 237532
rect 474372 237448 474424 237454
rect 474372 237390 474424 237396
rect 473820 204468 473872 204474
rect 473820 204410 473872 204416
rect 473832 204202 473860 204410
rect 473820 204196 473872 204202
rect 473820 204138 473872 204144
rect 474188 204060 474240 204066
rect 474188 204002 474240 204008
rect 471886 203280 471942 203289
rect 473266 203280 473322 203289
rect 471886 203215 471942 203224
rect 472900 203244 472952 203250
rect 473266 203215 473322 203224
rect 472900 203186 472952 203192
rect 471796 203108 471848 203114
rect 471796 203050 471848 203056
rect 471888 203108 471940 203114
rect 471888 203050 471940 203056
rect 471808 203017 471836 203050
rect 455380 203008 455382 203017
rect 455326 202943 455382 202952
rect 456614 203008 456670 203017
rect 456614 202943 456670 202952
rect 457994 203008 458050 203017
rect 457994 202943 458050 202952
rect 459006 203008 459062 203017
rect 459006 202943 459062 202952
rect 460570 203008 460626 203017
rect 460570 202943 460626 202952
rect 461398 203008 461454 203017
rect 461398 202943 461454 202952
rect 462410 203008 462466 203017
rect 462410 202943 462466 202952
rect 463606 203008 463662 203017
rect 463606 202943 463662 202952
rect 464986 203008 465042 203017
rect 464986 202943 465042 202952
rect 466366 203008 466422 203017
rect 466366 202943 466422 202952
rect 467286 203008 467342 203017
rect 467286 202943 467342 202952
rect 468482 203008 468538 203017
rect 468482 202943 468538 202952
rect 469402 203008 469458 203017
rect 469402 202943 469458 202952
rect 470690 203008 470746 203017
rect 470690 202943 470746 202952
rect 471610 203008 471666 203017
rect 471794 203008 471850 203017
rect 471666 202966 471744 202994
rect 471610 202943 471666 202952
rect 452568 202914 452620 202920
rect 456628 202910 456656 202943
rect 456616 202904 456668 202910
rect 456616 202846 456668 202852
rect 471716 202858 471744 202966
rect 471794 202943 471850 202952
rect 471900 202858 471928 203050
rect 472912 203017 472940 203186
rect 474200 203017 474228 204002
rect 475568 203312 475620 203318
rect 476040 203289 476068 237526
rect 476776 204066 476804 237798
rect 476868 204105 476896 240094
rect 477040 238740 477092 238746
rect 477040 238682 477092 238688
rect 477224 238740 477276 238746
rect 477224 238682 477276 238688
rect 476948 237516 477000 237522
rect 476948 237458 477000 237464
rect 476960 207777 476988 237458
rect 476946 207768 477002 207777
rect 476946 207703 477002 207712
rect 477052 204270 477080 238682
rect 477132 238060 477184 238066
rect 477132 238002 477184 238008
rect 477040 204264 477092 204270
rect 477040 204206 477092 204212
rect 476854 204096 476910 204105
rect 476672 204060 476724 204066
rect 476672 204002 476724 204008
rect 476764 204060 476816 204066
rect 476854 204031 476910 204040
rect 476764 204002 476816 204008
rect 476684 203969 476712 204002
rect 476670 203960 476726 203969
rect 476670 203895 476726 203904
rect 477144 203454 477172 238002
rect 477236 204474 477264 238682
rect 478236 238128 478288 238134
rect 478236 238070 478288 238076
rect 478144 237788 478196 237794
rect 478144 237730 478196 237736
rect 477592 237652 477644 237658
rect 477592 237594 477644 237600
rect 477500 237448 477552 237454
rect 477500 237390 477552 237396
rect 477224 204468 477276 204474
rect 477224 204410 477276 204416
rect 477512 204241 477540 237390
rect 477498 204232 477554 204241
rect 477498 204167 477554 204176
rect 477604 204105 477632 237594
rect 478156 204241 478184 237730
rect 478142 204232 478198 204241
rect 478248 204202 478276 238070
rect 478328 238060 478380 238066
rect 478328 238002 478380 238008
rect 478142 204167 478198 204176
rect 478236 204196 478288 204202
rect 478236 204138 478288 204144
rect 477590 204096 477646 204105
rect 477590 204031 477646 204040
rect 477682 203960 477738 203969
rect 477682 203895 477738 203904
rect 477592 203516 477644 203522
rect 477592 203458 477644 203464
rect 477132 203448 477184 203454
rect 477604 203425 477632 203458
rect 477132 203390 477184 203396
rect 477590 203416 477646 203425
rect 476120 203380 476172 203386
rect 476120 203322 476172 203328
rect 477500 203380 477552 203386
rect 477696 203386 477724 203895
rect 478340 203658 478368 238002
rect 479444 237590 479472 240108
rect 479524 238672 479576 238678
rect 479524 238614 479576 238620
rect 479432 237584 479484 237590
rect 479432 237526 479484 237532
rect 479536 203658 479564 238614
rect 482020 237522 482048 240108
rect 484596 237930 484624 240108
rect 487172 237998 487200 240108
rect 488552 240094 489762 240122
rect 491312 240094 492338 240122
rect 494072 240094 494914 240122
rect 487160 237992 487212 237998
rect 487160 237934 487212 237940
rect 484584 237924 484636 237930
rect 484584 237866 484636 237872
rect 482008 237516 482060 237522
rect 482008 237458 482060 237464
rect 488552 205222 488580 240094
rect 488540 205216 488592 205222
rect 488540 205158 488592 205164
rect 491312 205086 491340 240094
rect 491300 205080 491352 205086
rect 491300 205022 491352 205028
rect 494072 205018 494100 240094
rect 497476 238746 497504 240108
rect 497464 238740 497516 238746
rect 497464 238682 497516 238688
rect 496360 238196 496412 238202
rect 496360 238138 496412 238144
rect 494060 205012 494112 205018
rect 494060 204954 494112 204960
rect 490196 204944 490248 204950
rect 490196 204886 490248 204892
rect 481640 204264 481692 204270
rect 481638 204232 481640 204241
rect 490208 204241 490236 204886
rect 481692 204232 481694 204241
rect 490194 204232 490250 204241
rect 481638 204167 481694 204176
rect 485780 204196 485832 204202
rect 490194 204167 490250 204176
rect 485780 204138 485832 204144
rect 485792 204105 485820 204138
rect 485778 204096 485834 204105
rect 480444 204060 480496 204066
rect 485778 204031 485834 204040
rect 480444 204002 480496 204008
rect 480456 203969 480484 204002
rect 480442 203960 480498 203969
rect 480442 203895 480498 203904
rect 483020 203720 483072 203726
rect 483018 203688 483020 203697
rect 483072 203688 483074 203697
rect 478328 203652 478380 203658
rect 478328 203594 478380 203600
rect 479524 203652 479576 203658
rect 483018 203623 483074 203632
rect 484400 203652 484452 203658
rect 479524 203594 479576 203600
rect 484400 203594 484452 203600
rect 484412 203561 484440 203594
rect 484398 203552 484454 203561
rect 484398 203487 484454 203496
rect 485780 203448 485832 203454
rect 485780 203390 485832 203396
rect 477590 203351 477646 203360
rect 477684 203380 477736 203386
rect 477500 203322 477552 203328
rect 477684 203322 477736 203328
rect 475568 203254 475620 203260
rect 476026 203280 476082 203289
rect 475580 203017 475608 203254
rect 476026 203215 476082 203224
rect 476132 203017 476160 203322
rect 477512 203289 477540 203322
rect 483020 203312 483072 203318
rect 477498 203280 477554 203289
rect 485792 203289 485820 203390
rect 483020 203254 483072 203260
rect 485778 203280 485834 203289
rect 477498 203215 477554 203224
rect 481640 203176 481692 203182
rect 481640 203118 481692 203124
rect 478880 203108 478932 203114
rect 478880 203050 478932 203056
rect 480628 203108 480680 203114
rect 480628 203050 480680 203056
rect 478892 203017 478920 203050
rect 480640 203017 480668 203050
rect 481652 203017 481680 203118
rect 483032 203017 483060 203254
rect 484400 203244 484452 203250
rect 485778 203215 485834 203224
rect 484400 203186 484452 203192
rect 484412 203017 484440 203186
rect 472898 203008 472954 203017
rect 472898 202943 472954 202952
rect 474186 203008 474242 203017
rect 474186 202943 474242 202952
rect 475566 203008 475622 203017
rect 475566 202943 475622 202952
rect 476118 203008 476174 203017
rect 476118 202943 476174 202952
rect 478878 203008 478934 203017
rect 478878 202943 478934 202952
rect 480626 203008 480682 203017
rect 480626 202943 480682 202952
rect 481638 203008 481694 203017
rect 481638 202943 481694 202952
rect 483018 203008 483074 203017
rect 483018 202943 483074 202952
rect 484398 203008 484454 203017
rect 484398 202943 484454 202952
rect 471716 202830 471928 202858
rect 448426 201512 448482 201521
rect 448426 201447 448482 201456
rect 447784 201204 447836 201210
rect 447784 201146 447836 201152
rect 496372 181370 496400 238138
rect 500052 238066 500080 240108
rect 502352 240094 502642 240122
rect 500040 238060 500092 238066
rect 500040 238002 500092 238008
rect 502352 203794 502380 240094
rect 505204 238610 505232 240108
rect 506492 240094 507794 240122
rect 509252 240094 510278 240122
rect 505192 238604 505244 238610
rect 505192 238546 505244 238552
rect 506492 203862 506520 240094
rect 509252 203930 509280 240094
rect 512840 238542 512868 240108
rect 514772 240094 515430 240122
rect 512828 238536 512880 238542
rect 512828 238478 512880 238484
rect 514772 203998 514800 240094
rect 517992 238474 518020 240108
rect 520292 240094 520582 240122
rect 517980 238468 518032 238474
rect 517980 238410 518032 238416
rect 514760 203992 514812 203998
rect 514760 203934 514812 203940
rect 509240 203924 509292 203930
rect 509240 203866 509292 203872
rect 506480 203856 506532 203862
rect 506480 203798 506532 203804
rect 502340 203788 502392 203794
rect 502340 203730 502392 203736
rect 520292 202910 520320 240094
rect 523144 238406 523172 240108
rect 524432 240094 525734 240122
rect 523132 238400 523184 238406
rect 523132 238342 523184 238348
rect 524432 203046 524460 240094
rect 528296 238338 528324 240108
rect 529952 240094 530886 240122
rect 528284 238332 528336 238338
rect 528284 238274 528336 238280
rect 524420 203040 524472 203046
rect 524420 202982 524472 202988
rect 529952 202978 529980 240094
rect 533448 238270 533476 240108
rect 535472 240094 536038 240122
rect 538232 240094 538614 240122
rect 533436 238264 533488 238270
rect 533436 238206 533488 238212
rect 535472 204134 535500 240094
rect 535460 204128 535512 204134
rect 535460 204070 535512 204076
rect 538232 203833 538260 240094
rect 540440 237386 540468 447335
rect 540532 405249 540560 479470
rect 540624 413681 540652 480218
rect 540888 479188 540940 479194
rect 540888 479130 540940 479136
rect 540796 479120 540848 479126
rect 540796 479062 540848 479068
rect 540704 478576 540756 478582
rect 540704 478518 540756 478524
rect 540716 417897 540744 478518
rect 540808 426329 540836 479062
rect 540900 428369 540928 479130
rect 540886 428360 540942 428369
rect 540886 428295 540942 428304
rect 540794 426320 540850 426329
rect 540794 426255 540850 426264
rect 540794 418432 540850 418441
rect 540794 418367 540850 418376
rect 540702 417888 540758 417897
rect 540702 417823 540758 417832
rect 540610 413672 540666 413681
rect 540610 413607 540666 413616
rect 540808 413574 540836 418367
rect 540992 415857 541020 495450
rect 540978 415848 541034 415857
rect 540978 415783 541034 415792
rect 540612 413568 540664 413574
rect 540612 413510 540664 413516
rect 540796 413568 540848 413574
rect 540796 413510 540848 413516
rect 540518 405240 540574 405249
rect 540518 405175 540574 405184
rect 540624 405090 540652 413510
rect 540532 405062 540652 405090
rect 540532 398585 540560 405062
rect 540610 399120 540666 399129
rect 540610 399055 540666 399064
rect 540518 398576 540574 398585
rect 540518 398511 540574 398520
rect 540624 395457 540652 399055
rect 540610 395448 540666 395457
rect 540610 395383 540666 395392
rect 541084 386345 541112 700266
rect 543476 688650 543504 703520
rect 559668 700330 559696 703520
rect 549904 700324 549956 700330
rect 549904 700266 549956 700272
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 543476 688622 543596 688650
rect 541164 681760 541216 681766
rect 541164 681702 541216 681708
rect 541176 392601 541204 681702
rect 543568 676190 543596 688622
rect 543280 676184 543332 676190
rect 543280 676126 543332 676132
rect 543556 676184 543608 676190
rect 543556 676126 543608 676132
rect 543292 669202 543320 676126
rect 547144 673532 547196 673538
rect 547144 673474 547196 673480
rect 543292 669174 543504 669202
rect 541256 667956 541308 667962
rect 541256 667898 541308 667904
rect 541268 396817 541296 667898
rect 543476 659682 543504 669174
rect 543476 659654 543596 659682
rect 543568 647290 543596 659654
rect 543464 647284 543516 647290
rect 543464 647226 543516 647232
rect 543556 647284 543608 647290
rect 543556 647226 543608 647232
rect 543476 640422 543504 647226
rect 543464 640416 543516 640422
rect 543464 640358 543516 640364
rect 543556 640416 543608 640422
rect 543556 640358 543608 640364
rect 543568 630698 543596 640358
rect 543372 630692 543424 630698
rect 543372 630634 543424 630640
rect 543556 630692 543608 630698
rect 543556 630634 543608 630640
rect 543384 630578 543412 630634
rect 543384 630550 543504 630578
rect 543476 621058 543504 630550
rect 545764 626612 545816 626618
rect 545764 626554 545816 626560
rect 543476 621030 543596 621058
rect 543568 611386 543596 621030
rect 543372 611380 543424 611386
rect 543372 611322 543424 611328
rect 543556 611380 543608 611386
rect 543556 611322 543608 611328
rect 543384 611266 543412 611322
rect 543384 611238 543504 611266
rect 541348 610836 541400 610842
rect 541348 610778 541400 610784
rect 541254 396808 541310 396817
rect 541254 396743 541310 396752
rect 541162 392592 541218 392601
rect 541162 392527 541218 392536
rect 541070 386336 541126 386345
rect 541070 386271 541126 386280
rect 541360 342145 541388 610778
rect 541440 610700 541492 610706
rect 541440 610642 541492 610648
rect 541452 348401 541480 610642
rect 541532 610632 541584 610638
rect 541532 610574 541584 610580
rect 541544 354793 541572 610574
rect 541716 610360 541768 610366
rect 541716 610302 541768 610308
rect 541622 449440 541678 449449
rect 541622 449375 541678 449384
rect 541530 354784 541586 354793
rect 541530 354719 541586 354728
rect 541438 348392 541494 348401
rect 541438 348327 541494 348336
rect 541346 342136 541402 342145
rect 541346 342071 541402 342080
rect 541164 280152 541216 280158
rect 541164 280094 541216 280100
rect 541176 279449 541204 280094
rect 541162 279440 541218 279449
rect 541162 279375 541218 279384
rect 540428 237380 540480 237386
rect 540428 237322 540480 237328
rect 538310 222864 538366 222873
rect 538310 222799 538366 222808
rect 538324 205465 538352 222799
rect 539966 216064 540022 216073
rect 539966 215999 540022 216008
rect 538310 205456 538366 205465
rect 538310 205391 538366 205400
rect 538218 203824 538274 203833
rect 538218 203759 538274 203768
rect 539980 203017 540008 215999
rect 541636 208350 541664 449375
rect 541728 403209 541756 610302
rect 543476 601746 543504 611238
rect 543476 601718 543596 601746
rect 543568 592074 543596 601718
rect 543372 592068 543424 592074
rect 543372 592010 543424 592016
rect 543556 592068 543608 592074
rect 543556 592010 543608 592016
rect 543384 591954 543412 592010
rect 543384 591926 543504 591954
rect 543476 582434 543504 591926
rect 543476 582406 543596 582434
rect 543568 572762 543596 582406
rect 544384 579692 544436 579698
rect 544384 579634 544436 579640
rect 543372 572756 543424 572762
rect 543372 572698 543424 572704
rect 543556 572756 543608 572762
rect 543556 572698 543608 572704
rect 543384 572642 543412 572698
rect 543384 572614 543504 572642
rect 543476 563122 543504 572614
rect 543476 563094 543596 563122
rect 543568 553450 543596 563094
rect 543372 553444 543424 553450
rect 543372 553386 543424 553392
rect 543556 553444 543608 553450
rect 543556 553386 543608 553392
rect 543384 553330 543412 553386
rect 543384 553302 543504 553330
rect 543476 543810 543504 553302
rect 543476 543782 543596 543810
rect 543568 534138 543596 543782
rect 543372 534132 543424 534138
rect 543372 534074 543424 534080
rect 543556 534132 543608 534138
rect 543556 534074 543608 534080
rect 543384 534018 543412 534074
rect 543384 533990 543504 534018
rect 543476 524498 543504 533990
rect 543476 524470 543596 524498
rect 543568 514826 543596 524470
rect 543372 514820 543424 514826
rect 543372 514762 543424 514768
rect 543556 514820 543608 514826
rect 543556 514762 543608 514768
rect 543384 514706 543412 514762
rect 543384 514678 543504 514706
rect 543476 512009 543504 514678
rect 543278 512000 543334 512009
rect 543278 511935 543334 511944
rect 543462 512000 543518 512009
rect 543462 511935 543518 511944
rect 543292 502382 543320 511935
rect 543280 502376 543332 502382
rect 543280 502318 543332 502324
rect 543556 502376 543608 502382
rect 543556 502318 543608 502324
rect 543568 492658 543596 502318
rect 543280 492652 543332 492658
rect 543280 492594 543332 492600
rect 543556 492652 543608 492658
rect 543556 492594 543608 492600
rect 543292 483041 543320 492594
rect 543278 483032 543334 483041
rect 543278 482967 543334 482976
rect 543462 483032 543518 483041
rect 543462 482967 543518 482976
rect 543476 480978 543504 482967
rect 543384 480950 543504 480978
rect 541808 479868 541860 479874
rect 541808 479810 541860 479816
rect 541714 403200 541770 403209
rect 541714 403135 541770 403144
rect 541820 337929 541848 479810
rect 541900 479800 541952 479806
rect 541900 479742 541952 479748
rect 541912 361049 541940 479742
rect 541992 479732 542044 479738
rect 541992 479674 542044 479680
rect 542004 367305 542032 479674
rect 542084 479664 542136 479670
rect 542084 479606 542136 479612
rect 542096 373697 542124 479606
rect 542176 479596 542228 479602
rect 542176 479538 542228 479544
rect 542188 379953 542216 479538
rect 542452 478984 542504 478990
rect 542452 478926 542504 478932
rect 542266 466304 542322 466313
rect 542266 466239 542322 466248
rect 542174 379944 542230 379953
rect 542174 379879 542230 379888
rect 542082 373688 542138 373697
rect 542082 373623 542138 373632
rect 541990 367296 542046 367305
rect 541990 367231 542046 367240
rect 541898 361040 541954 361049
rect 541898 360975 541954 360984
rect 541806 337920 541862 337929
rect 541806 337855 541862 337864
rect 542174 241496 542230 241505
rect 542174 241431 542230 241440
rect 542188 234666 542216 241431
rect 542176 234660 542228 234666
rect 542176 234602 542228 234608
rect 541624 208344 541676 208350
rect 541624 208286 541676 208292
rect 539966 203008 540022 203017
rect 529940 202972 529992 202978
rect 539966 202943 540022 202952
rect 529940 202914 529992 202920
rect 520280 202904 520332 202910
rect 520280 202846 520332 202852
rect 500224 202224 500276 202230
rect 500224 202166 500276 202172
rect 499764 202156 499816 202162
rect 499764 202098 499816 202104
rect 499672 201204 499724 201210
rect 499672 201146 499724 201152
rect 496450 181384 496506 181393
rect 496372 181342 496450 181370
rect 496450 181319 496506 181328
rect 417422 180568 417478 180577
rect 417422 180503 417478 180512
rect 418066 171728 418122 171737
rect 418066 171663 418122 171672
rect 393964 115932 394016 115938
rect 393964 115874 394016 115880
rect 380808 115864 380860 115870
rect 380806 115832 380808 115841
rect 391204 115864 391256 115870
rect 380860 115832 380862 115841
rect 391204 115806 391256 115812
rect 380806 115767 380862 115776
rect 380714 114744 380770 114753
rect 380714 114679 380770 114688
rect 300766 111344 300822 111353
rect 300766 111279 300822 111288
rect 416778 111344 416834 111353
rect 416778 111279 416834 111288
rect 300780 110974 300808 111279
rect 416792 110974 416820 111279
rect 300768 110968 300820 110974
rect 300768 110910 300820 110916
rect 416780 110968 416832 110974
rect 416780 110910 416832 110916
rect 303618 109032 303674 109041
rect 303618 108967 303674 108976
rect 307758 109032 307814 109041
rect 307758 108967 307814 108976
rect 303632 108934 303660 108967
rect 307772 108934 307800 108967
rect 418080 108934 418108 171663
rect 499684 115841 499712 201146
rect 499776 118153 499804 202098
rect 499856 201136 499908 201142
rect 499856 201078 499908 201084
rect 499868 118697 499896 201078
rect 499948 201068 500000 201074
rect 499948 201010 500000 201016
rect 499960 120873 499988 201010
rect 500040 201000 500092 201006
rect 500040 200942 500092 200948
rect 500052 122097 500080 200942
rect 500132 200932 500184 200938
rect 500132 200874 500184 200880
rect 500144 123729 500172 200874
rect 500130 123720 500186 123729
rect 500130 123655 500186 123664
rect 500038 122088 500094 122097
rect 500038 122023 500094 122032
rect 499946 120864 500002 120873
rect 499946 120799 500002 120808
rect 499854 118688 499910 118697
rect 499854 118623 499910 118632
rect 499762 118144 499818 118153
rect 499762 118079 499818 118088
rect 499670 115832 499726 115841
rect 499670 115767 499726 115776
rect 500236 115297 500264 202166
rect 500316 201612 500368 201618
rect 500316 201554 500368 201560
rect 500328 183161 500356 201554
rect 539966 193216 540022 193225
rect 539966 193151 540022 193160
rect 539980 183705 540008 193151
rect 539966 183696 540022 183705
rect 539966 183631 540022 183640
rect 500314 183152 500370 183161
rect 500314 183087 500370 183096
rect 540150 167104 540206 167113
rect 540150 167039 540206 167048
rect 540164 164257 540192 167039
rect 540150 164248 540206 164257
rect 540150 164183 540206 164192
rect 539966 162616 540022 162625
rect 539966 162551 540022 162560
rect 539980 153241 540008 162551
rect 539966 153232 540022 153241
rect 539966 153167 540022 153176
rect 539966 147792 540022 147801
rect 539966 147727 540022 147736
rect 539980 144945 540008 147727
rect 539966 144936 540022 144945
rect 539966 144871 540022 144880
rect 539966 120728 540022 120737
rect 539966 120663 540022 120672
rect 539980 115977 540008 120663
rect 539966 115968 540022 115977
rect 539966 115903 540022 115912
rect 500222 115288 500278 115297
rect 500222 115223 500278 115232
rect 424230 109032 424286 109041
rect 424230 108967 424286 108976
rect 427818 109032 427874 109041
rect 542280 109002 542308 466239
rect 542360 451988 542412 451994
rect 542360 451930 542412 451936
rect 542372 445330 542400 451930
rect 542360 445324 542412 445330
rect 542360 445266 542412 445272
rect 542358 445224 542414 445233
rect 542358 445159 542414 445168
rect 542372 223582 542400 445159
rect 542464 441017 542492 478926
rect 543188 478916 543240 478922
rect 543188 478858 543240 478864
rect 542728 478508 542780 478514
rect 542728 478450 542780 478456
rect 542636 478440 542688 478446
rect 542636 478382 542688 478388
rect 542542 451616 542598 451625
rect 542542 451551 542598 451560
rect 542450 441008 542506 441017
rect 542450 440943 542506 440952
rect 542450 438968 542506 438977
rect 542450 438903 542506 438912
rect 542464 243234 542492 438903
rect 542452 243228 542504 243234
rect 542452 243170 542504 243176
rect 542450 243128 542506 243137
rect 542450 243063 542506 243072
rect 542464 242962 542492 243063
rect 542452 242956 542504 242962
rect 542452 242898 542504 242904
rect 542450 241088 542506 241097
rect 542450 241023 542506 241032
rect 542464 240174 542492 241023
rect 542452 240168 542504 240174
rect 542452 240110 542504 240116
rect 542360 223576 542412 223582
rect 542360 223518 542412 223524
rect 542556 200802 542584 451551
rect 542648 430545 542676 478382
rect 542634 430536 542690 430545
rect 542634 430471 542690 430480
rect 542740 424153 542768 478450
rect 542912 478304 542964 478310
rect 542912 478246 542964 478252
rect 542820 478236 542872 478242
rect 542820 478178 542872 478184
rect 542726 424144 542782 424153
rect 542726 424079 542782 424088
rect 542832 401033 542860 478178
rect 542924 407425 542952 478246
rect 543004 478168 543056 478174
rect 543004 478110 543056 478116
rect 543016 409465 543044 478110
rect 543096 478100 543148 478106
rect 543096 478042 543148 478048
rect 543108 420073 543136 478042
rect 543200 422113 543228 478858
rect 543280 478032 543332 478038
rect 543280 477974 543332 477980
rect 543292 436801 543320 477974
rect 543384 476134 543412 480950
rect 543464 479052 543516 479058
rect 543464 478994 543516 479000
rect 543372 476128 543424 476134
rect 543372 476070 543424 476076
rect 543372 460964 543424 460970
rect 543372 460906 543424 460912
rect 543384 451994 543412 460906
rect 543372 451988 543424 451994
rect 543372 451930 543424 451936
rect 543372 441652 543424 441658
rect 543372 441594 543424 441600
rect 543384 437442 543412 441594
rect 543372 437436 543424 437442
rect 543372 437378 543424 437384
rect 543278 436792 543334 436801
rect 543278 436727 543334 436736
rect 543280 436688 543332 436694
rect 543280 436630 543332 436636
rect 543292 427854 543320 436630
rect 543476 434761 543504 478994
rect 543556 478372 543608 478378
rect 543556 478314 543608 478320
rect 543462 434752 543518 434761
rect 543462 434687 543518 434696
rect 543568 432585 543596 478314
rect 543648 476128 543700 476134
rect 543648 476070 543700 476076
rect 543660 460970 543688 476070
rect 543648 460964 543700 460970
rect 543648 460906 543700 460912
rect 543646 453656 543702 453665
rect 543646 453591 543702 453600
rect 543554 432576 543610 432585
rect 543554 432511 543610 432520
rect 543280 427848 543332 427854
rect 543280 427790 543332 427796
rect 543372 427780 543424 427786
rect 543372 427722 543424 427728
rect 543186 422104 543242 422113
rect 543186 422039 543242 422048
rect 543094 420064 543150 420073
rect 543094 419999 543150 420008
rect 543384 418198 543412 427722
rect 543372 418192 543424 418198
rect 543372 418134 543424 418140
rect 543464 418056 543516 418062
rect 543464 417998 543516 418004
rect 543002 409456 543058 409465
rect 543002 409391 543058 409400
rect 542910 407416 542966 407425
rect 542910 407351 542966 407360
rect 543476 404530 543504 417998
rect 543464 404524 543516 404530
rect 543464 404466 543516 404472
rect 543464 404388 543516 404394
rect 543464 404330 543516 404336
rect 542818 401024 542874 401033
rect 542818 400959 542874 400968
rect 543476 399537 543504 404330
rect 543462 399528 543518 399537
rect 543462 399463 543518 399472
rect 543462 389056 543518 389065
rect 543462 388991 543518 389000
rect 543476 386374 543504 388991
rect 543188 386368 543240 386374
rect 543188 386310 543240 386316
rect 543464 386368 543516 386374
rect 543464 386310 543516 386316
rect 543200 376786 543228 386310
rect 543188 376780 543240 376786
rect 543188 376722 543240 376728
rect 543372 376780 543424 376786
rect 543372 376722 543424 376728
rect 543384 376689 543412 376722
rect 543370 376680 543426 376689
rect 543370 376615 543426 376624
rect 543462 369744 543518 369753
rect 543462 369679 543518 369688
rect 543476 367062 543504 369679
rect 543188 367056 543240 367062
rect 543188 366998 543240 367004
rect 543464 367056 543516 367062
rect 543464 366998 543516 367004
rect 543200 357474 543228 366998
rect 543188 357468 543240 357474
rect 543188 357410 543240 357416
rect 543372 357468 543424 357474
rect 543372 357410 543424 357416
rect 543384 357377 543412 357410
rect 543370 357368 543426 357377
rect 543370 357303 543426 357312
rect 543462 350432 543518 350441
rect 543462 350367 543518 350376
rect 543476 339969 543504 350367
rect 543462 339960 543518 339969
rect 543462 339895 543518 339904
rect 542636 336252 542688 336258
rect 542636 336194 542688 336200
rect 542648 335753 542676 336194
rect 542634 335744 542690 335753
rect 542634 335679 542690 335688
rect 542636 333940 542688 333946
rect 542636 333882 542688 333888
rect 542648 333713 542676 333882
rect 542634 333704 542690 333713
rect 542634 333639 542690 333648
rect 542636 332580 542688 332586
rect 542636 332522 542688 332528
rect 542648 331537 542676 332522
rect 542634 331528 542690 331537
rect 542634 331463 542690 331472
rect 542634 329488 542690 329497
rect 542634 329423 542690 329432
rect 542648 328914 542676 329423
rect 542636 328908 542688 328914
rect 542636 328850 542688 328856
rect 542636 328432 542688 328438
rect 542636 328374 542688 328380
rect 542648 327321 542676 328374
rect 542634 327312 542690 327321
rect 542634 327247 542690 327256
rect 542636 325644 542688 325650
rect 542636 325586 542688 325592
rect 542648 325281 542676 325586
rect 542634 325272 542690 325281
rect 542634 325207 542690 325216
rect 542636 324216 542688 324222
rect 542636 324158 542688 324164
rect 542648 323105 542676 324158
rect 542634 323096 542690 323105
rect 542634 323031 542690 323040
rect 542636 321564 542688 321570
rect 542636 321506 542688 321512
rect 542648 321065 542676 321506
rect 542634 321056 542690 321065
rect 542634 320991 542690 321000
rect 542636 320136 542688 320142
rect 542636 320078 542688 320084
rect 542648 318889 542676 320078
rect 542634 318880 542690 318889
rect 542634 318815 542690 318824
rect 542636 316940 542688 316946
rect 542636 316882 542688 316888
rect 542648 316849 542676 316882
rect 542634 316840 542690 316849
rect 542634 316775 542690 316784
rect 542634 314664 542690 314673
rect 542634 314599 542636 314608
rect 542688 314599 542690 314608
rect 542636 314570 542688 314576
rect 542636 313268 542688 313274
rect 542636 313210 542688 313216
rect 542648 312633 542676 313210
rect 542634 312624 542690 312633
rect 542634 312559 542690 312568
rect 542634 310448 542690 310457
rect 542634 310383 542690 310392
rect 542648 310010 542676 310383
rect 542636 310004 542688 310010
rect 542636 309946 542688 309952
rect 542636 309120 542688 309126
rect 542636 309062 542688 309068
rect 542648 308417 542676 309062
rect 542634 308408 542690 308417
rect 542634 308343 542690 308352
rect 542636 306332 542688 306338
rect 542636 306274 542688 306280
rect 542648 306241 542676 306274
rect 542634 306232 542690 306241
rect 542634 306167 542690 306176
rect 542636 304904 542688 304910
rect 542636 304846 542688 304852
rect 542648 304201 542676 304846
rect 542634 304192 542690 304201
rect 542634 304127 542690 304136
rect 542636 302184 542688 302190
rect 542636 302126 542688 302132
rect 542648 302025 542676 302126
rect 542634 302016 542690 302025
rect 542634 301951 542690 301960
rect 542636 300824 542688 300830
rect 542636 300766 542688 300772
rect 542648 299985 542676 300766
rect 542634 299976 542690 299985
rect 542634 299911 542690 299920
rect 542636 298104 542688 298110
rect 542636 298046 542688 298052
rect 542648 297945 542676 298046
rect 542634 297936 542690 297945
rect 542634 297871 542690 297880
rect 542636 296676 542688 296682
rect 542636 296618 542688 296624
rect 542648 295769 542676 296618
rect 542634 295760 542690 295769
rect 542634 295695 542690 295704
rect 542636 293956 542688 293962
rect 542636 293898 542688 293904
rect 542648 293729 542676 293898
rect 542634 293720 542690 293729
rect 542634 293655 542690 293664
rect 542634 291544 542690 291553
rect 542634 291479 542690 291488
rect 542648 291310 542676 291479
rect 542636 291304 542688 291310
rect 542636 291246 542688 291252
rect 542636 289808 542688 289814
rect 542636 289750 542688 289756
rect 542648 289513 542676 289750
rect 542634 289504 542690 289513
rect 542634 289439 542690 289448
rect 542636 288380 542688 288386
rect 542636 288322 542688 288328
rect 542648 287337 542676 288322
rect 542634 287328 542690 287337
rect 542634 287263 542690 287272
rect 542636 285660 542688 285666
rect 542636 285602 542688 285608
rect 542648 285297 542676 285602
rect 542634 285288 542690 285297
rect 542634 285223 542690 285232
rect 542636 284300 542688 284306
rect 542636 284242 542688 284248
rect 542648 283121 542676 284242
rect 542634 283112 542690 283121
rect 542634 283047 542690 283056
rect 542636 281512 542688 281518
rect 542636 281454 542688 281460
rect 542648 281081 542676 281454
rect 542634 281072 542690 281081
rect 542634 281007 542690 281016
rect 543094 276856 543150 276865
rect 543094 276791 543150 276800
rect 542636 275324 542688 275330
rect 542636 275266 542688 275272
rect 542648 274689 542676 275266
rect 542634 274680 542690 274689
rect 542634 274615 542690 274624
rect 543002 272640 543058 272649
rect 543002 272575 543058 272584
rect 542634 257816 542690 257825
rect 542634 257751 542690 257760
rect 542648 256766 542676 257751
rect 542636 256760 542688 256766
rect 542636 256702 542688 256708
rect 542634 255776 542690 255785
rect 542634 255711 542690 255720
rect 542648 255338 542676 255711
rect 542636 255332 542688 255338
rect 542636 255274 542688 255280
rect 542634 253600 542690 253609
rect 542634 253535 542690 253544
rect 542648 252618 542676 253535
rect 542636 252612 542688 252618
rect 542636 252554 542688 252560
rect 543016 252550 543044 272575
rect 543108 264926 543136 276791
rect 543462 270464 543518 270473
rect 543462 270399 543518 270408
rect 543370 266248 543426 266257
rect 543370 266183 543426 266192
rect 543096 264920 543148 264926
rect 543096 264862 543148 264868
rect 543278 262032 543334 262041
rect 543278 261967 543334 261976
rect 543094 259992 543150 260001
rect 543094 259927 543150 259936
rect 543004 252544 543056 252550
rect 543004 252486 543056 252492
rect 543108 251682 543136 259927
rect 543108 251654 543228 251682
rect 543094 251560 543150 251569
rect 543094 251495 543150 251504
rect 542634 249384 542690 249393
rect 542634 249319 542690 249328
rect 542648 248470 542676 249319
rect 542636 248464 542688 248470
rect 542636 248406 542688 248412
rect 542634 247344 542690 247353
rect 542634 247279 542690 247288
rect 542648 247110 542676 247279
rect 542636 247104 542688 247110
rect 542636 247046 542688 247052
rect 542910 245168 542966 245177
rect 542910 245103 542966 245112
rect 542728 243228 542780 243234
rect 542728 243170 542780 243176
rect 542740 241126 542768 243170
rect 542924 241505 542952 245103
rect 542910 241496 542966 241505
rect 542910 241431 542966 241440
rect 542728 241120 542780 241126
rect 542728 241062 542780 241068
rect 542820 234660 542872 234666
rect 542820 234602 542872 234608
rect 542832 231810 542860 234602
rect 542636 231804 542688 231810
rect 542636 231746 542688 231752
rect 542820 231804 542872 231810
rect 542820 231746 542872 231752
rect 542648 222222 542676 231746
rect 542636 222216 542688 222222
rect 542636 222158 542688 222164
rect 542912 222216 542964 222222
rect 542912 222158 542964 222164
rect 542924 215422 542952 222158
rect 542912 215416 542964 215422
rect 542912 215358 542964 215364
rect 542820 215280 542872 215286
rect 542820 215222 542872 215228
rect 542832 212498 542860 215222
rect 542728 212492 542780 212498
rect 542728 212434 542780 212440
rect 542820 212492 542872 212498
rect 542820 212434 542872 212440
rect 542740 202910 542768 212434
rect 542728 202904 542780 202910
rect 542728 202846 542780 202852
rect 542912 202904 542964 202910
rect 542912 202846 542964 202852
rect 542544 200796 542596 200802
rect 542544 200738 542596 200744
rect 542924 196110 542952 202846
rect 542912 196104 542964 196110
rect 542912 196046 542964 196052
rect 542820 195968 542872 195974
rect 542820 195910 542872 195916
rect 542832 186266 542860 195910
rect 542832 186238 542952 186266
rect 542924 178786 542952 186238
rect 542832 178758 542952 178786
rect 542832 173942 542860 178758
rect 542820 173936 542872 173942
rect 543004 173936 543056 173942
rect 542820 173878 542872 173884
rect 543002 173904 543004 173913
rect 543056 173904 543058 173913
rect 543002 173839 543058 173848
rect 543002 164248 543058 164257
rect 543002 164183 543058 164192
rect 543016 162858 543044 164183
rect 542820 162852 542872 162858
rect 542820 162794 542872 162800
rect 543004 162852 543056 162858
rect 543004 162794 543056 162800
rect 542832 153270 542860 162794
rect 542820 153264 542872 153270
rect 542820 153206 542872 153212
rect 543004 153264 543056 153270
rect 543004 153206 543056 153212
rect 543016 143546 543044 153206
rect 543004 143540 543056 143546
rect 543004 143482 543056 143488
rect 543004 133952 543056 133958
rect 543004 133894 543056 133900
rect 543016 124166 543044 133894
rect 543004 124160 543056 124166
rect 543004 124102 543056 124108
rect 543108 109138 543136 251495
rect 543200 158710 543228 251654
rect 543292 182170 543320 261967
rect 543384 205630 543412 266183
rect 543476 218006 543504 270399
rect 543554 268424 543610 268433
rect 543554 268359 543610 268368
rect 543568 229090 543596 268359
rect 543556 229084 543608 229090
rect 543556 229026 543608 229032
rect 543464 218000 543516 218006
rect 543464 217942 543516 217948
rect 543372 205624 543424 205630
rect 543372 205566 543424 205572
rect 543660 200870 543688 453591
rect 543740 445324 543792 445330
rect 543740 445266 543792 445272
rect 543752 441658 543780 445266
rect 543740 441652 543792 441658
rect 543740 441594 543792 441600
rect 544396 316946 544424 579634
rect 544476 532772 544528 532778
rect 544476 532714 544528 532720
rect 544384 316940 544436 316946
rect 544384 316882 544436 316888
rect 544488 310010 544516 532714
rect 544568 485852 544620 485858
rect 544568 485794 544620 485800
rect 544476 310004 544528 310010
rect 544476 309946 544528 309952
rect 544580 304910 544608 485794
rect 544660 392012 544712 392018
rect 544660 391954 544712 391960
rect 544568 304904 544620 304910
rect 544568 304846 544620 304852
rect 544672 291310 544700 391954
rect 545776 324222 545804 626554
rect 547156 328914 547184 673474
rect 549916 336258 549944 700266
rect 580170 698048 580226 698057
rect 580170 697983 580226 697992
rect 580184 696998 580212 697983
rect 563704 696992 563756 696998
rect 563704 696934 563756 696940
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 554044 685908 554096 685914
rect 554044 685850 554096 685856
rect 549996 404388 550048 404394
rect 549996 404330 550048 404336
rect 549904 336252 549956 336258
rect 549904 336194 549956 336200
rect 547144 328908 547196 328914
rect 547144 328850 547196 328856
rect 545764 324216 545816 324222
rect 545764 324158 545816 324164
rect 550008 296682 550036 404330
rect 554056 333946 554084 685850
rect 560944 650072 560996 650078
rect 560944 650014 560996 650020
rect 558184 603152 558236 603158
rect 558184 603094 558236 603100
rect 556804 556232 556856 556238
rect 556804 556174 556856 556180
rect 555424 509312 555476 509318
rect 555424 509254 555476 509260
rect 554136 438932 554188 438938
rect 554136 438874 554188 438880
rect 554044 333940 554096 333946
rect 554044 333882 554096 333888
rect 554148 298110 554176 438874
rect 555436 306338 555464 509254
rect 556816 313274 556844 556174
rect 558196 320142 558224 603094
rect 560956 325650 560984 650014
rect 563716 332586 563744 696934
rect 580170 686352 580226 686361
rect 580170 686287 580226 686296
rect 580184 685914 580212 686287
rect 580172 685908 580224 685914
rect 580172 685850 580224 685856
rect 580170 674656 580226 674665
rect 580170 674591 580226 674600
rect 580184 673538 580212 674591
rect 580172 673532 580224 673538
rect 580172 673474 580224 673480
rect 580170 651128 580226 651137
rect 580170 651063 580226 651072
rect 580184 650078 580212 651063
rect 580172 650072 580224 650078
rect 580172 650014 580224 650020
rect 580170 639432 580226 639441
rect 580170 639367 580226 639376
rect 580184 638994 580212 639367
rect 565084 638988 565136 638994
rect 565084 638930 565136 638936
rect 580172 638988 580224 638994
rect 580172 638930 580224 638936
rect 563796 451308 563848 451314
rect 563796 451250 563848 451256
rect 563704 332580 563756 332586
rect 563704 332522 563756 332528
rect 560944 325644 560996 325650
rect 560944 325586 560996 325592
rect 558184 320136 558236 320142
rect 558184 320078 558236 320084
rect 556804 313268 556856 313274
rect 556804 313210 556856 313216
rect 555424 306332 555476 306338
rect 555424 306274 555476 306280
rect 563808 302190 563836 451250
rect 565096 328438 565124 638930
rect 580170 627736 580226 627745
rect 580170 627671 580226 627680
rect 580184 626618 580212 627671
rect 580172 626612 580224 626618
rect 580172 626554 580224 626560
rect 580170 604208 580226 604217
rect 580170 604143 580226 604152
rect 580184 603158 580212 604143
rect 580172 603152 580224 603158
rect 580172 603094 580224 603100
rect 580170 592512 580226 592521
rect 580170 592447 580226 592456
rect 580184 592074 580212 592447
rect 574744 592068 574796 592074
rect 574744 592010 574796 592016
rect 580172 592068 580224 592074
rect 580172 592010 580224 592016
rect 573364 545148 573416 545154
rect 573364 545090 573416 545096
rect 571984 498228 572036 498234
rect 571984 498170 572036 498176
rect 567844 462392 567896 462398
rect 567844 462334 567896 462340
rect 565176 415472 565228 415478
rect 565176 415414 565228 415420
rect 565084 328432 565136 328438
rect 565084 328374 565136 328380
rect 563796 302184 563848 302190
rect 563796 302126 563848 302132
rect 554136 298104 554188 298110
rect 554136 298046 554188 298052
rect 549996 296676 550048 296682
rect 549996 296618 550048 296624
rect 565188 293962 565216 415414
rect 567856 300830 567884 462334
rect 571996 309126 572024 498170
rect 573376 314634 573404 545090
rect 574756 321570 574784 592010
rect 580170 580816 580226 580825
rect 580170 580751 580226 580760
rect 580184 579698 580212 580751
rect 580172 579692 580224 579698
rect 580172 579634 580224 579640
rect 580170 557288 580226 557297
rect 580170 557223 580226 557232
rect 580184 556238 580212 557223
rect 580172 556232 580224 556238
rect 580172 556174 580224 556180
rect 580170 545592 580226 545601
rect 580170 545527 580226 545536
rect 580184 545154 580212 545527
rect 580172 545148 580224 545154
rect 580172 545090 580224 545096
rect 580170 533896 580226 533905
rect 580170 533831 580226 533840
rect 580184 532778 580212 533831
rect 580172 532772 580224 532778
rect 580172 532714 580224 532720
rect 580170 510368 580226 510377
rect 580170 510303 580226 510312
rect 580184 509318 580212 510303
rect 580172 509312 580224 509318
rect 580172 509254 580224 509260
rect 580170 498672 580226 498681
rect 580170 498607 580226 498616
rect 580184 498234 580212 498607
rect 580172 498228 580224 498234
rect 580172 498170 580224 498176
rect 580170 486840 580226 486849
rect 580170 486775 580226 486784
rect 580184 485858 580212 486775
rect 580172 485852 580224 485858
rect 580172 485794 580224 485800
rect 580170 463448 580226 463457
rect 580170 463383 580226 463392
rect 580184 462398 580212 463383
rect 580172 462392 580224 462398
rect 580172 462334 580224 462340
rect 580170 451752 580226 451761
rect 580170 451687 580226 451696
rect 580184 451314 580212 451687
rect 580172 451308 580224 451314
rect 580172 451250 580224 451256
rect 580170 439920 580226 439929
rect 580170 439855 580226 439864
rect 580184 438938 580212 439855
rect 580172 438932 580224 438938
rect 580172 438874 580224 438880
rect 580170 416528 580226 416537
rect 580170 416463 580226 416472
rect 580184 415478 580212 416463
rect 580172 415472 580224 415478
rect 580172 415414 580224 415420
rect 580170 404832 580226 404841
rect 580170 404767 580226 404776
rect 580184 404394 580212 404767
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 580170 393000 580226 393009
rect 580170 392935 580226 392944
rect 580184 392018 580212 392935
rect 580172 392012 580224 392018
rect 580172 391954 580224 391960
rect 580262 369608 580318 369617
rect 580262 369543 580318 369552
rect 574744 321564 574796 321570
rect 574744 321506 574796 321512
rect 573364 314628 573416 314634
rect 573364 314570 573416 314576
rect 571984 309120 572036 309126
rect 571984 309062 572036 309068
rect 567844 300824 567896 300830
rect 567844 300766 567896 300772
rect 565176 293956 565228 293962
rect 565176 293898 565228 293904
rect 544660 291304 544712 291310
rect 544660 291246 544712 291252
rect 580276 288386 580304 369543
rect 580354 357912 580410 357921
rect 580354 357847 580410 357856
rect 580368 289814 580396 357847
rect 580446 346080 580502 346089
rect 580446 346015 580502 346024
rect 580356 289808 580408 289814
rect 580356 289750 580408 289756
rect 580264 288380 580316 288386
rect 580264 288322 580316 288328
rect 580460 285666 580488 346015
rect 580538 322688 580594 322697
rect 580538 322623 580594 322632
rect 580448 285660 580500 285666
rect 580448 285602 580500 285608
rect 580552 281518 580580 322623
rect 580630 310856 580686 310865
rect 580630 310791 580686 310800
rect 580644 284306 580672 310791
rect 580722 299160 580778 299169
rect 580722 299095 580778 299104
rect 580632 284300 580684 284306
rect 580632 284242 580684 284248
rect 580540 281512 580592 281518
rect 580540 281454 580592 281460
rect 580736 280158 580764 299095
rect 580724 280152 580776 280158
rect 580724 280094 580776 280100
rect 580170 275768 580226 275777
rect 580170 275703 580226 275712
rect 580184 275330 580212 275703
rect 580172 275324 580224 275330
rect 580172 275266 580224 275272
rect 580172 264920 580224 264926
rect 580172 264862 580224 264868
rect 544382 264208 544438 264217
rect 544382 264143 544438 264152
rect 543648 200864 543700 200870
rect 543648 200806 543700 200812
rect 543280 182164 543332 182170
rect 543280 182106 543332 182112
rect 544396 171086 544424 264143
rect 580184 263945 580212 264862
rect 580170 263936 580226 263945
rect 580170 263871 580226 263880
rect 558184 256760 558236 256766
rect 558184 256702 558236 256708
rect 556804 255332 556856 255338
rect 556804 255274 556856 255280
rect 549904 252612 549956 252618
rect 549904 252554 549956 252560
rect 547144 247104 547196 247110
rect 547144 247046 547196 247052
rect 545764 240168 545816 240174
rect 545764 240110 545816 240116
rect 544384 171080 544436 171086
rect 544384 171022 544436 171028
rect 543188 158704 543240 158710
rect 543188 158646 543240 158652
rect 543188 143540 543240 143546
rect 543188 143482 543240 143488
rect 543200 133958 543228 143482
rect 543188 133952 543240 133958
rect 543188 133894 543240 133900
rect 543372 124160 543424 124166
rect 543372 124102 543424 124108
rect 543096 109132 543148 109138
rect 543096 109074 543148 109080
rect 427818 108967 427874 108976
rect 542268 108996 542320 109002
rect 424244 108934 424272 108967
rect 427832 108934 427860 108967
rect 542268 108938 542320 108944
rect 543096 108996 543148 109002
rect 543096 108938 543148 108944
rect 297916 108928 297968 108934
rect 297916 108870 297968 108876
rect 303620 108928 303672 108934
rect 303620 108870 303672 108876
rect 305644 108928 305696 108934
rect 305644 108870 305696 108876
rect 307760 108928 307812 108934
rect 307760 108870 307812 108876
rect 418068 108928 418120 108934
rect 418068 108870 418120 108876
rect 424232 108928 424284 108934
rect 424232 108870 424284 108876
rect 427820 108928 427872 108934
rect 427820 108870 427872 108876
rect 257436 3528 257488 3534
rect 257436 3470 257488 3476
rect 257344 3460 257396 3466
rect 257344 3402 257396 3408
rect 305656 2854 305684 108870
rect 543016 99414 543044 99445
rect 543004 99408 543056 99414
rect 542924 99356 543004 99362
rect 542924 99350 543056 99356
rect 542924 99334 543044 99350
rect 542924 96626 542952 99334
rect 542820 96620 542872 96626
rect 542820 96562 542872 96568
rect 542912 96620 542964 96626
rect 542912 96562 542964 96568
rect 542832 89758 542860 96562
rect 542820 89752 542872 89758
rect 542820 89694 542872 89700
rect 542912 89684 542964 89690
rect 542912 89626 542964 89632
rect 542924 86986 542952 89626
rect 542832 86970 542952 86986
rect 542820 86964 542952 86970
rect 542872 86958 542952 86964
rect 542820 86906 542872 86912
rect 542910 77208 542966 77217
rect 543108 77178 543136 108938
rect 543384 106321 543412 124102
rect 543186 106312 543242 106321
rect 543186 106247 543242 106256
rect 543370 106312 543426 106321
rect 543370 106247 543426 106256
rect 543200 99414 543228 106247
rect 543188 99408 543240 99414
rect 543188 99350 543240 99356
rect 543280 86964 543332 86970
rect 543280 86906 543332 86912
rect 543292 77330 543320 86906
rect 543200 77302 543320 77330
rect 543200 77217 543228 77302
rect 543186 77208 543242 77217
rect 542910 77143 542966 77152
rect 543096 77172 543148 77178
rect 542924 67658 542952 77143
rect 543186 77143 543242 77152
rect 543096 77114 543148 77120
rect 542912 67652 542964 67658
rect 542912 67594 542964 67600
rect 543096 67652 543148 67658
rect 543096 67594 543148 67600
rect 543108 60790 543136 67594
rect 543096 60784 543148 60790
rect 543096 60726 543148 60732
rect 542820 60716 542872 60722
rect 542820 60658 542872 60664
rect 542832 51066 542860 60658
rect 542820 51060 542872 51066
rect 542820 51002 542872 51008
rect 543004 51060 543056 51066
rect 543004 51002 543056 51008
rect 543016 48278 543044 51002
rect 543004 48272 543056 48278
rect 543004 48214 543056 48220
rect 543280 48272 543332 48278
rect 543280 48214 543332 48220
rect 543292 38690 543320 48214
rect 543096 38684 543148 38690
rect 543096 38626 543148 38632
rect 543280 38684 543332 38690
rect 543280 38626 543332 38632
rect 543108 30326 543136 38626
rect 543096 30320 543148 30326
rect 543096 30262 543148 30268
rect 545776 17950 545804 240110
rect 547156 64870 547184 247046
rect 549916 111790 549944 252554
rect 555424 248464 555476 248470
rect 555424 248406 555476 248412
rect 554044 242956 554096 242962
rect 554044 242898 554096 242904
rect 549904 111784 549956 111790
rect 549904 111726 549956 111732
rect 547144 64864 547196 64870
rect 547144 64806 547196 64812
rect 554056 41410 554084 242898
rect 555436 88330 555464 248406
rect 556816 135250 556844 255274
rect 556804 135244 556856 135250
rect 556804 135186 556856 135192
rect 558196 124166 558224 256702
rect 579804 252544 579856 252550
rect 579804 252486 579856 252492
rect 579816 252249 579844 252486
rect 579802 252240 579858 252249
rect 579802 252175 579858 252184
rect 580172 229084 580224 229090
rect 580172 229026 580224 229032
rect 580184 228857 580212 229026
rect 580170 228848 580226 228857
rect 580170 228783 580226 228792
rect 580172 218000 580224 218006
rect 580172 217942 580224 217948
rect 580184 217025 580212 217942
rect 580170 217016 580226 217025
rect 580170 216951 580226 216960
rect 579804 205624 579856 205630
rect 579804 205566 579856 205572
rect 579816 205329 579844 205566
rect 579802 205320 579858 205329
rect 579802 205255 579858 205264
rect 580172 182164 580224 182170
rect 580172 182106 580224 182112
rect 580184 181937 580212 182106
rect 580170 181928 580226 181937
rect 580170 181863 580226 181872
rect 580172 171080 580224 171086
rect 580172 171022 580224 171028
rect 580184 170105 580212 171022
rect 580170 170096 580226 170105
rect 580170 170031 580226 170040
rect 579804 158704 579856 158710
rect 579804 158646 579856 158652
rect 579816 158409 579844 158646
rect 579802 158400 579858 158409
rect 579802 158335 579858 158344
rect 580172 135244 580224 135250
rect 580172 135186 580224 135192
rect 580184 134881 580212 135186
rect 580170 134872 580226 134881
rect 580170 134807 580226 134816
rect 558184 124160 558236 124166
rect 558184 124102 558236 124108
rect 580172 124160 580224 124166
rect 580172 124102 580224 124108
rect 580184 123185 580212 124102
rect 580170 123176 580226 123185
rect 580170 123111 580226 123120
rect 579804 111784 579856 111790
rect 579804 111726 579856 111732
rect 579816 111489 579844 111726
rect 579802 111480 579858 111489
rect 579802 111415 579858 111424
rect 555424 88324 555476 88330
rect 555424 88266 555476 88272
rect 580172 88324 580224 88330
rect 580172 88266 580224 88272
rect 580184 87961 580212 88266
rect 580170 87952 580226 87961
rect 580170 87887 580226 87896
rect 580172 77240 580224 77246
rect 580172 77182 580224 77188
rect 580184 76265 580212 77182
rect 580170 76256 580226 76265
rect 580170 76191 580226 76200
rect 579804 64864 579856 64870
rect 579804 64806 579856 64812
rect 579816 64569 579844 64806
rect 579802 64560 579858 64569
rect 579802 64495 579858 64504
rect 554044 41404 554096 41410
rect 554044 41346 554096 41352
rect 580172 41404 580224 41410
rect 580172 41346 580224 41352
rect 580184 41041 580212 41346
rect 580170 41032 580226 41041
rect 580170 40967 580226 40976
rect 580172 30320 580224 30326
rect 580172 30262 580224 30268
rect 580184 29345 580212 30262
rect 580170 29336 580226 29345
rect 580170 29271 580226 29280
rect 545764 17944 545816 17950
rect 545764 17886 545816 17892
rect 579804 17944 579856 17950
rect 579804 17886 579856 17892
rect 579816 17649 579844 17886
rect 579802 17640 579858 17649
rect 579802 17575 579858 17584
rect 142068 2848 142120 2854
rect 142068 2790 142120 2796
rect 145656 2848 145708 2854
rect 145656 2790 145708 2796
rect 149244 2848 149296 2854
rect 149244 2790 149296 2796
rect 152740 2848 152792 2854
rect 152740 2790 152792 2796
rect 156328 2848 156380 2854
rect 156328 2790 156380 2796
rect 159916 2848 159968 2854
rect 159916 2790 159968 2796
rect 163504 2848 163556 2854
rect 163504 2790 163556 2796
rect 167092 2848 167144 2854
rect 167092 2790 167144 2796
rect 170588 2848 170640 2854
rect 170588 2790 170640 2796
rect 174176 2848 174228 2854
rect 174176 2790 174228 2796
rect 177764 2848 177816 2854
rect 177764 2790 177816 2796
rect 181352 2848 181404 2854
rect 181352 2790 181404 2796
rect 184848 2848 184900 2854
rect 184848 2790 184900 2796
rect 188436 2848 188488 2854
rect 188436 2790 188488 2796
rect 192024 2848 192076 2854
rect 192024 2790 192076 2796
rect 195612 2848 195664 2854
rect 195612 2790 195664 2796
rect 199200 2848 199252 2854
rect 199200 2790 199252 2796
rect 202696 2848 202748 2854
rect 202696 2790 202748 2796
rect 206284 2848 206336 2854
rect 206284 2790 206336 2796
rect 209872 2848 209924 2854
rect 209872 2790 209924 2796
rect 213460 2848 213512 2854
rect 213460 2790 213512 2796
rect 217048 2848 217100 2854
rect 217048 2790 217100 2796
rect 220544 2848 220596 2854
rect 220544 2790 220596 2796
rect 224132 2848 224184 2854
rect 224132 2790 224184 2796
rect 227720 2848 227772 2854
rect 227720 2790 227772 2796
rect 231308 2848 231360 2854
rect 231308 2790 231360 2796
rect 234804 2848 234856 2854
rect 234804 2790 234856 2796
rect 238392 2848 238444 2854
rect 238392 2790 238444 2796
rect 241980 2848 242032 2854
rect 241980 2790 242032 2796
rect 245568 2848 245620 2854
rect 245568 2790 245620 2796
rect 249156 2848 249208 2854
rect 249156 2790 249208 2796
rect 252652 2848 252704 2854
rect 252652 2790 252704 2796
rect 256240 2848 256292 2854
rect 256240 2790 256292 2796
rect 259828 2848 259880 2854
rect 259828 2790 259880 2796
rect 263416 2848 263468 2854
rect 263416 2790 263468 2796
rect 267004 2848 267056 2854
rect 267004 2790 267056 2796
rect 270500 2848 270552 2854
rect 270500 2790 270552 2796
rect 274088 2848 274140 2854
rect 274088 2790 274140 2796
rect 277676 2848 277728 2854
rect 277676 2790 277728 2796
rect 281264 2848 281316 2854
rect 281264 2790 281316 2796
rect 284760 2848 284812 2854
rect 284760 2790 284812 2796
rect 288348 2848 288400 2854
rect 288348 2790 288400 2796
rect 291936 2848 291988 2854
rect 291936 2790 291988 2796
rect 295524 2848 295576 2854
rect 295524 2790 295576 2796
rect 299112 2848 299164 2854
rect 299112 2790 299164 2796
rect 302608 2848 302660 2854
rect 302608 2790 302660 2796
rect 305644 2848 305696 2854
rect 305644 2790 305696 2796
rect 306196 2848 306248 2854
rect 306196 2790 306248 2796
rect 309784 2848 309836 2854
rect 309784 2790 309836 2796
rect 313372 2848 313424 2854
rect 313372 2790 313424 2796
rect 316960 2848 317012 2854
rect 316960 2790 317012 2796
rect 320456 2848 320508 2854
rect 320456 2790 320508 2796
rect 324044 2848 324096 2854
rect 324044 2790 324096 2796
rect 327632 2848 327684 2854
rect 327632 2790 327684 2796
rect 331220 2848 331272 2854
rect 331220 2790 331272 2796
rect 334716 2848 334768 2854
rect 334716 2790 334768 2796
rect 338304 2848 338356 2854
rect 338304 2790 338356 2796
rect 341892 2848 341944 2854
rect 341892 2790 341944 2796
rect 345480 2848 345532 2854
rect 345480 2790 345532 2796
rect 349068 2848 349120 2854
rect 349068 2790 349120 2796
rect 352564 2848 352616 2854
rect 352564 2790 352616 2796
rect 356152 2848 356204 2854
rect 356152 2790 356204 2796
rect 359740 2848 359792 2854
rect 359740 2790 359792 2796
rect 363328 2848 363380 2854
rect 363328 2790 363380 2796
rect 366916 2848 366968 2854
rect 366916 2790 366968 2796
rect 370412 2848 370464 2854
rect 370412 2790 370464 2796
rect 374000 2848 374052 2854
rect 374000 2790 374052 2796
rect 377588 2848 377640 2854
rect 377588 2790 377640 2796
rect 381176 2848 381228 2854
rect 381176 2790 381228 2796
rect 384672 2848 384724 2854
rect 384672 2790 384724 2796
rect 388260 2848 388312 2854
rect 388260 2790 388312 2796
rect 391848 2848 391900 2854
rect 391848 2790 391900 2796
rect 395436 2848 395488 2854
rect 395436 2790 395488 2796
rect 399024 2848 399076 2854
rect 399024 2790 399076 2796
rect 402520 2848 402572 2854
rect 402520 2790 402572 2796
rect 406108 2848 406160 2854
rect 406108 2790 406160 2796
rect 409696 2848 409748 2854
rect 409696 2790 409748 2796
rect 413284 2848 413336 2854
rect 413284 2790 413336 2796
rect 416872 2848 416924 2854
rect 416872 2790 416924 2796
rect 420368 2848 420420 2854
rect 420368 2790 420420 2796
rect 423956 2848 424008 2854
rect 423956 2790 424008 2796
rect 427544 2848 427596 2854
rect 427544 2790 427596 2796
rect 431132 2848 431184 2854
rect 431132 2790 431184 2796
rect 434628 2848 434680 2854
rect 434628 2790 434680 2796
rect 438216 2848 438268 2854
rect 438216 2790 438268 2796
rect 441804 2848 441856 2854
rect 441804 2790 441856 2796
rect 445392 2848 445444 2854
rect 445392 2790 445444 2796
rect 448980 2848 449032 2854
rect 448980 2790 449032 2796
rect 452476 2848 452528 2854
rect 452476 2790 452528 2796
rect 456064 2848 456116 2854
rect 456064 2790 456116 2796
rect 459652 2848 459704 2854
rect 459652 2790 459704 2796
rect 463240 2848 463292 2854
rect 463240 2790 463292 2796
rect 466828 2848 466880 2854
rect 466828 2790 466880 2796
rect 470324 2848 470376 2854
rect 470324 2790 470376 2796
rect 473912 2848 473964 2854
rect 473912 2790 473964 2796
rect 477500 2848 477552 2854
rect 477500 2790 477552 2796
rect 481088 2848 481140 2854
rect 481088 2790 481140 2796
rect 484584 2848 484636 2854
rect 484584 2790 484636 2796
rect 488172 2848 488224 2854
rect 488172 2790 488224 2796
rect 491760 2848 491812 2854
rect 491760 2790 491812 2796
rect 495348 2848 495400 2854
rect 495348 2790 495400 2796
rect 498936 2848 498988 2854
rect 498936 2790 498988 2796
rect 502432 2848 502484 2854
rect 502432 2790 502484 2796
rect 506020 2848 506072 2854
rect 506020 2790 506072 2796
rect 509608 2848 509660 2854
rect 509608 2790 509660 2796
rect 513196 2848 513248 2854
rect 513196 2790 513248 2796
rect 516784 2848 516836 2854
rect 516784 2790 516836 2796
rect 520280 2848 520332 2854
rect 520280 2790 520332 2796
rect 523868 2848 523920 2854
rect 523868 2790 523920 2796
rect 527456 2848 527508 2854
rect 527456 2790 527508 2796
rect 531044 2848 531096 2854
rect 531044 2790 531096 2796
rect 534540 2848 534592 2854
rect 534540 2790 534592 2796
rect 538128 2848 538180 2854
rect 538128 2790 538180 2796
rect 541716 2848 541768 2854
rect 541716 2790 541768 2796
rect 545304 2848 545356 2854
rect 545304 2790 545356 2796
rect 548892 2848 548944 2854
rect 548892 2790 548944 2796
rect 552388 2848 552440 2854
rect 552388 2790 552440 2796
rect 555976 2848 556028 2854
rect 555976 2790 556028 2796
rect 559564 2848 559616 2854
rect 559564 2790 559616 2796
rect 563152 2848 563204 2854
rect 563152 2790 563204 2796
rect 566740 2848 566792 2854
rect 566740 2790 566792 2796
rect 570236 2848 570288 2854
rect 570236 2790 570288 2796
rect 573824 2848 573876 2854
rect 573824 2790 573876 2796
rect 577412 2848 577464 2854
rect 577412 2790 577464 2796
rect 581000 2848 581052 2854
rect 581000 2790 581052 2796
rect 134904 598 135208 626
rect 142080 610 142108 2790
rect 138480 604 138532 610
rect 134904 480 134932 598
rect 138480 546 138532 552
rect 142068 604 142120 610
rect 142068 546 142120 552
rect 138492 480 138520 546
rect 142080 480 142108 546
rect 145668 480 145696 2790
rect 149256 480 149284 2790
rect 152752 480 152780 2790
rect 156340 480 156368 2790
rect 159928 480 159956 2790
rect 163516 480 163544 2790
rect 167104 480 167132 2790
rect 170600 480 170628 2790
rect 174188 480 174216 2790
rect 177776 480 177804 2790
rect 181364 480 181392 2790
rect 184860 480 184888 2790
rect 188448 480 188476 2790
rect 192036 480 192064 2790
rect 195624 480 195652 2790
rect 199212 480 199240 2790
rect 202708 480 202736 2790
rect 206296 480 206324 2790
rect 209884 480 209912 2790
rect 213472 480 213500 2790
rect 217060 480 217088 2790
rect 220556 480 220584 2790
rect 224144 480 224172 2790
rect 227732 480 227760 2790
rect 231320 480 231348 2790
rect 234816 480 234844 2790
rect 238404 480 238432 2790
rect 241992 480 242020 2790
rect 245580 480 245608 2790
rect 249168 480 249196 2790
rect 252664 480 252692 2790
rect 256252 480 256280 2790
rect 259840 480 259868 2790
rect 263428 480 263456 2790
rect 267016 480 267044 2790
rect 270512 480 270540 2790
rect 274100 480 274128 2790
rect 277688 480 277716 2790
rect 281276 480 281304 2790
rect 284772 480 284800 2790
rect 288360 480 288388 2790
rect 291948 480 291976 2790
rect 295536 480 295564 2790
rect 299124 480 299152 2790
rect 302620 480 302648 2790
rect 306208 480 306236 2790
rect 309796 480 309824 2790
rect 313384 480 313412 2790
rect 316972 480 317000 2790
rect 320468 480 320496 2790
rect 324056 480 324084 2790
rect 327644 480 327672 2790
rect 331232 480 331260 2790
rect 334728 480 334756 2790
rect 338316 480 338344 2790
rect 341904 480 341932 2790
rect 345492 480 345520 2790
rect 349080 480 349108 2790
rect 352576 480 352604 2790
rect 356164 480 356192 2790
rect 359752 480 359780 2790
rect 363340 480 363368 2790
rect 366928 480 366956 2790
rect 370424 480 370452 2790
rect 374012 480 374040 2790
rect 377600 480 377628 2790
rect 381188 480 381216 2790
rect 384684 480 384712 2790
rect 388272 480 388300 2790
rect 391860 480 391888 2790
rect 395448 480 395476 2790
rect 399036 480 399064 2790
rect 402532 480 402560 2790
rect 406120 480 406148 2790
rect 409708 480 409736 2790
rect 413296 480 413324 2790
rect 416884 480 416912 2790
rect 420380 480 420408 2790
rect 423968 480 423996 2790
rect 427556 480 427584 2790
rect 431144 480 431172 2790
rect 434640 480 434668 2790
rect 438228 480 438256 2790
rect 441816 480 441844 2790
rect 445404 480 445432 2790
rect 448992 480 449020 2790
rect 452488 480 452516 2790
rect 456076 480 456104 2790
rect 459664 480 459692 2790
rect 463252 480 463280 2790
rect 466840 480 466868 2790
rect 470336 480 470364 2790
rect 473924 480 473952 2790
rect 477512 480 477540 2790
rect 481100 480 481128 2790
rect 484596 480 484624 2790
rect 488184 480 488212 2790
rect 491772 480 491800 2790
rect 495360 480 495388 2790
rect 498948 480 498976 2790
rect 502444 480 502472 2790
rect 506032 480 506060 2790
rect 509620 480 509648 2790
rect 513208 480 513236 2790
rect 516796 480 516824 2790
rect 520292 480 520320 2790
rect 523880 480 523908 2790
rect 527468 480 527496 2790
rect 531056 480 531084 2790
rect 534552 480 534580 2790
rect 538140 480 538168 2790
rect 541728 480 541756 2790
rect 545316 480 545344 2790
rect 548904 480 548932 2790
rect 552400 480 552428 2790
rect 555988 480 556016 2790
rect 559576 480 559604 2790
rect 563164 480 563192 2790
rect 566752 480 566780 2790
rect 570248 480 570276 2790
rect 573836 480 573864 2790
rect 577424 480 577452 2790
rect 581012 480 581040 2790
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 13606 -960 13718 480
rect 14802 -960 14914 480
rect 15998 -960 16110 480
rect 17194 -960 17306 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 27866 -960 27978 480
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44518 -960 44630 480
rect 45714 -960 45826 480
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49302 -960 49414 480
rect 50498 -960 50610 480
rect 51602 -960 51714 480
rect 52798 -960 52910 480
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 56386 -960 56498 480
rect 57582 -960 57694 480
rect 58778 -960 58890 480
rect 59974 -960 60086 480
rect 61170 -960 61282 480
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64758 -960 64870 480
rect 65954 -960 66066 480
rect 67150 -960 67262 480
rect 68254 -960 68366 480
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 73038 -960 73150 480
rect 74234 -960 74346 480
rect 75430 -960 75542 480
rect 76626 -960 76738 480
rect 77822 -960 77934 480
rect 79018 -960 79130 480
rect 80214 -960 80326 480
rect 81410 -960 81522 480
rect 82606 -960 82718 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 88494 -960 88606 480
rect 89690 -960 89802 480
rect 90886 -960 90998 480
rect 92082 -960 92194 480
rect 93278 -960 93390 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 107538 -960 107650 480
rect 108734 -960 108846 480
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 151514 -960 151626 480
rect 152710 -960 152822 480
rect 153906 -960 154018 480
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157494 -960 157606 480
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 162278 -960 162390 480
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 189602 -960 189714 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197974 -960 198086 480
rect 199170 -960 199282 480
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246734 -960 246846 480
rect 247930 -960 248042 480
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 252622 -960 252734 480
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259798 -960 259910 480
rect 260994 -960 261106 480
rect 262190 -960 262302 480
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 268078 -960 268190 480
rect 269274 -960 269386 480
rect 270470 -960 270582 480
rect 271666 -960 271778 480
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 280038 -960 280150 480
rect 281234 -960 281346 480
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 289514 -960 289626 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436990 -960 437102 480
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441774 -960 441886 480
rect 442970 -960 443082 480
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 459622 -960 459734 480
rect 460818 -960 460930 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509578 -960 509690 480
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528622 -960 528734 480
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 569010 -960 569122 480
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 24306 700440 24362 700496
rect 8114 700304 8170 700360
rect 89166 700576 89222 700632
rect 137834 700712 137890 700768
rect 3514 682216 3570 682272
rect 3422 667956 3478 667992
rect 3422 667936 3424 667956
rect 3424 667936 3476 667956
rect 3476 667936 3478 667956
rect 3054 653520 3110 653576
rect 3422 624824 3478 624880
rect 3422 623736 3478 623792
rect 3422 610408 3478 610464
rect 3422 595992 3478 596048
rect 3238 509904 3294 509960
rect 3330 495508 3386 495544
rect 3330 495488 3332 495508
rect 3332 495488 3384 495508
rect 3384 495488 3386 495508
rect 3146 481072 3202 481128
rect 3514 567296 3570 567352
rect 3606 553016 3662 553072
rect 3698 538600 3754 538656
rect 298006 606600 298062 606656
rect 297914 605376 297970 605432
rect 297822 603744 297878 603800
rect 297730 602520 297786 602576
rect 297638 600888 297694 600944
rect 297546 599800 297602 599856
rect 297454 598032 297510 598088
rect 297362 540232 297418 540288
rect 297270 538464 297326 538520
rect 256698 478916 256754 478952
rect 256698 478896 256700 478916
rect 256700 478896 256752 478916
rect 256752 478896 256754 478916
rect 3422 452376 3478 452432
rect 3146 437960 3202 438016
rect 3238 423680 3294 423736
rect 3146 394984 3202 395040
rect 3238 380568 3294 380624
rect 3146 366152 3202 366208
rect 3422 337456 3478 337512
rect 3238 323040 3294 323096
rect 3330 308760 3386 308816
rect 3422 294344 3478 294400
rect 3422 280100 3424 280120
rect 3424 280100 3476 280120
rect 3476 280100 3478 280120
rect 3422 280064 3478 280100
rect 3422 265648 3478 265704
rect 3514 251232 3570 251288
rect 3514 240760 3570 240816
rect 3422 236952 3478 237008
rect 3146 222536 3202 222592
rect 3422 208120 3478 208176
rect 3974 201048 4030 201104
rect 3422 200912 3478 200968
rect 3790 200776 3846 200832
rect 3606 200640 3662 200696
rect 3514 179424 3570 179480
rect 4066 193840 4122 193896
rect 3974 165008 4030 165064
rect 3790 150728 3846 150784
rect 3606 136312 3662 136368
rect 3422 122032 3478 122088
rect 3238 107616 3294 107672
rect 3422 80008 3478 80064
rect 3422 78920 3478 78976
rect 3330 50904 3386 50960
rect 3330 50088 3386 50144
rect 3422 8200 3478 8256
rect 3422 7112 3478 7168
rect 38658 93508 38660 93528
rect 38660 93508 38712 93528
rect 38712 93508 38714 93528
rect 38658 93472 38714 93508
rect 48134 93608 48190 93664
rect 72422 93880 72478 93936
rect 72422 93608 72478 93664
rect 91742 93880 91798 93936
rect 91742 93608 91798 93664
rect 111062 93880 111118 93936
rect 111062 93608 111118 93664
rect 130382 93880 130438 93936
rect 130382 93608 130438 93664
rect 256698 476720 256754 476776
rect 256698 474680 256754 474736
rect 256698 472504 256754 472560
rect 256698 470328 256754 470384
rect 256698 468288 256754 468344
rect 256698 466112 256754 466168
rect 256698 464072 256754 464128
rect 256698 461896 256754 461952
rect 256698 459720 256754 459776
rect 256698 457680 256754 457736
rect 256698 455504 256754 455560
rect 256698 453328 256754 453384
rect 256698 451308 256754 451344
rect 256698 451288 256700 451308
rect 256700 451288 256752 451308
rect 256752 451288 256754 451308
rect 256698 449112 256754 449168
rect 256698 447072 256754 447128
rect 256698 444896 256754 444952
rect 256698 442720 256754 442776
rect 256698 440680 256754 440736
rect 256698 438504 256754 438560
rect 256698 436328 256754 436384
rect 256698 434288 256754 434344
rect 256698 432112 256754 432168
rect 256698 430072 256754 430128
rect 256698 427896 256754 427952
rect 256698 425720 256754 425776
rect 256698 423700 256754 423736
rect 256698 423680 256700 423700
rect 256700 423680 256752 423700
rect 256752 423680 256754 423700
rect 256698 421504 256754 421560
rect 256698 419464 256754 419520
rect 256698 417288 256754 417344
rect 256698 415112 256754 415168
rect 256698 413072 256754 413128
rect 256698 410896 256754 410952
rect 256698 408720 256754 408776
rect 256698 406680 256754 406736
rect 256698 404504 256754 404560
rect 256698 402464 256754 402520
rect 256698 400288 256754 400344
rect 256698 398112 256754 398168
rect 256698 396092 256754 396128
rect 256698 396072 256700 396092
rect 256700 396072 256752 396092
rect 256752 396072 256754 396092
rect 256698 393896 256754 393952
rect 256698 391720 256754 391776
rect 256698 389680 256754 389736
rect 256698 387504 256754 387560
rect 256698 385464 256754 385520
rect 256698 383288 256754 383344
rect 256698 381112 256754 381168
rect 256698 379072 256754 379128
rect 256698 376896 256754 376952
rect 256698 374856 256754 374912
rect 256698 372680 256754 372736
rect 256698 370504 256754 370560
rect 256698 368500 256700 368520
rect 256700 368500 256752 368520
rect 256752 368500 256754 368520
rect 256698 368464 256754 368500
rect 256698 366288 256754 366344
rect 256698 364112 256754 364168
rect 256698 362072 256754 362128
rect 256698 359896 256754 359952
rect 256698 357856 256754 357912
rect 256698 355680 256754 355736
rect 256698 353504 256754 353560
rect 256698 351464 256754 351520
rect 256698 349288 256754 349344
rect 256698 347112 256754 347168
rect 256698 345092 256754 345128
rect 256698 345072 256700 345092
rect 256700 345072 256752 345092
rect 256752 345072 256754 345092
rect 256698 342896 256754 342952
rect 256698 340892 256700 340912
rect 256700 340892 256752 340912
rect 256752 340892 256754 340912
rect 256698 340856 256754 340892
rect 256698 338680 256754 338736
rect 256698 336504 256754 336560
rect 256698 334464 256754 334520
rect 256698 332288 256754 332344
rect 256698 330248 256754 330304
rect 256698 328072 256754 328128
rect 256698 325896 256754 325952
rect 256698 323856 256754 323912
rect 256698 321680 256754 321736
rect 256698 319504 256754 319560
rect 256698 317484 256754 317520
rect 256698 317464 256700 317484
rect 256700 317464 256752 317484
rect 256752 317464 256754 317484
rect 256698 315288 256754 315344
rect 256698 313284 256700 313304
rect 256700 313284 256752 313304
rect 256752 313284 256754 313304
rect 256698 313248 256754 313284
rect 256698 311072 256754 311128
rect 256698 308896 256754 308952
rect 256698 306856 256754 306912
rect 256698 304680 256754 304736
rect 256698 302504 256754 302560
rect 256698 300464 256754 300520
rect 256698 298288 256754 298344
rect 256698 296248 256754 296304
rect 256698 294072 256754 294128
rect 256698 291896 256754 291952
rect 256698 289876 256754 289912
rect 256698 289856 256700 289876
rect 256700 289856 256752 289876
rect 256752 289856 256754 289876
rect 256698 287680 256754 287736
rect 256698 285676 256700 285696
rect 256700 285676 256752 285696
rect 256752 285676 256754 285696
rect 256698 285640 256754 285676
rect 256698 283464 256754 283520
rect 256698 281288 256754 281344
rect 256698 279248 256754 279304
rect 256698 277072 256754 277128
rect 256698 274896 256754 274952
rect 256698 272856 256754 272912
rect 256698 270680 256754 270736
rect 256698 268640 256754 268696
rect 256698 266464 256754 266520
rect 256698 264288 256754 264344
rect 256698 262268 256754 262304
rect 256698 262248 256700 262268
rect 256700 262248 256752 262268
rect 256752 262248 256754 262268
rect 256698 260072 256754 260128
rect 256698 257896 256754 257952
rect 256698 255856 256754 255912
rect 256698 253680 256754 253736
rect 256698 251640 256754 251696
rect 256698 249464 256754 249520
rect 257342 247288 257398 247344
rect 256974 243072 257030 243128
rect 154486 93744 154542 93800
rect 140042 93608 140098 93664
rect 144918 93644 144920 93664
rect 144920 93644 144972 93664
rect 144972 93644 144974 93664
rect 144918 93608 144974 93644
rect 140042 93200 140098 93256
rect 257434 245248 257490 245304
rect 257986 241032 258042 241088
rect 263690 482160 263746 482216
rect 373630 612756 373632 612776
rect 373632 612756 373684 612776
rect 373684 612756 373686 612776
rect 373630 612720 373686 612756
rect 314566 518744 314622 518800
rect 320086 518744 320142 518800
rect 322938 518780 322940 518800
rect 322940 518780 322992 518800
rect 322992 518780 322994 518800
rect 322938 518744 322994 518780
rect 324318 518744 324374 518800
rect 325422 518744 325478 518800
rect 326434 518744 326490 518800
rect 327354 518780 327356 518800
rect 327356 518780 327408 518800
rect 327408 518780 327410 518800
rect 327354 518744 327410 518780
rect 328918 518744 328974 518800
rect 303618 518220 303674 518256
rect 303618 518200 303620 518220
rect 303620 518200 303672 518220
rect 303672 518200 303674 518220
rect 307574 517520 307630 517576
rect 313186 518608 313242 518664
rect 317234 518608 317290 518664
rect 318706 518628 318762 518664
rect 318706 518608 318708 518628
rect 318708 518608 318760 518628
rect 318760 518608 318762 518628
rect 314658 518472 314714 518528
rect 316038 518492 316094 518528
rect 316038 518472 316040 518492
rect 316040 518472 316092 518492
rect 316092 518472 316094 518492
rect 313278 518336 313334 518392
rect 321098 518608 321154 518664
rect 323122 518644 323124 518664
rect 323124 518644 323176 518664
rect 323176 518644 323178 518664
rect 323122 518608 323178 518644
rect 317326 518492 317382 518528
rect 317326 518472 317328 518492
rect 317328 518472 317380 518492
rect 317380 518472 317382 518492
rect 317510 518472 317566 518528
rect 315946 518084 316002 518120
rect 315946 518064 315948 518084
rect 315948 518064 316000 518084
rect 316000 518064 316002 518084
rect 317418 517928 317474 517984
rect 318798 518356 318854 518392
rect 318798 518336 318800 518356
rect 318800 518336 318852 518356
rect 318852 518336 318854 518356
rect 320178 518336 320234 518392
rect 321742 518200 321798 518256
rect 318798 518064 318854 518120
rect 325514 518472 325570 518528
rect 330114 518744 330170 518800
rect 331310 518764 331366 518800
rect 331310 518744 331312 518764
rect 331312 518744 331364 518764
rect 331364 518744 331366 518764
rect 332414 518744 332470 518800
rect 333794 518744 333850 518800
rect 334714 518744 334770 518800
rect 335818 518744 335874 518800
rect 336922 518780 336924 518800
rect 336924 518780 336976 518800
rect 336976 518780 336978 518800
rect 336922 518744 336978 518780
rect 338118 518744 338174 518800
rect 339498 518744 339554 518800
rect 340602 518764 340658 518800
rect 340602 518744 340604 518764
rect 340604 518744 340656 518764
rect 340656 518744 340658 518764
rect 331402 518608 331458 518664
rect 329838 518472 329894 518528
rect 312174 517792 312230 517848
rect 310242 517656 310298 517712
rect 309046 517520 309102 517576
rect 310334 517520 310390 517576
rect 311806 517520 311862 517576
rect 320178 482044 320234 482080
rect 320178 482024 320180 482044
rect 320180 482024 320232 482044
rect 320232 482024 320234 482044
rect 321558 482044 321614 482080
rect 321558 482024 321560 482044
rect 321560 482024 321612 482044
rect 321612 482024 321614 482044
rect 324502 517656 324558 517712
rect 324410 517520 324466 517576
rect 325698 517656 325754 517712
rect 327170 517656 327226 517712
rect 328458 517656 328514 517712
rect 332690 518200 332746 518256
rect 332598 517656 332654 517712
rect 336738 518336 336794 518392
rect 341522 518744 341578 518800
rect 345294 518780 345296 518800
rect 345296 518780 345348 518800
rect 345348 518780 345350 518800
rect 345294 518744 345350 518780
rect 346582 518764 346638 518800
rect 346582 518744 346584 518764
rect 346584 518744 346636 518764
rect 346636 518744 346638 518764
rect 339590 518608 339646 518664
rect 338118 518336 338174 518392
rect 339498 518336 339554 518392
rect 340878 518200 340934 518256
rect 342994 518472 343050 518528
rect 348974 518744 349030 518800
rect 343730 518336 343786 518392
rect 347686 518628 347742 518664
rect 347686 518608 347688 518628
rect 347688 518608 347740 518628
rect 347740 518608 347742 518628
rect 347778 518472 347834 518528
rect 333978 517812 334034 517848
rect 333978 517792 333980 517812
rect 333980 517792 334032 517812
rect 334032 517792 334034 517812
rect 342258 517792 342314 517848
rect 335358 517656 335414 517712
rect 343638 517676 343694 517712
rect 343638 517656 343640 517676
rect 343640 517656 343692 517676
rect 343692 517656 343694 517676
rect 345202 517656 345258 517712
rect 346398 517656 346454 517712
rect 347870 517792 347926 517848
rect 379702 609592 379758 609648
rect 379978 609592 380034 609648
rect 379610 549344 379666 549400
rect 379794 540912 379850 540968
rect 379702 482160 379758 482216
rect 488538 612756 488540 612776
rect 488540 612756 488592 612776
rect 488592 612756 488594 612776
rect 488538 612720 488594 612756
rect 493966 612756 493968 612776
rect 493968 612756 494020 612776
rect 494020 612756 494022 612776
rect 493966 612720 494022 612756
rect 496450 609864 496506 609920
rect 416778 606056 416834 606112
rect 416778 604832 416834 604888
rect 416778 603200 416834 603256
rect 416778 601976 416834 602032
rect 416778 600480 416834 600536
rect 417422 599256 417478 599312
rect 416962 539688 417018 539744
rect 416778 538328 416834 538384
rect 417514 597624 417570 597680
rect 499578 549480 499634 549536
rect 499578 542000 499634 542056
rect 499578 540912 499634 540968
rect 425334 519696 425390 519752
rect 434166 519696 434222 519752
rect 423678 518220 423734 518256
rect 423678 518200 423680 518220
rect 423680 518200 423732 518220
rect 423732 518200 423734 518220
rect 429290 518608 429346 518664
rect 426438 518472 426494 518528
rect 430578 518356 430634 518392
rect 430578 518336 430580 518356
rect 430580 518336 430632 518356
rect 430632 518336 430634 518356
rect 429198 518200 429254 518256
rect 432602 517792 432658 517848
rect 433246 517656 433302 517712
rect 443182 518744 443238 518800
rect 442538 518608 442594 518664
rect 435362 518336 435418 518392
rect 435914 518356 435970 518392
rect 435914 518336 435916 518356
rect 435916 518336 435968 518356
rect 435968 518336 435970 518356
rect 434626 517656 434682 517712
rect 434074 495488 434130 495544
rect 433890 492652 433946 492688
rect 433890 492632 433892 492652
rect 433892 492632 433944 492652
rect 433944 492632 433946 492652
rect 433614 482976 433670 483032
rect 433798 482976 433854 483032
rect 436926 518220 436982 518256
rect 436926 518200 436928 518220
rect 436928 518200 436980 518220
rect 436980 518200 436982 518220
rect 440882 518200 440938 518256
rect 436006 517656 436062 517712
rect 437294 517792 437350 517848
rect 437386 517656 437442 517712
rect 438674 517656 438730 517712
rect 438122 517520 438178 517576
rect 438766 517520 438822 517576
rect 439502 517520 439558 517576
rect 440146 517520 440202 517576
rect 441526 517520 441582 517576
rect 442906 517520 442962 517576
rect 444286 518608 444342 518664
rect 445390 518608 445446 518664
rect 446402 518608 446458 518664
rect 444102 518472 444158 518528
rect 445482 518472 445538 518528
rect 445574 518336 445630 518392
rect 447138 518472 447194 518528
rect 447966 518492 448022 518528
rect 447966 518472 447968 518492
rect 447968 518472 448020 518492
rect 448020 518472 448022 518492
rect 447046 518336 447102 518392
rect 448334 518200 448390 518256
rect 451278 518764 451334 518800
rect 451278 518744 451280 518764
rect 451280 518744 451332 518764
rect 451332 518744 451334 518764
rect 452566 518744 452622 518800
rect 448702 518472 448758 518528
rect 449806 517520 449862 517576
rect 450174 518336 450230 518392
rect 451186 517520 451242 517576
rect 452566 517520 452622 517576
rect 453762 518472 453818 518528
rect 455326 518472 455382 518528
rect 453854 517656 453910 517712
rect 453946 517520 454002 517576
rect 455326 517520 455382 517576
rect 458362 518780 458364 518800
rect 458364 518780 458416 518800
rect 458416 518780 458418 518800
rect 458362 518744 458418 518780
rect 459558 518764 459614 518800
rect 459558 518744 459560 518764
rect 459560 518744 459612 518764
rect 459612 518744 459614 518764
rect 457074 518644 457076 518664
rect 457076 518644 457128 518664
rect 457128 518644 457130 518664
rect 457074 518608 457130 518644
rect 456062 518472 456118 518528
rect 466458 518744 466514 518800
rect 461030 518608 461086 518664
rect 462318 518472 462374 518528
rect 463698 518472 463754 518528
rect 466458 518492 466514 518528
rect 466458 518472 466460 518492
rect 466460 518472 466512 518492
rect 466512 518472 466514 518492
rect 459558 518336 459614 518392
rect 465078 518336 465134 518392
rect 467838 518220 467894 518256
rect 467838 518200 467840 518220
rect 467840 518200 467892 518220
rect 467892 518200 467894 518220
rect 460846 517656 460902 517712
rect 469034 517656 469090 517712
rect 456706 517520 456762 517576
rect 458086 517520 458142 517576
rect 459466 517520 459522 517576
rect 460754 517520 460810 517576
rect 462226 517520 462282 517576
rect 463606 517520 463662 517576
rect 464986 517520 465042 517576
rect 466366 517520 466422 517576
rect 467746 517520 467802 517576
rect 466366 482432 466422 482488
rect 469126 517520 469182 517576
rect 469034 482296 469090 482352
rect 469126 482160 469182 482216
rect 471242 481752 471298 481808
rect 477222 481772 477278 481808
rect 477222 481752 477224 481772
rect 477224 481752 477276 481772
rect 477276 481752 477278 481772
rect 530858 482432 530914 482488
rect 536010 482296 536066 482352
rect 538586 482160 538642 482216
rect 539322 357312 539378 357368
rect 539506 412120 539562 412176
rect 539506 406408 539562 406464
rect 539506 405728 539562 405784
rect 539506 402192 539562 402248
rect 539506 391312 539562 391368
rect 539506 388592 539562 388648
rect 539506 373224 539562 373280
rect 539506 365644 539508 365664
rect 539508 365644 539560 365664
rect 539560 365644 539562 365664
rect 539506 365608 539562 365644
rect 539414 350648 539470 350704
rect 540242 394712 540298 394768
rect 540150 382064 540206 382120
rect 540058 377984 540114 378040
rect 539966 372000 540022 372056
rect 539874 369552 539930 369608
rect 540426 447344 540482 447400
rect 540334 363024 540390 363080
rect 539782 359488 539838 359544
rect 539690 353096 539746 353152
rect 539966 348880 540022 348936
rect 539598 346432 539654 346488
rect 539322 344256 539378 344312
rect 539782 331200 539838 331256
rect 539322 292712 539378 292768
rect 539322 292032 539378 292088
rect 539874 291896 539930 291952
rect 539322 286592 539378 286648
rect 539874 279112 539930 279168
rect 539782 273400 539838 273456
rect 539322 264968 539378 265024
rect 539782 264968 539838 265024
rect 357438 240660 357440 240680
rect 357440 240660 357492 240680
rect 357492 240660 357494 240680
rect 357438 240624 357494 240660
rect 366914 240624 366970 240680
rect 277306 204176 277362 204232
rect 274546 204040 274602 204096
rect 271786 203904 271842 203960
rect 269026 203768 269082 203824
rect 328366 203632 328422 203688
rect 329746 203632 329802 203688
rect 331126 203632 331182 203688
rect 328366 203396 328368 203416
rect 328368 203396 328420 203416
rect 328420 203396 328422 203416
rect 328366 203360 328422 203396
rect 331126 203260 331128 203280
rect 331128 203260 331180 203280
rect 331180 203260 331182 203280
rect 331126 203224 331182 203260
rect 329746 203088 329802 203144
rect 332414 203360 332470 203416
rect 333886 203360 333942 203416
rect 332506 203224 332562 203280
rect 334070 203632 334126 203688
rect 335174 203496 335230 203552
rect 333978 203224 334034 203280
rect 335358 203224 335414 203280
rect 333886 203088 333942 203144
rect 335266 203088 335322 203144
rect 336646 203380 336702 203416
rect 336646 203360 336648 203380
rect 336648 203360 336700 203380
rect 336700 203360 336702 203380
rect 336738 203224 336794 203280
rect 338118 203360 338174 203416
rect 339590 203516 339646 203552
rect 339590 203496 339592 203516
rect 339592 203496 339644 203516
rect 339644 203496 339646 203516
rect 340878 203496 340934 203552
rect 339498 203224 339554 203280
rect 342258 203668 342260 203688
rect 342260 203668 342312 203688
rect 342312 203668 342314 203688
rect 342258 203632 342314 203668
rect 343638 203632 343694 203688
rect 342166 203088 342222 203144
rect 336646 202952 336702 203008
rect 337934 202952 337990 203008
rect 339222 202952 339278 203008
rect 345018 203224 345074 203280
rect 346398 203088 346454 203144
rect 349158 203632 349214 203688
rect 351090 203632 351146 203688
rect 347778 203088 347834 203144
rect 349066 203496 349122 203552
rect 349158 203224 349214 203280
rect 342258 202952 342314 203008
rect 342442 202952 342498 203008
rect 343638 202952 343694 203008
rect 344926 202952 344982 203008
rect 345938 202952 345994 203008
rect 347134 202952 347190 203008
rect 348330 202952 348386 203008
rect 349250 202952 349306 203008
rect 351826 203632 351882 203688
rect 351918 203088 351974 203144
rect 353206 203088 353262 203144
rect 350998 202952 351054 203008
rect 351734 202952 351790 203008
rect 354678 203088 354734 203144
rect 356058 203124 356060 203144
rect 356060 203124 356112 203144
rect 356112 203124 356114 203144
rect 356058 203088 356114 203124
rect 357438 203360 357494 203416
rect 357806 203088 357862 203144
rect 366362 204176 366418 204232
rect 371146 204176 371202 204232
rect 367098 204040 367154 204096
rect 365718 203904 365774 203960
rect 364338 203768 364394 203824
rect 368478 203224 368534 203280
rect 353298 202988 353300 203008
rect 353300 202988 353352 203008
rect 353352 202988 353354 203008
rect 353298 202952 353354 202988
rect 354310 202952 354366 203008
rect 355598 202952 355654 203008
rect 356426 202952 356482 203008
rect 357438 202972 357494 203008
rect 357438 202952 357440 202972
rect 357440 202952 357492 202972
rect 357492 202952 357494 202972
rect 358634 202952 358690 203008
rect 360014 202952 360070 203008
rect 361302 202952 361358 203008
rect 362498 202952 362554 203008
rect 363510 202952 363566 203008
rect 364706 202952 364762 203008
rect 373262 203088 373318 203144
rect 379794 182688 379850 182744
rect 297914 180240 297970 180296
rect 297914 171808 297970 171864
rect 297822 111696 297878 111752
rect 379794 125568 379850 125624
rect 379978 125568 380034 125624
rect 380438 180920 380494 180976
rect 380806 123120 380862 123176
rect 380346 122032 380402 122088
rect 380254 120264 380310 120320
rect 379978 119176 380034 119232
rect 380806 118088 380862 118144
rect 449806 204076 449808 204096
rect 449808 204076 449860 204096
rect 449860 204076 449862 204096
rect 449806 204040 449862 204076
rect 449162 203360 449218 203416
rect 450542 203360 450598 203416
rect 451922 203360 451978 203416
rect 453302 203360 453358 203416
rect 451186 203224 451242 203280
rect 456614 204212 456616 204232
rect 456616 204212 456668 204232
rect 456668 204212 456670 204232
rect 456614 204176 456670 204212
rect 456154 203396 456156 203416
rect 456156 203396 456208 203416
rect 456208 203396 456210 203416
rect 456154 203360 456210 203396
rect 453946 203224 454002 203280
rect 454682 203224 454738 203280
rect 455050 203224 455106 203280
rect 455234 203224 455290 203280
rect 452566 202972 452622 203008
rect 452566 202952 452568 202972
rect 452568 202952 452620 202972
rect 452620 202952 452622 202972
rect 458086 203224 458142 203280
rect 459466 203360 459522 203416
rect 460846 203224 460902 203280
rect 462134 203360 462190 203416
rect 463514 203360 463570 203416
rect 463606 203224 463662 203280
rect 464618 203260 464620 203280
rect 464620 203260 464672 203280
rect 464672 203260 464674 203280
rect 464618 203224 464674 203260
rect 469126 204176 469182 204232
rect 470506 204176 470562 204232
rect 467746 204040 467802 204096
rect 470414 204040 470470 204096
rect 465078 203224 465134 203280
rect 466550 203260 466552 203280
rect 466552 203260 466604 203280
rect 466604 203260 466606 203280
rect 466550 203224 466606 203260
rect 471886 203224 471942 203280
rect 473266 203224 473322 203280
rect 455326 202988 455328 203008
rect 455328 202988 455380 203008
rect 455380 202988 455382 203008
rect 455326 202952 455382 202988
rect 456614 202952 456670 203008
rect 457994 202952 458050 203008
rect 459006 202952 459062 203008
rect 460570 202952 460626 203008
rect 461398 202952 461454 203008
rect 462410 202952 462466 203008
rect 463606 202952 463662 203008
rect 464986 202952 465042 203008
rect 466366 202952 466422 203008
rect 467286 202952 467342 203008
rect 468482 202952 468538 203008
rect 469402 202952 469458 203008
rect 470690 202952 470746 203008
rect 471610 202952 471666 203008
rect 471794 202952 471850 203008
rect 476946 207712 477002 207768
rect 476854 204040 476910 204096
rect 476670 203904 476726 203960
rect 477498 204176 477554 204232
rect 478142 204176 478198 204232
rect 477590 204040 477646 204096
rect 477682 203904 477738 203960
rect 477590 203360 477646 203416
rect 481638 204212 481640 204232
rect 481640 204212 481692 204232
rect 481692 204212 481694 204232
rect 481638 204176 481694 204212
rect 490194 204176 490250 204232
rect 485778 204040 485834 204096
rect 480442 203904 480498 203960
rect 483018 203668 483020 203688
rect 483020 203668 483072 203688
rect 483072 203668 483074 203688
rect 483018 203632 483074 203668
rect 484398 203496 484454 203552
rect 476026 203224 476082 203280
rect 477498 203224 477554 203280
rect 485778 203224 485834 203280
rect 472898 202952 472954 203008
rect 474186 202952 474242 203008
rect 475566 202952 475622 203008
rect 476118 202952 476174 203008
rect 478878 202952 478934 203008
rect 480626 202952 480682 203008
rect 481638 202952 481694 203008
rect 483018 202952 483074 203008
rect 484398 202952 484454 203008
rect 448426 201456 448482 201512
rect 540886 428304 540942 428360
rect 540794 426264 540850 426320
rect 540794 418376 540850 418432
rect 540702 417832 540758 417888
rect 540610 413616 540666 413672
rect 540978 415792 541034 415848
rect 540518 405184 540574 405240
rect 540610 399064 540666 399120
rect 540518 398520 540574 398576
rect 540610 395392 540666 395448
rect 541254 396752 541310 396808
rect 541162 392536 541218 392592
rect 541070 386280 541126 386336
rect 541622 449384 541678 449440
rect 541530 354728 541586 354784
rect 541438 348336 541494 348392
rect 541346 342080 541402 342136
rect 541162 279384 541218 279440
rect 538310 222808 538366 222864
rect 539966 216008 540022 216064
rect 538310 205400 538366 205456
rect 538218 203768 538274 203824
rect 543278 511944 543334 512000
rect 543462 511944 543518 512000
rect 543278 482976 543334 483032
rect 543462 482976 543518 483032
rect 541714 403144 541770 403200
rect 542266 466248 542322 466304
rect 542174 379888 542230 379944
rect 542082 373632 542138 373688
rect 541990 367240 542046 367296
rect 541898 360984 541954 361040
rect 541806 337864 541862 337920
rect 542174 241440 542230 241496
rect 539966 202952 540022 203008
rect 496450 181328 496506 181384
rect 417422 180512 417478 180568
rect 418066 171672 418122 171728
rect 380806 115812 380808 115832
rect 380808 115812 380860 115832
rect 380860 115812 380862 115832
rect 380806 115776 380862 115812
rect 380714 114688 380770 114744
rect 300766 111288 300822 111344
rect 416778 111288 416834 111344
rect 303618 108976 303674 109032
rect 307758 108976 307814 109032
rect 500130 123664 500186 123720
rect 500038 122032 500094 122088
rect 499946 120808 500002 120864
rect 499854 118632 499910 118688
rect 499762 118088 499818 118144
rect 499670 115776 499726 115832
rect 539966 193160 540022 193216
rect 539966 183640 540022 183696
rect 500314 183096 500370 183152
rect 540150 167048 540206 167104
rect 540150 164192 540206 164248
rect 539966 162560 540022 162616
rect 539966 153176 540022 153232
rect 539966 147736 540022 147792
rect 539966 144880 540022 144936
rect 539966 120672 540022 120728
rect 539966 115912 540022 115968
rect 500222 115232 500278 115288
rect 424230 108976 424286 109032
rect 427818 108976 427874 109032
rect 542358 445168 542414 445224
rect 542542 451560 542598 451616
rect 542450 440952 542506 441008
rect 542450 438912 542506 438968
rect 542450 243072 542506 243128
rect 542450 241032 542506 241088
rect 542634 430480 542690 430536
rect 542726 424088 542782 424144
rect 543278 436736 543334 436792
rect 543462 434696 543518 434752
rect 543646 453600 543702 453656
rect 543554 432520 543610 432576
rect 543186 422048 543242 422104
rect 543094 420008 543150 420064
rect 543002 409400 543058 409456
rect 542910 407360 542966 407416
rect 542818 400968 542874 401024
rect 543462 399472 543518 399528
rect 543462 389000 543518 389056
rect 543370 376624 543426 376680
rect 543462 369688 543518 369744
rect 543370 357312 543426 357368
rect 543462 350376 543518 350432
rect 543462 339904 543518 339960
rect 542634 335688 542690 335744
rect 542634 333648 542690 333704
rect 542634 331472 542690 331528
rect 542634 329432 542690 329488
rect 542634 327256 542690 327312
rect 542634 325216 542690 325272
rect 542634 323040 542690 323096
rect 542634 321000 542690 321056
rect 542634 318824 542690 318880
rect 542634 316784 542690 316840
rect 542634 314628 542690 314664
rect 542634 314608 542636 314628
rect 542636 314608 542688 314628
rect 542688 314608 542690 314628
rect 542634 312568 542690 312624
rect 542634 310392 542690 310448
rect 542634 308352 542690 308408
rect 542634 306176 542690 306232
rect 542634 304136 542690 304192
rect 542634 301960 542690 302016
rect 542634 299920 542690 299976
rect 542634 297880 542690 297936
rect 542634 295704 542690 295760
rect 542634 293664 542690 293720
rect 542634 291488 542690 291544
rect 542634 289448 542690 289504
rect 542634 287272 542690 287328
rect 542634 285232 542690 285288
rect 542634 283056 542690 283112
rect 542634 281016 542690 281072
rect 543094 276800 543150 276856
rect 542634 274624 542690 274680
rect 543002 272584 543058 272640
rect 542634 257760 542690 257816
rect 542634 255720 542690 255776
rect 542634 253544 542690 253600
rect 543462 270408 543518 270464
rect 543370 266192 543426 266248
rect 543278 261976 543334 262032
rect 543094 259936 543150 259992
rect 543094 251504 543150 251560
rect 542634 249328 542690 249384
rect 542634 247288 542690 247344
rect 542910 245112 542966 245168
rect 542910 241440 542966 241496
rect 543002 173884 543004 173904
rect 543004 173884 543056 173904
rect 543056 173884 543058 173904
rect 543002 173848 543058 173884
rect 543002 164192 543058 164248
rect 543554 268368 543610 268424
rect 580170 697992 580226 698048
rect 580170 686296 580226 686352
rect 580170 674600 580226 674656
rect 580170 651072 580226 651128
rect 580170 639376 580226 639432
rect 580170 627680 580226 627736
rect 580170 604152 580226 604208
rect 580170 592456 580226 592512
rect 580170 580760 580226 580816
rect 580170 557232 580226 557288
rect 580170 545536 580226 545592
rect 580170 533840 580226 533896
rect 580170 510312 580226 510368
rect 580170 498616 580226 498672
rect 580170 486784 580226 486840
rect 580170 463392 580226 463448
rect 580170 451696 580226 451752
rect 580170 439864 580226 439920
rect 580170 416472 580226 416528
rect 580170 404776 580226 404832
rect 580170 392944 580226 393000
rect 580262 369552 580318 369608
rect 580354 357856 580410 357912
rect 580446 346024 580502 346080
rect 580538 322632 580594 322688
rect 580630 310800 580686 310856
rect 580722 299104 580778 299160
rect 580170 275712 580226 275768
rect 544382 264152 544438 264208
rect 580170 263880 580226 263936
rect 542910 77152 542966 77208
rect 543186 106256 543242 106312
rect 543370 106256 543426 106312
rect 543186 77152 543242 77208
rect 579802 252184 579858 252240
rect 580170 228792 580226 228848
rect 580170 216960 580226 217016
rect 579802 205264 579858 205320
rect 580170 181872 580226 181928
rect 580170 170040 580226 170096
rect 579802 158344 579858 158400
rect 580170 134816 580226 134872
rect 580170 123120 580226 123176
rect 579802 111424 579858 111480
rect 580170 87896 580226 87952
rect 580170 76200 580226 76256
rect 579802 64504 579858 64560
rect 580170 40976 580226 41032
rect 580170 29280 580226 29336
rect 579802 17584 579858 17640
<< metal3 >>
rect 137829 700770 137895 700773
rect 538254 700770 538260 700772
rect 137829 700768 538260 700770
rect 137829 700712 137834 700768
rect 137890 700712 538260 700768
rect 137829 700710 538260 700712
rect 137829 700707 137895 700710
rect 538254 700708 538260 700710
rect 538324 700708 538330 700772
rect 89161 700634 89227 700637
rect 538438 700634 538444 700636
rect 89161 700632 538444 700634
rect 89161 700576 89166 700632
rect 89222 700576 538444 700632
rect 89161 700574 538444 700576
rect 89161 700571 89227 700574
rect 538438 700572 538444 700574
rect 538508 700572 538514 700636
rect 24301 700498 24367 700501
rect 540094 700498 540100 700500
rect 24301 700496 540100 700498
rect 24301 700440 24306 700496
rect 24362 700440 540100 700496
rect 24301 700438 540100 700440
rect 24301 700435 24367 700438
rect 540094 700436 540100 700438
rect 540164 700436 540170 700500
rect 8109 700362 8175 700365
rect 539910 700362 539916 700364
rect 8109 700360 539916 700362
rect 8109 700304 8114 700360
rect 8170 700304 539916 700360
rect 8109 700302 539916 700304
rect 8109 700299 8175 700302
rect 539910 700300 539916 700302
rect 539980 700300 539986 700364
rect 580165 698050 580231 698053
rect 583520 698050 584960 698140
rect 580165 698048 584960 698050
rect 580165 697992 580170 698048
rect 580226 697992 584960 698048
rect 580165 697990 584960 697992
rect 580165 697987 580231 697990
rect 583520 697900 584960 697990
rect -960 696540 480 696780
rect 580165 686354 580231 686357
rect 583520 686354 584960 686444
rect 580165 686352 584960 686354
rect 580165 686296 580170 686352
rect 580226 686296 584960 686352
rect 580165 686294 584960 686296
rect 580165 686291 580231 686294
rect 583520 686204 584960 686294
rect -960 682274 480 682364
rect 3509 682274 3575 682277
rect -960 682272 3575 682274
rect -960 682216 3514 682272
rect 3570 682216 3575 682272
rect -960 682214 3575 682216
rect -960 682124 480 682214
rect 3509 682211 3575 682214
rect 580165 674658 580231 674661
rect 583520 674658 584960 674748
rect 580165 674656 584960 674658
rect 580165 674600 580170 674656
rect 580226 674600 584960 674656
rect 580165 674598 584960 674600
rect 580165 674595 580231 674598
rect 583520 674508 584960 674598
rect -960 667994 480 668084
rect 3417 667994 3483 667997
rect -960 667992 3483 667994
rect -960 667936 3422 667992
rect 3478 667936 3483 667992
rect -960 667934 3483 667936
rect -960 667844 480 667934
rect 3417 667931 3483 667934
rect 583520 662676 584960 662916
rect -960 653578 480 653668
rect 3049 653578 3115 653581
rect -960 653576 3115 653578
rect -960 653520 3054 653576
rect 3110 653520 3115 653576
rect -960 653518 3115 653520
rect -960 653428 480 653518
rect 3049 653515 3115 653518
rect 580165 651130 580231 651133
rect 583520 651130 584960 651220
rect 580165 651128 584960 651130
rect 580165 651072 580170 651128
rect 580226 651072 584960 651128
rect 580165 651070 584960 651072
rect 580165 651067 580231 651070
rect 583520 650980 584960 651070
rect 580165 639434 580231 639437
rect 583520 639434 584960 639524
rect 580165 639432 584960 639434
rect 580165 639376 580170 639432
rect 580226 639376 584960 639432
rect 580165 639374 584960 639376
rect 580165 639371 580231 639374
rect 583520 639284 584960 639374
rect -960 639012 480 639252
rect 580165 627738 580231 627741
rect 583520 627738 584960 627828
rect 580165 627736 584960 627738
rect 580165 627680 580170 627736
rect 580226 627680 584960 627736
rect 580165 627678 584960 627680
rect 580165 627675 580231 627678
rect 583520 627588 584960 627678
rect -960 624882 480 624972
rect 3417 624882 3483 624885
rect -960 624880 3483 624882
rect -960 624824 3422 624880
rect 3478 624824 3483 624880
rect -960 624822 3483 624824
rect -960 624732 480 624822
rect 3417 624819 3483 624822
rect 3417 623794 3483 623797
rect 538806 623794 538812 623796
rect 3417 623792 538812 623794
rect 3417 623736 3422 623792
rect 3478 623736 538812 623792
rect 3417 623734 538812 623736
rect 3417 623731 3483 623734
rect 538806 623732 538812 623734
rect 538876 623732 538882 623796
rect 583520 615756 584960 615996
rect 373625 612780 373691 612781
rect 373574 612716 373580 612780
rect 373644 612778 373691 612780
rect 488533 612780 488599 612781
rect 493961 612780 494027 612781
rect 373644 612776 373736 612778
rect 373686 612720 373736 612776
rect 373644 612718 373736 612720
rect 488533 612776 488580 612780
rect 488644 612778 488650 612780
rect 493910 612778 493916 612780
rect 488533 612720 488538 612776
rect 373644 612716 373691 612718
rect 373625 612715 373691 612716
rect 488533 612716 488580 612720
rect 488644 612718 488690 612778
rect 493870 612718 493916 612778
rect 493980 612776 494027 612780
rect 494022 612720 494027 612776
rect 488644 612716 488650 612718
rect 493910 612716 493916 612718
rect 493980 612716 494027 612720
rect 488533 612715 488599 612716
rect 493961 612715 494027 612716
rect 369158 610948 369164 611012
rect 369228 611010 369234 611012
rect 373022 611010 373028 611012
rect 369228 610950 373028 611010
rect 369228 610948 369234 610950
rect 373022 610948 373028 610950
rect 373092 610948 373098 611012
rect -960 610466 480 610556
rect 3417 610466 3483 610469
rect -960 610464 3483 610466
rect -960 610408 3422 610464
rect 3478 610408 3483 610464
rect -960 610406 3483 610408
rect -960 610316 480 610406
rect 3417 610403 3483 610406
rect 496445 609922 496511 609925
rect 496445 609920 496554 609922
rect 496445 609864 496450 609920
rect 496506 609864 496554 609920
rect 496445 609859 496554 609864
rect 377292 609653 377874 609713
rect 496494 609683 496554 609859
rect 377814 609650 377874 609653
rect 379697 609650 379763 609653
rect 379973 609650 380039 609653
rect 377814 609648 380039 609650
rect 377814 609592 379702 609648
rect 379758 609592 379978 609648
rect 380034 609592 380039 609648
rect 377814 609590 380039 609592
rect 379697 609587 379763 609590
rect 379973 609587 380039 609590
rect 298001 606658 298067 606661
rect 298001 606656 299490 606658
rect 298001 606600 298006 606656
rect 298062 606617 299490 606656
rect 298062 606600 300012 606617
rect 298001 606598 300012 606600
rect 298001 606595 298067 606598
rect 299430 606557 300012 606598
rect 416773 606114 416839 606117
rect 420134 606114 420194 606587
rect 416773 606112 420194 606114
rect 416773 606056 416778 606112
rect 416834 606056 420194 606112
rect 416773 606054 420194 606056
rect 416773 606051 416839 606054
rect 297909 605434 297975 605437
rect 299430 605434 300012 605489
rect 297909 605432 300012 605434
rect 297909 605376 297914 605432
rect 297970 605429 300012 605432
rect 297970 605376 299490 605429
rect 297909 605374 299490 605376
rect 297909 605371 297975 605374
rect 416773 604890 416839 604893
rect 420134 604890 420194 605459
rect 416773 604888 420194 604890
rect 416773 604832 416778 604888
rect 416834 604832 420194 604888
rect 416773 604830 420194 604832
rect 416773 604827 416839 604830
rect 580165 604210 580231 604213
rect 583520 604210 584960 604300
rect 580165 604208 584960 604210
rect 580165 604152 580170 604208
rect 580226 604152 584960 604208
rect 580165 604150 584960 604152
rect 580165 604147 580231 604150
rect 583520 604060 584960 604150
rect 297817 603802 297883 603805
rect 297817 603800 299490 603802
rect 297817 603744 297822 603800
rect 297878 603789 299490 603800
rect 297878 603744 300012 603789
rect 297817 603742 300012 603744
rect 297817 603739 297883 603742
rect 299430 603729 300012 603742
rect 416773 603258 416839 603261
rect 420134 603258 420194 603759
rect 416773 603256 420194 603258
rect 416773 603200 416778 603256
rect 416834 603200 420194 603256
rect 416773 603198 420194 603200
rect 416773 603195 416839 603198
rect 299430 602601 300012 602661
rect 297725 602578 297791 602581
rect 299430 602578 299490 602601
rect 297725 602576 299490 602578
rect 297725 602520 297730 602576
rect 297786 602520 299490 602576
rect 297725 602518 299490 602520
rect 297725 602515 297791 602518
rect 416773 602034 416839 602037
rect 420134 602034 420194 602631
rect 416773 602032 420194 602034
rect 416773 601976 416778 602032
rect 416834 601976 420194 602032
rect 416773 601974 420194 601976
rect 416773 601971 416839 601974
rect 297633 600946 297699 600949
rect 299430 600946 300012 600961
rect 297633 600944 300012 600946
rect 297633 600888 297638 600944
rect 297694 600901 300012 600944
rect 297694 600888 299490 600901
rect 297633 600886 299490 600888
rect 297633 600883 297699 600886
rect 416773 600538 416839 600541
rect 420134 600538 420194 600931
rect 416773 600536 420194 600538
rect 416773 600480 416778 600536
rect 416834 600480 420194 600536
rect 416773 600478 420194 600480
rect 416773 600475 416839 600478
rect 297541 599858 297607 599861
rect 297541 599856 299490 599858
rect 297541 599800 297546 599856
rect 297602 599833 299490 599856
rect 297602 599800 300012 599833
rect 297541 599798 300012 599800
rect 297541 599795 297607 599798
rect 299430 599773 300012 599798
rect 417417 599314 417483 599317
rect 420134 599314 420194 599803
rect 417417 599312 420194 599314
rect 417417 599256 417422 599312
rect 417478 599256 420194 599312
rect 417417 599254 420194 599256
rect 417417 599251 417483 599254
rect 297449 598090 297515 598093
rect 299430 598090 300012 598133
rect 297449 598088 300012 598090
rect 297449 598032 297454 598088
rect 297510 598073 300012 598088
rect 297510 598032 299490 598073
rect 297449 598030 299490 598032
rect 297449 598027 297515 598030
rect 417509 597682 417575 597685
rect 420134 597682 420194 598103
rect 417509 597680 420194 597682
rect 417509 597624 417514 597680
rect 417570 597624 420194 597680
rect 417509 597622 420194 597624
rect 417509 597619 417575 597622
rect -960 596050 480 596140
rect 3417 596050 3483 596053
rect -960 596048 3483 596050
rect -960 595992 3422 596048
rect 3478 595992 3483 596048
rect -960 595990 3483 595992
rect -960 595900 480 595990
rect 3417 595987 3483 595990
rect 580165 592514 580231 592517
rect 583520 592514 584960 592604
rect 580165 592512 584960 592514
rect 580165 592456 580170 592512
rect 580226 592456 584960 592512
rect 580165 592454 584960 592456
rect 580165 592451 580231 592454
rect 583520 592364 584960 592454
rect -960 581620 480 581860
rect 580165 580818 580231 580821
rect 583520 580818 584960 580908
rect 580165 580816 584960 580818
rect 580165 580760 580170 580816
rect 580226 580760 584960 580816
rect 580165 580758 584960 580760
rect 580165 580755 580231 580758
rect 583520 580668 584960 580758
rect 583520 568836 584960 569076
rect -960 567354 480 567444
rect 3509 567354 3575 567357
rect -960 567352 3575 567354
rect -960 567296 3514 567352
rect 3570 567296 3575 567352
rect -960 567294 3575 567296
rect -960 567204 480 567294
rect 3509 567291 3575 567294
rect 580165 557290 580231 557293
rect 583520 557290 584960 557380
rect 580165 557288 584960 557290
rect 580165 557232 580170 557288
rect 580226 557232 584960 557288
rect 580165 557230 584960 557232
rect 580165 557227 580231 557230
rect 583520 557140 584960 557230
rect -960 553074 480 553164
rect 3601 553074 3667 553077
rect -960 553072 3667 553074
rect -960 553016 3606 553072
rect 3662 553016 3667 553072
rect -960 553014 3667 553016
rect -960 552924 480 553014
rect 3601 553011 3667 553014
rect 499573 549538 499639 549541
rect 497782 549536 499639 549538
rect 497782 549480 499578 549536
rect 499634 549480 499639 549536
rect 497782 549478 499639 549480
rect 497782 549442 497842 549478
rect 499573 549475 499639 549478
rect 377108 549412 377874 549442
rect 497076 549412 497842 549442
rect 377078 549402 377874 549412
rect 379605 549402 379671 549405
rect 377078 549400 379671 549402
rect 377078 549382 379610 549400
rect 377078 540958 377138 549382
rect 377814 549344 379610 549382
rect 379666 549344 379671 549400
rect 377814 549342 379671 549344
rect 379605 549339 379671 549342
rect 497046 549382 497842 549412
rect 497046 547906 497106 549382
rect 497046 547846 497290 547906
rect 497230 542058 497290 547846
rect 580165 545594 580231 545597
rect 583520 545594 584960 545684
rect 580165 545592 584960 545594
rect 580165 545536 580170 545592
rect 580226 545536 584960 545592
rect 580165 545534 584960 545536
rect 580165 545531 580231 545534
rect 583520 545444 584960 545534
rect 499573 542058 499639 542061
rect 497230 542056 499639 542058
rect 497230 542000 499578 542056
rect 499634 542000 499639 542056
rect 497230 541998 499639 542000
rect 499573 541995 499639 541998
rect 379789 540970 379855 540973
rect 499573 540970 499639 540973
rect 377446 540968 379855 540970
rect 377446 540958 379794 540968
rect 377078 540928 379794 540958
rect 377108 540912 379794 540928
rect 379850 540912 379855 540968
rect 377108 540910 379855 540912
rect 497230 540968 499639 540970
rect 497230 540912 499578 540968
rect 499634 540912 499639 540968
rect 497230 540910 499639 540912
rect 377108 540898 377506 540910
rect 379789 540907 379855 540910
rect 499573 540907 499639 540910
rect 297357 540290 297423 540293
rect 297357 540288 299490 540290
rect 297357 540232 297362 540288
rect 297418 540285 299490 540288
rect 297418 540232 300012 540285
rect 297357 540230 300012 540232
rect 297357 540227 297423 540230
rect 299430 540225 300012 540230
rect 416957 539746 417023 539749
rect 420134 539746 420194 540255
rect 416957 539744 420194 539746
rect 416957 539688 416962 539744
rect 417018 539688 420194 539744
rect 416957 539686 420194 539688
rect 416957 539683 417023 539686
rect -960 538658 480 538748
rect 3693 538658 3759 538661
rect -960 538656 3759 538658
rect -960 538600 3698 538656
rect 3754 538600 3759 538656
rect -960 538598 3759 538600
rect -960 538508 480 538598
rect 3693 538595 3759 538598
rect 299430 538525 300012 538585
rect 297265 538522 297331 538525
rect 299430 538522 299490 538525
rect 297265 538520 299490 538522
rect 297265 538464 297270 538520
rect 297326 538464 299490 538520
rect 297265 538462 299490 538464
rect 297265 538459 297331 538462
rect 416773 538386 416839 538389
rect 420134 538386 420194 538555
rect 416773 538384 420194 538386
rect 416773 538328 416778 538384
rect 416834 538328 420194 538384
rect 416773 538326 420194 538328
rect 416773 538323 416839 538326
rect 580165 533898 580231 533901
rect 583520 533898 584960 533988
rect 580165 533896 584960 533898
rect 580165 533840 580170 533896
rect 580226 533840 584960 533896
rect 580165 533838 584960 533840
rect 580165 533835 580231 533838
rect 583520 533748 584960 533838
rect -960 524092 480 524332
rect 583520 521916 584960 522156
rect 425329 519754 425395 519757
rect 427962 519754 427968 519756
rect 425329 519752 427968 519754
rect 425329 519696 425334 519752
rect 425390 519696 427968 519752
rect 425329 519694 427968 519696
rect 425329 519691 425395 519694
rect 427962 519692 427968 519694
rect 428032 519692 428038 519756
rect 433802 519692 433808 519756
rect 433872 519754 433878 519756
rect 434161 519754 434227 519757
rect 433872 519752 434227 519754
rect 433872 519696 434166 519752
rect 434222 519696 434227 519752
rect 433872 519694 434227 519696
rect 433872 519692 433878 519694
rect 434161 519691 434227 519694
rect 313774 518740 313780 518804
rect 313844 518802 313850 518804
rect 314561 518802 314627 518805
rect 313844 518800 314627 518802
rect 313844 518744 314566 518800
rect 314622 518744 314627 518800
rect 313844 518742 314627 518744
rect 313844 518740 313850 518742
rect 314561 518739 314627 518742
rect 319662 518740 319668 518804
rect 319732 518802 319738 518804
rect 320081 518802 320147 518805
rect 319732 518800 320147 518802
rect 319732 518744 320086 518800
rect 320142 518744 320147 518800
rect 319732 518742 320147 518744
rect 319732 518740 319738 518742
rect 320081 518739 320147 518742
rect 322933 518802 322999 518805
rect 324313 518804 324379 518805
rect 323526 518802 323532 518804
rect 322933 518800 323532 518802
rect 322933 518744 322938 518800
rect 322994 518744 323532 518800
rect 322933 518742 323532 518744
rect 322933 518739 322999 518742
rect 323526 518740 323532 518742
rect 323596 518740 323602 518804
rect 324262 518802 324268 518804
rect 324222 518742 324268 518802
rect 324332 518800 324379 518804
rect 324374 518744 324379 518800
rect 324262 518740 324268 518742
rect 324332 518740 324379 518744
rect 325182 518740 325188 518804
rect 325252 518802 325258 518804
rect 325417 518802 325483 518805
rect 325252 518800 325483 518802
rect 325252 518744 325422 518800
rect 325478 518744 325483 518800
rect 325252 518742 325483 518744
rect 325252 518740 325258 518742
rect 324313 518739 324379 518740
rect 325417 518739 325483 518742
rect 326429 518804 326495 518805
rect 327349 518804 327415 518805
rect 328913 518804 328979 518805
rect 326429 518800 326476 518804
rect 326540 518802 326546 518804
rect 326429 518744 326434 518800
rect 326429 518740 326476 518744
rect 326540 518742 326586 518802
rect 327349 518800 327396 518804
rect 327460 518802 327466 518804
rect 328862 518802 328868 518804
rect 327349 518744 327354 518800
rect 326540 518740 326546 518742
rect 327349 518740 327396 518744
rect 327460 518742 327506 518802
rect 328822 518742 328868 518802
rect 328932 518800 328979 518804
rect 328974 518744 328979 518800
rect 327460 518740 327466 518742
rect 328862 518740 328868 518742
rect 328932 518740 328979 518744
rect 326429 518739 326495 518740
rect 327349 518739 327415 518740
rect 328913 518739 328979 518740
rect 330109 518804 330175 518805
rect 330109 518800 330156 518804
rect 330220 518802 330226 518804
rect 331305 518802 331371 518805
rect 332409 518804 332475 518805
rect 331622 518802 331628 518804
rect 330109 518744 330114 518800
rect 330109 518740 330156 518744
rect 330220 518742 330266 518802
rect 331305 518800 331628 518802
rect 331305 518744 331310 518800
rect 331366 518744 331628 518800
rect 331305 518742 331628 518744
rect 330220 518740 330226 518742
rect 330109 518739 330175 518740
rect 331305 518739 331371 518742
rect 331622 518740 331628 518742
rect 331692 518740 331698 518804
rect 332358 518802 332364 518804
rect 332318 518742 332364 518802
rect 332428 518800 332475 518804
rect 332470 518744 332475 518800
rect 332358 518740 332364 518742
rect 332428 518740 332475 518744
rect 333646 518740 333652 518804
rect 333716 518802 333722 518804
rect 333789 518802 333855 518805
rect 333716 518800 333855 518802
rect 333716 518744 333794 518800
rect 333850 518744 333855 518800
rect 333716 518742 333855 518744
rect 333716 518740 333722 518742
rect 332409 518739 332475 518740
rect 333789 518739 333855 518742
rect 334566 518740 334572 518804
rect 334636 518802 334642 518804
rect 334709 518802 334775 518805
rect 334636 518800 334775 518802
rect 334636 518744 334714 518800
rect 334770 518744 334775 518800
rect 334636 518742 334775 518744
rect 334636 518740 334642 518742
rect 334709 518739 334775 518742
rect 335813 518804 335879 518805
rect 336917 518804 336983 518805
rect 338113 518804 338179 518805
rect 335813 518800 335860 518804
rect 335924 518802 335930 518804
rect 335813 518744 335818 518800
rect 335813 518740 335860 518744
rect 335924 518742 335970 518802
rect 336917 518800 336964 518804
rect 337028 518802 337034 518804
rect 338062 518802 338068 518804
rect 336917 518744 336922 518800
rect 335924 518740 335930 518742
rect 336917 518740 336964 518744
rect 337028 518742 337074 518802
rect 338022 518742 338068 518802
rect 338132 518800 338179 518804
rect 338174 518744 338179 518800
rect 337028 518740 337034 518742
rect 338062 518740 338068 518742
rect 338132 518740 338179 518744
rect 335813 518739 335879 518740
rect 336917 518739 336983 518740
rect 338113 518739 338179 518740
rect 339493 518804 339559 518805
rect 339493 518800 339540 518804
rect 339604 518802 339610 518804
rect 339493 518744 339498 518800
rect 339493 518740 339540 518744
rect 339604 518742 339650 518802
rect 339604 518740 339610 518742
rect 340454 518740 340460 518804
rect 340524 518802 340530 518804
rect 340597 518802 340663 518805
rect 340524 518800 340663 518802
rect 340524 518744 340602 518800
rect 340658 518744 340663 518800
rect 340524 518742 340663 518744
rect 340524 518740 340530 518742
rect 339493 518739 339559 518740
rect 340597 518739 340663 518742
rect 341517 518804 341583 518805
rect 341517 518800 341564 518804
rect 341628 518802 341634 518804
rect 341517 518744 341522 518800
rect 341517 518740 341564 518744
rect 341628 518742 341674 518802
rect 341628 518740 341634 518742
rect 345054 518740 345060 518804
rect 345124 518802 345130 518804
rect 345289 518802 345355 518805
rect 346577 518804 346643 518805
rect 348969 518804 349035 518805
rect 443177 518804 443243 518805
rect 451273 518804 451339 518805
rect 452561 518804 452627 518805
rect 346526 518802 346532 518804
rect 345124 518800 345355 518802
rect 345124 518744 345294 518800
rect 345350 518744 345355 518800
rect 345124 518742 345355 518744
rect 346486 518742 346532 518802
rect 346596 518800 346643 518804
rect 348918 518802 348924 518804
rect 346638 518744 346643 518800
rect 345124 518740 345130 518742
rect 341517 518739 341583 518740
rect 345289 518739 345355 518742
rect 346526 518740 346532 518742
rect 346596 518740 346643 518744
rect 348878 518742 348924 518802
rect 348988 518800 349035 518804
rect 443126 518802 443132 518804
rect 349030 518744 349035 518800
rect 348918 518740 348924 518742
rect 348988 518740 349035 518744
rect 443086 518742 443132 518802
rect 443196 518800 443243 518804
rect 443238 518744 443243 518800
rect 443126 518740 443132 518742
rect 443196 518740 443243 518744
rect 451222 518740 451228 518804
rect 451292 518802 451339 518804
rect 452510 518802 452516 518804
rect 451292 518800 451384 518802
rect 451334 518744 451384 518800
rect 451292 518742 451384 518744
rect 452470 518742 452516 518802
rect 452580 518800 452627 518804
rect 452622 518744 452627 518800
rect 451292 518740 451339 518742
rect 452510 518740 452516 518742
rect 452580 518740 452627 518744
rect 346577 518739 346643 518740
rect 348969 518739 349035 518740
rect 443177 518739 443243 518740
rect 451273 518739 451339 518740
rect 452561 518739 452627 518740
rect 458357 518804 458423 518805
rect 458357 518800 458404 518804
rect 458468 518802 458474 518804
rect 459553 518802 459619 518805
rect 466453 518804 466519 518805
rect 460422 518802 460428 518804
rect 458357 518744 458362 518800
rect 458357 518740 458404 518744
rect 458468 518742 458514 518802
rect 459553 518800 460428 518802
rect 459553 518744 459558 518800
rect 459614 518744 460428 518800
rect 459553 518742 460428 518744
rect 458468 518740 458474 518742
rect 458357 518739 458423 518740
rect 459553 518739 459619 518742
rect 460422 518740 460428 518742
rect 460492 518740 460498 518804
rect 466453 518802 466500 518804
rect 466408 518800 466500 518802
rect 466408 518744 466458 518800
rect 466408 518742 466500 518744
rect 466453 518740 466500 518742
rect 466564 518740 466570 518804
rect 466453 518739 466519 518740
rect 312486 518604 312492 518668
rect 312556 518666 312562 518668
rect 313181 518666 313247 518669
rect 312556 518664 313247 518666
rect 312556 518608 313186 518664
rect 313242 518608 313247 518664
rect 312556 518606 313247 518608
rect 312556 518604 312562 518606
rect 313181 518603 313247 518606
rect 316166 518604 316172 518668
rect 316236 518666 316242 518668
rect 317229 518666 317295 518669
rect 316236 518664 317295 518666
rect 316236 518608 317234 518664
rect 317290 518608 317295 518664
rect 316236 518606 317295 518608
rect 316236 518604 316242 518606
rect 317229 518603 317295 518606
rect 318558 518604 318564 518668
rect 318628 518666 318634 518668
rect 318701 518666 318767 518669
rect 318628 518664 318767 518666
rect 318628 518608 318706 518664
rect 318762 518608 318767 518664
rect 318628 518606 318767 518608
rect 318628 518604 318634 518606
rect 318701 518603 318767 518606
rect 320766 518604 320772 518668
rect 320836 518666 320842 518668
rect 321093 518666 321159 518669
rect 320836 518664 321159 518666
rect 320836 518608 321098 518664
rect 321154 518608 321159 518664
rect 320836 518606 321159 518608
rect 320836 518604 320842 518606
rect 321093 518603 321159 518606
rect 323117 518668 323183 518669
rect 323117 518664 323164 518668
rect 323228 518666 323234 518668
rect 323117 518608 323122 518664
rect 323117 518604 323164 518608
rect 323228 518606 323274 518666
rect 323228 518604 323234 518606
rect 331254 518604 331260 518668
rect 331324 518666 331330 518668
rect 331397 518666 331463 518669
rect 331324 518664 331463 518666
rect 331324 518608 331402 518664
rect 331458 518608 331463 518664
rect 331324 518606 331463 518608
rect 331324 518604 331330 518606
rect 323117 518603 323183 518604
rect 331397 518603 331463 518606
rect 339585 518666 339651 518669
rect 347681 518668 347747 518669
rect 340638 518666 340644 518668
rect 339585 518664 340644 518666
rect 339585 518608 339590 518664
rect 339646 518608 340644 518664
rect 339585 518606 340644 518608
rect 339585 518603 339651 518606
rect 340638 518604 340644 518606
rect 340708 518604 340714 518668
rect 347630 518666 347636 518668
rect 347590 518606 347636 518666
rect 347700 518664 347747 518668
rect 347742 518608 347747 518664
rect 347630 518604 347636 518606
rect 347700 518604 347747 518608
rect 347681 518603 347747 518604
rect 429285 518666 429351 518669
rect 429694 518666 429700 518668
rect 429285 518664 429700 518666
rect 429285 518608 429290 518664
rect 429346 518608 429700 518664
rect 429285 518606 429700 518608
rect 429285 518603 429351 518606
rect 429694 518604 429700 518606
rect 429764 518604 429770 518668
rect 441654 518604 441660 518668
rect 441724 518666 441730 518668
rect 442533 518666 442599 518669
rect 441724 518664 442599 518666
rect 441724 518608 442538 518664
rect 442594 518608 442599 518664
rect 441724 518606 442599 518608
rect 441724 518604 441730 518606
rect 442533 518603 442599 518606
rect 444046 518604 444052 518668
rect 444116 518666 444122 518668
rect 444281 518666 444347 518669
rect 445385 518668 445451 518669
rect 445334 518666 445340 518668
rect 444116 518664 444347 518666
rect 444116 518608 444286 518664
rect 444342 518608 444347 518664
rect 444116 518606 444347 518608
rect 445294 518606 445340 518666
rect 445404 518664 445451 518668
rect 445446 518608 445451 518664
rect 444116 518604 444122 518606
rect 444281 518603 444347 518606
rect 445334 518604 445340 518606
rect 445404 518604 445451 518608
rect 445385 518603 445451 518604
rect 446397 518666 446463 518669
rect 457069 518668 457135 518669
rect 446622 518666 446628 518668
rect 446397 518664 446628 518666
rect 446397 518608 446402 518664
rect 446458 518608 446628 518664
rect 446397 518606 446628 518608
rect 446397 518603 446463 518606
rect 446622 518604 446628 518606
rect 446692 518604 446698 518668
rect 457069 518664 457116 518668
rect 457180 518666 457186 518668
rect 461025 518666 461091 518669
rect 461158 518666 461164 518668
rect 457069 518608 457074 518664
rect 457069 518604 457116 518608
rect 457180 518606 457226 518666
rect 461025 518664 461164 518666
rect 461025 518608 461030 518664
rect 461086 518608 461164 518664
rect 461025 518606 461164 518608
rect 457180 518604 457186 518606
rect 457069 518603 457135 518604
rect 461025 518603 461091 518606
rect 461158 518604 461164 518606
rect 461228 518604 461234 518668
rect 314653 518530 314719 518533
rect 315062 518530 315068 518532
rect 314653 518528 315068 518530
rect 314653 518472 314658 518528
rect 314714 518472 315068 518528
rect 314653 518470 315068 518472
rect 314653 518467 314719 518470
rect 315062 518468 315068 518470
rect 315132 518468 315138 518532
rect 316033 518530 316099 518533
rect 317321 518532 317387 518533
rect 316534 518530 316540 518532
rect 316033 518528 316540 518530
rect 316033 518472 316038 518528
rect 316094 518472 316540 518528
rect 316033 518470 316540 518472
rect 316033 518467 316099 518470
rect 316534 518468 316540 518470
rect 316604 518468 316610 518532
rect 317270 518468 317276 518532
rect 317340 518530 317387 518532
rect 317505 518530 317571 518533
rect 318558 518530 318564 518532
rect 317340 518528 317432 518530
rect 317382 518472 317432 518528
rect 317340 518470 317432 518472
rect 317505 518528 318564 518530
rect 317505 518472 317510 518528
rect 317566 518472 318564 518528
rect 317505 518470 318564 518472
rect 317340 518468 317387 518470
rect 317321 518467 317387 518468
rect 317505 518467 317571 518470
rect 318558 518468 318564 518470
rect 318628 518468 318634 518532
rect 321686 518530 321692 518532
rect 318796 518470 321692 518530
rect 318796 518397 318856 518470
rect 321686 518468 321692 518470
rect 321756 518530 321762 518532
rect 325509 518530 325575 518533
rect 321756 518528 325575 518530
rect 321756 518472 325514 518528
rect 325570 518472 325575 518528
rect 321756 518470 325575 518472
rect 321756 518468 321762 518470
rect 325509 518467 325575 518470
rect 329833 518530 329899 518533
rect 342989 518532 343055 518533
rect 330334 518530 330340 518532
rect 329833 518528 330340 518530
rect 329833 518472 329838 518528
rect 329894 518472 330340 518528
rect 329833 518470 330340 518472
rect 329833 518467 329899 518470
rect 330334 518468 330340 518470
rect 330404 518468 330410 518532
rect 342989 518528 343036 518532
rect 343100 518530 343106 518532
rect 347773 518530 347839 518533
rect 348918 518530 348924 518532
rect 342989 518472 342994 518528
rect 342989 518468 343036 518472
rect 343100 518470 343146 518530
rect 347773 518528 348924 518530
rect 347773 518472 347778 518528
rect 347834 518472 348924 518528
rect 347773 518470 348924 518472
rect 343100 518468 343106 518470
rect 342989 518467 343055 518468
rect 347773 518467 347839 518470
rect 348918 518468 348924 518470
rect 348988 518468 348994 518532
rect 426433 518530 426499 518533
rect 426566 518530 426572 518532
rect 426433 518528 426572 518530
rect 426433 518472 426438 518528
rect 426494 518472 426572 518528
rect 426433 518470 426572 518472
rect 426433 518467 426499 518470
rect 426566 518468 426572 518470
rect 426636 518468 426642 518532
rect 443862 518468 443868 518532
rect 443932 518530 443938 518532
rect 444097 518530 444163 518533
rect 443932 518528 444163 518530
rect 443932 518472 444102 518528
rect 444158 518472 444163 518528
rect 443932 518470 444163 518472
rect 443932 518468 443938 518470
rect 444097 518467 444163 518470
rect 444966 518468 444972 518532
rect 445036 518530 445042 518532
rect 445477 518530 445543 518533
rect 445036 518528 445543 518530
rect 445036 518472 445482 518528
rect 445538 518472 445543 518528
rect 445036 518470 445543 518472
rect 445036 518468 445042 518470
rect 445477 518467 445543 518470
rect 447133 518530 447199 518533
rect 447726 518530 447732 518532
rect 447133 518528 447732 518530
rect 447133 518472 447138 518528
rect 447194 518472 447732 518528
rect 447133 518470 447732 518472
rect 447133 518467 447199 518470
rect 447726 518468 447732 518470
rect 447796 518530 447802 518532
rect 447961 518530 448027 518533
rect 447796 518528 448027 518530
rect 447796 518472 447966 518528
rect 448022 518472 448027 518528
rect 447796 518470 448027 518472
rect 447796 518468 447802 518470
rect 447961 518467 448027 518470
rect 448697 518530 448763 518533
rect 448830 518530 448836 518532
rect 448697 518528 448836 518530
rect 448697 518472 448702 518528
rect 448758 518472 448836 518528
rect 448697 518470 448836 518472
rect 448697 518467 448763 518470
rect 448830 518468 448836 518470
rect 448900 518468 448906 518532
rect 453614 518468 453620 518532
rect 453684 518530 453690 518532
rect 453757 518530 453823 518533
rect 453684 518528 453823 518530
rect 453684 518472 453762 518528
rect 453818 518472 453823 518528
rect 453684 518470 453823 518472
rect 453684 518468 453690 518470
rect 453757 518467 453823 518470
rect 454718 518468 454724 518532
rect 454788 518530 454794 518532
rect 455321 518530 455387 518533
rect 456057 518532 456123 518533
rect 456006 518530 456012 518532
rect 454788 518528 455387 518530
rect 454788 518472 455326 518528
rect 455382 518472 455387 518528
rect 454788 518470 455387 518472
rect 455966 518470 456012 518530
rect 456076 518528 456123 518532
rect 456118 518472 456123 518528
rect 454788 518468 454794 518470
rect 455321 518467 455387 518470
rect 456006 518468 456012 518470
rect 456076 518468 456123 518472
rect 456057 518467 456123 518468
rect 462313 518530 462379 518533
rect 462446 518530 462452 518532
rect 462313 518528 462452 518530
rect 462313 518472 462318 518528
rect 462374 518472 462452 518528
rect 462313 518470 462452 518472
rect 462313 518467 462379 518470
rect 462446 518468 462452 518470
rect 462516 518468 462522 518532
rect 463693 518530 463759 518533
rect 463918 518530 463924 518532
rect 463693 518528 463924 518530
rect 463693 518472 463698 518528
rect 463754 518472 463924 518528
rect 463693 518470 463924 518472
rect 463693 518467 463759 518470
rect 463918 518468 463924 518470
rect 463988 518468 463994 518532
rect 466453 518530 466519 518533
rect 467414 518530 467420 518532
rect 466453 518528 467420 518530
rect 466453 518472 466458 518528
rect 466514 518472 467420 518528
rect 466453 518470 467420 518472
rect 466453 518467 466519 518470
rect 467414 518468 467420 518470
rect 467484 518468 467490 518532
rect 313273 518394 313339 518397
rect 313958 518394 313964 518396
rect 313273 518392 313964 518394
rect 313273 518336 313278 518392
rect 313334 518336 313964 518392
rect 313273 518334 313964 518336
rect 313273 518331 313339 518334
rect 313958 518332 313964 518334
rect 314028 518332 314034 518396
rect 318793 518392 318859 518397
rect 318793 518336 318798 518392
rect 318854 518336 318859 518392
rect 318793 518331 318859 518336
rect 320173 518394 320239 518397
rect 320950 518394 320956 518396
rect 320173 518392 320956 518394
rect 320173 518336 320178 518392
rect 320234 518336 320956 518392
rect 320173 518334 320956 518336
rect 320173 518331 320239 518334
rect 320950 518332 320956 518334
rect 321020 518332 321026 518396
rect 336733 518394 336799 518397
rect 337326 518394 337332 518396
rect 336733 518392 337332 518394
rect 336733 518336 336738 518392
rect 336794 518336 337332 518392
rect 336733 518334 337332 518336
rect 336733 518331 336799 518334
rect 337326 518332 337332 518334
rect 337396 518332 337402 518396
rect 338113 518394 338179 518397
rect 338430 518394 338436 518396
rect 338113 518392 338436 518394
rect 338113 518336 338118 518392
rect 338174 518336 338436 518392
rect 338113 518334 338436 518336
rect 338113 518331 338179 518334
rect 338430 518332 338436 518334
rect 338500 518332 338506 518396
rect 339493 518394 339559 518397
rect 343725 518396 343791 518397
rect 339902 518394 339908 518396
rect 339493 518392 339908 518394
rect 339493 518336 339498 518392
rect 339554 518336 339908 518392
rect 339493 518334 339908 518336
rect 339493 518331 339559 518334
rect 339902 518332 339908 518334
rect 339972 518332 339978 518396
rect 343725 518392 343772 518396
rect 343836 518394 343842 518396
rect 430573 518394 430639 518397
rect 430798 518394 430804 518396
rect 343725 518336 343730 518392
rect 343725 518332 343772 518336
rect 343836 518334 343882 518394
rect 430573 518392 430804 518394
rect 430573 518336 430578 518392
rect 430634 518336 430804 518392
rect 430573 518334 430804 518336
rect 343836 518332 343842 518334
rect 343725 518331 343791 518332
rect 430573 518331 430639 518334
rect 430798 518332 430804 518334
rect 430868 518332 430874 518396
rect 435030 518332 435036 518396
rect 435100 518394 435106 518396
rect 435357 518394 435423 518397
rect 435909 518394 435975 518397
rect 445569 518396 445635 518397
rect 447041 518396 447107 518397
rect 450169 518396 450235 518397
rect 459553 518396 459619 518397
rect 445518 518394 445524 518396
rect 435100 518392 435975 518394
rect 435100 518336 435362 518392
rect 435418 518336 435914 518392
rect 435970 518336 435975 518392
rect 435100 518334 435975 518336
rect 445478 518334 445524 518394
rect 445588 518392 445635 518396
rect 446990 518394 446996 518396
rect 445630 518336 445635 518392
rect 435100 518332 435106 518334
rect 435357 518331 435423 518334
rect 435909 518331 435975 518334
rect 445518 518332 445524 518334
rect 445588 518332 445635 518336
rect 446950 518334 446996 518394
rect 447060 518392 447107 518396
rect 450118 518394 450124 518396
rect 447102 518336 447107 518392
rect 446990 518332 446996 518334
rect 447060 518332 447107 518336
rect 450078 518334 450124 518394
rect 450188 518392 450235 518396
rect 459502 518394 459508 518396
rect 450230 518336 450235 518392
rect 450118 518332 450124 518334
rect 450188 518332 450235 518336
rect 459462 518334 459508 518394
rect 459572 518392 459619 518396
rect 459614 518336 459619 518392
rect 459502 518332 459508 518334
rect 459572 518332 459619 518336
rect 445569 518331 445635 518332
rect 447041 518331 447107 518332
rect 450169 518331 450235 518332
rect 459553 518331 459619 518332
rect 465073 518394 465139 518397
rect 465206 518394 465212 518396
rect 465073 518392 465212 518394
rect 465073 518336 465078 518392
rect 465134 518336 465212 518392
rect 465073 518334 465212 518336
rect 465073 518331 465139 518334
rect 465206 518332 465212 518334
rect 465276 518332 465282 518396
rect 303613 518260 303679 518261
rect 303613 518256 303660 518260
rect 303724 518258 303730 518260
rect 321737 518258 321803 518261
rect 322054 518258 322060 518260
rect 303613 518200 303618 518256
rect 303613 518196 303660 518200
rect 303724 518198 303770 518258
rect 321737 518256 322060 518258
rect 321737 518200 321742 518256
rect 321798 518200 322060 518256
rect 321737 518198 322060 518200
rect 303724 518196 303730 518198
rect 303613 518195 303679 518196
rect 321737 518195 321803 518198
rect 322054 518196 322060 518198
rect 322124 518196 322130 518260
rect 332685 518258 332751 518261
rect 333830 518258 333836 518260
rect 332685 518256 333836 518258
rect 332685 518200 332690 518256
rect 332746 518200 333836 518256
rect 332685 518198 333836 518200
rect 332685 518195 332751 518198
rect 333830 518196 333836 518198
rect 333900 518196 333906 518260
rect 340873 518258 340939 518261
rect 341926 518258 341932 518260
rect 340873 518256 341932 518258
rect 340873 518200 340878 518256
rect 340934 518200 341932 518256
rect 340873 518198 341932 518200
rect 340873 518195 340939 518198
rect 341926 518196 341932 518198
rect 341996 518196 342002 518260
rect 423673 518258 423739 518261
rect 429193 518260 429259 518261
rect 423806 518258 423812 518260
rect 423673 518256 423812 518258
rect 423673 518200 423678 518256
rect 423734 518200 423812 518256
rect 423673 518198 423812 518200
rect 423673 518195 423739 518198
rect 423806 518196 423812 518198
rect 423876 518196 423882 518260
rect 429142 518196 429148 518260
rect 429212 518258 429259 518260
rect 429212 518256 429304 518258
rect 429254 518200 429304 518256
rect 429212 518198 429304 518200
rect 429212 518196 429259 518198
rect 436134 518196 436140 518260
rect 436204 518258 436210 518260
rect 436921 518258 436987 518261
rect 436204 518256 436987 518258
rect 436204 518200 436926 518256
rect 436982 518200 436987 518256
rect 436204 518198 436987 518200
rect 436204 518196 436210 518198
rect 429193 518195 429259 518196
rect 436921 518195 436987 518198
rect 440734 518196 440740 518260
rect 440804 518258 440810 518260
rect 440877 518258 440943 518261
rect 448329 518260 448395 518261
rect 448278 518258 448284 518260
rect 440804 518256 440943 518258
rect 440804 518200 440882 518256
rect 440938 518200 440943 518256
rect 440804 518198 440943 518200
rect 448238 518198 448284 518258
rect 448348 518256 448395 518260
rect 448390 518200 448395 518256
rect 440804 518196 440810 518198
rect 440877 518195 440943 518198
rect 448278 518196 448284 518198
rect 448348 518196 448395 518200
rect 448329 518195 448395 518196
rect 467833 518258 467899 518261
rect 468518 518258 468524 518260
rect 467833 518256 468524 518258
rect 467833 518200 467838 518256
rect 467894 518200 468524 518256
rect 467833 518198 468524 518200
rect 467833 518195 467899 518198
rect 468518 518196 468524 518198
rect 468588 518196 468594 518260
rect 314694 518060 314700 518124
rect 314764 518122 314770 518124
rect 315941 518122 316007 518125
rect 314764 518120 316007 518122
rect 314764 518064 315946 518120
rect 316002 518064 316007 518120
rect 314764 518062 316007 518064
rect 314764 518060 314770 518062
rect 315941 518059 316007 518062
rect 318793 518122 318859 518125
rect 320030 518122 320036 518124
rect 318793 518120 320036 518122
rect 318793 518064 318798 518120
rect 318854 518064 320036 518120
rect 318793 518062 320036 518064
rect 318793 518059 318859 518062
rect 320030 518060 320036 518062
rect 320100 518060 320106 518124
rect 317413 517988 317479 517989
rect 317413 517986 317460 517988
rect 317368 517984 317460 517986
rect 317368 517928 317418 517984
rect 317368 517926 317460 517928
rect 317413 517924 317460 517926
rect 317524 517924 317530 517988
rect 317413 517923 317479 517924
rect 312169 517850 312235 517853
rect 312670 517850 312676 517852
rect 312169 517848 312676 517850
rect 312169 517792 312174 517848
rect 312230 517792 312676 517848
rect 312169 517790 312676 517792
rect 312169 517787 312235 517790
rect 312670 517788 312676 517790
rect 312740 517788 312746 517852
rect 333973 517850 334039 517853
rect 334934 517850 334940 517852
rect 333973 517848 334940 517850
rect 333973 517792 333978 517848
rect 334034 517792 334940 517848
rect 333973 517790 334940 517792
rect 333973 517787 334039 517790
rect 334934 517788 334940 517790
rect 335004 517788 335010 517852
rect 342253 517850 342319 517853
rect 347865 517852 347931 517853
rect 343398 517850 343404 517852
rect 342253 517848 343404 517850
rect 342253 517792 342258 517848
rect 342314 517792 343404 517848
rect 342253 517790 343404 517792
rect 342253 517787 342319 517790
rect 343398 517788 343404 517790
rect 343468 517788 343474 517852
rect 347814 517788 347820 517852
rect 347884 517850 347931 517852
rect 432597 517852 432663 517853
rect 437289 517852 437355 517853
rect 432597 517850 432644 517852
rect 347884 517848 347976 517850
rect 347926 517792 347976 517848
rect 347884 517790 347976 517792
rect 432552 517848 432644 517850
rect 432552 517792 432602 517848
rect 432552 517790 432644 517792
rect 347884 517788 347931 517790
rect 347865 517787 347931 517788
rect 432597 517788 432644 517790
rect 432708 517788 432714 517852
rect 437238 517788 437244 517852
rect 437308 517850 437355 517852
rect 437308 517848 437400 517850
rect 437350 517792 437400 517848
rect 437308 517790 437400 517792
rect 437308 517788 437355 517790
rect 432597 517787 432663 517788
rect 437289 517787 437355 517788
rect 309726 517652 309732 517716
rect 309796 517714 309802 517716
rect 310237 517714 310303 517717
rect 324497 517716 324563 517717
rect 309796 517712 310303 517714
rect 309796 517656 310242 517712
rect 310298 517656 310303 517712
rect 309796 517654 310303 517656
rect 309796 517652 309802 517654
rect 310237 517651 310303 517654
rect 324446 517652 324452 517716
rect 324516 517714 324563 517716
rect 325693 517714 325759 517717
rect 326654 517714 326660 517716
rect 324516 517712 324608 517714
rect 324558 517656 324608 517712
rect 324516 517654 324608 517656
rect 325693 517712 326660 517714
rect 325693 517656 325698 517712
rect 325754 517656 326660 517712
rect 325693 517654 326660 517656
rect 324516 517652 324563 517654
rect 324497 517651 324563 517652
rect 325693 517651 325759 517654
rect 326654 517652 326660 517654
rect 326724 517652 326730 517716
rect 327165 517714 327231 517717
rect 327942 517714 327948 517716
rect 327165 517712 327948 517714
rect 327165 517656 327170 517712
rect 327226 517656 327948 517712
rect 327165 517654 327948 517656
rect 327165 517651 327231 517654
rect 327942 517652 327948 517654
rect 328012 517652 328018 517716
rect 328453 517714 328519 517717
rect 332593 517716 332659 517717
rect 329046 517714 329052 517716
rect 328453 517712 329052 517714
rect 328453 517656 328458 517712
rect 328514 517656 329052 517712
rect 328453 517654 329052 517656
rect 328453 517651 328519 517654
rect 329046 517652 329052 517654
rect 329116 517652 329122 517716
rect 332542 517652 332548 517716
rect 332612 517714 332659 517716
rect 335353 517714 335419 517717
rect 336038 517714 336044 517716
rect 332612 517712 332704 517714
rect 332654 517656 332704 517712
rect 332612 517654 332704 517656
rect 335353 517712 336044 517714
rect 335353 517656 335358 517712
rect 335414 517656 336044 517712
rect 335353 517654 336044 517656
rect 332612 517652 332659 517654
rect 332593 517651 332659 517652
rect 335353 517651 335419 517654
rect 336038 517652 336044 517654
rect 336108 517652 336114 517716
rect 343633 517714 343699 517717
rect 344318 517714 344324 517716
rect 343633 517712 344324 517714
rect 343633 517656 343638 517712
rect 343694 517656 344324 517712
rect 343633 517654 344324 517656
rect 343633 517651 343699 517654
rect 344318 517652 344324 517654
rect 344388 517652 344394 517716
rect 345197 517714 345263 517717
rect 345422 517714 345428 517716
rect 345197 517712 345428 517714
rect 345197 517656 345202 517712
rect 345258 517656 345428 517712
rect 345197 517654 345428 517656
rect 345197 517651 345263 517654
rect 345422 517652 345428 517654
rect 345492 517652 345498 517716
rect 346393 517714 346459 517717
rect 346710 517714 346716 517716
rect 346393 517712 346716 517714
rect 346393 517656 346398 517712
rect 346454 517656 346716 517712
rect 346393 517654 346716 517656
rect 346393 517651 346459 517654
rect 346710 517652 346716 517654
rect 346780 517652 346786 517716
rect 433006 517652 433012 517716
rect 433076 517714 433082 517716
rect 433241 517714 433307 517717
rect 433076 517712 433307 517714
rect 433076 517656 433246 517712
rect 433302 517656 433307 517712
rect 433076 517654 433307 517656
rect 433076 517652 433082 517654
rect 433241 517651 433307 517654
rect 433926 517652 433932 517716
rect 433996 517714 434002 517716
rect 434621 517714 434687 517717
rect 433996 517712 434687 517714
rect 433996 517656 434626 517712
rect 434682 517656 434687 517712
rect 433996 517654 434687 517656
rect 433996 517652 434002 517654
rect 434621 517651 434687 517654
rect 435766 517652 435772 517716
rect 435836 517714 435842 517716
rect 436001 517714 436067 517717
rect 435836 517712 436067 517714
rect 435836 517656 436006 517712
rect 436062 517656 436067 517712
rect 435836 517654 436067 517656
rect 435836 517652 435842 517654
rect 436001 517651 436067 517654
rect 436870 517652 436876 517716
rect 436940 517714 436946 517716
rect 437381 517714 437447 517717
rect 436940 517712 437447 517714
rect 436940 517656 437386 517712
rect 437442 517656 437447 517712
rect 436940 517654 437447 517656
rect 436940 517652 436946 517654
rect 437381 517651 437447 517654
rect 437974 517652 437980 517716
rect 438044 517714 438050 517716
rect 438669 517714 438735 517717
rect 438044 517712 438735 517714
rect 438044 517656 438674 517712
rect 438730 517656 438735 517712
rect 438044 517654 438735 517656
rect 438044 517652 438050 517654
rect 438669 517651 438735 517654
rect 453246 517652 453252 517716
rect 453316 517714 453322 517716
rect 453849 517714 453915 517717
rect 453316 517712 453915 517714
rect 453316 517656 453854 517712
rect 453910 517656 453915 517712
rect 453316 517654 453915 517656
rect 453316 517652 453322 517654
rect 453849 517651 453915 517654
rect 460238 517652 460244 517716
rect 460308 517714 460314 517716
rect 460841 517714 460907 517717
rect 460308 517712 460907 517714
rect 460308 517656 460846 517712
rect 460902 517656 460907 517712
rect 460308 517654 460907 517656
rect 460308 517652 460314 517654
rect 460841 517651 460907 517654
rect 468334 517652 468340 517716
rect 468404 517714 468410 517716
rect 469029 517714 469095 517717
rect 468404 517712 469095 517714
rect 468404 517656 469034 517712
rect 469090 517656 469095 517712
rect 468404 517654 469095 517656
rect 468404 517652 468410 517654
rect 469029 517651 469095 517654
rect 307334 517516 307340 517580
rect 307404 517578 307410 517580
rect 307569 517578 307635 517581
rect 307404 517576 307635 517578
rect 307404 517520 307574 517576
rect 307630 517520 307635 517576
rect 307404 517518 307635 517520
rect 307404 517516 307410 517518
rect 307569 517515 307635 517518
rect 308622 517516 308628 517580
rect 308692 517578 308698 517580
rect 309041 517578 309107 517581
rect 310329 517580 310395 517581
rect 311801 517580 311867 517581
rect 310278 517578 310284 517580
rect 308692 517576 309107 517578
rect 308692 517520 309046 517576
rect 309102 517520 309107 517576
rect 308692 517518 309107 517520
rect 310238 517518 310284 517578
rect 310348 517576 310395 517580
rect 311750 517578 311756 517580
rect 310390 517520 310395 517576
rect 308692 517516 308698 517518
rect 309041 517515 309107 517518
rect 310278 517516 310284 517518
rect 310348 517516 310395 517520
rect 311710 517518 311756 517578
rect 311820 517576 311867 517580
rect 311862 517520 311867 517576
rect 311750 517516 311756 517518
rect 311820 517516 311867 517520
rect 310329 517515 310395 517516
rect 311801 517515 311867 517516
rect 324405 517578 324471 517581
rect 325550 517578 325556 517580
rect 324405 517576 325556 517578
rect 324405 517520 324410 517576
rect 324466 517520 325556 517576
rect 324405 517518 325556 517520
rect 324405 517515 324471 517518
rect 325550 517516 325556 517518
rect 325620 517516 325626 517580
rect 438117 517578 438183 517581
rect 438761 517580 438827 517581
rect 438342 517578 438348 517580
rect 438117 517576 438348 517578
rect 438117 517520 438122 517576
rect 438178 517520 438348 517576
rect 438117 517518 438348 517520
rect 438117 517515 438183 517518
rect 438342 517516 438348 517518
rect 438412 517516 438418 517580
rect 438710 517578 438716 517580
rect 438670 517518 438716 517578
rect 438780 517576 438827 517580
rect 438822 517520 438827 517576
rect 438710 517516 438716 517518
rect 438780 517516 438827 517520
rect 438761 517515 438827 517516
rect 439497 517578 439563 517581
rect 439630 517578 439636 517580
rect 439497 517576 439636 517578
rect 439497 517520 439502 517576
rect 439558 517520 439636 517576
rect 439497 517518 439636 517520
rect 439497 517515 439563 517518
rect 439630 517516 439636 517518
rect 439700 517516 439706 517580
rect 439998 517516 440004 517580
rect 440068 517578 440074 517580
rect 440141 517578 440207 517581
rect 441521 517580 441587 517581
rect 441470 517578 441476 517580
rect 440068 517576 440207 517578
rect 440068 517520 440146 517576
rect 440202 517520 440207 517576
rect 440068 517518 440207 517520
rect 441430 517518 441476 517578
rect 441540 517576 441587 517580
rect 441582 517520 441587 517576
rect 440068 517516 440074 517518
rect 440141 517515 440207 517518
rect 441470 517516 441476 517518
rect 441540 517516 441587 517520
rect 442758 517516 442764 517580
rect 442828 517578 442834 517580
rect 442901 517578 442967 517581
rect 449801 517580 449867 517581
rect 449750 517578 449756 517580
rect 442828 517576 442967 517578
rect 442828 517520 442906 517576
rect 442962 517520 442967 517576
rect 442828 517518 442967 517520
rect 449710 517518 449756 517578
rect 449820 517576 449867 517580
rect 449862 517520 449867 517576
rect 442828 517516 442834 517518
rect 441521 517515 441587 517516
rect 442901 517515 442967 517518
rect 449750 517516 449756 517518
rect 449820 517516 449867 517520
rect 450854 517516 450860 517580
rect 450924 517578 450930 517580
rect 451181 517578 451247 517581
rect 450924 517576 451247 517578
rect 450924 517520 451186 517576
rect 451242 517520 451247 517576
rect 450924 517518 451247 517520
rect 450924 517516 450930 517518
rect 449801 517515 449867 517516
rect 451181 517515 451247 517518
rect 451958 517516 451964 517580
rect 452028 517578 452034 517580
rect 452561 517578 452627 517581
rect 452028 517576 452627 517578
rect 452028 517520 452566 517576
rect 452622 517520 452627 517576
rect 452028 517518 452627 517520
rect 452028 517516 452034 517518
rect 452561 517515 452627 517518
rect 453798 517516 453804 517580
rect 453868 517578 453874 517580
rect 453941 517578 454007 517581
rect 455321 517580 455387 517581
rect 455270 517578 455276 517580
rect 453868 517576 454007 517578
rect 453868 517520 453946 517576
rect 454002 517520 454007 517576
rect 453868 517518 454007 517520
rect 455230 517518 455276 517578
rect 455340 517576 455387 517580
rect 455382 517520 455387 517576
rect 453868 517516 453874 517518
rect 453941 517515 454007 517518
rect 455270 517516 455276 517518
rect 455340 517516 455387 517520
rect 456374 517516 456380 517580
rect 456444 517578 456450 517580
rect 456701 517578 456767 517581
rect 456444 517576 456767 517578
rect 456444 517520 456706 517576
rect 456762 517520 456767 517576
rect 456444 517518 456767 517520
rect 456444 517516 456450 517518
rect 455321 517515 455387 517516
rect 456701 517515 456767 517518
rect 457846 517516 457852 517580
rect 457916 517578 457922 517580
rect 458081 517578 458147 517581
rect 457916 517576 458147 517578
rect 457916 517520 458086 517576
rect 458142 517520 458147 517576
rect 457916 517518 458147 517520
rect 457916 517516 457922 517518
rect 458081 517515 458147 517518
rect 459134 517516 459140 517580
rect 459204 517578 459210 517580
rect 459461 517578 459527 517581
rect 460749 517580 460815 517581
rect 460749 517578 460796 517580
rect 459204 517576 459527 517578
rect 459204 517520 459466 517576
rect 459522 517520 459527 517576
rect 459204 517518 459527 517520
rect 460704 517576 460796 517578
rect 460704 517520 460754 517576
rect 460704 517518 460796 517520
rect 459204 517516 459210 517518
rect 459461 517515 459527 517518
rect 460749 517516 460796 517518
rect 460860 517516 460866 517580
rect 462078 517516 462084 517580
rect 462148 517578 462154 517580
rect 462221 517578 462287 517581
rect 463601 517580 463667 517581
rect 463550 517578 463556 517580
rect 462148 517576 462287 517578
rect 462148 517520 462226 517576
rect 462282 517520 462287 517576
rect 462148 517518 462287 517520
rect 463510 517518 463556 517578
rect 463620 517576 463667 517580
rect 463662 517520 463667 517576
rect 462148 517516 462154 517518
rect 460749 517515 460815 517516
rect 462221 517515 462287 517518
rect 463550 517516 463556 517518
rect 463620 517516 463667 517520
rect 464838 517516 464844 517580
rect 464908 517578 464914 517580
rect 464981 517578 465047 517581
rect 464908 517576 465047 517578
rect 464908 517520 464986 517576
rect 465042 517520 465047 517576
rect 464908 517518 465047 517520
rect 464908 517516 464914 517518
rect 463601 517515 463667 517516
rect 464981 517515 465047 517518
rect 466126 517516 466132 517580
rect 466196 517578 466202 517580
rect 466361 517578 466427 517581
rect 466196 517576 466427 517578
rect 466196 517520 466366 517576
rect 466422 517520 466427 517576
rect 466196 517518 466427 517520
rect 466196 517516 466202 517518
rect 466361 517515 466427 517518
rect 467230 517516 467236 517580
rect 467300 517578 467306 517580
rect 467741 517578 467807 517581
rect 469121 517580 469187 517581
rect 469070 517578 469076 517580
rect 467300 517576 467807 517578
rect 467300 517520 467746 517576
rect 467802 517520 467807 517576
rect 467300 517518 467807 517520
rect 469030 517518 469076 517578
rect 469140 517576 469187 517580
rect 469182 517520 469187 517576
rect 467300 517516 467306 517518
rect 467741 517515 467807 517518
rect 469070 517516 469076 517518
rect 469140 517516 469187 517520
rect 469121 517515 469187 517516
rect 543273 512002 543339 512005
rect 543457 512002 543523 512005
rect 543273 512000 543523 512002
rect 543273 511944 543278 512000
rect 543334 511944 543462 512000
rect 543518 511944 543523 512000
rect 543273 511942 543523 511944
rect 543273 511939 543339 511942
rect 543457 511939 543523 511942
rect 580165 510370 580231 510373
rect 583520 510370 584960 510460
rect 580165 510368 584960 510370
rect 580165 510312 580170 510368
rect 580226 510312 584960 510368
rect 580165 510310 584960 510312
rect 580165 510307 580231 510310
rect 583520 510220 584960 510310
rect -960 509962 480 510052
rect 3233 509962 3299 509965
rect -960 509960 3299 509962
rect -960 509904 3238 509960
rect 3294 509904 3299 509960
rect -960 509902 3299 509904
rect -960 509812 480 509902
rect 3233 509899 3299 509902
rect 580165 498674 580231 498677
rect 583520 498674 584960 498764
rect 580165 498672 584960 498674
rect 580165 498616 580170 498672
rect 580226 498616 584960 498672
rect 580165 498614 584960 498616
rect 580165 498611 580231 498614
rect 583520 498524 584960 498614
rect -960 495546 480 495636
rect 3325 495546 3391 495549
rect -960 495544 3391 495546
rect -960 495488 3330 495544
rect 3386 495488 3391 495544
rect -960 495486 3391 495488
rect -960 495396 480 495486
rect 3325 495483 3391 495486
rect 433926 495484 433932 495548
rect 433996 495546 434002 495548
rect 434069 495546 434135 495549
rect 433996 495544 434135 495546
rect 433996 495488 434074 495544
rect 434130 495488 434135 495544
rect 433996 495486 434135 495488
rect 433996 495484 434002 495486
rect 434069 495483 434135 495486
rect 433885 492692 433951 492693
rect 433885 492688 433932 492692
rect 433996 492690 434002 492692
rect 433885 492632 433890 492688
rect 433885 492628 433932 492632
rect 433996 492630 434042 492690
rect 433996 492628 434002 492630
rect 433885 492627 433951 492628
rect 580165 486842 580231 486845
rect 583520 486842 584960 486932
rect 580165 486840 584960 486842
rect 580165 486784 580170 486840
rect 580226 486784 584960 486840
rect 580165 486782 584960 486784
rect 580165 486779 580231 486782
rect 583520 486692 584960 486782
rect 433609 483034 433675 483037
rect 433793 483034 433859 483037
rect 433609 483032 433859 483034
rect 433609 482976 433614 483032
rect 433670 482976 433798 483032
rect 433854 482976 433859 483032
rect 433609 482974 433859 482976
rect 433609 482971 433675 482974
rect 433793 482971 433859 482974
rect 543273 483034 543339 483037
rect 543457 483034 543523 483037
rect 543273 483032 543523 483034
rect 543273 482976 543278 483032
rect 543334 482976 543462 483032
rect 543518 482976 543523 483032
rect 543273 482974 543523 482976
rect 543273 482971 543339 482974
rect 543457 482971 543523 482974
rect 466361 482490 466427 482493
rect 530853 482490 530919 482493
rect 466361 482488 530919 482490
rect 466361 482432 466366 482488
rect 466422 482432 530858 482488
rect 530914 482432 530919 482488
rect 466361 482430 530919 482432
rect 466361 482427 466427 482430
rect 530853 482427 530919 482430
rect 469029 482354 469095 482357
rect 536005 482354 536071 482357
rect 469029 482352 536071 482354
rect 469029 482296 469034 482352
rect 469090 482296 536010 482352
rect 536066 482296 536071 482352
rect 469029 482294 536071 482296
rect 469029 482291 469095 482294
rect 536005 482291 536071 482294
rect 263685 482218 263751 482221
rect 379697 482218 379763 482221
rect 263685 482216 379763 482218
rect 263685 482160 263690 482216
rect 263746 482160 379702 482216
rect 379758 482160 379763 482216
rect 263685 482158 379763 482160
rect 263685 482155 263751 482158
rect 379697 482155 379763 482158
rect 469121 482218 469187 482221
rect 538581 482218 538647 482221
rect 469121 482216 538647 482218
rect 469121 482160 469126 482216
rect 469182 482160 538586 482216
rect 538642 482160 538647 482216
rect 469121 482158 538647 482160
rect 469121 482155 469187 482158
rect 538581 482155 538647 482158
rect 320173 482082 320239 482085
rect 321553 482082 321619 482085
rect 320173 482080 321619 482082
rect 320173 482024 320178 482080
rect 320234 482024 321558 482080
rect 321614 482024 321619 482080
rect 320173 482022 321619 482024
rect 320173 482019 320239 482022
rect 321553 482019 321619 482022
rect 471237 481810 471303 481813
rect 477217 481810 477283 481813
rect 471237 481808 477283 481810
rect 471237 481752 471242 481808
rect 471298 481752 477222 481808
rect 477278 481752 477283 481808
rect 471237 481750 477283 481752
rect 471237 481747 471303 481750
rect 477217 481747 477283 481750
rect -960 481130 480 481220
rect 3141 481130 3207 481133
rect -960 481128 3207 481130
rect -960 481072 3146 481128
rect 3202 481072 3207 481128
rect -960 481070 3207 481072
rect -960 480980 480 481070
rect 3141 481067 3207 481070
rect 256693 478954 256759 478957
rect 542486 478954 542492 478956
rect 256693 478952 260084 478954
rect 256693 478896 256698 478952
rect 256754 478896 260084 478952
rect 256693 478894 260084 478896
rect 539948 478894 542492 478954
rect 256693 478891 256759 478894
rect 542486 478892 542492 478894
rect 542556 478892 542562 478956
rect 542302 476914 542308 476916
rect 539948 476854 542308 476914
rect 542302 476852 542308 476854
rect 542372 476852 542378 476916
rect 256693 476778 256759 476781
rect 256693 476776 260084 476778
rect 256693 476720 256698 476776
rect 256754 476720 260084 476776
rect 256693 476718 260084 476720
rect 256693 476715 256759 476718
rect 583520 474996 584960 475236
rect 256693 474738 256759 474741
rect 542670 474738 542676 474740
rect 256693 474736 260084 474738
rect 256693 474680 256698 474736
rect 256754 474680 260084 474736
rect 256693 474678 260084 474680
rect 539948 474678 542676 474738
rect 256693 474675 256759 474678
rect 542670 474676 542676 474678
rect 542740 474676 542746 474740
rect 541566 472698 541572 472700
rect 539948 472638 541572 472698
rect 541566 472636 541572 472638
rect 541636 472636 541642 472700
rect 256693 472562 256759 472565
rect 256693 472560 260084 472562
rect 256693 472504 256698 472560
rect 256754 472504 260084 472560
rect 256693 472502 260084 472504
rect 256693 472499 256759 472502
rect 256693 470386 256759 470389
rect 256693 470384 260084 470386
rect 256693 470328 256698 470384
rect 256754 470328 260084 470384
rect 256693 470326 260084 470328
rect 256693 470323 256759 470326
rect 539550 469980 539610 470492
rect 539542 469916 539548 469980
rect 539612 469916 539618 469980
rect 542854 468482 542860 468484
rect 539948 468422 542860 468482
rect 542854 468420 542860 468422
rect 542924 468420 542930 468484
rect 256693 468346 256759 468349
rect 256693 468344 260084 468346
rect 256693 468288 256698 468344
rect 256754 468288 260084 468344
rect 256693 468286 260084 468288
rect 256693 468283 256759 468286
rect -960 466700 480 466940
rect 542261 466306 542327 466309
rect 539948 466304 542327 466306
rect 539948 466248 542266 466304
rect 542322 466248 542327 466304
rect 539948 466246 542327 466248
rect 542261 466243 542327 466246
rect 256693 466170 256759 466173
rect 256693 466168 260084 466170
rect 256693 466112 256698 466168
rect 256754 466112 260084 466168
rect 256693 466110 260084 466112
rect 256693 466107 256759 466110
rect 256693 464130 256759 464133
rect 256693 464128 260084 464130
rect 256693 464072 256698 464128
rect 256754 464072 260084 464128
rect 256693 464070 260084 464072
rect 256693 464067 256759 464070
rect 539734 463724 539794 464236
rect 539726 463660 539732 463724
rect 539796 463660 539802 463724
rect 580165 463450 580231 463453
rect 583520 463450 584960 463540
rect 580165 463448 584960 463450
rect 580165 463392 580170 463448
rect 580226 463392 584960 463448
rect 580165 463390 584960 463392
rect 580165 463387 580231 463390
rect 583520 463300 584960 463390
rect 540278 462090 540284 462092
rect 539948 462030 540284 462090
rect 540278 462028 540284 462030
rect 540348 462028 540354 462092
rect 256693 461954 256759 461957
rect 256693 461952 260084 461954
rect 256693 461896 256698 461952
rect 256754 461896 260084 461952
rect 256693 461894 260084 461896
rect 256693 461891 256759 461894
rect 543038 460050 543044 460052
rect 539948 459990 543044 460050
rect 543038 459988 543044 459990
rect 543108 459988 543114 460052
rect 256693 459778 256759 459781
rect 256693 459776 260084 459778
rect 256693 459720 256698 459776
rect 256754 459720 260084 459776
rect 256693 459718 260084 459720
rect 256693 459715 256759 459718
rect 543222 457874 543228 457876
rect 539948 457814 543228 457874
rect 543222 457812 543228 457814
rect 543292 457812 543298 457876
rect 256693 457738 256759 457741
rect 256693 457736 260084 457738
rect 256693 457680 256698 457736
rect 256754 457680 260084 457736
rect 256693 457678 260084 457680
rect 256693 457675 256759 457678
rect 256693 455562 256759 455565
rect 256693 455560 260084 455562
rect 256693 455504 256698 455560
rect 256754 455504 260084 455560
rect 256693 455502 260084 455504
rect 256693 455499 256759 455502
rect 539366 455292 539426 455804
rect 539358 455228 539364 455292
rect 539428 455228 539434 455292
rect 543641 453658 543707 453661
rect 539948 453656 543707 453658
rect 539948 453600 543646 453656
rect 543702 453600 543707 453656
rect 539948 453598 543707 453600
rect 543641 453595 543707 453598
rect 256693 453386 256759 453389
rect 256693 453384 260084 453386
rect 256693 453328 256698 453384
rect 256754 453328 260084 453384
rect 256693 453326 260084 453328
rect 256693 453323 256759 453326
rect -960 452434 480 452524
rect 3417 452434 3483 452437
rect -960 452432 3483 452434
rect -960 452376 3422 452432
rect 3478 452376 3483 452432
rect -960 452374 3483 452376
rect -960 452284 480 452374
rect 3417 452371 3483 452374
rect 539726 451964 539732 452028
rect 539796 452026 539802 452028
rect 540462 452026 540468 452028
rect 539796 451966 540468 452026
rect 539796 451964 539802 451966
rect 540462 451964 540468 451966
rect 540532 451964 540538 452028
rect 580165 451754 580231 451757
rect 583520 451754 584960 451844
rect 580165 451752 584960 451754
rect 580165 451696 580170 451752
rect 580226 451696 584960 451752
rect 580165 451694 584960 451696
rect 580165 451691 580231 451694
rect 542537 451618 542603 451621
rect 539948 451616 542603 451618
rect 539948 451560 542542 451616
rect 542598 451560 542603 451616
rect 583520 451604 584960 451694
rect 539948 451558 542603 451560
rect 542537 451555 542603 451558
rect 256693 451346 256759 451349
rect 256693 451344 260084 451346
rect 256693 451288 256698 451344
rect 256754 451288 260084 451344
rect 256693 451286 260084 451288
rect 256693 451283 256759 451286
rect 539358 451148 539364 451212
rect 539428 451210 539434 451212
rect 539726 451210 539732 451212
rect 539428 451150 539732 451210
rect 539428 451148 539434 451150
rect 539726 451148 539732 451150
rect 539796 451148 539802 451212
rect 541617 449442 541683 449445
rect 539948 449440 541683 449442
rect 539948 449384 541622 449440
rect 541678 449384 541683 449440
rect 539948 449382 541683 449384
rect 541617 449379 541683 449382
rect 256693 449170 256759 449173
rect 256693 449168 260084 449170
rect 256693 449112 256698 449168
rect 256754 449112 260084 449168
rect 256693 449110 260084 449112
rect 256693 449107 256759 449110
rect 540421 447402 540487 447405
rect 539948 447400 540487 447402
rect 539948 447344 540426 447400
rect 540482 447344 540487 447400
rect 539948 447342 540487 447344
rect 540421 447339 540487 447342
rect 256693 447130 256759 447133
rect 256693 447128 260084 447130
rect 256693 447072 256698 447128
rect 256754 447072 260084 447128
rect 256693 447070 260084 447072
rect 256693 447067 256759 447070
rect 542353 445226 542419 445229
rect 539948 445224 542419 445226
rect 539948 445168 542358 445224
rect 542414 445168 542419 445224
rect 539948 445166 542419 445168
rect 542353 445163 542419 445166
rect 256693 444954 256759 444957
rect 256693 444952 260084 444954
rect 256693 444896 256698 444952
rect 256754 444896 260084 444952
rect 256693 444894 260084 444896
rect 256693 444891 256759 444894
rect 256693 442778 256759 442781
rect 256693 442776 260084 442778
rect 256693 442720 256698 442776
rect 256754 442720 260084 442776
rect 256693 442718 260084 442720
rect 256693 442715 256759 442718
rect 539366 442644 539426 443156
rect 539358 442580 539364 442644
rect 539428 442580 539434 442644
rect 539726 442506 539732 442508
rect 539550 442446 539732 442506
rect 539358 442172 539364 442236
rect 539428 442234 539434 442236
rect 539550 442234 539610 442446
rect 539726 442444 539732 442446
rect 539796 442444 539802 442508
rect 539726 442308 539732 442372
rect 539796 442370 539802 442372
rect 540462 442370 540468 442372
rect 539796 442310 540468 442370
rect 539796 442308 539802 442310
rect 540462 442308 540468 442310
rect 540532 442308 540538 442372
rect 539428 442174 539610 442234
rect 539428 442172 539434 442174
rect 542445 441010 542511 441013
rect 539948 441008 542511 441010
rect 539948 440952 542450 441008
rect 542506 440952 542511 441008
rect 539948 440950 542511 440952
rect 542445 440947 542511 440950
rect 256693 440738 256759 440741
rect 256693 440736 260084 440738
rect 256693 440680 256698 440736
rect 256754 440680 260084 440736
rect 256693 440678 260084 440680
rect 256693 440675 256759 440678
rect 580165 439922 580231 439925
rect 583520 439922 584960 440012
rect 580165 439920 584960 439922
rect 580165 439864 580170 439920
rect 580226 439864 584960 439920
rect 580165 439862 584960 439864
rect 580165 439859 580231 439862
rect 583520 439772 584960 439862
rect 542445 438970 542511 438973
rect 539948 438968 542511 438970
rect 539948 438912 542450 438968
rect 542506 438912 542511 438968
rect 539948 438910 542511 438912
rect 542445 438907 542511 438910
rect 256693 438562 256759 438565
rect 256693 438560 260084 438562
rect 256693 438504 256698 438560
rect 256754 438504 260084 438560
rect 256693 438502 260084 438504
rect 256693 438499 256759 438502
rect -960 438018 480 438108
rect 3141 438018 3207 438021
rect -960 438016 3207 438018
rect -960 437960 3146 438016
rect 3202 437960 3207 438016
rect -960 437958 3207 437960
rect -960 437868 480 437958
rect 3141 437955 3207 437958
rect 543273 436794 543339 436797
rect 539948 436792 543339 436794
rect 539948 436736 543278 436792
rect 543334 436736 543339 436792
rect 539948 436734 543339 436736
rect 543273 436731 543339 436734
rect 256693 436386 256759 436389
rect 256693 436384 260084 436386
rect 256693 436328 256698 436384
rect 256754 436328 260084 436384
rect 256693 436326 260084 436328
rect 256693 436323 256759 436326
rect 543457 434754 543523 434757
rect 539948 434752 543523 434754
rect 539948 434696 543462 434752
rect 543518 434696 543523 434752
rect 539948 434694 543523 434696
rect 543457 434691 543523 434694
rect 256693 434346 256759 434349
rect 256693 434344 260084 434346
rect 256693 434288 256698 434344
rect 256754 434288 260084 434344
rect 256693 434286 260084 434288
rect 256693 434283 256759 434286
rect 539726 432652 539732 432716
rect 539796 432714 539802 432716
rect 540462 432714 540468 432716
rect 539796 432654 540468 432714
rect 539796 432652 539802 432654
rect 540462 432652 540468 432654
rect 540532 432652 540538 432716
rect 543549 432578 543615 432581
rect 539948 432576 543615 432578
rect 539948 432520 543554 432576
rect 543610 432520 543615 432576
rect 539948 432518 543615 432520
rect 543549 432515 543615 432518
rect 256693 432170 256759 432173
rect 256693 432168 260084 432170
rect 256693 432112 256698 432168
rect 256754 432112 260084 432168
rect 256693 432110 260084 432112
rect 256693 432107 256759 432110
rect 542629 430538 542695 430541
rect 539948 430536 542695 430538
rect 539948 430480 542634 430536
rect 542690 430480 542695 430536
rect 539948 430478 542695 430480
rect 542629 430475 542695 430478
rect 256693 430130 256759 430133
rect 256693 430128 260084 430130
rect 256693 430072 256698 430128
rect 256754 430072 260084 430128
rect 256693 430070 260084 430072
rect 256693 430067 256759 430070
rect 540881 428362 540947 428365
rect 539948 428360 540947 428362
rect 539948 428304 540886 428360
rect 540942 428304 540947 428360
rect 539948 428302 540947 428304
rect 540881 428299 540947 428302
rect 583520 428076 584960 428316
rect 256693 427954 256759 427957
rect 256693 427952 260084 427954
rect 256693 427896 256698 427952
rect 256754 427896 260084 427952
rect 256693 427894 260084 427896
rect 256693 427891 256759 427894
rect 540789 426322 540855 426325
rect 539948 426320 540855 426322
rect 539948 426264 540794 426320
rect 540850 426264 540855 426320
rect 539948 426262 540855 426264
rect 540789 426259 540855 426262
rect 256693 425778 256759 425781
rect 256693 425776 260084 425778
rect 256693 425720 256698 425776
rect 256754 425720 260084 425776
rect 256693 425718 260084 425720
rect 256693 425715 256759 425718
rect 542721 424146 542787 424149
rect 539948 424144 542787 424146
rect 539948 424088 542726 424144
rect 542782 424088 542787 424144
rect 539948 424086 542787 424088
rect 542721 424083 542787 424086
rect -960 423738 480 423828
rect 3233 423738 3299 423741
rect -960 423736 3299 423738
rect -960 423680 3238 423736
rect 3294 423680 3299 423736
rect -960 423678 3299 423680
rect -960 423588 480 423678
rect 3233 423675 3299 423678
rect 256693 423738 256759 423741
rect 256693 423736 260084 423738
rect 256693 423680 256698 423736
rect 256754 423680 260084 423736
rect 256693 423678 260084 423680
rect 256693 423675 256759 423678
rect 543181 422106 543247 422109
rect 539948 422104 543247 422106
rect 539948 422048 543186 422104
rect 543242 422048 543247 422104
rect 539948 422046 543247 422048
rect 543181 422043 543247 422046
rect 256693 421562 256759 421565
rect 256693 421560 260084 421562
rect 256693 421504 256698 421560
rect 256754 421504 260084 421560
rect 256693 421502 260084 421504
rect 256693 421499 256759 421502
rect 543089 420066 543155 420069
rect 539948 420064 543155 420066
rect 539948 420008 543094 420064
rect 543150 420008 543155 420064
rect 539948 420006 543155 420008
rect 543089 420003 543155 420006
rect 256693 419522 256759 419525
rect 256693 419520 260084 419522
rect 256693 419464 256698 419520
rect 256754 419464 260084 419520
rect 256693 419462 260084 419464
rect 256693 419459 256759 419462
rect 539542 418372 539548 418436
rect 539612 418434 539618 418436
rect 540789 418434 540855 418437
rect 539612 418432 540855 418434
rect 539612 418376 540794 418432
rect 540850 418376 540855 418432
rect 539612 418374 540855 418376
rect 539612 418372 539618 418374
rect 540789 418371 540855 418374
rect 540697 417890 540763 417893
rect 539948 417888 540763 417890
rect 539948 417832 540702 417888
rect 540758 417832 540763 417888
rect 539948 417830 540763 417832
rect 540697 417827 540763 417830
rect 256693 417346 256759 417349
rect 256693 417344 260084 417346
rect 256693 417288 256698 417344
rect 256754 417288 260084 417344
rect 256693 417286 260084 417288
rect 256693 417283 256759 417286
rect 580165 416530 580231 416533
rect 583520 416530 584960 416620
rect 580165 416528 584960 416530
rect 580165 416472 580170 416528
rect 580226 416472 584960 416528
rect 580165 416470 584960 416472
rect 580165 416467 580231 416470
rect 583520 416380 584960 416470
rect 540973 415850 541039 415853
rect 539948 415848 541039 415850
rect 539948 415792 540978 415848
rect 541034 415792 541039 415848
rect 539948 415790 541039 415792
rect 540973 415787 541039 415790
rect 256693 415170 256759 415173
rect 256693 415168 260084 415170
rect 256693 415112 256698 415168
rect 256754 415112 260084 415168
rect 256693 415110 260084 415112
rect 256693 415107 256759 415110
rect 539358 414972 539364 415036
rect 539428 415034 539434 415036
rect 539428 414974 539978 415034
rect 539428 414972 539434 414974
rect 539358 414428 539364 414492
rect 539428 414490 539434 414492
rect 539726 414490 539732 414492
rect 539428 414430 539732 414490
rect 539428 414428 539434 414430
rect 539726 414428 539732 414430
rect 539796 414428 539802 414492
rect 539358 413748 539364 413812
rect 539428 413810 539434 413812
rect 539918 413810 539978 414974
rect 539428 413750 539978 413810
rect 539428 413748 539434 413750
rect 540605 413674 540671 413677
rect 539948 413672 540671 413674
rect 539948 413616 540610 413672
rect 540666 413616 540671 413672
rect 539948 413614 540671 413616
rect 540605 413611 540671 413614
rect 539726 413340 539732 413404
rect 539796 413402 539802 413404
rect 540462 413402 540468 413404
rect 539796 413342 540468 413402
rect 539796 413340 539802 413342
rect 540462 413340 540468 413342
rect 540532 413340 540538 413404
rect 256693 413130 256759 413133
rect 256693 413128 260084 413130
rect 256693 413072 256698 413128
rect 256754 413072 260084 413128
rect 256693 413070 260084 413072
rect 256693 413067 256759 413070
rect 539501 412178 539567 412181
rect 539501 412176 539610 412178
rect 539501 412120 539506 412176
rect 539562 412120 539610 412176
rect 539501 412115 539610 412120
rect 539550 411604 539610 412115
rect 256693 410954 256759 410957
rect 256693 410952 260084 410954
rect 256693 410896 256698 410952
rect 256754 410896 260084 410952
rect 256693 410894 260084 410896
rect 256693 410891 256759 410894
rect 542997 409458 543063 409461
rect 539948 409456 543063 409458
rect -960 409172 480 409412
rect 539948 409400 543002 409456
rect 543058 409400 543063 409456
rect 539948 409398 543063 409400
rect 542997 409395 543063 409398
rect 256693 408778 256759 408781
rect 256693 408776 260084 408778
rect 256693 408720 256698 408776
rect 256754 408720 260084 408776
rect 256693 408718 260084 408720
rect 256693 408715 256759 408718
rect 542905 407418 542971 407421
rect 539948 407416 542971 407418
rect 539948 407360 542910 407416
rect 542966 407360 542971 407416
rect 539948 407358 542971 407360
rect 542905 407355 542971 407358
rect 256693 406738 256759 406741
rect 256693 406736 260084 406738
rect 256693 406680 256698 406736
rect 256754 406680 260084 406736
rect 256693 406678 260084 406680
rect 256693 406675 256759 406678
rect 539501 406468 539567 406469
rect 539501 406466 539548 406468
rect 539456 406464 539548 406466
rect 539456 406408 539506 406464
rect 539456 406406 539548 406408
rect 539501 406404 539548 406406
rect 539612 406404 539618 406468
rect 539501 406403 539567 406404
rect 539358 405724 539364 405788
rect 539428 405786 539434 405788
rect 539501 405786 539567 405789
rect 539428 405784 539567 405786
rect 539428 405728 539506 405784
rect 539562 405728 539567 405784
rect 539428 405726 539567 405728
rect 539428 405724 539434 405726
rect 539501 405723 539567 405726
rect 540513 405242 540579 405245
rect 539948 405240 540579 405242
rect 539948 405184 540518 405240
rect 540574 405184 540579 405240
rect 539948 405182 540579 405184
rect 540513 405179 540579 405182
rect 580165 404834 580231 404837
rect 583520 404834 584960 404924
rect 580165 404832 584960 404834
rect 580165 404776 580170 404832
rect 580226 404776 584960 404832
rect 580165 404774 584960 404776
rect 580165 404771 580231 404774
rect 583520 404684 584960 404774
rect 256693 404562 256759 404565
rect 256693 404560 260084 404562
rect 256693 404504 256698 404560
rect 256754 404504 260084 404560
rect 256693 404502 260084 404504
rect 256693 404499 256759 404502
rect 539726 403684 539732 403748
rect 539796 403746 539802 403748
rect 540462 403746 540468 403748
rect 539796 403686 540468 403746
rect 539796 403684 539802 403686
rect 540462 403684 540468 403686
rect 540532 403684 540538 403748
rect 541709 403202 541775 403205
rect 539948 403200 541775 403202
rect 539948 403144 541714 403200
rect 541770 403144 541775 403200
rect 539948 403142 541775 403144
rect 541709 403139 541775 403142
rect 256693 402522 256759 402525
rect 256693 402520 260084 402522
rect 256693 402464 256698 402520
rect 256754 402464 260084 402520
rect 256693 402462 260084 402464
rect 256693 402459 256759 402462
rect 539358 402188 539364 402252
rect 539428 402250 539434 402252
rect 539501 402250 539567 402253
rect 539428 402248 539567 402250
rect 539428 402192 539506 402248
rect 539562 402192 539567 402248
rect 539428 402190 539567 402192
rect 539428 402188 539434 402190
rect 539501 402187 539567 402190
rect 542813 401026 542879 401029
rect 539948 401024 542879 401026
rect 539948 400968 542818 401024
rect 542874 400968 542879 401024
rect 539948 400966 542879 400968
rect 542813 400963 542879 400966
rect 256693 400346 256759 400349
rect 256693 400344 260084 400346
rect 256693 400288 256698 400344
rect 256754 400288 260084 400344
rect 256693 400286 260084 400288
rect 256693 400283 256759 400286
rect 543457 399532 543523 399533
rect 539358 399468 539364 399532
rect 539428 399468 539434 399532
rect 543406 399530 543412 399532
rect 543366 399470 543412 399530
rect 543476 399528 543523 399532
rect 543518 399472 543523 399528
rect 543406 399468 543412 399470
rect 543476 399468 543523 399472
rect 539366 398956 539426 399468
rect 543457 399467 543523 399468
rect 539542 399060 539548 399124
rect 539612 399122 539618 399124
rect 540605 399122 540671 399125
rect 539612 399120 540671 399122
rect 539612 399064 540610 399120
rect 540666 399064 540671 399120
rect 539612 399062 540671 399064
rect 539612 399060 539618 399062
rect 540605 399059 540671 399062
rect 539542 398516 539548 398580
rect 539612 398578 539618 398580
rect 540513 398578 540579 398581
rect 539612 398576 540579 398578
rect 539612 398520 540518 398576
rect 540574 398520 540579 398576
rect 539612 398518 540579 398520
rect 539612 398516 539618 398518
rect 540513 398515 540579 398518
rect 256693 398170 256759 398173
rect 256693 398168 260084 398170
rect 256693 398112 256698 398168
rect 256754 398112 260084 398168
rect 256693 398110 260084 398112
rect 256693 398107 256759 398110
rect 541249 396810 541315 396813
rect 539948 396808 541315 396810
rect 539948 396752 541254 396808
rect 541310 396752 541315 396808
rect 539948 396750 541315 396752
rect 541249 396747 541315 396750
rect 256693 396130 256759 396133
rect 256693 396128 260084 396130
rect 256693 396072 256698 396128
rect 256754 396072 260084 396128
rect 256693 396070 260084 396072
rect 256693 396067 256759 396070
rect 539358 395388 539364 395452
rect 539428 395450 539434 395452
rect 540605 395450 540671 395453
rect 539428 395448 540671 395450
rect 539428 395392 540610 395448
rect 540666 395392 540671 395448
rect 539428 395390 540671 395392
rect 539428 395388 539434 395390
rect 540605 395387 540671 395390
rect -960 395042 480 395132
rect 3141 395042 3207 395045
rect -960 395040 3207 395042
rect -960 394984 3146 395040
rect 3202 394984 3207 395040
rect -960 394982 3207 394984
rect -960 394892 480 394982
rect 3141 394979 3207 394982
rect 540237 394770 540303 394773
rect 539948 394768 540303 394770
rect 539948 394712 540242 394768
rect 540298 394712 540303 394768
rect 539948 394710 540303 394712
rect 540237 394707 540303 394710
rect 256693 393954 256759 393957
rect 256693 393952 260084 393954
rect 256693 393896 256698 393952
rect 256754 393896 260084 393952
rect 256693 393894 260084 393896
rect 256693 393891 256759 393894
rect 580165 393002 580231 393005
rect 583520 393002 584960 393092
rect 580165 393000 584960 393002
rect 580165 392944 580170 393000
rect 580226 392944 584960 393000
rect 580165 392942 584960 392944
rect 580165 392939 580231 392942
rect 583520 392852 584960 392942
rect 541157 392594 541223 392597
rect 539948 392592 541223 392594
rect 539948 392536 541162 392592
rect 541218 392536 541223 392592
rect 539948 392534 541223 392536
rect 541157 392531 541223 392534
rect 256693 391778 256759 391781
rect 256693 391776 260084 391778
rect 256693 391720 256698 391776
rect 256754 391720 260084 391776
rect 256693 391718 260084 391720
rect 256693 391715 256759 391718
rect 539358 391308 539364 391372
rect 539428 391370 539434 391372
rect 539501 391370 539567 391373
rect 539428 391368 539567 391370
rect 539428 391312 539506 391368
rect 539562 391312 539567 391368
rect 539428 391310 539567 391312
rect 539428 391308 539434 391310
rect 539501 391307 539567 391310
rect 540094 390554 540100 390556
rect 539948 390494 540100 390554
rect 540094 390492 540100 390494
rect 540164 390492 540170 390556
rect 256693 389738 256759 389741
rect 256693 389736 260084 389738
rect 256693 389680 256698 389736
rect 256754 389680 260084 389736
rect 256693 389678 260084 389680
rect 256693 389675 256759 389678
rect 543457 389060 543523 389061
rect 543406 389058 543412 389060
rect 543366 388998 543412 389058
rect 543476 389056 543523 389060
rect 543518 389000 543523 389056
rect 543406 388996 543412 388998
rect 543476 388996 543523 389000
rect 543457 388995 543523 388996
rect 539358 388588 539364 388652
rect 539428 388650 539434 388652
rect 539501 388650 539567 388653
rect 539428 388648 539567 388650
rect 539428 388592 539506 388648
rect 539562 388592 539567 388648
rect 539428 388590 539567 388592
rect 539428 388588 539434 388590
rect 539501 388587 539567 388590
rect 539358 388452 539364 388516
rect 539428 388514 539434 388516
rect 539726 388514 539732 388516
rect 539428 388454 539732 388514
rect 539428 388452 539434 388454
rect 539726 388452 539732 388454
rect 539796 388452 539802 388516
rect 539910 388452 539916 388516
rect 539980 388452 539986 388516
rect 539918 388348 539978 388452
rect 256693 387562 256759 387565
rect 256693 387560 260084 387562
rect 256693 387504 256698 387560
rect 256754 387504 260084 387560
rect 256693 387502 260084 387504
rect 256693 387499 256759 387502
rect 541065 386338 541131 386341
rect 539948 386336 541131 386338
rect 539948 386280 541070 386336
rect 541126 386280 541131 386336
rect 539948 386278 541131 386280
rect 541065 386275 541131 386278
rect 256693 385522 256759 385525
rect 256693 385520 260084 385522
rect 256693 385464 256698 385520
rect 256754 385464 260084 385520
rect 256693 385462 260084 385464
rect 256693 385459 256759 385462
rect 539358 384508 539364 384572
rect 539428 384508 539434 384572
rect 539366 384132 539426 384508
rect 539358 383420 539364 383484
rect 539428 383482 539434 383484
rect 539726 383482 539732 383484
rect 539428 383422 539732 383482
rect 539428 383420 539434 383422
rect 539726 383420 539732 383422
rect 539796 383420 539802 383484
rect 256693 383346 256759 383349
rect 256693 383344 260084 383346
rect 256693 383288 256698 383344
rect 256754 383288 260084 383344
rect 256693 383286 260084 383288
rect 256693 383283 256759 383286
rect 540145 382122 540211 382125
rect 539948 382120 540211 382122
rect 539948 382064 540150 382120
rect 540206 382064 540211 382120
rect 539948 382062 540211 382064
rect 540145 382059 540211 382062
rect 256693 381170 256759 381173
rect 256693 381168 260084 381170
rect 256693 381112 256698 381168
rect 256754 381112 260084 381168
rect 583520 381156 584960 381396
rect 256693 381110 260084 381112
rect 256693 381107 256759 381110
rect 539726 380972 539732 381036
rect 539796 381034 539802 381036
rect 540462 381034 540468 381036
rect 539796 380974 540468 381034
rect 539796 380972 539802 380974
rect 540462 380972 540468 380974
rect 540532 380972 540538 381036
rect -960 380626 480 380716
rect 3233 380626 3299 380629
rect -960 380624 3299 380626
rect -960 380568 3238 380624
rect 3294 380568 3299 380624
rect -960 380566 3299 380568
rect -960 380476 480 380566
rect 3233 380563 3299 380566
rect 542169 379946 542235 379949
rect 539948 379944 542235 379946
rect 539948 379888 542174 379944
rect 542230 379888 542235 379944
rect 539948 379886 542235 379888
rect 542169 379883 542235 379886
rect 256693 379130 256759 379133
rect 256693 379128 260084 379130
rect 256693 379072 256698 379128
rect 256754 379072 260084 379128
rect 256693 379070 260084 379072
rect 256693 379067 256759 379070
rect 540053 378042 540119 378045
rect 539918 378040 540119 378042
rect 539918 377984 540058 378040
rect 540114 377984 540119 378040
rect 539918 377982 540119 377984
rect 539918 377876 539978 377982
rect 540053 377979 540119 377982
rect 256693 376954 256759 376957
rect 256693 376952 260084 376954
rect 256693 376896 256698 376952
rect 256754 376896 260084 376952
rect 256693 376894 260084 376896
rect 256693 376891 256759 376894
rect 543365 376684 543431 376685
rect 543365 376680 543412 376684
rect 543476 376682 543482 376684
rect 543365 376624 543370 376680
rect 543365 376620 543412 376624
rect 543476 376622 543522 376682
rect 543476 376620 543482 376622
rect 543365 376619 543431 376620
rect 539358 376348 539364 376412
rect 539428 376410 539434 376412
rect 539726 376410 539732 376412
rect 539428 376350 539732 376410
rect 539428 376348 539434 376350
rect 539726 376348 539732 376350
rect 539796 376348 539802 376412
rect 539358 376212 539364 376276
rect 539428 376212 539434 376276
rect 539366 375700 539426 376212
rect 256693 374914 256759 374917
rect 256693 374912 260084 374914
rect 256693 374856 256698 374912
rect 256754 374856 260084 374912
rect 256693 374854 260084 374856
rect 256693 374851 256759 374854
rect 539358 374580 539364 374644
rect 539428 374642 539434 374644
rect 539726 374642 539732 374644
rect 539428 374582 539732 374642
rect 539428 374580 539434 374582
rect 539726 374580 539732 374582
rect 539796 374580 539802 374644
rect 542077 373690 542143 373693
rect 539948 373688 542143 373690
rect 539948 373632 542082 373688
rect 542138 373632 542143 373688
rect 539948 373630 542143 373632
rect 542077 373627 542143 373630
rect 539501 373282 539567 373285
rect 539726 373282 539732 373284
rect 539501 373280 539732 373282
rect 539501 373224 539506 373280
rect 539562 373224 539732 373280
rect 539501 373222 539732 373224
rect 539501 373219 539567 373222
rect 539726 373220 539732 373222
rect 539796 373220 539802 373284
rect 256693 372738 256759 372741
rect 256693 372736 260084 372738
rect 256693 372680 256698 372736
rect 256754 372680 260084 372736
rect 256693 372678 260084 372680
rect 256693 372675 256759 372678
rect 539961 372058 540027 372061
rect 539918 372056 540027 372058
rect 539918 372000 539966 372056
rect 540022 372000 540027 372056
rect 539918 371995 540027 372000
rect 539918 371484 539978 371995
rect 256693 370562 256759 370565
rect 256693 370560 260084 370562
rect 256693 370504 256698 370560
rect 256754 370504 260084 370560
rect 256693 370502 260084 370504
rect 256693 370499 256759 370502
rect 543457 369748 543523 369749
rect 543406 369746 543412 369748
rect 543366 369686 543412 369746
rect 543476 369744 543523 369748
rect 543518 369688 543523 369744
rect 543406 369684 543412 369686
rect 543476 369684 543523 369688
rect 543457 369683 543523 369684
rect 539869 369610 539935 369613
rect 580257 369610 580323 369613
rect 583520 369610 584960 369700
rect 539869 369608 539978 369610
rect 539869 369552 539874 369608
rect 539930 369552 539978 369608
rect 539869 369547 539978 369552
rect 580257 369608 584960 369610
rect 580257 369552 580262 369608
rect 580318 369552 584960 369608
rect 580257 369550 584960 369552
rect 580257 369547 580323 369550
rect 539918 369444 539978 369547
rect 583520 369460 584960 369550
rect 256693 368522 256759 368525
rect 256693 368520 260084 368522
rect 256693 368464 256698 368520
rect 256754 368464 260084 368520
rect 256693 368462 260084 368464
rect 256693 368459 256759 368462
rect 541985 367298 542051 367301
rect 539948 367296 542051 367298
rect 539948 367240 541990 367296
rect 542046 367240 542051 367296
rect 539948 367238 542051 367240
rect 541985 367235 542051 367238
rect 256693 366346 256759 366349
rect 256693 366344 260084 366346
rect -960 366210 480 366300
rect 256693 366288 256698 366344
rect 256754 366288 260084 366344
rect 256693 366286 260084 366288
rect 256693 366283 256759 366286
rect 3141 366210 3207 366213
rect -960 366208 3207 366210
rect -960 366152 3146 366208
rect 3202 366152 3207 366208
rect -960 366150 3207 366152
rect -960 366060 480 366150
rect 3141 366147 3207 366150
rect 539501 365666 539567 365669
rect 539420 365664 539610 365666
rect 539420 365608 539506 365664
rect 539562 365608 539610 365664
rect 539420 365606 539610 365608
rect 539501 365603 539610 365606
rect 539550 365228 539610 365603
rect 256693 364170 256759 364173
rect 256693 364168 260084 364170
rect 256693 364112 256698 364168
rect 256754 364112 260084 364168
rect 256693 364110 260084 364112
rect 256693 364107 256759 364110
rect 539358 364108 539364 364172
rect 539428 364170 539434 364172
rect 539726 364170 539732 364172
rect 539428 364110 539732 364170
rect 539428 364108 539434 364110
rect 539726 364108 539732 364110
rect 539796 364108 539802 364172
rect 540329 363082 540395 363085
rect 539948 363080 540395 363082
rect 539948 363024 540334 363080
rect 540390 363024 540395 363080
rect 539948 363022 540395 363024
rect 540329 363019 540395 363022
rect 256693 362130 256759 362133
rect 256693 362128 260084 362130
rect 256693 362072 256698 362128
rect 256754 362072 260084 362128
rect 256693 362070 260084 362072
rect 256693 362067 256759 362070
rect 541893 361042 541959 361045
rect 539948 361040 541959 361042
rect 539948 360984 541898 361040
rect 541954 360984 541959 361040
rect 539948 360982 541959 360984
rect 541893 360979 541959 360982
rect 256693 359954 256759 359957
rect 256693 359952 260084 359954
rect 256693 359896 256698 359952
rect 256754 359896 260084 359952
rect 256693 359894 260084 359896
rect 256693 359891 256759 359894
rect 539542 359484 539548 359548
rect 539612 359484 539618 359548
rect 539777 359546 539843 359549
rect 539734 359544 539843 359546
rect 539734 359488 539782 359544
rect 539838 359488 539843 359544
rect 539550 359412 539610 359484
rect 539734 359483 539843 359488
rect 539542 359348 539548 359412
rect 539612 359348 539618 359412
rect 539734 358972 539794 359483
rect 256693 357914 256759 357917
rect 580349 357914 580415 357917
rect 583520 357914 584960 358004
rect 256693 357912 260084 357914
rect 256693 357856 256698 357912
rect 256754 357856 260084 357912
rect 256693 357854 260084 357856
rect 580349 357912 584960 357914
rect 580349 357856 580354 357912
rect 580410 357856 584960 357912
rect 580349 357854 584960 357856
rect 256693 357851 256759 357854
rect 580349 357851 580415 357854
rect 583520 357764 584960 357854
rect 539317 357370 539383 357373
rect 543365 357372 543431 357373
rect 539317 357368 539610 357370
rect 539317 357312 539322 357368
rect 539378 357312 539610 357368
rect 539317 357310 539610 357312
rect 539317 357307 539383 357310
rect 539550 356796 539610 357310
rect 543365 357368 543412 357372
rect 543476 357370 543482 357372
rect 543365 357312 543370 357368
rect 543365 357308 543412 357312
rect 543476 357310 543522 357370
rect 543476 357308 543482 357310
rect 543365 357307 543431 357308
rect 256693 355738 256759 355741
rect 256693 355736 260084 355738
rect 256693 355680 256698 355736
rect 256754 355680 260084 355736
rect 256693 355678 260084 355680
rect 256693 355675 256759 355678
rect 541525 354786 541591 354789
rect 539948 354784 541591 354786
rect 539948 354728 541530 354784
rect 541586 354728 541591 354784
rect 539948 354726 541591 354728
rect 541525 354723 541591 354726
rect 256693 353562 256759 353565
rect 256693 353560 260084 353562
rect 256693 353504 256698 353560
rect 256754 353504 260084 353560
rect 256693 353502 260084 353504
rect 256693 353499 256759 353502
rect 539685 353154 539751 353157
rect 539685 353152 539794 353154
rect 539685 353096 539690 353152
rect 539746 353096 539794 353152
rect 539685 353091 539794 353096
rect 539734 352580 539794 353091
rect -960 351780 480 352020
rect 256693 351522 256759 351525
rect 256693 351520 260084 351522
rect 256693 351464 256698 351520
rect 256754 351464 260084 351520
rect 256693 351462 260084 351464
rect 256693 351459 256759 351462
rect 539409 350706 539475 350709
rect 539366 350704 539475 350706
rect 539366 350648 539414 350704
rect 539470 350648 539475 350704
rect 539366 350643 539475 350648
rect 539366 350540 539426 350643
rect 543457 350436 543523 350437
rect 543406 350434 543412 350436
rect 543366 350374 543412 350434
rect 543476 350432 543523 350436
rect 543518 350376 543523 350432
rect 543406 350372 543412 350374
rect 543476 350372 543523 350376
rect 543457 350371 543523 350372
rect 256693 349346 256759 349349
rect 256693 349344 260084 349346
rect 256693 349288 256698 349344
rect 256754 349288 260084 349344
rect 256693 349286 260084 349288
rect 256693 349283 256759 349286
rect 539726 349012 539732 349076
rect 539796 349012 539802 349076
rect 539734 348938 539794 349012
rect 539961 348938 540027 348941
rect 539734 348936 540027 348938
rect 539734 348880 539966 348936
rect 540022 348880 540027 348936
rect 539734 348878 540027 348880
rect 539961 348875 540027 348878
rect 541433 348394 541499 348397
rect 539948 348392 541499 348394
rect 539948 348336 541438 348392
rect 541494 348336 541499 348392
rect 539948 348334 541499 348336
rect 541433 348331 541499 348334
rect 256693 347170 256759 347173
rect 256693 347168 260084 347170
rect 256693 347112 256698 347168
rect 256754 347112 260084 347168
rect 256693 347110 260084 347112
rect 256693 347107 256759 347110
rect 539593 346490 539659 346493
rect 539550 346488 539659 346490
rect 539550 346432 539598 346488
rect 539654 346432 539659 346488
rect 539550 346427 539659 346432
rect 539550 346324 539610 346427
rect 580441 346082 580507 346085
rect 583520 346082 584960 346172
rect 580441 346080 584960 346082
rect 580441 346024 580446 346080
rect 580502 346024 584960 346080
rect 580441 346022 584960 346024
rect 580441 346019 580507 346022
rect 583520 345932 584960 346022
rect 256693 345130 256759 345133
rect 256693 345128 260084 345130
rect 256693 345072 256698 345128
rect 256754 345072 260084 345128
rect 256693 345070 260084 345072
rect 256693 345067 256759 345070
rect 539317 344314 539383 344317
rect 539317 344312 539426 344314
rect 539317 344256 539322 344312
rect 539378 344256 539426 344312
rect 539317 344251 539426 344256
rect 539366 344148 539426 344251
rect 256693 342954 256759 342957
rect 256693 342952 260084 342954
rect 256693 342896 256698 342952
rect 256754 342896 260084 342952
rect 256693 342894 260084 342896
rect 256693 342891 256759 342894
rect 541341 342138 541407 342141
rect 539948 342136 541407 342138
rect 539948 342080 541346 342136
rect 541402 342080 541407 342136
rect 539948 342078 541407 342080
rect 541341 342075 541407 342078
rect 256693 340914 256759 340917
rect 256693 340912 260084 340914
rect 256693 340856 256698 340912
rect 256754 340856 260084 340912
rect 256693 340854 260084 340856
rect 256693 340851 256759 340854
rect 543457 339962 543523 339965
rect 539948 339960 543523 339962
rect 539948 339904 543462 339960
rect 543518 339904 543523 339960
rect 539948 339902 543523 339904
rect 543457 339899 543523 339902
rect 256693 338738 256759 338741
rect 256693 338736 260084 338738
rect 256693 338680 256698 338736
rect 256754 338680 260084 338736
rect 256693 338678 260084 338680
rect 256693 338675 256759 338678
rect 541801 337922 541867 337925
rect 539948 337920 541867 337922
rect 539948 337864 541806 337920
rect 541862 337864 541867 337920
rect 539948 337862 541867 337864
rect 541801 337859 541867 337862
rect -960 337514 480 337604
rect 3417 337514 3483 337517
rect -960 337512 3483 337514
rect -960 337456 3422 337512
rect 3478 337456 3483 337512
rect -960 337454 3483 337456
rect -960 337364 480 337454
rect 3417 337451 3483 337454
rect 256693 336562 256759 336565
rect 256693 336560 260084 336562
rect 256693 336504 256698 336560
rect 256754 336504 260084 336560
rect 256693 336502 260084 336504
rect 256693 336499 256759 336502
rect 542629 335746 542695 335749
rect 539948 335744 542695 335746
rect 539948 335688 542634 335744
rect 542690 335688 542695 335744
rect 539948 335686 542695 335688
rect 542629 335683 542695 335686
rect 256693 334522 256759 334525
rect 256693 334520 260084 334522
rect 256693 334464 256698 334520
rect 256754 334464 260084 334520
rect 256693 334462 260084 334464
rect 256693 334459 256759 334462
rect 583520 334236 584960 334476
rect 542629 333706 542695 333709
rect 539948 333704 542695 333706
rect 539948 333648 542634 333704
rect 542690 333648 542695 333704
rect 539948 333646 542695 333648
rect 542629 333643 542695 333646
rect 256693 332346 256759 332349
rect 256693 332344 260084 332346
rect 256693 332288 256698 332344
rect 256754 332288 260084 332344
rect 256693 332286 260084 332288
rect 256693 332283 256759 332286
rect 542629 331530 542695 331533
rect 539948 331528 542695 331530
rect 539948 331472 542634 331528
rect 542690 331472 542695 331528
rect 539948 331470 542695 331472
rect 542629 331467 542695 331470
rect 539777 331258 539843 331261
rect 539910 331258 539916 331260
rect 539777 331256 539916 331258
rect 539777 331200 539782 331256
rect 539838 331200 539916 331256
rect 539777 331198 539916 331200
rect 539777 331195 539843 331198
rect 539910 331196 539916 331198
rect 539980 331196 539986 331260
rect 256693 330306 256759 330309
rect 256693 330304 260084 330306
rect 256693 330248 256698 330304
rect 256754 330248 260084 330304
rect 256693 330246 260084 330248
rect 256693 330243 256759 330246
rect 542629 329490 542695 329493
rect 539948 329488 542695 329490
rect 539948 329432 542634 329488
rect 542690 329432 542695 329488
rect 539948 329430 542695 329432
rect 542629 329427 542695 329430
rect 256693 328130 256759 328133
rect 256693 328128 260084 328130
rect 256693 328072 256698 328128
rect 256754 328072 260084 328128
rect 256693 328070 260084 328072
rect 256693 328067 256759 328070
rect 542629 327314 542695 327317
rect 539948 327312 542695 327314
rect 539948 327256 542634 327312
rect 542690 327256 542695 327312
rect 539948 327254 542695 327256
rect 542629 327251 542695 327254
rect 256693 325954 256759 325957
rect 256693 325952 260084 325954
rect 256693 325896 256698 325952
rect 256754 325896 260084 325952
rect 256693 325894 260084 325896
rect 256693 325891 256759 325894
rect 542629 325274 542695 325277
rect 539948 325272 542695 325274
rect 539948 325216 542634 325272
rect 542690 325216 542695 325272
rect 539948 325214 542695 325216
rect 542629 325211 542695 325214
rect 256693 323914 256759 323917
rect 256693 323912 260084 323914
rect 256693 323856 256698 323912
rect 256754 323856 260084 323912
rect 256693 323854 260084 323856
rect 256693 323851 256759 323854
rect -960 323098 480 323188
rect 3233 323098 3299 323101
rect 542629 323098 542695 323101
rect -960 323096 3299 323098
rect -960 323040 3238 323096
rect 3294 323040 3299 323096
rect -960 323038 3299 323040
rect 539948 323096 542695 323098
rect 539948 323040 542634 323096
rect 542690 323040 542695 323096
rect 539948 323038 542695 323040
rect -960 322948 480 323038
rect 3233 323035 3299 323038
rect 542629 323035 542695 323038
rect 580533 322690 580599 322693
rect 583520 322690 584960 322780
rect 580533 322688 584960 322690
rect 580533 322632 580538 322688
rect 580594 322632 584960 322688
rect 580533 322630 584960 322632
rect 580533 322627 580599 322630
rect 583520 322540 584960 322630
rect 256693 321738 256759 321741
rect 256693 321736 260084 321738
rect 256693 321680 256698 321736
rect 256754 321680 260084 321736
rect 256693 321678 260084 321680
rect 256693 321675 256759 321678
rect 542629 321058 542695 321061
rect 539948 321056 542695 321058
rect 539948 321000 542634 321056
rect 542690 321000 542695 321056
rect 539948 320998 542695 321000
rect 542629 320995 542695 320998
rect 256693 319562 256759 319565
rect 256693 319560 260084 319562
rect 256693 319504 256698 319560
rect 256754 319504 260084 319560
rect 256693 319502 260084 319504
rect 256693 319499 256759 319502
rect 542629 318882 542695 318885
rect 539948 318880 542695 318882
rect 539948 318824 542634 318880
rect 542690 318824 542695 318880
rect 539948 318822 542695 318824
rect 542629 318819 542695 318822
rect 256693 317522 256759 317525
rect 256693 317520 260084 317522
rect 256693 317464 256698 317520
rect 256754 317464 260084 317520
rect 256693 317462 260084 317464
rect 256693 317459 256759 317462
rect 542629 316842 542695 316845
rect 539948 316840 542695 316842
rect 539948 316784 542634 316840
rect 542690 316784 542695 316840
rect 539948 316782 542695 316784
rect 542629 316779 542695 316782
rect 256693 315346 256759 315349
rect 256693 315344 260084 315346
rect 256693 315288 256698 315344
rect 256754 315288 260084 315344
rect 256693 315286 260084 315288
rect 256693 315283 256759 315286
rect 542629 314666 542695 314669
rect 539948 314664 542695 314666
rect 539948 314608 542634 314664
rect 542690 314608 542695 314664
rect 539948 314606 542695 314608
rect 542629 314603 542695 314606
rect 256693 313306 256759 313309
rect 256693 313304 260084 313306
rect 256693 313248 256698 313304
rect 256754 313248 260084 313304
rect 256693 313246 260084 313248
rect 256693 313243 256759 313246
rect 542629 312626 542695 312629
rect 539948 312624 542695 312626
rect 539948 312568 542634 312624
rect 542690 312568 542695 312624
rect 539948 312566 542695 312568
rect 542629 312563 542695 312566
rect 256693 311130 256759 311133
rect 256693 311128 260084 311130
rect 256693 311072 256698 311128
rect 256754 311072 260084 311128
rect 256693 311070 260084 311072
rect 256693 311067 256759 311070
rect 580625 310858 580691 310861
rect 583520 310858 584960 310948
rect 580625 310856 584960 310858
rect 580625 310800 580630 310856
rect 580686 310800 584960 310856
rect 580625 310798 584960 310800
rect 580625 310795 580691 310798
rect 583520 310708 584960 310798
rect 542629 310450 542695 310453
rect 539948 310448 542695 310450
rect 539948 310392 542634 310448
rect 542690 310392 542695 310448
rect 539948 310390 542695 310392
rect 542629 310387 542695 310390
rect 256693 308954 256759 308957
rect 256693 308952 260084 308954
rect -960 308818 480 308908
rect 256693 308896 256698 308952
rect 256754 308896 260084 308952
rect 256693 308894 260084 308896
rect 256693 308891 256759 308894
rect 3325 308818 3391 308821
rect -960 308816 3391 308818
rect -960 308760 3330 308816
rect 3386 308760 3391 308816
rect -960 308758 3391 308760
rect -960 308668 480 308758
rect 3325 308755 3391 308758
rect 542629 308410 542695 308413
rect 539948 308408 542695 308410
rect 539948 308352 542634 308408
rect 542690 308352 542695 308408
rect 539948 308350 542695 308352
rect 542629 308347 542695 308350
rect 256693 306914 256759 306917
rect 256693 306912 260084 306914
rect 256693 306856 256698 306912
rect 256754 306856 260084 306912
rect 256693 306854 260084 306856
rect 256693 306851 256759 306854
rect 542629 306234 542695 306237
rect 539948 306232 542695 306234
rect 539948 306176 542634 306232
rect 542690 306176 542695 306232
rect 539948 306174 542695 306176
rect 542629 306171 542695 306174
rect 256693 304738 256759 304741
rect 256693 304736 260084 304738
rect 256693 304680 256698 304736
rect 256754 304680 260084 304736
rect 256693 304678 260084 304680
rect 256693 304675 256759 304678
rect 542629 304194 542695 304197
rect 539948 304192 542695 304194
rect 539948 304136 542634 304192
rect 542690 304136 542695 304192
rect 539948 304134 542695 304136
rect 542629 304131 542695 304134
rect 256693 302562 256759 302565
rect 256693 302560 260084 302562
rect 256693 302504 256698 302560
rect 256754 302504 260084 302560
rect 256693 302502 260084 302504
rect 256693 302499 256759 302502
rect 539910 302364 539916 302428
rect 539980 302364 539986 302428
rect 539918 302154 539978 302364
rect 540094 302154 540100 302156
rect 539918 302094 540100 302154
rect 540094 302092 540100 302094
rect 540164 302092 540170 302156
rect 542629 302018 542695 302021
rect 539948 302016 542695 302018
rect 539948 301960 542634 302016
rect 542690 301960 542695 302016
rect 539948 301958 542695 301960
rect 542629 301955 542695 301958
rect 256693 300522 256759 300525
rect 256693 300520 260084 300522
rect 256693 300464 256698 300520
rect 256754 300464 260084 300520
rect 256693 300462 260084 300464
rect 256693 300459 256759 300462
rect 542629 299978 542695 299981
rect 539948 299976 542695 299978
rect 539948 299920 542634 299976
rect 542690 299920 542695 299976
rect 539948 299918 542695 299920
rect 542629 299915 542695 299918
rect 580717 299162 580783 299165
rect 583520 299162 584960 299252
rect 580717 299160 584960 299162
rect 580717 299104 580722 299160
rect 580778 299104 584960 299160
rect 580717 299102 584960 299104
rect 580717 299099 580783 299102
rect 583520 299012 584960 299102
rect 256693 298346 256759 298349
rect 256693 298344 260084 298346
rect 256693 298288 256698 298344
rect 256754 298288 260084 298344
rect 256693 298286 260084 298288
rect 256693 298283 256759 298286
rect 542629 297938 542695 297941
rect 539948 297936 542695 297938
rect 539948 297880 542634 297936
rect 542690 297880 542695 297936
rect 539948 297878 542695 297880
rect 542629 297875 542695 297878
rect 256693 296306 256759 296309
rect 256693 296304 260084 296306
rect 256693 296248 256698 296304
rect 256754 296248 260084 296304
rect 256693 296246 260084 296248
rect 256693 296243 256759 296246
rect 542629 295762 542695 295765
rect 539948 295760 542695 295762
rect 539948 295704 542634 295760
rect 542690 295704 542695 295760
rect 539948 295702 542695 295704
rect 542629 295699 542695 295702
rect -960 294402 480 294492
rect 3417 294402 3483 294405
rect -960 294400 3483 294402
rect -960 294344 3422 294400
rect 3478 294344 3483 294400
rect -960 294342 3483 294344
rect -960 294252 480 294342
rect 3417 294339 3483 294342
rect 256693 294130 256759 294133
rect 256693 294128 260084 294130
rect 256693 294072 256698 294128
rect 256754 294072 260084 294128
rect 256693 294070 260084 294072
rect 256693 294067 256759 294070
rect 542629 293722 542695 293725
rect 539948 293720 542695 293722
rect 539948 293664 542634 293720
rect 542690 293664 542695 293720
rect 539948 293662 542695 293664
rect 542629 293659 542695 293662
rect 539317 292772 539383 292773
rect 539317 292770 539364 292772
rect 539272 292768 539364 292770
rect 539272 292712 539322 292768
rect 539272 292710 539364 292712
rect 539317 292708 539364 292710
rect 539428 292708 539434 292772
rect 539317 292707 539383 292708
rect 539317 292092 539383 292093
rect 539317 292088 539364 292092
rect 539428 292090 539434 292092
rect 539317 292032 539322 292088
rect 539317 292028 539364 292032
rect 539428 292030 539474 292090
rect 539428 292028 539434 292030
rect 539317 292027 539383 292028
rect 256693 291954 256759 291957
rect 539869 291954 539935 291957
rect 540094 291954 540100 291956
rect 256693 291952 260084 291954
rect 256693 291896 256698 291952
rect 256754 291896 260084 291952
rect 256693 291894 260084 291896
rect 539869 291952 540100 291954
rect 539869 291896 539874 291952
rect 539930 291896 540100 291952
rect 539869 291894 540100 291896
rect 256693 291891 256759 291894
rect 539869 291891 539935 291894
rect 540094 291892 540100 291894
rect 540164 291892 540170 291956
rect 542629 291546 542695 291549
rect 539948 291544 542695 291546
rect 539948 291488 542634 291544
rect 542690 291488 542695 291544
rect 539948 291486 542695 291488
rect 542629 291483 542695 291486
rect 256693 289914 256759 289917
rect 256693 289912 260084 289914
rect 256693 289856 256698 289912
rect 256754 289856 260084 289912
rect 256693 289854 260084 289856
rect 256693 289851 256759 289854
rect 542629 289506 542695 289509
rect 539948 289504 542695 289506
rect 539948 289448 542634 289504
rect 542690 289448 542695 289504
rect 539948 289446 542695 289448
rect 542629 289443 542695 289446
rect 256693 287738 256759 287741
rect 256693 287736 260084 287738
rect 256693 287680 256698 287736
rect 256754 287680 260084 287736
rect 256693 287678 260084 287680
rect 256693 287675 256759 287678
rect 542629 287330 542695 287333
rect 539948 287328 542695 287330
rect 539948 287272 542634 287328
rect 542690 287272 542695 287328
rect 583520 287316 584960 287556
rect 539948 287270 542695 287272
rect 542629 287267 542695 287270
rect 539317 286652 539383 286653
rect 539317 286648 539364 286652
rect 539428 286650 539434 286652
rect 539317 286592 539322 286648
rect 539317 286588 539364 286592
rect 539428 286590 539474 286650
rect 539428 286588 539434 286590
rect 539317 286587 539383 286588
rect 256693 285698 256759 285701
rect 256693 285696 260084 285698
rect 256693 285640 256698 285696
rect 256754 285640 260084 285696
rect 256693 285638 260084 285640
rect 256693 285635 256759 285638
rect 542629 285290 542695 285293
rect 539948 285288 542695 285290
rect 539948 285232 542634 285288
rect 542690 285232 542695 285288
rect 539948 285230 542695 285232
rect 542629 285227 542695 285230
rect 256693 283522 256759 283525
rect 256693 283520 260084 283522
rect 256693 283464 256698 283520
rect 256754 283464 260084 283520
rect 256693 283462 260084 283464
rect 256693 283459 256759 283462
rect 542629 283114 542695 283117
rect 539948 283112 542695 283114
rect 539948 283056 542634 283112
rect 542690 283056 542695 283112
rect 539948 283054 542695 283056
rect 542629 283051 542695 283054
rect 256693 281346 256759 281349
rect 256693 281344 260084 281346
rect 256693 281288 256698 281344
rect 256754 281288 260084 281344
rect 256693 281286 260084 281288
rect 256693 281283 256759 281286
rect 542629 281074 542695 281077
rect 539948 281072 542695 281074
rect 539948 281016 542634 281072
rect 542690 281016 542695 281072
rect 539948 281014 542695 281016
rect 542629 281011 542695 281014
rect -960 280122 480 280212
rect 3417 280122 3483 280125
rect -960 280120 3483 280122
rect -960 280064 3422 280120
rect 3478 280064 3483 280120
rect -960 280062 3483 280064
rect -960 279972 480 280062
rect 3417 280059 3483 280062
rect 541157 279442 541223 279445
rect 539734 279440 541223 279442
rect 539734 279384 541162 279440
rect 541218 279384 541223 279440
rect 539734 279382 541223 279384
rect 256693 279306 256759 279309
rect 256693 279304 260084 279306
rect 256693 279248 256698 279304
rect 256754 279248 260084 279304
rect 256693 279246 260084 279248
rect 256693 279243 256759 279246
rect 539734 278868 539794 279382
rect 541157 279379 541223 279382
rect 539869 279170 539935 279173
rect 540094 279170 540100 279172
rect 539869 279168 540100 279170
rect 539869 279112 539874 279168
rect 539930 279112 540100 279168
rect 539869 279110 540100 279112
rect 539869 279107 539935 279110
rect 540094 279108 540100 279110
rect 540164 279108 540170 279172
rect 256693 277130 256759 277133
rect 256693 277128 260084 277130
rect 256693 277072 256698 277128
rect 256754 277072 260084 277128
rect 256693 277070 260084 277072
rect 256693 277067 256759 277070
rect 543089 276858 543155 276861
rect 539948 276856 543155 276858
rect 539948 276800 543094 276856
rect 543150 276800 543155 276856
rect 539948 276798 543155 276800
rect 543089 276795 543155 276798
rect 580165 275770 580231 275773
rect 583520 275770 584960 275860
rect 580165 275768 584960 275770
rect 580165 275712 580170 275768
rect 580226 275712 584960 275768
rect 580165 275710 584960 275712
rect 580165 275707 580231 275710
rect 583520 275620 584960 275710
rect 256693 274954 256759 274957
rect 256693 274952 260084 274954
rect 256693 274896 256698 274952
rect 256754 274896 260084 274952
rect 256693 274894 260084 274896
rect 256693 274891 256759 274894
rect 542629 274682 542695 274685
rect 539948 274680 542695 274682
rect 539948 274624 542634 274680
rect 542690 274624 542695 274680
rect 539948 274622 542695 274624
rect 542629 274619 542695 274622
rect 539777 273458 539843 273461
rect 540094 273458 540100 273460
rect 539777 273456 540100 273458
rect 539777 273400 539782 273456
rect 539838 273400 540100 273456
rect 539777 273398 540100 273400
rect 539777 273395 539843 273398
rect 540094 273396 540100 273398
rect 540164 273396 540170 273460
rect 256693 272914 256759 272917
rect 256693 272912 260084 272914
rect 256693 272856 256698 272912
rect 256754 272856 260084 272912
rect 256693 272854 260084 272856
rect 256693 272851 256759 272854
rect 542997 272642 543063 272645
rect 539948 272640 543063 272642
rect 539948 272584 543002 272640
rect 543058 272584 543063 272640
rect 539948 272582 543063 272584
rect 542997 272579 543063 272582
rect 256693 270738 256759 270741
rect 256693 270736 260084 270738
rect 256693 270680 256698 270736
rect 256754 270680 260084 270736
rect 256693 270678 260084 270680
rect 256693 270675 256759 270678
rect 543457 270466 543523 270469
rect 539948 270464 543523 270466
rect 539948 270408 543462 270464
rect 543518 270408 543523 270464
rect 539948 270406 543523 270408
rect 543457 270403 543523 270406
rect 256693 268698 256759 268701
rect 256693 268696 260084 268698
rect 256693 268640 256698 268696
rect 256754 268640 260084 268696
rect 256693 268638 260084 268640
rect 256693 268635 256759 268638
rect 543549 268426 543615 268429
rect 539948 268424 543615 268426
rect 539948 268368 543554 268424
rect 543610 268368 543615 268424
rect 539948 268366 543615 268368
rect 543549 268363 543615 268366
rect 256693 266522 256759 266525
rect 256693 266520 260084 266522
rect 256693 266464 256698 266520
rect 256754 266464 260084 266520
rect 256693 266462 260084 266464
rect 256693 266459 256759 266462
rect 543365 266250 543431 266253
rect 539948 266248 543431 266250
rect 539948 266192 543370 266248
rect 543426 266192 543431 266248
rect 539948 266190 543431 266192
rect 543365 266187 543431 266190
rect -960 265706 480 265796
rect 3417 265706 3483 265709
rect -960 265704 3483 265706
rect -960 265648 3422 265704
rect 3478 265648 3483 265704
rect -960 265646 3483 265648
rect -960 265556 480 265646
rect 3417 265643 3483 265646
rect 539317 265028 539383 265029
rect 539777 265028 539843 265029
rect 539317 265026 539364 265028
rect 539272 265024 539364 265026
rect 539272 264968 539322 265024
rect 539272 264966 539364 264968
rect 539317 264964 539364 264966
rect 539428 264964 539434 265028
rect 539726 265026 539732 265028
rect 539686 264966 539732 265026
rect 539796 265024 539843 265028
rect 539838 264968 539843 265024
rect 539726 264964 539732 264966
rect 539796 264964 539843 264968
rect 539317 264963 539383 264964
rect 539777 264963 539843 264964
rect 256693 264346 256759 264349
rect 256693 264344 260084 264346
rect 256693 264288 256698 264344
rect 256754 264288 260084 264344
rect 256693 264286 260084 264288
rect 256693 264283 256759 264286
rect 544377 264210 544443 264213
rect 539948 264208 544443 264210
rect 539948 264152 544382 264208
rect 544438 264152 544443 264208
rect 539948 264150 544443 264152
rect 544377 264147 544443 264150
rect 580165 263938 580231 263941
rect 583520 263938 584960 264028
rect 580165 263936 584960 263938
rect 580165 263880 580170 263936
rect 580226 263880 584960 263936
rect 580165 263878 584960 263880
rect 580165 263875 580231 263878
rect 583520 263788 584960 263878
rect 539726 263604 539732 263668
rect 539796 263666 539802 263668
rect 539796 263606 539978 263666
rect 539796 263604 539802 263606
rect 539918 263532 539978 263606
rect 539910 263468 539916 263532
rect 539980 263468 539986 263532
rect 256693 262306 256759 262309
rect 256693 262304 260084 262306
rect 256693 262248 256698 262304
rect 256754 262248 260084 262304
rect 256693 262246 260084 262248
rect 256693 262243 256759 262246
rect 543273 262034 543339 262037
rect 539948 262032 543339 262034
rect 539948 261976 543278 262032
rect 543334 261976 543339 262032
rect 539948 261974 543339 261976
rect 543273 261971 543339 261974
rect 256693 260130 256759 260133
rect 256693 260128 260084 260130
rect 256693 260072 256698 260128
rect 256754 260072 260084 260128
rect 256693 260070 260084 260072
rect 256693 260067 256759 260070
rect 543089 259994 543155 259997
rect 539948 259992 543155 259994
rect 539948 259936 543094 259992
rect 543150 259936 543155 259992
rect 539948 259934 543155 259936
rect 543089 259931 543155 259934
rect 256693 257954 256759 257957
rect 256693 257952 260084 257954
rect 256693 257896 256698 257952
rect 256754 257896 260084 257952
rect 256693 257894 260084 257896
rect 256693 257891 256759 257894
rect 542629 257818 542695 257821
rect 539948 257816 542695 257818
rect 539948 257760 542634 257816
rect 542690 257760 542695 257816
rect 539948 257758 542695 257760
rect 542629 257755 542695 257758
rect 539358 256804 539364 256868
rect 539428 256804 539434 256868
rect 539366 256732 539426 256804
rect 539358 256668 539364 256732
rect 539428 256668 539434 256732
rect 256693 255914 256759 255917
rect 256693 255912 260084 255914
rect 256693 255856 256698 255912
rect 256754 255856 260084 255912
rect 256693 255854 260084 255856
rect 256693 255851 256759 255854
rect 542629 255778 542695 255781
rect 539948 255776 542695 255778
rect 539948 255720 542634 255776
rect 542690 255720 542695 255776
rect 539948 255718 542695 255720
rect 542629 255715 542695 255718
rect 256693 253738 256759 253741
rect 256693 253736 260084 253738
rect 256693 253680 256698 253736
rect 256754 253680 260084 253736
rect 256693 253678 260084 253680
rect 256693 253675 256759 253678
rect 542629 253602 542695 253605
rect 539948 253600 542695 253602
rect 539948 253544 542634 253600
rect 542690 253544 542695 253600
rect 539948 253542 542695 253544
rect 542629 253539 542695 253542
rect 579797 252242 579863 252245
rect 583520 252242 584960 252332
rect 579797 252240 584960 252242
rect 579797 252184 579802 252240
rect 579858 252184 584960 252240
rect 579797 252182 584960 252184
rect 579797 252179 579863 252182
rect 583520 252092 584960 252182
rect 256693 251698 256759 251701
rect 256693 251696 260084 251698
rect 256693 251640 256698 251696
rect 256754 251640 260084 251696
rect 256693 251638 260084 251640
rect 256693 251635 256759 251638
rect 543089 251562 543155 251565
rect 539948 251560 543155 251562
rect 539948 251504 543094 251560
rect 543150 251504 543155 251560
rect 539948 251502 543155 251504
rect 543089 251499 543155 251502
rect -960 251290 480 251380
rect 3509 251290 3575 251293
rect -960 251288 3575 251290
rect -960 251232 3514 251288
rect 3570 251232 3575 251288
rect -960 251230 3575 251232
rect -960 251140 480 251230
rect 3509 251227 3575 251230
rect 256693 249522 256759 249525
rect 256693 249520 260084 249522
rect 256693 249464 256698 249520
rect 256754 249464 260084 249520
rect 256693 249462 260084 249464
rect 256693 249459 256759 249462
rect 542629 249386 542695 249389
rect 539948 249384 542695 249386
rect 539948 249328 542634 249384
rect 542690 249328 542695 249384
rect 539948 249326 542695 249328
rect 542629 249323 542695 249326
rect 257337 247346 257403 247349
rect 542629 247346 542695 247349
rect 257337 247344 260084 247346
rect 257337 247288 257342 247344
rect 257398 247288 260084 247344
rect 257337 247286 260084 247288
rect 539948 247344 542695 247346
rect 539948 247288 542634 247344
rect 542690 247288 542695 247344
rect 539948 247286 542695 247288
rect 257337 247283 257403 247286
rect 542629 247283 542695 247286
rect 257429 245306 257495 245309
rect 257429 245304 260084 245306
rect 257429 245248 257434 245304
rect 257490 245248 260084 245304
rect 257429 245246 260084 245248
rect 257429 245243 257495 245246
rect 542905 245170 542971 245173
rect 539948 245168 542971 245170
rect 539948 245112 542910 245168
rect 542966 245112 542971 245168
rect 539948 245110 542971 245112
rect 542905 245107 542971 245110
rect 256969 243130 257035 243133
rect 542445 243130 542511 243133
rect 256969 243128 260084 243130
rect 256969 243072 256974 243128
rect 257030 243072 260084 243128
rect 256969 243070 260084 243072
rect 539948 243128 542511 243130
rect 539948 243072 542450 243128
rect 542506 243072 542511 243128
rect 539948 243070 542511 243072
rect 256969 243067 257035 243070
rect 542445 243067 542511 243070
rect 542169 241498 542235 241501
rect 542905 241498 542971 241501
rect 542169 241496 542971 241498
rect 542169 241440 542174 241496
rect 542230 241440 542910 241496
rect 542966 241440 542971 241496
rect 542169 241438 542971 241440
rect 542169 241435 542235 241438
rect 542905 241435 542971 241438
rect 257981 241090 258047 241093
rect 542445 241090 542511 241093
rect 257981 241088 260084 241090
rect 257981 241032 257986 241088
rect 258042 241032 260084 241088
rect 257981 241030 260084 241032
rect 539948 241088 542511 241090
rect 539948 241032 542450 241088
rect 542506 241032 542511 241088
rect 539948 241030 542511 241032
rect 257981 241027 258047 241030
rect 542445 241027 542511 241030
rect 3509 240818 3575 240821
rect 538990 240818 538996 240820
rect 3509 240816 538996 240818
rect 3509 240760 3514 240816
rect 3570 240760 538996 240816
rect 3509 240758 538996 240760
rect 3509 240755 3575 240758
rect 538990 240756 538996 240758
rect 539060 240756 539066 240820
rect 357433 240682 357499 240685
rect 366909 240682 366975 240685
rect 357433 240680 366975 240682
rect 357433 240624 357438 240680
rect 357494 240624 366914 240680
rect 366970 240624 366975 240680
rect 357433 240622 366975 240624
rect 357433 240619 357499 240622
rect 366909 240619 366975 240622
rect 583520 240396 584960 240636
rect -960 237010 480 237100
rect 3417 237010 3483 237013
rect -960 237008 3483 237010
rect -960 236952 3422 237008
rect 3478 236952 3483 237008
rect -960 236950 3483 236952
rect -960 236860 480 236950
rect 3417 236947 3483 236950
rect 580165 228850 580231 228853
rect 583520 228850 584960 228940
rect 580165 228848 584960 228850
rect 580165 228792 580170 228848
rect 580226 228792 584960 228848
rect 580165 228790 584960 228792
rect 580165 228787 580231 228790
rect 583520 228700 584960 228790
rect 538438 227700 538444 227764
rect 538508 227762 538514 227764
rect 538622 227762 538628 227764
rect 538508 227702 538628 227762
rect 538508 227700 538514 227702
rect 538622 227700 538628 227702
rect 538692 227700 538698 227764
rect 538305 222866 538371 222869
rect 538622 222866 538628 222868
rect 538305 222864 538628 222866
rect 538305 222808 538310 222864
rect 538366 222808 538628 222864
rect 538305 222806 538628 222808
rect 538305 222803 538371 222806
rect 538622 222804 538628 222806
rect 538692 222804 538698 222868
rect -960 222594 480 222684
rect 3141 222594 3207 222597
rect -960 222592 3207 222594
rect -960 222536 3146 222592
rect 3202 222536 3207 222592
rect -960 222534 3207 222536
rect -960 222444 480 222534
rect 3141 222531 3207 222534
rect 580165 217018 580231 217021
rect 583520 217018 584960 217108
rect 580165 217016 584960 217018
rect 580165 216960 580170 217016
rect 580226 216960 584960 217016
rect 580165 216958 584960 216960
rect 580165 216955 580231 216958
rect 583520 216868 584960 216958
rect 539961 216066 540027 216069
rect 540094 216066 540100 216068
rect 539961 216064 540100 216066
rect 539961 216008 539966 216064
rect 540022 216008 540100 216064
rect 539961 216006 540100 216008
rect 539961 216003 540027 216006
rect 540094 216004 540100 216006
rect 540164 216004 540170 216068
rect -960 208178 480 208268
rect 3417 208178 3483 208181
rect -960 208176 3483 208178
rect -960 208120 3422 208176
rect 3478 208120 3483 208176
rect -960 208118 3483 208120
rect -960 208028 480 208118
rect 3417 208115 3483 208118
rect 474038 207708 474044 207772
rect 474108 207770 474114 207772
rect 476941 207770 477007 207773
rect 474108 207768 477007 207770
rect 474108 207712 476946 207768
rect 477002 207712 477007 207768
rect 474108 207710 477007 207712
rect 474108 207708 474114 207710
rect 476941 207707 477007 207710
rect 538305 205460 538371 205461
rect 538254 205458 538260 205460
rect 538214 205398 538260 205458
rect 538324 205456 538371 205460
rect 538366 205400 538371 205456
rect 538254 205396 538260 205398
rect 538324 205396 538371 205400
rect 538305 205395 538371 205396
rect 579797 205322 579863 205325
rect 583520 205322 584960 205412
rect 579797 205320 584960 205322
rect 579797 205264 579802 205320
rect 579858 205264 584960 205320
rect 579797 205262 584960 205264
rect 579797 205259 579863 205262
rect 583520 205172 584960 205262
rect 277301 204234 277367 204237
rect 359222 204234 359228 204236
rect 277301 204232 359228 204234
rect 277301 204176 277306 204232
rect 277362 204176 359228 204232
rect 277301 204174 359228 204176
rect 277301 204171 277367 204174
rect 359222 204172 359228 204174
rect 359292 204172 359298 204236
rect 366030 204172 366036 204236
rect 366100 204234 366106 204236
rect 366357 204234 366423 204237
rect 366100 204232 366423 204234
rect 366100 204176 366362 204232
rect 366418 204176 366423 204232
rect 366100 204174 366423 204176
rect 366100 204172 366106 204174
rect 366357 204171 366423 204174
rect 370998 204172 371004 204236
rect 371068 204234 371074 204236
rect 371141 204234 371207 204237
rect 456609 204236 456675 204237
rect 371068 204232 371207 204234
rect 371068 204176 371146 204232
rect 371202 204176 371207 204232
rect 371068 204174 371207 204176
rect 371068 204172 371074 204174
rect 371141 204171 371207 204174
rect 456558 204172 456564 204236
rect 456628 204234 456675 204236
rect 456628 204232 456720 204234
rect 456670 204176 456720 204232
rect 456628 204174 456720 204176
rect 456628 204172 456675 204174
rect 468150 204172 468156 204236
rect 468220 204234 468226 204236
rect 469121 204234 469187 204237
rect 468220 204232 469187 204234
rect 468220 204176 469126 204232
rect 469182 204176 469187 204232
rect 468220 204174 469187 204176
rect 468220 204172 468226 204174
rect 456609 204171 456675 204172
rect 469121 204171 469187 204174
rect 470358 204172 470364 204236
rect 470428 204234 470434 204236
rect 470501 204234 470567 204237
rect 477493 204236 477559 204237
rect 477493 204234 477540 204236
rect 470428 204232 470567 204234
rect 470428 204176 470506 204232
rect 470562 204176 470567 204232
rect 470428 204174 470567 204176
rect 477448 204232 477540 204234
rect 477448 204176 477498 204232
rect 477448 204174 477540 204176
rect 470428 204172 470434 204174
rect 470501 204171 470567 204174
rect 477493 204172 477540 204174
rect 477604 204172 477610 204236
rect 478137 204234 478203 204237
rect 479190 204234 479196 204236
rect 478137 204232 479196 204234
rect 478137 204176 478142 204232
rect 478198 204176 479196 204232
rect 478137 204174 479196 204176
rect 477493 204171 477559 204172
rect 478137 204171 478203 204174
rect 479190 204172 479196 204174
rect 479260 204172 479266 204236
rect 481633 204234 481699 204237
rect 490189 204236 490255 204237
rect 481766 204234 481772 204236
rect 481633 204232 481772 204234
rect 481633 204176 481638 204232
rect 481694 204176 481772 204232
rect 481633 204174 481772 204176
rect 481633 204171 481699 204174
rect 481766 204172 481772 204174
rect 481836 204172 481842 204236
rect 490189 204234 490236 204236
rect 490144 204232 490236 204234
rect 490144 204176 490194 204232
rect 490144 204174 490236 204176
rect 490189 204172 490236 204174
rect 490300 204172 490306 204236
rect 490189 204171 490255 204172
rect 274541 204098 274607 204101
rect 360326 204098 360332 204100
rect 274541 204096 360332 204098
rect 274541 204040 274546 204096
rect 274602 204040 360332 204096
rect 274541 204038 360332 204040
rect 274541 204035 274607 204038
rect 360326 204036 360332 204038
rect 360396 204036 360402 204100
rect 367093 204098 367159 204101
rect 367502 204098 367508 204100
rect 367093 204096 367508 204098
rect 367093 204040 367098 204096
rect 367154 204040 367508 204096
rect 367093 204038 367508 204040
rect 367093 204035 367159 204038
rect 367502 204036 367508 204038
rect 367572 204036 367578 204100
rect 449382 204036 449388 204100
rect 449452 204098 449458 204100
rect 449801 204098 449867 204101
rect 449452 204096 449867 204098
rect 449452 204040 449806 204096
rect 449862 204040 449867 204096
rect 449452 204038 449867 204040
rect 449452 204036 449458 204038
rect 449801 204035 449867 204038
rect 467046 204036 467052 204100
rect 467116 204098 467122 204100
rect 467741 204098 467807 204101
rect 467116 204096 467807 204098
rect 467116 204040 467746 204096
rect 467802 204040 467807 204096
rect 467116 204038 467807 204040
rect 467116 204036 467122 204038
rect 467741 204035 467807 204038
rect 469254 204036 469260 204100
rect 469324 204098 469330 204100
rect 470409 204098 470475 204101
rect 469324 204096 470475 204098
rect 469324 204040 470414 204096
rect 470470 204040 470475 204096
rect 469324 204038 470475 204040
rect 469324 204036 469330 204038
rect 470409 204035 470475 204038
rect 476246 204036 476252 204100
rect 476316 204098 476322 204100
rect 476849 204098 476915 204101
rect 476316 204096 476915 204098
rect 476316 204040 476854 204096
rect 476910 204040 476915 204096
rect 476316 204038 476915 204040
rect 476316 204036 476322 204038
rect 476849 204035 476915 204038
rect 477585 204098 477651 204101
rect 485773 204100 485839 204101
rect 478086 204098 478092 204100
rect 477585 204096 478092 204098
rect 477585 204040 477590 204096
rect 477646 204040 478092 204096
rect 477585 204038 478092 204040
rect 477585 204035 477651 204038
rect 478086 204036 478092 204038
rect 478156 204036 478162 204100
rect 485773 204098 485820 204100
rect 485728 204096 485820 204098
rect 485728 204040 485778 204096
rect 485728 204038 485820 204040
rect 485773 204036 485820 204038
rect 485884 204036 485890 204100
rect 485773 204035 485839 204036
rect 271781 203962 271847 203965
rect 361614 203962 361620 203964
rect 271781 203960 361620 203962
rect 271781 203904 271786 203960
rect 271842 203904 361620 203960
rect 271781 203902 361620 203904
rect 271781 203899 271847 203902
rect 361614 203900 361620 203902
rect 361684 203900 361690 203964
rect 365713 203962 365779 203965
rect 366398 203962 366404 203964
rect 365713 203960 366404 203962
rect 365713 203904 365718 203960
rect 365774 203904 366404 203960
rect 365713 203902 366404 203904
rect 365713 203899 365779 203902
rect 366398 203900 366404 203902
rect 366468 203900 366474 203964
rect 476665 203962 476731 203965
rect 477677 203962 477743 203965
rect 480437 203964 480503 203965
rect 480437 203962 480484 203964
rect 476665 203960 477743 203962
rect 476665 203904 476670 203960
rect 476726 203904 477682 203960
rect 477738 203904 477743 203960
rect 476665 203902 477743 203904
rect 480392 203960 480484 203962
rect 480392 203904 480442 203960
rect 480392 203902 480484 203904
rect 476665 203899 476731 203902
rect 477677 203899 477743 203902
rect 480437 203900 480484 203902
rect 480548 203900 480554 203964
rect 480437 203899 480503 203900
rect 269021 203826 269087 203829
rect 364333 203828 364399 203829
rect 362902 203826 362908 203828
rect 269021 203824 362908 203826
rect 269021 203768 269026 203824
rect 269082 203768 362908 203824
rect 269021 203766 362908 203768
rect 269021 203763 269087 203766
rect 362902 203764 362908 203766
rect 362972 203764 362978 203828
rect 364333 203824 364380 203828
rect 364444 203826 364450 203828
rect 364333 203768 364338 203824
rect 364333 203764 364380 203768
rect 364444 203766 364490 203826
rect 364444 203764 364450 203766
rect 448278 203764 448284 203828
rect 448348 203826 448354 203828
rect 538213 203826 538279 203829
rect 448348 203824 538279 203826
rect 448348 203768 538218 203824
rect 538274 203768 538279 203824
rect 448348 203766 538279 203768
rect 448348 203764 448354 203766
rect 364333 203763 364399 203764
rect 538213 203763 538279 203766
rect 328126 203628 328132 203692
rect 328196 203690 328202 203692
rect 328361 203690 328427 203693
rect 328196 203688 328427 203690
rect 328196 203632 328366 203688
rect 328422 203632 328427 203688
rect 328196 203630 328427 203632
rect 328196 203628 328202 203630
rect 328361 203627 328427 203630
rect 329414 203628 329420 203692
rect 329484 203690 329490 203692
rect 329741 203690 329807 203693
rect 329484 203688 329807 203690
rect 329484 203632 329746 203688
rect 329802 203632 329807 203688
rect 329484 203630 329807 203632
rect 329484 203628 329490 203630
rect 329741 203627 329807 203630
rect 330702 203628 330708 203692
rect 330772 203690 330778 203692
rect 331121 203690 331187 203693
rect 330772 203688 331187 203690
rect 330772 203632 331126 203688
rect 331182 203632 331187 203688
rect 330772 203630 331187 203632
rect 330772 203628 330778 203630
rect 331121 203627 331187 203630
rect 334065 203690 334131 203693
rect 334934 203690 334940 203692
rect 334065 203688 334940 203690
rect 334065 203632 334070 203688
rect 334126 203632 334940 203688
rect 334065 203630 334940 203632
rect 334065 203627 334131 203630
rect 334934 203628 334940 203630
rect 335004 203628 335010 203692
rect 342253 203690 342319 203693
rect 342846 203690 342852 203692
rect 342253 203688 342852 203690
rect 342253 203632 342258 203688
rect 342314 203632 342852 203688
rect 342253 203630 342852 203632
rect 342253 203627 342319 203630
rect 342846 203628 342852 203630
rect 342916 203628 342922 203692
rect 343633 203690 343699 203693
rect 349153 203692 349219 203693
rect 343950 203690 343956 203692
rect 343633 203688 343956 203690
rect 343633 203632 343638 203688
rect 343694 203632 343956 203688
rect 343633 203630 343956 203632
rect 343633 203627 343699 203630
rect 343950 203628 343956 203630
rect 344020 203628 344026 203692
rect 349102 203628 349108 203692
rect 349172 203690 349219 203692
rect 351085 203692 351151 203693
rect 351085 203690 351132 203692
rect 349172 203688 349264 203690
rect 349214 203632 349264 203688
rect 349172 203630 349264 203632
rect 351040 203688 351132 203690
rect 351040 203632 351090 203688
rect 351040 203630 351132 203632
rect 349172 203628 349219 203630
rect 349153 203627 349219 203628
rect 351085 203628 351132 203630
rect 351196 203628 351202 203692
rect 351821 203690 351887 203693
rect 483013 203692 483079 203693
rect 483013 203690 483060 203692
rect 351821 203688 482754 203690
rect 351821 203632 351826 203688
rect 351882 203632 482754 203688
rect 351821 203630 482754 203632
rect 482968 203688 483060 203690
rect 482968 203632 483018 203688
rect 482968 203630 483060 203632
rect 351085 203627 351151 203628
rect 351821 203627 351887 203630
rect 335169 203554 335235 203557
rect 339585 203554 339651 203557
rect 340873 203556 340939 203557
rect 340086 203554 340092 203556
rect 335169 203552 340092 203554
rect 335169 203496 335174 203552
rect 335230 203496 339590 203552
rect 339646 203496 340092 203552
rect 335169 203494 340092 203496
rect 335169 203491 335235 203494
rect 339585 203491 339651 203494
rect 340086 203492 340092 203494
rect 340156 203492 340162 203556
rect 340822 203492 340828 203556
rect 340892 203554 340939 203556
rect 349061 203554 349127 203557
rect 482694 203554 482754 203630
rect 483013 203628 483060 203630
rect 483124 203628 483130 203692
rect 487470 203690 487476 203692
rect 483246 203630 487476 203690
rect 483013 203627 483079 203628
rect 483246 203554 483306 203630
rect 487470 203628 487476 203630
rect 487540 203628 487546 203692
rect 484393 203556 484459 203557
rect 340892 203552 340984 203554
rect 340934 203496 340984 203552
rect 340892 203494 340984 203496
rect 349061 203552 482570 203554
rect 349061 203496 349066 203552
rect 349122 203496 482570 203552
rect 349061 203494 482570 203496
rect 482694 203494 483306 203554
rect 340892 203492 340939 203494
rect 340873 203491 340939 203492
rect 349061 203491 349127 203494
rect 328361 203420 328427 203421
rect 332409 203420 332475 203421
rect 328310 203356 328316 203420
rect 328380 203418 328427 203420
rect 328380 203416 328472 203418
rect 328422 203360 328472 203416
rect 328380 203358 328472 203360
rect 328380 203356 328427 203358
rect 332358 203356 332364 203420
rect 332428 203418 332475 203420
rect 332428 203416 332520 203418
rect 332470 203360 332520 203416
rect 332428 203358 332520 203360
rect 332428 203356 332475 203358
rect 332910 203356 332916 203420
rect 332980 203418 332986 203420
rect 333881 203418 333947 203421
rect 336641 203420 336707 203421
rect 332980 203416 333947 203418
rect 332980 203360 333886 203416
rect 333942 203360 333947 203416
rect 332980 203358 333947 203360
rect 332980 203356 332986 203358
rect 328361 203355 328427 203356
rect 332409 203355 332475 203356
rect 333881 203355 333947 203358
rect 336590 203356 336596 203420
rect 336660 203418 336707 203420
rect 338113 203418 338179 203421
rect 357433 203420 357499 203421
rect 338246 203418 338252 203420
rect 336660 203416 336752 203418
rect 336702 203360 336752 203416
rect 336660 203358 336752 203360
rect 338113 203416 338252 203418
rect 338113 203360 338118 203416
rect 338174 203360 338252 203416
rect 338113 203358 338252 203360
rect 336660 203356 336707 203358
rect 336641 203355 336707 203356
rect 338113 203355 338179 203358
rect 338246 203356 338252 203358
rect 338316 203356 338322 203420
rect 357382 203356 357388 203420
rect 357452 203418 357499 203420
rect 449157 203418 449223 203421
rect 449566 203418 449572 203420
rect 357452 203416 357544 203418
rect 357494 203360 357544 203416
rect 357452 203358 357544 203360
rect 449157 203416 449572 203418
rect 449157 203360 449162 203416
rect 449218 203360 449572 203416
rect 449157 203358 449572 203360
rect 357452 203356 357499 203358
rect 357433 203355 357499 203356
rect 449157 203355 449223 203358
rect 449566 203356 449572 203358
rect 449636 203356 449642 203420
rect 450537 203418 450603 203421
rect 450854 203418 450860 203420
rect 450537 203416 450860 203418
rect 450537 203360 450542 203416
rect 450598 203360 450860 203416
rect 450537 203358 450860 203360
rect 450537 203355 450603 203358
rect 450854 203356 450860 203358
rect 450924 203356 450930 203420
rect 451917 203418 451983 203421
rect 453297 203420 453363 203421
rect 452142 203418 452148 203420
rect 451917 203416 452148 203418
rect 451917 203360 451922 203416
rect 451978 203360 452148 203416
rect 451917 203358 452148 203360
rect 451917 203355 451983 203358
rect 452142 203356 452148 203358
rect 452212 203356 452218 203420
rect 453246 203356 453252 203420
rect 453316 203418 453363 203420
rect 453316 203416 453408 203418
rect 453358 203360 453408 203416
rect 453316 203358 453408 203360
rect 453316 203356 453363 203358
rect 456006 203356 456012 203420
rect 456076 203418 456082 203420
rect 456149 203418 456215 203421
rect 456076 203416 456215 203418
rect 456076 203360 456154 203416
rect 456210 203360 456215 203416
rect 456076 203358 456215 203360
rect 456076 203356 456082 203358
rect 453297 203355 453363 203356
rect 456149 203355 456215 203358
rect 458766 203356 458772 203420
rect 458836 203418 458842 203420
rect 459461 203418 459527 203421
rect 458836 203416 459527 203418
rect 458836 203360 459466 203416
rect 459522 203360 459527 203416
rect 458836 203358 459527 203360
rect 458836 203356 458842 203358
rect 459461 203355 459527 203358
rect 460974 203356 460980 203420
rect 461044 203418 461050 203420
rect 462129 203418 462195 203421
rect 461044 203416 462195 203418
rect 461044 203360 462134 203416
rect 462190 203360 462195 203416
rect 461044 203358 462195 203360
rect 461044 203356 461050 203358
rect 462129 203355 462195 203358
rect 462262 203356 462268 203420
rect 462332 203418 462338 203420
rect 463509 203418 463575 203421
rect 462332 203416 463575 203418
rect 462332 203360 463514 203416
rect 463570 203360 463575 203416
rect 462332 203358 463575 203360
rect 462332 203356 462338 203358
rect 463509 203355 463575 203358
rect 477585 203418 477651 203421
rect 478638 203418 478644 203420
rect 477585 203416 478644 203418
rect 477585 203360 477590 203416
rect 477646 203360 478644 203416
rect 477585 203358 478644 203360
rect 477585 203355 477651 203358
rect 478638 203356 478644 203358
rect 478708 203356 478714 203420
rect 331121 203284 331187 203285
rect 331070 203220 331076 203284
rect 331140 203282 331187 203284
rect 331140 203280 331232 203282
rect 331182 203224 331232 203280
rect 331140 203222 331232 203224
rect 331140 203220 331187 203222
rect 331622 203220 331628 203284
rect 331692 203282 331698 203284
rect 332501 203282 332567 203285
rect 333973 203284 334039 203285
rect 333973 203282 334020 203284
rect 331692 203280 332567 203282
rect 331692 203224 332506 203280
rect 332562 203224 332567 203280
rect 331692 203222 332567 203224
rect 333928 203280 334020 203282
rect 333928 203224 333978 203280
rect 333928 203222 334020 203224
rect 331692 203220 331698 203222
rect 331121 203219 331187 203220
rect 332501 203219 332567 203222
rect 333973 203220 334020 203222
rect 334084 203220 334090 203284
rect 335353 203282 335419 203285
rect 336222 203282 336228 203284
rect 335353 203280 336228 203282
rect 335353 203224 335358 203280
rect 335414 203224 336228 203280
rect 335353 203222 336228 203224
rect 333973 203219 334039 203220
rect 335353 203219 335419 203222
rect 336222 203220 336228 203222
rect 336292 203220 336298 203284
rect 336733 203282 336799 203285
rect 339493 203284 339559 203285
rect 336958 203282 336964 203284
rect 336733 203280 336964 203282
rect 336733 203224 336738 203280
rect 336794 203224 336964 203280
rect 336733 203222 336964 203224
rect 336733 203219 336799 203222
rect 336958 203220 336964 203222
rect 337028 203220 337034 203284
rect 339493 203282 339540 203284
rect 339448 203280 339540 203282
rect 339448 203224 339498 203280
rect 339448 203222 339540 203224
rect 339493 203220 339540 203222
rect 339604 203220 339610 203284
rect 345013 203282 345079 203285
rect 345238 203282 345244 203284
rect 345013 203280 345244 203282
rect 345013 203224 345018 203280
rect 345074 203224 345244 203280
rect 345013 203222 345244 203224
rect 339493 203219 339559 203220
rect 345013 203219 345079 203222
rect 345238 203220 345244 203222
rect 345308 203220 345314 203284
rect 349153 203282 349219 203285
rect 349838 203282 349844 203284
rect 349153 203280 349844 203282
rect 349153 203224 349158 203280
rect 349214 203224 349844 203280
rect 349153 203222 349844 203224
rect 349153 203219 349219 203222
rect 349838 203220 349844 203222
rect 349908 203220 349914 203284
rect 368473 203282 368539 203285
rect 368606 203282 368612 203284
rect 368473 203280 368612 203282
rect 368473 203224 368478 203280
rect 368534 203224 368612 203280
rect 368473 203222 368612 203224
rect 368473 203219 368539 203222
rect 368606 203220 368612 203222
rect 368676 203220 368682 203284
rect 450670 203220 450676 203284
rect 450740 203282 450746 203284
rect 451181 203282 451247 203285
rect 450740 203280 451247 203282
rect 450740 203224 451186 203280
rect 451242 203224 451247 203280
rect 450740 203222 451247 203224
rect 450740 203220 450746 203222
rect 451181 203219 451247 203222
rect 452878 203220 452884 203284
rect 452948 203282 452954 203284
rect 453941 203282 454007 203285
rect 452948 203280 454007 203282
rect 452948 203224 453946 203280
rect 454002 203224 454007 203280
rect 452948 203222 454007 203224
rect 452948 203220 452954 203222
rect 453941 203219 454007 203222
rect 454677 203282 454743 203285
rect 454902 203282 454908 203284
rect 454677 203280 454908 203282
rect 454677 203224 454682 203280
rect 454738 203224 454908 203280
rect 454677 203222 454908 203224
rect 454677 203219 454743 203222
rect 454902 203220 454908 203222
rect 454972 203282 454978 203284
rect 455045 203282 455111 203285
rect 455229 203284 455295 203285
rect 455229 203282 455276 203284
rect 454972 203280 455111 203282
rect 454972 203224 455050 203280
rect 455106 203224 455111 203280
rect 454972 203222 455111 203224
rect 455184 203280 455276 203282
rect 455184 203224 455234 203280
rect 455184 203222 455276 203224
rect 454972 203220 454978 203222
rect 455045 203219 455111 203222
rect 455229 203220 455276 203222
rect 455340 203220 455346 203284
rect 457478 203220 457484 203284
rect 457548 203282 457554 203284
rect 458081 203282 458147 203285
rect 457548 203280 458147 203282
rect 457548 203224 458086 203280
rect 458142 203224 458147 203280
rect 457548 203222 458147 203224
rect 457548 203220 457554 203222
rect 455229 203219 455295 203220
rect 458081 203219 458147 203222
rect 460054 203220 460060 203284
rect 460124 203282 460130 203284
rect 460841 203282 460907 203285
rect 460124 203280 460907 203282
rect 460124 203224 460846 203280
rect 460902 203224 460907 203280
rect 460124 203222 460907 203224
rect 460124 203220 460130 203222
rect 460841 203219 460907 203222
rect 463182 203220 463188 203284
rect 463252 203282 463258 203284
rect 463601 203282 463667 203285
rect 463252 203280 463667 203282
rect 463252 203224 463606 203280
rect 463662 203224 463667 203280
rect 463252 203222 463667 203224
rect 463252 203220 463258 203222
rect 463601 203219 463667 203222
rect 464613 203284 464679 203285
rect 464613 203280 464660 203284
rect 464724 203282 464730 203284
rect 465073 203282 465139 203285
rect 465942 203282 465948 203284
rect 464613 203224 464618 203280
rect 464613 203220 464660 203224
rect 464724 203222 464770 203282
rect 465073 203280 465948 203282
rect 465073 203224 465078 203280
rect 465134 203224 465948 203280
rect 465073 203222 465948 203224
rect 464724 203220 464730 203222
rect 464613 203219 464679 203220
rect 465073 203219 465139 203222
rect 465942 203220 465948 203222
rect 466012 203282 466018 203284
rect 466545 203282 466611 203285
rect 466012 203280 466611 203282
rect 466012 203224 466550 203280
rect 466606 203224 466611 203280
rect 466012 203222 466611 203224
rect 466012 203220 466018 203222
rect 466545 203219 466611 203222
rect 471646 203220 471652 203284
rect 471716 203282 471722 203284
rect 471881 203282 471947 203285
rect 471716 203280 471947 203282
rect 471716 203224 471886 203280
rect 471942 203224 471947 203280
rect 471716 203222 471947 203224
rect 471716 203220 471722 203222
rect 471881 203219 471947 203222
rect 472750 203220 472756 203284
rect 472820 203282 472826 203284
rect 473261 203282 473327 203285
rect 472820 203280 473327 203282
rect 472820 203224 473266 203280
rect 473322 203224 473327 203280
rect 472820 203222 473327 203224
rect 472820 203220 472826 203222
rect 473261 203219 473327 203222
rect 475142 203220 475148 203284
rect 475212 203282 475218 203284
rect 476021 203282 476087 203285
rect 475212 203280 476087 203282
rect 475212 203224 476026 203280
rect 476082 203224 476087 203280
rect 475212 203222 476087 203224
rect 475212 203220 475218 203222
rect 476021 203219 476087 203222
rect 477493 203282 477559 203285
rect 477718 203282 477724 203284
rect 477493 203280 477724 203282
rect 477493 203224 477498 203280
rect 477554 203224 477724 203280
rect 477493 203222 477724 203224
rect 477493 203219 477559 203222
rect 477718 203220 477724 203222
rect 477788 203220 477794 203284
rect 482510 203282 482570 203494
rect 484342 203492 484348 203556
rect 484412 203554 484459 203556
rect 488574 203554 488580 203556
rect 484412 203552 484504 203554
rect 484454 203496 484504 203552
rect 484412 203494 484504 203496
rect 484594 203494 488580 203554
rect 484412 203492 484459 203494
rect 484393 203491 484459 203492
rect 484594 203282 484654 203494
rect 488574 203492 488580 203494
rect 488644 203492 488650 203556
rect 482510 203222 484654 203282
rect 485773 203282 485839 203285
rect 486366 203282 486372 203284
rect 485773 203280 486372 203282
rect 485773 203224 485778 203280
rect 485834 203224 486372 203280
rect 485773 203222 486372 203224
rect 485773 203219 485839 203222
rect 486366 203220 486372 203222
rect 486436 203220 486442 203284
rect 329598 203084 329604 203148
rect 329668 203146 329674 203148
rect 329741 203146 329807 203149
rect 329668 203144 329807 203146
rect 329668 203088 329746 203144
rect 329802 203088 329807 203144
rect 329668 203086 329807 203088
rect 329668 203084 329674 203086
rect 329741 203083 329807 203086
rect 333646 203084 333652 203148
rect 333716 203146 333722 203148
rect 333881 203146 333947 203149
rect 333716 203144 333947 203146
rect 333716 203088 333886 203144
rect 333942 203088 333947 203144
rect 333716 203086 333947 203088
rect 333716 203084 333722 203086
rect 333881 203083 333947 203086
rect 334750 203084 334756 203148
rect 334820 203146 334826 203148
rect 335261 203146 335327 203149
rect 334820 203144 335327 203146
rect 334820 203088 335266 203144
rect 335322 203088 335327 203144
rect 334820 203086 335327 203088
rect 334820 203084 334826 203086
rect 335261 203083 335327 203086
rect 341742 203084 341748 203148
rect 341812 203146 341818 203148
rect 342161 203146 342227 203149
rect 341812 203144 342227 203146
rect 341812 203088 342166 203144
rect 342222 203088 342227 203144
rect 341812 203086 342227 203088
rect 341812 203084 341818 203086
rect 342161 203083 342227 203086
rect 346393 203146 346459 203149
rect 347773 203148 347839 203149
rect 346526 203146 346532 203148
rect 346393 203144 346532 203146
rect 346393 203088 346398 203144
rect 346454 203088 346532 203144
rect 346393 203086 346532 203088
rect 346393 203083 346459 203086
rect 346526 203084 346532 203086
rect 346596 203084 346602 203148
rect 347773 203146 347820 203148
rect 347728 203144 347820 203146
rect 347728 203088 347778 203144
rect 347728 203086 347820 203088
rect 347773 203084 347820 203086
rect 347884 203084 347890 203148
rect 351913 203146 351979 203149
rect 353201 203148 353267 203149
rect 352782 203146 352788 203148
rect 351913 203144 352788 203146
rect 351913 203088 351918 203144
rect 351974 203088 352788 203144
rect 351913 203086 352788 203088
rect 347773 203083 347839 203084
rect 351913 203083 351979 203086
rect 352782 203084 352788 203086
rect 352852 203084 352858 203148
rect 353150 203146 353156 203148
rect 353110 203086 353156 203146
rect 353220 203144 353267 203148
rect 353262 203088 353267 203144
rect 353150 203084 353156 203086
rect 353220 203084 353267 203088
rect 353201 203083 353267 203084
rect 354673 203146 354739 203149
rect 356053 203148 356119 203149
rect 357801 203148 357867 203149
rect 354806 203146 354812 203148
rect 354673 203144 354812 203146
rect 354673 203088 354678 203144
rect 354734 203088 354812 203144
rect 354673 203086 354812 203088
rect 354673 203083 354739 203086
rect 354806 203084 354812 203086
rect 354876 203084 354882 203148
rect 356053 203146 356100 203148
rect 356008 203144 356100 203146
rect 356008 203088 356058 203144
rect 356008 203086 356100 203088
rect 356053 203084 356100 203086
rect 356164 203084 356170 203148
rect 357750 203146 357756 203148
rect 357710 203086 357756 203146
rect 357820 203144 357867 203148
rect 357862 203088 357867 203144
rect 357750 203084 357756 203086
rect 357820 203084 357867 203088
rect 356053 203083 356119 203084
rect 357801 203083 357867 203084
rect 373257 203146 373323 203149
rect 373390 203146 373396 203148
rect 373257 203144 373396 203146
rect 373257 203088 373262 203144
rect 373318 203088 373396 203144
rect 373257 203086 373396 203088
rect 373257 203083 373323 203086
rect 373390 203084 373396 203086
rect 373460 203146 373466 203148
rect 492806 203146 492812 203148
rect 373460 203086 492812 203146
rect 373460 203084 373466 203086
rect 492806 203084 492812 203086
rect 492876 203084 492882 203148
rect 336038 202948 336044 203012
rect 336108 203010 336114 203012
rect 336641 203010 336707 203013
rect 337929 203012 337995 203013
rect 339217 203012 339283 203013
rect 337878 203010 337884 203012
rect 336108 203008 336707 203010
rect 336108 202952 336646 203008
rect 336702 202952 336707 203008
rect 336108 202950 336707 202952
rect 337838 202950 337884 203010
rect 337948 203008 337995 203012
rect 339166 203010 339172 203012
rect 337990 202952 337995 203008
rect 336108 202948 336114 202950
rect 336641 202947 336707 202950
rect 337878 202948 337884 202950
rect 337948 202948 337995 202952
rect 339126 202950 339172 203010
rect 339236 203008 339283 203012
rect 342253 203012 342319 203013
rect 342437 203012 342503 203013
rect 343633 203012 343699 203013
rect 344921 203012 344987 203013
rect 342253 203010 342300 203012
rect 339278 202952 339283 203008
rect 339166 202948 339172 202950
rect 339236 202948 339283 202952
rect 342208 203008 342300 203010
rect 342208 202952 342258 203008
rect 342208 202950 342300 202952
rect 337929 202947 337995 202948
rect 339217 202947 339283 202948
rect 342253 202948 342300 202950
rect 342364 202948 342370 203012
rect 342437 203008 342484 203012
rect 342548 203010 342554 203012
rect 343582 203010 343588 203012
rect 342437 202952 342442 203008
rect 342437 202948 342484 202952
rect 342548 202950 342594 203010
rect 343542 202950 343588 203010
rect 343652 203008 343699 203012
rect 344870 203010 344876 203012
rect 343694 202952 343699 203008
rect 342548 202948 342554 202950
rect 343582 202948 343588 202950
rect 343652 202948 343699 202952
rect 344830 202950 344876 203010
rect 344940 203008 344987 203012
rect 344982 202952 344987 203008
rect 344870 202948 344876 202950
rect 344940 202948 344987 202952
rect 342253 202947 342319 202948
rect 342437 202947 342503 202948
rect 343633 202947 343699 202948
rect 344921 202947 344987 202948
rect 345933 203012 345999 203013
rect 347129 203012 347195 203013
rect 345933 203008 345980 203012
rect 346044 203010 346050 203012
rect 347078 203010 347084 203012
rect 345933 202952 345938 203008
rect 345933 202948 345980 202952
rect 346044 202950 346090 203010
rect 347038 202950 347084 203010
rect 347148 203008 347195 203012
rect 347190 202952 347195 203008
rect 346044 202948 346050 202950
rect 347078 202948 347084 202950
rect 347148 202948 347195 202952
rect 345933 202947 345999 202948
rect 347129 202947 347195 202948
rect 348325 203012 348391 203013
rect 348325 203008 348372 203012
rect 348436 203010 348442 203012
rect 349245 203010 349311 203013
rect 350993 203012 351059 203013
rect 351729 203012 351795 203013
rect 349654 203010 349660 203012
rect 348325 202952 348330 203008
rect 348325 202948 348372 202952
rect 348436 202950 348482 203010
rect 349245 203008 349660 203010
rect 349245 202952 349250 203008
rect 349306 202952 349660 203008
rect 349245 202950 349660 202952
rect 348436 202948 348442 202950
rect 348325 202947 348391 202948
rect 349245 202947 349311 202950
rect 349654 202948 349660 202950
rect 349724 202948 349730 203012
rect 350942 203010 350948 203012
rect 350902 202950 350948 203010
rect 351012 203008 351059 203012
rect 351678 203010 351684 203012
rect 351054 202952 351059 203008
rect 350942 202948 350948 202950
rect 351012 202948 351059 202952
rect 351638 202950 351684 203010
rect 351748 203008 351795 203012
rect 353293 203012 353359 203013
rect 354305 203012 354371 203013
rect 355593 203012 355659 203013
rect 353293 203010 353340 203012
rect 351790 202952 351795 203008
rect 351678 202948 351684 202950
rect 351748 202948 351795 202952
rect 353248 203008 353340 203010
rect 353248 202952 353298 203008
rect 353248 202950 353340 202952
rect 350993 202947 351059 202948
rect 351729 202947 351795 202948
rect 353293 202948 353340 202950
rect 353404 202948 353410 203012
rect 354254 203010 354260 203012
rect 354214 202950 354260 203010
rect 354324 203008 354371 203012
rect 355542 203010 355548 203012
rect 354366 202952 354371 203008
rect 354254 202948 354260 202950
rect 354324 202948 354371 202952
rect 355502 202950 355548 203010
rect 355612 203008 355659 203012
rect 355654 202952 355659 203008
rect 355542 202948 355548 202950
rect 355612 202948 355659 202952
rect 353293 202947 353359 202948
rect 354305 202947 354371 202948
rect 355593 202947 355659 202948
rect 356421 203012 356487 203013
rect 356421 203008 356468 203012
rect 356532 203010 356538 203012
rect 357433 203010 357499 203013
rect 358629 203012 358695 203013
rect 360009 203012 360075 203013
rect 361297 203012 361363 203013
rect 357934 203010 357940 203012
rect 356421 202952 356426 203008
rect 356421 202948 356468 202952
rect 356532 202950 356578 203010
rect 357433 203008 357940 203010
rect 357433 202952 357438 203008
rect 357494 202952 357940 203008
rect 357433 202950 357940 202952
rect 356532 202948 356538 202950
rect 356421 202947 356487 202948
rect 357433 202947 357499 202950
rect 357934 202948 357940 202950
rect 358004 202948 358010 203012
rect 358629 203008 358676 203012
rect 358740 203010 358746 203012
rect 359958 203010 359964 203012
rect 358629 202952 358634 203008
rect 358629 202948 358676 202952
rect 358740 202950 358786 203010
rect 359918 202950 359964 203010
rect 360028 203008 360075 203012
rect 361246 203010 361252 203012
rect 360070 202952 360075 203008
rect 358740 202948 358746 202950
rect 359958 202948 359964 202950
rect 360028 202948 360075 202952
rect 361206 202950 361252 203010
rect 361316 203008 361363 203012
rect 361358 202952 361363 203008
rect 361246 202948 361252 202950
rect 361316 202948 361363 202952
rect 358629 202947 358695 202948
rect 360009 202947 360075 202948
rect 361297 202947 361363 202948
rect 362493 203012 362559 203013
rect 363505 203012 363571 203013
rect 362493 203008 362540 203012
rect 362604 203010 362610 203012
rect 363454 203010 363460 203012
rect 362493 202952 362498 203008
rect 362493 202948 362540 202952
rect 362604 202950 362650 203010
rect 363414 202950 363460 203010
rect 363524 203008 363571 203012
rect 363566 202952 363571 203008
rect 362604 202948 362610 202950
rect 363454 202948 363460 202950
rect 363524 202948 363571 202952
rect 362493 202947 362559 202948
rect 363505 202947 363571 202948
rect 364701 203012 364767 203013
rect 364701 203008 364748 203012
rect 364812 203010 364818 203012
rect 364701 202952 364706 203008
rect 364701 202948 364748 202952
rect 364812 202950 364858 203010
rect 364812 202948 364818 202950
rect 451774 202948 451780 203012
rect 451844 203010 451850 203012
rect 452561 203010 452627 203013
rect 451844 203008 452627 203010
rect 451844 202952 452566 203008
rect 452622 202952 452627 203008
rect 451844 202950 452627 202952
rect 451844 202948 451850 202950
rect 364701 202947 364767 202948
rect 452561 202947 452627 202950
rect 454166 202948 454172 203012
rect 454236 203010 454242 203012
rect 455321 203010 455387 203013
rect 454236 203008 455387 203010
rect 454236 202952 455326 203008
rect 455382 202952 455387 203008
rect 454236 202950 455387 202952
rect 454236 202948 454242 202950
rect 455321 202947 455387 202950
rect 456374 202948 456380 203012
rect 456444 203010 456450 203012
rect 456609 203010 456675 203013
rect 456444 203008 456675 203010
rect 456444 202952 456614 203008
rect 456670 202952 456675 203008
rect 456444 202950 456675 202952
rect 456444 202948 456450 202950
rect 456609 202947 456675 202950
rect 457846 202948 457852 203012
rect 457916 203010 457922 203012
rect 457989 203010 458055 203013
rect 459001 203012 459067 203013
rect 458950 203010 458956 203012
rect 457916 203008 458055 203010
rect 457916 202952 457994 203008
rect 458050 202952 458055 203008
rect 457916 202950 458055 202952
rect 458910 202950 458956 203010
rect 459020 203008 459067 203012
rect 459062 202952 459067 203008
rect 457916 202948 457922 202950
rect 457989 202947 458055 202950
rect 458950 202948 458956 202950
rect 459020 202948 459067 202952
rect 460422 202948 460428 203012
rect 460492 203010 460498 203012
rect 460565 203010 460631 203013
rect 460492 203008 460631 203010
rect 460492 202952 460570 203008
rect 460626 202952 460631 203008
rect 460492 202950 460631 202952
rect 460492 202948 460498 202950
rect 459001 202947 459067 202948
rect 460565 202947 460631 202950
rect 461393 203010 461459 203013
rect 462405 203012 462471 203013
rect 463601 203012 463667 203013
rect 461526 203010 461532 203012
rect 461393 203008 461532 203010
rect 461393 202952 461398 203008
rect 461454 202952 461532 203008
rect 461393 202950 461532 202952
rect 461393 202947 461459 202950
rect 461526 202948 461532 202950
rect 461596 202948 461602 203012
rect 462405 203008 462452 203012
rect 462516 203010 462522 203012
rect 463550 203010 463556 203012
rect 462405 202952 462410 203008
rect 462405 202948 462452 202952
rect 462516 202950 462562 203010
rect 463510 202950 463556 203010
rect 463620 203008 463667 203012
rect 463662 202952 463667 203008
rect 462516 202948 462522 202950
rect 463550 202948 463556 202950
rect 463620 202948 463667 202952
rect 464470 202948 464476 203012
rect 464540 203010 464546 203012
rect 464981 203010 465047 203013
rect 464540 203008 465047 203010
rect 464540 202952 464986 203008
rect 465042 202952 465047 203008
rect 464540 202950 465047 202952
rect 464540 202948 464546 202950
rect 462405 202947 462471 202948
rect 463601 202947 463667 202948
rect 464981 202947 465047 202950
rect 465758 202948 465764 203012
rect 465828 203010 465834 203012
rect 466361 203010 466427 203013
rect 467281 203012 467347 203013
rect 467230 203010 467236 203012
rect 465828 203008 466427 203010
rect 465828 202952 466366 203008
rect 466422 202952 466427 203008
rect 465828 202950 466427 202952
rect 467190 202950 467236 203010
rect 467300 203008 467347 203012
rect 467342 202952 467347 203008
rect 465828 202948 465834 202950
rect 466361 202947 466427 202950
rect 467230 202948 467236 202950
rect 467300 202948 467347 202952
rect 467281 202947 467347 202948
rect 468477 203012 468543 203013
rect 469397 203012 469463 203013
rect 470685 203012 470751 203013
rect 468477 203008 468524 203012
rect 468588 203010 468594 203012
rect 468477 202952 468482 203008
rect 468477 202948 468524 202952
rect 468588 202950 468634 203010
rect 469397 203008 469444 203012
rect 469508 203010 469514 203012
rect 469397 202952 469402 203008
rect 468588 202948 468594 202950
rect 469397 202948 469444 202952
rect 469508 202950 469554 203010
rect 470685 203008 470732 203012
rect 470796 203010 470802 203012
rect 471605 203010 471671 203013
rect 470796 203008 471671 203010
rect 470685 202952 470690 203008
rect 470796 202952 471610 203008
rect 471666 202952 471671 203008
rect 469508 202948 469514 202950
rect 470685 202948 470732 202952
rect 470796 202950 471671 202952
rect 470796 202948 470802 202950
rect 468477 202947 468543 202948
rect 469397 202947 469463 202948
rect 470685 202947 470751 202948
rect 471605 202947 471671 202950
rect 471789 203012 471855 203013
rect 472893 203012 472959 203013
rect 474181 203012 474247 203013
rect 475561 203012 475627 203013
rect 471789 203008 471836 203012
rect 471900 203010 471906 203012
rect 471789 202952 471794 203008
rect 471789 202948 471836 202952
rect 471900 202950 471946 203010
rect 472893 203008 472940 203012
rect 473004 203010 473010 203012
rect 472893 202952 472898 203008
rect 471900 202948 471906 202950
rect 472893 202948 472940 202952
rect 473004 202950 473050 203010
rect 474181 203008 474228 203012
rect 474292 203010 474298 203012
rect 475510 203010 475516 203012
rect 474181 202952 474186 203008
rect 473004 202948 473010 202950
rect 474181 202948 474228 202952
rect 474292 202950 474338 203010
rect 475470 202950 475516 203010
rect 475580 203008 475627 203012
rect 475622 202952 475627 203008
rect 474292 202948 474298 202950
rect 475510 202948 475516 202950
rect 475580 202948 475627 202952
rect 471789 202947 471855 202948
rect 472893 202947 472959 202948
rect 474181 202947 474247 202948
rect 475561 202947 475627 202948
rect 476113 203010 476179 203013
rect 476430 203010 476436 203012
rect 476113 203008 476436 203010
rect 476113 202952 476118 203008
rect 476174 202952 476436 203008
rect 476113 202950 476436 202952
rect 476113 202947 476179 202950
rect 476430 202948 476436 202950
rect 476500 202948 476506 203012
rect 478873 203010 478939 203013
rect 479926 203010 479932 203012
rect 478873 203008 479932 203010
rect 478873 202952 478878 203008
rect 478934 202952 479932 203008
rect 478873 202950 479932 202952
rect 478873 202947 478939 202950
rect 479926 202948 479932 202950
rect 479996 202948 480002 203012
rect 480621 203010 480687 203013
rect 481214 203010 481220 203012
rect 480621 203008 481220 203010
rect 480621 202952 480626 203008
rect 480682 202952 481220 203008
rect 480621 202950 481220 202952
rect 480621 202947 480687 202950
rect 481214 202948 481220 202950
rect 481284 202948 481290 203012
rect 481633 203010 481699 203013
rect 482134 203010 482140 203012
rect 481633 203008 482140 203010
rect 481633 202952 481638 203008
rect 481694 202952 482140 203008
rect 481633 202950 482140 202952
rect 481633 202947 481699 202950
rect 482134 202948 482140 202950
rect 482204 202948 482210 203012
rect 483013 203010 483079 203013
rect 483422 203010 483428 203012
rect 483013 203008 483428 203010
rect 483013 202952 483018 203008
rect 483074 202952 483428 203008
rect 483013 202950 483428 202952
rect 483013 202947 483079 202950
rect 483422 202948 483428 202950
rect 483492 202948 483498 203012
rect 484393 203010 484459 203013
rect 539961 203012 540027 203013
rect 484710 203010 484716 203012
rect 484393 203008 484716 203010
rect 484393 202952 484398 203008
rect 484454 202952 484716 203008
rect 484393 202950 484716 202952
rect 484393 202947 484459 202950
rect 484710 202948 484716 202950
rect 484780 202948 484786 203012
rect 539910 203010 539916 203012
rect 539870 202950 539916 203010
rect 539980 203008 540027 203012
rect 540022 202952 540027 203008
rect 539910 202948 539916 202950
rect 539980 202948 540027 202952
rect 539961 202947 540027 202948
rect 342294 201724 342300 201788
rect 342364 201724 342370 201788
rect 342302 201516 342362 201724
rect 448421 201516 448487 201517
rect 342270 201452 342276 201516
rect 342340 201454 342362 201516
rect 448378 201514 448384 201516
rect 448330 201454 448384 201514
rect 448448 201512 448487 201516
rect 448482 201456 448487 201512
rect 342340 201452 342346 201454
rect 448378 201452 448384 201454
rect 448448 201452 448487 201456
rect 448421 201451 448487 201452
rect 3969 201106 4035 201109
rect 538254 201106 538260 201108
rect 3969 201104 538260 201106
rect 3969 201048 3974 201104
rect 4030 201048 538260 201104
rect 3969 201046 538260 201048
rect 3969 201043 4035 201046
rect 538254 201044 538260 201046
rect 538324 201044 538330 201108
rect 3417 200970 3483 200973
rect 540278 200970 540284 200972
rect 3417 200968 540284 200970
rect 3417 200912 3422 200968
rect 3478 200912 540284 200968
rect 3417 200910 540284 200912
rect 3417 200907 3483 200910
rect 540278 200908 540284 200910
rect 540348 200908 540354 200972
rect 3785 200834 3851 200837
rect 543038 200834 543044 200836
rect 3785 200832 543044 200834
rect 3785 200776 3790 200832
rect 3846 200776 543044 200832
rect 3785 200774 543044 200776
rect 3785 200771 3851 200774
rect 543038 200772 543044 200774
rect 543108 200772 543114 200836
rect 3601 200698 3667 200701
rect 543222 200698 543228 200700
rect 3601 200696 543228 200698
rect 3601 200640 3606 200696
rect 3662 200640 543228 200696
rect 3601 200638 543228 200640
rect 3601 200635 3667 200638
rect 543222 200636 543228 200638
rect 543292 200636 543298 200700
rect 539910 196012 539916 196076
rect 539980 196012 539986 196076
rect 539918 195802 539978 196012
rect 540094 195802 540100 195804
rect 539918 195742 540100 195802
rect 540094 195740 540100 195742
rect 540164 195740 540170 195804
rect -960 193898 480 193988
rect 4061 193898 4127 193901
rect -960 193896 4127 193898
rect -960 193840 4066 193896
rect 4122 193840 4127 193896
rect -960 193838 4127 193840
rect -960 193748 480 193838
rect 4061 193835 4127 193838
rect 583520 193476 584960 193716
rect 539961 193218 540027 193221
rect 540094 193218 540100 193220
rect 539961 193216 540100 193218
rect 539961 193160 539966 193216
rect 540022 193160 540100 193216
rect 539961 193158 540100 193160
rect 539961 193155 540027 193158
rect 540094 193156 540100 193158
rect 540164 193156 540170 193220
rect 539961 183700 540027 183701
rect 539910 183698 539916 183700
rect 539870 183638 539916 183698
rect 539980 183696 540027 183700
rect 540022 183640 540027 183696
rect 539910 183636 539916 183638
rect 539980 183636 540027 183640
rect 539961 183635 540027 183636
rect 500309 183154 500375 183157
rect 497230 183152 500375 183154
rect 497230 183096 500314 183152
rect 500370 183096 500375 183152
rect 497230 183094 500375 183096
rect 379789 182746 379855 182749
rect 377814 182744 379855 182746
rect 377814 182722 379794 182744
rect 377292 182688 379794 182722
rect 379850 182688 379855 182744
rect 497230 182692 497290 183094
rect 500309 183091 500375 183094
rect 377292 182686 379855 182688
rect 377292 182662 377874 182686
rect 379789 182683 379855 182686
rect 580165 181930 580231 181933
rect 583520 181930 584960 182020
rect 580165 181928 584960 181930
rect 580165 181872 580170 181928
rect 580226 181872 584960 181928
rect 580165 181870 584960 181872
rect 580165 181867 580231 181870
rect 583520 181780 584960 181870
rect 496445 181386 496511 181389
rect 496445 181384 496554 181386
rect 496445 181328 496450 181384
rect 496506 181328 496554 181384
rect 496445 181323 496554 181328
rect 377292 180978 377874 181022
rect 496494 180992 496554 181323
rect 380433 180978 380499 180981
rect 377292 180976 380499 180978
rect 377292 180962 380438 180976
rect 377814 180920 380438 180962
rect 380494 180920 380499 180976
rect 377814 180918 380499 180920
rect 380433 180915 380499 180918
rect 417417 180570 417483 180573
rect 417417 180568 420378 180570
rect 417417 180512 417422 180568
rect 417478 180512 420378 180568
rect 417417 180510 420378 180512
rect 417417 180507 417483 180510
rect 297909 180298 297975 180301
rect 300166 180298 300226 180319
rect 297909 180296 300226 180298
rect 297909 180240 297914 180296
rect 297970 180240 300226 180296
rect 297909 180238 300226 180240
rect 297909 180235 297975 180238
rect -960 179482 480 179572
rect 3509 179482 3575 179485
rect -960 179480 3575 179482
rect -960 179424 3514 179480
rect 3570 179424 3575 179480
rect -960 179422 3575 179424
rect -960 179332 480 179422
rect 3509 179419 3575 179422
rect 297909 171866 297975 171869
rect 297909 171865 299674 171866
rect 300166 171865 300226 180238
rect 420318 171865 420378 180510
rect 539910 176700 539916 176764
rect 539980 176700 539986 176764
rect 539918 176490 539978 176700
rect 540094 176490 540100 176492
rect 539918 176430 540100 176490
rect 540094 176428 540100 176430
rect 540164 176428 540170 176492
rect 542997 173908 543063 173909
rect 542997 173904 543044 173908
rect 543108 173906 543114 173908
rect 542997 173848 543002 173904
rect 542997 173844 543044 173848
rect 543108 173846 543154 173906
rect 543108 173844 543114 173846
rect 542997 173843 543063 173844
rect 297909 171864 300226 171865
rect 297909 171808 297914 171864
rect 297970 171835 300226 171864
rect 420164 171835 420378 171865
rect 297970 171808 300196 171835
rect 297909 171806 300196 171808
rect 297909 171803 297975 171806
rect 299614 171805 300196 171806
rect 420134 171805 420348 171835
rect 418061 171730 418127 171733
rect 420134 171730 420194 171805
rect 418061 171728 420194 171730
rect 418061 171672 418066 171728
rect 418122 171672 420194 171728
rect 418061 171670 420194 171672
rect 418061 171667 418127 171670
rect 580165 170098 580231 170101
rect 583520 170098 584960 170188
rect 580165 170096 584960 170098
rect 580165 170040 580170 170096
rect 580226 170040 584960 170096
rect 580165 170038 584960 170040
rect 580165 170035 580231 170038
rect 583520 169948 584960 170038
rect 540145 167108 540211 167109
rect 540094 167044 540100 167108
rect 540164 167106 540211 167108
rect 540164 167104 540256 167106
rect 540206 167048 540256 167104
rect 540164 167046 540256 167048
rect 540164 167044 540211 167046
rect 540145 167043 540211 167044
rect -960 165066 480 165156
rect 3969 165066 4035 165069
rect -960 165064 4035 165066
rect -960 165008 3974 165064
rect 4030 165008 4035 165064
rect -960 165006 4035 165008
rect -960 164916 480 165006
rect 3969 165003 4035 165006
rect 540145 164252 540211 164253
rect 540094 164250 540100 164252
rect 540054 164190 540100 164250
rect 540164 164248 540211 164252
rect 540206 164192 540211 164248
rect 540094 164188 540100 164190
rect 540164 164188 540211 164192
rect 540145 164187 540211 164188
rect 542997 164252 543063 164253
rect 542997 164248 543044 164252
rect 543108 164250 543114 164252
rect 542997 164192 543002 164248
rect 542997 164188 543044 164192
rect 543108 164190 543154 164250
rect 543108 164188 543114 164190
rect 542997 164187 543063 164188
rect 539910 162692 539916 162756
rect 539980 162692 539986 162756
rect 539918 162621 539978 162692
rect 539918 162616 540027 162621
rect 539918 162560 539966 162616
rect 540022 162560 540027 162616
rect 539918 162558 540027 162560
rect 539961 162555 540027 162558
rect 579797 158402 579863 158405
rect 583520 158402 584960 158492
rect 579797 158400 584960 158402
rect 579797 158344 579802 158400
rect 579858 158344 584960 158400
rect 579797 158342 584960 158344
rect 579797 158339 579863 158342
rect 583520 158252 584960 158342
rect 539961 153234 540027 153237
rect 540094 153234 540100 153236
rect 539961 153232 540100 153234
rect 539961 153176 539966 153232
rect 540022 153176 540100 153232
rect 539961 153174 540100 153176
rect 539961 153171 540027 153174
rect 540094 153172 540100 153174
rect 540164 153172 540170 153236
rect -960 150786 480 150876
rect 3785 150786 3851 150789
rect -960 150784 3851 150786
rect -960 150728 3790 150784
rect 3846 150728 3851 150784
rect -960 150726 3851 150728
rect -960 150636 480 150726
rect 3785 150723 3851 150726
rect 539961 147794 540027 147797
rect 540094 147794 540100 147796
rect 539961 147792 540100 147794
rect 539961 147736 539966 147792
rect 540022 147736 540100 147792
rect 539961 147734 540100 147736
rect 539961 147731 540027 147734
rect 540094 147732 540100 147734
rect 540164 147732 540170 147796
rect 583520 146556 584960 146796
rect 539726 144876 539732 144940
rect 539796 144938 539802 144940
rect 539961 144938 540027 144941
rect 539796 144936 540027 144938
rect 539796 144880 539966 144936
rect 540022 144880 540027 144936
rect 539796 144878 540027 144880
rect 539796 144876 539802 144878
rect 539961 144875 540027 144878
rect -960 136370 480 136460
rect 3601 136370 3667 136373
rect -960 136368 3667 136370
rect -960 136312 3606 136368
rect 3662 136312 3667 136368
rect -960 136310 3667 136312
rect -960 136220 480 136310
rect 3601 136307 3667 136310
rect 580165 134874 580231 134877
rect 583520 134874 584960 134964
rect 580165 134872 584960 134874
rect 580165 134816 580170 134872
rect 580226 134816 584960 134872
rect 580165 134814 584960 134816
rect 580165 134811 580231 134814
rect 583520 134724 584960 134814
rect 379789 125626 379855 125629
rect 379973 125626 380039 125629
rect 379789 125624 380039 125626
rect 379789 125568 379794 125624
rect 379850 125568 379978 125624
rect 380034 125568 380039 125624
rect 379789 125566 380039 125568
rect 379789 125563 379855 125566
rect 379973 125563 380039 125566
rect 500125 123722 500191 123725
rect 497230 123720 500191 123722
rect 497230 123664 500130 123720
rect 500186 123664 500191 123720
rect 497230 123662 500191 123664
rect 380801 123178 380867 123181
rect 377814 123176 380867 123178
rect 377814 123174 380806 123176
rect 377292 123120 380806 123174
rect 380862 123120 380867 123176
rect 497230 123144 497290 123662
rect 500125 123659 500191 123662
rect 580165 123178 580231 123181
rect 583520 123178 584960 123268
rect 580165 123176 584960 123178
rect 377292 123118 380867 123120
rect 377292 123114 377874 123118
rect 380801 123115 380867 123118
rect 580165 123120 580170 123176
rect 580226 123120 584960 123176
rect 580165 123118 584960 123120
rect 580165 123115 580231 123118
rect 583520 123028 584960 123118
rect -960 122090 480 122180
rect 3417 122090 3483 122093
rect 380341 122090 380407 122093
rect 500033 122090 500099 122093
rect -960 122088 3483 122090
rect -960 122032 3422 122088
rect 3478 122032 3483 122088
rect -960 122030 3483 122032
rect -960 121940 480 122030
rect 3417 122027 3483 122030
rect 377078 122088 380407 122090
rect 377078 122032 380346 122088
rect 380402 122032 380407 122088
rect 377078 122030 380407 122032
rect 377078 121444 377138 122030
rect 380341 122027 380407 122030
rect 497230 122088 500099 122090
rect 497230 122032 500038 122088
rect 500094 122032 500099 122088
rect 497230 122030 500099 122032
rect 497230 121444 497290 122030
rect 500033 122027 500099 122030
rect 499941 120866 500007 120869
rect 497230 120864 500007 120866
rect 497230 120808 499946 120864
rect 500002 120808 500007 120864
rect 497230 120806 500007 120808
rect 377292 120322 377874 120346
rect 380249 120322 380315 120325
rect 377292 120320 380315 120322
rect 377292 120286 380254 120320
rect 377814 120264 380254 120286
rect 380310 120264 380315 120320
rect 497230 120316 497290 120806
rect 499941 120803 500007 120806
rect 539961 120732 540027 120733
rect 539910 120730 539916 120732
rect 539870 120670 539916 120730
rect 539980 120728 540027 120732
rect 540022 120672 540027 120728
rect 539910 120668 539916 120670
rect 539980 120668 540027 120672
rect 539961 120667 540027 120668
rect 377814 120262 380315 120264
rect 380249 120259 380315 120262
rect 379973 119234 380039 119237
rect 377078 119232 380039 119234
rect 377078 119176 379978 119232
rect 380034 119176 380039 119232
rect 377078 119174 380039 119176
rect 377078 118616 377138 119174
rect 379973 119171 380039 119174
rect 499849 118690 499915 118693
rect 497230 118688 499915 118690
rect 497230 118632 499854 118688
rect 499910 118632 499915 118688
rect 497230 118630 499915 118632
rect 497230 118616 497290 118630
rect 499849 118627 499915 118630
rect 380801 118146 380867 118149
rect 499757 118146 499823 118149
rect 377078 118144 380867 118146
rect 377078 118088 380806 118144
rect 380862 118088 380867 118144
rect 377078 118086 380867 118088
rect 377078 117488 377138 118086
rect 380801 118083 380867 118086
rect 497230 118144 499823 118146
rect 497230 118088 499762 118144
rect 499818 118088 499823 118144
rect 497230 118086 499823 118088
rect 497230 117488 497290 118086
rect 499757 118083 499823 118086
rect 539961 115970 540027 115973
rect 540094 115970 540100 115972
rect 539961 115968 540100 115970
rect 539961 115912 539966 115968
rect 540022 115912 540100 115968
rect 539961 115910 540100 115912
rect 539961 115907 540027 115910
rect 540094 115908 540100 115910
rect 540164 115908 540170 115972
rect 380801 115834 380867 115837
rect 499665 115834 499731 115837
rect 377814 115832 380867 115834
rect 377814 115818 380806 115832
rect 377292 115776 380806 115818
rect 380862 115776 380867 115832
rect 377292 115774 380867 115776
rect 497230 115832 499731 115834
rect 497230 115776 499670 115832
rect 499726 115776 499731 115832
rect 497230 115774 499731 115776
rect 377292 115758 377874 115774
rect 380801 115771 380867 115774
rect 499665 115771 499731 115774
rect 500217 115290 500283 115293
rect 497230 115288 500283 115290
rect 497230 115232 500222 115288
rect 500278 115232 500283 115288
rect 497230 115230 500283 115232
rect 380709 114746 380775 114749
rect 377814 114744 380775 114746
rect 377814 114690 380714 114744
rect 377292 114688 380714 114690
rect 380770 114688 380775 114744
rect 377292 114686 380775 114688
rect 377292 114630 377874 114686
rect 380709 114683 380775 114686
rect 497230 114660 497290 115230
rect 500217 115227 500283 115230
rect 297817 111754 297883 111757
rect 297817 111752 300778 111754
rect 297817 111696 297822 111752
rect 297878 111696 300778 111752
rect 297817 111694 300778 111696
rect 297817 111691 297883 111694
rect 300718 111349 300778 111694
rect 300718 111344 300827 111349
rect 300718 111288 300766 111344
rect 300822 111288 300827 111344
rect 300718 111286 300827 111288
rect 300761 111283 300827 111286
rect 416773 111346 416839 111349
rect 420134 111346 420194 111564
rect 579797 111482 579863 111485
rect 583520 111482 584960 111572
rect 579797 111480 584960 111482
rect 579797 111424 579802 111480
rect 579858 111424 584960 111480
rect 579797 111422 584960 111424
rect 579797 111419 579863 111422
rect 416773 111344 420194 111346
rect 416773 111288 416778 111344
rect 416834 111288 420194 111344
rect 583520 111332 584960 111422
rect 416773 111286 420194 111288
rect 416773 111283 416839 111286
rect 303613 109036 303679 109037
rect 303613 109032 303660 109036
rect 303724 109034 303730 109036
rect 307753 109034 307819 109037
rect 424225 109036 424291 109037
rect 308070 109034 308076 109036
rect 303613 108976 303618 109032
rect 303613 108972 303660 108976
rect 303724 108974 303770 109034
rect 307753 109032 308076 109034
rect 307753 108976 307758 109032
rect 307814 108976 308076 109032
rect 307753 108974 308076 108976
rect 303724 108972 303730 108974
rect 303613 108971 303679 108972
rect 307753 108971 307819 108974
rect 308070 108972 308076 108974
rect 308140 108972 308146 109036
rect 424174 109034 424180 109036
rect 424134 108974 424180 109034
rect 424244 109032 424291 109036
rect 424286 108976 424291 109032
rect 424174 108972 424180 108974
rect 424244 108972 424291 108976
rect 424225 108971 424291 108972
rect 427813 109034 427879 109037
rect 428038 109034 428044 109036
rect 427813 109032 428044 109034
rect 427813 108976 427818 109032
rect 427874 108976 428044 109032
rect 427813 108974 428044 108976
rect 427813 108971 427879 108974
rect 428038 108972 428044 108974
rect 428108 108972 428114 109036
rect -960 107674 480 107764
rect 3233 107674 3299 107677
rect -960 107672 3299 107674
rect -960 107616 3238 107672
rect 3294 107616 3299 107672
rect -960 107614 3299 107616
rect -960 107524 480 107614
rect 3233 107611 3299 107614
rect 543181 106314 543247 106317
rect 543365 106314 543431 106317
rect 543181 106312 543431 106314
rect 543181 106256 543186 106312
rect 543242 106256 543370 106312
rect 543426 106256 543431 106312
rect 543181 106254 543431 106256
rect 543181 106251 543247 106254
rect 543365 106251 543431 106254
rect 583520 99636 584960 99876
rect 67582 93876 67588 93940
rect 67652 93938 67658 93940
rect 72417 93938 72483 93941
rect 67652 93936 72483 93938
rect 67652 93880 72422 93936
rect 72478 93880 72483 93936
rect 67652 93878 72483 93880
rect 67652 93876 67658 93878
rect 72417 93875 72483 93878
rect 86902 93876 86908 93940
rect 86972 93938 86978 93940
rect 91737 93938 91803 93941
rect 86972 93936 91803 93938
rect 86972 93880 91742 93936
rect 91798 93880 91803 93936
rect 86972 93878 91803 93880
rect 86972 93876 86978 93878
rect 91737 93875 91803 93878
rect 106222 93876 106228 93940
rect 106292 93938 106298 93940
rect 111057 93938 111123 93941
rect 106292 93936 111123 93938
rect 106292 93880 111062 93936
rect 111118 93880 111123 93936
rect 106292 93878 111123 93880
rect 106292 93876 106298 93878
rect 111057 93875 111123 93878
rect 125542 93876 125548 93940
rect 125612 93938 125618 93940
rect 130377 93938 130443 93941
rect 125612 93936 130443 93938
rect 125612 93880 130382 93936
rect 130438 93880 130443 93936
rect 125612 93878 130443 93880
rect 125612 93876 125618 93878
rect 130377 93875 130443 93878
rect 9622 93740 9628 93804
rect 9692 93802 9698 93804
rect 154481 93802 154547 93805
rect 9692 93742 19258 93802
rect 9692 93740 9698 93742
rect 19198 93530 19258 93742
rect 21958 93742 22202 93802
rect 21958 93530 22018 93742
rect 22142 93666 22202 93742
rect 60598 93742 60842 93802
rect 28942 93666 28948 93668
rect 22142 93606 28948 93666
rect 28942 93604 28948 93606
rect 29012 93604 29018 93668
rect 48129 93666 48195 93669
rect 48262 93666 48268 93668
rect 48129 93664 48268 93666
rect 48129 93608 48134 93664
rect 48190 93608 48268 93664
rect 48129 93606 48268 93608
rect 48129 93603 48195 93606
rect 48262 93604 48268 93606
rect 48332 93604 48338 93668
rect 38653 93530 38719 93533
rect 19198 93470 22018 93530
rect 38518 93528 38719 93530
rect 38518 93472 38658 93528
rect 38714 93472 38719 93528
rect 38518 93470 38719 93472
rect 9622 93394 9628 93396
rect -960 93258 480 93348
rect 4846 93334 9628 93394
rect 4846 93258 4906 93334
rect 9622 93332 9628 93334
rect 9692 93332 9698 93396
rect -960 93198 4906 93258
rect -960 93108 480 93198
rect 28942 93196 28948 93260
rect 29012 93258 29018 93260
rect 38518 93258 38578 93470
rect 38653 93467 38719 93470
rect 57830 93468 57836 93532
rect 57900 93530 57906 93532
rect 60598 93530 60658 93742
rect 60782 93666 60842 93742
rect 79918 93742 80162 93802
rect 67582 93666 67588 93668
rect 60782 93606 67588 93666
rect 67582 93604 67588 93606
rect 67652 93604 67658 93668
rect 72417 93666 72483 93669
rect 72417 93664 77218 93666
rect 72417 93608 72422 93664
rect 72478 93608 77218 93664
rect 72417 93606 77218 93608
rect 72417 93603 72483 93606
rect 57900 93470 60658 93530
rect 77158 93530 77218 93606
rect 79918 93530 79978 93742
rect 80102 93666 80162 93742
rect 99238 93742 99482 93802
rect 86902 93666 86908 93668
rect 80102 93606 86908 93666
rect 86902 93604 86908 93606
rect 86972 93604 86978 93668
rect 91737 93666 91803 93669
rect 91737 93664 96538 93666
rect 91737 93608 91742 93664
rect 91798 93608 96538 93664
rect 91737 93606 96538 93608
rect 91737 93603 91803 93606
rect 77158 93470 79978 93530
rect 96478 93530 96538 93606
rect 99238 93530 99298 93742
rect 99422 93666 99482 93742
rect 118558 93742 118802 93802
rect 106222 93666 106228 93668
rect 99422 93606 106228 93666
rect 106222 93604 106228 93606
rect 106292 93604 106298 93668
rect 111057 93666 111123 93669
rect 111057 93664 115858 93666
rect 111057 93608 111062 93664
rect 111118 93608 115858 93664
rect 111057 93606 115858 93608
rect 111057 93603 111123 93606
rect 96478 93470 99298 93530
rect 115798 93530 115858 93606
rect 118558 93530 118618 93742
rect 118742 93666 118802 93742
rect 154481 93800 161490 93802
rect 154481 93744 154486 93800
rect 154542 93744 161490 93800
rect 154481 93742 161490 93744
rect 154481 93739 154547 93742
rect 125542 93666 125548 93668
rect 118742 93606 125548 93666
rect 125542 93604 125548 93606
rect 125612 93604 125618 93668
rect 130377 93666 130443 93669
rect 140037 93666 140103 93669
rect 144913 93666 144979 93669
rect 130377 93664 135178 93666
rect 130377 93608 130382 93664
rect 130438 93608 135178 93664
rect 130377 93606 135178 93608
rect 130377 93603 130443 93606
rect 115798 93470 118618 93530
rect 135118 93530 135178 93606
rect 140037 93664 144979 93666
rect 140037 93608 140042 93664
rect 140098 93608 144918 93664
rect 144974 93608 144979 93664
rect 140037 93606 144979 93608
rect 140037 93603 140103 93606
rect 144913 93603 144979 93606
rect 161430 93530 161490 93742
rect 170998 93742 180810 93802
rect 170998 93530 171058 93742
rect 135118 93470 135362 93530
rect 161430 93470 171058 93530
rect 180750 93530 180810 93742
rect 190318 93742 200130 93802
rect 190318 93530 190378 93742
rect 180750 93470 190378 93530
rect 200070 93530 200130 93742
rect 209638 93742 219450 93802
rect 209638 93530 209698 93742
rect 200070 93470 209698 93530
rect 219390 93530 219450 93742
rect 228958 93742 238770 93802
rect 228958 93530 229018 93742
rect 219390 93470 229018 93530
rect 238710 93530 238770 93742
rect 248278 93742 258090 93802
rect 248278 93530 248338 93742
rect 238710 93470 248338 93530
rect 258030 93530 258090 93742
rect 267598 93742 277410 93802
rect 267598 93530 267658 93742
rect 258030 93470 267658 93530
rect 277350 93530 277410 93742
rect 286918 93742 296730 93802
rect 286918 93530 286978 93742
rect 277350 93470 286978 93530
rect 296670 93530 296730 93742
rect 306238 93742 316050 93802
rect 306238 93530 306298 93742
rect 296670 93470 306298 93530
rect 315990 93530 316050 93742
rect 325558 93742 335370 93802
rect 325558 93530 325618 93742
rect 315990 93470 325618 93530
rect 335310 93530 335370 93742
rect 344878 93742 354690 93802
rect 344878 93530 344938 93742
rect 335310 93470 344938 93530
rect 354630 93530 354690 93742
rect 364198 93742 374010 93802
rect 364198 93530 364258 93742
rect 354630 93470 364258 93530
rect 373950 93530 374010 93742
rect 383518 93742 393330 93802
rect 383518 93530 383578 93742
rect 373950 93470 383578 93530
rect 393270 93530 393330 93742
rect 402838 93742 412650 93802
rect 402838 93530 402898 93742
rect 393270 93470 402898 93530
rect 412590 93530 412650 93742
rect 422158 93742 431970 93802
rect 422158 93530 422218 93742
rect 412590 93470 422218 93530
rect 431910 93530 431970 93742
rect 441478 93742 451290 93802
rect 441478 93530 441538 93742
rect 431910 93470 441538 93530
rect 451230 93530 451290 93742
rect 460798 93742 470610 93802
rect 460798 93530 460858 93742
rect 451230 93470 460858 93530
rect 470550 93530 470610 93742
rect 480118 93742 489930 93802
rect 480118 93530 480178 93742
rect 470550 93470 480178 93530
rect 489870 93530 489930 93742
rect 499438 93742 509250 93802
rect 499438 93530 499498 93742
rect 489870 93470 499498 93530
rect 509190 93530 509250 93742
rect 518758 93742 528570 93802
rect 518758 93530 518818 93742
rect 509190 93470 518818 93530
rect 528510 93530 528570 93742
rect 540094 93530 540100 93532
rect 528510 93470 540100 93530
rect 57900 93468 57906 93470
rect 29012 93198 38578 93258
rect 29012 93196 29018 93198
rect 48262 93196 48268 93260
rect 48332 93258 48338 93260
rect 57830 93258 57836 93260
rect 48332 93198 57836 93258
rect 48332 93196 48338 93198
rect 57830 93196 57836 93198
rect 57900 93196 57906 93260
rect 135302 93258 135362 93470
rect 540094 93468 540100 93470
rect 540164 93468 540170 93532
rect 140037 93258 140103 93261
rect 135302 93256 140103 93258
rect 135302 93200 140042 93256
rect 140098 93200 140103 93256
rect 135302 93198 140103 93200
rect 140037 93195 140103 93198
rect 580165 87954 580231 87957
rect 583520 87954 584960 88044
rect 580165 87952 584960 87954
rect 580165 87896 580170 87952
rect 580226 87896 584960 87952
rect 580165 87894 584960 87896
rect 580165 87891 580231 87894
rect 583520 87804 584960 87894
rect 3417 80066 3483 80069
rect 542854 80066 542860 80068
rect 3417 80064 542860 80066
rect 3417 80008 3422 80064
rect 3478 80008 542860 80064
rect 3417 80006 542860 80008
rect 3417 80003 3483 80006
rect 542854 80004 542860 80006
rect 542924 80004 542930 80068
rect -960 78978 480 79068
rect 3417 78978 3483 78981
rect -960 78976 3483 78978
rect -960 78920 3422 78976
rect 3478 78920 3483 78976
rect -960 78918 3483 78920
rect -960 78828 480 78918
rect 3417 78915 3483 78918
rect 542905 77210 542971 77213
rect 543181 77210 543247 77213
rect 542905 77208 543247 77210
rect 542905 77152 542910 77208
rect 542966 77152 543186 77208
rect 543242 77152 543247 77208
rect 542905 77150 543247 77152
rect 542905 77147 542971 77150
rect 543181 77147 543247 77150
rect 580165 76258 580231 76261
rect 583520 76258 584960 76348
rect 580165 76256 584960 76258
rect 580165 76200 580170 76256
rect 580226 76200 584960 76256
rect 580165 76198 584960 76200
rect 580165 76195 580231 76198
rect 583520 76108 584960 76198
rect 541566 64834 541572 64836
rect 614 64774 541572 64834
rect -960 64562 480 64652
rect 614 64562 674 64774
rect 541566 64772 541572 64774
rect 541636 64772 541642 64836
rect -960 64502 674 64562
rect 579797 64562 579863 64565
rect 583520 64562 584960 64652
rect 579797 64560 584960 64562
rect 579797 64504 579802 64560
rect 579858 64504 584960 64560
rect 579797 64502 584960 64504
rect -960 64412 480 64502
rect 579797 64499 579863 64502
rect 583520 64412 584960 64502
rect 583520 52716 584960 52956
rect 3325 50962 3391 50965
rect 539542 50962 539548 50964
rect 3325 50960 539548 50962
rect 3325 50904 3330 50960
rect 3386 50904 539548 50960
rect 3325 50902 539548 50904
rect 3325 50899 3391 50902
rect 539542 50900 539548 50902
rect 539612 50900 539618 50964
rect -960 50146 480 50236
rect 3325 50146 3391 50149
rect -960 50144 3391 50146
rect -960 50088 3330 50144
rect 3386 50088 3391 50144
rect -960 50086 3391 50088
rect -960 49996 480 50086
rect 3325 50083 3391 50086
rect 580165 41034 580231 41037
rect 583520 41034 584960 41124
rect 580165 41032 584960 41034
rect 580165 40976 580170 41032
rect 580226 40976 584960 41032
rect 580165 40974 584960 40976
rect 580165 40971 580231 40974
rect 583520 40884 584960 40974
rect -960 35866 480 35956
rect 542670 35866 542676 35868
rect -960 35806 542676 35866
rect -960 35716 480 35806
rect 542670 35804 542676 35806
rect 542740 35804 542746 35868
rect 580165 29338 580231 29341
rect 583520 29338 584960 29428
rect 580165 29336 584960 29338
rect 580165 29280 580170 29336
rect 580226 29280 584960 29336
rect 580165 29278 584960 29280
rect 580165 29275 580231 29278
rect 583520 29188 584960 29278
rect 542486 21994 542492 21996
rect 614 21934 542492 21994
rect -960 21450 480 21540
rect 614 21450 674 21934
rect 542486 21932 542492 21934
rect 542556 21932 542562 21996
rect -960 21390 674 21450
rect -960 21300 480 21390
rect 579797 17642 579863 17645
rect 583520 17642 584960 17732
rect 579797 17640 584960 17642
rect 579797 17584 579802 17640
rect 579858 17584 584960 17640
rect 579797 17582 584960 17584
rect 579797 17579 579863 17582
rect 583520 17492 584960 17582
rect 3417 8258 3483 8261
rect 542302 8258 542308 8260
rect 3417 8256 542308 8258
rect 3417 8200 3422 8256
rect 3478 8200 542308 8256
rect 3417 8198 542308 8200
rect 3417 8195 3483 8198
rect 542302 8196 542308 8198
rect 542372 8196 542378 8260
rect -960 7170 480 7260
rect 3417 7170 3483 7173
rect -960 7168 3483 7170
rect -960 7112 3422 7168
rect 3478 7112 3483 7168
rect -960 7110 3483 7112
rect -960 7020 480 7110
rect 3417 7107 3483 7110
rect 583520 5796 584960 6036
<< via3 >>
rect 538260 700708 538324 700772
rect 538444 700572 538508 700636
rect 540100 700436 540164 700500
rect 539916 700300 539980 700364
rect 538812 623732 538876 623796
rect 373580 612776 373644 612780
rect 373580 612720 373630 612776
rect 373630 612720 373644 612776
rect 373580 612716 373644 612720
rect 488580 612776 488644 612780
rect 488580 612720 488594 612776
rect 488594 612720 488644 612776
rect 488580 612716 488644 612720
rect 493916 612776 493980 612780
rect 493916 612720 493966 612776
rect 493966 612720 493980 612776
rect 493916 612716 493980 612720
rect 369164 610948 369228 611012
rect 373028 610948 373092 611012
rect 427968 519692 428032 519756
rect 433808 519692 433872 519756
rect 313780 518740 313844 518804
rect 319668 518740 319732 518804
rect 323532 518740 323596 518804
rect 324268 518800 324332 518804
rect 324268 518744 324318 518800
rect 324318 518744 324332 518800
rect 324268 518740 324332 518744
rect 325188 518740 325252 518804
rect 326476 518800 326540 518804
rect 326476 518744 326490 518800
rect 326490 518744 326540 518800
rect 326476 518740 326540 518744
rect 327396 518800 327460 518804
rect 327396 518744 327410 518800
rect 327410 518744 327460 518800
rect 327396 518740 327460 518744
rect 328868 518800 328932 518804
rect 328868 518744 328918 518800
rect 328918 518744 328932 518800
rect 328868 518740 328932 518744
rect 330156 518800 330220 518804
rect 330156 518744 330170 518800
rect 330170 518744 330220 518800
rect 330156 518740 330220 518744
rect 331628 518740 331692 518804
rect 332364 518800 332428 518804
rect 332364 518744 332414 518800
rect 332414 518744 332428 518800
rect 332364 518740 332428 518744
rect 333652 518740 333716 518804
rect 334572 518740 334636 518804
rect 335860 518800 335924 518804
rect 335860 518744 335874 518800
rect 335874 518744 335924 518800
rect 335860 518740 335924 518744
rect 336964 518800 337028 518804
rect 336964 518744 336978 518800
rect 336978 518744 337028 518800
rect 336964 518740 337028 518744
rect 338068 518800 338132 518804
rect 338068 518744 338118 518800
rect 338118 518744 338132 518800
rect 338068 518740 338132 518744
rect 339540 518800 339604 518804
rect 339540 518744 339554 518800
rect 339554 518744 339604 518800
rect 339540 518740 339604 518744
rect 340460 518740 340524 518804
rect 341564 518800 341628 518804
rect 341564 518744 341578 518800
rect 341578 518744 341628 518800
rect 341564 518740 341628 518744
rect 345060 518740 345124 518804
rect 346532 518800 346596 518804
rect 346532 518744 346582 518800
rect 346582 518744 346596 518800
rect 346532 518740 346596 518744
rect 348924 518800 348988 518804
rect 348924 518744 348974 518800
rect 348974 518744 348988 518800
rect 348924 518740 348988 518744
rect 443132 518800 443196 518804
rect 443132 518744 443182 518800
rect 443182 518744 443196 518800
rect 443132 518740 443196 518744
rect 451228 518800 451292 518804
rect 451228 518744 451278 518800
rect 451278 518744 451292 518800
rect 451228 518740 451292 518744
rect 452516 518800 452580 518804
rect 452516 518744 452566 518800
rect 452566 518744 452580 518800
rect 452516 518740 452580 518744
rect 458404 518800 458468 518804
rect 458404 518744 458418 518800
rect 458418 518744 458468 518800
rect 458404 518740 458468 518744
rect 460428 518740 460492 518804
rect 466500 518800 466564 518804
rect 466500 518744 466514 518800
rect 466514 518744 466564 518800
rect 466500 518740 466564 518744
rect 312492 518604 312556 518668
rect 316172 518604 316236 518668
rect 318564 518604 318628 518668
rect 320772 518604 320836 518668
rect 323164 518664 323228 518668
rect 323164 518608 323178 518664
rect 323178 518608 323228 518664
rect 323164 518604 323228 518608
rect 331260 518604 331324 518668
rect 340644 518604 340708 518668
rect 347636 518664 347700 518668
rect 347636 518608 347686 518664
rect 347686 518608 347700 518664
rect 347636 518604 347700 518608
rect 429700 518604 429764 518668
rect 441660 518604 441724 518668
rect 444052 518604 444116 518668
rect 445340 518664 445404 518668
rect 445340 518608 445390 518664
rect 445390 518608 445404 518664
rect 445340 518604 445404 518608
rect 446628 518604 446692 518668
rect 457116 518664 457180 518668
rect 457116 518608 457130 518664
rect 457130 518608 457180 518664
rect 457116 518604 457180 518608
rect 461164 518604 461228 518668
rect 315068 518468 315132 518532
rect 316540 518468 316604 518532
rect 317276 518528 317340 518532
rect 317276 518472 317326 518528
rect 317326 518472 317340 518528
rect 317276 518468 317340 518472
rect 318564 518468 318628 518532
rect 321692 518468 321756 518532
rect 330340 518468 330404 518532
rect 343036 518528 343100 518532
rect 343036 518472 343050 518528
rect 343050 518472 343100 518528
rect 343036 518468 343100 518472
rect 348924 518468 348988 518532
rect 426572 518468 426636 518532
rect 443868 518468 443932 518532
rect 444972 518468 445036 518532
rect 447732 518468 447796 518532
rect 448836 518468 448900 518532
rect 453620 518468 453684 518532
rect 454724 518468 454788 518532
rect 456012 518528 456076 518532
rect 456012 518472 456062 518528
rect 456062 518472 456076 518528
rect 456012 518468 456076 518472
rect 462452 518468 462516 518532
rect 463924 518468 463988 518532
rect 467420 518468 467484 518532
rect 313964 518332 314028 518396
rect 320956 518332 321020 518396
rect 337332 518332 337396 518396
rect 338436 518332 338500 518396
rect 339908 518332 339972 518396
rect 343772 518392 343836 518396
rect 343772 518336 343786 518392
rect 343786 518336 343836 518392
rect 343772 518332 343836 518336
rect 430804 518332 430868 518396
rect 435036 518332 435100 518396
rect 445524 518392 445588 518396
rect 445524 518336 445574 518392
rect 445574 518336 445588 518392
rect 445524 518332 445588 518336
rect 446996 518392 447060 518396
rect 446996 518336 447046 518392
rect 447046 518336 447060 518392
rect 446996 518332 447060 518336
rect 450124 518392 450188 518396
rect 450124 518336 450174 518392
rect 450174 518336 450188 518392
rect 450124 518332 450188 518336
rect 459508 518392 459572 518396
rect 459508 518336 459558 518392
rect 459558 518336 459572 518392
rect 459508 518332 459572 518336
rect 465212 518332 465276 518396
rect 303660 518256 303724 518260
rect 303660 518200 303674 518256
rect 303674 518200 303724 518256
rect 303660 518196 303724 518200
rect 322060 518196 322124 518260
rect 333836 518196 333900 518260
rect 341932 518196 341996 518260
rect 423812 518196 423876 518260
rect 429148 518256 429212 518260
rect 429148 518200 429198 518256
rect 429198 518200 429212 518256
rect 429148 518196 429212 518200
rect 436140 518196 436204 518260
rect 440740 518196 440804 518260
rect 448284 518256 448348 518260
rect 448284 518200 448334 518256
rect 448334 518200 448348 518256
rect 448284 518196 448348 518200
rect 468524 518196 468588 518260
rect 314700 518060 314764 518124
rect 320036 518060 320100 518124
rect 317460 517984 317524 517988
rect 317460 517928 317474 517984
rect 317474 517928 317524 517984
rect 317460 517924 317524 517928
rect 312676 517788 312740 517852
rect 334940 517788 335004 517852
rect 343404 517788 343468 517852
rect 347820 517848 347884 517852
rect 347820 517792 347870 517848
rect 347870 517792 347884 517848
rect 347820 517788 347884 517792
rect 432644 517848 432708 517852
rect 432644 517792 432658 517848
rect 432658 517792 432708 517848
rect 432644 517788 432708 517792
rect 437244 517848 437308 517852
rect 437244 517792 437294 517848
rect 437294 517792 437308 517848
rect 437244 517788 437308 517792
rect 309732 517652 309796 517716
rect 324452 517712 324516 517716
rect 324452 517656 324502 517712
rect 324502 517656 324516 517712
rect 324452 517652 324516 517656
rect 326660 517652 326724 517716
rect 327948 517652 328012 517716
rect 329052 517652 329116 517716
rect 332548 517712 332612 517716
rect 332548 517656 332598 517712
rect 332598 517656 332612 517712
rect 332548 517652 332612 517656
rect 336044 517652 336108 517716
rect 344324 517652 344388 517716
rect 345428 517652 345492 517716
rect 346716 517652 346780 517716
rect 433012 517652 433076 517716
rect 433932 517652 433996 517716
rect 435772 517652 435836 517716
rect 436876 517652 436940 517716
rect 437980 517652 438044 517716
rect 453252 517652 453316 517716
rect 460244 517652 460308 517716
rect 468340 517652 468404 517716
rect 307340 517516 307404 517580
rect 308628 517516 308692 517580
rect 310284 517576 310348 517580
rect 310284 517520 310334 517576
rect 310334 517520 310348 517576
rect 310284 517516 310348 517520
rect 311756 517576 311820 517580
rect 311756 517520 311806 517576
rect 311806 517520 311820 517576
rect 311756 517516 311820 517520
rect 325556 517516 325620 517580
rect 438348 517516 438412 517580
rect 438716 517576 438780 517580
rect 438716 517520 438766 517576
rect 438766 517520 438780 517576
rect 438716 517516 438780 517520
rect 439636 517516 439700 517580
rect 440004 517516 440068 517580
rect 441476 517576 441540 517580
rect 441476 517520 441526 517576
rect 441526 517520 441540 517576
rect 441476 517516 441540 517520
rect 442764 517516 442828 517580
rect 449756 517576 449820 517580
rect 449756 517520 449806 517576
rect 449806 517520 449820 517576
rect 449756 517516 449820 517520
rect 450860 517516 450924 517580
rect 451964 517516 452028 517580
rect 453804 517516 453868 517580
rect 455276 517576 455340 517580
rect 455276 517520 455326 517576
rect 455326 517520 455340 517576
rect 455276 517516 455340 517520
rect 456380 517516 456444 517580
rect 457852 517516 457916 517580
rect 459140 517516 459204 517580
rect 460796 517576 460860 517580
rect 460796 517520 460810 517576
rect 460810 517520 460860 517576
rect 460796 517516 460860 517520
rect 462084 517516 462148 517580
rect 463556 517576 463620 517580
rect 463556 517520 463606 517576
rect 463606 517520 463620 517576
rect 463556 517516 463620 517520
rect 464844 517516 464908 517580
rect 466132 517516 466196 517580
rect 467236 517516 467300 517580
rect 469076 517576 469140 517580
rect 469076 517520 469126 517576
rect 469126 517520 469140 517576
rect 469076 517516 469140 517520
rect 433932 495484 433996 495548
rect 433932 492688 433996 492692
rect 433932 492632 433946 492688
rect 433946 492632 433996 492688
rect 433932 492628 433996 492632
rect 542492 478892 542556 478956
rect 542308 476852 542372 476916
rect 542676 474676 542740 474740
rect 541572 472636 541636 472700
rect 539548 469916 539612 469980
rect 542860 468420 542924 468484
rect 539732 463660 539796 463724
rect 540284 462028 540348 462092
rect 543044 459988 543108 460052
rect 543228 457812 543292 457876
rect 539364 455228 539428 455292
rect 539732 451964 539796 452028
rect 540468 451964 540532 452028
rect 539364 451148 539428 451212
rect 539732 451148 539796 451212
rect 539364 442580 539428 442644
rect 539364 442172 539428 442236
rect 539732 442444 539796 442508
rect 539732 442308 539796 442372
rect 540468 442308 540532 442372
rect 539732 432652 539796 432716
rect 540468 432652 540532 432716
rect 539548 418372 539612 418436
rect 539364 414972 539428 415036
rect 539364 414428 539428 414492
rect 539732 414428 539796 414492
rect 539364 413748 539428 413812
rect 539732 413340 539796 413404
rect 540468 413340 540532 413404
rect 539548 406464 539612 406468
rect 539548 406408 539562 406464
rect 539562 406408 539612 406464
rect 539548 406404 539612 406408
rect 539364 405724 539428 405788
rect 539732 403684 539796 403748
rect 540468 403684 540532 403748
rect 539364 402188 539428 402252
rect 539364 399468 539428 399532
rect 543412 399528 543476 399532
rect 543412 399472 543462 399528
rect 543462 399472 543476 399528
rect 543412 399468 543476 399472
rect 539548 399060 539612 399124
rect 539548 398516 539612 398580
rect 539364 395388 539428 395452
rect 539364 391308 539428 391372
rect 540100 390492 540164 390556
rect 543412 389056 543476 389060
rect 543412 389000 543462 389056
rect 543462 389000 543476 389056
rect 543412 388996 543476 389000
rect 539364 388588 539428 388652
rect 539364 388452 539428 388516
rect 539732 388452 539796 388516
rect 539916 388452 539980 388516
rect 539364 384508 539428 384572
rect 539364 383420 539428 383484
rect 539732 383420 539796 383484
rect 539732 380972 539796 381036
rect 540468 380972 540532 381036
rect 543412 376680 543476 376684
rect 543412 376624 543426 376680
rect 543426 376624 543476 376680
rect 543412 376620 543476 376624
rect 539364 376348 539428 376412
rect 539732 376348 539796 376412
rect 539364 376212 539428 376276
rect 539364 374580 539428 374644
rect 539732 374580 539796 374644
rect 539732 373220 539796 373284
rect 543412 369744 543476 369748
rect 543412 369688 543462 369744
rect 543462 369688 543476 369744
rect 543412 369684 543476 369688
rect 539364 364108 539428 364172
rect 539732 364108 539796 364172
rect 539548 359484 539612 359548
rect 539548 359348 539612 359412
rect 543412 357368 543476 357372
rect 543412 357312 543426 357368
rect 543426 357312 543476 357368
rect 543412 357308 543476 357312
rect 543412 350432 543476 350436
rect 543412 350376 543462 350432
rect 543462 350376 543476 350432
rect 543412 350372 543476 350376
rect 539732 349012 539796 349076
rect 539916 331196 539980 331260
rect 539916 302364 539980 302428
rect 540100 302092 540164 302156
rect 539364 292768 539428 292772
rect 539364 292712 539378 292768
rect 539378 292712 539428 292768
rect 539364 292708 539428 292712
rect 539364 292088 539428 292092
rect 539364 292032 539378 292088
rect 539378 292032 539428 292088
rect 539364 292028 539428 292032
rect 540100 291892 540164 291956
rect 539364 286648 539428 286652
rect 539364 286592 539378 286648
rect 539378 286592 539428 286648
rect 539364 286588 539428 286592
rect 540100 279108 540164 279172
rect 540100 273396 540164 273460
rect 539364 265024 539428 265028
rect 539364 264968 539378 265024
rect 539378 264968 539428 265024
rect 539364 264964 539428 264968
rect 539732 265024 539796 265028
rect 539732 264968 539782 265024
rect 539782 264968 539796 265024
rect 539732 264964 539796 264968
rect 539732 263604 539796 263668
rect 539916 263468 539980 263532
rect 539364 256804 539428 256868
rect 539364 256668 539428 256732
rect 538996 240756 539060 240820
rect 538444 227700 538508 227764
rect 538628 227700 538692 227764
rect 538628 222804 538692 222868
rect 540100 216004 540164 216068
rect 474044 207708 474108 207772
rect 538260 205456 538324 205460
rect 538260 205400 538310 205456
rect 538310 205400 538324 205456
rect 538260 205396 538324 205400
rect 359228 204172 359292 204236
rect 366036 204172 366100 204236
rect 371004 204172 371068 204236
rect 456564 204232 456628 204236
rect 456564 204176 456614 204232
rect 456614 204176 456628 204232
rect 456564 204172 456628 204176
rect 468156 204172 468220 204236
rect 470364 204172 470428 204236
rect 477540 204232 477604 204236
rect 477540 204176 477554 204232
rect 477554 204176 477604 204232
rect 477540 204172 477604 204176
rect 479196 204172 479260 204236
rect 481772 204172 481836 204236
rect 490236 204232 490300 204236
rect 490236 204176 490250 204232
rect 490250 204176 490300 204232
rect 490236 204172 490300 204176
rect 360332 204036 360396 204100
rect 367508 204036 367572 204100
rect 449388 204036 449452 204100
rect 467052 204036 467116 204100
rect 469260 204036 469324 204100
rect 476252 204036 476316 204100
rect 478092 204036 478156 204100
rect 485820 204096 485884 204100
rect 485820 204040 485834 204096
rect 485834 204040 485884 204096
rect 485820 204036 485884 204040
rect 361620 203900 361684 203964
rect 366404 203900 366468 203964
rect 480484 203960 480548 203964
rect 480484 203904 480498 203960
rect 480498 203904 480548 203960
rect 480484 203900 480548 203904
rect 362908 203764 362972 203828
rect 364380 203824 364444 203828
rect 364380 203768 364394 203824
rect 364394 203768 364444 203824
rect 364380 203764 364444 203768
rect 448284 203764 448348 203828
rect 328132 203628 328196 203692
rect 329420 203628 329484 203692
rect 330708 203628 330772 203692
rect 334940 203628 335004 203692
rect 342852 203628 342916 203692
rect 343956 203628 344020 203692
rect 349108 203688 349172 203692
rect 349108 203632 349158 203688
rect 349158 203632 349172 203688
rect 349108 203628 349172 203632
rect 351132 203688 351196 203692
rect 351132 203632 351146 203688
rect 351146 203632 351196 203688
rect 351132 203628 351196 203632
rect 483060 203688 483124 203692
rect 483060 203632 483074 203688
rect 483074 203632 483124 203688
rect 340092 203492 340156 203556
rect 340828 203552 340892 203556
rect 483060 203628 483124 203632
rect 487476 203628 487540 203692
rect 340828 203496 340878 203552
rect 340878 203496 340892 203552
rect 340828 203492 340892 203496
rect 328316 203416 328380 203420
rect 328316 203360 328366 203416
rect 328366 203360 328380 203416
rect 328316 203356 328380 203360
rect 332364 203416 332428 203420
rect 332364 203360 332414 203416
rect 332414 203360 332428 203416
rect 332364 203356 332428 203360
rect 332916 203356 332980 203420
rect 336596 203416 336660 203420
rect 336596 203360 336646 203416
rect 336646 203360 336660 203416
rect 336596 203356 336660 203360
rect 338252 203356 338316 203420
rect 357388 203416 357452 203420
rect 357388 203360 357438 203416
rect 357438 203360 357452 203416
rect 357388 203356 357452 203360
rect 449572 203356 449636 203420
rect 450860 203356 450924 203420
rect 452148 203356 452212 203420
rect 453252 203416 453316 203420
rect 453252 203360 453302 203416
rect 453302 203360 453316 203416
rect 453252 203356 453316 203360
rect 456012 203356 456076 203420
rect 458772 203356 458836 203420
rect 460980 203356 461044 203420
rect 462268 203356 462332 203420
rect 478644 203356 478708 203420
rect 331076 203280 331140 203284
rect 331076 203224 331126 203280
rect 331126 203224 331140 203280
rect 331076 203220 331140 203224
rect 331628 203220 331692 203284
rect 334020 203280 334084 203284
rect 334020 203224 334034 203280
rect 334034 203224 334084 203280
rect 334020 203220 334084 203224
rect 336228 203220 336292 203284
rect 336964 203220 337028 203284
rect 339540 203280 339604 203284
rect 339540 203224 339554 203280
rect 339554 203224 339604 203280
rect 339540 203220 339604 203224
rect 345244 203220 345308 203284
rect 349844 203220 349908 203284
rect 368612 203220 368676 203284
rect 450676 203220 450740 203284
rect 452884 203220 452948 203284
rect 454908 203220 454972 203284
rect 455276 203280 455340 203284
rect 455276 203224 455290 203280
rect 455290 203224 455340 203280
rect 455276 203220 455340 203224
rect 457484 203220 457548 203284
rect 460060 203220 460124 203284
rect 463188 203220 463252 203284
rect 464660 203280 464724 203284
rect 464660 203224 464674 203280
rect 464674 203224 464724 203280
rect 464660 203220 464724 203224
rect 465948 203220 466012 203284
rect 471652 203220 471716 203284
rect 472756 203220 472820 203284
rect 475148 203220 475212 203284
rect 477724 203220 477788 203284
rect 484348 203552 484412 203556
rect 484348 203496 484398 203552
rect 484398 203496 484412 203552
rect 484348 203492 484412 203496
rect 488580 203492 488644 203556
rect 486372 203220 486436 203284
rect 329604 203084 329668 203148
rect 333652 203084 333716 203148
rect 334756 203084 334820 203148
rect 341748 203084 341812 203148
rect 346532 203084 346596 203148
rect 347820 203144 347884 203148
rect 347820 203088 347834 203144
rect 347834 203088 347884 203144
rect 347820 203084 347884 203088
rect 352788 203084 352852 203148
rect 353156 203144 353220 203148
rect 353156 203088 353206 203144
rect 353206 203088 353220 203144
rect 353156 203084 353220 203088
rect 354812 203084 354876 203148
rect 356100 203144 356164 203148
rect 356100 203088 356114 203144
rect 356114 203088 356164 203144
rect 356100 203084 356164 203088
rect 357756 203144 357820 203148
rect 357756 203088 357806 203144
rect 357806 203088 357820 203144
rect 357756 203084 357820 203088
rect 373396 203084 373460 203148
rect 492812 203084 492876 203148
rect 336044 202948 336108 203012
rect 337884 203008 337948 203012
rect 337884 202952 337934 203008
rect 337934 202952 337948 203008
rect 337884 202948 337948 202952
rect 339172 203008 339236 203012
rect 339172 202952 339222 203008
rect 339222 202952 339236 203008
rect 339172 202948 339236 202952
rect 342300 203008 342364 203012
rect 342300 202952 342314 203008
rect 342314 202952 342364 203008
rect 342300 202948 342364 202952
rect 342484 203008 342548 203012
rect 342484 202952 342498 203008
rect 342498 202952 342548 203008
rect 342484 202948 342548 202952
rect 343588 203008 343652 203012
rect 343588 202952 343638 203008
rect 343638 202952 343652 203008
rect 343588 202948 343652 202952
rect 344876 203008 344940 203012
rect 344876 202952 344926 203008
rect 344926 202952 344940 203008
rect 344876 202948 344940 202952
rect 345980 203008 346044 203012
rect 345980 202952 345994 203008
rect 345994 202952 346044 203008
rect 345980 202948 346044 202952
rect 347084 203008 347148 203012
rect 347084 202952 347134 203008
rect 347134 202952 347148 203008
rect 347084 202948 347148 202952
rect 348372 203008 348436 203012
rect 348372 202952 348386 203008
rect 348386 202952 348436 203008
rect 348372 202948 348436 202952
rect 349660 202948 349724 203012
rect 350948 203008 351012 203012
rect 350948 202952 350998 203008
rect 350998 202952 351012 203008
rect 350948 202948 351012 202952
rect 351684 203008 351748 203012
rect 351684 202952 351734 203008
rect 351734 202952 351748 203008
rect 351684 202948 351748 202952
rect 353340 203008 353404 203012
rect 353340 202952 353354 203008
rect 353354 202952 353404 203008
rect 353340 202948 353404 202952
rect 354260 203008 354324 203012
rect 354260 202952 354310 203008
rect 354310 202952 354324 203008
rect 354260 202948 354324 202952
rect 355548 203008 355612 203012
rect 355548 202952 355598 203008
rect 355598 202952 355612 203008
rect 355548 202948 355612 202952
rect 356468 203008 356532 203012
rect 356468 202952 356482 203008
rect 356482 202952 356532 203008
rect 356468 202948 356532 202952
rect 357940 202948 358004 203012
rect 358676 203008 358740 203012
rect 358676 202952 358690 203008
rect 358690 202952 358740 203008
rect 358676 202948 358740 202952
rect 359964 203008 360028 203012
rect 359964 202952 360014 203008
rect 360014 202952 360028 203008
rect 359964 202948 360028 202952
rect 361252 203008 361316 203012
rect 361252 202952 361302 203008
rect 361302 202952 361316 203008
rect 361252 202948 361316 202952
rect 362540 203008 362604 203012
rect 362540 202952 362554 203008
rect 362554 202952 362604 203008
rect 362540 202948 362604 202952
rect 363460 203008 363524 203012
rect 363460 202952 363510 203008
rect 363510 202952 363524 203008
rect 363460 202948 363524 202952
rect 364748 203008 364812 203012
rect 364748 202952 364762 203008
rect 364762 202952 364812 203008
rect 364748 202948 364812 202952
rect 451780 202948 451844 203012
rect 454172 202948 454236 203012
rect 456380 202948 456444 203012
rect 457852 202948 457916 203012
rect 458956 203008 459020 203012
rect 458956 202952 459006 203008
rect 459006 202952 459020 203008
rect 458956 202948 459020 202952
rect 460428 202948 460492 203012
rect 461532 202948 461596 203012
rect 462452 203008 462516 203012
rect 462452 202952 462466 203008
rect 462466 202952 462516 203008
rect 462452 202948 462516 202952
rect 463556 203008 463620 203012
rect 463556 202952 463606 203008
rect 463606 202952 463620 203008
rect 463556 202948 463620 202952
rect 464476 202948 464540 203012
rect 465764 202948 465828 203012
rect 467236 203008 467300 203012
rect 467236 202952 467286 203008
rect 467286 202952 467300 203008
rect 467236 202948 467300 202952
rect 468524 203008 468588 203012
rect 468524 202952 468538 203008
rect 468538 202952 468588 203008
rect 468524 202948 468588 202952
rect 469444 203008 469508 203012
rect 469444 202952 469458 203008
rect 469458 202952 469508 203008
rect 469444 202948 469508 202952
rect 470732 203008 470796 203012
rect 470732 202952 470746 203008
rect 470746 202952 470796 203008
rect 470732 202948 470796 202952
rect 471836 203008 471900 203012
rect 471836 202952 471850 203008
rect 471850 202952 471900 203008
rect 471836 202948 471900 202952
rect 472940 203008 473004 203012
rect 472940 202952 472954 203008
rect 472954 202952 473004 203008
rect 472940 202948 473004 202952
rect 474228 203008 474292 203012
rect 474228 202952 474242 203008
rect 474242 202952 474292 203008
rect 474228 202948 474292 202952
rect 475516 203008 475580 203012
rect 475516 202952 475566 203008
rect 475566 202952 475580 203008
rect 475516 202948 475580 202952
rect 476436 202948 476500 203012
rect 479932 202948 479996 203012
rect 481220 202948 481284 203012
rect 482140 202948 482204 203012
rect 483428 202948 483492 203012
rect 484716 202948 484780 203012
rect 539916 203008 539980 203012
rect 539916 202952 539966 203008
rect 539966 202952 539980 203008
rect 539916 202948 539980 202952
rect 342300 201724 342364 201788
rect 342276 201452 342340 201516
rect 448384 201512 448448 201516
rect 448384 201456 448426 201512
rect 448426 201456 448448 201512
rect 448384 201452 448448 201456
rect 538260 201044 538324 201108
rect 540284 200908 540348 200972
rect 543044 200772 543108 200836
rect 543228 200636 543292 200700
rect 539916 196012 539980 196076
rect 540100 195740 540164 195804
rect 540100 193156 540164 193220
rect 539916 183696 539980 183700
rect 539916 183640 539966 183696
rect 539966 183640 539980 183696
rect 539916 183636 539980 183640
rect 539916 176700 539980 176764
rect 540100 176428 540164 176492
rect 543044 173904 543108 173908
rect 543044 173848 543058 173904
rect 543058 173848 543108 173904
rect 543044 173844 543108 173848
rect 540100 167104 540164 167108
rect 540100 167048 540150 167104
rect 540150 167048 540164 167104
rect 540100 167044 540164 167048
rect 540100 164248 540164 164252
rect 540100 164192 540150 164248
rect 540150 164192 540164 164248
rect 540100 164188 540164 164192
rect 543044 164248 543108 164252
rect 543044 164192 543058 164248
rect 543058 164192 543108 164248
rect 543044 164188 543108 164192
rect 539916 162692 539980 162756
rect 540100 153172 540164 153236
rect 540100 147732 540164 147796
rect 539732 144876 539796 144940
rect 539916 120728 539980 120732
rect 539916 120672 539966 120728
rect 539966 120672 539980 120728
rect 539916 120668 539980 120672
rect 540100 115908 540164 115972
rect 303660 109032 303724 109036
rect 303660 108976 303674 109032
rect 303674 108976 303724 109032
rect 303660 108972 303724 108976
rect 308076 108972 308140 109036
rect 424180 109032 424244 109036
rect 424180 108976 424230 109032
rect 424230 108976 424244 109032
rect 424180 108972 424244 108976
rect 428044 108972 428108 109036
rect 67588 93876 67652 93940
rect 86908 93876 86972 93940
rect 106228 93876 106292 93940
rect 125548 93876 125612 93940
rect 9628 93740 9692 93804
rect 28948 93604 29012 93668
rect 48268 93604 48332 93668
rect 9628 93332 9692 93396
rect 28948 93196 29012 93260
rect 57836 93468 57900 93532
rect 67588 93604 67652 93668
rect 86908 93604 86972 93668
rect 106228 93604 106292 93668
rect 125548 93604 125612 93668
rect 48268 93196 48332 93260
rect 57836 93196 57900 93260
rect 540100 93468 540164 93532
rect 542860 80004 542924 80068
rect 541572 64772 541636 64836
rect 539548 50900 539612 50964
rect 542676 35804 542740 35868
rect 542492 21932 542556 21996
rect 542308 8196 542372 8260
<< metal4 >>
rect -8576 711418 -7976 711440
rect -8576 711182 -8394 711418
rect -8158 711182 -7976 711418
rect -8576 711098 -7976 711182
rect -8576 710862 -8394 711098
rect -8158 710862 -7976 711098
rect -8576 679254 -7976 710862
rect -8576 679018 -8394 679254
rect -8158 679018 -7976 679254
rect -8576 678934 -7976 679018
rect -8576 678698 -8394 678934
rect -8158 678698 -7976 678934
rect -8576 643254 -7976 678698
rect -8576 643018 -8394 643254
rect -8158 643018 -7976 643254
rect -8576 642934 -7976 643018
rect -8576 642698 -8394 642934
rect -8158 642698 -7976 642934
rect -8576 607254 -7976 642698
rect -8576 607018 -8394 607254
rect -8158 607018 -7976 607254
rect -8576 606934 -7976 607018
rect -8576 606698 -8394 606934
rect -8158 606698 -7976 606934
rect -8576 571254 -7976 606698
rect -8576 571018 -8394 571254
rect -8158 571018 -7976 571254
rect -8576 570934 -7976 571018
rect -8576 570698 -8394 570934
rect -8158 570698 -7976 570934
rect -8576 535254 -7976 570698
rect -8576 535018 -8394 535254
rect -8158 535018 -7976 535254
rect -8576 534934 -7976 535018
rect -8576 534698 -8394 534934
rect -8158 534698 -7976 534934
rect -8576 499254 -7976 534698
rect -8576 499018 -8394 499254
rect -8158 499018 -7976 499254
rect -8576 498934 -7976 499018
rect -8576 498698 -8394 498934
rect -8158 498698 -7976 498934
rect -8576 463254 -7976 498698
rect -8576 463018 -8394 463254
rect -8158 463018 -7976 463254
rect -8576 462934 -7976 463018
rect -8576 462698 -8394 462934
rect -8158 462698 -7976 462934
rect -8576 427254 -7976 462698
rect -8576 427018 -8394 427254
rect -8158 427018 -7976 427254
rect -8576 426934 -7976 427018
rect -8576 426698 -8394 426934
rect -8158 426698 -7976 426934
rect -8576 391254 -7976 426698
rect -8576 391018 -8394 391254
rect -8158 391018 -7976 391254
rect -8576 390934 -7976 391018
rect -8576 390698 -8394 390934
rect -8158 390698 -7976 390934
rect -8576 355254 -7976 390698
rect -8576 355018 -8394 355254
rect -8158 355018 -7976 355254
rect -8576 354934 -7976 355018
rect -8576 354698 -8394 354934
rect -8158 354698 -7976 354934
rect -8576 319254 -7976 354698
rect -8576 319018 -8394 319254
rect -8158 319018 -7976 319254
rect -8576 318934 -7976 319018
rect -8576 318698 -8394 318934
rect -8158 318698 -7976 318934
rect -8576 283254 -7976 318698
rect -8576 283018 -8394 283254
rect -8158 283018 -7976 283254
rect -8576 282934 -7976 283018
rect -8576 282698 -8394 282934
rect -8158 282698 -7976 282934
rect -8576 247254 -7976 282698
rect -8576 247018 -8394 247254
rect -8158 247018 -7976 247254
rect -8576 246934 -7976 247018
rect -8576 246698 -8394 246934
rect -8158 246698 -7976 246934
rect -8576 211254 -7976 246698
rect -8576 211018 -8394 211254
rect -8158 211018 -7976 211254
rect -8576 210934 -7976 211018
rect -8576 210698 -8394 210934
rect -8158 210698 -7976 210934
rect -8576 175254 -7976 210698
rect -8576 175018 -8394 175254
rect -8158 175018 -7976 175254
rect -8576 174934 -7976 175018
rect -8576 174698 -8394 174934
rect -8158 174698 -7976 174934
rect -8576 139254 -7976 174698
rect -8576 139018 -8394 139254
rect -8158 139018 -7976 139254
rect -8576 138934 -7976 139018
rect -8576 138698 -8394 138934
rect -8158 138698 -7976 138934
rect -8576 103254 -7976 138698
rect -8576 103018 -8394 103254
rect -8158 103018 -7976 103254
rect -8576 102934 -7976 103018
rect -8576 102698 -8394 102934
rect -8158 102698 -7976 102934
rect -8576 67254 -7976 102698
rect -8576 67018 -8394 67254
rect -8158 67018 -7976 67254
rect -8576 66934 -7976 67018
rect -8576 66698 -8394 66934
rect -8158 66698 -7976 66934
rect -8576 31254 -7976 66698
rect -8576 31018 -8394 31254
rect -8158 31018 -7976 31254
rect -8576 30934 -7976 31018
rect -8576 30698 -8394 30934
rect -8158 30698 -7976 30934
rect -8576 -6926 -7976 30698
rect -7636 710478 -7036 710500
rect -7636 710242 -7454 710478
rect -7218 710242 -7036 710478
rect -7636 710158 -7036 710242
rect -7636 709922 -7454 710158
rect -7218 709922 -7036 710158
rect -7636 697254 -7036 709922
rect 11604 710478 12204 711440
rect 11604 710242 11786 710478
rect 12022 710242 12204 710478
rect 11604 710158 12204 710242
rect 11604 709922 11786 710158
rect 12022 709922 12204 710158
rect -7636 697018 -7454 697254
rect -7218 697018 -7036 697254
rect -7636 696934 -7036 697018
rect -7636 696698 -7454 696934
rect -7218 696698 -7036 696934
rect -7636 661254 -7036 696698
rect -7636 661018 -7454 661254
rect -7218 661018 -7036 661254
rect -7636 660934 -7036 661018
rect -7636 660698 -7454 660934
rect -7218 660698 -7036 660934
rect -7636 625254 -7036 660698
rect -7636 625018 -7454 625254
rect -7218 625018 -7036 625254
rect -7636 624934 -7036 625018
rect -7636 624698 -7454 624934
rect -7218 624698 -7036 624934
rect -7636 589254 -7036 624698
rect -7636 589018 -7454 589254
rect -7218 589018 -7036 589254
rect -7636 588934 -7036 589018
rect -7636 588698 -7454 588934
rect -7218 588698 -7036 588934
rect -7636 553254 -7036 588698
rect -7636 553018 -7454 553254
rect -7218 553018 -7036 553254
rect -7636 552934 -7036 553018
rect -7636 552698 -7454 552934
rect -7218 552698 -7036 552934
rect -7636 517254 -7036 552698
rect -7636 517018 -7454 517254
rect -7218 517018 -7036 517254
rect -7636 516934 -7036 517018
rect -7636 516698 -7454 516934
rect -7218 516698 -7036 516934
rect -7636 481254 -7036 516698
rect -7636 481018 -7454 481254
rect -7218 481018 -7036 481254
rect -7636 480934 -7036 481018
rect -7636 480698 -7454 480934
rect -7218 480698 -7036 480934
rect -7636 445254 -7036 480698
rect -7636 445018 -7454 445254
rect -7218 445018 -7036 445254
rect -7636 444934 -7036 445018
rect -7636 444698 -7454 444934
rect -7218 444698 -7036 444934
rect -7636 409254 -7036 444698
rect -7636 409018 -7454 409254
rect -7218 409018 -7036 409254
rect -7636 408934 -7036 409018
rect -7636 408698 -7454 408934
rect -7218 408698 -7036 408934
rect -7636 373254 -7036 408698
rect -7636 373018 -7454 373254
rect -7218 373018 -7036 373254
rect -7636 372934 -7036 373018
rect -7636 372698 -7454 372934
rect -7218 372698 -7036 372934
rect -7636 337254 -7036 372698
rect -7636 337018 -7454 337254
rect -7218 337018 -7036 337254
rect -7636 336934 -7036 337018
rect -7636 336698 -7454 336934
rect -7218 336698 -7036 336934
rect -7636 301254 -7036 336698
rect -7636 301018 -7454 301254
rect -7218 301018 -7036 301254
rect -7636 300934 -7036 301018
rect -7636 300698 -7454 300934
rect -7218 300698 -7036 300934
rect -7636 265254 -7036 300698
rect -7636 265018 -7454 265254
rect -7218 265018 -7036 265254
rect -7636 264934 -7036 265018
rect -7636 264698 -7454 264934
rect -7218 264698 -7036 264934
rect -7636 229254 -7036 264698
rect -7636 229018 -7454 229254
rect -7218 229018 -7036 229254
rect -7636 228934 -7036 229018
rect -7636 228698 -7454 228934
rect -7218 228698 -7036 228934
rect -7636 193254 -7036 228698
rect -7636 193018 -7454 193254
rect -7218 193018 -7036 193254
rect -7636 192934 -7036 193018
rect -7636 192698 -7454 192934
rect -7218 192698 -7036 192934
rect -7636 157254 -7036 192698
rect -7636 157018 -7454 157254
rect -7218 157018 -7036 157254
rect -7636 156934 -7036 157018
rect -7636 156698 -7454 156934
rect -7218 156698 -7036 156934
rect -7636 121254 -7036 156698
rect -7636 121018 -7454 121254
rect -7218 121018 -7036 121254
rect -7636 120934 -7036 121018
rect -7636 120698 -7454 120934
rect -7218 120698 -7036 120934
rect -7636 85254 -7036 120698
rect -7636 85018 -7454 85254
rect -7218 85018 -7036 85254
rect -7636 84934 -7036 85018
rect -7636 84698 -7454 84934
rect -7218 84698 -7036 84934
rect -7636 49254 -7036 84698
rect -7636 49018 -7454 49254
rect -7218 49018 -7036 49254
rect -7636 48934 -7036 49018
rect -7636 48698 -7454 48934
rect -7218 48698 -7036 48934
rect -7636 13254 -7036 48698
rect -7636 13018 -7454 13254
rect -7218 13018 -7036 13254
rect -7636 12934 -7036 13018
rect -7636 12698 -7454 12934
rect -7218 12698 -7036 12934
rect -7636 -5986 -7036 12698
rect -6696 709538 -6096 709560
rect -6696 709302 -6514 709538
rect -6278 709302 -6096 709538
rect -6696 709218 -6096 709302
rect -6696 708982 -6514 709218
rect -6278 708982 -6096 709218
rect -6696 675654 -6096 708982
rect -6696 675418 -6514 675654
rect -6278 675418 -6096 675654
rect -6696 675334 -6096 675418
rect -6696 675098 -6514 675334
rect -6278 675098 -6096 675334
rect -6696 639654 -6096 675098
rect -6696 639418 -6514 639654
rect -6278 639418 -6096 639654
rect -6696 639334 -6096 639418
rect -6696 639098 -6514 639334
rect -6278 639098 -6096 639334
rect -6696 603654 -6096 639098
rect -6696 603418 -6514 603654
rect -6278 603418 -6096 603654
rect -6696 603334 -6096 603418
rect -6696 603098 -6514 603334
rect -6278 603098 -6096 603334
rect -6696 567654 -6096 603098
rect -6696 567418 -6514 567654
rect -6278 567418 -6096 567654
rect -6696 567334 -6096 567418
rect -6696 567098 -6514 567334
rect -6278 567098 -6096 567334
rect -6696 531654 -6096 567098
rect -6696 531418 -6514 531654
rect -6278 531418 -6096 531654
rect -6696 531334 -6096 531418
rect -6696 531098 -6514 531334
rect -6278 531098 -6096 531334
rect -6696 495654 -6096 531098
rect -6696 495418 -6514 495654
rect -6278 495418 -6096 495654
rect -6696 495334 -6096 495418
rect -6696 495098 -6514 495334
rect -6278 495098 -6096 495334
rect -6696 459654 -6096 495098
rect -6696 459418 -6514 459654
rect -6278 459418 -6096 459654
rect -6696 459334 -6096 459418
rect -6696 459098 -6514 459334
rect -6278 459098 -6096 459334
rect -6696 423654 -6096 459098
rect -6696 423418 -6514 423654
rect -6278 423418 -6096 423654
rect -6696 423334 -6096 423418
rect -6696 423098 -6514 423334
rect -6278 423098 -6096 423334
rect -6696 387654 -6096 423098
rect -6696 387418 -6514 387654
rect -6278 387418 -6096 387654
rect -6696 387334 -6096 387418
rect -6696 387098 -6514 387334
rect -6278 387098 -6096 387334
rect -6696 351654 -6096 387098
rect -6696 351418 -6514 351654
rect -6278 351418 -6096 351654
rect -6696 351334 -6096 351418
rect -6696 351098 -6514 351334
rect -6278 351098 -6096 351334
rect -6696 315654 -6096 351098
rect -6696 315418 -6514 315654
rect -6278 315418 -6096 315654
rect -6696 315334 -6096 315418
rect -6696 315098 -6514 315334
rect -6278 315098 -6096 315334
rect -6696 279654 -6096 315098
rect -6696 279418 -6514 279654
rect -6278 279418 -6096 279654
rect -6696 279334 -6096 279418
rect -6696 279098 -6514 279334
rect -6278 279098 -6096 279334
rect -6696 243654 -6096 279098
rect -6696 243418 -6514 243654
rect -6278 243418 -6096 243654
rect -6696 243334 -6096 243418
rect -6696 243098 -6514 243334
rect -6278 243098 -6096 243334
rect -6696 207654 -6096 243098
rect -6696 207418 -6514 207654
rect -6278 207418 -6096 207654
rect -6696 207334 -6096 207418
rect -6696 207098 -6514 207334
rect -6278 207098 -6096 207334
rect -6696 171654 -6096 207098
rect -6696 171418 -6514 171654
rect -6278 171418 -6096 171654
rect -6696 171334 -6096 171418
rect -6696 171098 -6514 171334
rect -6278 171098 -6096 171334
rect -6696 135654 -6096 171098
rect -6696 135418 -6514 135654
rect -6278 135418 -6096 135654
rect -6696 135334 -6096 135418
rect -6696 135098 -6514 135334
rect -6278 135098 -6096 135334
rect -6696 99654 -6096 135098
rect -6696 99418 -6514 99654
rect -6278 99418 -6096 99654
rect -6696 99334 -6096 99418
rect -6696 99098 -6514 99334
rect -6278 99098 -6096 99334
rect -6696 63654 -6096 99098
rect -6696 63418 -6514 63654
rect -6278 63418 -6096 63654
rect -6696 63334 -6096 63418
rect -6696 63098 -6514 63334
rect -6278 63098 -6096 63334
rect -6696 27654 -6096 63098
rect -6696 27418 -6514 27654
rect -6278 27418 -6096 27654
rect -6696 27334 -6096 27418
rect -6696 27098 -6514 27334
rect -6278 27098 -6096 27334
rect -6696 -5046 -6096 27098
rect -5756 708598 -5156 708620
rect -5756 708362 -5574 708598
rect -5338 708362 -5156 708598
rect -5756 708278 -5156 708362
rect -5756 708042 -5574 708278
rect -5338 708042 -5156 708278
rect -5756 693654 -5156 708042
rect 8004 708598 8604 709560
rect 8004 708362 8186 708598
rect 8422 708362 8604 708598
rect 8004 708278 8604 708362
rect 8004 708042 8186 708278
rect 8422 708042 8604 708278
rect -5756 693418 -5574 693654
rect -5338 693418 -5156 693654
rect -5756 693334 -5156 693418
rect -5756 693098 -5574 693334
rect -5338 693098 -5156 693334
rect -5756 657654 -5156 693098
rect -5756 657418 -5574 657654
rect -5338 657418 -5156 657654
rect -5756 657334 -5156 657418
rect -5756 657098 -5574 657334
rect -5338 657098 -5156 657334
rect -5756 621654 -5156 657098
rect -5756 621418 -5574 621654
rect -5338 621418 -5156 621654
rect -5756 621334 -5156 621418
rect -5756 621098 -5574 621334
rect -5338 621098 -5156 621334
rect -5756 585654 -5156 621098
rect -5756 585418 -5574 585654
rect -5338 585418 -5156 585654
rect -5756 585334 -5156 585418
rect -5756 585098 -5574 585334
rect -5338 585098 -5156 585334
rect -5756 549654 -5156 585098
rect -5756 549418 -5574 549654
rect -5338 549418 -5156 549654
rect -5756 549334 -5156 549418
rect -5756 549098 -5574 549334
rect -5338 549098 -5156 549334
rect -5756 513654 -5156 549098
rect -5756 513418 -5574 513654
rect -5338 513418 -5156 513654
rect -5756 513334 -5156 513418
rect -5756 513098 -5574 513334
rect -5338 513098 -5156 513334
rect -5756 477654 -5156 513098
rect -5756 477418 -5574 477654
rect -5338 477418 -5156 477654
rect -5756 477334 -5156 477418
rect -5756 477098 -5574 477334
rect -5338 477098 -5156 477334
rect -5756 441654 -5156 477098
rect -5756 441418 -5574 441654
rect -5338 441418 -5156 441654
rect -5756 441334 -5156 441418
rect -5756 441098 -5574 441334
rect -5338 441098 -5156 441334
rect -5756 405654 -5156 441098
rect -5756 405418 -5574 405654
rect -5338 405418 -5156 405654
rect -5756 405334 -5156 405418
rect -5756 405098 -5574 405334
rect -5338 405098 -5156 405334
rect -5756 369654 -5156 405098
rect -5756 369418 -5574 369654
rect -5338 369418 -5156 369654
rect -5756 369334 -5156 369418
rect -5756 369098 -5574 369334
rect -5338 369098 -5156 369334
rect -5756 333654 -5156 369098
rect -5756 333418 -5574 333654
rect -5338 333418 -5156 333654
rect -5756 333334 -5156 333418
rect -5756 333098 -5574 333334
rect -5338 333098 -5156 333334
rect -5756 297654 -5156 333098
rect -5756 297418 -5574 297654
rect -5338 297418 -5156 297654
rect -5756 297334 -5156 297418
rect -5756 297098 -5574 297334
rect -5338 297098 -5156 297334
rect -5756 261654 -5156 297098
rect -5756 261418 -5574 261654
rect -5338 261418 -5156 261654
rect -5756 261334 -5156 261418
rect -5756 261098 -5574 261334
rect -5338 261098 -5156 261334
rect -5756 225654 -5156 261098
rect -5756 225418 -5574 225654
rect -5338 225418 -5156 225654
rect -5756 225334 -5156 225418
rect -5756 225098 -5574 225334
rect -5338 225098 -5156 225334
rect -5756 189654 -5156 225098
rect -5756 189418 -5574 189654
rect -5338 189418 -5156 189654
rect -5756 189334 -5156 189418
rect -5756 189098 -5574 189334
rect -5338 189098 -5156 189334
rect -5756 153654 -5156 189098
rect -5756 153418 -5574 153654
rect -5338 153418 -5156 153654
rect -5756 153334 -5156 153418
rect -5756 153098 -5574 153334
rect -5338 153098 -5156 153334
rect -5756 117654 -5156 153098
rect -5756 117418 -5574 117654
rect -5338 117418 -5156 117654
rect -5756 117334 -5156 117418
rect -5756 117098 -5574 117334
rect -5338 117098 -5156 117334
rect -5756 81654 -5156 117098
rect -5756 81418 -5574 81654
rect -5338 81418 -5156 81654
rect -5756 81334 -5156 81418
rect -5756 81098 -5574 81334
rect -5338 81098 -5156 81334
rect -5756 45654 -5156 81098
rect -5756 45418 -5574 45654
rect -5338 45418 -5156 45654
rect -5756 45334 -5156 45418
rect -5756 45098 -5574 45334
rect -5338 45098 -5156 45334
rect -5756 9654 -5156 45098
rect -5756 9418 -5574 9654
rect -5338 9418 -5156 9654
rect -5756 9334 -5156 9418
rect -5756 9098 -5574 9334
rect -5338 9098 -5156 9334
rect -5756 -4106 -5156 9098
rect -4816 707658 -4216 707680
rect -4816 707422 -4634 707658
rect -4398 707422 -4216 707658
rect -4816 707338 -4216 707422
rect -4816 707102 -4634 707338
rect -4398 707102 -4216 707338
rect -4816 672054 -4216 707102
rect -4816 671818 -4634 672054
rect -4398 671818 -4216 672054
rect -4816 671734 -4216 671818
rect -4816 671498 -4634 671734
rect -4398 671498 -4216 671734
rect -4816 636054 -4216 671498
rect -4816 635818 -4634 636054
rect -4398 635818 -4216 636054
rect -4816 635734 -4216 635818
rect -4816 635498 -4634 635734
rect -4398 635498 -4216 635734
rect -4816 600054 -4216 635498
rect -4816 599818 -4634 600054
rect -4398 599818 -4216 600054
rect -4816 599734 -4216 599818
rect -4816 599498 -4634 599734
rect -4398 599498 -4216 599734
rect -4816 564054 -4216 599498
rect -4816 563818 -4634 564054
rect -4398 563818 -4216 564054
rect -4816 563734 -4216 563818
rect -4816 563498 -4634 563734
rect -4398 563498 -4216 563734
rect -4816 528054 -4216 563498
rect -4816 527818 -4634 528054
rect -4398 527818 -4216 528054
rect -4816 527734 -4216 527818
rect -4816 527498 -4634 527734
rect -4398 527498 -4216 527734
rect -4816 492054 -4216 527498
rect -4816 491818 -4634 492054
rect -4398 491818 -4216 492054
rect -4816 491734 -4216 491818
rect -4816 491498 -4634 491734
rect -4398 491498 -4216 491734
rect -4816 456054 -4216 491498
rect -4816 455818 -4634 456054
rect -4398 455818 -4216 456054
rect -4816 455734 -4216 455818
rect -4816 455498 -4634 455734
rect -4398 455498 -4216 455734
rect -4816 420054 -4216 455498
rect -4816 419818 -4634 420054
rect -4398 419818 -4216 420054
rect -4816 419734 -4216 419818
rect -4816 419498 -4634 419734
rect -4398 419498 -4216 419734
rect -4816 384054 -4216 419498
rect -4816 383818 -4634 384054
rect -4398 383818 -4216 384054
rect -4816 383734 -4216 383818
rect -4816 383498 -4634 383734
rect -4398 383498 -4216 383734
rect -4816 348054 -4216 383498
rect -4816 347818 -4634 348054
rect -4398 347818 -4216 348054
rect -4816 347734 -4216 347818
rect -4816 347498 -4634 347734
rect -4398 347498 -4216 347734
rect -4816 312054 -4216 347498
rect -4816 311818 -4634 312054
rect -4398 311818 -4216 312054
rect -4816 311734 -4216 311818
rect -4816 311498 -4634 311734
rect -4398 311498 -4216 311734
rect -4816 276054 -4216 311498
rect -4816 275818 -4634 276054
rect -4398 275818 -4216 276054
rect -4816 275734 -4216 275818
rect -4816 275498 -4634 275734
rect -4398 275498 -4216 275734
rect -4816 240054 -4216 275498
rect -4816 239818 -4634 240054
rect -4398 239818 -4216 240054
rect -4816 239734 -4216 239818
rect -4816 239498 -4634 239734
rect -4398 239498 -4216 239734
rect -4816 204054 -4216 239498
rect -4816 203818 -4634 204054
rect -4398 203818 -4216 204054
rect -4816 203734 -4216 203818
rect -4816 203498 -4634 203734
rect -4398 203498 -4216 203734
rect -4816 168054 -4216 203498
rect -4816 167818 -4634 168054
rect -4398 167818 -4216 168054
rect -4816 167734 -4216 167818
rect -4816 167498 -4634 167734
rect -4398 167498 -4216 167734
rect -4816 132054 -4216 167498
rect -4816 131818 -4634 132054
rect -4398 131818 -4216 132054
rect -4816 131734 -4216 131818
rect -4816 131498 -4634 131734
rect -4398 131498 -4216 131734
rect -4816 96054 -4216 131498
rect -4816 95818 -4634 96054
rect -4398 95818 -4216 96054
rect -4816 95734 -4216 95818
rect -4816 95498 -4634 95734
rect -4398 95498 -4216 95734
rect -4816 60054 -4216 95498
rect -4816 59818 -4634 60054
rect -4398 59818 -4216 60054
rect -4816 59734 -4216 59818
rect -4816 59498 -4634 59734
rect -4398 59498 -4216 59734
rect -4816 24054 -4216 59498
rect -4816 23818 -4634 24054
rect -4398 23818 -4216 24054
rect -4816 23734 -4216 23818
rect -4816 23498 -4634 23734
rect -4398 23498 -4216 23734
rect -4816 -3166 -4216 23498
rect -3876 706718 -3276 706740
rect -3876 706482 -3694 706718
rect -3458 706482 -3276 706718
rect -3876 706398 -3276 706482
rect -3876 706162 -3694 706398
rect -3458 706162 -3276 706398
rect -3876 690054 -3276 706162
rect 4404 706718 5004 707680
rect 4404 706482 4586 706718
rect 4822 706482 5004 706718
rect 4404 706398 5004 706482
rect 4404 706162 4586 706398
rect 4822 706162 5004 706398
rect -3876 689818 -3694 690054
rect -3458 689818 -3276 690054
rect -3876 689734 -3276 689818
rect -3876 689498 -3694 689734
rect -3458 689498 -3276 689734
rect -3876 654054 -3276 689498
rect -3876 653818 -3694 654054
rect -3458 653818 -3276 654054
rect -3876 653734 -3276 653818
rect -3876 653498 -3694 653734
rect -3458 653498 -3276 653734
rect -3876 618054 -3276 653498
rect -3876 617818 -3694 618054
rect -3458 617818 -3276 618054
rect -3876 617734 -3276 617818
rect -3876 617498 -3694 617734
rect -3458 617498 -3276 617734
rect -3876 582054 -3276 617498
rect -3876 581818 -3694 582054
rect -3458 581818 -3276 582054
rect -3876 581734 -3276 581818
rect -3876 581498 -3694 581734
rect -3458 581498 -3276 581734
rect -3876 546054 -3276 581498
rect -3876 545818 -3694 546054
rect -3458 545818 -3276 546054
rect -3876 545734 -3276 545818
rect -3876 545498 -3694 545734
rect -3458 545498 -3276 545734
rect -3876 510054 -3276 545498
rect -3876 509818 -3694 510054
rect -3458 509818 -3276 510054
rect -3876 509734 -3276 509818
rect -3876 509498 -3694 509734
rect -3458 509498 -3276 509734
rect -3876 474054 -3276 509498
rect -3876 473818 -3694 474054
rect -3458 473818 -3276 474054
rect -3876 473734 -3276 473818
rect -3876 473498 -3694 473734
rect -3458 473498 -3276 473734
rect -3876 438054 -3276 473498
rect -3876 437818 -3694 438054
rect -3458 437818 -3276 438054
rect -3876 437734 -3276 437818
rect -3876 437498 -3694 437734
rect -3458 437498 -3276 437734
rect -3876 402054 -3276 437498
rect -3876 401818 -3694 402054
rect -3458 401818 -3276 402054
rect -3876 401734 -3276 401818
rect -3876 401498 -3694 401734
rect -3458 401498 -3276 401734
rect -3876 366054 -3276 401498
rect -3876 365818 -3694 366054
rect -3458 365818 -3276 366054
rect -3876 365734 -3276 365818
rect -3876 365498 -3694 365734
rect -3458 365498 -3276 365734
rect -3876 330054 -3276 365498
rect -3876 329818 -3694 330054
rect -3458 329818 -3276 330054
rect -3876 329734 -3276 329818
rect -3876 329498 -3694 329734
rect -3458 329498 -3276 329734
rect -3876 294054 -3276 329498
rect -3876 293818 -3694 294054
rect -3458 293818 -3276 294054
rect -3876 293734 -3276 293818
rect -3876 293498 -3694 293734
rect -3458 293498 -3276 293734
rect -3876 258054 -3276 293498
rect -3876 257818 -3694 258054
rect -3458 257818 -3276 258054
rect -3876 257734 -3276 257818
rect -3876 257498 -3694 257734
rect -3458 257498 -3276 257734
rect -3876 222054 -3276 257498
rect -3876 221818 -3694 222054
rect -3458 221818 -3276 222054
rect -3876 221734 -3276 221818
rect -3876 221498 -3694 221734
rect -3458 221498 -3276 221734
rect -3876 186054 -3276 221498
rect -3876 185818 -3694 186054
rect -3458 185818 -3276 186054
rect -3876 185734 -3276 185818
rect -3876 185498 -3694 185734
rect -3458 185498 -3276 185734
rect -3876 150054 -3276 185498
rect -3876 149818 -3694 150054
rect -3458 149818 -3276 150054
rect -3876 149734 -3276 149818
rect -3876 149498 -3694 149734
rect -3458 149498 -3276 149734
rect -3876 114054 -3276 149498
rect -3876 113818 -3694 114054
rect -3458 113818 -3276 114054
rect -3876 113734 -3276 113818
rect -3876 113498 -3694 113734
rect -3458 113498 -3276 113734
rect -3876 78054 -3276 113498
rect -3876 77818 -3694 78054
rect -3458 77818 -3276 78054
rect -3876 77734 -3276 77818
rect -3876 77498 -3694 77734
rect -3458 77498 -3276 77734
rect -3876 42054 -3276 77498
rect -3876 41818 -3694 42054
rect -3458 41818 -3276 42054
rect -3876 41734 -3276 41818
rect -3876 41498 -3694 41734
rect -3458 41498 -3276 41734
rect -3876 6054 -3276 41498
rect -3876 5818 -3694 6054
rect -3458 5818 -3276 6054
rect -3876 5734 -3276 5818
rect -3876 5498 -3694 5734
rect -3458 5498 -3276 5734
rect -3876 -2226 -3276 5498
rect -2936 705778 -2336 705800
rect -2936 705542 -2754 705778
rect -2518 705542 -2336 705778
rect -2936 705458 -2336 705542
rect -2936 705222 -2754 705458
rect -2518 705222 -2336 705458
rect -2936 668454 -2336 705222
rect -2936 668218 -2754 668454
rect -2518 668218 -2336 668454
rect -2936 668134 -2336 668218
rect -2936 667898 -2754 668134
rect -2518 667898 -2336 668134
rect -2936 632454 -2336 667898
rect -2936 632218 -2754 632454
rect -2518 632218 -2336 632454
rect -2936 632134 -2336 632218
rect -2936 631898 -2754 632134
rect -2518 631898 -2336 632134
rect -2936 596454 -2336 631898
rect -2936 596218 -2754 596454
rect -2518 596218 -2336 596454
rect -2936 596134 -2336 596218
rect -2936 595898 -2754 596134
rect -2518 595898 -2336 596134
rect -2936 560454 -2336 595898
rect -2936 560218 -2754 560454
rect -2518 560218 -2336 560454
rect -2936 560134 -2336 560218
rect -2936 559898 -2754 560134
rect -2518 559898 -2336 560134
rect -2936 524454 -2336 559898
rect -2936 524218 -2754 524454
rect -2518 524218 -2336 524454
rect -2936 524134 -2336 524218
rect -2936 523898 -2754 524134
rect -2518 523898 -2336 524134
rect -2936 488454 -2336 523898
rect -2936 488218 -2754 488454
rect -2518 488218 -2336 488454
rect -2936 488134 -2336 488218
rect -2936 487898 -2754 488134
rect -2518 487898 -2336 488134
rect -2936 452454 -2336 487898
rect -2936 452218 -2754 452454
rect -2518 452218 -2336 452454
rect -2936 452134 -2336 452218
rect -2936 451898 -2754 452134
rect -2518 451898 -2336 452134
rect -2936 416454 -2336 451898
rect -2936 416218 -2754 416454
rect -2518 416218 -2336 416454
rect -2936 416134 -2336 416218
rect -2936 415898 -2754 416134
rect -2518 415898 -2336 416134
rect -2936 380454 -2336 415898
rect -2936 380218 -2754 380454
rect -2518 380218 -2336 380454
rect -2936 380134 -2336 380218
rect -2936 379898 -2754 380134
rect -2518 379898 -2336 380134
rect -2936 344454 -2336 379898
rect -2936 344218 -2754 344454
rect -2518 344218 -2336 344454
rect -2936 344134 -2336 344218
rect -2936 343898 -2754 344134
rect -2518 343898 -2336 344134
rect -2936 308454 -2336 343898
rect -2936 308218 -2754 308454
rect -2518 308218 -2336 308454
rect -2936 308134 -2336 308218
rect -2936 307898 -2754 308134
rect -2518 307898 -2336 308134
rect -2936 272454 -2336 307898
rect -2936 272218 -2754 272454
rect -2518 272218 -2336 272454
rect -2936 272134 -2336 272218
rect -2936 271898 -2754 272134
rect -2518 271898 -2336 272134
rect -2936 236454 -2336 271898
rect -2936 236218 -2754 236454
rect -2518 236218 -2336 236454
rect -2936 236134 -2336 236218
rect -2936 235898 -2754 236134
rect -2518 235898 -2336 236134
rect -2936 200454 -2336 235898
rect -2936 200218 -2754 200454
rect -2518 200218 -2336 200454
rect -2936 200134 -2336 200218
rect -2936 199898 -2754 200134
rect -2518 199898 -2336 200134
rect -2936 164454 -2336 199898
rect -2936 164218 -2754 164454
rect -2518 164218 -2336 164454
rect -2936 164134 -2336 164218
rect -2936 163898 -2754 164134
rect -2518 163898 -2336 164134
rect -2936 128454 -2336 163898
rect -2936 128218 -2754 128454
rect -2518 128218 -2336 128454
rect -2936 128134 -2336 128218
rect -2936 127898 -2754 128134
rect -2518 127898 -2336 128134
rect -2936 92454 -2336 127898
rect -2936 92218 -2754 92454
rect -2518 92218 -2336 92454
rect -2936 92134 -2336 92218
rect -2936 91898 -2754 92134
rect -2518 91898 -2336 92134
rect -2936 56454 -2336 91898
rect -2936 56218 -2754 56454
rect -2518 56218 -2336 56454
rect -2936 56134 -2336 56218
rect -2936 55898 -2754 56134
rect -2518 55898 -2336 56134
rect -2936 20454 -2336 55898
rect -2936 20218 -2754 20454
rect -2518 20218 -2336 20454
rect -2936 20134 -2336 20218
rect -2936 19898 -2754 20134
rect -2518 19898 -2336 20134
rect -2936 -1286 -2336 19898
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 686454 -1396 704282
rect -1996 686218 -1814 686454
rect -1578 686218 -1396 686454
rect -1996 686134 -1396 686218
rect -1996 685898 -1814 686134
rect -1578 685898 -1396 686134
rect -1996 650454 -1396 685898
rect -1996 650218 -1814 650454
rect -1578 650218 -1396 650454
rect -1996 650134 -1396 650218
rect -1996 649898 -1814 650134
rect -1578 649898 -1396 650134
rect -1996 614454 -1396 649898
rect -1996 614218 -1814 614454
rect -1578 614218 -1396 614454
rect -1996 614134 -1396 614218
rect -1996 613898 -1814 614134
rect -1578 613898 -1396 614134
rect -1996 578454 -1396 613898
rect -1996 578218 -1814 578454
rect -1578 578218 -1396 578454
rect -1996 578134 -1396 578218
rect -1996 577898 -1814 578134
rect -1578 577898 -1396 578134
rect -1996 542454 -1396 577898
rect -1996 542218 -1814 542454
rect -1578 542218 -1396 542454
rect -1996 542134 -1396 542218
rect -1996 541898 -1814 542134
rect -1578 541898 -1396 542134
rect -1996 506454 -1396 541898
rect -1996 506218 -1814 506454
rect -1578 506218 -1396 506454
rect -1996 506134 -1396 506218
rect -1996 505898 -1814 506134
rect -1578 505898 -1396 506134
rect -1996 470454 -1396 505898
rect -1996 470218 -1814 470454
rect -1578 470218 -1396 470454
rect -1996 470134 -1396 470218
rect -1996 469898 -1814 470134
rect -1578 469898 -1396 470134
rect -1996 434454 -1396 469898
rect -1996 434218 -1814 434454
rect -1578 434218 -1396 434454
rect -1996 434134 -1396 434218
rect -1996 433898 -1814 434134
rect -1578 433898 -1396 434134
rect -1996 398454 -1396 433898
rect -1996 398218 -1814 398454
rect -1578 398218 -1396 398454
rect -1996 398134 -1396 398218
rect -1996 397898 -1814 398134
rect -1578 397898 -1396 398134
rect -1996 362454 -1396 397898
rect -1996 362218 -1814 362454
rect -1578 362218 -1396 362454
rect -1996 362134 -1396 362218
rect -1996 361898 -1814 362134
rect -1578 361898 -1396 362134
rect -1996 326454 -1396 361898
rect -1996 326218 -1814 326454
rect -1578 326218 -1396 326454
rect -1996 326134 -1396 326218
rect -1996 325898 -1814 326134
rect -1578 325898 -1396 326134
rect -1996 290454 -1396 325898
rect -1996 290218 -1814 290454
rect -1578 290218 -1396 290454
rect -1996 290134 -1396 290218
rect -1996 289898 -1814 290134
rect -1578 289898 -1396 290134
rect -1996 254454 -1396 289898
rect -1996 254218 -1814 254454
rect -1578 254218 -1396 254454
rect -1996 254134 -1396 254218
rect -1996 253898 -1814 254134
rect -1578 253898 -1396 254134
rect -1996 218454 -1396 253898
rect -1996 218218 -1814 218454
rect -1578 218218 -1396 218454
rect -1996 218134 -1396 218218
rect -1996 217898 -1814 218134
rect -1578 217898 -1396 218134
rect -1996 182454 -1396 217898
rect -1996 182218 -1814 182454
rect -1578 182218 -1396 182454
rect -1996 182134 -1396 182218
rect -1996 181898 -1814 182134
rect -1578 181898 -1396 182134
rect -1996 146454 -1396 181898
rect -1996 146218 -1814 146454
rect -1578 146218 -1396 146454
rect -1996 146134 -1396 146218
rect -1996 145898 -1814 146134
rect -1578 145898 -1396 146134
rect -1996 110454 -1396 145898
rect -1996 110218 -1814 110454
rect -1578 110218 -1396 110454
rect -1996 110134 -1396 110218
rect -1996 109898 -1814 110134
rect -1578 109898 -1396 110134
rect -1996 74454 -1396 109898
rect -1996 74218 -1814 74454
rect -1578 74218 -1396 74454
rect -1996 74134 -1396 74218
rect -1996 73898 -1814 74134
rect -1578 73898 -1396 74134
rect -1996 38454 -1396 73898
rect -1996 38218 -1814 38454
rect -1578 38218 -1396 38454
rect -1996 38134 -1396 38218
rect -1996 37898 -1814 38134
rect -1578 37898 -1396 38134
rect -1996 2454 -1396 37898
rect -1996 2218 -1814 2454
rect -1578 2218 -1396 2454
rect -1996 2134 -1396 2218
rect -1996 1898 -1814 2134
rect -1578 1898 -1396 2134
rect -1996 -346 -1396 1898
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 804 704838 1404 705800
rect 804 704602 986 704838
rect 1222 704602 1404 704838
rect 804 704518 1404 704602
rect 804 704282 986 704518
rect 1222 704282 1404 704518
rect 804 686454 1404 704282
rect 804 686218 986 686454
rect 1222 686218 1404 686454
rect 804 686134 1404 686218
rect 804 685898 986 686134
rect 1222 685898 1404 686134
rect 804 650454 1404 685898
rect 804 650218 986 650454
rect 1222 650218 1404 650454
rect 804 650134 1404 650218
rect 804 649898 986 650134
rect 1222 649898 1404 650134
rect 804 614454 1404 649898
rect 804 614218 986 614454
rect 1222 614218 1404 614454
rect 804 614134 1404 614218
rect 804 613898 986 614134
rect 1222 613898 1404 614134
rect 804 578454 1404 613898
rect 804 578218 986 578454
rect 1222 578218 1404 578454
rect 804 578134 1404 578218
rect 804 577898 986 578134
rect 1222 577898 1404 578134
rect 804 542454 1404 577898
rect 804 542218 986 542454
rect 1222 542218 1404 542454
rect 804 542134 1404 542218
rect 804 541898 986 542134
rect 1222 541898 1404 542134
rect 804 506454 1404 541898
rect 804 506218 986 506454
rect 1222 506218 1404 506454
rect 804 506134 1404 506218
rect 804 505898 986 506134
rect 1222 505898 1404 506134
rect 804 470454 1404 505898
rect 804 470218 986 470454
rect 1222 470218 1404 470454
rect 804 470134 1404 470218
rect 804 469898 986 470134
rect 1222 469898 1404 470134
rect 804 434454 1404 469898
rect 804 434218 986 434454
rect 1222 434218 1404 434454
rect 804 434134 1404 434218
rect 804 433898 986 434134
rect 1222 433898 1404 434134
rect 804 398454 1404 433898
rect 804 398218 986 398454
rect 1222 398218 1404 398454
rect 804 398134 1404 398218
rect 804 397898 986 398134
rect 1222 397898 1404 398134
rect 804 362454 1404 397898
rect 804 362218 986 362454
rect 1222 362218 1404 362454
rect 804 362134 1404 362218
rect 804 361898 986 362134
rect 1222 361898 1404 362134
rect 804 326454 1404 361898
rect 804 326218 986 326454
rect 1222 326218 1404 326454
rect 804 326134 1404 326218
rect 804 325898 986 326134
rect 1222 325898 1404 326134
rect 804 290454 1404 325898
rect 804 290218 986 290454
rect 1222 290218 1404 290454
rect 804 290134 1404 290218
rect 804 289898 986 290134
rect 1222 289898 1404 290134
rect 804 254454 1404 289898
rect 804 254218 986 254454
rect 1222 254218 1404 254454
rect 804 254134 1404 254218
rect 804 253898 986 254134
rect 1222 253898 1404 254134
rect 804 218454 1404 253898
rect 804 218218 986 218454
rect 1222 218218 1404 218454
rect 804 218134 1404 218218
rect 804 217898 986 218134
rect 1222 217898 1404 218134
rect 804 182454 1404 217898
rect 804 182218 986 182454
rect 1222 182218 1404 182454
rect 804 182134 1404 182218
rect 804 181898 986 182134
rect 1222 181898 1404 182134
rect 804 146454 1404 181898
rect 804 146218 986 146454
rect 1222 146218 1404 146454
rect 804 146134 1404 146218
rect 804 145898 986 146134
rect 1222 145898 1404 146134
rect 804 110454 1404 145898
rect 804 110218 986 110454
rect 1222 110218 1404 110454
rect 804 110134 1404 110218
rect 804 109898 986 110134
rect 1222 109898 1404 110134
rect 804 74454 1404 109898
rect 804 74218 986 74454
rect 1222 74218 1404 74454
rect 804 74134 1404 74218
rect 804 73898 986 74134
rect 1222 73898 1404 74134
rect 804 38454 1404 73898
rect 804 38218 986 38454
rect 1222 38218 1404 38454
rect 804 38134 1404 38218
rect 804 37898 986 38134
rect 1222 37898 1404 38134
rect 804 2454 1404 37898
rect 804 2218 986 2454
rect 1222 2218 1404 2454
rect 804 2134 1404 2218
rect 804 1898 986 2134
rect 1222 1898 1404 2134
rect 804 -346 1404 1898
rect 804 -582 986 -346
rect 1222 -582 1404 -346
rect 804 -666 1404 -582
rect 804 -902 986 -666
rect 1222 -902 1404 -666
rect -2936 -1522 -2754 -1286
rect -2518 -1522 -2336 -1286
rect -2936 -1606 -2336 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 -2336 -1606
rect -2936 -1864 -2336 -1842
rect 804 -1864 1404 -902
rect 4404 690054 5004 706162
rect 4404 689818 4586 690054
rect 4822 689818 5004 690054
rect 4404 689734 5004 689818
rect 4404 689498 4586 689734
rect 4822 689498 5004 689734
rect 4404 654054 5004 689498
rect 4404 653818 4586 654054
rect 4822 653818 5004 654054
rect 4404 653734 5004 653818
rect 4404 653498 4586 653734
rect 4822 653498 5004 653734
rect 4404 618054 5004 653498
rect 4404 617818 4586 618054
rect 4822 617818 5004 618054
rect 4404 617734 5004 617818
rect 4404 617498 4586 617734
rect 4822 617498 5004 617734
rect 4404 582054 5004 617498
rect 4404 581818 4586 582054
rect 4822 581818 5004 582054
rect 4404 581734 5004 581818
rect 4404 581498 4586 581734
rect 4822 581498 5004 581734
rect 4404 546054 5004 581498
rect 4404 545818 4586 546054
rect 4822 545818 5004 546054
rect 4404 545734 5004 545818
rect 4404 545498 4586 545734
rect 4822 545498 5004 545734
rect 4404 510054 5004 545498
rect 4404 509818 4586 510054
rect 4822 509818 5004 510054
rect 4404 509734 5004 509818
rect 4404 509498 4586 509734
rect 4822 509498 5004 509734
rect 4404 474054 5004 509498
rect 4404 473818 4586 474054
rect 4822 473818 5004 474054
rect 4404 473734 5004 473818
rect 4404 473498 4586 473734
rect 4822 473498 5004 473734
rect 4404 438054 5004 473498
rect 4404 437818 4586 438054
rect 4822 437818 5004 438054
rect 4404 437734 5004 437818
rect 4404 437498 4586 437734
rect 4822 437498 5004 437734
rect 4404 402054 5004 437498
rect 4404 401818 4586 402054
rect 4822 401818 5004 402054
rect 4404 401734 5004 401818
rect 4404 401498 4586 401734
rect 4822 401498 5004 401734
rect 4404 366054 5004 401498
rect 4404 365818 4586 366054
rect 4822 365818 5004 366054
rect 4404 365734 5004 365818
rect 4404 365498 4586 365734
rect 4822 365498 5004 365734
rect 4404 330054 5004 365498
rect 4404 329818 4586 330054
rect 4822 329818 5004 330054
rect 4404 329734 5004 329818
rect 4404 329498 4586 329734
rect 4822 329498 5004 329734
rect 4404 294054 5004 329498
rect 4404 293818 4586 294054
rect 4822 293818 5004 294054
rect 4404 293734 5004 293818
rect 4404 293498 4586 293734
rect 4822 293498 5004 293734
rect 4404 258054 5004 293498
rect 4404 257818 4586 258054
rect 4822 257818 5004 258054
rect 4404 257734 5004 257818
rect 4404 257498 4586 257734
rect 4822 257498 5004 257734
rect 4404 222054 5004 257498
rect 4404 221818 4586 222054
rect 4822 221818 5004 222054
rect 4404 221734 5004 221818
rect 4404 221498 4586 221734
rect 4822 221498 5004 221734
rect 4404 186054 5004 221498
rect 4404 185818 4586 186054
rect 4822 185818 5004 186054
rect 4404 185734 5004 185818
rect 4404 185498 4586 185734
rect 4822 185498 5004 185734
rect 4404 150054 5004 185498
rect 4404 149818 4586 150054
rect 4822 149818 5004 150054
rect 4404 149734 5004 149818
rect 4404 149498 4586 149734
rect 4822 149498 5004 149734
rect 4404 114054 5004 149498
rect 4404 113818 4586 114054
rect 4822 113818 5004 114054
rect 4404 113734 5004 113818
rect 4404 113498 4586 113734
rect 4822 113498 5004 113734
rect 4404 78054 5004 113498
rect 4404 77818 4586 78054
rect 4822 77818 5004 78054
rect 4404 77734 5004 77818
rect 4404 77498 4586 77734
rect 4822 77498 5004 77734
rect 4404 42054 5004 77498
rect 4404 41818 4586 42054
rect 4822 41818 5004 42054
rect 4404 41734 5004 41818
rect 4404 41498 4586 41734
rect 4822 41498 5004 41734
rect 4404 6054 5004 41498
rect 4404 5818 4586 6054
rect 4822 5818 5004 6054
rect 4404 5734 5004 5818
rect 4404 5498 4586 5734
rect 4822 5498 5004 5734
rect -3876 -2462 -3694 -2226
rect -3458 -2462 -3276 -2226
rect -3876 -2546 -3276 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 -3276 -2546
rect -3876 -2804 -3276 -2782
rect 4404 -2226 5004 5498
rect 4404 -2462 4586 -2226
rect 4822 -2462 5004 -2226
rect 4404 -2546 5004 -2462
rect 4404 -2782 4586 -2546
rect 4822 -2782 5004 -2546
rect -4816 -3402 -4634 -3166
rect -4398 -3402 -4216 -3166
rect -4816 -3486 -4216 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 -4216 -3486
rect -4816 -3744 -4216 -3722
rect 4404 -3744 5004 -2782
rect 8004 693654 8604 708042
rect 8004 693418 8186 693654
rect 8422 693418 8604 693654
rect 8004 693334 8604 693418
rect 8004 693098 8186 693334
rect 8422 693098 8604 693334
rect 8004 657654 8604 693098
rect 8004 657418 8186 657654
rect 8422 657418 8604 657654
rect 8004 657334 8604 657418
rect 8004 657098 8186 657334
rect 8422 657098 8604 657334
rect 8004 621654 8604 657098
rect 8004 621418 8186 621654
rect 8422 621418 8604 621654
rect 8004 621334 8604 621418
rect 8004 621098 8186 621334
rect 8422 621098 8604 621334
rect 8004 585654 8604 621098
rect 8004 585418 8186 585654
rect 8422 585418 8604 585654
rect 8004 585334 8604 585418
rect 8004 585098 8186 585334
rect 8422 585098 8604 585334
rect 8004 549654 8604 585098
rect 8004 549418 8186 549654
rect 8422 549418 8604 549654
rect 8004 549334 8604 549418
rect 8004 549098 8186 549334
rect 8422 549098 8604 549334
rect 8004 513654 8604 549098
rect 8004 513418 8186 513654
rect 8422 513418 8604 513654
rect 8004 513334 8604 513418
rect 8004 513098 8186 513334
rect 8422 513098 8604 513334
rect 8004 477654 8604 513098
rect 8004 477418 8186 477654
rect 8422 477418 8604 477654
rect 8004 477334 8604 477418
rect 8004 477098 8186 477334
rect 8422 477098 8604 477334
rect 8004 441654 8604 477098
rect 8004 441418 8186 441654
rect 8422 441418 8604 441654
rect 8004 441334 8604 441418
rect 8004 441098 8186 441334
rect 8422 441098 8604 441334
rect 8004 405654 8604 441098
rect 8004 405418 8186 405654
rect 8422 405418 8604 405654
rect 8004 405334 8604 405418
rect 8004 405098 8186 405334
rect 8422 405098 8604 405334
rect 8004 369654 8604 405098
rect 8004 369418 8186 369654
rect 8422 369418 8604 369654
rect 8004 369334 8604 369418
rect 8004 369098 8186 369334
rect 8422 369098 8604 369334
rect 8004 333654 8604 369098
rect 8004 333418 8186 333654
rect 8422 333418 8604 333654
rect 8004 333334 8604 333418
rect 8004 333098 8186 333334
rect 8422 333098 8604 333334
rect 8004 297654 8604 333098
rect 8004 297418 8186 297654
rect 8422 297418 8604 297654
rect 8004 297334 8604 297418
rect 8004 297098 8186 297334
rect 8422 297098 8604 297334
rect 8004 261654 8604 297098
rect 8004 261418 8186 261654
rect 8422 261418 8604 261654
rect 8004 261334 8604 261418
rect 8004 261098 8186 261334
rect 8422 261098 8604 261334
rect 8004 225654 8604 261098
rect 8004 225418 8186 225654
rect 8422 225418 8604 225654
rect 8004 225334 8604 225418
rect 8004 225098 8186 225334
rect 8422 225098 8604 225334
rect 8004 189654 8604 225098
rect 8004 189418 8186 189654
rect 8422 189418 8604 189654
rect 8004 189334 8604 189418
rect 8004 189098 8186 189334
rect 8422 189098 8604 189334
rect 8004 153654 8604 189098
rect 8004 153418 8186 153654
rect 8422 153418 8604 153654
rect 8004 153334 8604 153418
rect 8004 153098 8186 153334
rect 8422 153098 8604 153334
rect 8004 117654 8604 153098
rect 8004 117418 8186 117654
rect 8422 117418 8604 117654
rect 8004 117334 8604 117418
rect 8004 117098 8186 117334
rect 8422 117098 8604 117334
rect 8004 81654 8604 117098
rect 11604 697254 12204 709922
rect 29604 711418 30204 711440
rect 29604 711182 29786 711418
rect 30022 711182 30204 711418
rect 29604 711098 30204 711182
rect 29604 710862 29786 711098
rect 30022 710862 30204 711098
rect 26004 709538 26604 709560
rect 26004 709302 26186 709538
rect 26422 709302 26604 709538
rect 26004 709218 26604 709302
rect 26004 708982 26186 709218
rect 26422 708982 26604 709218
rect 22404 707658 23004 707680
rect 22404 707422 22586 707658
rect 22822 707422 23004 707658
rect 22404 707338 23004 707422
rect 22404 707102 22586 707338
rect 22822 707102 23004 707338
rect 11604 697018 11786 697254
rect 12022 697018 12204 697254
rect 11604 696934 12204 697018
rect 11604 696698 11786 696934
rect 12022 696698 12204 696934
rect 11604 661254 12204 696698
rect 11604 661018 11786 661254
rect 12022 661018 12204 661254
rect 11604 660934 12204 661018
rect 11604 660698 11786 660934
rect 12022 660698 12204 660934
rect 11604 625254 12204 660698
rect 11604 625018 11786 625254
rect 12022 625018 12204 625254
rect 11604 624934 12204 625018
rect 11604 624698 11786 624934
rect 12022 624698 12204 624934
rect 11604 589254 12204 624698
rect 11604 589018 11786 589254
rect 12022 589018 12204 589254
rect 11604 588934 12204 589018
rect 11604 588698 11786 588934
rect 12022 588698 12204 588934
rect 11604 553254 12204 588698
rect 11604 553018 11786 553254
rect 12022 553018 12204 553254
rect 11604 552934 12204 553018
rect 11604 552698 11786 552934
rect 12022 552698 12204 552934
rect 11604 517254 12204 552698
rect 11604 517018 11786 517254
rect 12022 517018 12204 517254
rect 11604 516934 12204 517018
rect 11604 516698 11786 516934
rect 12022 516698 12204 516934
rect 11604 481254 12204 516698
rect 11604 481018 11786 481254
rect 12022 481018 12204 481254
rect 11604 480934 12204 481018
rect 11604 480698 11786 480934
rect 12022 480698 12204 480934
rect 11604 445254 12204 480698
rect 11604 445018 11786 445254
rect 12022 445018 12204 445254
rect 11604 444934 12204 445018
rect 11604 444698 11786 444934
rect 12022 444698 12204 444934
rect 11604 409254 12204 444698
rect 11604 409018 11786 409254
rect 12022 409018 12204 409254
rect 11604 408934 12204 409018
rect 11604 408698 11786 408934
rect 12022 408698 12204 408934
rect 11604 373254 12204 408698
rect 11604 373018 11786 373254
rect 12022 373018 12204 373254
rect 11604 372934 12204 373018
rect 11604 372698 11786 372934
rect 12022 372698 12204 372934
rect 11604 337254 12204 372698
rect 11604 337018 11786 337254
rect 12022 337018 12204 337254
rect 11604 336934 12204 337018
rect 11604 336698 11786 336934
rect 12022 336698 12204 336934
rect 11604 301254 12204 336698
rect 11604 301018 11786 301254
rect 12022 301018 12204 301254
rect 11604 300934 12204 301018
rect 11604 300698 11786 300934
rect 12022 300698 12204 300934
rect 11604 265254 12204 300698
rect 11604 265018 11786 265254
rect 12022 265018 12204 265254
rect 11604 264934 12204 265018
rect 11604 264698 11786 264934
rect 12022 264698 12204 264934
rect 11604 229254 12204 264698
rect 11604 229018 11786 229254
rect 12022 229018 12204 229254
rect 11604 228934 12204 229018
rect 11604 228698 11786 228934
rect 12022 228698 12204 228934
rect 11604 193254 12204 228698
rect 11604 193018 11786 193254
rect 12022 193018 12204 193254
rect 11604 192934 12204 193018
rect 11604 192698 11786 192934
rect 12022 192698 12204 192934
rect 11604 157254 12204 192698
rect 11604 157018 11786 157254
rect 12022 157018 12204 157254
rect 11604 156934 12204 157018
rect 11604 156698 11786 156934
rect 12022 156698 12204 156934
rect 11604 121254 12204 156698
rect 11604 121018 11786 121254
rect 12022 121018 12204 121254
rect 11604 120934 12204 121018
rect 11604 120698 11786 120934
rect 12022 120698 12204 120934
rect 9627 93804 9693 93805
rect 9627 93740 9628 93804
rect 9692 93740 9693 93804
rect 9627 93739 9693 93740
rect 9630 93397 9690 93739
rect 9627 93396 9693 93397
rect 9627 93332 9628 93396
rect 9692 93332 9693 93396
rect 9627 93331 9693 93332
rect 8004 81418 8186 81654
rect 8422 81418 8604 81654
rect 8004 81334 8604 81418
rect 8004 81098 8186 81334
rect 8422 81098 8604 81334
rect 8004 45654 8604 81098
rect 8004 45418 8186 45654
rect 8422 45418 8604 45654
rect 8004 45334 8604 45418
rect 8004 45098 8186 45334
rect 8422 45098 8604 45334
rect 8004 9654 8604 45098
rect 8004 9418 8186 9654
rect 8422 9418 8604 9654
rect 8004 9334 8604 9418
rect 8004 9098 8186 9334
rect 8422 9098 8604 9334
rect -5756 -4342 -5574 -4106
rect -5338 -4342 -5156 -4106
rect -5756 -4426 -5156 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 -5156 -4426
rect -5756 -4684 -5156 -4662
rect 8004 -4106 8604 9098
rect 8004 -4342 8186 -4106
rect 8422 -4342 8604 -4106
rect 8004 -4426 8604 -4342
rect 8004 -4662 8186 -4426
rect 8422 -4662 8604 -4426
rect -6696 -5282 -6514 -5046
rect -6278 -5282 -6096 -5046
rect -6696 -5366 -6096 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 -6096 -5366
rect -6696 -5624 -6096 -5602
rect 8004 -5624 8604 -4662
rect 11604 85254 12204 120698
rect 11604 85018 11786 85254
rect 12022 85018 12204 85254
rect 11604 84934 12204 85018
rect 11604 84698 11786 84934
rect 12022 84698 12204 84934
rect 11604 49254 12204 84698
rect 11604 49018 11786 49254
rect 12022 49018 12204 49254
rect 11604 48934 12204 49018
rect 11604 48698 11786 48934
rect 12022 48698 12204 48934
rect 11604 13254 12204 48698
rect 11604 13018 11786 13254
rect 12022 13018 12204 13254
rect 11604 12934 12204 13018
rect 11604 12698 11786 12934
rect 12022 12698 12204 12934
rect -7636 -6222 -7454 -5986
rect -7218 -6222 -7036 -5986
rect -7636 -6306 -7036 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 -7036 -6306
rect -7636 -6564 -7036 -6542
rect 11604 -5986 12204 12698
rect 18804 705778 19404 705800
rect 18804 705542 18986 705778
rect 19222 705542 19404 705778
rect 18804 705458 19404 705542
rect 18804 705222 18986 705458
rect 19222 705222 19404 705458
rect 18804 668454 19404 705222
rect 18804 668218 18986 668454
rect 19222 668218 19404 668454
rect 18804 668134 19404 668218
rect 18804 667898 18986 668134
rect 19222 667898 19404 668134
rect 18804 632454 19404 667898
rect 18804 632218 18986 632454
rect 19222 632218 19404 632454
rect 18804 632134 19404 632218
rect 18804 631898 18986 632134
rect 19222 631898 19404 632134
rect 18804 596454 19404 631898
rect 18804 596218 18986 596454
rect 19222 596218 19404 596454
rect 18804 596134 19404 596218
rect 18804 595898 18986 596134
rect 19222 595898 19404 596134
rect 18804 560454 19404 595898
rect 18804 560218 18986 560454
rect 19222 560218 19404 560454
rect 18804 560134 19404 560218
rect 18804 559898 18986 560134
rect 19222 559898 19404 560134
rect 18804 524454 19404 559898
rect 18804 524218 18986 524454
rect 19222 524218 19404 524454
rect 18804 524134 19404 524218
rect 18804 523898 18986 524134
rect 19222 523898 19404 524134
rect 18804 488454 19404 523898
rect 18804 488218 18986 488454
rect 19222 488218 19404 488454
rect 18804 488134 19404 488218
rect 18804 487898 18986 488134
rect 19222 487898 19404 488134
rect 18804 452454 19404 487898
rect 18804 452218 18986 452454
rect 19222 452218 19404 452454
rect 18804 452134 19404 452218
rect 18804 451898 18986 452134
rect 19222 451898 19404 452134
rect 18804 416454 19404 451898
rect 18804 416218 18986 416454
rect 19222 416218 19404 416454
rect 18804 416134 19404 416218
rect 18804 415898 18986 416134
rect 19222 415898 19404 416134
rect 18804 380454 19404 415898
rect 18804 380218 18986 380454
rect 19222 380218 19404 380454
rect 18804 380134 19404 380218
rect 18804 379898 18986 380134
rect 19222 379898 19404 380134
rect 18804 344454 19404 379898
rect 18804 344218 18986 344454
rect 19222 344218 19404 344454
rect 18804 344134 19404 344218
rect 18804 343898 18986 344134
rect 19222 343898 19404 344134
rect 18804 308454 19404 343898
rect 18804 308218 18986 308454
rect 19222 308218 19404 308454
rect 18804 308134 19404 308218
rect 18804 307898 18986 308134
rect 19222 307898 19404 308134
rect 18804 272454 19404 307898
rect 18804 272218 18986 272454
rect 19222 272218 19404 272454
rect 18804 272134 19404 272218
rect 18804 271898 18986 272134
rect 19222 271898 19404 272134
rect 18804 236454 19404 271898
rect 18804 236218 18986 236454
rect 19222 236218 19404 236454
rect 18804 236134 19404 236218
rect 18804 235898 18986 236134
rect 19222 235898 19404 236134
rect 18804 200454 19404 235898
rect 18804 200218 18986 200454
rect 19222 200218 19404 200454
rect 18804 200134 19404 200218
rect 18804 199898 18986 200134
rect 19222 199898 19404 200134
rect 18804 164454 19404 199898
rect 18804 164218 18986 164454
rect 19222 164218 19404 164454
rect 18804 164134 19404 164218
rect 18804 163898 18986 164134
rect 19222 163898 19404 164134
rect 18804 128454 19404 163898
rect 18804 128218 18986 128454
rect 19222 128218 19404 128454
rect 18804 128134 19404 128218
rect 18804 127898 18986 128134
rect 19222 127898 19404 128134
rect 18804 92454 19404 127898
rect 18804 92218 18986 92454
rect 19222 92218 19404 92454
rect 18804 92134 19404 92218
rect 18804 91898 18986 92134
rect 19222 91898 19404 92134
rect 18804 56454 19404 91898
rect 18804 56218 18986 56454
rect 19222 56218 19404 56454
rect 18804 56134 19404 56218
rect 18804 55898 18986 56134
rect 19222 55898 19404 56134
rect 18804 20454 19404 55898
rect 18804 20218 18986 20454
rect 19222 20218 19404 20454
rect 18804 20134 19404 20218
rect 18804 19898 18986 20134
rect 19222 19898 19404 20134
rect 18804 -1286 19404 19898
rect 18804 -1522 18986 -1286
rect 19222 -1522 19404 -1286
rect 18804 -1606 19404 -1522
rect 18804 -1842 18986 -1606
rect 19222 -1842 19404 -1606
rect 18804 -1864 19404 -1842
rect 22404 672054 23004 707102
rect 22404 671818 22586 672054
rect 22822 671818 23004 672054
rect 22404 671734 23004 671818
rect 22404 671498 22586 671734
rect 22822 671498 23004 671734
rect 22404 636054 23004 671498
rect 22404 635818 22586 636054
rect 22822 635818 23004 636054
rect 22404 635734 23004 635818
rect 22404 635498 22586 635734
rect 22822 635498 23004 635734
rect 22404 600054 23004 635498
rect 22404 599818 22586 600054
rect 22822 599818 23004 600054
rect 22404 599734 23004 599818
rect 22404 599498 22586 599734
rect 22822 599498 23004 599734
rect 22404 564054 23004 599498
rect 22404 563818 22586 564054
rect 22822 563818 23004 564054
rect 22404 563734 23004 563818
rect 22404 563498 22586 563734
rect 22822 563498 23004 563734
rect 22404 528054 23004 563498
rect 22404 527818 22586 528054
rect 22822 527818 23004 528054
rect 22404 527734 23004 527818
rect 22404 527498 22586 527734
rect 22822 527498 23004 527734
rect 22404 492054 23004 527498
rect 22404 491818 22586 492054
rect 22822 491818 23004 492054
rect 22404 491734 23004 491818
rect 22404 491498 22586 491734
rect 22822 491498 23004 491734
rect 22404 456054 23004 491498
rect 22404 455818 22586 456054
rect 22822 455818 23004 456054
rect 22404 455734 23004 455818
rect 22404 455498 22586 455734
rect 22822 455498 23004 455734
rect 22404 420054 23004 455498
rect 22404 419818 22586 420054
rect 22822 419818 23004 420054
rect 22404 419734 23004 419818
rect 22404 419498 22586 419734
rect 22822 419498 23004 419734
rect 22404 384054 23004 419498
rect 22404 383818 22586 384054
rect 22822 383818 23004 384054
rect 22404 383734 23004 383818
rect 22404 383498 22586 383734
rect 22822 383498 23004 383734
rect 22404 348054 23004 383498
rect 22404 347818 22586 348054
rect 22822 347818 23004 348054
rect 22404 347734 23004 347818
rect 22404 347498 22586 347734
rect 22822 347498 23004 347734
rect 22404 312054 23004 347498
rect 22404 311818 22586 312054
rect 22822 311818 23004 312054
rect 22404 311734 23004 311818
rect 22404 311498 22586 311734
rect 22822 311498 23004 311734
rect 22404 276054 23004 311498
rect 22404 275818 22586 276054
rect 22822 275818 23004 276054
rect 22404 275734 23004 275818
rect 22404 275498 22586 275734
rect 22822 275498 23004 275734
rect 22404 240054 23004 275498
rect 22404 239818 22586 240054
rect 22822 239818 23004 240054
rect 22404 239734 23004 239818
rect 22404 239498 22586 239734
rect 22822 239498 23004 239734
rect 22404 204054 23004 239498
rect 22404 203818 22586 204054
rect 22822 203818 23004 204054
rect 22404 203734 23004 203818
rect 22404 203498 22586 203734
rect 22822 203498 23004 203734
rect 22404 168054 23004 203498
rect 22404 167818 22586 168054
rect 22822 167818 23004 168054
rect 22404 167734 23004 167818
rect 22404 167498 22586 167734
rect 22822 167498 23004 167734
rect 22404 132054 23004 167498
rect 22404 131818 22586 132054
rect 22822 131818 23004 132054
rect 22404 131734 23004 131818
rect 22404 131498 22586 131734
rect 22822 131498 23004 131734
rect 22404 96054 23004 131498
rect 22404 95818 22586 96054
rect 22822 95818 23004 96054
rect 22404 95734 23004 95818
rect 22404 95498 22586 95734
rect 22822 95498 23004 95734
rect 22404 60054 23004 95498
rect 22404 59818 22586 60054
rect 22822 59818 23004 60054
rect 22404 59734 23004 59818
rect 22404 59498 22586 59734
rect 22822 59498 23004 59734
rect 22404 24054 23004 59498
rect 22404 23818 22586 24054
rect 22822 23818 23004 24054
rect 22404 23734 23004 23818
rect 22404 23498 22586 23734
rect 22822 23498 23004 23734
rect 22404 -3166 23004 23498
rect 22404 -3402 22586 -3166
rect 22822 -3402 23004 -3166
rect 22404 -3486 23004 -3402
rect 22404 -3722 22586 -3486
rect 22822 -3722 23004 -3486
rect 22404 -3744 23004 -3722
rect 26004 675654 26604 708982
rect 26004 675418 26186 675654
rect 26422 675418 26604 675654
rect 26004 675334 26604 675418
rect 26004 675098 26186 675334
rect 26422 675098 26604 675334
rect 26004 639654 26604 675098
rect 26004 639418 26186 639654
rect 26422 639418 26604 639654
rect 26004 639334 26604 639418
rect 26004 639098 26186 639334
rect 26422 639098 26604 639334
rect 26004 603654 26604 639098
rect 26004 603418 26186 603654
rect 26422 603418 26604 603654
rect 26004 603334 26604 603418
rect 26004 603098 26186 603334
rect 26422 603098 26604 603334
rect 26004 567654 26604 603098
rect 26004 567418 26186 567654
rect 26422 567418 26604 567654
rect 26004 567334 26604 567418
rect 26004 567098 26186 567334
rect 26422 567098 26604 567334
rect 26004 531654 26604 567098
rect 26004 531418 26186 531654
rect 26422 531418 26604 531654
rect 26004 531334 26604 531418
rect 26004 531098 26186 531334
rect 26422 531098 26604 531334
rect 26004 495654 26604 531098
rect 26004 495418 26186 495654
rect 26422 495418 26604 495654
rect 26004 495334 26604 495418
rect 26004 495098 26186 495334
rect 26422 495098 26604 495334
rect 26004 459654 26604 495098
rect 26004 459418 26186 459654
rect 26422 459418 26604 459654
rect 26004 459334 26604 459418
rect 26004 459098 26186 459334
rect 26422 459098 26604 459334
rect 26004 423654 26604 459098
rect 26004 423418 26186 423654
rect 26422 423418 26604 423654
rect 26004 423334 26604 423418
rect 26004 423098 26186 423334
rect 26422 423098 26604 423334
rect 26004 387654 26604 423098
rect 26004 387418 26186 387654
rect 26422 387418 26604 387654
rect 26004 387334 26604 387418
rect 26004 387098 26186 387334
rect 26422 387098 26604 387334
rect 26004 351654 26604 387098
rect 26004 351418 26186 351654
rect 26422 351418 26604 351654
rect 26004 351334 26604 351418
rect 26004 351098 26186 351334
rect 26422 351098 26604 351334
rect 26004 315654 26604 351098
rect 26004 315418 26186 315654
rect 26422 315418 26604 315654
rect 26004 315334 26604 315418
rect 26004 315098 26186 315334
rect 26422 315098 26604 315334
rect 26004 279654 26604 315098
rect 26004 279418 26186 279654
rect 26422 279418 26604 279654
rect 26004 279334 26604 279418
rect 26004 279098 26186 279334
rect 26422 279098 26604 279334
rect 26004 243654 26604 279098
rect 26004 243418 26186 243654
rect 26422 243418 26604 243654
rect 26004 243334 26604 243418
rect 26004 243098 26186 243334
rect 26422 243098 26604 243334
rect 26004 207654 26604 243098
rect 26004 207418 26186 207654
rect 26422 207418 26604 207654
rect 26004 207334 26604 207418
rect 26004 207098 26186 207334
rect 26422 207098 26604 207334
rect 26004 171654 26604 207098
rect 26004 171418 26186 171654
rect 26422 171418 26604 171654
rect 26004 171334 26604 171418
rect 26004 171098 26186 171334
rect 26422 171098 26604 171334
rect 26004 135654 26604 171098
rect 26004 135418 26186 135654
rect 26422 135418 26604 135654
rect 26004 135334 26604 135418
rect 26004 135098 26186 135334
rect 26422 135098 26604 135334
rect 26004 99654 26604 135098
rect 26004 99418 26186 99654
rect 26422 99418 26604 99654
rect 26004 99334 26604 99418
rect 26004 99098 26186 99334
rect 26422 99098 26604 99334
rect 26004 63654 26604 99098
rect 29604 679254 30204 710862
rect 47604 710478 48204 711440
rect 47604 710242 47786 710478
rect 48022 710242 48204 710478
rect 47604 710158 48204 710242
rect 47604 709922 47786 710158
rect 48022 709922 48204 710158
rect 44004 708598 44604 709560
rect 44004 708362 44186 708598
rect 44422 708362 44604 708598
rect 44004 708278 44604 708362
rect 44004 708042 44186 708278
rect 44422 708042 44604 708278
rect 40404 706718 41004 707680
rect 40404 706482 40586 706718
rect 40822 706482 41004 706718
rect 40404 706398 41004 706482
rect 40404 706162 40586 706398
rect 40822 706162 41004 706398
rect 29604 679018 29786 679254
rect 30022 679018 30204 679254
rect 29604 678934 30204 679018
rect 29604 678698 29786 678934
rect 30022 678698 30204 678934
rect 29604 643254 30204 678698
rect 29604 643018 29786 643254
rect 30022 643018 30204 643254
rect 29604 642934 30204 643018
rect 29604 642698 29786 642934
rect 30022 642698 30204 642934
rect 29604 607254 30204 642698
rect 29604 607018 29786 607254
rect 30022 607018 30204 607254
rect 29604 606934 30204 607018
rect 29604 606698 29786 606934
rect 30022 606698 30204 606934
rect 29604 571254 30204 606698
rect 29604 571018 29786 571254
rect 30022 571018 30204 571254
rect 29604 570934 30204 571018
rect 29604 570698 29786 570934
rect 30022 570698 30204 570934
rect 29604 535254 30204 570698
rect 29604 535018 29786 535254
rect 30022 535018 30204 535254
rect 29604 534934 30204 535018
rect 29604 534698 29786 534934
rect 30022 534698 30204 534934
rect 29604 499254 30204 534698
rect 29604 499018 29786 499254
rect 30022 499018 30204 499254
rect 29604 498934 30204 499018
rect 29604 498698 29786 498934
rect 30022 498698 30204 498934
rect 29604 463254 30204 498698
rect 29604 463018 29786 463254
rect 30022 463018 30204 463254
rect 29604 462934 30204 463018
rect 29604 462698 29786 462934
rect 30022 462698 30204 462934
rect 29604 427254 30204 462698
rect 29604 427018 29786 427254
rect 30022 427018 30204 427254
rect 29604 426934 30204 427018
rect 29604 426698 29786 426934
rect 30022 426698 30204 426934
rect 29604 391254 30204 426698
rect 29604 391018 29786 391254
rect 30022 391018 30204 391254
rect 29604 390934 30204 391018
rect 29604 390698 29786 390934
rect 30022 390698 30204 390934
rect 29604 355254 30204 390698
rect 29604 355018 29786 355254
rect 30022 355018 30204 355254
rect 29604 354934 30204 355018
rect 29604 354698 29786 354934
rect 30022 354698 30204 354934
rect 29604 319254 30204 354698
rect 29604 319018 29786 319254
rect 30022 319018 30204 319254
rect 29604 318934 30204 319018
rect 29604 318698 29786 318934
rect 30022 318698 30204 318934
rect 29604 283254 30204 318698
rect 29604 283018 29786 283254
rect 30022 283018 30204 283254
rect 29604 282934 30204 283018
rect 29604 282698 29786 282934
rect 30022 282698 30204 282934
rect 29604 247254 30204 282698
rect 29604 247018 29786 247254
rect 30022 247018 30204 247254
rect 29604 246934 30204 247018
rect 29604 246698 29786 246934
rect 30022 246698 30204 246934
rect 29604 211254 30204 246698
rect 29604 211018 29786 211254
rect 30022 211018 30204 211254
rect 29604 210934 30204 211018
rect 29604 210698 29786 210934
rect 30022 210698 30204 210934
rect 29604 175254 30204 210698
rect 29604 175018 29786 175254
rect 30022 175018 30204 175254
rect 29604 174934 30204 175018
rect 29604 174698 29786 174934
rect 30022 174698 30204 174934
rect 29604 139254 30204 174698
rect 29604 139018 29786 139254
rect 30022 139018 30204 139254
rect 29604 138934 30204 139018
rect 29604 138698 29786 138934
rect 30022 138698 30204 138934
rect 29604 103254 30204 138698
rect 29604 103018 29786 103254
rect 30022 103018 30204 103254
rect 29604 102934 30204 103018
rect 29604 102698 29786 102934
rect 30022 102698 30204 102934
rect 28947 93668 29013 93669
rect 28947 93604 28948 93668
rect 29012 93604 29013 93668
rect 28947 93603 29013 93604
rect 28950 93261 29010 93603
rect 28947 93260 29013 93261
rect 28947 93196 28948 93260
rect 29012 93196 29013 93260
rect 28947 93195 29013 93196
rect 26004 63418 26186 63654
rect 26422 63418 26604 63654
rect 26004 63334 26604 63418
rect 26004 63098 26186 63334
rect 26422 63098 26604 63334
rect 26004 27654 26604 63098
rect 26004 27418 26186 27654
rect 26422 27418 26604 27654
rect 26004 27334 26604 27418
rect 26004 27098 26186 27334
rect 26422 27098 26604 27334
rect 26004 -5046 26604 27098
rect 26004 -5282 26186 -5046
rect 26422 -5282 26604 -5046
rect 26004 -5366 26604 -5282
rect 26004 -5602 26186 -5366
rect 26422 -5602 26604 -5366
rect 26004 -5624 26604 -5602
rect 29604 67254 30204 102698
rect 29604 67018 29786 67254
rect 30022 67018 30204 67254
rect 29604 66934 30204 67018
rect 29604 66698 29786 66934
rect 30022 66698 30204 66934
rect 29604 31254 30204 66698
rect 29604 31018 29786 31254
rect 30022 31018 30204 31254
rect 29604 30934 30204 31018
rect 29604 30698 29786 30934
rect 30022 30698 30204 30934
rect 11604 -6222 11786 -5986
rect 12022 -6222 12204 -5986
rect 11604 -6306 12204 -6222
rect 11604 -6542 11786 -6306
rect 12022 -6542 12204 -6306
rect -8576 -7162 -8394 -6926
rect -8158 -7162 -7976 -6926
rect -8576 -7246 -7976 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 -7976 -7246
rect -8576 -7504 -7976 -7482
rect 11604 -7504 12204 -6542
rect 29604 -6926 30204 30698
rect 36804 704838 37404 705800
rect 36804 704602 36986 704838
rect 37222 704602 37404 704838
rect 36804 704518 37404 704602
rect 36804 704282 36986 704518
rect 37222 704282 37404 704518
rect 36804 686454 37404 704282
rect 36804 686218 36986 686454
rect 37222 686218 37404 686454
rect 36804 686134 37404 686218
rect 36804 685898 36986 686134
rect 37222 685898 37404 686134
rect 36804 650454 37404 685898
rect 36804 650218 36986 650454
rect 37222 650218 37404 650454
rect 36804 650134 37404 650218
rect 36804 649898 36986 650134
rect 37222 649898 37404 650134
rect 36804 614454 37404 649898
rect 36804 614218 36986 614454
rect 37222 614218 37404 614454
rect 36804 614134 37404 614218
rect 36804 613898 36986 614134
rect 37222 613898 37404 614134
rect 36804 578454 37404 613898
rect 36804 578218 36986 578454
rect 37222 578218 37404 578454
rect 36804 578134 37404 578218
rect 36804 577898 36986 578134
rect 37222 577898 37404 578134
rect 36804 542454 37404 577898
rect 36804 542218 36986 542454
rect 37222 542218 37404 542454
rect 36804 542134 37404 542218
rect 36804 541898 36986 542134
rect 37222 541898 37404 542134
rect 36804 506454 37404 541898
rect 36804 506218 36986 506454
rect 37222 506218 37404 506454
rect 36804 506134 37404 506218
rect 36804 505898 36986 506134
rect 37222 505898 37404 506134
rect 36804 470454 37404 505898
rect 36804 470218 36986 470454
rect 37222 470218 37404 470454
rect 36804 470134 37404 470218
rect 36804 469898 36986 470134
rect 37222 469898 37404 470134
rect 36804 434454 37404 469898
rect 36804 434218 36986 434454
rect 37222 434218 37404 434454
rect 36804 434134 37404 434218
rect 36804 433898 36986 434134
rect 37222 433898 37404 434134
rect 36804 398454 37404 433898
rect 36804 398218 36986 398454
rect 37222 398218 37404 398454
rect 36804 398134 37404 398218
rect 36804 397898 36986 398134
rect 37222 397898 37404 398134
rect 36804 362454 37404 397898
rect 36804 362218 36986 362454
rect 37222 362218 37404 362454
rect 36804 362134 37404 362218
rect 36804 361898 36986 362134
rect 37222 361898 37404 362134
rect 36804 326454 37404 361898
rect 36804 326218 36986 326454
rect 37222 326218 37404 326454
rect 36804 326134 37404 326218
rect 36804 325898 36986 326134
rect 37222 325898 37404 326134
rect 36804 290454 37404 325898
rect 36804 290218 36986 290454
rect 37222 290218 37404 290454
rect 36804 290134 37404 290218
rect 36804 289898 36986 290134
rect 37222 289898 37404 290134
rect 36804 254454 37404 289898
rect 36804 254218 36986 254454
rect 37222 254218 37404 254454
rect 36804 254134 37404 254218
rect 36804 253898 36986 254134
rect 37222 253898 37404 254134
rect 36804 218454 37404 253898
rect 36804 218218 36986 218454
rect 37222 218218 37404 218454
rect 36804 218134 37404 218218
rect 36804 217898 36986 218134
rect 37222 217898 37404 218134
rect 36804 182454 37404 217898
rect 36804 182218 36986 182454
rect 37222 182218 37404 182454
rect 36804 182134 37404 182218
rect 36804 181898 36986 182134
rect 37222 181898 37404 182134
rect 36804 146454 37404 181898
rect 36804 146218 36986 146454
rect 37222 146218 37404 146454
rect 36804 146134 37404 146218
rect 36804 145898 36986 146134
rect 37222 145898 37404 146134
rect 36804 110454 37404 145898
rect 36804 110218 36986 110454
rect 37222 110218 37404 110454
rect 36804 110134 37404 110218
rect 36804 109898 36986 110134
rect 37222 109898 37404 110134
rect 36804 74454 37404 109898
rect 36804 74218 36986 74454
rect 37222 74218 37404 74454
rect 36804 74134 37404 74218
rect 36804 73898 36986 74134
rect 37222 73898 37404 74134
rect 36804 38454 37404 73898
rect 36804 38218 36986 38454
rect 37222 38218 37404 38454
rect 36804 38134 37404 38218
rect 36804 37898 36986 38134
rect 37222 37898 37404 38134
rect 36804 2454 37404 37898
rect 36804 2218 36986 2454
rect 37222 2218 37404 2454
rect 36804 2134 37404 2218
rect 36804 1898 36986 2134
rect 37222 1898 37404 2134
rect 36804 -346 37404 1898
rect 36804 -582 36986 -346
rect 37222 -582 37404 -346
rect 36804 -666 37404 -582
rect 36804 -902 36986 -666
rect 37222 -902 37404 -666
rect 36804 -1864 37404 -902
rect 40404 690054 41004 706162
rect 40404 689818 40586 690054
rect 40822 689818 41004 690054
rect 40404 689734 41004 689818
rect 40404 689498 40586 689734
rect 40822 689498 41004 689734
rect 40404 654054 41004 689498
rect 40404 653818 40586 654054
rect 40822 653818 41004 654054
rect 40404 653734 41004 653818
rect 40404 653498 40586 653734
rect 40822 653498 41004 653734
rect 40404 618054 41004 653498
rect 40404 617818 40586 618054
rect 40822 617818 41004 618054
rect 40404 617734 41004 617818
rect 40404 617498 40586 617734
rect 40822 617498 41004 617734
rect 40404 582054 41004 617498
rect 40404 581818 40586 582054
rect 40822 581818 41004 582054
rect 40404 581734 41004 581818
rect 40404 581498 40586 581734
rect 40822 581498 41004 581734
rect 40404 546054 41004 581498
rect 40404 545818 40586 546054
rect 40822 545818 41004 546054
rect 40404 545734 41004 545818
rect 40404 545498 40586 545734
rect 40822 545498 41004 545734
rect 40404 510054 41004 545498
rect 40404 509818 40586 510054
rect 40822 509818 41004 510054
rect 40404 509734 41004 509818
rect 40404 509498 40586 509734
rect 40822 509498 41004 509734
rect 40404 474054 41004 509498
rect 40404 473818 40586 474054
rect 40822 473818 41004 474054
rect 40404 473734 41004 473818
rect 40404 473498 40586 473734
rect 40822 473498 41004 473734
rect 40404 438054 41004 473498
rect 40404 437818 40586 438054
rect 40822 437818 41004 438054
rect 40404 437734 41004 437818
rect 40404 437498 40586 437734
rect 40822 437498 41004 437734
rect 40404 402054 41004 437498
rect 40404 401818 40586 402054
rect 40822 401818 41004 402054
rect 40404 401734 41004 401818
rect 40404 401498 40586 401734
rect 40822 401498 41004 401734
rect 40404 366054 41004 401498
rect 40404 365818 40586 366054
rect 40822 365818 41004 366054
rect 40404 365734 41004 365818
rect 40404 365498 40586 365734
rect 40822 365498 41004 365734
rect 40404 330054 41004 365498
rect 40404 329818 40586 330054
rect 40822 329818 41004 330054
rect 40404 329734 41004 329818
rect 40404 329498 40586 329734
rect 40822 329498 41004 329734
rect 40404 294054 41004 329498
rect 40404 293818 40586 294054
rect 40822 293818 41004 294054
rect 40404 293734 41004 293818
rect 40404 293498 40586 293734
rect 40822 293498 41004 293734
rect 40404 258054 41004 293498
rect 40404 257818 40586 258054
rect 40822 257818 41004 258054
rect 40404 257734 41004 257818
rect 40404 257498 40586 257734
rect 40822 257498 41004 257734
rect 40404 222054 41004 257498
rect 40404 221818 40586 222054
rect 40822 221818 41004 222054
rect 40404 221734 41004 221818
rect 40404 221498 40586 221734
rect 40822 221498 41004 221734
rect 40404 186054 41004 221498
rect 40404 185818 40586 186054
rect 40822 185818 41004 186054
rect 40404 185734 41004 185818
rect 40404 185498 40586 185734
rect 40822 185498 41004 185734
rect 40404 150054 41004 185498
rect 40404 149818 40586 150054
rect 40822 149818 41004 150054
rect 40404 149734 41004 149818
rect 40404 149498 40586 149734
rect 40822 149498 41004 149734
rect 40404 114054 41004 149498
rect 40404 113818 40586 114054
rect 40822 113818 41004 114054
rect 40404 113734 41004 113818
rect 40404 113498 40586 113734
rect 40822 113498 41004 113734
rect 40404 78054 41004 113498
rect 40404 77818 40586 78054
rect 40822 77818 41004 78054
rect 40404 77734 41004 77818
rect 40404 77498 40586 77734
rect 40822 77498 41004 77734
rect 40404 42054 41004 77498
rect 40404 41818 40586 42054
rect 40822 41818 41004 42054
rect 40404 41734 41004 41818
rect 40404 41498 40586 41734
rect 40822 41498 41004 41734
rect 40404 6054 41004 41498
rect 40404 5818 40586 6054
rect 40822 5818 41004 6054
rect 40404 5734 41004 5818
rect 40404 5498 40586 5734
rect 40822 5498 41004 5734
rect 40404 -2226 41004 5498
rect 40404 -2462 40586 -2226
rect 40822 -2462 41004 -2226
rect 40404 -2546 41004 -2462
rect 40404 -2782 40586 -2546
rect 40822 -2782 41004 -2546
rect 40404 -3744 41004 -2782
rect 44004 693654 44604 708042
rect 44004 693418 44186 693654
rect 44422 693418 44604 693654
rect 44004 693334 44604 693418
rect 44004 693098 44186 693334
rect 44422 693098 44604 693334
rect 44004 657654 44604 693098
rect 44004 657418 44186 657654
rect 44422 657418 44604 657654
rect 44004 657334 44604 657418
rect 44004 657098 44186 657334
rect 44422 657098 44604 657334
rect 44004 621654 44604 657098
rect 44004 621418 44186 621654
rect 44422 621418 44604 621654
rect 44004 621334 44604 621418
rect 44004 621098 44186 621334
rect 44422 621098 44604 621334
rect 44004 585654 44604 621098
rect 44004 585418 44186 585654
rect 44422 585418 44604 585654
rect 44004 585334 44604 585418
rect 44004 585098 44186 585334
rect 44422 585098 44604 585334
rect 44004 549654 44604 585098
rect 44004 549418 44186 549654
rect 44422 549418 44604 549654
rect 44004 549334 44604 549418
rect 44004 549098 44186 549334
rect 44422 549098 44604 549334
rect 44004 513654 44604 549098
rect 44004 513418 44186 513654
rect 44422 513418 44604 513654
rect 44004 513334 44604 513418
rect 44004 513098 44186 513334
rect 44422 513098 44604 513334
rect 44004 477654 44604 513098
rect 44004 477418 44186 477654
rect 44422 477418 44604 477654
rect 44004 477334 44604 477418
rect 44004 477098 44186 477334
rect 44422 477098 44604 477334
rect 44004 441654 44604 477098
rect 44004 441418 44186 441654
rect 44422 441418 44604 441654
rect 44004 441334 44604 441418
rect 44004 441098 44186 441334
rect 44422 441098 44604 441334
rect 44004 405654 44604 441098
rect 44004 405418 44186 405654
rect 44422 405418 44604 405654
rect 44004 405334 44604 405418
rect 44004 405098 44186 405334
rect 44422 405098 44604 405334
rect 44004 369654 44604 405098
rect 44004 369418 44186 369654
rect 44422 369418 44604 369654
rect 44004 369334 44604 369418
rect 44004 369098 44186 369334
rect 44422 369098 44604 369334
rect 44004 333654 44604 369098
rect 44004 333418 44186 333654
rect 44422 333418 44604 333654
rect 44004 333334 44604 333418
rect 44004 333098 44186 333334
rect 44422 333098 44604 333334
rect 44004 297654 44604 333098
rect 44004 297418 44186 297654
rect 44422 297418 44604 297654
rect 44004 297334 44604 297418
rect 44004 297098 44186 297334
rect 44422 297098 44604 297334
rect 44004 261654 44604 297098
rect 44004 261418 44186 261654
rect 44422 261418 44604 261654
rect 44004 261334 44604 261418
rect 44004 261098 44186 261334
rect 44422 261098 44604 261334
rect 44004 225654 44604 261098
rect 44004 225418 44186 225654
rect 44422 225418 44604 225654
rect 44004 225334 44604 225418
rect 44004 225098 44186 225334
rect 44422 225098 44604 225334
rect 44004 189654 44604 225098
rect 44004 189418 44186 189654
rect 44422 189418 44604 189654
rect 44004 189334 44604 189418
rect 44004 189098 44186 189334
rect 44422 189098 44604 189334
rect 44004 153654 44604 189098
rect 44004 153418 44186 153654
rect 44422 153418 44604 153654
rect 44004 153334 44604 153418
rect 44004 153098 44186 153334
rect 44422 153098 44604 153334
rect 44004 117654 44604 153098
rect 44004 117418 44186 117654
rect 44422 117418 44604 117654
rect 44004 117334 44604 117418
rect 44004 117098 44186 117334
rect 44422 117098 44604 117334
rect 44004 81654 44604 117098
rect 44004 81418 44186 81654
rect 44422 81418 44604 81654
rect 44004 81334 44604 81418
rect 44004 81098 44186 81334
rect 44422 81098 44604 81334
rect 44004 45654 44604 81098
rect 44004 45418 44186 45654
rect 44422 45418 44604 45654
rect 44004 45334 44604 45418
rect 44004 45098 44186 45334
rect 44422 45098 44604 45334
rect 44004 9654 44604 45098
rect 44004 9418 44186 9654
rect 44422 9418 44604 9654
rect 44004 9334 44604 9418
rect 44004 9098 44186 9334
rect 44422 9098 44604 9334
rect 44004 -4106 44604 9098
rect 44004 -4342 44186 -4106
rect 44422 -4342 44604 -4106
rect 44004 -4426 44604 -4342
rect 44004 -4662 44186 -4426
rect 44422 -4662 44604 -4426
rect 44004 -5624 44604 -4662
rect 47604 697254 48204 709922
rect 65604 711418 66204 711440
rect 65604 711182 65786 711418
rect 66022 711182 66204 711418
rect 65604 711098 66204 711182
rect 65604 710862 65786 711098
rect 66022 710862 66204 711098
rect 62004 709538 62604 709560
rect 62004 709302 62186 709538
rect 62422 709302 62604 709538
rect 62004 709218 62604 709302
rect 62004 708982 62186 709218
rect 62422 708982 62604 709218
rect 58404 707658 59004 707680
rect 58404 707422 58586 707658
rect 58822 707422 59004 707658
rect 58404 707338 59004 707422
rect 58404 707102 58586 707338
rect 58822 707102 59004 707338
rect 47604 697018 47786 697254
rect 48022 697018 48204 697254
rect 47604 696934 48204 697018
rect 47604 696698 47786 696934
rect 48022 696698 48204 696934
rect 47604 661254 48204 696698
rect 47604 661018 47786 661254
rect 48022 661018 48204 661254
rect 47604 660934 48204 661018
rect 47604 660698 47786 660934
rect 48022 660698 48204 660934
rect 47604 625254 48204 660698
rect 47604 625018 47786 625254
rect 48022 625018 48204 625254
rect 47604 624934 48204 625018
rect 47604 624698 47786 624934
rect 48022 624698 48204 624934
rect 47604 589254 48204 624698
rect 47604 589018 47786 589254
rect 48022 589018 48204 589254
rect 47604 588934 48204 589018
rect 47604 588698 47786 588934
rect 48022 588698 48204 588934
rect 47604 553254 48204 588698
rect 47604 553018 47786 553254
rect 48022 553018 48204 553254
rect 47604 552934 48204 553018
rect 47604 552698 47786 552934
rect 48022 552698 48204 552934
rect 47604 517254 48204 552698
rect 47604 517018 47786 517254
rect 48022 517018 48204 517254
rect 47604 516934 48204 517018
rect 47604 516698 47786 516934
rect 48022 516698 48204 516934
rect 47604 481254 48204 516698
rect 47604 481018 47786 481254
rect 48022 481018 48204 481254
rect 47604 480934 48204 481018
rect 47604 480698 47786 480934
rect 48022 480698 48204 480934
rect 47604 445254 48204 480698
rect 47604 445018 47786 445254
rect 48022 445018 48204 445254
rect 47604 444934 48204 445018
rect 47604 444698 47786 444934
rect 48022 444698 48204 444934
rect 47604 409254 48204 444698
rect 47604 409018 47786 409254
rect 48022 409018 48204 409254
rect 47604 408934 48204 409018
rect 47604 408698 47786 408934
rect 48022 408698 48204 408934
rect 47604 373254 48204 408698
rect 47604 373018 47786 373254
rect 48022 373018 48204 373254
rect 47604 372934 48204 373018
rect 47604 372698 47786 372934
rect 48022 372698 48204 372934
rect 47604 337254 48204 372698
rect 47604 337018 47786 337254
rect 48022 337018 48204 337254
rect 47604 336934 48204 337018
rect 47604 336698 47786 336934
rect 48022 336698 48204 336934
rect 47604 301254 48204 336698
rect 47604 301018 47786 301254
rect 48022 301018 48204 301254
rect 47604 300934 48204 301018
rect 47604 300698 47786 300934
rect 48022 300698 48204 300934
rect 47604 265254 48204 300698
rect 47604 265018 47786 265254
rect 48022 265018 48204 265254
rect 47604 264934 48204 265018
rect 47604 264698 47786 264934
rect 48022 264698 48204 264934
rect 47604 229254 48204 264698
rect 47604 229018 47786 229254
rect 48022 229018 48204 229254
rect 47604 228934 48204 229018
rect 47604 228698 47786 228934
rect 48022 228698 48204 228934
rect 47604 193254 48204 228698
rect 47604 193018 47786 193254
rect 48022 193018 48204 193254
rect 47604 192934 48204 193018
rect 47604 192698 47786 192934
rect 48022 192698 48204 192934
rect 47604 157254 48204 192698
rect 47604 157018 47786 157254
rect 48022 157018 48204 157254
rect 47604 156934 48204 157018
rect 47604 156698 47786 156934
rect 48022 156698 48204 156934
rect 47604 121254 48204 156698
rect 47604 121018 47786 121254
rect 48022 121018 48204 121254
rect 47604 120934 48204 121018
rect 47604 120698 47786 120934
rect 48022 120698 48204 120934
rect 47604 85254 48204 120698
rect 54804 705778 55404 705800
rect 54804 705542 54986 705778
rect 55222 705542 55404 705778
rect 54804 705458 55404 705542
rect 54804 705222 54986 705458
rect 55222 705222 55404 705458
rect 54804 668454 55404 705222
rect 54804 668218 54986 668454
rect 55222 668218 55404 668454
rect 54804 668134 55404 668218
rect 54804 667898 54986 668134
rect 55222 667898 55404 668134
rect 54804 632454 55404 667898
rect 54804 632218 54986 632454
rect 55222 632218 55404 632454
rect 54804 632134 55404 632218
rect 54804 631898 54986 632134
rect 55222 631898 55404 632134
rect 54804 596454 55404 631898
rect 54804 596218 54986 596454
rect 55222 596218 55404 596454
rect 54804 596134 55404 596218
rect 54804 595898 54986 596134
rect 55222 595898 55404 596134
rect 54804 560454 55404 595898
rect 54804 560218 54986 560454
rect 55222 560218 55404 560454
rect 54804 560134 55404 560218
rect 54804 559898 54986 560134
rect 55222 559898 55404 560134
rect 54804 524454 55404 559898
rect 54804 524218 54986 524454
rect 55222 524218 55404 524454
rect 54804 524134 55404 524218
rect 54804 523898 54986 524134
rect 55222 523898 55404 524134
rect 54804 488454 55404 523898
rect 54804 488218 54986 488454
rect 55222 488218 55404 488454
rect 54804 488134 55404 488218
rect 54804 487898 54986 488134
rect 55222 487898 55404 488134
rect 54804 452454 55404 487898
rect 54804 452218 54986 452454
rect 55222 452218 55404 452454
rect 54804 452134 55404 452218
rect 54804 451898 54986 452134
rect 55222 451898 55404 452134
rect 54804 416454 55404 451898
rect 54804 416218 54986 416454
rect 55222 416218 55404 416454
rect 54804 416134 55404 416218
rect 54804 415898 54986 416134
rect 55222 415898 55404 416134
rect 54804 380454 55404 415898
rect 54804 380218 54986 380454
rect 55222 380218 55404 380454
rect 54804 380134 55404 380218
rect 54804 379898 54986 380134
rect 55222 379898 55404 380134
rect 54804 344454 55404 379898
rect 54804 344218 54986 344454
rect 55222 344218 55404 344454
rect 54804 344134 55404 344218
rect 54804 343898 54986 344134
rect 55222 343898 55404 344134
rect 54804 308454 55404 343898
rect 54804 308218 54986 308454
rect 55222 308218 55404 308454
rect 54804 308134 55404 308218
rect 54804 307898 54986 308134
rect 55222 307898 55404 308134
rect 54804 272454 55404 307898
rect 54804 272218 54986 272454
rect 55222 272218 55404 272454
rect 54804 272134 55404 272218
rect 54804 271898 54986 272134
rect 55222 271898 55404 272134
rect 54804 236454 55404 271898
rect 54804 236218 54986 236454
rect 55222 236218 55404 236454
rect 54804 236134 55404 236218
rect 54804 235898 54986 236134
rect 55222 235898 55404 236134
rect 54804 200454 55404 235898
rect 54804 200218 54986 200454
rect 55222 200218 55404 200454
rect 54804 200134 55404 200218
rect 54804 199898 54986 200134
rect 55222 199898 55404 200134
rect 54804 164454 55404 199898
rect 54804 164218 54986 164454
rect 55222 164218 55404 164454
rect 54804 164134 55404 164218
rect 54804 163898 54986 164134
rect 55222 163898 55404 164134
rect 54804 128454 55404 163898
rect 54804 128218 54986 128454
rect 55222 128218 55404 128454
rect 54804 128134 55404 128218
rect 54804 127898 54986 128134
rect 55222 127898 55404 128134
rect 48267 93668 48333 93669
rect 48267 93604 48268 93668
rect 48332 93604 48333 93668
rect 48267 93603 48333 93604
rect 48270 93261 48330 93603
rect 48267 93260 48333 93261
rect 48267 93196 48268 93260
rect 48332 93196 48333 93260
rect 48267 93195 48333 93196
rect 47604 85018 47786 85254
rect 48022 85018 48204 85254
rect 47604 84934 48204 85018
rect 47604 84698 47786 84934
rect 48022 84698 48204 84934
rect 47604 49254 48204 84698
rect 47604 49018 47786 49254
rect 48022 49018 48204 49254
rect 47604 48934 48204 49018
rect 47604 48698 47786 48934
rect 48022 48698 48204 48934
rect 47604 13254 48204 48698
rect 47604 13018 47786 13254
rect 48022 13018 48204 13254
rect 47604 12934 48204 13018
rect 47604 12698 47786 12934
rect 48022 12698 48204 12934
rect 29604 -7162 29786 -6926
rect 30022 -7162 30204 -6926
rect 29604 -7246 30204 -7162
rect 29604 -7482 29786 -7246
rect 30022 -7482 30204 -7246
rect 29604 -7504 30204 -7482
rect 47604 -5986 48204 12698
rect 54804 92454 55404 127898
rect 58404 672054 59004 707102
rect 58404 671818 58586 672054
rect 58822 671818 59004 672054
rect 58404 671734 59004 671818
rect 58404 671498 58586 671734
rect 58822 671498 59004 671734
rect 58404 636054 59004 671498
rect 58404 635818 58586 636054
rect 58822 635818 59004 636054
rect 58404 635734 59004 635818
rect 58404 635498 58586 635734
rect 58822 635498 59004 635734
rect 58404 600054 59004 635498
rect 58404 599818 58586 600054
rect 58822 599818 59004 600054
rect 58404 599734 59004 599818
rect 58404 599498 58586 599734
rect 58822 599498 59004 599734
rect 58404 564054 59004 599498
rect 58404 563818 58586 564054
rect 58822 563818 59004 564054
rect 58404 563734 59004 563818
rect 58404 563498 58586 563734
rect 58822 563498 59004 563734
rect 58404 528054 59004 563498
rect 58404 527818 58586 528054
rect 58822 527818 59004 528054
rect 58404 527734 59004 527818
rect 58404 527498 58586 527734
rect 58822 527498 59004 527734
rect 58404 492054 59004 527498
rect 58404 491818 58586 492054
rect 58822 491818 59004 492054
rect 58404 491734 59004 491818
rect 58404 491498 58586 491734
rect 58822 491498 59004 491734
rect 58404 456054 59004 491498
rect 58404 455818 58586 456054
rect 58822 455818 59004 456054
rect 58404 455734 59004 455818
rect 58404 455498 58586 455734
rect 58822 455498 59004 455734
rect 58404 420054 59004 455498
rect 58404 419818 58586 420054
rect 58822 419818 59004 420054
rect 58404 419734 59004 419818
rect 58404 419498 58586 419734
rect 58822 419498 59004 419734
rect 58404 384054 59004 419498
rect 58404 383818 58586 384054
rect 58822 383818 59004 384054
rect 58404 383734 59004 383818
rect 58404 383498 58586 383734
rect 58822 383498 59004 383734
rect 58404 348054 59004 383498
rect 58404 347818 58586 348054
rect 58822 347818 59004 348054
rect 58404 347734 59004 347818
rect 58404 347498 58586 347734
rect 58822 347498 59004 347734
rect 58404 312054 59004 347498
rect 58404 311818 58586 312054
rect 58822 311818 59004 312054
rect 58404 311734 59004 311818
rect 58404 311498 58586 311734
rect 58822 311498 59004 311734
rect 58404 276054 59004 311498
rect 58404 275818 58586 276054
rect 58822 275818 59004 276054
rect 58404 275734 59004 275818
rect 58404 275498 58586 275734
rect 58822 275498 59004 275734
rect 58404 240054 59004 275498
rect 58404 239818 58586 240054
rect 58822 239818 59004 240054
rect 58404 239734 59004 239818
rect 58404 239498 58586 239734
rect 58822 239498 59004 239734
rect 58404 204054 59004 239498
rect 58404 203818 58586 204054
rect 58822 203818 59004 204054
rect 58404 203734 59004 203818
rect 58404 203498 58586 203734
rect 58822 203498 59004 203734
rect 58404 168054 59004 203498
rect 58404 167818 58586 168054
rect 58822 167818 59004 168054
rect 58404 167734 59004 167818
rect 58404 167498 58586 167734
rect 58822 167498 59004 167734
rect 58404 132054 59004 167498
rect 58404 131818 58586 132054
rect 58822 131818 59004 132054
rect 58404 131734 59004 131818
rect 58404 131498 58586 131734
rect 58822 131498 59004 131734
rect 58404 96054 59004 131498
rect 58404 95818 58586 96054
rect 58822 95818 59004 96054
rect 58404 95734 59004 95818
rect 58404 95498 58586 95734
rect 58822 95498 59004 95734
rect 57835 93532 57901 93533
rect 57835 93468 57836 93532
rect 57900 93468 57901 93532
rect 57835 93467 57901 93468
rect 57838 93261 57898 93467
rect 57835 93260 57901 93261
rect 57835 93196 57836 93260
rect 57900 93196 57901 93260
rect 57835 93195 57901 93196
rect 54804 92218 54986 92454
rect 55222 92218 55404 92454
rect 54804 92134 55404 92218
rect 54804 91898 54986 92134
rect 55222 91898 55404 92134
rect 54804 56454 55404 91898
rect 54804 56218 54986 56454
rect 55222 56218 55404 56454
rect 54804 56134 55404 56218
rect 54804 55898 54986 56134
rect 55222 55898 55404 56134
rect 54804 20454 55404 55898
rect 54804 20218 54986 20454
rect 55222 20218 55404 20454
rect 54804 20134 55404 20218
rect 54804 19898 54986 20134
rect 55222 19898 55404 20134
rect 54804 -1286 55404 19898
rect 54804 -1522 54986 -1286
rect 55222 -1522 55404 -1286
rect 54804 -1606 55404 -1522
rect 54804 -1842 54986 -1606
rect 55222 -1842 55404 -1606
rect 54804 -1864 55404 -1842
rect 58404 60054 59004 95498
rect 58404 59818 58586 60054
rect 58822 59818 59004 60054
rect 58404 59734 59004 59818
rect 58404 59498 58586 59734
rect 58822 59498 59004 59734
rect 58404 24054 59004 59498
rect 58404 23818 58586 24054
rect 58822 23818 59004 24054
rect 58404 23734 59004 23818
rect 58404 23498 58586 23734
rect 58822 23498 59004 23734
rect 58404 -3166 59004 23498
rect 58404 -3402 58586 -3166
rect 58822 -3402 59004 -3166
rect 58404 -3486 59004 -3402
rect 58404 -3722 58586 -3486
rect 58822 -3722 59004 -3486
rect 58404 -3744 59004 -3722
rect 62004 675654 62604 708982
rect 62004 675418 62186 675654
rect 62422 675418 62604 675654
rect 62004 675334 62604 675418
rect 62004 675098 62186 675334
rect 62422 675098 62604 675334
rect 62004 639654 62604 675098
rect 62004 639418 62186 639654
rect 62422 639418 62604 639654
rect 62004 639334 62604 639418
rect 62004 639098 62186 639334
rect 62422 639098 62604 639334
rect 62004 603654 62604 639098
rect 62004 603418 62186 603654
rect 62422 603418 62604 603654
rect 62004 603334 62604 603418
rect 62004 603098 62186 603334
rect 62422 603098 62604 603334
rect 62004 567654 62604 603098
rect 62004 567418 62186 567654
rect 62422 567418 62604 567654
rect 62004 567334 62604 567418
rect 62004 567098 62186 567334
rect 62422 567098 62604 567334
rect 62004 531654 62604 567098
rect 62004 531418 62186 531654
rect 62422 531418 62604 531654
rect 62004 531334 62604 531418
rect 62004 531098 62186 531334
rect 62422 531098 62604 531334
rect 62004 495654 62604 531098
rect 62004 495418 62186 495654
rect 62422 495418 62604 495654
rect 62004 495334 62604 495418
rect 62004 495098 62186 495334
rect 62422 495098 62604 495334
rect 62004 459654 62604 495098
rect 62004 459418 62186 459654
rect 62422 459418 62604 459654
rect 62004 459334 62604 459418
rect 62004 459098 62186 459334
rect 62422 459098 62604 459334
rect 62004 423654 62604 459098
rect 62004 423418 62186 423654
rect 62422 423418 62604 423654
rect 62004 423334 62604 423418
rect 62004 423098 62186 423334
rect 62422 423098 62604 423334
rect 62004 387654 62604 423098
rect 62004 387418 62186 387654
rect 62422 387418 62604 387654
rect 62004 387334 62604 387418
rect 62004 387098 62186 387334
rect 62422 387098 62604 387334
rect 62004 351654 62604 387098
rect 62004 351418 62186 351654
rect 62422 351418 62604 351654
rect 62004 351334 62604 351418
rect 62004 351098 62186 351334
rect 62422 351098 62604 351334
rect 62004 315654 62604 351098
rect 62004 315418 62186 315654
rect 62422 315418 62604 315654
rect 62004 315334 62604 315418
rect 62004 315098 62186 315334
rect 62422 315098 62604 315334
rect 62004 279654 62604 315098
rect 62004 279418 62186 279654
rect 62422 279418 62604 279654
rect 62004 279334 62604 279418
rect 62004 279098 62186 279334
rect 62422 279098 62604 279334
rect 62004 243654 62604 279098
rect 62004 243418 62186 243654
rect 62422 243418 62604 243654
rect 62004 243334 62604 243418
rect 62004 243098 62186 243334
rect 62422 243098 62604 243334
rect 62004 207654 62604 243098
rect 62004 207418 62186 207654
rect 62422 207418 62604 207654
rect 62004 207334 62604 207418
rect 62004 207098 62186 207334
rect 62422 207098 62604 207334
rect 62004 171654 62604 207098
rect 62004 171418 62186 171654
rect 62422 171418 62604 171654
rect 62004 171334 62604 171418
rect 62004 171098 62186 171334
rect 62422 171098 62604 171334
rect 62004 135654 62604 171098
rect 62004 135418 62186 135654
rect 62422 135418 62604 135654
rect 62004 135334 62604 135418
rect 62004 135098 62186 135334
rect 62422 135098 62604 135334
rect 62004 99654 62604 135098
rect 62004 99418 62186 99654
rect 62422 99418 62604 99654
rect 62004 99334 62604 99418
rect 62004 99098 62186 99334
rect 62422 99098 62604 99334
rect 62004 63654 62604 99098
rect 62004 63418 62186 63654
rect 62422 63418 62604 63654
rect 62004 63334 62604 63418
rect 62004 63098 62186 63334
rect 62422 63098 62604 63334
rect 62004 27654 62604 63098
rect 62004 27418 62186 27654
rect 62422 27418 62604 27654
rect 62004 27334 62604 27418
rect 62004 27098 62186 27334
rect 62422 27098 62604 27334
rect 62004 -5046 62604 27098
rect 62004 -5282 62186 -5046
rect 62422 -5282 62604 -5046
rect 62004 -5366 62604 -5282
rect 62004 -5602 62186 -5366
rect 62422 -5602 62604 -5366
rect 62004 -5624 62604 -5602
rect 65604 679254 66204 710862
rect 83604 710478 84204 711440
rect 83604 710242 83786 710478
rect 84022 710242 84204 710478
rect 83604 710158 84204 710242
rect 83604 709922 83786 710158
rect 84022 709922 84204 710158
rect 80004 708598 80604 709560
rect 80004 708362 80186 708598
rect 80422 708362 80604 708598
rect 80004 708278 80604 708362
rect 80004 708042 80186 708278
rect 80422 708042 80604 708278
rect 76404 706718 77004 707680
rect 76404 706482 76586 706718
rect 76822 706482 77004 706718
rect 76404 706398 77004 706482
rect 76404 706162 76586 706398
rect 76822 706162 77004 706398
rect 65604 679018 65786 679254
rect 66022 679018 66204 679254
rect 65604 678934 66204 679018
rect 65604 678698 65786 678934
rect 66022 678698 66204 678934
rect 65604 643254 66204 678698
rect 65604 643018 65786 643254
rect 66022 643018 66204 643254
rect 65604 642934 66204 643018
rect 65604 642698 65786 642934
rect 66022 642698 66204 642934
rect 65604 607254 66204 642698
rect 65604 607018 65786 607254
rect 66022 607018 66204 607254
rect 65604 606934 66204 607018
rect 65604 606698 65786 606934
rect 66022 606698 66204 606934
rect 65604 571254 66204 606698
rect 65604 571018 65786 571254
rect 66022 571018 66204 571254
rect 65604 570934 66204 571018
rect 65604 570698 65786 570934
rect 66022 570698 66204 570934
rect 65604 535254 66204 570698
rect 65604 535018 65786 535254
rect 66022 535018 66204 535254
rect 65604 534934 66204 535018
rect 65604 534698 65786 534934
rect 66022 534698 66204 534934
rect 65604 499254 66204 534698
rect 65604 499018 65786 499254
rect 66022 499018 66204 499254
rect 65604 498934 66204 499018
rect 65604 498698 65786 498934
rect 66022 498698 66204 498934
rect 65604 463254 66204 498698
rect 65604 463018 65786 463254
rect 66022 463018 66204 463254
rect 65604 462934 66204 463018
rect 65604 462698 65786 462934
rect 66022 462698 66204 462934
rect 65604 427254 66204 462698
rect 65604 427018 65786 427254
rect 66022 427018 66204 427254
rect 65604 426934 66204 427018
rect 65604 426698 65786 426934
rect 66022 426698 66204 426934
rect 65604 391254 66204 426698
rect 65604 391018 65786 391254
rect 66022 391018 66204 391254
rect 65604 390934 66204 391018
rect 65604 390698 65786 390934
rect 66022 390698 66204 390934
rect 65604 355254 66204 390698
rect 65604 355018 65786 355254
rect 66022 355018 66204 355254
rect 65604 354934 66204 355018
rect 65604 354698 65786 354934
rect 66022 354698 66204 354934
rect 65604 319254 66204 354698
rect 65604 319018 65786 319254
rect 66022 319018 66204 319254
rect 65604 318934 66204 319018
rect 65604 318698 65786 318934
rect 66022 318698 66204 318934
rect 65604 283254 66204 318698
rect 65604 283018 65786 283254
rect 66022 283018 66204 283254
rect 65604 282934 66204 283018
rect 65604 282698 65786 282934
rect 66022 282698 66204 282934
rect 65604 247254 66204 282698
rect 65604 247018 65786 247254
rect 66022 247018 66204 247254
rect 65604 246934 66204 247018
rect 65604 246698 65786 246934
rect 66022 246698 66204 246934
rect 65604 211254 66204 246698
rect 65604 211018 65786 211254
rect 66022 211018 66204 211254
rect 65604 210934 66204 211018
rect 65604 210698 65786 210934
rect 66022 210698 66204 210934
rect 65604 175254 66204 210698
rect 65604 175018 65786 175254
rect 66022 175018 66204 175254
rect 65604 174934 66204 175018
rect 65604 174698 65786 174934
rect 66022 174698 66204 174934
rect 65604 139254 66204 174698
rect 65604 139018 65786 139254
rect 66022 139018 66204 139254
rect 65604 138934 66204 139018
rect 65604 138698 65786 138934
rect 66022 138698 66204 138934
rect 65604 103254 66204 138698
rect 65604 103018 65786 103254
rect 66022 103018 66204 103254
rect 65604 102934 66204 103018
rect 65604 102698 65786 102934
rect 66022 102698 66204 102934
rect 65604 67254 66204 102698
rect 72804 704838 73404 705800
rect 72804 704602 72986 704838
rect 73222 704602 73404 704838
rect 72804 704518 73404 704602
rect 72804 704282 72986 704518
rect 73222 704282 73404 704518
rect 72804 686454 73404 704282
rect 72804 686218 72986 686454
rect 73222 686218 73404 686454
rect 72804 686134 73404 686218
rect 72804 685898 72986 686134
rect 73222 685898 73404 686134
rect 72804 650454 73404 685898
rect 72804 650218 72986 650454
rect 73222 650218 73404 650454
rect 72804 650134 73404 650218
rect 72804 649898 72986 650134
rect 73222 649898 73404 650134
rect 72804 614454 73404 649898
rect 72804 614218 72986 614454
rect 73222 614218 73404 614454
rect 72804 614134 73404 614218
rect 72804 613898 72986 614134
rect 73222 613898 73404 614134
rect 72804 578454 73404 613898
rect 72804 578218 72986 578454
rect 73222 578218 73404 578454
rect 72804 578134 73404 578218
rect 72804 577898 72986 578134
rect 73222 577898 73404 578134
rect 72804 542454 73404 577898
rect 72804 542218 72986 542454
rect 73222 542218 73404 542454
rect 72804 542134 73404 542218
rect 72804 541898 72986 542134
rect 73222 541898 73404 542134
rect 72804 506454 73404 541898
rect 72804 506218 72986 506454
rect 73222 506218 73404 506454
rect 72804 506134 73404 506218
rect 72804 505898 72986 506134
rect 73222 505898 73404 506134
rect 72804 470454 73404 505898
rect 72804 470218 72986 470454
rect 73222 470218 73404 470454
rect 72804 470134 73404 470218
rect 72804 469898 72986 470134
rect 73222 469898 73404 470134
rect 72804 434454 73404 469898
rect 72804 434218 72986 434454
rect 73222 434218 73404 434454
rect 72804 434134 73404 434218
rect 72804 433898 72986 434134
rect 73222 433898 73404 434134
rect 72804 398454 73404 433898
rect 72804 398218 72986 398454
rect 73222 398218 73404 398454
rect 72804 398134 73404 398218
rect 72804 397898 72986 398134
rect 73222 397898 73404 398134
rect 72804 362454 73404 397898
rect 72804 362218 72986 362454
rect 73222 362218 73404 362454
rect 72804 362134 73404 362218
rect 72804 361898 72986 362134
rect 73222 361898 73404 362134
rect 72804 326454 73404 361898
rect 72804 326218 72986 326454
rect 73222 326218 73404 326454
rect 72804 326134 73404 326218
rect 72804 325898 72986 326134
rect 73222 325898 73404 326134
rect 72804 290454 73404 325898
rect 72804 290218 72986 290454
rect 73222 290218 73404 290454
rect 72804 290134 73404 290218
rect 72804 289898 72986 290134
rect 73222 289898 73404 290134
rect 72804 254454 73404 289898
rect 72804 254218 72986 254454
rect 73222 254218 73404 254454
rect 72804 254134 73404 254218
rect 72804 253898 72986 254134
rect 73222 253898 73404 254134
rect 72804 218454 73404 253898
rect 72804 218218 72986 218454
rect 73222 218218 73404 218454
rect 72804 218134 73404 218218
rect 72804 217898 72986 218134
rect 73222 217898 73404 218134
rect 72804 182454 73404 217898
rect 72804 182218 72986 182454
rect 73222 182218 73404 182454
rect 72804 182134 73404 182218
rect 72804 181898 72986 182134
rect 73222 181898 73404 182134
rect 72804 146454 73404 181898
rect 72804 146218 72986 146454
rect 73222 146218 73404 146454
rect 72804 146134 73404 146218
rect 72804 145898 72986 146134
rect 73222 145898 73404 146134
rect 72804 110454 73404 145898
rect 72804 110218 72986 110454
rect 73222 110218 73404 110454
rect 72804 110134 73404 110218
rect 72804 109898 72986 110134
rect 73222 109898 73404 110134
rect 67587 93940 67653 93941
rect 67587 93876 67588 93940
rect 67652 93876 67653 93940
rect 67587 93875 67653 93876
rect 67590 93669 67650 93875
rect 67587 93668 67653 93669
rect 67587 93604 67588 93668
rect 67652 93604 67653 93668
rect 67587 93603 67653 93604
rect 65604 67018 65786 67254
rect 66022 67018 66204 67254
rect 65604 66934 66204 67018
rect 65604 66698 65786 66934
rect 66022 66698 66204 66934
rect 65604 31254 66204 66698
rect 65604 31018 65786 31254
rect 66022 31018 66204 31254
rect 65604 30934 66204 31018
rect 65604 30698 65786 30934
rect 66022 30698 66204 30934
rect 47604 -6222 47786 -5986
rect 48022 -6222 48204 -5986
rect 47604 -6306 48204 -6222
rect 47604 -6542 47786 -6306
rect 48022 -6542 48204 -6306
rect 47604 -7504 48204 -6542
rect 65604 -6926 66204 30698
rect 72804 74454 73404 109898
rect 72804 74218 72986 74454
rect 73222 74218 73404 74454
rect 72804 74134 73404 74218
rect 72804 73898 72986 74134
rect 73222 73898 73404 74134
rect 72804 38454 73404 73898
rect 72804 38218 72986 38454
rect 73222 38218 73404 38454
rect 72804 38134 73404 38218
rect 72804 37898 72986 38134
rect 73222 37898 73404 38134
rect 72804 2454 73404 37898
rect 72804 2218 72986 2454
rect 73222 2218 73404 2454
rect 72804 2134 73404 2218
rect 72804 1898 72986 2134
rect 73222 1898 73404 2134
rect 72804 -346 73404 1898
rect 72804 -582 72986 -346
rect 73222 -582 73404 -346
rect 72804 -666 73404 -582
rect 72804 -902 72986 -666
rect 73222 -902 73404 -666
rect 72804 -1864 73404 -902
rect 76404 690054 77004 706162
rect 76404 689818 76586 690054
rect 76822 689818 77004 690054
rect 76404 689734 77004 689818
rect 76404 689498 76586 689734
rect 76822 689498 77004 689734
rect 76404 654054 77004 689498
rect 76404 653818 76586 654054
rect 76822 653818 77004 654054
rect 76404 653734 77004 653818
rect 76404 653498 76586 653734
rect 76822 653498 77004 653734
rect 76404 618054 77004 653498
rect 76404 617818 76586 618054
rect 76822 617818 77004 618054
rect 76404 617734 77004 617818
rect 76404 617498 76586 617734
rect 76822 617498 77004 617734
rect 76404 582054 77004 617498
rect 76404 581818 76586 582054
rect 76822 581818 77004 582054
rect 76404 581734 77004 581818
rect 76404 581498 76586 581734
rect 76822 581498 77004 581734
rect 76404 546054 77004 581498
rect 76404 545818 76586 546054
rect 76822 545818 77004 546054
rect 76404 545734 77004 545818
rect 76404 545498 76586 545734
rect 76822 545498 77004 545734
rect 76404 510054 77004 545498
rect 76404 509818 76586 510054
rect 76822 509818 77004 510054
rect 76404 509734 77004 509818
rect 76404 509498 76586 509734
rect 76822 509498 77004 509734
rect 76404 474054 77004 509498
rect 76404 473818 76586 474054
rect 76822 473818 77004 474054
rect 76404 473734 77004 473818
rect 76404 473498 76586 473734
rect 76822 473498 77004 473734
rect 76404 438054 77004 473498
rect 76404 437818 76586 438054
rect 76822 437818 77004 438054
rect 76404 437734 77004 437818
rect 76404 437498 76586 437734
rect 76822 437498 77004 437734
rect 76404 402054 77004 437498
rect 76404 401818 76586 402054
rect 76822 401818 77004 402054
rect 76404 401734 77004 401818
rect 76404 401498 76586 401734
rect 76822 401498 77004 401734
rect 76404 366054 77004 401498
rect 76404 365818 76586 366054
rect 76822 365818 77004 366054
rect 76404 365734 77004 365818
rect 76404 365498 76586 365734
rect 76822 365498 77004 365734
rect 76404 330054 77004 365498
rect 76404 329818 76586 330054
rect 76822 329818 77004 330054
rect 76404 329734 77004 329818
rect 76404 329498 76586 329734
rect 76822 329498 77004 329734
rect 76404 294054 77004 329498
rect 76404 293818 76586 294054
rect 76822 293818 77004 294054
rect 76404 293734 77004 293818
rect 76404 293498 76586 293734
rect 76822 293498 77004 293734
rect 76404 258054 77004 293498
rect 76404 257818 76586 258054
rect 76822 257818 77004 258054
rect 76404 257734 77004 257818
rect 76404 257498 76586 257734
rect 76822 257498 77004 257734
rect 76404 222054 77004 257498
rect 76404 221818 76586 222054
rect 76822 221818 77004 222054
rect 76404 221734 77004 221818
rect 76404 221498 76586 221734
rect 76822 221498 77004 221734
rect 76404 186054 77004 221498
rect 76404 185818 76586 186054
rect 76822 185818 77004 186054
rect 76404 185734 77004 185818
rect 76404 185498 76586 185734
rect 76822 185498 77004 185734
rect 76404 150054 77004 185498
rect 76404 149818 76586 150054
rect 76822 149818 77004 150054
rect 76404 149734 77004 149818
rect 76404 149498 76586 149734
rect 76822 149498 77004 149734
rect 76404 114054 77004 149498
rect 76404 113818 76586 114054
rect 76822 113818 77004 114054
rect 76404 113734 77004 113818
rect 76404 113498 76586 113734
rect 76822 113498 77004 113734
rect 76404 78054 77004 113498
rect 76404 77818 76586 78054
rect 76822 77818 77004 78054
rect 76404 77734 77004 77818
rect 76404 77498 76586 77734
rect 76822 77498 77004 77734
rect 76404 42054 77004 77498
rect 76404 41818 76586 42054
rect 76822 41818 77004 42054
rect 76404 41734 77004 41818
rect 76404 41498 76586 41734
rect 76822 41498 77004 41734
rect 76404 6054 77004 41498
rect 76404 5818 76586 6054
rect 76822 5818 77004 6054
rect 76404 5734 77004 5818
rect 76404 5498 76586 5734
rect 76822 5498 77004 5734
rect 76404 -2226 77004 5498
rect 76404 -2462 76586 -2226
rect 76822 -2462 77004 -2226
rect 76404 -2546 77004 -2462
rect 76404 -2782 76586 -2546
rect 76822 -2782 77004 -2546
rect 76404 -3744 77004 -2782
rect 80004 693654 80604 708042
rect 80004 693418 80186 693654
rect 80422 693418 80604 693654
rect 80004 693334 80604 693418
rect 80004 693098 80186 693334
rect 80422 693098 80604 693334
rect 80004 657654 80604 693098
rect 80004 657418 80186 657654
rect 80422 657418 80604 657654
rect 80004 657334 80604 657418
rect 80004 657098 80186 657334
rect 80422 657098 80604 657334
rect 80004 621654 80604 657098
rect 80004 621418 80186 621654
rect 80422 621418 80604 621654
rect 80004 621334 80604 621418
rect 80004 621098 80186 621334
rect 80422 621098 80604 621334
rect 80004 585654 80604 621098
rect 80004 585418 80186 585654
rect 80422 585418 80604 585654
rect 80004 585334 80604 585418
rect 80004 585098 80186 585334
rect 80422 585098 80604 585334
rect 80004 549654 80604 585098
rect 80004 549418 80186 549654
rect 80422 549418 80604 549654
rect 80004 549334 80604 549418
rect 80004 549098 80186 549334
rect 80422 549098 80604 549334
rect 80004 513654 80604 549098
rect 80004 513418 80186 513654
rect 80422 513418 80604 513654
rect 80004 513334 80604 513418
rect 80004 513098 80186 513334
rect 80422 513098 80604 513334
rect 80004 477654 80604 513098
rect 80004 477418 80186 477654
rect 80422 477418 80604 477654
rect 80004 477334 80604 477418
rect 80004 477098 80186 477334
rect 80422 477098 80604 477334
rect 80004 441654 80604 477098
rect 80004 441418 80186 441654
rect 80422 441418 80604 441654
rect 80004 441334 80604 441418
rect 80004 441098 80186 441334
rect 80422 441098 80604 441334
rect 80004 405654 80604 441098
rect 80004 405418 80186 405654
rect 80422 405418 80604 405654
rect 80004 405334 80604 405418
rect 80004 405098 80186 405334
rect 80422 405098 80604 405334
rect 80004 369654 80604 405098
rect 80004 369418 80186 369654
rect 80422 369418 80604 369654
rect 80004 369334 80604 369418
rect 80004 369098 80186 369334
rect 80422 369098 80604 369334
rect 80004 333654 80604 369098
rect 80004 333418 80186 333654
rect 80422 333418 80604 333654
rect 80004 333334 80604 333418
rect 80004 333098 80186 333334
rect 80422 333098 80604 333334
rect 80004 297654 80604 333098
rect 80004 297418 80186 297654
rect 80422 297418 80604 297654
rect 80004 297334 80604 297418
rect 80004 297098 80186 297334
rect 80422 297098 80604 297334
rect 80004 261654 80604 297098
rect 80004 261418 80186 261654
rect 80422 261418 80604 261654
rect 80004 261334 80604 261418
rect 80004 261098 80186 261334
rect 80422 261098 80604 261334
rect 80004 225654 80604 261098
rect 80004 225418 80186 225654
rect 80422 225418 80604 225654
rect 80004 225334 80604 225418
rect 80004 225098 80186 225334
rect 80422 225098 80604 225334
rect 80004 189654 80604 225098
rect 80004 189418 80186 189654
rect 80422 189418 80604 189654
rect 80004 189334 80604 189418
rect 80004 189098 80186 189334
rect 80422 189098 80604 189334
rect 80004 153654 80604 189098
rect 80004 153418 80186 153654
rect 80422 153418 80604 153654
rect 80004 153334 80604 153418
rect 80004 153098 80186 153334
rect 80422 153098 80604 153334
rect 80004 117654 80604 153098
rect 80004 117418 80186 117654
rect 80422 117418 80604 117654
rect 80004 117334 80604 117418
rect 80004 117098 80186 117334
rect 80422 117098 80604 117334
rect 80004 81654 80604 117098
rect 80004 81418 80186 81654
rect 80422 81418 80604 81654
rect 80004 81334 80604 81418
rect 80004 81098 80186 81334
rect 80422 81098 80604 81334
rect 80004 45654 80604 81098
rect 80004 45418 80186 45654
rect 80422 45418 80604 45654
rect 80004 45334 80604 45418
rect 80004 45098 80186 45334
rect 80422 45098 80604 45334
rect 80004 9654 80604 45098
rect 80004 9418 80186 9654
rect 80422 9418 80604 9654
rect 80004 9334 80604 9418
rect 80004 9098 80186 9334
rect 80422 9098 80604 9334
rect 80004 -4106 80604 9098
rect 80004 -4342 80186 -4106
rect 80422 -4342 80604 -4106
rect 80004 -4426 80604 -4342
rect 80004 -4662 80186 -4426
rect 80422 -4662 80604 -4426
rect 80004 -5624 80604 -4662
rect 83604 697254 84204 709922
rect 101604 711418 102204 711440
rect 101604 711182 101786 711418
rect 102022 711182 102204 711418
rect 101604 711098 102204 711182
rect 101604 710862 101786 711098
rect 102022 710862 102204 711098
rect 98004 709538 98604 709560
rect 98004 709302 98186 709538
rect 98422 709302 98604 709538
rect 98004 709218 98604 709302
rect 98004 708982 98186 709218
rect 98422 708982 98604 709218
rect 94404 707658 95004 707680
rect 94404 707422 94586 707658
rect 94822 707422 95004 707658
rect 94404 707338 95004 707422
rect 94404 707102 94586 707338
rect 94822 707102 95004 707338
rect 83604 697018 83786 697254
rect 84022 697018 84204 697254
rect 83604 696934 84204 697018
rect 83604 696698 83786 696934
rect 84022 696698 84204 696934
rect 83604 661254 84204 696698
rect 83604 661018 83786 661254
rect 84022 661018 84204 661254
rect 83604 660934 84204 661018
rect 83604 660698 83786 660934
rect 84022 660698 84204 660934
rect 83604 625254 84204 660698
rect 83604 625018 83786 625254
rect 84022 625018 84204 625254
rect 83604 624934 84204 625018
rect 83604 624698 83786 624934
rect 84022 624698 84204 624934
rect 83604 589254 84204 624698
rect 83604 589018 83786 589254
rect 84022 589018 84204 589254
rect 83604 588934 84204 589018
rect 83604 588698 83786 588934
rect 84022 588698 84204 588934
rect 83604 553254 84204 588698
rect 83604 553018 83786 553254
rect 84022 553018 84204 553254
rect 83604 552934 84204 553018
rect 83604 552698 83786 552934
rect 84022 552698 84204 552934
rect 83604 517254 84204 552698
rect 83604 517018 83786 517254
rect 84022 517018 84204 517254
rect 83604 516934 84204 517018
rect 83604 516698 83786 516934
rect 84022 516698 84204 516934
rect 83604 481254 84204 516698
rect 83604 481018 83786 481254
rect 84022 481018 84204 481254
rect 83604 480934 84204 481018
rect 83604 480698 83786 480934
rect 84022 480698 84204 480934
rect 83604 445254 84204 480698
rect 83604 445018 83786 445254
rect 84022 445018 84204 445254
rect 83604 444934 84204 445018
rect 83604 444698 83786 444934
rect 84022 444698 84204 444934
rect 83604 409254 84204 444698
rect 83604 409018 83786 409254
rect 84022 409018 84204 409254
rect 83604 408934 84204 409018
rect 83604 408698 83786 408934
rect 84022 408698 84204 408934
rect 83604 373254 84204 408698
rect 83604 373018 83786 373254
rect 84022 373018 84204 373254
rect 83604 372934 84204 373018
rect 83604 372698 83786 372934
rect 84022 372698 84204 372934
rect 83604 337254 84204 372698
rect 83604 337018 83786 337254
rect 84022 337018 84204 337254
rect 83604 336934 84204 337018
rect 83604 336698 83786 336934
rect 84022 336698 84204 336934
rect 83604 301254 84204 336698
rect 83604 301018 83786 301254
rect 84022 301018 84204 301254
rect 83604 300934 84204 301018
rect 83604 300698 83786 300934
rect 84022 300698 84204 300934
rect 83604 265254 84204 300698
rect 83604 265018 83786 265254
rect 84022 265018 84204 265254
rect 83604 264934 84204 265018
rect 83604 264698 83786 264934
rect 84022 264698 84204 264934
rect 83604 229254 84204 264698
rect 83604 229018 83786 229254
rect 84022 229018 84204 229254
rect 83604 228934 84204 229018
rect 83604 228698 83786 228934
rect 84022 228698 84204 228934
rect 83604 193254 84204 228698
rect 83604 193018 83786 193254
rect 84022 193018 84204 193254
rect 83604 192934 84204 193018
rect 83604 192698 83786 192934
rect 84022 192698 84204 192934
rect 83604 157254 84204 192698
rect 83604 157018 83786 157254
rect 84022 157018 84204 157254
rect 83604 156934 84204 157018
rect 83604 156698 83786 156934
rect 84022 156698 84204 156934
rect 83604 121254 84204 156698
rect 83604 121018 83786 121254
rect 84022 121018 84204 121254
rect 83604 120934 84204 121018
rect 83604 120698 83786 120934
rect 84022 120698 84204 120934
rect 83604 85254 84204 120698
rect 90804 705778 91404 705800
rect 90804 705542 90986 705778
rect 91222 705542 91404 705778
rect 90804 705458 91404 705542
rect 90804 705222 90986 705458
rect 91222 705222 91404 705458
rect 90804 668454 91404 705222
rect 90804 668218 90986 668454
rect 91222 668218 91404 668454
rect 90804 668134 91404 668218
rect 90804 667898 90986 668134
rect 91222 667898 91404 668134
rect 90804 632454 91404 667898
rect 90804 632218 90986 632454
rect 91222 632218 91404 632454
rect 90804 632134 91404 632218
rect 90804 631898 90986 632134
rect 91222 631898 91404 632134
rect 90804 596454 91404 631898
rect 90804 596218 90986 596454
rect 91222 596218 91404 596454
rect 90804 596134 91404 596218
rect 90804 595898 90986 596134
rect 91222 595898 91404 596134
rect 90804 560454 91404 595898
rect 90804 560218 90986 560454
rect 91222 560218 91404 560454
rect 90804 560134 91404 560218
rect 90804 559898 90986 560134
rect 91222 559898 91404 560134
rect 90804 524454 91404 559898
rect 90804 524218 90986 524454
rect 91222 524218 91404 524454
rect 90804 524134 91404 524218
rect 90804 523898 90986 524134
rect 91222 523898 91404 524134
rect 90804 488454 91404 523898
rect 90804 488218 90986 488454
rect 91222 488218 91404 488454
rect 90804 488134 91404 488218
rect 90804 487898 90986 488134
rect 91222 487898 91404 488134
rect 90804 452454 91404 487898
rect 90804 452218 90986 452454
rect 91222 452218 91404 452454
rect 90804 452134 91404 452218
rect 90804 451898 90986 452134
rect 91222 451898 91404 452134
rect 90804 416454 91404 451898
rect 90804 416218 90986 416454
rect 91222 416218 91404 416454
rect 90804 416134 91404 416218
rect 90804 415898 90986 416134
rect 91222 415898 91404 416134
rect 90804 380454 91404 415898
rect 90804 380218 90986 380454
rect 91222 380218 91404 380454
rect 90804 380134 91404 380218
rect 90804 379898 90986 380134
rect 91222 379898 91404 380134
rect 90804 344454 91404 379898
rect 90804 344218 90986 344454
rect 91222 344218 91404 344454
rect 90804 344134 91404 344218
rect 90804 343898 90986 344134
rect 91222 343898 91404 344134
rect 90804 308454 91404 343898
rect 90804 308218 90986 308454
rect 91222 308218 91404 308454
rect 90804 308134 91404 308218
rect 90804 307898 90986 308134
rect 91222 307898 91404 308134
rect 90804 272454 91404 307898
rect 90804 272218 90986 272454
rect 91222 272218 91404 272454
rect 90804 272134 91404 272218
rect 90804 271898 90986 272134
rect 91222 271898 91404 272134
rect 90804 236454 91404 271898
rect 90804 236218 90986 236454
rect 91222 236218 91404 236454
rect 90804 236134 91404 236218
rect 90804 235898 90986 236134
rect 91222 235898 91404 236134
rect 90804 200454 91404 235898
rect 90804 200218 90986 200454
rect 91222 200218 91404 200454
rect 90804 200134 91404 200218
rect 90804 199898 90986 200134
rect 91222 199898 91404 200134
rect 90804 164454 91404 199898
rect 90804 164218 90986 164454
rect 91222 164218 91404 164454
rect 90804 164134 91404 164218
rect 90804 163898 90986 164134
rect 91222 163898 91404 164134
rect 90804 128454 91404 163898
rect 90804 128218 90986 128454
rect 91222 128218 91404 128454
rect 90804 128134 91404 128218
rect 90804 127898 90986 128134
rect 91222 127898 91404 128134
rect 86907 93940 86973 93941
rect 86907 93876 86908 93940
rect 86972 93876 86973 93940
rect 86907 93875 86973 93876
rect 86910 93669 86970 93875
rect 86907 93668 86973 93669
rect 86907 93604 86908 93668
rect 86972 93604 86973 93668
rect 86907 93603 86973 93604
rect 83604 85018 83786 85254
rect 84022 85018 84204 85254
rect 83604 84934 84204 85018
rect 83604 84698 83786 84934
rect 84022 84698 84204 84934
rect 83604 49254 84204 84698
rect 83604 49018 83786 49254
rect 84022 49018 84204 49254
rect 83604 48934 84204 49018
rect 83604 48698 83786 48934
rect 84022 48698 84204 48934
rect 83604 13254 84204 48698
rect 83604 13018 83786 13254
rect 84022 13018 84204 13254
rect 83604 12934 84204 13018
rect 83604 12698 83786 12934
rect 84022 12698 84204 12934
rect 65604 -7162 65786 -6926
rect 66022 -7162 66204 -6926
rect 65604 -7246 66204 -7162
rect 65604 -7482 65786 -7246
rect 66022 -7482 66204 -7246
rect 65604 -7504 66204 -7482
rect 83604 -5986 84204 12698
rect 90804 92454 91404 127898
rect 90804 92218 90986 92454
rect 91222 92218 91404 92454
rect 90804 92134 91404 92218
rect 90804 91898 90986 92134
rect 91222 91898 91404 92134
rect 90804 56454 91404 91898
rect 90804 56218 90986 56454
rect 91222 56218 91404 56454
rect 90804 56134 91404 56218
rect 90804 55898 90986 56134
rect 91222 55898 91404 56134
rect 90804 20454 91404 55898
rect 90804 20218 90986 20454
rect 91222 20218 91404 20454
rect 90804 20134 91404 20218
rect 90804 19898 90986 20134
rect 91222 19898 91404 20134
rect 90804 -1286 91404 19898
rect 90804 -1522 90986 -1286
rect 91222 -1522 91404 -1286
rect 90804 -1606 91404 -1522
rect 90804 -1842 90986 -1606
rect 91222 -1842 91404 -1606
rect 90804 -1864 91404 -1842
rect 94404 672054 95004 707102
rect 94404 671818 94586 672054
rect 94822 671818 95004 672054
rect 94404 671734 95004 671818
rect 94404 671498 94586 671734
rect 94822 671498 95004 671734
rect 94404 636054 95004 671498
rect 94404 635818 94586 636054
rect 94822 635818 95004 636054
rect 94404 635734 95004 635818
rect 94404 635498 94586 635734
rect 94822 635498 95004 635734
rect 94404 600054 95004 635498
rect 94404 599818 94586 600054
rect 94822 599818 95004 600054
rect 94404 599734 95004 599818
rect 94404 599498 94586 599734
rect 94822 599498 95004 599734
rect 94404 564054 95004 599498
rect 94404 563818 94586 564054
rect 94822 563818 95004 564054
rect 94404 563734 95004 563818
rect 94404 563498 94586 563734
rect 94822 563498 95004 563734
rect 94404 528054 95004 563498
rect 94404 527818 94586 528054
rect 94822 527818 95004 528054
rect 94404 527734 95004 527818
rect 94404 527498 94586 527734
rect 94822 527498 95004 527734
rect 94404 492054 95004 527498
rect 94404 491818 94586 492054
rect 94822 491818 95004 492054
rect 94404 491734 95004 491818
rect 94404 491498 94586 491734
rect 94822 491498 95004 491734
rect 94404 456054 95004 491498
rect 94404 455818 94586 456054
rect 94822 455818 95004 456054
rect 94404 455734 95004 455818
rect 94404 455498 94586 455734
rect 94822 455498 95004 455734
rect 94404 420054 95004 455498
rect 94404 419818 94586 420054
rect 94822 419818 95004 420054
rect 94404 419734 95004 419818
rect 94404 419498 94586 419734
rect 94822 419498 95004 419734
rect 94404 384054 95004 419498
rect 94404 383818 94586 384054
rect 94822 383818 95004 384054
rect 94404 383734 95004 383818
rect 94404 383498 94586 383734
rect 94822 383498 95004 383734
rect 94404 348054 95004 383498
rect 94404 347818 94586 348054
rect 94822 347818 95004 348054
rect 94404 347734 95004 347818
rect 94404 347498 94586 347734
rect 94822 347498 95004 347734
rect 94404 312054 95004 347498
rect 94404 311818 94586 312054
rect 94822 311818 95004 312054
rect 94404 311734 95004 311818
rect 94404 311498 94586 311734
rect 94822 311498 95004 311734
rect 94404 276054 95004 311498
rect 94404 275818 94586 276054
rect 94822 275818 95004 276054
rect 94404 275734 95004 275818
rect 94404 275498 94586 275734
rect 94822 275498 95004 275734
rect 94404 240054 95004 275498
rect 94404 239818 94586 240054
rect 94822 239818 95004 240054
rect 94404 239734 95004 239818
rect 94404 239498 94586 239734
rect 94822 239498 95004 239734
rect 94404 204054 95004 239498
rect 94404 203818 94586 204054
rect 94822 203818 95004 204054
rect 94404 203734 95004 203818
rect 94404 203498 94586 203734
rect 94822 203498 95004 203734
rect 94404 168054 95004 203498
rect 94404 167818 94586 168054
rect 94822 167818 95004 168054
rect 94404 167734 95004 167818
rect 94404 167498 94586 167734
rect 94822 167498 95004 167734
rect 94404 132054 95004 167498
rect 94404 131818 94586 132054
rect 94822 131818 95004 132054
rect 94404 131734 95004 131818
rect 94404 131498 94586 131734
rect 94822 131498 95004 131734
rect 94404 96054 95004 131498
rect 94404 95818 94586 96054
rect 94822 95818 95004 96054
rect 94404 95734 95004 95818
rect 94404 95498 94586 95734
rect 94822 95498 95004 95734
rect 94404 60054 95004 95498
rect 94404 59818 94586 60054
rect 94822 59818 95004 60054
rect 94404 59734 95004 59818
rect 94404 59498 94586 59734
rect 94822 59498 95004 59734
rect 94404 24054 95004 59498
rect 94404 23818 94586 24054
rect 94822 23818 95004 24054
rect 94404 23734 95004 23818
rect 94404 23498 94586 23734
rect 94822 23498 95004 23734
rect 94404 -3166 95004 23498
rect 94404 -3402 94586 -3166
rect 94822 -3402 95004 -3166
rect 94404 -3486 95004 -3402
rect 94404 -3722 94586 -3486
rect 94822 -3722 95004 -3486
rect 94404 -3744 95004 -3722
rect 98004 675654 98604 708982
rect 98004 675418 98186 675654
rect 98422 675418 98604 675654
rect 98004 675334 98604 675418
rect 98004 675098 98186 675334
rect 98422 675098 98604 675334
rect 98004 639654 98604 675098
rect 98004 639418 98186 639654
rect 98422 639418 98604 639654
rect 98004 639334 98604 639418
rect 98004 639098 98186 639334
rect 98422 639098 98604 639334
rect 98004 603654 98604 639098
rect 98004 603418 98186 603654
rect 98422 603418 98604 603654
rect 98004 603334 98604 603418
rect 98004 603098 98186 603334
rect 98422 603098 98604 603334
rect 98004 567654 98604 603098
rect 98004 567418 98186 567654
rect 98422 567418 98604 567654
rect 98004 567334 98604 567418
rect 98004 567098 98186 567334
rect 98422 567098 98604 567334
rect 98004 531654 98604 567098
rect 98004 531418 98186 531654
rect 98422 531418 98604 531654
rect 98004 531334 98604 531418
rect 98004 531098 98186 531334
rect 98422 531098 98604 531334
rect 98004 495654 98604 531098
rect 98004 495418 98186 495654
rect 98422 495418 98604 495654
rect 98004 495334 98604 495418
rect 98004 495098 98186 495334
rect 98422 495098 98604 495334
rect 98004 459654 98604 495098
rect 98004 459418 98186 459654
rect 98422 459418 98604 459654
rect 98004 459334 98604 459418
rect 98004 459098 98186 459334
rect 98422 459098 98604 459334
rect 98004 423654 98604 459098
rect 98004 423418 98186 423654
rect 98422 423418 98604 423654
rect 98004 423334 98604 423418
rect 98004 423098 98186 423334
rect 98422 423098 98604 423334
rect 98004 387654 98604 423098
rect 98004 387418 98186 387654
rect 98422 387418 98604 387654
rect 98004 387334 98604 387418
rect 98004 387098 98186 387334
rect 98422 387098 98604 387334
rect 98004 351654 98604 387098
rect 98004 351418 98186 351654
rect 98422 351418 98604 351654
rect 98004 351334 98604 351418
rect 98004 351098 98186 351334
rect 98422 351098 98604 351334
rect 98004 315654 98604 351098
rect 98004 315418 98186 315654
rect 98422 315418 98604 315654
rect 98004 315334 98604 315418
rect 98004 315098 98186 315334
rect 98422 315098 98604 315334
rect 98004 279654 98604 315098
rect 98004 279418 98186 279654
rect 98422 279418 98604 279654
rect 98004 279334 98604 279418
rect 98004 279098 98186 279334
rect 98422 279098 98604 279334
rect 98004 243654 98604 279098
rect 98004 243418 98186 243654
rect 98422 243418 98604 243654
rect 98004 243334 98604 243418
rect 98004 243098 98186 243334
rect 98422 243098 98604 243334
rect 98004 207654 98604 243098
rect 98004 207418 98186 207654
rect 98422 207418 98604 207654
rect 98004 207334 98604 207418
rect 98004 207098 98186 207334
rect 98422 207098 98604 207334
rect 98004 171654 98604 207098
rect 98004 171418 98186 171654
rect 98422 171418 98604 171654
rect 98004 171334 98604 171418
rect 98004 171098 98186 171334
rect 98422 171098 98604 171334
rect 98004 135654 98604 171098
rect 98004 135418 98186 135654
rect 98422 135418 98604 135654
rect 98004 135334 98604 135418
rect 98004 135098 98186 135334
rect 98422 135098 98604 135334
rect 98004 99654 98604 135098
rect 98004 99418 98186 99654
rect 98422 99418 98604 99654
rect 98004 99334 98604 99418
rect 98004 99098 98186 99334
rect 98422 99098 98604 99334
rect 98004 63654 98604 99098
rect 98004 63418 98186 63654
rect 98422 63418 98604 63654
rect 98004 63334 98604 63418
rect 98004 63098 98186 63334
rect 98422 63098 98604 63334
rect 98004 27654 98604 63098
rect 98004 27418 98186 27654
rect 98422 27418 98604 27654
rect 98004 27334 98604 27418
rect 98004 27098 98186 27334
rect 98422 27098 98604 27334
rect 98004 -5046 98604 27098
rect 98004 -5282 98186 -5046
rect 98422 -5282 98604 -5046
rect 98004 -5366 98604 -5282
rect 98004 -5602 98186 -5366
rect 98422 -5602 98604 -5366
rect 98004 -5624 98604 -5602
rect 101604 679254 102204 710862
rect 119604 710478 120204 711440
rect 119604 710242 119786 710478
rect 120022 710242 120204 710478
rect 119604 710158 120204 710242
rect 119604 709922 119786 710158
rect 120022 709922 120204 710158
rect 116004 708598 116604 709560
rect 116004 708362 116186 708598
rect 116422 708362 116604 708598
rect 116004 708278 116604 708362
rect 116004 708042 116186 708278
rect 116422 708042 116604 708278
rect 112404 706718 113004 707680
rect 112404 706482 112586 706718
rect 112822 706482 113004 706718
rect 112404 706398 113004 706482
rect 112404 706162 112586 706398
rect 112822 706162 113004 706398
rect 101604 679018 101786 679254
rect 102022 679018 102204 679254
rect 101604 678934 102204 679018
rect 101604 678698 101786 678934
rect 102022 678698 102204 678934
rect 101604 643254 102204 678698
rect 101604 643018 101786 643254
rect 102022 643018 102204 643254
rect 101604 642934 102204 643018
rect 101604 642698 101786 642934
rect 102022 642698 102204 642934
rect 101604 607254 102204 642698
rect 101604 607018 101786 607254
rect 102022 607018 102204 607254
rect 101604 606934 102204 607018
rect 101604 606698 101786 606934
rect 102022 606698 102204 606934
rect 101604 571254 102204 606698
rect 101604 571018 101786 571254
rect 102022 571018 102204 571254
rect 101604 570934 102204 571018
rect 101604 570698 101786 570934
rect 102022 570698 102204 570934
rect 101604 535254 102204 570698
rect 101604 535018 101786 535254
rect 102022 535018 102204 535254
rect 101604 534934 102204 535018
rect 101604 534698 101786 534934
rect 102022 534698 102204 534934
rect 101604 499254 102204 534698
rect 101604 499018 101786 499254
rect 102022 499018 102204 499254
rect 101604 498934 102204 499018
rect 101604 498698 101786 498934
rect 102022 498698 102204 498934
rect 101604 463254 102204 498698
rect 101604 463018 101786 463254
rect 102022 463018 102204 463254
rect 101604 462934 102204 463018
rect 101604 462698 101786 462934
rect 102022 462698 102204 462934
rect 101604 427254 102204 462698
rect 101604 427018 101786 427254
rect 102022 427018 102204 427254
rect 101604 426934 102204 427018
rect 101604 426698 101786 426934
rect 102022 426698 102204 426934
rect 101604 391254 102204 426698
rect 101604 391018 101786 391254
rect 102022 391018 102204 391254
rect 101604 390934 102204 391018
rect 101604 390698 101786 390934
rect 102022 390698 102204 390934
rect 101604 355254 102204 390698
rect 101604 355018 101786 355254
rect 102022 355018 102204 355254
rect 101604 354934 102204 355018
rect 101604 354698 101786 354934
rect 102022 354698 102204 354934
rect 101604 319254 102204 354698
rect 101604 319018 101786 319254
rect 102022 319018 102204 319254
rect 101604 318934 102204 319018
rect 101604 318698 101786 318934
rect 102022 318698 102204 318934
rect 101604 283254 102204 318698
rect 101604 283018 101786 283254
rect 102022 283018 102204 283254
rect 101604 282934 102204 283018
rect 101604 282698 101786 282934
rect 102022 282698 102204 282934
rect 101604 247254 102204 282698
rect 101604 247018 101786 247254
rect 102022 247018 102204 247254
rect 101604 246934 102204 247018
rect 101604 246698 101786 246934
rect 102022 246698 102204 246934
rect 101604 211254 102204 246698
rect 101604 211018 101786 211254
rect 102022 211018 102204 211254
rect 101604 210934 102204 211018
rect 101604 210698 101786 210934
rect 102022 210698 102204 210934
rect 101604 175254 102204 210698
rect 101604 175018 101786 175254
rect 102022 175018 102204 175254
rect 101604 174934 102204 175018
rect 101604 174698 101786 174934
rect 102022 174698 102204 174934
rect 101604 139254 102204 174698
rect 101604 139018 101786 139254
rect 102022 139018 102204 139254
rect 101604 138934 102204 139018
rect 101604 138698 101786 138934
rect 102022 138698 102204 138934
rect 101604 103254 102204 138698
rect 101604 103018 101786 103254
rect 102022 103018 102204 103254
rect 101604 102934 102204 103018
rect 101604 102698 101786 102934
rect 102022 102698 102204 102934
rect 101604 67254 102204 102698
rect 108804 704838 109404 705800
rect 108804 704602 108986 704838
rect 109222 704602 109404 704838
rect 108804 704518 109404 704602
rect 108804 704282 108986 704518
rect 109222 704282 109404 704518
rect 108804 686454 109404 704282
rect 108804 686218 108986 686454
rect 109222 686218 109404 686454
rect 108804 686134 109404 686218
rect 108804 685898 108986 686134
rect 109222 685898 109404 686134
rect 108804 650454 109404 685898
rect 108804 650218 108986 650454
rect 109222 650218 109404 650454
rect 108804 650134 109404 650218
rect 108804 649898 108986 650134
rect 109222 649898 109404 650134
rect 108804 614454 109404 649898
rect 108804 614218 108986 614454
rect 109222 614218 109404 614454
rect 108804 614134 109404 614218
rect 108804 613898 108986 614134
rect 109222 613898 109404 614134
rect 108804 578454 109404 613898
rect 108804 578218 108986 578454
rect 109222 578218 109404 578454
rect 108804 578134 109404 578218
rect 108804 577898 108986 578134
rect 109222 577898 109404 578134
rect 108804 542454 109404 577898
rect 108804 542218 108986 542454
rect 109222 542218 109404 542454
rect 108804 542134 109404 542218
rect 108804 541898 108986 542134
rect 109222 541898 109404 542134
rect 108804 506454 109404 541898
rect 108804 506218 108986 506454
rect 109222 506218 109404 506454
rect 108804 506134 109404 506218
rect 108804 505898 108986 506134
rect 109222 505898 109404 506134
rect 108804 470454 109404 505898
rect 108804 470218 108986 470454
rect 109222 470218 109404 470454
rect 108804 470134 109404 470218
rect 108804 469898 108986 470134
rect 109222 469898 109404 470134
rect 108804 434454 109404 469898
rect 108804 434218 108986 434454
rect 109222 434218 109404 434454
rect 108804 434134 109404 434218
rect 108804 433898 108986 434134
rect 109222 433898 109404 434134
rect 108804 398454 109404 433898
rect 108804 398218 108986 398454
rect 109222 398218 109404 398454
rect 108804 398134 109404 398218
rect 108804 397898 108986 398134
rect 109222 397898 109404 398134
rect 108804 362454 109404 397898
rect 108804 362218 108986 362454
rect 109222 362218 109404 362454
rect 108804 362134 109404 362218
rect 108804 361898 108986 362134
rect 109222 361898 109404 362134
rect 108804 326454 109404 361898
rect 108804 326218 108986 326454
rect 109222 326218 109404 326454
rect 108804 326134 109404 326218
rect 108804 325898 108986 326134
rect 109222 325898 109404 326134
rect 108804 290454 109404 325898
rect 108804 290218 108986 290454
rect 109222 290218 109404 290454
rect 108804 290134 109404 290218
rect 108804 289898 108986 290134
rect 109222 289898 109404 290134
rect 108804 254454 109404 289898
rect 108804 254218 108986 254454
rect 109222 254218 109404 254454
rect 108804 254134 109404 254218
rect 108804 253898 108986 254134
rect 109222 253898 109404 254134
rect 108804 218454 109404 253898
rect 108804 218218 108986 218454
rect 109222 218218 109404 218454
rect 108804 218134 109404 218218
rect 108804 217898 108986 218134
rect 109222 217898 109404 218134
rect 108804 182454 109404 217898
rect 108804 182218 108986 182454
rect 109222 182218 109404 182454
rect 108804 182134 109404 182218
rect 108804 181898 108986 182134
rect 109222 181898 109404 182134
rect 108804 146454 109404 181898
rect 108804 146218 108986 146454
rect 109222 146218 109404 146454
rect 108804 146134 109404 146218
rect 108804 145898 108986 146134
rect 109222 145898 109404 146134
rect 108804 110454 109404 145898
rect 108804 110218 108986 110454
rect 109222 110218 109404 110454
rect 108804 110134 109404 110218
rect 108804 109898 108986 110134
rect 109222 109898 109404 110134
rect 106227 93940 106293 93941
rect 106227 93876 106228 93940
rect 106292 93876 106293 93940
rect 106227 93875 106293 93876
rect 106230 93669 106290 93875
rect 106227 93668 106293 93669
rect 106227 93604 106228 93668
rect 106292 93604 106293 93668
rect 106227 93603 106293 93604
rect 101604 67018 101786 67254
rect 102022 67018 102204 67254
rect 101604 66934 102204 67018
rect 101604 66698 101786 66934
rect 102022 66698 102204 66934
rect 101604 31254 102204 66698
rect 101604 31018 101786 31254
rect 102022 31018 102204 31254
rect 101604 30934 102204 31018
rect 101604 30698 101786 30934
rect 102022 30698 102204 30934
rect 83604 -6222 83786 -5986
rect 84022 -6222 84204 -5986
rect 83604 -6306 84204 -6222
rect 83604 -6542 83786 -6306
rect 84022 -6542 84204 -6306
rect 83604 -7504 84204 -6542
rect 101604 -6926 102204 30698
rect 108804 74454 109404 109898
rect 108804 74218 108986 74454
rect 109222 74218 109404 74454
rect 108804 74134 109404 74218
rect 108804 73898 108986 74134
rect 109222 73898 109404 74134
rect 108804 38454 109404 73898
rect 108804 38218 108986 38454
rect 109222 38218 109404 38454
rect 108804 38134 109404 38218
rect 108804 37898 108986 38134
rect 109222 37898 109404 38134
rect 108804 2454 109404 37898
rect 108804 2218 108986 2454
rect 109222 2218 109404 2454
rect 108804 2134 109404 2218
rect 108804 1898 108986 2134
rect 109222 1898 109404 2134
rect 108804 -346 109404 1898
rect 108804 -582 108986 -346
rect 109222 -582 109404 -346
rect 108804 -666 109404 -582
rect 108804 -902 108986 -666
rect 109222 -902 109404 -666
rect 108804 -1864 109404 -902
rect 112404 690054 113004 706162
rect 112404 689818 112586 690054
rect 112822 689818 113004 690054
rect 112404 689734 113004 689818
rect 112404 689498 112586 689734
rect 112822 689498 113004 689734
rect 112404 654054 113004 689498
rect 112404 653818 112586 654054
rect 112822 653818 113004 654054
rect 112404 653734 113004 653818
rect 112404 653498 112586 653734
rect 112822 653498 113004 653734
rect 112404 618054 113004 653498
rect 112404 617818 112586 618054
rect 112822 617818 113004 618054
rect 112404 617734 113004 617818
rect 112404 617498 112586 617734
rect 112822 617498 113004 617734
rect 112404 582054 113004 617498
rect 112404 581818 112586 582054
rect 112822 581818 113004 582054
rect 112404 581734 113004 581818
rect 112404 581498 112586 581734
rect 112822 581498 113004 581734
rect 112404 546054 113004 581498
rect 112404 545818 112586 546054
rect 112822 545818 113004 546054
rect 112404 545734 113004 545818
rect 112404 545498 112586 545734
rect 112822 545498 113004 545734
rect 112404 510054 113004 545498
rect 112404 509818 112586 510054
rect 112822 509818 113004 510054
rect 112404 509734 113004 509818
rect 112404 509498 112586 509734
rect 112822 509498 113004 509734
rect 112404 474054 113004 509498
rect 112404 473818 112586 474054
rect 112822 473818 113004 474054
rect 112404 473734 113004 473818
rect 112404 473498 112586 473734
rect 112822 473498 113004 473734
rect 112404 438054 113004 473498
rect 112404 437818 112586 438054
rect 112822 437818 113004 438054
rect 112404 437734 113004 437818
rect 112404 437498 112586 437734
rect 112822 437498 113004 437734
rect 112404 402054 113004 437498
rect 112404 401818 112586 402054
rect 112822 401818 113004 402054
rect 112404 401734 113004 401818
rect 112404 401498 112586 401734
rect 112822 401498 113004 401734
rect 112404 366054 113004 401498
rect 112404 365818 112586 366054
rect 112822 365818 113004 366054
rect 112404 365734 113004 365818
rect 112404 365498 112586 365734
rect 112822 365498 113004 365734
rect 112404 330054 113004 365498
rect 112404 329818 112586 330054
rect 112822 329818 113004 330054
rect 112404 329734 113004 329818
rect 112404 329498 112586 329734
rect 112822 329498 113004 329734
rect 112404 294054 113004 329498
rect 112404 293818 112586 294054
rect 112822 293818 113004 294054
rect 112404 293734 113004 293818
rect 112404 293498 112586 293734
rect 112822 293498 113004 293734
rect 112404 258054 113004 293498
rect 112404 257818 112586 258054
rect 112822 257818 113004 258054
rect 112404 257734 113004 257818
rect 112404 257498 112586 257734
rect 112822 257498 113004 257734
rect 112404 222054 113004 257498
rect 112404 221818 112586 222054
rect 112822 221818 113004 222054
rect 112404 221734 113004 221818
rect 112404 221498 112586 221734
rect 112822 221498 113004 221734
rect 112404 186054 113004 221498
rect 112404 185818 112586 186054
rect 112822 185818 113004 186054
rect 112404 185734 113004 185818
rect 112404 185498 112586 185734
rect 112822 185498 113004 185734
rect 112404 150054 113004 185498
rect 112404 149818 112586 150054
rect 112822 149818 113004 150054
rect 112404 149734 113004 149818
rect 112404 149498 112586 149734
rect 112822 149498 113004 149734
rect 112404 114054 113004 149498
rect 112404 113818 112586 114054
rect 112822 113818 113004 114054
rect 112404 113734 113004 113818
rect 112404 113498 112586 113734
rect 112822 113498 113004 113734
rect 112404 78054 113004 113498
rect 112404 77818 112586 78054
rect 112822 77818 113004 78054
rect 112404 77734 113004 77818
rect 112404 77498 112586 77734
rect 112822 77498 113004 77734
rect 112404 42054 113004 77498
rect 112404 41818 112586 42054
rect 112822 41818 113004 42054
rect 112404 41734 113004 41818
rect 112404 41498 112586 41734
rect 112822 41498 113004 41734
rect 112404 6054 113004 41498
rect 112404 5818 112586 6054
rect 112822 5818 113004 6054
rect 112404 5734 113004 5818
rect 112404 5498 112586 5734
rect 112822 5498 113004 5734
rect 112404 -2226 113004 5498
rect 112404 -2462 112586 -2226
rect 112822 -2462 113004 -2226
rect 112404 -2546 113004 -2462
rect 112404 -2782 112586 -2546
rect 112822 -2782 113004 -2546
rect 112404 -3744 113004 -2782
rect 116004 693654 116604 708042
rect 116004 693418 116186 693654
rect 116422 693418 116604 693654
rect 116004 693334 116604 693418
rect 116004 693098 116186 693334
rect 116422 693098 116604 693334
rect 116004 657654 116604 693098
rect 116004 657418 116186 657654
rect 116422 657418 116604 657654
rect 116004 657334 116604 657418
rect 116004 657098 116186 657334
rect 116422 657098 116604 657334
rect 116004 621654 116604 657098
rect 116004 621418 116186 621654
rect 116422 621418 116604 621654
rect 116004 621334 116604 621418
rect 116004 621098 116186 621334
rect 116422 621098 116604 621334
rect 116004 585654 116604 621098
rect 116004 585418 116186 585654
rect 116422 585418 116604 585654
rect 116004 585334 116604 585418
rect 116004 585098 116186 585334
rect 116422 585098 116604 585334
rect 116004 549654 116604 585098
rect 116004 549418 116186 549654
rect 116422 549418 116604 549654
rect 116004 549334 116604 549418
rect 116004 549098 116186 549334
rect 116422 549098 116604 549334
rect 116004 513654 116604 549098
rect 116004 513418 116186 513654
rect 116422 513418 116604 513654
rect 116004 513334 116604 513418
rect 116004 513098 116186 513334
rect 116422 513098 116604 513334
rect 116004 477654 116604 513098
rect 116004 477418 116186 477654
rect 116422 477418 116604 477654
rect 116004 477334 116604 477418
rect 116004 477098 116186 477334
rect 116422 477098 116604 477334
rect 116004 441654 116604 477098
rect 116004 441418 116186 441654
rect 116422 441418 116604 441654
rect 116004 441334 116604 441418
rect 116004 441098 116186 441334
rect 116422 441098 116604 441334
rect 116004 405654 116604 441098
rect 116004 405418 116186 405654
rect 116422 405418 116604 405654
rect 116004 405334 116604 405418
rect 116004 405098 116186 405334
rect 116422 405098 116604 405334
rect 116004 369654 116604 405098
rect 116004 369418 116186 369654
rect 116422 369418 116604 369654
rect 116004 369334 116604 369418
rect 116004 369098 116186 369334
rect 116422 369098 116604 369334
rect 116004 333654 116604 369098
rect 116004 333418 116186 333654
rect 116422 333418 116604 333654
rect 116004 333334 116604 333418
rect 116004 333098 116186 333334
rect 116422 333098 116604 333334
rect 116004 297654 116604 333098
rect 116004 297418 116186 297654
rect 116422 297418 116604 297654
rect 116004 297334 116604 297418
rect 116004 297098 116186 297334
rect 116422 297098 116604 297334
rect 116004 261654 116604 297098
rect 116004 261418 116186 261654
rect 116422 261418 116604 261654
rect 116004 261334 116604 261418
rect 116004 261098 116186 261334
rect 116422 261098 116604 261334
rect 116004 225654 116604 261098
rect 116004 225418 116186 225654
rect 116422 225418 116604 225654
rect 116004 225334 116604 225418
rect 116004 225098 116186 225334
rect 116422 225098 116604 225334
rect 116004 189654 116604 225098
rect 116004 189418 116186 189654
rect 116422 189418 116604 189654
rect 116004 189334 116604 189418
rect 116004 189098 116186 189334
rect 116422 189098 116604 189334
rect 116004 153654 116604 189098
rect 116004 153418 116186 153654
rect 116422 153418 116604 153654
rect 116004 153334 116604 153418
rect 116004 153098 116186 153334
rect 116422 153098 116604 153334
rect 116004 117654 116604 153098
rect 116004 117418 116186 117654
rect 116422 117418 116604 117654
rect 116004 117334 116604 117418
rect 116004 117098 116186 117334
rect 116422 117098 116604 117334
rect 116004 81654 116604 117098
rect 116004 81418 116186 81654
rect 116422 81418 116604 81654
rect 116004 81334 116604 81418
rect 116004 81098 116186 81334
rect 116422 81098 116604 81334
rect 116004 45654 116604 81098
rect 116004 45418 116186 45654
rect 116422 45418 116604 45654
rect 116004 45334 116604 45418
rect 116004 45098 116186 45334
rect 116422 45098 116604 45334
rect 116004 9654 116604 45098
rect 116004 9418 116186 9654
rect 116422 9418 116604 9654
rect 116004 9334 116604 9418
rect 116004 9098 116186 9334
rect 116422 9098 116604 9334
rect 116004 -4106 116604 9098
rect 116004 -4342 116186 -4106
rect 116422 -4342 116604 -4106
rect 116004 -4426 116604 -4342
rect 116004 -4662 116186 -4426
rect 116422 -4662 116604 -4426
rect 116004 -5624 116604 -4662
rect 119604 697254 120204 709922
rect 137604 711418 138204 711440
rect 137604 711182 137786 711418
rect 138022 711182 138204 711418
rect 137604 711098 138204 711182
rect 137604 710862 137786 711098
rect 138022 710862 138204 711098
rect 134004 709538 134604 709560
rect 134004 709302 134186 709538
rect 134422 709302 134604 709538
rect 134004 709218 134604 709302
rect 134004 708982 134186 709218
rect 134422 708982 134604 709218
rect 130404 707658 131004 707680
rect 130404 707422 130586 707658
rect 130822 707422 131004 707658
rect 130404 707338 131004 707422
rect 130404 707102 130586 707338
rect 130822 707102 131004 707338
rect 119604 697018 119786 697254
rect 120022 697018 120204 697254
rect 119604 696934 120204 697018
rect 119604 696698 119786 696934
rect 120022 696698 120204 696934
rect 119604 661254 120204 696698
rect 119604 661018 119786 661254
rect 120022 661018 120204 661254
rect 119604 660934 120204 661018
rect 119604 660698 119786 660934
rect 120022 660698 120204 660934
rect 119604 625254 120204 660698
rect 119604 625018 119786 625254
rect 120022 625018 120204 625254
rect 119604 624934 120204 625018
rect 119604 624698 119786 624934
rect 120022 624698 120204 624934
rect 119604 589254 120204 624698
rect 119604 589018 119786 589254
rect 120022 589018 120204 589254
rect 119604 588934 120204 589018
rect 119604 588698 119786 588934
rect 120022 588698 120204 588934
rect 119604 553254 120204 588698
rect 119604 553018 119786 553254
rect 120022 553018 120204 553254
rect 119604 552934 120204 553018
rect 119604 552698 119786 552934
rect 120022 552698 120204 552934
rect 119604 517254 120204 552698
rect 119604 517018 119786 517254
rect 120022 517018 120204 517254
rect 119604 516934 120204 517018
rect 119604 516698 119786 516934
rect 120022 516698 120204 516934
rect 119604 481254 120204 516698
rect 119604 481018 119786 481254
rect 120022 481018 120204 481254
rect 119604 480934 120204 481018
rect 119604 480698 119786 480934
rect 120022 480698 120204 480934
rect 119604 445254 120204 480698
rect 119604 445018 119786 445254
rect 120022 445018 120204 445254
rect 119604 444934 120204 445018
rect 119604 444698 119786 444934
rect 120022 444698 120204 444934
rect 119604 409254 120204 444698
rect 119604 409018 119786 409254
rect 120022 409018 120204 409254
rect 119604 408934 120204 409018
rect 119604 408698 119786 408934
rect 120022 408698 120204 408934
rect 119604 373254 120204 408698
rect 119604 373018 119786 373254
rect 120022 373018 120204 373254
rect 119604 372934 120204 373018
rect 119604 372698 119786 372934
rect 120022 372698 120204 372934
rect 119604 337254 120204 372698
rect 119604 337018 119786 337254
rect 120022 337018 120204 337254
rect 119604 336934 120204 337018
rect 119604 336698 119786 336934
rect 120022 336698 120204 336934
rect 119604 301254 120204 336698
rect 119604 301018 119786 301254
rect 120022 301018 120204 301254
rect 119604 300934 120204 301018
rect 119604 300698 119786 300934
rect 120022 300698 120204 300934
rect 119604 265254 120204 300698
rect 119604 265018 119786 265254
rect 120022 265018 120204 265254
rect 119604 264934 120204 265018
rect 119604 264698 119786 264934
rect 120022 264698 120204 264934
rect 119604 229254 120204 264698
rect 119604 229018 119786 229254
rect 120022 229018 120204 229254
rect 119604 228934 120204 229018
rect 119604 228698 119786 228934
rect 120022 228698 120204 228934
rect 119604 193254 120204 228698
rect 119604 193018 119786 193254
rect 120022 193018 120204 193254
rect 119604 192934 120204 193018
rect 119604 192698 119786 192934
rect 120022 192698 120204 192934
rect 119604 157254 120204 192698
rect 119604 157018 119786 157254
rect 120022 157018 120204 157254
rect 119604 156934 120204 157018
rect 119604 156698 119786 156934
rect 120022 156698 120204 156934
rect 119604 121254 120204 156698
rect 119604 121018 119786 121254
rect 120022 121018 120204 121254
rect 119604 120934 120204 121018
rect 119604 120698 119786 120934
rect 120022 120698 120204 120934
rect 119604 85254 120204 120698
rect 126804 705778 127404 705800
rect 126804 705542 126986 705778
rect 127222 705542 127404 705778
rect 126804 705458 127404 705542
rect 126804 705222 126986 705458
rect 127222 705222 127404 705458
rect 126804 668454 127404 705222
rect 126804 668218 126986 668454
rect 127222 668218 127404 668454
rect 126804 668134 127404 668218
rect 126804 667898 126986 668134
rect 127222 667898 127404 668134
rect 126804 632454 127404 667898
rect 126804 632218 126986 632454
rect 127222 632218 127404 632454
rect 126804 632134 127404 632218
rect 126804 631898 126986 632134
rect 127222 631898 127404 632134
rect 126804 596454 127404 631898
rect 126804 596218 126986 596454
rect 127222 596218 127404 596454
rect 126804 596134 127404 596218
rect 126804 595898 126986 596134
rect 127222 595898 127404 596134
rect 126804 560454 127404 595898
rect 126804 560218 126986 560454
rect 127222 560218 127404 560454
rect 126804 560134 127404 560218
rect 126804 559898 126986 560134
rect 127222 559898 127404 560134
rect 126804 524454 127404 559898
rect 126804 524218 126986 524454
rect 127222 524218 127404 524454
rect 126804 524134 127404 524218
rect 126804 523898 126986 524134
rect 127222 523898 127404 524134
rect 126804 488454 127404 523898
rect 126804 488218 126986 488454
rect 127222 488218 127404 488454
rect 126804 488134 127404 488218
rect 126804 487898 126986 488134
rect 127222 487898 127404 488134
rect 126804 452454 127404 487898
rect 126804 452218 126986 452454
rect 127222 452218 127404 452454
rect 126804 452134 127404 452218
rect 126804 451898 126986 452134
rect 127222 451898 127404 452134
rect 126804 416454 127404 451898
rect 126804 416218 126986 416454
rect 127222 416218 127404 416454
rect 126804 416134 127404 416218
rect 126804 415898 126986 416134
rect 127222 415898 127404 416134
rect 126804 380454 127404 415898
rect 126804 380218 126986 380454
rect 127222 380218 127404 380454
rect 126804 380134 127404 380218
rect 126804 379898 126986 380134
rect 127222 379898 127404 380134
rect 126804 344454 127404 379898
rect 126804 344218 126986 344454
rect 127222 344218 127404 344454
rect 126804 344134 127404 344218
rect 126804 343898 126986 344134
rect 127222 343898 127404 344134
rect 126804 308454 127404 343898
rect 126804 308218 126986 308454
rect 127222 308218 127404 308454
rect 126804 308134 127404 308218
rect 126804 307898 126986 308134
rect 127222 307898 127404 308134
rect 126804 272454 127404 307898
rect 126804 272218 126986 272454
rect 127222 272218 127404 272454
rect 126804 272134 127404 272218
rect 126804 271898 126986 272134
rect 127222 271898 127404 272134
rect 126804 236454 127404 271898
rect 126804 236218 126986 236454
rect 127222 236218 127404 236454
rect 126804 236134 127404 236218
rect 126804 235898 126986 236134
rect 127222 235898 127404 236134
rect 126804 200454 127404 235898
rect 126804 200218 126986 200454
rect 127222 200218 127404 200454
rect 126804 200134 127404 200218
rect 126804 199898 126986 200134
rect 127222 199898 127404 200134
rect 126804 164454 127404 199898
rect 126804 164218 126986 164454
rect 127222 164218 127404 164454
rect 126804 164134 127404 164218
rect 126804 163898 126986 164134
rect 127222 163898 127404 164134
rect 126804 128454 127404 163898
rect 126804 128218 126986 128454
rect 127222 128218 127404 128454
rect 126804 128134 127404 128218
rect 126804 127898 126986 128134
rect 127222 127898 127404 128134
rect 125547 93940 125613 93941
rect 125547 93876 125548 93940
rect 125612 93876 125613 93940
rect 125547 93875 125613 93876
rect 125550 93669 125610 93875
rect 125547 93668 125613 93669
rect 125547 93604 125548 93668
rect 125612 93604 125613 93668
rect 125547 93603 125613 93604
rect 119604 85018 119786 85254
rect 120022 85018 120204 85254
rect 119604 84934 120204 85018
rect 119604 84698 119786 84934
rect 120022 84698 120204 84934
rect 119604 49254 120204 84698
rect 119604 49018 119786 49254
rect 120022 49018 120204 49254
rect 119604 48934 120204 49018
rect 119604 48698 119786 48934
rect 120022 48698 120204 48934
rect 119604 13254 120204 48698
rect 119604 13018 119786 13254
rect 120022 13018 120204 13254
rect 119604 12934 120204 13018
rect 119604 12698 119786 12934
rect 120022 12698 120204 12934
rect 101604 -7162 101786 -6926
rect 102022 -7162 102204 -6926
rect 101604 -7246 102204 -7162
rect 101604 -7482 101786 -7246
rect 102022 -7482 102204 -7246
rect 101604 -7504 102204 -7482
rect 119604 -5986 120204 12698
rect 126804 92454 127404 127898
rect 126804 92218 126986 92454
rect 127222 92218 127404 92454
rect 126804 92134 127404 92218
rect 126804 91898 126986 92134
rect 127222 91898 127404 92134
rect 126804 56454 127404 91898
rect 126804 56218 126986 56454
rect 127222 56218 127404 56454
rect 126804 56134 127404 56218
rect 126804 55898 126986 56134
rect 127222 55898 127404 56134
rect 126804 20454 127404 55898
rect 126804 20218 126986 20454
rect 127222 20218 127404 20454
rect 126804 20134 127404 20218
rect 126804 19898 126986 20134
rect 127222 19898 127404 20134
rect 126804 -1286 127404 19898
rect 126804 -1522 126986 -1286
rect 127222 -1522 127404 -1286
rect 126804 -1606 127404 -1522
rect 126804 -1842 126986 -1606
rect 127222 -1842 127404 -1606
rect 126804 -1864 127404 -1842
rect 130404 672054 131004 707102
rect 130404 671818 130586 672054
rect 130822 671818 131004 672054
rect 130404 671734 131004 671818
rect 130404 671498 130586 671734
rect 130822 671498 131004 671734
rect 130404 636054 131004 671498
rect 130404 635818 130586 636054
rect 130822 635818 131004 636054
rect 130404 635734 131004 635818
rect 130404 635498 130586 635734
rect 130822 635498 131004 635734
rect 130404 600054 131004 635498
rect 130404 599818 130586 600054
rect 130822 599818 131004 600054
rect 130404 599734 131004 599818
rect 130404 599498 130586 599734
rect 130822 599498 131004 599734
rect 130404 564054 131004 599498
rect 130404 563818 130586 564054
rect 130822 563818 131004 564054
rect 130404 563734 131004 563818
rect 130404 563498 130586 563734
rect 130822 563498 131004 563734
rect 130404 528054 131004 563498
rect 130404 527818 130586 528054
rect 130822 527818 131004 528054
rect 130404 527734 131004 527818
rect 130404 527498 130586 527734
rect 130822 527498 131004 527734
rect 130404 492054 131004 527498
rect 130404 491818 130586 492054
rect 130822 491818 131004 492054
rect 130404 491734 131004 491818
rect 130404 491498 130586 491734
rect 130822 491498 131004 491734
rect 130404 456054 131004 491498
rect 130404 455818 130586 456054
rect 130822 455818 131004 456054
rect 130404 455734 131004 455818
rect 130404 455498 130586 455734
rect 130822 455498 131004 455734
rect 130404 420054 131004 455498
rect 130404 419818 130586 420054
rect 130822 419818 131004 420054
rect 130404 419734 131004 419818
rect 130404 419498 130586 419734
rect 130822 419498 131004 419734
rect 130404 384054 131004 419498
rect 130404 383818 130586 384054
rect 130822 383818 131004 384054
rect 130404 383734 131004 383818
rect 130404 383498 130586 383734
rect 130822 383498 131004 383734
rect 130404 348054 131004 383498
rect 130404 347818 130586 348054
rect 130822 347818 131004 348054
rect 130404 347734 131004 347818
rect 130404 347498 130586 347734
rect 130822 347498 131004 347734
rect 130404 312054 131004 347498
rect 130404 311818 130586 312054
rect 130822 311818 131004 312054
rect 130404 311734 131004 311818
rect 130404 311498 130586 311734
rect 130822 311498 131004 311734
rect 130404 276054 131004 311498
rect 130404 275818 130586 276054
rect 130822 275818 131004 276054
rect 130404 275734 131004 275818
rect 130404 275498 130586 275734
rect 130822 275498 131004 275734
rect 130404 240054 131004 275498
rect 130404 239818 130586 240054
rect 130822 239818 131004 240054
rect 130404 239734 131004 239818
rect 130404 239498 130586 239734
rect 130822 239498 131004 239734
rect 130404 204054 131004 239498
rect 130404 203818 130586 204054
rect 130822 203818 131004 204054
rect 130404 203734 131004 203818
rect 130404 203498 130586 203734
rect 130822 203498 131004 203734
rect 130404 168054 131004 203498
rect 130404 167818 130586 168054
rect 130822 167818 131004 168054
rect 130404 167734 131004 167818
rect 130404 167498 130586 167734
rect 130822 167498 131004 167734
rect 130404 132054 131004 167498
rect 130404 131818 130586 132054
rect 130822 131818 131004 132054
rect 130404 131734 131004 131818
rect 130404 131498 130586 131734
rect 130822 131498 131004 131734
rect 130404 96054 131004 131498
rect 130404 95818 130586 96054
rect 130822 95818 131004 96054
rect 130404 95734 131004 95818
rect 130404 95498 130586 95734
rect 130822 95498 131004 95734
rect 130404 60054 131004 95498
rect 130404 59818 130586 60054
rect 130822 59818 131004 60054
rect 130404 59734 131004 59818
rect 130404 59498 130586 59734
rect 130822 59498 131004 59734
rect 130404 24054 131004 59498
rect 130404 23818 130586 24054
rect 130822 23818 131004 24054
rect 130404 23734 131004 23818
rect 130404 23498 130586 23734
rect 130822 23498 131004 23734
rect 130404 -3166 131004 23498
rect 130404 -3402 130586 -3166
rect 130822 -3402 131004 -3166
rect 130404 -3486 131004 -3402
rect 130404 -3722 130586 -3486
rect 130822 -3722 131004 -3486
rect 130404 -3744 131004 -3722
rect 134004 675654 134604 708982
rect 134004 675418 134186 675654
rect 134422 675418 134604 675654
rect 134004 675334 134604 675418
rect 134004 675098 134186 675334
rect 134422 675098 134604 675334
rect 134004 639654 134604 675098
rect 134004 639418 134186 639654
rect 134422 639418 134604 639654
rect 134004 639334 134604 639418
rect 134004 639098 134186 639334
rect 134422 639098 134604 639334
rect 134004 603654 134604 639098
rect 134004 603418 134186 603654
rect 134422 603418 134604 603654
rect 134004 603334 134604 603418
rect 134004 603098 134186 603334
rect 134422 603098 134604 603334
rect 134004 567654 134604 603098
rect 134004 567418 134186 567654
rect 134422 567418 134604 567654
rect 134004 567334 134604 567418
rect 134004 567098 134186 567334
rect 134422 567098 134604 567334
rect 134004 531654 134604 567098
rect 134004 531418 134186 531654
rect 134422 531418 134604 531654
rect 134004 531334 134604 531418
rect 134004 531098 134186 531334
rect 134422 531098 134604 531334
rect 134004 495654 134604 531098
rect 134004 495418 134186 495654
rect 134422 495418 134604 495654
rect 134004 495334 134604 495418
rect 134004 495098 134186 495334
rect 134422 495098 134604 495334
rect 134004 459654 134604 495098
rect 134004 459418 134186 459654
rect 134422 459418 134604 459654
rect 134004 459334 134604 459418
rect 134004 459098 134186 459334
rect 134422 459098 134604 459334
rect 134004 423654 134604 459098
rect 134004 423418 134186 423654
rect 134422 423418 134604 423654
rect 134004 423334 134604 423418
rect 134004 423098 134186 423334
rect 134422 423098 134604 423334
rect 134004 387654 134604 423098
rect 134004 387418 134186 387654
rect 134422 387418 134604 387654
rect 134004 387334 134604 387418
rect 134004 387098 134186 387334
rect 134422 387098 134604 387334
rect 134004 351654 134604 387098
rect 134004 351418 134186 351654
rect 134422 351418 134604 351654
rect 134004 351334 134604 351418
rect 134004 351098 134186 351334
rect 134422 351098 134604 351334
rect 134004 315654 134604 351098
rect 134004 315418 134186 315654
rect 134422 315418 134604 315654
rect 134004 315334 134604 315418
rect 134004 315098 134186 315334
rect 134422 315098 134604 315334
rect 134004 279654 134604 315098
rect 134004 279418 134186 279654
rect 134422 279418 134604 279654
rect 134004 279334 134604 279418
rect 134004 279098 134186 279334
rect 134422 279098 134604 279334
rect 134004 243654 134604 279098
rect 134004 243418 134186 243654
rect 134422 243418 134604 243654
rect 134004 243334 134604 243418
rect 134004 243098 134186 243334
rect 134422 243098 134604 243334
rect 134004 207654 134604 243098
rect 134004 207418 134186 207654
rect 134422 207418 134604 207654
rect 134004 207334 134604 207418
rect 134004 207098 134186 207334
rect 134422 207098 134604 207334
rect 134004 171654 134604 207098
rect 134004 171418 134186 171654
rect 134422 171418 134604 171654
rect 134004 171334 134604 171418
rect 134004 171098 134186 171334
rect 134422 171098 134604 171334
rect 134004 135654 134604 171098
rect 134004 135418 134186 135654
rect 134422 135418 134604 135654
rect 134004 135334 134604 135418
rect 134004 135098 134186 135334
rect 134422 135098 134604 135334
rect 134004 99654 134604 135098
rect 134004 99418 134186 99654
rect 134422 99418 134604 99654
rect 134004 99334 134604 99418
rect 134004 99098 134186 99334
rect 134422 99098 134604 99334
rect 134004 63654 134604 99098
rect 134004 63418 134186 63654
rect 134422 63418 134604 63654
rect 134004 63334 134604 63418
rect 134004 63098 134186 63334
rect 134422 63098 134604 63334
rect 134004 27654 134604 63098
rect 134004 27418 134186 27654
rect 134422 27418 134604 27654
rect 134004 27334 134604 27418
rect 134004 27098 134186 27334
rect 134422 27098 134604 27334
rect 134004 -5046 134604 27098
rect 134004 -5282 134186 -5046
rect 134422 -5282 134604 -5046
rect 134004 -5366 134604 -5282
rect 134004 -5602 134186 -5366
rect 134422 -5602 134604 -5366
rect 134004 -5624 134604 -5602
rect 137604 679254 138204 710862
rect 155604 710478 156204 711440
rect 155604 710242 155786 710478
rect 156022 710242 156204 710478
rect 155604 710158 156204 710242
rect 155604 709922 155786 710158
rect 156022 709922 156204 710158
rect 152004 708598 152604 709560
rect 152004 708362 152186 708598
rect 152422 708362 152604 708598
rect 152004 708278 152604 708362
rect 152004 708042 152186 708278
rect 152422 708042 152604 708278
rect 148404 706718 149004 707680
rect 148404 706482 148586 706718
rect 148822 706482 149004 706718
rect 148404 706398 149004 706482
rect 148404 706162 148586 706398
rect 148822 706162 149004 706398
rect 137604 679018 137786 679254
rect 138022 679018 138204 679254
rect 137604 678934 138204 679018
rect 137604 678698 137786 678934
rect 138022 678698 138204 678934
rect 137604 643254 138204 678698
rect 137604 643018 137786 643254
rect 138022 643018 138204 643254
rect 137604 642934 138204 643018
rect 137604 642698 137786 642934
rect 138022 642698 138204 642934
rect 137604 607254 138204 642698
rect 137604 607018 137786 607254
rect 138022 607018 138204 607254
rect 137604 606934 138204 607018
rect 137604 606698 137786 606934
rect 138022 606698 138204 606934
rect 137604 571254 138204 606698
rect 137604 571018 137786 571254
rect 138022 571018 138204 571254
rect 137604 570934 138204 571018
rect 137604 570698 137786 570934
rect 138022 570698 138204 570934
rect 137604 535254 138204 570698
rect 137604 535018 137786 535254
rect 138022 535018 138204 535254
rect 137604 534934 138204 535018
rect 137604 534698 137786 534934
rect 138022 534698 138204 534934
rect 137604 499254 138204 534698
rect 137604 499018 137786 499254
rect 138022 499018 138204 499254
rect 137604 498934 138204 499018
rect 137604 498698 137786 498934
rect 138022 498698 138204 498934
rect 137604 463254 138204 498698
rect 137604 463018 137786 463254
rect 138022 463018 138204 463254
rect 137604 462934 138204 463018
rect 137604 462698 137786 462934
rect 138022 462698 138204 462934
rect 137604 427254 138204 462698
rect 137604 427018 137786 427254
rect 138022 427018 138204 427254
rect 137604 426934 138204 427018
rect 137604 426698 137786 426934
rect 138022 426698 138204 426934
rect 137604 391254 138204 426698
rect 137604 391018 137786 391254
rect 138022 391018 138204 391254
rect 137604 390934 138204 391018
rect 137604 390698 137786 390934
rect 138022 390698 138204 390934
rect 137604 355254 138204 390698
rect 137604 355018 137786 355254
rect 138022 355018 138204 355254
rect 137604 354934 138204 355018
rect 137604 354698 137786 354934
rect 138022 354698 138204 354934
rect 137604 319254 138204 354698
rect 137604 319018 137786 319254
rect 138022 319018 138204 319254
rect 137604 318934 138204 319018
rect 137604 318698 137786 318934
rect 138022 318698 138204 318934
rect 137604 283254 138204 318698
rect 137604 283018 137786 283254
rect 138022 283018 138204 283254
rect 137604 282934 138204 283018
rect 137604 282698 137786 282934
rect 138022 282698 138204 282934
rect 137604 247254 138204 282698
rect 137604 247018 137786 247254
rect 138022 247018 138204 247254
rect 137604 246934 138204 247018
rect 137604 246698 137786 246934
rect 138022 246698 138204 246934
rect 137604 211254 138204 246698
rect 137604 211018 137786 211254
rect 138022 211018 138204 211254
rect 137604 210934 138204 211018
rect 137604 210698 137786 210934
rect 138022 210698 138204 210934
rect 137604 175254 138204 210698
rect 137604 175018 137786 175254
rect 138022 175018 138204 175254
rect 137604 174934 138204 175018
rect 137604 174698 137786 174934
rect 138022 174698 138204 174934
rect 137604 139254 138204 174698
rect 137604 139018 137786 139254
rect 138022 139018 138204 139254
rect 137604 138934 138204 139018
rect 137604 138698 137786 138934
rect 138022 138698 138204 138934
rect 137604 103254 138204 138698
rect 137604 103018 137786 103254
rect 138022 103018 138204 103254
rect 137604 102934 138204 103018
rect 137604 102698 137786 102934
rect 138022 102698 138204 102934
rect 137604 67254 138204 102698
rect 137604 67018 137786 67254
rect 138022 67018 138204 67254
rect 137604 66934 138204 67018
rect 137604 66698 137786 66934
rect 138022 66698 138204 66934
rect 137604 31254 138204 66698
rect 137604 31018 137786 31254
rect 138022 31018 138204 31254
rect 137604 30934 138204 31018
rect 137604 30698 137786 30934
rect 138022 30698 138204 30934
rect 119604 -6222 119786 -5986
rect 120022 -6222 120204 -5986
rect 119604 -6306 120204 -6222
rect 119604 -6542 119786 -6306
rect 120022 -6542 120204 -6306
rect 119604 -7504 120204 -6542
rect 137604 -6926 138204 30698
rect 144804 704838 145404 705800
rect 144804 704602 144986 704838
rect 145222 704602 145404 704838
rect 144804 704518 145404 704602
rect 144804 704282 144986 704518
rect 145222 704282 145404 704518
rect 144804 686454 145404 704282
rect 144804 686218 144986 686454
rect 145222 686218 145404 686454
rect 144804 686134 145404 686218
rect 144804 685898 144986 686134
rect 145222 685898 145404 686134
rect 144804 650454 145404 685898
rect 144804 650218 144986 650454
rect 145222 650218 145404 650454
rect 144804 650134 145404 650218
rect 144804 649898 144986 650134
rect 145222 649898 145404 650134
rect 144804 614454 145404 649898
rect 144804 614218 144986 614454
rect 145222 614218 145404 614454
rect 144804 614134 145404 614218
rect 144804 613898 144986 614134
rect 145222 613898 145404 614134
rect 144804 578454 145404 613898
rect 144804 578218 144986 578454
rect 145222 578218 145404 578454
rect 144804 578134 145404 578218
rect 144804 577898 144986 578134
rect 145222 577898 145404 578134
rect 144804 542454 145404 577898
rect 144804 542218 144986 542454
rect 145222 542218 145404 542454
rect 144804 542134 145404 542218
rect 144804 541898 144986 542134
rect 145222 541898 145404 542134
rect 144804 506454 145404 541898
rect 144804 506218 144986 506454
rect 145222 506218 145404 506454
rect 144804 506134 145404 506218
rect 144804 505898 144986 506134
rect 145222 505898 145404 506134
rect 144804 470454 145404 505898
rect 144804 470218 144986 470454
rect 145222 470218 145404 470454
rect 144804 470134 145404 470218
rect 144804 469898 144986 470134
rect 145222 469898 145404 470134
rect 144804 434454 145404 469898
rect 144804 434218 144986 434454
rect 145222 434218 145404 434454
rect 144804 434134 145404 434218
rect 144804 433898 144986 434134
rect 145222 433898 145404 434134
rect 144804 398454 145404 433898
rect 144804 398218 144986 398454
rect 145222 398218 145404 398454
rect 144804 398134 145404 398218
rect 144804 397898 144986 398134
rect 145222 397898 145404 398134
rect 144804 362454 145404 397898
rect 144804 362218 144986 362454
rect 145222 362218 145404 362454
rect 144804 362134 145404 362218
rect 144804 361898 144986 362134
rect 145222 361898 145404 362134
rect 144804 326454 145404 361898
rect 144804 326218 144986 326454
rect 145222 326218 145404 326454
rect 144804 326134 145404 326218
rect 144804 325898 144986 326134
rect 145222 325898 145404 326134
rect 144804 290454 145404 325898
rect 144804 290218 144986 290454
rect 145222 290218 145404 290454
rect 144804 290134 145404 290218
rect 144804 289898 144986 290134
rect 145222 289898 145404 290134
rect 144804 254454 145404 289898
rect 144804 254218 144986 254454
rect 145222 254218 145404 254454
rect 144804 254134 145404 254218
rect 144804 253898 144986 254134
rect 145222 253898 145404 254134
rect 144804 218454 145404 253898
rect 144804 218218 144986 218454
rect 145222 218218 145404 218454
rect 144804 218134 145404 218218
rect 144804 217898 144986 218134
rect 145222 217898 145404 218134
rect 144804 182454 145404 217898
rect 144804 182218 144986 182454
rect 145222 182218 145404 182454
rect 144804 182134 145404 182218
rect 144804 181898 144986 182134
rect 145222 181898 145404 182134
rect 144804 146454 145404 181898
rect 144804 146218 144986 146454
rect 145222 146218 145404 146454
rect 144804 146134 145404 146218
rect 144804 145898 144986 146134
rect 145222 145898 145404 146134
rect 144804 110454 145404 145898
rect 144804 110218 144986 110454
rect 145222 110218 145404 110454
rect 144804 110134 145404 110218
rect 144804 109898 144986 110134
rect 145222 109898 145404 110134
rect 144804 74454 145404 109898
rect 144804 74218 144986 74454
rect 145222 74218 145404 74454
rect 144804 74134 145404 74218
rect 144804 73898 144986 74134
rect 145222 73898 145404 74134
rect 144804 38454 145404 73898
rect 144804 38218 144986 38454
rect 145222 38218 145404 38454
rect 144804 38134 145404 38218
rect 144804 37898 144986 38134
rect 145222 37898 145404 38134
rect 144804 2454 145404 37898
rect 144804 2218 144986 2454
rect 145222 2218 145404 2454
rect 144804 2134 145404 2218
rect 144804 1898 144986 2134
rect 145222 1898 145404 2134
rect 144804 -346 145404 1898
rect 144804 -582 144986 -346
rect 145222 -582 145404 -346
rect 144804 -666 145404 -582
rect 144804 -902 144986 -666
rect 145222 -902 145404 -666
rect 144804 -1864 145404 -902
rect 148404 690054 149004 706162
rect 148404 689818 148586 690054
rect 148822 689818 149004 690054
rect 148404 689734 149004 689818
rect 148404 689498 148586 689734
rect 148822 689498 149004 689734
rect 148404 654054 149004 689498
rect 148404 653818 148586 654054
rect 148822 653818 149004 654054
rect 148404 653734 149004 653818
rect 148404 653498 148586 653734
rect 148822 653498 149004 653734
rect 148404 618054 149004 653498
rect 148404 617818 148586 618054
rect 148822 617818 149004 618054
rect 148404 617734 149004 617818
rect 148404 617498 148586 617734
rect 148822 617498 149004 617734
rect 148404 582054 149004 617498
rect 148404 581818 148586 582054
rect 148822 581818 149004 582054
rect 148404 581734 149004 581818
rect 148404 581498 148586 581734
rect 148822 581498 149004 581734
rect 148404 546054 149004 581498
rect 148404 545818 148586 546054
rect 148822 545818 149004 546054
rect 148404 545734 149004 545818
rect 148404 545498 148586 545734
rect 148822 545498 149004 545734
rect 148404 510054 149004 545498
rect 148404 509818 148586 510054
rect 148822 509818 149004 510054
rect 148404 509734 149004 509818
rect 148404 509498 148586 509734
rect 148822 509498 149004 509734
rect 148404 474054 149004 509498
rect 148404 473818 148586 474054
rect 148822 473818 149004 474054
rect 148404 473734 149004 473818
rect 148404 473498 148586 473734
rect 148822 473498 149004 473734
rect 148404 438054 149004 473498
rect 148404 437818 148586 438054
rect 148822 437818 149004 438054
rect 148404 437734 149004 437818
rect 148404 437498 148586 437734
rect 148822 437498 149004 437734
rect 148404 402054 149004 437498
rect 148404 401818 148586 402054
rect 148822 401818 149004 402054
rect 148404 401734 149004 401818
rect 148404 401498 148586 401734
rect 148822 401498 149004 401734
rect 148404 366054 149004 401498
rect 148404 365818 148586 366054
rect 148822 365818 149004 366054
rect 148404 365734 149004 365818
rect 148404 365498 148586 365734
rect 148822 365498 149004 365734
rect 148404 330054 149004 365498
rect 148404 329818 148586 330054
rect 148822 329818 149004 330054
rect 148404 329734 149004 329818
rect 148404 329498 148586 329734
rect 148822 329498 149004 329734
rect 148404 294054 149004 329498
rect 148404 293818 148586 294054
rect 148822 293818 149004 294054
rect 148404 293734 149004 293818
rect 148404 293498 148586 293734
rect 148822 293498 149004 293734
rect 148404 258054 149004 293498
rect 148404 257818 148586 258054
rect 148822 257818 149004 258054
rect 148404 257734 149004 257818
rect 148404 257498 148586 257734
rect 148822 257498 149004 257734
rect 148404 222054 149004 257498
rect 148404 221818 148586 222054
rect 148822 221818 149004 222054
rect 148404 221734 149004 221818
rect 148404 221498 148586 221734
rect 148822 221498 149004 221734
rect 148404 186054 149004 221498
rect 148404 185818 148586 186054
rect 148822 185818 149004 186054
rect 148404 185734 149004 185818
rect 148404 185498 148586 185734
rect 148822 185498 149004 185734
rect 148404 150054 149004 185498
rect 148404 149818 148586 150054
rect 148822 149818 149004 150054
rect 148404 149734 149004 149818
rect 148404 149498 148586 149734
rect 148822 149498 149004 149734
rect 148404 114054 149004 149498
rect 148404 113818 148586 114054
rect 148822 113818 149004 114054
rect 148404 113734 149004 113818
rect 148404 113498 148586 113734
rect 148822 113498 149004 113734
rect 148404 78054 149004 113498
rect 148404 77818 148586 78054
rect 148822 77818 149004 78054
rect 148404 77734 149004 77818
rect 148404 77498 148586 77734
rect 148822 77498 149004 77734
rect 148404 42054 149004 77498
rect 148404 41818 148586 42054
rect 148822 41818 149004 42054
rect 148404 41734 149004 41818
rect 148404 41498 148586 41734
rect 148822 41498 149004 41734
rect 148404 6054 149004 41498
rect 148404 5818 148586 6054
rect 148822 5818 149004 6054
rect 148404 5734 149004 5818
rect 148404 5498 148586 5734
rect 148822 5498 149004 5734
rect 148404 -2226 149004 5498
rect 148404 -2462 148586 -2226
rect 148822 -2462 149004 -2226
rect 148404 -2546 149004 -2462
rect 148404 -2782 148586 -2546
rect 148822 -2782 149004 -2546
rect 148404 -3744 149004 -2782
rect 152004 693654 152604 708042
rect 152004 693418 152186 693654
rect 152422 693418 152604 693654
rect 152004 693334 152604 693418
rect 152004 693098 152186 693334
rect 152422 693098 152604 693334
rect 152004 657654 152604 693098
rect 152004 657418 152186 657654
rect 152422 657418 152604 657654
rect 152004 657334 152604 657418
rect 152004 657098 152186 657334
rect 152422 657098 152604 657334
rect 152004 621654 152604 657098
rect 152004 621418 152186 621654
rect 152422 621418 152604 621654
rect 152004 621334 152604 621418
rect 152004 621098 152186 621334
rect 152422 621098 152604 621334
rect 152004 585654 152604 621098
rect 152004 585418 152186 585654
rect 152422 585418 152604 585654
rect 152004 585334 152604 585418
rect 152004 585098 152186 585334
rect 152422 585098 152604 585334
rect 152004 549654 152604 585098
rect 152004 549418 152186 549654
rect 152422 549418 152604 549654
rect 152004 549334 152604 549418
rect 152004 549098 152186 549334
rect 152422 549098 152604 549334
rect 152004 513654 152604 549098
rect 152004 513418 152186 513654
rect 152422 513418 152604 513654
rect 152004 513334 152604 513418
rect 152004 513098 152186 513334
rect 152422 513098 152604 513334
rect 152004 477654 152604 513098
rect 152004 477418 152186 477654
rect 152422 477418 152604 477654
rect 152004 477334 152604 477418
rect 152004 477098 152186 477334
rect 152422 477098 152604 477334
rect 152004 441654 152604 477098
rect 152004 441418 152186 441654
rect 152422 441418 152604 441654
rect 152004 441334 152604 441418
rect 152004 441098 152186 441334
rect 152422 441098 152604 441334
rect 152004 405654 152604 441098
rect 152004 405418 152186 405654
rect 152422 405418 152604 405654
rect 152004 405334 152604 405418
rect 152004 405098 152186 405334
rect 152422 405098 152604 405334
rect 152004 369654 152604 405098
rect 152004 369418 152186 369654
rect 152422 369418 152604 369654
rect 152004 369334 152604 369418
rect 152004 369098 152186 369334
rect 152422 369098 152604 369334
rect 152004 333654 152604 369098
rect 152004 333418 152186 333654
rect 152422 333418 152604 333654
rect 152004 333334 152604 333418
rect 152004 333098 152186 333334
rect 152422 333098 152604 333334
rect 152004 297654 152604 333098
rect 152004 297418 152186 297654
rect 152422 297418 152604 297654
rect 152004 297334 152604 297418
rect 152004 297098 152186 297334
rect 152422 297098 152604 297334
rect 152004 261654 152604 297098
rect 152004 261418 152186 261654
rect 152422 261418 152604 261654
rect 152004 261334 152604 261418
rect 152004 261098 152186 261334
rect 152422 261098 152604 261334
rect 152004 225654 152604 261098
rect 152004 225418 152186 225654
rect 152422 225418 152604 225654
rect 152004 225334 152604 225418
rect 152004 225098 152186 225334
rect 152422 225098 152604 225334
rect 152004 189654 152604 225098
rect 152004 189418 152186 189654
rect 152422 189418 152604 189654
rect 152004 189334 152604 189418
rect 152004 189098 152186 189334
rect 152422 189098 152604 189334
rect 152004 153654 152604 189098
rect 152004 153418 152186 153654
rect 152422 153418 152604 153654
rect 152004 153334 152604 153418
rect 152004 153098 152186 153334
rect 152422 153098 152604 153334
rect 152004 117654 152604 153098
rect 152004 117418 152186 117654
rect 152422 117418 152604 117654
rect 152004 117334 152604 117418
rect 152004 117098 152186 117334
rect 152422 117098 152604 117334
rect 152004 81654 152604 117098
rect 152004 81418 152186 81654
rect 152422 81418 152604 81654
rect 152004 81334 152604 81418
rect 152004 81098 152186 81334
rect 152422 81098 152604 81334
rect 152004 45654 152604 81098
rect 152004 45418 152186 45654
rect 152422 45418 152604 45654
rect 152004 45334 152604 45418
rect 152004 45098 152186 45334
rect 152422 45098 152604 45334
rect 152004 9654 152604 45098
rect 152004 9418 152186 9654
rect 152422 9418 152604 9654
rect 152004 9334 152604 9418
rect 152004 9098 152186 9334
rect 152422 9098 152604 9334
rect 152004 -4106 152604 9098
rect 152004 -4342 152186 -4106
rect 152422 -4342 152604 -4106
rect 152004 -4426 152604 -4342
rect 152004 -4662 152186 -4426
rect 152422 -4662 152604 -4426
rect 152004 -5624 152604 -4662
rect 155604 697254 156204 709922
rect 173604 711418 174204 711440
rect 173604 711182 173786 711418
rect 174022 711182 174204 711418
rect 173604 711098 174204 711182
rect 173604 710862 173786 711098
rect 174022 710862 174204 711098
rect 170004 709538 170604 709560
rect 170004 709302 170186 709538
rect 170422 709302 170604 709538
rect 170004 709218 170604 709302
rect 170004 708982 170186 709218
rect 170422 708982 170604 709218
rect 166404 707658 167004 707680
rect 166404 707422 166586 707658
rect 166822 707422 167004 707658
rect 166404 707338 167004 707422
rect 166404 707102 166586 707338
rect 166822 707102 167004 707338
rect 155604 697018 155786 697254
rect 156022 697018 156204 697254
rect 155604 696934 156204 697018
rect 155604 696698 155786 696934
rect 156022 696698 156204 696934
rect 155604 661254 156204 696698
rect 155604 661018 155786 661254
rect 156022 661018 156204 661254
rect 155604 660934 156204 661018
rect 155604 660698 155786 660934
rect 156022 660698 156204 660934
rect 155604 625254 156204 660698
rect 155604 625018 155786 625254
rect 156022 625018 156204 625254
rect 155604 624934 156204 625018
rect 155604 624698 155786 624934
rect 156022 624698 156204 624934
rect 155604 589254 156204 624698
rect 155604 589018 155786 589254
rect 156022 589018 156204 589254
rect 155604 588934 156204 589018
rect 155604 588698 155786 588934
rect 156022 588698 156204 588934
rect 155604 553254 156204 588698
rect 155604 553018 155786 553254
rect 156022 553018 156204 553254
rect 155604 552934 156204 553018
rect 155604 552698 155786 552934
rect 156022 552698 156204 552934
rect 155604 517254 156204 552698
rect 155604 517018 155786 517254
rect 156022 517018 156204 517254
rect 155604 516934 156204 517018
rect 155604 516698 155786 516934
rect 156022 516698 156204 516934
rect 155604 481254 156204 516698
rect 155604 481018 155786 481254
rect 156022 481018 156204 481254
rect 155604 480934 156204 481018
rect 155604 480698 155786 480934
rect 156022 480698 156204 480934
rect 155604 445254 156204 480698
rect 155604 445018 155786 445254
rect 156022 445018 156204 445254
rect 155604 444934 156204 445018
rect 155604 444698 155786 444934
rect 156022 444698 156204 444934
rect 155604 409254 156204 444698
rect 155604 409018 155786 409254
rect 156022 409018 156204 409254
rect 155604 408934 156204 409018
rect 155604 408698 155786 408934
rect 156022 408698 156204 408934
rect 155604 373254 156204 408698
rect 155604 373018 155786 373254
rect 156022 373018 156204 373254
rect 155604 372934 156204 373018
rect 155604 372698 155786 372934
rect 156022 372698 156204 372934
rect 155604 337254 156204 372698
rect 155604 337018 155786 337254
rect 156022 337018 156204 337254
rect 155604 336934 156204 337018
rect 155604 336698 155786 336934
rect 156022 336698 156204 336934
rect 155604 301254 156204 336698
rect 155604 301018 155786 301254
rect 156022 301018 156204 301254
rect 155604 300934 156204 301018
rect 155604 300698 155786 300934
rect 156022 300698 156204 300934
rect 155604 265254 156204 300698
rect 155604 265018 155786 265254
rect 156022 265018 156204 265254
rect 155604 264934 156204 265018
rect 155604 264698 155786 264934
rect 156022 264698 156204 264934
rect 155604 229254 156204 264698
rect 155604 229018 155786 229254
rect 156022 229018 156204 229254
rect 155604 228934 156204 229018
rect 155604 228698 155786 228934
rect 156022 228698 156204 228934
rect 155604 193254 156204 228698
rect 155604 193018 155786 193254
rect 156022 193018 156204 193254
rect 155604 192934 156204 193018
rect 155604 192698 155786 192934
rect 156022 192698 156204 192934
rect 155604 157254 156204 192698
rect 155604 157018 155786 157254
rect 156022 157018 156204 157254
rect 155604 156934 156204 157018
rect 155604 156698 155786 156934
rect 156022 156698 156204 156934
rect 155604 121254 156204 156698
rect 155604 121018 155786 121254
rect 156022 121018 156204 121254
rect 155604 120934 156204 121018
rect 155604 120698 155786 120934
rect 156022 120698 156204 120934
rect 155604 85254 156204 120698
rect 155604 85018 155786 85254
rect 156022 85018 156204 85254
rect 155604 84934 156204 85018
rect 155604 84698 155786 84934
rect 156022 84698 156204 84934
rect 155604 49254 156204 84698
rect 155604 49018 155786 49254
rect 156022 49018 156204 49254
rect 155604 48934 156204 49018
rect 155604 48698 155786 48934
rect 156022 48698 156204 48934
rect 155604 13254 156204 48698
rect 155604 13018 155786 13254
rect 156022 13018 156204 13254
rect 155604 12934 156204 13018
rect 155604 12698 155786 12934
rect 156022 12698 156204 12934
rect 137604 -7162 137786 -6926
rect 138022 -7162 138204 -6926
rect 137604 -7246 138204 -7162
rect 137604 -7482 137786 -7246
rect 138022 -7482 138204 -7246
rect 137604 -7504 138204 -7482
rect 155604 -5986 156204 12698
rect 162804 705778 163404 705800
rect 162804 705542 162986 705778
rect 163222 705542 163404 705778
rect 162804 705458 163404 705542
rect 162804 705222 162986 705458
rect 163222 705222 163404 705458
rect 162804 668454 163404 705222
rect 162804 668218 162986 668454
rect 163222 668218 163404 668454
rect 162804 668134 163404 668218
rect 162804 667898 162986 668134
rect 163222 667898 163404 668134
rect 162804 632454 163404 667898
rect 162804 632218 162986 632454
rect 163222 632218 163404 632454
rect 162804 632134 163404 632218
rect 162804 631898 162986 632134
rect 163222 631898 163404 632134
rect 162804 596454 163404 631898
rect 162804 596218 162986 596454
rect 163222 596218 163404 596454
rect 162804 596134 163404 596218
rect 162804 595898 162986 596134
rect 163222 595898 163404 596134
rect 162804 560454 163404 595898
rect 162804 560218 162986 560454
rect 163222 560218 163404 560454
rect 162804 560134 163404 560218
rect 162804 559898 162986 560134
rect 163222 559898 163404 560134
rect 162804 524454 163404 559898
rect 162804 524218 162986 524454
rect 163222 524218 163404 524454
rect 162804 524134 163404 524218
rect 162804 523898 162986 524134
rect 163222 523898 163404 524134
rect 162804 488454 163404 523898
rect 162804 488218 162986 488454
rect 163222 488218 163404 488454
rect 162804 488134 163404 488218
rect 162804 487898 162986 488134
rect 163222 487898 163404 488134
rect 162804 452454 163404 487898
rect 162804 452218 162986 452454
rect 163222 452218 163404 452454
rect 162804 452134 163404 452218
rect 162804 451898 162986 452134
rect 163222 451898 163404 452134
rect 162804 416454 163404 451898
rect 162804 416218 162986 416454
rect 163222 416218 163404 416454
rect 162804 416134 163404 416218
rect 162804 415898 162986 416134
rect 163222 415898 163404 416134
rect 162804 380454 163404 415898
rect 162804 380218 162986 380454
rect 163222 380218 163404 380454
rect 162804 380134 163404 380218
rect 162804 379898 162986 380134
rect 163222 379898 163404 380134
rect 162804 344454 163404 379898
rect 162804 344218 162986 344454
rect 163222 344218 163404 344454
rect 162804 344134 163404 344218
rect 162804 343898 162986 344134
rect 163222 343898 163404 344134
rect 162804 308454 163404 343898
rect 162804 308218 162986 308454
rect 163222 308218 163404 308454
rect 162804 308134 163404 308218
rect 162804 307898 162986 308134
rect 163222 307898 163404 308134
rect 162804 272454 163404 307898
rect 162804 272218 162986 272454
rect 163222 272218 163404 272454
rect 162804 272134 163404 272218
rect 162804 271898 162986 272134
rect 163222 271898 163404 272134
rect 162804 236454 163404 271898
rect 162804 236218 162986 236454
rect 163222 236218 163404 236454
rect 162804 236134 163404 236218
rect 162804 235898 162986 236134
rect 163222 235898 163404 236134
rect 162804 200454 163404 235898
rect 162804 200218 162986 200454
rect 163222 200218 163404 200454
rect 162804 200134 163404 200218
rect 162804 199898 162986 200134
rect 163222 199898 163404 200134
rect 162804 164454 163404 199898
rect 162804 164218 162986 164454
rect 163222 164218 163404 164454
rect 162804 164134 163404 164218
rect 162804 163898 162986 164134
rect 163222 163898 163404 164134
rect 162804 128454 163404 163898
rect 162804 128218 162986 128454
rect 163222 128218 163404 128454
rect 162804 128134 163404 128218
rect 162804 127898 162986 128134
rect 163222 127898 163404 128134
rect 162804 92454 163404 127898
rect 162804 92218 162986 92454
rect 163222 92218 163404 92454
rect 162804 92134 163404 92218
rect 162804 91898 162986 92134
rect 163222 91898 163404 92134
rect 162804 56454 163404 91898
rect 162804 56218 162986 56454
rect 163222 56218 163404 56454
rect 162804 56134 163404 56218
rect 162804 55898 162986 56134
rect 163222 55898 163404 56134
rect 162804 20454 163404 55898
rect 162804 20218 162986 20454
rect 163222 20218 163404 20454
rect 162804 20134 163404 20218
rect 162804 19898 162986 20134
rect 163222 19898 163404 20134
rect 162804 -1286 163404 19898
rect 162804 -1522 162986 -1286
rect 163222 -1522 163404 -1286
rect 162804 -1606 163404 -1522
rect 162804 -1842 162986 -1606
rect 163222 -1842 163404 -1606
rect 162804 -1864 163404 -1842
rect 166404 672054 167004 707102
rect 166404 671818 166586 672054
rect 166822 671818 167004 672054
rect 166404 671734 167004 671818
rect 166404 671498 166586 671734
rect 166822 671498 167004 671734
rect 166404 636054 167004 671498
rect 166404 635818 166586 636054
rect 166822 635818 167004 636054
rect 166404 635734 167004 635818
rect 166404 635498 166586 635734
rect 166822 635498 167004 635734
rect 166404 600054 167004 635498
rect 166404 599818 166586 600054
rect 166822 599818 167004 600054
rect 166404 599734 167004 599818
rect 166404 599498 166586 599734
rect 166822 599498 167004 599734
rect 166404 564054 167004 599498
rect 166404 563818 166586 564054
rect 166822 563818 167004 564054
rect 166404 563734 167004 563818
rect 166404 563498 166586 563734
rect 166822 563498 167004 563734
rect 166404 528054 167004 563498
rect 166404 527818 166586 528054
rect 166822 527818 167004 528054
rect 166404 527734 167004 527818
rect 166404 527498 166586 527734
rect 166822 527498 167004 527734
rect 166404 492054 167004 527498
rect 166404 491818 166586 492054
rect 166822 491818 167004 492054
rect 166404 491734 167004 491818
rect 166404 491498 166586 491734
rect 166822 491498 167004 491734
rect 166404 456054 167004 491498
rect 166404 455818 166586 456054
rect 166822 455818 167004 456054
rect 166404 455734 167004 455818
rect 166404 455498 166586 455734
rect 166822 455498 167004 455734
rect 166404 420054 167004 455498
rect 166404 419818 166586 420054
rect 166822 419818 167004 420054
rect 166404 419734 167004 419818
rect 166404 419498 166586 419734
rect 166822 419498 167004 419734
rect 166404 384054 167004 419498
rect 166404 383818 166586 384054
rect 166822 383818 167004 384054
rect 166404 383734 167004 383818
rect 166404 383498 166586 383734
rect 166822 383498 167004 383734
rect 166404 348054 167004 383498
rect 166404 347818 166586 348054
rect 166822 347818 167004 348054
rect 166404 347734 167004 347818
rect 166404 347498 166586 347734
rect 166822 347498 167004 347734
rect 166404 312054 167004 347498
rect 166404 311818 166586 312054
rect 166822 311818 167004 312054
rect 166404 311734 167004 311818
rect 166404 311498 166586 311734
rect 166822 311498 167004 311734
rect 166404 276054 167004 311498
rect 166404 275818 166586 276054
rect 166822 275818 167004 276054
rect 166404 275734 167004 275818
rect 166404 275498 166586 275734
rect 166822 275498 167004 275734
rect 166404 240054 167004 275498
rect 166404 239818 166586 240054
rect 166822 239818 167004 240054
rect 166404 239734 167004 239818
rect 166404 239498 166586 239734
rect 166822 239498 167004 239734
rect 166404 204054 167004 239498
rect 166404 203818 166586 204054
rect 166822 203818 167004 204054
rect 166404 203734 167004 203818
rect 166404 203498 166586 203734
rect 166822 203498 167004 203734
rect 166404 168054 167004 203498
rect 166404 167818 166586 168054
rect 166822 167818 167004 168054
rect 166404 167734 167004 167818
rect 166404 167498 166586 167734
rect 166822 167498 167004 167734
rect 166404 132054 167004 167498
rect 166404 131818 166586 132054
rect 166822 131818 167004 132054
rect 166404 131734 167004 131818
rect 166404 131498 166586 131734
rect 166822 131498 167004 131734
rect 166404 96054 167004 131498
rect 166404 95818 166586 96054
rect 166822 95818 167004 96054
rect 166404 95734 167004 95818
rect 166404 95498 166586 95734
rect 166822 95498 167004 95734
rect 166404 60054 167004 95498
rect 166404 59818 166586 60054
rect 166822 59818 167004 60054
rect 166404 59734 167004 59818
rect 166404 59498 166586 59734
rect 166822 59498 167004 59734
rect 166404 24054 167004 59498
rect 166404 23818 166586 24054
rect 166822 23818 167004 24054
rect 166404 23734 167004 23818
rect 166404 23498 166586 23734
rect 166822 23498 167004 23734
rect 166404 -3166 167004 23498
rect 166404 -3402 166586 -3166
rect 166822 -3402 167004 -3166
rect 166404 -3486 167004 -3402
rect 166404 -3722 166586 -3486
rect 166822 -3722 167004 -3486
rect 166404 -3744 167004 -3722
rect 170004 675654 170604 708982
rect 170004 675418 170186 675654
rect 170422 675418 170604 675654
rect 170004 675334 170604 675418
rect 170004 675098 170186 675334
rect 170422 675098 170604 675334
rect 170004 639654 170604 675098
rect 170004 639418 170186 639654
rect 170422 639418 170604 639654
rect 170004 639334 170604 639418
rect 170004 639098 170186 639334
rect 170422 639098 170604 639334
rect 170004 603654 170604 639098
rect 170004 603418 170186 603654
rect 170422 603418 170604 603654
rect 170004 603334 170604 603418
rect 170004 603098 170186 603334
rect 170422 603098 170604 603334
rect 170004 567654 170604 603098
rect 170004 567418 170186 567654
rect 170422 567418 170604 567654
rect 170004 567334 170604 567418
rect 170004 567098 170186 567334
rect 170422 567098 170604 567334
rect 170004 531654 170604 567098
rect 170004 531418 170186 531654
rect 170422 531418 170604 531654
rect 170004 531334 170604 531418
rect 170004 531098 170186 531334
rect 170422 531098 170604 531334
rect 170004 495654 170604 531098
rect 170004 495418 170186 495654
rect 170422 495418 170604 495654
rect 170004 495334 170604 495418
rect 170004 495098 170186 495334
rect 170422 495098 170604 495334
rect 170004 459654 170604 495098
rect 170004 459418 170186 459654
rect 170422 459418 170604 459654
rect 170004 459334 170604 459418
rect 170004 459098 170186 459334
rect 170422 459098 170604 459334
rect 170004 423654 170604 459098
rect 170004 423418 170186 423654
rect 170422 423418 170604 423654
rect 170004 423334 170604 423418
rect 170004 423098 170186 423334
rect 170422 423098 170604 423334
rect 170004 387654 170604 423098
rect 170004 387418 170186 387654
rect 170422 387418 170604 387654
rect 170004 387334 170604 387418
rect 170004 387098 170186 387334
rect 170422 387098 170604 387334
rect 170004 351654 170604 387098
rect 170004 351418 170186 351654
rect 170422 351418 170604 351654
rect 170004 351334 170604 351418
rect 170004 351098 170186 351334
rect 170422 351098 170604 351334
rect 170004 315654 170604 351098
rect 170004 315418 170186 315654
rect 170422 315418 170604 315654
rect 170004 315334 170604 315418
rect 170004 315098 170186 315334
rect 170422 315098 170604 315334
rect 170004 279654 170604 315098
rect 170004 279418 170186 279654
rect 170422 279418 170604 279654
rect 170004 279334 170604 279418
rect 170004 279098 170186 279334
rect 170422 279098 170604 279334
rect 170004 243654 170604 279098
rect 170004 243418 170186 243654
rect 170422 243418 170604 243654
rect 170004 243334 170604 243418
rect 170004 243098 170186 243334
rect 170422 243098 170604 243334
rect 170004 207654 170604 243098
rect 170004 207418 170186 207654
rect 170422 207418 170604 207654
rect 170004 207334 170604 207418
rect 170004 207098 170186 207334
rect 170422 207098 170604 207334
rect 170004 171654 170604 207098
rect 170004 171418 170186 171654
rect 170422 171418 170604 171654
rect 170004 171334 170604 171418
rect 170004 171098 170186 171334
rect 170422 171098 170604 171334
rect 170004 135654 170604 171098
rect 170004 135418 170186 135654
rect 170422 135418 170604 135654
rect 170004 135334 170604 135418
rect 170004 135098 170186 135334
rect 170422 135098 170604 135334
rect 170004 99654 170604 135098
rect 170004 99418 170186 99654
rect 170422 99418 170604 99654
rect 170004 99334 170604 99418
rect 170004 99098 170186 99334
rect 170422 99098 170604 99334
rect 170004 63654 170604 99098
rect 170004 63418 170186 63654
rect 170422 63418 170604 63654
rect 170004 63334 170604 63418
rect 170004 63098 170186 63334
rect 170422 63098 170604 63334
rect 170004 27654 170604 63098
rect 170004 27418 170186 27654
rect 170422 27418 170604 27654
rect 170004 27334 170604 27418
rect 170004 27098 170186 27334
rect 170422 27098 170604 27334
rect 170004 -5046 170604 27098
rect 170004 -5282 170186 -5046
rect 170422 -5282 170604 -5046
rect 170004 -5366 170604 -5282
rect 170004 -5602 170186 -5366
rect 170422 -5602 170604 -5366
rect 170004 -5624 170604 -5602
rect 173604 679254 174204 710862
rect 191604 710478 192204 711440
rect 191604 710242 191786 710478
rect 192022 710242 192204 710478
rect 191604 710158 192204 710242
rect 191604 709922 191786 710158
rect 192022 709922 192204 710158
rect 188004 708598 188604 709560
rect 188004 708362 188186 708598
rect 188422 708362 188604 708598
rect 188004 708278 188604 708362
rect 188004 708042 188186 708278
rect 188422 708042 188604 708278
rect 184404 706718 185004 707680
rect 184404 706482 184586 706718
rect 184822 706482 185004 706718
rect 184404 706398 185004 706482
rect 184404 706162 184586 706398
rect 184822 706162 185004 706398
rect 173604 679018 173786 679254
rect 174022 679018 174204 679254
rect 173604 678934 174204 679018
rect 173604 678698 173786 678934
rect 174022 678698 174204 678934
rect 173604 643254 174204 678698
rect 173604 643018 173786 643254
rect 174022 643018 174204 643254
rect 173604 642934 174204 643018
rect 173604 642698 173786 642934
rect 174022 642698 174204 642934
rect 173604 607254 174204 642698
rect 173604 607018 173786 607254
rect 174022 607018 174204 607254
rect 173604 606934 174204 607018
rect 173604 606698 173786 606934
rect 174022 606698 174204 606934
rect 173604 571254 174204 606698
rect 173604 571018 173786 571254
rect 174022 571018 174204 571254
rect 173604 570934 174204 571018
rect 173604 570698 173786 570934
rect 174022 570698 174204 570934
rect 173604 535254 174204 570698
rect 173604 535018 173786 535254
rect 174022 535018 174204 535254
rect 173604 534934 174204 535018
rect 173604 534698 173786 534934
rect 174022 534698 174204 534934
rect 173604 499254 174204 534698
rect 173604 499018 173786 499254
rect 174022 499018 174204 499254
rect 173604 498934 174204 499018
rect 173604 498698 173786 498934
rect 174022 498698 174204 498934
rect 173604 463254 174204 498698
rect 173604 463018 173786 463254
rect 174022 463018 174204 463254
rect 173604 462934 174204 463018
rect 173604 462698 173786 462934
rect 174022 462698 174204 462934
rect 173604 427254 174204 462698
rect 173604 427018 173786 427254
rect 174022 427018 174204 427254
rect 173604 426934 174204 427018
rect 173604 426698 173786 426934
rect 174022 426698 174204 426934
rect 173604 391254 174204 426698
rect 173604 391018 173786 391254
rect 174022 391018 174204 391254
rect 173604 390934 174204 391018
rect 173604 390698 173786 390934
rect 174022 390698 174204 390934
rect 173604 355254 174204 390698
rect 173604 355018 173786 355254
rect 174022 355018 174204 355254
rect 173604 354934 174204 355018
rect 173604 354698 173786 354934
rect 174022 354698 174204 354934
rect 173604 319254 174204 354698
rect 173604 319018 173786 319254
rect 174022 319018 174204 319254
rect 173604 318934 174204 319018
rect 173604 318698 173786 318934
rect 174022 318698 174204 318934
rect 173604 283254 174204 318698
rect 173604 283018 173786 283254
rect 174022 283018 174204 283254
rect 173604 282934 174204 283018
rect 173604 282698 173786 282934
rect 174022 282698 174204 282934
rect 173604 247254 174204 282698
rect 173604 247018 173786 247254
rect 174022 247018 174204 247254
rect 173604 246934 174204 247018
rect 173604 246698 173786 246934
rect 174022 246698 174204 246934
rect 173604 211254 174204 246698
rect 173604 211018 173786 211254
rect 174022 211018 174204 211254
rect 173604 210934 174204 211018
rect 173604 210698 173786 210934
rect 174022 210698 174204 210934
rect 173604 175254 174204 210698
rect 173604 175018 173786 175254
rect 174022 175018 174204 175254
rect 173604 174934 174204 175018
rect 173604 174698 173786 174934
rect 174022 174698 174204 174934
rect 173604 139254 174204 174698
rect 173604 139018 173786 139254
rect 174022 139018 174204 139254
rect 173604 138934 174204 139018
rect 173604 138698 173786 138934
rect 174022 138698 174204 138934
rect 173604 103254 174204 138698
rect 173604 103018 173786 103254
rect 174022 103018 174204 103254
rect 173604 102934 174204 103018
rect 173604 102698 173786 102934
rect 174022 102698 174204 102934
rect 173604 67254 174204 102698
rect 173604 67018 173786 67254
rect 174022 67018 174204 67254
rect 173604 66934 174204 67018
rect 173604 66698 173786 66934
rect 174022 66698 174204 66934
rect 173604 31254 174204 66698
rect 173604 31018 173786 31254
rect 174022 31018 174204 31254
rect 173604 30934 174204 31018
rect 173604 30698 173786 30934
rect 174022 30698 174204 30934
rect 155604 -6222 155786 -5986
rect 156022 -6222 156204 -5986
rect 155604 -6306 156204 -6222
rect 155604 -6542 155786 -6306
rect 156022 -6542 156204 -6306
rect 155604 -7504 156204 -6542
rect 173604 -6926 174204 30698
rect 180804 704838 181404 705800
rect 180804 704602 180986 704838
rect 181222 704602 181404 704838
rect 180804 704518 181404 704602
rect 180804 704282 180986 704518
rect 181222 704282 181404 704518
rect 180804 686454 181404 704282
rect 180804 686218 180986 686454
rect 181222 686218 181404 686454
rect 180804 686134 181404 686218
rect 180804 685898 180986 686134
rect 181222 685898 181404 686134
rect 180804 650454 181404 685898
rect 180804 650218 180986 650454
rect 181222 650218 181404 650454
rect 180804 650134 181404 650218
rect 180804 649898 180986 650134
rect 181222 649898 181404 650134
rect 180804 614454 181404 649898
rect 180804 614218 180986 614454
rect 181222 614218 181404 614454
rect 180804 614134 181404 614218
rect 180804 613898 180986 614134
rect 181222 613898 181404 614134
rect 180804 578454 181404 613898
rect 180804 578218 180986 578454
rect 181222 578218 181404 578454
rect 180804 578134 181404 578218
rect 180804 577898 180986 578134
rect 181222 577898 181404 578134
rect 180804 542454 181404 577898
rect 180804 542218 180986 542454
rect 181222 542218 181404 542454
rect 180804 542134 181404 542218
rect 180804 541898 180986 542134
rect 181222 541898 181404 542134
rect 180804 506454 181404 541898
rect 180804 506218 180986 506454
rect 181222 506218 181404 506454
rect 180804 506134 181404 506218
rect 180804 505898 180986 506134
rect 181222 505898 181404 506134
rect 180804 470454 181404 505898
rect 180804 470218 180986 470454
rect 181222 470218 181404 470454
rect 180804 470134 181404 470218
rect 180804 469898 180986 470134
rect 181222 469898 181404 470134
rect 180804 434454 181404 469898
rect 180804 434218 180986 434454
rect 181222 434218 181404 434454
rect 180804 434134 181404 434218
rect 180804 433898 180986 434134
rect 181222 433898 181404 434134
rect 180804 398454 181404 433898
rect 180804 398218 180986 398454
rect 181222 398218 181404 398454
rect 180804 398134 181404 398218
rect 180804 397898 180986 398134
rect 181222 397898 181404 398134
rect 180804 362454 181404 397898
rect 180804 362218 180986 362454
rect 181222 362218 181404 362454
rect 180804 362134 181404 362218
rect 180804 361898 180986 362134
rect 181222 361898 181404 362134
rect 180804 326454 181404 361898
rect 180804 326218 180986 326454
rect 181222 326218 181404 326454
rect 180804 326134 181404 326218
rect 180804 325898 180986 326134
rect 181222 325898 181404 326134
rect 180804 290454 181404 325898
rect 180804 290218 180986 290454
rect 181222 290218 181404 290454
rect 180804 290134 181404 290218
rect 180804 289898 180986 290134
rect 181222 289898 181404 290134
rect 180804 254454 181404 289898
rect 180804 254218 180986 254454
rect 181222 254218 181404 254454
rect 180804 254134 181404 254218
rect 180804 253898 180986 254134
rect 181222 253898 181404 254134
rect 180804 218454 181404 253898
rect 180804 218218 180986 218454
rect 181222 218218 181404 218454
rect 180804 218134 181404 218218
rect 180804 217898 180986 218134
rect 181222 217898 181404 218134
rect 180804 182454 181404 217898
rect 180804 182218 180986 182454
rect 181222 182218 181404 182454
rect 180804 182134 181404 182218
rect 180804 181898 180986 182134
rect 181222 181898 181404 182134
rect 180804 146454 181404 181898
rect 180804 146218 180986 146454
rect 181222 146218 181404 146454
rect 180804 146134 181404 146218
rect 180804 145898 180986 146134
rect 181222 145898 181404 146134
rect 180804 110454 181404 145898
rect 180804 110218 180986 110454
rect 181222 110218 181404 110454
rect 180804 110134 181404 110218
rect 180804 109898 180986 110134
rect 181222 109898 181404 110134
rect 180804 74454 181404 109898
rect 180804 74218 180986 74454
rect 181222 74218 181404 74454
rect 180804 74134 181404 74218
rect 180804 73898 180986 74134
rect 181222 73898 181404 74134
rect 180804 38454 181404 73898
rect 180804 38218 180986 38454
rect 181222 38218 181404 38454
rect 180804 38134 181404 38218
rect 180804 37898 180986 38134
rect 181222 37898 181404 38134
rect 180804 2454 181404 37898
rect 180804 2218 180986 2454
rect 181222 2218 181404 2454
rect 180804 2134 181404 2218
rect 180804 1898 180986 2134
rect 181222 1898 181404 2134
rect 180804 -346 181404 1898
rect 180804 -582 180986 -346
rect 181222 -582 181404 -346
rect 180804 -666 181404 -582
rect 180804 -902 180986 -666
rect 181222 -902 181404 -666
rect 180804 -1864 181404 -902
rect 184404 690054 185004 706162
rect 184404 689818 184586 690054
rect 184822 689818 185004 690054
rect 184404 689734 185004 689818
rect 184404 689498 184586 689734
rect 184822 689498 185004 689734
rect 184404 654054 185004 689498
rect 184404 653818 184586 654054
rect 184822 653818 185004 654054
rect 184404 653734 185004 653818
rect 184404 653498 184586 653734
rect 184822 653498 185004 653734
rect 184404 618054 185004 653498
rect 184404 617818 184586 618054
rect 184822 617818 185004 618054
rect 184404 617734 185004 617818
rect 184404 617498 184586 617734
rect 184822 617498 185004 617734
rect 184404 582054 185004 617498
rect 184404 581818 184586 582054
rect 184822 581818 185004 582054
rect 184404 581734 185004 581818
rect 184404 581498 184586 581734
rect 184822 581498 185004 581734
rect 184404 546054 185004 581498
rect 184404 545818 184586 546054
rect 184822 545818 185004 546054
rect 184404 545734 185004 545818
rect 184404 545498 184586 545734
rect 184822 545498 185004 545734
rect 184404 510054 185004 545498
rect 184404 509818 184586 510054
rect 184822 509818 185004 510054
rect 184404 509734 185004 509818
rect 184404 509498 184586 509734
rect 184822 509498 185004 509734
rect 184404 474054 185004 509498
rect 184404 473818 184586 474054
rect 184822 473818 185004 474054
rect 184404 473734 185004 473818
rect 184404 473498 184586 473734
rect 184822 473498 185004 473734
rect 184404 438054 185004 473498
rect 184404 437818 184586 438054
rect 184822 437818 185004 438054
rect 184404 437734 185004 437818
rect 184404 437498 184586 437734
rect 184822 437498 185004 437734
rect 184404 402054 185004 437498
rect 184404 401818 184586 402054
rect 184822 401818 185004 402054
rect 184404 401734 185004 401818
rect 184404 401498 184586 401734
rect 184822 401498 185004 401734
rect 184404 366054 185004 401498
rect 184404 365818 184586 366054
rect 184822 365818 185004 366054
rect 184404 365734 185004 365818
rect 184404 365498 184586 365734
rect 184822 365498 185004 365734
rect 184404 330054 185004 365498
rect 184404 329818 184586 330054
rect 184822 329818 185004 330054
rect 184404 329734 185004 329818
rect 184404 329498 184586 329734
rect 184822 329498 185004 329734
rect 184404 294054 185004 329498
rect 184404 293818 184586 294054
rect 184822 293818 185004 294054
rect 184404 293734 185004 293818
rect 184404 293498 184586 293734
rect 184822 293498 185004 293734
rect 184404 258054 185004 293498
rect 184404 257818 184586 258054
rect 184822 257818 185004 258054
rect 184404 257734 185004 257818
rect 184404 257498 184586 257734
rect 184822 257498 185004 257734
rect 184404 222054 185004 257498
rect 184404 221818 184586 222054
rect 184822 221818 185004 222054
rect 184404 221734 185004 221818
rect 184404 221498 184586 221734
rect 184822 221498 185004 221734
rect 184404 186054 185004 221498
rect 184404 185818 184586 186054
rect 184822 185818 185004 186054
rect 184404 185734 185004 185818
rect 184404 185498 184586 185734
rect 184822 185498 185004 185734
rect 184404 150054 185004 185498
rect 184404 149818 184586 150054
rect 184822 149818 185004 150054
rect 184404 149734 185004 149818
rect 184404 149498 184586 149734
rect 184822 149498 185004 149734
rect 184404 114054 185004 149498
rect 184404 113818 184586 114054
rect 184822 113818 185004 114054
rect 184404 113734 185004 113818
rect 184404 113498 184586 113734
rect 184822 113498 185004 113734
rect 184404 78054 185004 113498
rect 184404 77818 184586 78054
rect 184822 77818 185004 78054
rect 184404 77734 185004 77818
rect 184404 77498 184586 77734
rect 184822 77498 185004 77734
rect 184404 42054 185004 77498
rect 184404 41818 184586 42054
rect 184822 41818 185004 42054
rect 184404 41734 185004 41818
rect 184404 41498 184586 41734
rect 184822 41498 185004 41734
rect 184404 6054 185004 41498
rect 184404 5818 184586 6054
rect 184822 5818 185004 6054
rect 184404 5734 185004 5818
rect 184404 5498 184586 5734
rect 184822 5498 185004 5734
rect 184404 -2226 185004 5498
rect 184404 -2462 184586 -2226
rect 184822 -2462 185004 -2226
rect 184404 -2546 185004 -2462
rect 184404 -2782 184586 -2546
rect 184822 -2782 185004 -2546
rect 184404 -3744 185004 -2782
rect 188004 693654 188604 708042
rect 188004 693418 188186 693654
rect 188422 693418 188604 693654
rect 188004 693334 188604 693418
rect 188004 693098 188186 693334
rect 188422 693098 188604 693334
rect 188004 657654 188604 693098
rect 188004 657418 188186 657654
rect 188422 657418 188604 657654
rect 188004 657334 188604 657418
rect 188004 657098 188186 657334
rect 188422 657098 188604 657334
rect 188004 621654 188604 657098
rect 188004 621418 188186 621654
rect 188422 621418 188604 621654
rect 188004 621334 188604 621418
rect 188004 621098 188186 621334
rect 188422 621098 188604 621334
rect 188004 585654 188604 621098
rect 188004 585418 188186 585654
rect 188422 585418 188604 585654
rect 188004 585334 188604 585418
rect 188004 585098 188186 585334
rect 188422 585098 188604 585334
rect 188004 549654 188604 585098
rect 188004 549418 188186 549654
rect 188422 549418 188604 549654
rect 188004 549334 188604 549418
rect 188004 549098 188186 549334
rect 188422 549098 188604 549334
rect 188004 513654 188604 549098
rect 188004 513418 188186 513654
rect 188422 513418 188604 513654
rect 188004 513334 188604 513418
rect 188004 513098 188186 513334
rect 188422 513098 188604 513334
rect 188004 477654 188604 513098
rect 188004 477418 188186 477654
rect 188422 477418 188604 477654
rect 188004 477334 188604 477418
rect 188004 477098 188186 477334
rect 188422 477098 188604 477334
rect 188004 441654 188604 477098
rect 188004 441418 188186 441654
rect 188422 441418 188604 441654
rect 188004 441334 188604 441418
rect 188004 441098 188186 441334
rect 188422 441098 188604 441334
rect 188004 405654 188604 441098
rect 188004 405418 188186 405654
rect 188422 405418 188604 405654
rect 188004 405334 188604 405418
rect 188004 405098 188186 405334
rect 188422 405098 188604 405334
rect 188004 369654 188604 405098
rect 188004 369418 188186 369654
rect 188422 369418 188604 369654
rect 188004 369334 188604 369418
rect 188004 369098 188186 369334
rect 188422 369098 188604 369334
rect 188004 333654 188604 369098
rect 188004 333418 188186 333654
rect 188422 333418 188604 333654
rect 188004 333334 188604 333418
rect 188004 333098 188186 333334
rect 188422 333098 188604 333334
rect 188004 297654 188604 333098
rect 188004 297418 188186 297654
rect 188422 297418 188604 297654
rect 188004 297334 188604 297418
rect 188004 297098 188186 297334
rect 188422 297098 188604 297334
rect 188004 261654 188604 297098
rect 188004 261418 188186 261654
rect 188422 261418 188604 261654
rect 188004 261334 188604 261418
rect 188004 261098 188186 261334
rect 188422 261098 188604 261334
rect 188004 225654 188604 261098
rect 188004 225418 188186 225654
rect 188422 225418 188604 225654
rect 188004 225334 188604 225418
rect 188004 225098 188186 225334
rect 188422 225098 188604 225334
rect 188004 189654 188604 225098
rect 188004 189418 188186 189654
rect 188422 189418 188604 189654
rect 188004 189334 188604 189418
rect 188004 189098 188186 189334
rect 188422 189098 188604 189334
rect 188004 153654 188604 189098
rect 188004 153418 188186 153654
rect 188422 153418 188604 153654
rect 188004 153334 188604 153418
rect 188004 153098 188186 153334
rect 188422 153098 188604 153334
rect 188004 117654 188604 153098
rect 188004 117418 188186 117654
rect 188422 117418 188604 117654
rect 188004 117334 188604 117418
rect 188004 117098 188186 117334
rect 188422 117098 188604 117334
rect 188004 81654 188604 117098
rect 188004 81418 188186 81654
rect 188422 81418 188604 81654
rect 188004 81334 188604 81418
rect 188004 81098 188186 81334
rect 188422 81098 188604 81334
rect 188004 45654 188604 81098
rect 188004 45418 188186 45654
rect 188422 45418 188604 45654
rect 188004 45334 188604 45418
rect 188004 45098 188186 45334
rect 188422 45098 188604 45334
rect 188004 9654 188604 45098
rect 188004 9418 188186 9654
rect 188422 9418 188604 9654
rect 188004 9334 188604 9418
rect 188004 9098 188186 9334
rect 188422 9098 188604 9334
rect 188004 -4106 188604 9098
rect 188004 -4342 188186 -4106
rect 188422 -4342 188604 -4106
rect 188004 -4426 188604 -4342
rect 188004 -4662 188186 -4426
rect 188422 -4662 188604 -4426
rect 188004 -5624 188604 -4662
rect 191604 697254 192204 709922
rect 209604 711418 210204 711440
rect 209604 711182 209786 711418
rect 210022 711182 210204 711418
rect 209604 711098 210204 711182
rect 209604 710862 209786 711098
rect 210022 710862 210204 711098
rect 206004 709538 206604 709560
rect 206004 709302 206186 709538
rect 206422 709302 206604 709538
rect 206004 709218 206604 709302
rect 206004 708982 206186 709218
rect 206422 708982 206604 709218
rect 202404 707658 203004 707680
rect 202404 707422 202586 707658
rect 202822 707422 203004 707658
rect 202404 707338 203004 707422
rect 202404 707102 202586 707338
rect 202822 707102 203004 707338
rect 191604 697018 191786 697254
rect 192022 697018 192204 697254
rect 191604 696934 192204 697018
rect 191604 696698 191786 696934
rect 192022 696698 192204 696934
rect 191604 661254 192204 696698
rect 191604 661018 191786 661254
rect 192022 661018 192204 661254
rect 191604 660934 192204 661018
rect 191604 660698 191786 660934
rect 192022 660698 192204 660934
rect 191604 625254 192204 660698
rect 191604 625018 191786 625254
rect 192022 625018 192204 625254
rect 191604 624934 192204 625018
rect 191604 624698 191786 624934
rect 192022 624698 192204 624934
rect 191604 589254 192204 624698
rect 191604 589018 191786 589254
rect 192022 589018 192204 589254
rect 191604 588934 192204 589018
rect 191604 588698 191786 588934
rect 192022 588698 192204 588934
rect 191604 553254 192204 588698
rect 191604 553018 191786 553254
rect 192022 553018 192204 553254
rect 191604 552934 192204 553018
rect 191604 552698 191786 552934
rect 192022 552698 192204 552934
rect 191604 517254 192204 552698
rect 191604 517018 191786 517254
rect 192022 517018 192204 517254
rect 191604 516934 192204 517018
rect 191604 516698 191786 516934
rect 192022 516698 192204 516934
rect 191604 481254 192204 516698
rect 191604 481018 191786 481254
rect 192022 481018 192204 481254
rect 191604 480934 192204 481018
rect 191604 480698 191786 480934
rect 192022 480698 192204 480934
rect 191604 445254 192204 480698
rect 191604 445018 191786 445254
rect 192022 445018 192204 445254
rect 191604 444934 192204 445018
rect 191604 444698 191786 444934
rect 192022 444698 192204 444934
rect 191604 409254 192204 444698
rect 191604 409018 191786 409254
rect 192022 409018 192204 409254
rect 191604 408934 192204 409018
rect 191604 408698 191786 408934
rect 192022 408698 192204 408934
rect 191604 373254 192204 408698
rect 191604 373018 191786 373254
rect 192022 373018 192204 373254
rect 191604 372934 192204 373018
rect 191604 372698 191786 372934
rect 192022 372698 192204 372934
rect 191604 337254 192204 372698
rect 191604 337018 191786 337254
rect 192022 337018 192204 337254
rect 191604 336934 192204 337018
rect 191604 336698 191786 336934
rect 192022 336698 192204 336934
rect 191604 301254 192204 336698
rect 191604 301018 191786 301254
rect 192022 301018 192204 301254
rect 191604 300934 192204 301018
rect 191604 300698 191786 300934
rect 192022 300698 192204 300934
rect 191604 265254 192204 300698
rect 191604 265018 191786 265254
rect 192022 265018 192204 265254
rect 191604 264934 192204 265018
rect 191604 264698 191786 264934
rect 192022 264698 192204 264934
rect 191604 229254 192204 264698
rect 191604 229018 191786 229254
rect 192022 229018 192204 229254
rect 191604 228934 192204 229018
rect 191604 228698 191786 228934
rect 192022 228698 192204 228934
rect 191604 193254 192204 228698
rect 191604 193018 191786 193254
rect 192022 193018 192204 193254
rect 191604 192934 192204 193018
rect 191604 192698 191786 192934
rect 192022 192698 192204 192934
rect 191604 157254 192204 192698
rect 191604 157018 191786 157254
rect 192022 157018 192204 157254
rect 191604 156934 192204 157018
rect 191604 156698 191786 156934
rect 192022 156698 192204 156934
rect 191604 121254 192204 156698
rect 191604 121018 191786 121254
rect 192022 121018 192204 121254
rect 191604 120934 192204 121018
rect 191604 120698 191786 120934
rect 192022 120698 192204 120934
rect 191604 85254 192204 120698
rect 191604 85018 191786 85254
rect 192022 85018 192204 85254
rect 191604 84934 192204 85018
rect 191604 84698 191786 84934
rect 192022 84698 192204 84934
rect 191604 49254 192204 84698
rect 191604 49018 191786 49254
rect 192022 49018 192204 49254
rect 191604 48934 192204 49018
rect 191604 48698 191786 48934
rect 192022 48698 192204 48934
rect 191604 13254 192204 48698
rect 191604 13018 191786 13254
rect 192022 13018 192204 13254
rect 191604 12934 192204 13018
rect 191604 12698 191786 12934
rect 192022 12698 192204 12934
rect 173604 -7162 173786 -6926
rect 174022 -7162 174204 -6926
rect 173604 -7246 174204 -7162
rect 173604 -7482 173786 -7246
rect 174022 -7482 174204 -7246
rect 173604 -7504 174204 -7482
rect 191604 -5986 192204 12698
rect 198804 705778 199404 705800
rect 198804 705542 198986 705778
rect 199222 705542 199404 705778
rect 198804 705458 199404 705542
rect 198804 705222 198986 705458
rect 199222 705222 199404 705458
rect 198804 668454 199404 705222
rect 198804 668218 198986 668454
rect 199222 668218 199404 668454
rect 198804 668134 199404 668218
rect 198804 667898 198986 668134
rect 199222 667898 199404 668134
rect 198804 632454 199404 667898
rect 198804 632218 198986 632454
rect 199222 632218 199404 632454
rect 198804 632134 199404 632218
rect 198804 631898 198986 632134
rect 199222 631898 199404 632134
rect 198804 596454 199404 631898
rect 198804 596218 198986 596454
rect 199222 596218 199404 596454
rect 198804 596134 199404 596218
rect 198804 595898 198986 596134
rect 199222 595898 199404 596134
rect 198804 560454 199404 595898
rect 198804 560218 198986 560454
rect 199222 560218 199404 560454
rect 198804 560134 199404 560218
rect 198804 559898 198986 560134
rect 199222 559898 199404 560134
rect 198804 524454 199404 559898
rect 198804 524218 198986 524454
rect 199222 524218 199404 524454
rect 198804 524134 199404 524218
rect 198804 523898 198986 524134
rect 199222 523898 199404 524134
rect 198804 488454 199404 523898
rect 198804 488218 198986 488454
rect 199222 488218 199404 488454
rect 198804 488134 199404 488218
rect 198804 487898 198986 488134
rect 199222 487898 199404 488134
rect 198804 452454 199404 487898
rect 198804 452218 198986 452454
rect 199222 452218 199404 452454
rect 198804 452134 199404 452218
rect 198804 451898 198986 452134
rect 199222 451898 199404 452134
rect 198804 416454 199404 451898
rect 198804 416218 198986 416454
rect 199222 416218 199404 416454
rect 198804 416134 199404 416218
rect 198804 415898 198986 416134
rect 199222 415898 199404 416134
rect 198804 380454 199404 415898
rect 198804 380218 198986 380454
rect 199222 380218 199404 380454
rect 198804 380134 199404 380218
rect 198804 379898 198986 380134
rect 199222 379898 199404 380134
rect 198804 344454 199404 379898
rect 198804 344218 198986 344454
rect 199222 344218 199404 344454
rect 198804 344134 199404 344218
rect 198804 343898 198986 344134
rect 199222 343898 199404 344134
rect 198804 308454 199404 343898
rect 198804 308218 198986 308454
rect 199222 308218 199404 308454
rect 198804 308134 199404 308218
rect 198804 307898 198986 308134
rect 199222 307898 199404 308134
rect 198804 272454 199404 307898
rect 198804 272218 198986 272454
rect 199222 272218 199404 272454
rect 198804 272134 199404 272218
rect 198804 271898 198986 272134
rect 199222 271898 199404 272134
rect 198804 236454 199404 271898
rect 198804 236218 198986 236454
rect 199222 236218 199404 236454
rect 198804 236134 199404 236218
rect 198804 235898 198986 236134
rect 199222 235898 199404 236134
rect 198804 200454 199404 235898
rect 198804 200218 198986 200454
rect 199222 200218 199404 200454
rect 198804 200134 199404 200218
rect 198804 199898 198986 200134
rect 199222 199898 199404 200134
rect 198804 164454 199404 199898
rect 198804 164218 198986 164454
rect 199222 164218 199404 164454
rect 198804 164134 199404 164218
rect 198804 163898 198986 164134
rect 199222 163898 199404 164134
rect 198804 128454 199404 163898
rect 198804 128218 198986 128454
rect 199222 128218 199404 128454
rect 198804 128134 199404 128218
rect 198804 127898 198986 128134
rect 199222 127898 199404 128134
rect 198804 92454 199404 127898
rect 198804 92218 198986 92454
rect 199222 92218 199404 92454
rect 198804 92134 199404 92218
rect 198804 91898 198986 92134
rect 199222 91898 199404 92134
rect 198804 56454 199404 91898
rect 198804 56218 198986 56454
rect 199222 56218 199404 56454
rect 198804 56134 199404 56218
rect 198804 55898 198986 56134
rect 199222 55898 199404 56134
rect 198804 20454 199404 55898
rect 198804 20218 198986 20454
rect 199222 20218 199404 20454
rect 198804 20134 199404 20218
rect 198804 19898 198986 20134
rect 199222 19898 199404 20134
rect 198804 -1286 199404 19898
rect 198804 -1522 198986 -1286
rect 199222 -1522 199404 -1286
rect 198804 -1606 199404 -1522
rect 198804 -1842 198986 -1606
rect 199222 -1842 199404 -1606
rect 198804 -1864 199404 -1842
rect 202404 672054 203004 707102
rect 202404 671818 202586 672054
rect 202822 671818 203004 672054
rect 202404 671734 203004 671818
rect 202404 671498 202586 671734
rect 202822 671498 203004 671734
rect 202404 636054 203004 671498
rect 202404 635818 202586 636054
rect 202822 635818 203004 636054
rect 202404 635734 203004 635818
rect 202404 635498 202586 635734
rect 202822 635498 203004 635734
rect 202404 600054 203004 635498
rect 202404 599818 202586 600054
rect 202822 599818 203004 600054
rect 202404 599734 203004 599818
rect 202404 599498 202586 599734
rect 202822 599498 203004 599734
rect 202404 564054 203004 599498
rect 202404 563818 202586 564054
rect 202822 563818 203004 564054
rect 202404 563734 203004 563818
rect 202404 563498 202586 563734
rect 202822 563498 203004 563734
rect 202404 528054 203004 563498
rect 202404 527818 202586 528054
rect 202822 527818 203004 528054
rect 202404 527734 203004 527818
rect 202404 527498 202586 527734
rect 202822 527498 203004 527734
rect 202404 492054 203004 527498
rect 202404 491818 202586 492054
rect 202822 491818 203004 492054
rect 202404 491734 203004 491818
rect 202404 491498 202586 491734
rect 202822 491498 203004 491734
rect 202404 456054 203004 491498
rect 202404 455818 202586 456054
rect 202822 455818 203004 456054
rect 202404 455734 203004 455818
rect 202404 455498 202586 455734
rect 202822 455498 203004 455734
rect 202404 420054 203004 455498
rect 202404 419818 202586 420054
rect 202822 419818 203004 420054
rect 202404 419734 203004 419818
rect 202404 419498 202586 419734
rect 202822 419498 203004 419734
rect 202404 384054 203004 419498
rect 202404 383818 202586 384054
rect 202822 383818 203004 384054
rect 202404 383734 203004 383818
rect 202404 383498 202586 383734
rect 202822 383498 203004 383734
rect 202404 348054 203004 383498
rect 202404 347818 202586 348054
rect 202822 347818 203004 348054
rect 202404 347734 203004 347818
rect 202404 347498 202586 347734
rect 202822 347498 203004 347734
rect 202404 312054 203004 347498
rect 202404 311818 202586 312054
rect 202822 311818 203004 312054
rect 202404 311734 203004 311818
rect 202404 311498 202586 311734
rect 202822 311498 203004 311734
rect 202404 276054 203004 311498
rect 202404 275818 202586 276054
rect 202822 275818 203004 276054
rect 202404 275734 203004 275818
rect 202404 275498 202586 275734
rect 202822 275498 203004 275734
rect 202404 240054 203004 275498
rect 202404 239818 202586 240054
rect 202822 239818 203004 240054
rect 202404 239734 203004 239818
rect 202404 239498 202586 239734
rect 202822 239498 203004 239734
rect 202404 204054 203004 239498
rect 202404 203818 202586 204054
rect 202822 203818 203004 204054
rect 202404 203734 203004 203818
rect 202404 203498 202586 203734
rect 202822 203498 203004 203734
rect 202404 168054 203004 203498
rect 202404 167818 202586 168054
rect 202822 167818 203004 168054
rect 202404 167734 203004 167818
rect 202404 167498 202586 167734
rect 202822 167498 203004 167734
rect 202404 132054 203004 167498
rect 202404 131818 202586 132054
rect 202822 131818 203004 132054
rect 202404 131734 203004 131818
rect 202404 131498 202586 131734
rect 202822 131498 203004 131734
rect 202404 96054 203004 131498
rect 202404 95818 202586 96054
rect 202822 95818 203004 96054
rect 202404 95734 203004 95818
rect 202404 95498 202586 95734
rect 202822 95498 203004 95734
rect 202404 60054 203004 95498
rect 202404 59818 202586 60054
rect 202822 59818 203004 60054
rect 202404 59734 203004 59818
rect 202404 59498 202586 59734
rect 202822 59498 203004 59734
rect 202404 24054 203004 59498
rect 202404 23818 202586 24054
rect 202822 23818 203004 24054
rect 202404 23734 203004 23818
rect 202404 23498 202586 23734
rect 202822 23498 203004 23734
rect 202404 -3166 203004 23498
rect 202404 -3402 202586 -3166
rect 202822 -3402 203004 -3166
rect 202404 -3486 203004 -3402
rect 202404 -3722 202586 -3486
rect 202822 -3722 203004 -3486
rect 202404 -3744 203004 -3722
rect 206004 675654 206604 708982
rect 206004 675418 206186 675654
rect 206422 675418 206604 675654
rect 206004 675334 206604 675418
rect 206004 675098 206186 675334
rect 206422 675098 206604 675334
rect 206004 639654 206604 675098
rect 206004 639418 206186 639654
rect 206422 639418 206604 639654
rect 206004 639334 206604 639418
rect 206004 639098 206186 639334
rect 206422 639098 206604 639334
rect 206004 603654 206604 639098
rect 206004 603418 206186 603654
rect 206422 603418 206604 603654
rect 206004 603334 206604 603418
rect 206004 603098 206186 603334
rect 206422 603098 206604 603334
rect 206004 567654 206604 603098
rect 206004 567418 206186 567654
rect 206422 567418 206604 567654
rect 206004 567334 206604 567418
rect 206004 567098 206186 567334
rect 206422 567098 206604 567334
rect 206004 531654 206604 567098
rect 206004 531418 206186 531654
rect 206422 531418 206604 531654
rect 206004 531334 206604 531418
rect 206004 531098 206186 531334
rect 206422 531098 206604 531334
rect 206004 495654 206604 531098
rect 206004 495418 206186 495654
rect 206422 495418 206604 495654
rect 206004 495334 206604 495418
rect 206004 495098 206186 495334
rect 206422 495098 206604 495334
rect 206004 459654 206604 495098
rect 206004 459418 206186 459654
rect 206422 459418 206604 459654
rect 206004 459334 206604 459418
rect 206004 459098 206186 459334
rect 206422 459098 206604 459334
rect 206004 423654 206604 459098
rect 206004 423418 206186 423654
rect 206422 423418 206604 423654
rect 206004 423334 206604 423418
rect 206004 423098 206186 423334
rect 206422 423098 206604 423334
rect 206004 387654 206604 423098
rect 206004 387418 206186 387654
rect 206422 387418 206604 387654
rect 206004 387334 206604 387418
rect 206004 387098 206186 387334
rect 206422 387098 206604 387334
rect 206004 351654 206604 387098
rect 206004 351418 206186 351654
rect 206422 351418 206604 351654
rect 206004 351334 206604 351418
rect 206004 351098 206186 351334
rect 206422 351098 206604 351334
rect 206004 315654 206604 351098
rect 206004 315418 206186 315654
rect 206422 315418 206604 315654
rect 206004 315334 206604 315418
rect 206004 315098 206186 315334
rect 206422 315098 206604 315334
rect 206004 279654 206604 315098
rect 206004 279418 206186 279654
rect 206422 279418 206604 279654
rect 206004 279334 206604 279418
rect 206004 279098 206186 279334
rect 206422 279098 206604 279334
rect 206004 243654 206604 279098
rect 206004 243418 206186 243654
rect 206422 243418 206604 243654
rect 206004 243334 206604 243418
rect 206004 243098 206186 243334
rect 206422 243098 206604 243334
rect 206004 207654 206604 243098
rect 206004 207418 206186 207654
rect 206422 207418 206604 207654
rect 206004 207334 206604 207418
rect 206004 207098 206186 207334
rect 206422 207098 206604 207334
rect 206004 171654 206604 207098
rect 206004 171418 206186 171654
rect 206422 171418 206604 171654
rect 206004 171334 206604 171418
rect 206004 171098 206186 171334
rect 206422 171098 206604 171334
rect 206004 135654 206604 171098
rect 206004 135418 206186 135654
rect 206422 135418 206604 135654
rect 206004 135334 206604 135418
rect 206004 135098 206186 135334
rect 206422 135098 206604 135334
rect 206004 99654 206604 135098
rect 206004 99418 206186 99654
rect 206422 99418 206604 99654
rect 206004 99334 206604 99418
rect 206004 99098 206186 99334
rect 206422 99098 206604 99334
rect 206004 63654 206604 99098
rect 206004 63418 206186 63654
rect 206422 63418 206604 63654
rect 206004 63334 206604 63418
rect 206004 63098 206186 63334
rect 206422 63098 206604 63334
rect 206004 27654 206604 63098
rect 206004 27418 206186 27654
rect 206422 27418 206604 27654
rect 206004 27334 206604 27418
rect 206004 27098 206186 27334
rect 206422 27098 206604 27334
rect 206004 -5046 206604 27098
rect 206004 -5282 206186 -5046
rect 206422 -5282 206604 -5046
rect 206004 -5366 206604 -5282
rect 206004 -5602 206186 -5366
rect 206422 -5602 206604 -5366
rect 206004 -5624 206604 -5602
rect 209604 679254 210204 710862
rect 227604 710478 228204 711440
rect 227604 710242 227786 710478
rect 228022 710242 228204 710478
rect 227604 710158 228204 710242
rect 227604 709922 227786 710158
rect 228022 709922 228204 710158
rect 224004 708598 224604 709560
rect 224004 708362 224186 708598
rect 224422 708362 224604 708598
rect 224004 708278 224604 708362
rect 224004 708042 224186 708278
rect 224422 708042 224604 708278
rect 220404 706718 221004 707680
rect 220404 706482 220586 706718
rect 220822 706482 221004 706718
rect 220404 706398 221004 706482
rect 220404 706162 220586 706398
rect 220822 706162 221004 706398
rect 209604 679018 209786 679254
rect 210022 679018 210204 679254
rect 209604 678934 210204 679018
rect 209604 678698 209786 678934
rect 210022 678698 210204 678934
rect 209604 643254 210204 678698
rect 209604 643018 209786 643254
rect 210022 643018 210204 643254
rect 209604 642934 210204 643018
rect 209604 642698 209786 642934
rect 210022 642698 210204 642934
rect 209604 607254 210204 642698
rect 209604 607018 209786 607254
rect 210022 607018 210204 607254
rect 209604 606934 210204 607018
rect 209604 606698 209786 606934
rect 210022 606698 210204 606934
rect 209604 571254 210204 606698
rect 209604 571018 209786 571254
rect 210022 571018 210204 571254
rect 209604 570934 210204 571018
rect 209604 570698 209786 570934
rect 210022 570698 210204 570934
rect 209604 535254 210204 570698
rect 209604 535018 209786 535254
rect 210022 535018 210204 535254
rect 209604 534934 210204 535018
rect 209604 534698 209786 534934
rect 210022 534698 210204 534934
rect 209604 499254 210204 534698
rect 209604 499018 209786 499254
rect 210022 499018 210204 499254
rect 209604 498934 210204 499018
rect 209604 498698 209786 498934
rect 210022 498698 210204 498934
rect 209604 463254 210204 498698
rect 209604 463018 209786 463254
rect 210022 463018 210204 463254
rect 209604 462934 210204 463018
rect 209604 462698 209786 462934
rect 210022 462698 210204 462934
rect 209604 427254 210204 462698
rect 209604 427018 209786 427254
rect 210022 427018 210204 427254
rect 209604 426934 210204 427018
rect 209604 426698 209786 426934
rect 210022 426698 210204 426934
rect 209604 391254 210204 426698
rect 209604 391018 209786 391254
rect 210022 391018 210204 391254
rect 209604 390934 210204 391018
rect 209604 390698 209786 390934
rect 210022 390698 210204 390934
rect 209604 355254 210204 390698
rect 209604 355018 209786 355254
rect 210022 355018 210204 355254
rect 209604 354934 210204 355018
rect 209604 354698 209786 354934
rect 210022 354698 210204 354934
rect 209604 319254 210204 354698
rect 209604 319018 209786 319254
rect 210022 319018 210204 319254
rect 209604 318934 210204 319018
rect 209604 318698 209786 318934
rect 210022 318698 210204 318934
rect 209604 283254 210204 318698
rect 209604 283018 209786 283254
rect 210022 283018 210204 283254
rect 209604 282934 210204 283018
rect 209604 282698 209786 282934
rect 210022 282698 210204 282934
rect 209604 247254 210204 282698
rect 209604 247018 209786 247254
rect 210022 247018 210204 247254
rect 209604 246934 210204 247018
rect 209604 246698 209786 246934
rect 210022 246698 210204 246934
rect 209604 211254 210204 246698
rect 209604 211018 209786 211254
rect 210022 211018 210204 211254
rect 209604 210934 210204 211018
rect 209604 210698 209786 210934
rect 210022 210698 210204 210934
rect 209604 175254 210204 210698
rect 209604 175018 209786 175254
rect 210022 175018 210204 175254
rect 209604 174934 210204 175018
rect 209604 174698 209786 174934
rect 210022 174698 210204 174934
rect 209604 139254 210204 174698
rect 209604 139018 209786 139254
rect 210022 139018 210204 139254
rect 209604 138934 210204 139018
rect 209604 138698 209786 138934
rect 210022 138698 210204 138934
rect 209604 103254 210204 138698
rect 209604 103018 209786 103254
rect 210022 103018 210204 103254
rect 209604 102934 210204 103018
rect 209604 102698 209786 102934
rect 210022 102698 210204 102934
rect 209604 67254 210204 102698
rect 209604 67018 209786 67254
rect 210022 67018 210204 67254
rect 209604 66934 210204 67018
rect 209604 66698 209786 66934
rect 210022 66698 210204 66934
rect 209604 31254 210204 66698
rect 209604 31018 209786 31254
rect 210022 31018 210204 31254
rect 209604 30934 210204 31018
rect 209604 30698 209786 30934
rect 210022 30698 210204 30934
rect 191604 -6222 191786 -5986
rect 192022 -6222 192204 -5986
rect 191604 -6306 192204 -6222
rect 191604 -6542 191786 -6306
rect 192022 -6542 192204 -6306
rect 191604 -7504 192204 -6542
rect 209604 -6926 210204 30698
rect 216804 704838 217404 705800
rect 216804 704602 216986 704838
rect 217222 704602 217404 704838
rect 216804 704518 217404 704602
rect 216804 704282 216986 704518
rect 217222 704282 217404 704518
rect 216804 686454 217404 704282
rect 216804 686218 216986 686454
rect 217222 686218 217404 686454
rect 216804 686134 217404 686218
rect 216804 685898 216986 686134
rect 217222 685898 217404 686134
rect 216804 650454 217404 685898
rect 216804 650218 216986 650454
rect 217222 650218 217404 650454
rect 216804 650134 217404 650218
rect 216804 649898 216986 650134
rect 217222 649898 217404 650134
rect 216804 614454 217404 649898
rect 216804 614218 216986 614454
rect 217222 614218 217404 614454
rect 216804 614134 217404 614218
rect 216804 613898 216986 614134
rect 217222 613898 217404 614134
rect 216804 578454 217404 613898
rect 216804 578218 216986 578454
rect 217222 578218 217404 578454
rect 216804 578134 217404 578218
rect 216804 577898 216986 578134
rect 217222 577898 217404 578134
rect 216804 542454 217404 577898
rect 216804 542218 216986 542454
rect 217222 542218 217404 542454
rect 216804 542134 217404 542218
rect 216804 541898 216986 542134
rect 217222 541898 217404 542134
rect 216804 506454 217404 541898
rect 216804 506218 216986 506454
rect 217222 506218 217404 506454
rect 216804 506134 217404 506218
rect 216804 505898 216986 506134
rect 217222 505898 217404 506134
rect 216804 470454 217404 505898
rect 216804 470218 216986 470454
rect 217222 470218 217404 470454
rect 216804 470134 217404 470218
rect 216804 469898 216986 470134
rect 217222 469898 217404 470134
rect 216804 434454 217404 469898
rect 216804 434218 216986 434454
rect 217222 434218 217404 434454
rect 216804 434134 217404 434218
rect 216804 433898 216986 434134
rect 217222 433898 217404 434134
rect 216804 398454 217404 433898
rect 216804 398218 216986 398454
rect 217222 398218 217404 398454
rect 216804 398134 217404 398218
rect 216804 397898 216986 398134
rect 217222 397898 217404 398134
rect 216804 362454 217404 397898
rect 216804 362218 216986 362454
rect 217222 362218 217404 362454
rect 216804 362134 217404 362218
rect 216804 361898 216986 362134
rect 217222 361898 217404 362134
rect 216804 326454 217404 361898
rect 216804 326218 216986 326454
rect 217222 326218 217404 326454
rect 216804 326134 217404 326218
rect 216804 325898 216986 326134
rect 217222 325898 217404 326134
rect 216804 290454 217404 325898
rect 216804 290218 216986 290454
rect 217222 290218 217404 290454
rect 216804 290134 217404 290218
rect 216804 289898 216986 290134
rect 217222 289898 217404 290134
rect 216804 254454 217404 289898
rect 216804 254218 216986 254454
rect 217222 254218 217404 254454
rect 216804 254134 217404 254218
rect 216804 253898 216986 254134
rect 217222 253898 217404 254134
rect 216804 218454 217404 253898
rect 216804 218218 216986 218454
rect 217222 218218 217404 218454
rect 216804 218134 217404 218218
rect 216804 217898 216986 218134
rect 217222 217898 217404 218134
rect 216804 182454 217404 217898
rect 216804 182218 216986 182454
rect 217222 182218 217404 182454
rect 216804 182134 217404 182218
rect 216804 181898 216986 182134
rect 217222 181898 217404 182134
rect 216804 146454 217404 181898
rect 216804 146218 216986 146454
rect 217222 146218 217404 146454
rect 216804 146134 217404 146218
rect 216804 145898 216986 146134
rect 217222 145898 217404 146134
rect 216804 110454 217404 145898
rect 216804 110218 216986 110454
rect 217222 110218 217404 110454
rect 216804 110134 217404 110218
rect 216804 109898 216986 110134
rect 217222 109898 217404 110134
rect 216804 74454 217404 109898
rect 216804 74218 216986 74454
rect 217222 74218 217404 74454
rect 216804 74134 217404 74218
rect 216804 73898 216986 74134
rect 217222 73898 217404 74134
rect 216804 38454 217404 73898
rect 216804 38218 216986 38454
rect 217222 38218 217404 38454
rect 216804 38134 217404 38218
rect 216804 37898 216986 38134
rect 217222 37898 217404 38134
rect 216804 2454 217404 37898
rect 216804 2218 216986 2454
rect 217222 2218 217404 2454
rect 216804 2134 217404 2218
rect 216804 1898 216986 2134
rect 217222 1898 217404 2134
rect 216804 -346 217404 1898
rect 216804 -582 216986 -346
rect 217222 -582 217404 -346
rect 216804 -666 217404 -582
rect 216804 -902 216986 -666
rect 217222 -902 217404 -666
rect 216804 -1864 217404 -902
rect 220404 690054 221004 706162
rect 220404 689818 220586 690054
rect 220822 689818 221004 690054
rect 220404 689734 221004 689818
rect 220404 689498 220586 689734
rect 220822 689498 221004 689734
rect 220404 654054 221004 689498
rect 220404 653818 220586 654054
rect 220822 653818 221004 654054
rect 220404 653734 221004 653818
rect 220404 653498 220586 653734
rect 220822 653498 221004 653734
rect 220404 618054 221004 653498
rect 220404 617818 220586 618054
rect 220822 617818 221004 618054
rect 220404 617734 221004 617818
rect 220404 617498 220586 617734
rect 220822 617498 221004 617734
rect 220404 582054 221004 617498
rect 220404 581818 220586 582054
rect 220822 581818 221004 582054
rect 220404 581734 221004 581818
rect 220404 581498 220586 581734
rect 220822 581498 221004 581734
rect 220404 546054 221004 581498
rect 220404 545818 220586 546054
rect 220822 545818 221004 546054
rect 220404 545734 221004 545818
rect 220404 545498 220586 545734
rect 220822 545498 221004 545734
rect 220404 510054 221004 545498
rect 220404 509818 220586 510054
rect 220822 509818 221004 510054
rect 220404 509734 221004 509818
rect 220404 509498 220586 509734
rect 220822 509498 221004 509734
rect 220404 474054 221004 509498
rect 220404 473818 220586 474054
rect 220822 473818 221004 474054
rect 220404 473734 221004 473818
rect 220404 473498 220586 473734
rect 220822 473498 221004 473734
rect 220404 438054 221004 473498
rect 220404 437818 220586 438054
rect 220822 437818 221004 438054
rect 220404 437734 221004 437818
rect 220404 437498 220586 437734
rect 220822 437498 221004 437734
rect 220404 402054 221004 437498
rect 220404 401818 220586 402054
rect 220822 401818 221004 402054
rect 220404 401734 221004 401818
rect 220404 401498 220586 401734
rect 220822 401498 221004 401734
rect 220404 366054 221004 401498
rect 220404 365818 220586 366054
rect 220822 365818 221004 366054
rect 220404 365734 221004 365818
rect 220404 365498 220586 365734
rect 220822 365498 221004 365734
rect 220404 330054 221004 365498
rect 220404 329818 220586 330054
rect 220822 329818 221004 330054
rect 220404 329734 221004 329818
rect 220404 329498 220586 329734
rect 220822 329498 221004 329734
rect 220404 294054 221004 329498
rect 220404 293818 220586 294054
rect 220822 293818 221004 294054
rect 220404 293734 221004 293818
rect 220404 293498 220586 293734
rect 220822 293498 221004 293734
rect 220404 258054 221004 293498
rect 220404 257818 220586 258054
rect 220822 257818 221004 258054
rect 220404 257734 221004 257818
rect 220404 257498 220586 257734
rect 220822 257498 221004 257734
rect 220404 222054 221004 257498
rect 220404 221818 220586 222054
rect 220822 221818 221004 222054
rect 220404 221734 221004 221818
rect 220404 221498 220586 221734
rect 220822 221498 221004 221734
rect 220404 186054 221004 221498
rect 220404 185818 220586 186054
rect 220822 185818 221004 186054
rect 220404 185734 221004 185818
rect 220404 185498 220586 185734
rect 220822 185498 221004 185734
rect 220404 150054 221004 185498
rect 220404 149818 220586 150054
rect 220822 149818 221004 150054
rect 220404 149734 221004 149818
rect 220404 149498 220586 149734
rect 220822 149498 221004 149734
rect 220404 114054 221004 149498
rect 220404 113818 220586 114054
rect 220822 113818 221004 114054
rect 220404 113734 221004 113818
rect 220404 113498 220586 113734
rect 220822 113498 221004 113734
rect 220404 78054 221004 113498
rect 220404 77818 220586 78054
rect 220822 77818 221004 78054
rect 220404 77734 221004 77818
rect 220404 77498 220586 77734
rect 220822 77498 221004 77734
rect 220404 42054 221004 77498
rect 220404 41818 220586 42054
rect 220822 41818 221004 42054
rect 220404 41734 221004 41818
rect 220404 41498 220586 41734
rect 220822 41498 221004 41734
rect 220404 6054 221004 41498
rect 220404 5818 220586 6054
rect 220822 5818 221004 6054
rect 220404 5734 221004 5818
rect 220404 5498 220586 5734
rect 220822 5498 221004 5734
rect 220404 -2226 221004 5498
rect 220404 -2462 220586 -2226
rect 220822 -2462 221004 -2226
rect 220404 -2546 221004 -2462
rect 220404 -2782 220586 -2546
rect 220822 -2782 221004 -2546
rect 220404 -3744 221004 -2782
rect 224004 693654 224604 708042
rect 224004 693418 224186 693654
rect 224422 693418 224604 693654
rect 224004 693334 224604 693418
rect 224004 693098 224186 693334
rect 224422 693098 224604 693334
rect 224004 657654 224604 693098
rect 224004 657418 224186 657654
rect 224422 657418 224604 657654
rect 224004 657334 224604 657418
rect 224004 657098 224186 657334
rect 224422 657098 224604 657334
rect 224004 621654 224604 657098
rect 224004 621418 224186 621654
rect 224422 621418 224604 621654
rect 224004 621334 224604 621418
rect 224004 621098 224186 621334
rect 224422 621098 224604 621334
rect 224004 585654 224604 621098
rect 224004 585418 224186 585654
rect 224422 585418 224604 585654
rect 224004 585334 224604 585418
rect 224004 585098 224186 585334
rect 224422 585098 224604 585334
rect 224004 549654 224604 585098
rect 224004 549418 224186 549654
rect 224422 549418 224604 549654
rect 224004 549334 224604 549418
rect 224004 549098 224186 549334
rect 224422 549098 224604 549334
rect 224004 513654 224604 549098
rect 224004 513418 224186 513654
rect 224422 513418 224604 513654
rect 224004 513334 224604 513418
rect 224004 513098 224186 513334
rect 224422 513098 224604 513334
rect 224004 477654 224604 513098
rect 224004 477418 224186 477654
rect 224422 477418 224604 477654
rect 224004 477334 224604 477418
rect 224004 477098 224186 477334
rect 224422 477098 224604 477334
rect 224004 441654 224604 477098
rect 224004 441418 224186 441654
rect 224422 441418 224604 441654
rect 224004 441334 224604 441418
rect 224004 441098 224186 441334
rect 224422 441098 224604 441334
rect 224004 405654 224604 441098
rect 224004 405418 224186 405654
rect 224422 405418 224604 405654
rect 224004 405334 224604 405418
rect 224004 405098 224186 405334
rect 224422 405098 224604 405334
rect 224004 369654 224604 405098
rect 224004 369418 224186 369654
rect 224422 369418 224604 369654
rect 224004 369334 224604 369418
rect 224004 369098 224186 369334
rect 224422 369098 224604 369334
rect 224004 333654 224604 369098
rect 224004 333418 224186 333654
rect 224422 333418 224604 333654
rect 224004 333334 224604 333418
rect 224004 333098 224186 333334
rect 224422 333098 224604 333334
rect 224004 297654 224604 333098
rect 224004 297418 224186 297654
rect 224422 297418 224604 297654
rect 224004 297334 224604 297418
rect 224004 297098 224186 297334
rect 224422 297098 224604 297334
rect 224004 261654 224604 297098
rect 224004 261418 224186 261654
rect 224422 261418 224604 261654
rect 224004 261334 224604 261418
rect 224004 261098 224186 261334
rect 224422 261098 224604 261334
rect 224004 225654 224604 261098
rect 224004 225418 224186 225654
rect 224422 225418 224604 225654
rect 224004 225334 224604 225418
rect 224004 225098 224186 225334
rect 224422 225098 224604 225334
rect 224004 189654 224604 225098
rect 224004 189418 224186 189654
rect 224422 189418 224604 189654
rect 224004 189334 224604 189418
rect 224004 189098 224186 189334
rect 224422 189098 224604 189334
rect 224004 153654 224604 189098
rect 224004 153418 224186 153654
rect 224422 153418 224604 153654
rect 224004 153334 224604 153418
rect 224004 153098 224186 153334
rect 224422 153098 224604 153334
rect 224004 117654 224604 153098
rect 224004 117418 224186 117654
rect 224422 117418 224604 117654
rect 224004 117334 224604 117418
rect 224004 117098 224186 117334
rect 224422 117098 224604 117334
rect 224004 81654 224604 117098
rect 224004 81418 224186 81654
rect 224422 81418 224604 81654
rect 224004 81334 224604 81418
rect 224004 81098 224186 81334
rect 224422 81098 224604 81334
rect 224004 45654 224604 81098
rect 224004 45418 224186 45654
rect 224422 45418 224604 45654
rect 224004 45334 224604 45418
rect 224004 45098 224186 45334
rect 224422 45098 224604 45334
rect 224004 9654 224604 45098
rect 224004 9418 224186 9654
rect 224422 9418 224604 9654
rect 224004 9334 224604 9418
rect 224004 9098 224186 9334
rect 224422 9098 224604 9334
rect 224004 -4106 224604 9098
rect 224004 -4342 224186 -4106
rect 224422 -4342 224604 -4106
rect 224004 -4426 224604 -4342
rect 224004 -4662 224186 -4426
rect 224422 -4662 224604 -4426
rect 224004 -5624 224604 -4662
rect 227604 697254 228204 709922
rect 245604 711418 246204 711440
rect 245604 711182 245786 711418
rect 246022 711182 246204 711418
rect 245604 711098 246204 711182
rect 245604 710862 245786 711098
rect 246022 710862 246204 711098
rect 242004 709538 242604 709560
rect 242004 709302 242186 709538
rect 242422 709302 242604 709538
rect 242004 709218 242604 709302
rect 242004 708982 242186 709218
rect 242422 708982 242604 709218
rect 238404 707658 239004 707680
rect 238404 707422 238586 707658
rect 238822 707422 239004 707658
rect 238404 707338 239004 707422
rect 238404 707102 238586 707338
rect 238822 707102 239004 707338
rect 227604 697018 227786 697254
rect 228022 697018 228204 697254
rect 227604 696934 228204 697018
rect 227604 696698 227786 696934
rect 228022 696698 228204 696934
rect 227604 661254 228204 696698
rect 227604 661018 227786 661254
rect 228022 661018 228204 661254
rect 227604 660934 228204 661018
rect 227604 660698 227786 660934
rect 228022 660698 228204 660934
rect 227604 625254 228204 660698
rect 227604 625018 227786 625254
rect 228022 625018 228204 625254
rect 227604 624934 228204 625018
rect 227604 624698 227786 624934
rect 228022 624698 228204 624934
rect 227604 589254 228204 624698
rect 227604 589018 227786 589254
rect 228022 589018 228204 589254
rect 227604 588934 228204 589018
rect 227604 588698 227786 588934
rect 228022 588698 228204 588934
rect 227604 553254 228204 588698
rect 227604 553018 227786 553254
rect 228022 553018 228204 553254
rect 227604 552934 228204 553018
rect 227604 552698 227786 552934
rect 228022 552698 228204 552934
rect 227604 517254 228204 552698
rect 227604 517018 227786 517254
rect 228022 517018 228204 517254
rect 227604 516934 228204 517018
rect 227604 516698 227786 516934
rect 228022 516698 228204 516934
rect 227604 481254 228204 516698
rect 227604 481018 227786 481254
rect 228022 481018 228204 481254
rect 227604 480934 228204 481018
rect 227604 480698 227786 480934
rect 228022 480698 228204 480934
rect 227604 445254 228204 480698
rect 227604 445018 227786 445254
rect 228022 445018 228204 445254
rect 227604 444934 228204 445018
rect 227604 444698 227786 444934
rect 228022 444698 228204 444934
rect 227604 409254 228204 444698
rect 227604 409018 227786 409254
rect 228022 409018 228204 409254
rect 227604 408934 228204 409018
rect 227604 408698 227786 408934
rect 228022 408698 228204 408934
rect 227604 373254 228204 408698
rect 227604 373018 227786 373254
rect 228022 373018 228204 373254
rect 227604 372934 228204 373018
rect 227604 372698 227786 372934
rect 228022 372698 228204 372934
rect 227604 337254 228204 372698
rect 227604 337018 227786 337254
rect 228022 337018 228204 337254
rect 227604 336934 228204 337018
rect 227604 336698 227786 336934
rect 228022 336698 228204 336934
rect 227604 301254 228204 336698
rect 227604 301018 227786 301254
rect 228022 301018 228204 301254
rect 227604 300934 228204 301018
rect 227604 300698 227786 300934
rect 228022 300698 228204 300934
rect 227604 265254 228204 300698
rect 227604 265018 227786 265254
rect 228022 265018 228204 265254
rect 227604 264934 228204 265018
rect 227604 264698 227786 264934
rect 228022 264698 228204 264934
rect 227604 229254 228204 264698
rect 227604 229018 227786 229254
rect 228022 229018 228204 229254
rect 227604 228934 228204 229018
rect 227604 228698 227786 228934
rect 228022 228698 228204 228934
rect 227604 193254 228204 228698
rect 227604 193018 227786 193254
rect 228022 193018 228204 193254
rect 227604 192934 228204 193018
rect 227604 192698 227786 192934
rect 228022 192698 228204 192934
rect 227604 157254 228204 192698
rect 227604 157018 227786 157254
rect 228022 157018 228204 157254
rect 227604 156934 228204 157018
rect 227604 156698 227786 156934
rect 228022 156698 228204 156934
rect 227604 121254 228204 156698
rect 227604 121018 227786 121254
rect 228022 121018 228204 121254
rect 227604 120934 228204 121018
rect 227604 120698 227786 120934
rect 228022 120698 228204 120934
rect 227604 85254 228204 120698
rect 227604 85018 227786 85254
rect 228022 85018 228204 85254
rect 227604 84934 228204 85018
rect 227604 84698 227786 84934
rect 228022 84698 228204 84934
rect 227604 49254 228204 84698
rect 227604 49018 227786 49254
rect 228022 49018 228204 49254
rect 227604 48934 228204 49018
rect 227604 48698 227786 48934
rect 228022 48698 228204 48934
rect 227604 13254 228204 48698
rect 227604 13018 227786 13254
rect 228022 13018 228204 13254
rect 227604 12934 228204 13018
rect 227604 12698 227786 12934
rect 228022 12698 228204 12934
rect 209604 -7162 209786 -6926
rect 210022 -7162 210204 -6926
rect 209604 -7246 210204 -7162
rect 209604 -7482 209786 -7246
rect 210022 -7482 210204 -7246
rect 209604 -7504 210204 -7482
rect 227604 -5986 228204 12698
rect 234804 705778 235404 705800
rect 234804 705542 234986 705778
rect 235222 705542 235404 705778
rect 234804 705458 235404 705542
rect 234804 705222 234986 705458
rect 235222 705222 235404 705458
rect 234804 668454 235404 705222
rect 234804 668218 234986 668454
rect 235222 668218 235404 668454
rect 234804 668134 235404 668218
rect 234804 667898 234986 668134
rect 235222 667898 235404 668134
rect 234804 632454 235404 667898
rect 234804 632218 234986 632454
rect 235222 632218 235404 632454
rect 234804 632134 235404 632218
rect 234804 631898 234986 632134
rect 235222 631898 235404 632134
rect 234804 596454 235404 631898
rect 234804 596218 234986 596454
rect 235222 596218 235404 596454
rect 234804 596134 235404 596218
rect 234804 595898 234986 596134
rect 235222 595898 235404 596134
rect 234804 560454 235404 595898
rect 234804 560218 234986 560454
rect 235222 560218 235404 560454
rect 234804 560134 235404 560218
rect 234804 559898 234986 560134
rect 235222 559898 235404 560134
rect 234804 524454 235404 559898
rect 234804 524218 234986 524454
rect 235222 524218 235404 524454
rect 234804 524134 235404 524218
rect 234804 523898 234986 524134
rect 235222 523898 235404 524134
rect 234804 488454 235404 523898
rect 234804 488218 234986 488454
rect 235222 488218 235404 488454
rect 234804 488134 235404 488218
rect 234804 487898 234986 488134
rect 235222 487898 235404 488134
rect 234804 452454 235404 487898
rect 234804 452218 234986 452454
rect 235222 452218 235404 452454
rect 234804 452134 235404 452218
rect 234804 451898 234986 452134
rect 235222 451898 235404 452134
rect 234804 416454 235404 451898
rect 234804 416218 234986 416454
rect 235222 416218 235404 416454
rect 234804 416134 235404 416218
rect 234804 415898 234986 416134
rect 235222 415898 235404 416134
rect 234804 380454 235404 415898
rect 234804 380218 234986 380454
rect 235222 380218 235404 380454
rect 234804 380134 235404 380218
rect 234804 379898 234986 380134
rect 235222 379898 235404 380134
rect 234804 344454 235404 379898
rect 234804 344218 234986 344454
rect 235222 344218 235404 344454
rect 234804 344134 235404 344218
rect 234804 343898 234986 344134
rect 235222 343898 235404 344134
rect 234804 308454 235404 343898
rect 234804 308218 234986 308454
rect 235222 308218 235404 308454
rect 234804 308134 235404 308218
rect 234804 307898 234986 308134
rect 235222 307898 235404 308134
rect 234804 272454 235404 307898
rect 234804 272218 234986 272454
rect 235222 272218 235404 272454
rect 234804 272134 235404 272218
rect 234804 271898 234986 272134
rect 235222 271898 235404 272134
rect 234804 236454 235404 271898
rect 234804 236218 234986 236454
rect 235222 236218 235404 236454
rect 234804 236134 235404 236218
rect 234804 235898 234986 236134
rect 235222 235898 235404 236134
rect 234804 200454 235404 235898
rect 234804 200218 234986 200454
rect 235222 200218 235404 200454
rect 234804 200134 235404 200218
rect 234804 199898 234986 200134
rect 235222 199898 235404 200134
rect 234804 164454 235404 199898
rect 234804 164218 234986 164454
rect 235222 164218 235404 164454
rect 234804 164134 235404 164218
rect 234804 163898 234986 164134
rect 235222 163898 235404 164134
rect 234804 128454 235404 163898
rect 234804 128218 234986 128454
rect 235222 128218 235404 128454
rect 234804 128134 235404 128218
rect 234804 127898 234986 128134
rect 235222 127898 235404 128134
rect 234804 92454 235404 127898
rect 234804 92218 234986 92454
rect 235222 92218 235404 92454
rect 234804 92134 235404 92218
rect 234804 91898 234986 92134
rect 235222 91898 235404 92134
rect 234804 56454 235404 91898
rect 234804 56218 234986 56454
rect 235222 56218 235404 56454
rect 234804 56134 235404 56218
rect 234804 55898 234986 56134
rect 235222 55898 235404 56134
rect 234804 20454 235404 55898
rect 234804 20218 234986 20454
rect 235222 20218 235404 20454
rect 234804 20134 235404 20218
rect 234804 19898 234986 20134
rect 235222 19898 235404 20134
rect 234804 -1286 235404 19898
rect 234804 -1522 234986 -1286
rect 235222 -1522 235404 -1286
rect 234804 -1606 235404 -1522
rect 234804 -1842 234986 -1606
rect 235222 -1842 235404 -1606
rect 234804 -1864 235404 -1842
rect 238404 672054 239004 707102
rect 238404 671818 238586 672054
rect 238822 671818 239004 672054
rect 238404 671734 239004 671818
rect 238404 671498 238586 671734
rect 238822 671498 239004 671734
rect 238404 636054 239004 671498
rect 238404 635818 238586 636054
rect 238822 635818 239004 636054
rect 238404 635734 239004 635818
rect 238404 635498 238586 635734
rect 238822 635498 239004 635734
rect 238404 600054 239004 635498
rect 238404 599818 238586 600054
rect 238822 599818 239004 600054
rect 238404 599734 239004 599818
rect 238404 599498 238586 599734
rect 238822 599498 239004 599734
rect 238404 564054 239004 599498
rect 238404 563818 238586 564054
rect 238822 563818 239004 564054
rect 238404 563734 239004 563818
rect 238404 563498 238586 563734
rect 238822 563498 239004 563734
rect 238404 528054 239004 563498
rect 238404 527818 238586 528054
rect 238822 527818 239004 528054
rect 238404 527734 239004 527818
rect 238404 527498 238586 527734
rect 238822 527498 239004 527734
rect 238404 492054 239004 527498
rect 238404 491818 238586 492054
rect 238822 491818 239004 492054
rect 238404 491734 239004 491818
rect 238404 491498 238586 491734
rect 238822 491498 239004 491734
rect 238404 456054 239004 491498
rect 238404 455818 238586 456054
rect 238822 455818 239004 456054
rect 238404 455734 239004 455818
rect 238404 455498 238586 455734
rect 238822 455498 239004 455734
rect 238404 420054 239004 455498
rect 238404 419818 238586 420054
rect 238822 419818 239004 420054
rect 238404 419734 239004 419818
rect 238404 419498 238586 419734
rect 238822 419498 239004 419734
rect 238404 384054 239004 419498
rect 238404 383818 238586 384054
rect 238822 383818 239004 384054
rect 238404 383734 239004 383818
rect 238404 383498 238586 383734
rect 238822 383498 239004 383734
rect 238404 348054 239004 383498
rect 238404 347818 238586 348054
rect 238822 347818 239004 348054
rect 238404 347734 239004 347818
rect 238404 347498 238586 347734
rect 238822 347498 239004 347734
rect 238404 312054 239004 347498
rect 238404 311818 238586 312054
rect 238822 311818 239004 312054
rect 238404 311734 239004 311818
rect 238404 311498 238586 311734
rect 238822 311498 239004 311734
rect 238404 276054 239004 311498
rect 238404 275818 238586 276054
rect 238822 275818 239004 276054
rect 238404 275734 239004 275818
rect 238404 275498 238586 275734
rect 238822 275498 239004 275734
rect 238404 240054 239004 275498
rect 238404 239818 238586 240054
rect 238822 239818 239004 240054
rect 238404 239734 239004 239818
rect 238404 239498 238586 239734
rect 238822 239498 239004 239734
rect 238404 204054 239004 239498
rect 238404 203818 238586 204054
rect 238822 203818 239004 204054
rect 238404 203734 239004 203818
rect 238404 203498 238586 203734
rect 238822 203498 239004 203734
rect 238404 168054 239004 203498
rect 238404 167818 238586 168054
rect 238822 167818 239004 168054
rect 238404 167734 239004 167818
rect 238404 167498 238586 167734
rect 238822 167498 239004 167734
rect 238404 132054 239004 167498
rect 238404 131818 238586 132054
rect 238822 131818 239004 132054
rect 238404 131734 239004 131818
rect 238404 131498 238586 131734
rect 238822 131498 239004 131734
rect 238404 96054 239004 131498
rect 238404 95818 238586 96054
rect 238822 95818 239004 96054
rect 238404 95734 239004 95818
rect 238404 95498 238586 95734
rect 238822 95498 239004 95734
rect 238404 60054 239004 95498
rect 238404 59818 238586 60054
rect 238822 59818 239004 60054
rect 238404 59734 239004 59818
rect 238404 59498 238586 59734
rect 238822 59498 239004 59734
rect 238404 24054 239004 59498
rect 238404 23818 238586 24054
rect 238822 23818 239004 24054
rect 238404 23734 239004 23818
rect 238404 23498 238586 23734
rect 238822 23498 239004 23734
rect 238404 -3166 239004 23498
rect 238404 -3402 238586 -3166
rect 238822 -3402 239004 -3166
rect 238404 -3486 239004 -3402
rect 238404 -3722 238586 -3486
rect 238822 -3722 239004 -3486
rect 238404 -3744 239004 -3722
rect 242004 675654 242604 708982
rect 242004 675418 242186 675654
rect 242422 675418 242604 675654
rect 242004 675334 242604 675418
rect 242004 675098 242186 675334
rect 242422 675098 242604 675334
rect 242004 639654 242604 675098
rect 242004 639418 242186 639654
rect 242422 639418 242604 639654
rect 242004 639334 242604 639418
rect 242004 639098 242186 639334
rect 242422 639098 242604 639334
rect 242004 603654 242604 639098
rect 242004 603418 242186 603654
rect 242422 603418 242604 603654
rect 242004 603334 242604 603418
rect 242004 603098 242186 603334
rect 242422 603098 242604 603334
rect 242004 567654 242604 603098
rect 242004 567418 242186 567654
rect 242422 567418 242604 567654
rect 242004 567334 242604 567418
rect 242004 567098 242186 567334
rect 242422 567098 242604 567334
rect 242004 531654 242604 567098
rect 242004 531418 242186 531654
rect 242422 531418 242604 531654
rect 242004 531334 242604 531418
rect 242004 531098 242186 531334
rect 242422 531098 242604 531334
rect 242004 495654 242604 531098
rect 242004 495418 242186 495654
rect 242422 495418 242604 495654
rect 242004 495334 242604 495418
rect 242004 495098 242186 495334
rect 242422 495098 242604 495334
rect 242004 459654 242604 495098
rect 242004 459418 242186 459654
rect 242422 459418 242604 459654
rect 242004 459334 242604 459418
rect 242004 459098 242186 459334
rect 242422 459098 242604 459334
rect 242004 423654 242604 459098
rect 242004 423418 242186 423654
rect 242422 423418 242604 423654
rect 242004 423334 242604 423418
rect 242004 423098 242186 423334
rect 242422 423098 242604 423334
rect 242004 387654 242604 423098
rect 242004 387418 242186 387654
rect 242422 387418 242604 387654
rect 242004 387334 242604 387418
rect 242004 387098 242186 387334
rect 242422 387098 242604 387334
rect 242004 351654 242604 387098
rect 242004 351418 242186 351654
rect 242422 351418 242604 351654
rect 242004 351334 242604 351418
rect 242004 351098 242186 351334
rect 242422 351098 242604 351334
rect 242004 315654 242604 351098
rect 242004 315418 242186 315654
rect 242422 315418 242604 315654
rect 242004 315334 242604 315418
rect 242004 315098 242186 315334
rect 242422 315098 242604 315334
rect 242004 279654 242604 315098
rect 242004 279418 242186 279654
rect 242422 279418 242604 279654
rect 242004 279334 242604 279418
rect 242004 279098 242186 279334
rect 242422 279098 242604 279334
rect 242004 243654 242604 279098
rect 242004 243418 242186 243654
rect 242422 243418 242604 243654
rect 242004 243334 242604 243418
rect 242004 243098 242186 243334
rect 242422 243098 242604 243334
rect 242004 207654 242604 243098
rect 242004 207418 242186 207654
rect 242422 207418 242604 207654
rect 242004 207334 242604 207418
rect 242004 207098 242186 207334
rect 242422 207098 242604 207334
rect 242004 171654 242604 207098
rect 242004 171418 242186 171654
rect 242422 171418 242604 171654
rect 242004 171334 242604 171418
rect 242004 171098 242186 171334
rect 242422 171098 242604 171334
rect 242004 135654 242604 171098
rect 242004 135418 242186 135654
rect 242422 135418 242604 135654
rect 242004 135334 242604 135418
rect 242004 135098 242186 135334
rect 242422 135098 242604 135334
rect 242004 99654 242604 135098
rect 242004 99418 242186 99654
rect 242422 99418 242604 99654
rect 242004 99334 242604 99418
rect 242004 99098 242186 99334
rect 242422 99098 242604 99334
rect 242004 63654 242604 99098
rect 242004 63418 242186 63654
rect 242422 63418 242604 63654
rect 242004 63334 242604 63418
rect 242004 63098 242186 63334
rect 242422 63098 242604 63334
rect 242004 27654 242604 63098
rect 242004 27418 242186 27654
rect 242422 27418 242604 27654
rect 242004 27334 242604 27418
rect 242004 27098 242186 27334
rect 242422 27098 242604 27334
rect 242004 -5046 242604 27098
rect 242004 -5282 242186 -5046
rect 242422 -5282 242604 -5046
rect 242004 -5366 242604 -5282
rect 242004 -5602 242186 -5366
rect 242422 -5602 242604 -5366
rect 242004 -5624 242604 -5602
rect 245604 679254 246204 710862
rect 263604 710478 264204 711440
rect 263604 710242 263786 710478
rect 264022 710242 264204 710478
rect 263604 710158 264204 710242
rect 263604 709922 263786 710158
rect 264022 709922 264204 710158
rect 260004 708598 260604 709560
rect 260004 708362 260186 708598
rect 260422 708362 260604 708598
rect 260004 708278 260604 708362
rect 260004 708042 260186 708278
rect 260422 708042 260604 708278
rect 256404 706718 257004 707680
rect 256404 706482 256586 706718
rect 256822 706482 257004 706718
rect 256404 706398 257004 706482
rect 256404 706162 256586 706398
rect 256822 706162 257004 706398
rect 245604 679018 245786 679254
rect 246022 679018 246204 679254
rect 245604 678934 246204 679018
rect 245604 678698 245786 678934
rect 246022 678698 246204 678934
rect 245604 643254 246204 678698
rect 245604 643018 245786 643254
rect 246022 643018 246204 643254
rect 245604 642934 246204 643018
rect 245604 642698 245786 642934
rect 246022 642698 246204 642934
rect 245604 607254 246204 642698
rect 245604 607018 245786 607254
rect 246022 607018 246204 607254
rect 245604 606934 246204 607018
rect 245604 606698 245786 606934
rect 246022 606698 246204 606934
rect 245604 571254 246204 606698
rect 245604 571018 245786 571254
rect 246022 571018 246204 571254
rect 245604 570934 246204 571018
rect 245604 570698 245786 570934
rect 246022 570698 246204 570934
rect 245604 535254 246204 570698
rect 245604 535018 245786 535254
rect 246022 535018 246204 535254
rect 245604 534934 246204 535018
rect 245604 534698 245786 534934
rect 246022 534698 246204 534934
rect 245604 499254 246204 534698
rect 245604 499018 245786 499254
rect 246022 499018 246204 499254
rect 245604 498934 246204 499018
rect 245604 498698 245786 498934
rect 246022 498698 246204 498934
rect 245604 463254 246204 498698
rect 245604 463018 245786 463254
rect 246022 463018 246204 463254
rect 245604 462934 246204 463018
rect 245604 462698 245786 462934
rect 246022 462698 246204 462934
rect 245604 427254 246204 462698
rect 245604 427018 245786 427254
rect 246022 427018 246204 427254
rect 245604 426934 246204 427018
rect 245604 426698 245786 426934
rect 246022 426698 246204 426934
rect 245604 391254 246204 426698
rect 245604 391018 245786 391254
rect 246022 391018 246204 391254
rect 245604 390934 246204 391018
rect 245604 390698 245786 390934
rect 246022 390698 246204 390934
rect 245604 355254 246204 390698
rect 245604 355018 245786 355254
rect 246022 355018 246204 355254
rect 245604 354934 246204 355018
rect 245604 354698 245786 354934
rect 246022 354698 246204 354934
rect 245604 319254 246204 354698
rect 245604 319018 245786 319254
rect 246022 319018 246204 319254
rect 245604 318934 246204 319018
rect 245604 318698 245786 318934
rect 246022 318698 246204 318934
rect 245604 283254 246204 318698
rect 245604 283018 245786 283254
rect 246022 283018 246204 283254
rect 245604 282934 246204 283018
rect 245604 282698 245786 282934
rect 246022 282698 246204 282934
rect 245604 247254 246204 282698
rect 245604 247018 245786 247254
rect 246022 247018 246204 247254
rect 245604 246934 246204 247018
rect 245604 246698 245786 246934
rect 246022 246698 246204 246934
rect 245604 211254 246204 246698
rect 245604 211018 245786 211254
rect 246022 211018 246204 211254
rect 245604 210934 246204 211018
rect 245604 210698 245786 210934
rect 246022 210698 246204 210934
rect 245604 175254 246204 210698
rect 245604 175018 245786 175254
rect 246022 175018 246204 175254
rect 245604 174934 246204 175018
rect 245604 174698 245786 174934
rect 246022 174698 246204 174934
rect 245604 139254 246204 174698
rect 245604 139018 245786 139254
rect 246022 139018 246204 139254
rect 245604 138934 246204 139018
rect 245604 138698 245786 138934
rect 246022 138698 246204 138934
rect 245604 103254 246204 138698
rect 245604 103018 245786 103254
rect 246022 103018 246204 103254
rect 245604 102934 246204 103018
rect 245604 102698 245786 102934
rect 246022 102698 246204 102934
rect 245604 67254 246204 102698
rect 245604 67018 245786 67254
rect 246022 67018 246204 67254
rect 245604 66934 246204 67018
rect 245604 66698 245786 66934
rect 246022 66698 246204 66934
rect 245604 31254 246204 66698
rect 245604 31018 245786 31254
rect 246022 31018 246204 31254
rect 245604 30934 246204 31018
rect 245604 30698 245786 30934
rect 246022 30698 246204 30934
rect 227604 -6222 227786 -5986
rect 228022 -6222 228204 -5986
rect 227604 -6306 228204 -6222
rect 227604 -6542 227786 -6306
rect 228022 -6542 228204 -6306
rect 227604 -7504 228204 -6542
rect 245604 -6926 246204 30698
rect 252804 704838 253404 705800
rect 252804 704602 252986 704838
rect 253222 704602 253404 704838
rect 252804 704518 253404 704602
rect 252804 704282 252986 704518
rect 253222 704282 253404 704518
rect 252804 686454 253404 704282
rect 252804 686218 252986 686454
rect 253222 686218 253404 686454
rect 252804 686134 253404 686218
rect 252804 685898 252986 686134
rect 253222 685898 253404 686134
rect 252804 650454 253404 685898
rect 252804 650218 252986 650454
rect 253222 650218 253404 650454
rect 252804 650134 253404 650218
rect 252804 649898 252986 650134
rect 253222 649898 253404 650134
rect 252804 614454 253404 649898
rect 252804 614218 252986 614454
rect 253222 614218 253404 614454
rect 252804 614134 253404 614218
rect 252804 613898 252986 614134
rect 253222 613898 253404 614134
rect 252804 578454 253404 613898
rect 252804 578218 252986 578454
rect 253222 578218 253404 578454
rect 252804 578134 253404 578218
rect 252804 577898 252986 578134
rect 253222 577898 253404 578134
rect 252804 542454 253404 577898
rect 252804 542218 252986 542454
rect 253222 542218 253404 542454
rect 252804 542134 253404 542218
rect 252804 541898 252986 542134
rect 253222 541898 253404 542134
rect 252804 506454 253404 541898
rect 252804 506218 252986 506454
rect 253222 506218 253404 506454
rect 252804 506134 253404 506218
rect 252804 505898 252986 506134
rect 253222 505898 253404 506134
rect 252804 470454 253404 505898
rect 256404 690054 257004 706162
rect 256404 689818 256586 690054
rect 256822 689818 257004 690054
rect 256404 689734 257004 689818
rect 256404 689498 256586 689734
rect 256822 689498 257004 689734
rect 256404 654054 257004 689498
rect 256404 653818 256586 654054
rect 256822 653818 257004 654054
rect 256404 653734 257004 653818
rect 256404 653498 256586 653734
rect 256822 653498 257004 653734
rect 256404 618054 257004 653498
rect 256404 617818 256586 618054
rect 256822 617818 257004 618054
rect 256404 617734 257004 617818
rect 256404 617498 256586 617734
rect 256822 617498 257004 617734
rect 256404 582054 257004 617498
rect 256404 581818 256586 582054
rect 256822 581818 257004 582054
rect 256404 581734 257004 581818
rect 256404 581498 256586 581734
rect 256822 581498 257004 581734
rect 256404 546054 257004 581498
rect 256404 545818 256586 546054
rect 256822 545818 257004 546054
rect 256404 545734 257004 545818
rect 256404 545498 256586 545734
rect 256822 545498 257004 545734
rect 256404 510054 257004 545498
rect 256404 509818 256586 510054
rect 256822 509818 257004 510054
rect 256404 509734 257004 509818
rect 256404 509498 256586 509734
rect 256822 509498 257004 509734
rect 256404 483000 257004 509498
rect 260004 693654 260604 708042
rect 260004 693418 260186 693654
rect 260422 693418 260604 693654
rect 260004 693334 260604 693418
rect 260004 693098 260186 693334
rect 260422 693098 260604 693334
rect 260004 657654 260604 693098
rect 260004 657418 260186 657654
rect 260422 657418 260604 657654
rect 260004 657334 260604 657418
rect 260004 657098 260186 657334
rect 260422 657098 260604 657334
rect 260004 621654 260604 657098
rect 260004 621418 260186 621654
rect 260422 621418 260604 621654
rect 260004 621334 260604 621418
rect 260004 621098 260186 621334
rect 260422 621098 260604 621334
rect 260004 585654 260604 621098
rect 260004 585418 260186 585654
rect 260422 585418 260604 585654
rect 260004 585334 260604 585418
rect 260004 585098 260186 585334
rect 260422 585098 260604 585334
rect 260004 549654 260604 585098
rect 260004 549418 260186 549654
rect 260422 549418 260604 549654
rect 260004 549334 260604 549418
rect 260004 549098 260186 549334
rect 260422 549098 260604 549334
rect 260004 513654 260604 549098
rect 260004 513418 260186 513654
rect 260422 513418 260604 513654
rect 260004 513334 260604 513418
rect 260004 513098 260186 513334
rect 260422 513098 260604 513334
rect 260004 483000 260604 513098
rect 263604 697254 264204 709922
rect 281604 711418 282204 711440
rect 281604 711182 281786 711418
rect 282022 711182 282204 711418
rect 281604 711098 282204 711182
rect 281604 710862 281786 711098
rect 282022 710862 282204 711098
rect 278004 709538 278604 709560
rect 278004 709302 278186 709538
rect 278422 709302 278604 709538
rect 278004 709218 278604 709302
rect 278004 708982 278186 709218
rect 278422 708982 278604 709218
rect 274404 707658 275004 707680
rect 274404 707422 274586 707658
rect 274822 707422 275004 707658
rect 274404 707338 275004 707422
rect 274404 707102 274586 707338
rect 274822 707102 275004 707338
rect 263604 697018 263786 697254
rect 264022 697018 264204 697254
rect 263604 696934 264204 697018
rect 263604 696698 263786 696934
rect 264022 696698 264204 696934
rect 263604 661254 264204 696698
rect 263604 661018 263786 661254
rect 264022 661018 264204 661254
rect 263604 660934 264204 661018
rect 263604 660698 263786 660934
rect 264022 660698 264204 660934
rect 263604 625254 264204 660698
rect 263604 625018 263786 625254
rect 264022 625018 264204 625254
rect 263604 624934 264204 625018
rect 263604 624698 263786 624934
rect 264022 624698 264204 624934
rect 263604 589254 264204 624698
rect 263604 589018 263786 589254
rect 264022 589018 264204 589254
rect 263604 588934 264204 589018
rect 263604 588698 263786 588934
rect 264022 588698 264204 588934
rect 263604 553254 264204 588698
rect 263604 553018 263786 553254
rect 264022 553018 264204 553254
rect 263604 552934 264204 553018
rect 263604 552698 263786 552934
rect 264022 552698 264204 552934
rect 263604 517254 264204 552698
rect 263604 517018 263786 517254
rect 264022 517018 264204 517254
rect 263604 516934 264204 517018
rect 263604 516698 263786 516934
rect 264022 516698 264204 516934
rect 263604 483000 264204 516698
rect 270804 705778 271404 705800
rect 270804 705542 270986 705778
rect 271222 705542 271404 705778
rect 270804 705458 271404 705542
rect 270804 705222 270986 705458
rect 271222 705222 271404 705458
rect 270804 668454 271404 705222
rect 270804 668218 270986 668454
rect 271222 668218 271404 668454
rect 270804 668134 271404 668218
rect 270804 667898 270986 668134
rect 271222 667898 271404 668134
rect 270804 632454 271404 667898
rect 270804 632218 270986 632454
rect 271222 632218 271404 632454
rect 270804 632134 271404 632218
rect 270804 631898 270986 632134
rect 271222 631898 271404 632134
rect 270804 596454 271404 631898
rect 270804 596218 270986 596454
rect 271222 596218 271404 596454
rect 270804 596134 271404 596218
rect 270804 595898 270986 596134
rect 271222 595898 271404 596134
rect 270804 560454 271404 595898
rect 270804 560218 270986 560454
rect 271222 560218 271404 560454
rect 270804 560134 271404 560218
rect 270804 559898 270986 560134
rect 271222 559898 271404 560134
rect 270804 524454 271404 559898
rect 270804 524218 270986 524454
rect 271222 524218 271404 524454
rect 270804 524134 271404 524218
rect 270804 523898 270986 524134
rect 271222 523898 271404 524134
rect 270804 488454 271404 523898
rect 270804 488218 270986 488454
rect 271222 488218 271404 488454
rect 270804 488134 271404 488218
rect 270804 487898 270986 488134
rect 271222 487898 271404 488134
rect 270804 483000 271404 487898
rect 274404 672054 275004 707102
rect 274404 671818 274586 672054
rect 274822 671818 275004 672054
rect 274404 671734 275004 671818
rect 274404 671498 274586 671734
rect 274822 671498 275004 671734
rect 274404 636054 275004 671498
rect 274404 635818 274586 636054
rect 274822 635818 275004 636054
rect 274404 635734 275004 635818
rect 274404 635498 274586 635734
rect 274822 635498 275004 635734
rect 274404 600054 275004 635498
rect 274404 599818 274586 600054
rect 274822 599818 275004 600054
rect 274404 599734 275004 599818
rect 274404 599498 274586 599734
rect 274822 599498 275004 599734
rect 274404 564054 275004 599498
rect 274404 563818 274586 564054
rect 274822 563818 275004 564054
rect 274404 563734 275004 563818
rect 274404 563498 274586 563734
rect 274822 563498 275004 563734
rect 274404 528054 275004 563498
rect 274404 527818 274586 528054
rect 274822 527818 275004 528054
rect 274404 527734 275004 527818
rect 274404 527498 274586 527734
rect 274822 527498 275004 527734
rect 274404 492054 275004 527498
rect 274404 491818 274586 492054
rect 274822 491818 275004 492054
rect 274404 491734 275004 491818
rect 274404 491498 274586 491734
rect 274822 491498 275004 491734
rect 274404 483000 275004 491498
rect 278004 675654 278604 708982
rect 278004 675418 278186 675654
rect 278422 675418 278604 675654
rect 278004 675334 278604 675418
rect 278004 675098 278186 675334
rect 278422 675098 278604 675334
rect 278004 639654 278604 675098
rect 278004 639418 278186 639654
rect 278422 639418 278604 639654
rect 278004 639334 278604 639418
rect 278004 639098 278186 639334
rect 278422 639098 278604 639334
rect 278004 603654 278604 639098
rect 278004 603418 278186 603654
rect 278422 603418 278604 603654
rect 278004 603334 278604 603418
rect 278004 603098 278186 603334
rect 278422 603098 278604 603334
rect 278004 567654 278604 603098
rect 278004 567418 278186 567654
rect 278422 567418 278604 567654
rect 278004 567334 278604 567418
rect 278004 567098 278186 567334
rect 278422 567098 278604 567334
rect 278004 531654 278604 567098
rect 278004 531418 278186 531654
rect 278422 531418 278604 531654
rect 278004 531334 278604 531418
rect 278004 531098 278186 531334
rect 278422 531098 278604 531334
rect 278004 495654 278604 531098
rect 278004 495418 278186 495654
rect 278422 495418 278604 495654
rect 278004 495334 278604 495418
rect 278004 495098 278186 495334
rect 278422 495098 278604 495334
rect 278004 483000 278604 495098
rect 281604 679254 282204 710862
rect 299604 710478 300204 711440
rect 299604 710242 299786 710478
rect 300022 710242 300204 710478
rect 299604 710158 300204 710242
rect 299604 709922 299786 710158
rect 300022 709922 300204 710158
rect 296004 708598 296604 709560
rect 296004 708362 296186 708598
rect 296422 708362 296604 708598
rect 296004 708278 296604 708362
rect 296004 708042 296186 708278
rect 296422 708042 296604 708278
rect 292404 706718 293004 707680
rect 292404 706482 292586 706718
rect 292822 706482 293004 706718
rect 292404 706398 293004 706482
rect 292404 706162 292586 706398
rect 292822 706162 293004 706398
rect 281604 679018 281786 679254
rect 282022 679018 282204 679254
rect 281604 678934 282204 679018
rect 281604 678698 281786 678934
rect 282022 678698 282204 678934
rect 281604 643254 282204 678698
rect 281604 643018 281786 643254
rect 282022 643018 282204 643254
rect 281604 642934 282204 643018
rect 281604 642698 281786 642934
rect 282022 642698 282204 642934
rect 281604 607254 282204 642698
rect 281604 607018 281786 607254
rect 282022 607018 282204 607254
rect 281604 606934 282204 607018
rect 281604 606698 281786 606934
rect 282022 606698 282204 606934
rect 281604 571254 282204 606698
rect 281604 571018 281786 571254
rect 282022 571018 282204 571254
rect 281604 570934 282204 571018
rect 281604 570698 281786 570934
rect 282022 570698 282204 570934
rect 281604 535254 282204 570698
rect 281604 535018 281786 535254
rect 282022 535018 282204 535254
rect 281604 534934 282204 535018
rect 281604 534698 281786 534934
rect 282022 534698 282204 534934
rect 281604 499254 282204 534698
rect 281604 499018 281786 499254
rect 282022 499018 282204 499254
rect 281604 498934 282204 499018
rect 281604 498698 281786 498934
rect 282022 498698 282204 498934
rect 281604 483000 282204 498698
rect 288804 704838 289404 705800
rect 288804 704602 288986 704838
rect 289222 704602 289404 704838
rect 288804 704518 289404 704602
rect 288804 704282 288986 704518
rect 289222 704282 289404 704518
rect 288804 686454 289404 704282
rect 288804 686218 288986 686454
rect 289222 686218 289404 686454
rect 288804 686134 289404 686218
rect 288804 685898 288986 686134
rect 289222 685898 289404 686134
rect 288804 650454 289404 685898
rect 288804 650218 288986 650454
rect 289222 650218 289404 650454
rect 288804 650134 289404 650218
rect 288804 649898 288986 650134
rect 289222 649898 289404 650134
rect 288804 614454 289404 649898
rect 288804 614218 288986 614454
rect 289222 614218 289404 614454
rect 288804 614134 289404 614218
rect 288804 613898 288986 614134
rect 289222 613898 289404 614134
rect 288804 578454 289404 613898
rect 288804 578218 288986 578454
rect 289222 578218 289404 578454
rect 288804 578134 289404 578218
rect 288804 577898 288986 578134
rect 289222 577898 289404 578134
rect 288804 542454 289404 577898
rect 288804 542218 288986 542454
rect 289222 542218 289404 542454
rect 288804 542134 289404 542218
rect 288804 541898 288986 542134
rect 289222 541898 289404 542134
rect 288804 506454 289404 541898
rect 288804 506218 288986 506454
rect 289222 506218 289404 506454
rect 288804 506134 289404 506218
rect 288804 505898 288986 506134
rect 289222 505898 289404 506134
rect 288804 483000 289404 505898
rect 292404 690054 293004 706162
rect 292404 689818 292586 690054
rect 292822 689818 293004 690054
rect 292404 689734 293004 689818
rect 292404 689498 292586 689734
rect 292822 689498 293004 689734
rect 292404 654054 293004 689498
rect 292404 653818 292586 654054
rect 292822 653818 293004 654054
rect 292404 653734 293004 653818
rect 292404 653498 292586 653734
rect 292822 653498 293004 653734
rect 292404 618054 293004 653498
rect 292404 617818 292586 618054
rect 292822 617818 293004 618054
rect 292404 617734 293004 617818
rect 292404 617498 292586 617734
rect 292822 617498 293004 617734
rect 292404 582054 293004 617498
rect 292404 581818 292586 582054
rect 292822 581818 293004 582054
rect 292404 581734 293004 581818
rect 292404 581498 292586 581734
rect 292822 581498 293004 581734
rect 292404 546054 293004 581498
rect 292404 545818 292586 546054
rect 292822 545818 293004 546054
rect 292404 545734 293004 545818
rect 292404 545498 292586 545734
rect 292822 545498 293004 545734
rect 292404 510054 293004 545498
rect 292404 509818 292586 510054
rect 292822 509818 293004 510054
rect 292404 509734 293004 509818
rect 292404 509498 292586 509734
rect 292822 509498 293004 509734
rect 292404 483000 293004 509498
rect 296004 693654 296604 708042
rect 296004 693418 296186 693654
rect 296422 693418 296604 693654
rect 296004 693334 296604 693418
rect 296004 693098 296186 693334
rect 296422 693098 296604 693334
rect 296004 657654 296604 693098
rect 296004 657418 296186 657654
rect 296422 657418 296604 657654
rect 296004 657334 296604 657418
rect 296004 657098 296186 657334
rect 296422 657098 296604 657334
rect 296004 621654 296604 657098
rect 296004 621418 296186 621654
rect 296422 621418 296604 621654
rect 296004 621334 296604 621418
rect 296004 621098 296186 621334
rect 296422 621098 296604 621334
rect 296004 585654 296604 621098
rect 299604 697254 300204 709922
rect 317604 711418 318204 711440
rect 317604 711182 317786 711418
rect 318022 711182 318204 711418
rect 317604 711098 318204 711182
rect 317604 710862 317786 711098
rect 318022 710862 318204 711098
rect 314004 709538 314604 709560
rect 314004 709302 314186 709538
rect 314422 709302 314604 709538
rect 314004 709218 314604 709302
rect 314004 708982 314186 709218
rect 314422 708982 314604 709218
rect 310404 707658 311004 707680
rect 310404 707422 310586 707658
rect 310822 707422 311004 707658
rect 310404 707338 311004 707422
rect 310404 707102 310586 707338
rect 310822 707102 311004 707338
rect 299604 697018 299786 697254
rect 300022 697018 300204 697254
rect 299604 696934 300204 697018
rect 299604 696698 299786 696934
rect 300022 696698 300204 696934
rect 299604 661254 300204 696698
rect 299604 661018 299786 661254
rect 300022 661018 300204 661254
rect 299604 660934 300204 661018
rect 299604 660698 299786 660934
rect 300022 660698 300204 660934
rect 299604 625254 300204 660698
rect 299604 625018 299786 625254
rect 300022 625018 300204 625254
rect 299604 624934 300204 625018
rect 299604 624698 299786 624934
rect 300022 624698 300204 624934
rect 299604 614247 300204 624698
rect 306804 705778 307404 705800
rect 306804 705542 306986 705778
rect 307222 705542 307404 705778
rect 306804 705458 307404 705542
rect 306804 705222 306986 705458
rect 307222 705222 307404 705458
rect 306804 668454 307404 705222
rect 306804 668218 306986 668454
rect 307222 668218 307404 668454
rect 306804 668134 307404 668218
rect 306804 667898 306986 668134
rect 307222 667898 307404 668134
rect 306804 632454 307404 667898
rect 306804 632218 306986 632454
rect 307222 632218 307404 632454
rect 306804 632134 307404 632218
rect 306804 631898 306986 632134
rect 307222 631898 307404 632134
rect 306804 614247 307404 631898
rect 310404 672054 311004 707102
rect 310404 671818 310586 672054
rect 310822 671818 311004 672054
rect 310404 671734 311004 671818
rect 310404 671498 310586 671734
rect 310822 671498 311004 671734
rect 310404 636054 311004 671498
rect 310404 635818 310586 636054
rect 310822 635818 311004 636054
rect 310404 635734 311004 635818
rect 310404 635498 310586 635734
rect 310822 635498 311004 635734
rect 310404 614247 311004 635498
rect 314004 675654 314604 708982
rect 314004 675418 314186 675654
rect 314422 675418 314604 675654
rect 314004 675334 314604 675418
rect 314004 675098 314186 675334
rect 314422 675098 314604 675334
rect 314004 639654 314604 675098
rect 314004 639418 314186 639654
rect 314422 639418 314604 639654
rect 314004 639334 314604 639418
rect 314004 639098 314186 639334
rect 314422 639098 314604 639334
rect 314004 614247 314604 639098
rect 317604 679254 318204 710862
rect 335604 710478 336204 711440
rect 335604 710242 335786 710478
rect 336022 710242 336204 710478
rect 335604 710158 336204 710242
rect 335604 709922 335786 710158
rect 336022 709922 336204 710158
rect 332004 708598 332604 709560
rect 332004 708362 332186 708598
rect 332422 708362 332604 708598
rect 332004 708278 332604 708362
rect 332004 708042 332186 708278
rect 332422 708042 332604 708278
rect 328404 706718 329004 707680
rect 328404 706482 328586 706718
rect 328822 706482 329004 706718
rect 328404 706398 329004 706482
rect 328404 706162 328586 706398
rect 328822 706162 329004 706398
rect 317604 679018 317786 679254
rect 318022 679018 318204 679254
rect 317604 678934 318204 679018
rect 317604 678698 317786 678934
rect 318022 678698 318204 678934
rect 317604 643254 318204 678698
rect 317604 643018 317786 643254
rect 318022 643018 318204 643254
rect 317604 642934 318204 643018
rect 317604 642698 317786 642934
rect 318022 642698 318204 642934
rect 317604 614247 318204 642698
rect 324804 704838 325404 705800
rect 324804 704602 324986 704838
rect 325222 704602 325404 704838
rect 324804 704518 325404 704602
rect 324804 704282 324986 704518
rect 325222 704282 325404 704518
rect 324804 686454 325404 704282
rect 324804 686218 324986 686454
rect 325222 686218 325404 686454
rect 324804 686134 325404 686218
rect 324804 685898 324986 686134
rect 325222 685898 325404 686134
rect 324804 650454 325404 685898
rect 324804 650218 324986 650454
rect 325222 650218 325404 650454
rect 324804 650134 325404 650218
rect 324804 649898 324986 650134
rect 325222 649898 325404 650134
rect 324804 614247 325404 649898
rect 328404 690054 329004 706162
rect 328404 689818 328586 690054
rect 328822 689818 329004 690054
rect 328404 689734 329004 689818
rect 328404 689498 328586 689734
rect 328822 689498 329004 689734
rect 328404 654054 329004 689498
rect 328404 653818 328586 654054
rect 328822 653818 329004 654054
rect 328404 653734 329004 653818
rect 328404 653498 328586 653734
rect 328822 653498 329004 653734
rect 328404 618054 329004 653498
rect 328404 617818 328586 618054
rect 328822 617818 329004 618054
rect 328404 617734 329004 617818
rect 328404 617498 328586 617734
rect 328822 617498 329004 617734
rect 328404 614247 329004 617498
rect 332004 693654 332604 708042
rect 332004 693418 332186 693654
rect 332422 693418 332604 693654
rect 332004 693334 332604 693418
rect 332004 693098 332186 693334
rect 332422 693098 332604 693334
rect 332004 657654 332604 693098
rect 332004 657418 332186 657654
rect 332422 657418 332604 657654
rect 332004 657334 332604 657418
rect 332004 657098 332186 657334
rect 332422 657098 332604 657334
rect 332004 621654 332604 657098
rect 332004 621418 332186 621654
rect 332422 621418 332604 621654
rect 332004 621334 332604 621418
rect 332004 621098 332186 621334
rect 332422 621098 332604 621334
rect 332004 614247 332604 621098
rect 335604 697254 336204 709922
rect 353604 711418 354204 711440
rect 353604 711182 353786 711418
rect 354022 711182 354204 711418
rect 353604 711098 354204 711182
rect 353604 710862 353786 711098
rect 354022 710862 354204 711098
rect 350004 709538 350604 709560
rect 350004 709302 350186 709538
rect 350422 709302 350604 709538
rect 350004 709218 350604 709302
rect 350004 708982 350186 709218
rect 350422 708982 350604 709218
rect 346404 707658 347004 707680
rect 346404 707422 346586 707658
rect 346822 707422 347004 707658
rect 346404 707338 347004 707422
rect 346404 707102 346586 707338
rect 346822 707102 347004 707338
rect 335604 697018 335786 697254
rect 336022 697018 336204 697254
rect 335604 696934 336204 697018
rect 335604 696698 335786 696934
rect 336022 696698 336204 696934
rect 335604 661254 336204 696698
rect 335604 661018 335786 661254
rect 336022 661018 336204 661254
rect 335604 660934 336204 661018
rect 335604 660698 335786 660934
rect 336022 660698 336204 660934
rect 335604 625254 336204 660698
rect 335604 625018 335786 625254
rect 336022 625018 336204 625254
rect 335604 624934 336204 625018
rect 335604 624698 335786 624934
rect 336022 624698 336204 624934
rect 335604 614247 336204 624698
rect 342804 705778 343404 705800
rect 342804 705542 342986 705778
rect 343222 705542 343404 705778
rect 342804 705458 343404 705542
rect 342804 705222 342986 705458
rect 343222 705222 343404 705458
rect 342804 668454 343404 705222
rect 342804 668218 342986 668454
rect 343222 668218 343404 668454
rect 342804 668134 343404 668218
rect 342804 667898 342986 668134
rect 343222 667898 343404 668134
rect 342804 632454 343404 667898
rect 342804 632218 342986 632454
rect 343222 632218 343404 632454
rect 342804 632134 343404 632218
rect 342804 631898 342986 632134
rect 343222 631898 343404 632134
rect 342804 614247 343404 631898
rect 346404 672054 347004 707102
rect 346404 671818 346586 672054
rect 346822 671818 347004 672054
rect 346404 671734 347004 671818
rect 346404 671498 346586 671734
rect 346822 671498 347004 671734
rect 346404 636054 347004 671498
rect 346404 635818 346586 636054
rect 346822 635818 347004 636054
rect 346404 635734 347004 635818
rect 346404 635498 346586 635734
rect 346822 635498 347004 635734
rect 346404 614247 347004 635498
rect 350004 675654 350604 708982
rect 350004 675418 350186 675654
rect 350422 675418 350604 675654
rect 350004 675334 350604 675418
rect 350004 675098 350186 675334
rect 350422 675098 350604 675334
rect 350004 639654 350604 675098
rect 350004 639418 350186 639654
rect 350422 639418 350604 639654
rect 350004 639334 350604 639418
rect 350004 639098 350186 639334
rect 350422 639098 350604 639334
rect 350004 614247 350604 639098
rect 353604 679254 354204 710862
rect 371604 710478 372204 711440
rect 371604 710242 371786 710478
rect 372022 710242 372204 710478
rect 371604 710158 372204 710242
rect 371604 709922 371786 710158
rect 372022 709922 372204 710158
rect 368004 708598 368604 709560
rect 368004 708362 368186 708598
rect 368422 708362 368604 708598
rect 368004 708278 368604 708362
rect 368004 708042 368186 708278
rect 368422 708042 368604 708278
rect 364404 706718 365004 707680
rect 364404 706482 364586 706718
rect 364822 706482 365004 706718
rect 364404 706398 365004 706482
rect 364404 706162 364586 706398
rect 364822 706162 365004 706398
rect 353604 679018 353786 679254
rect 354022 679018 354204 679254
rect 353604 678934 354204 679018
rect 353604 678698 353786 678934
rect 354022 678698 354204 678934
rect 353604 643254 354204 678698
rect 353604 643018 353786 643254
rect 354022 643018 354204 643254
rect 353604 642934 354204 643018
rect 353604 642698 353786 642934
rect 354022 642698 354204 642934
rect 353604 614247 354204 642698
rect 360804 704838 361404 705800
rect 360804 704602 360986 704838
rect 361222 704602 361404 704838
rect 360804 704518 361404 704602
rect 360804 704282 360986 704518
rect 361222 704282 361404 704518
rect 360804 686454 361404 704282
rect 360804 686218 360986 686454
rect 361222 686218 361404 686454
rect 360804 686134 361404 686218
rect 360804 685898 360986 686134
rect 361222 685898 361404 686134
rect 360804 650454 361404 685898
rect 360804 650218 360986 650454
rect 361222 650218 361404 650454
rect 360804 650134 361404 650218
rect 360804 649898 360986 650134
rect 361222 649898 361404 650134
rect 360804 614247 361404 649898
rect 364404 690054 365004 706162
rect 364404 689818 364586 690054
rect 364822 689818 365004 690054
rect 364404 689734 365004 689818
rect 364404 689498 364586 689734
rect 364822 689498 365004 689734
rect 364404 654054 365004 689498
rect 364404 653818 364586 654054
rect 364822 653818 365004 654054
rect 364404 653734 365004 653818
rect 364404 653498 364586 653734
rect 364822 653498 365004 653734
rect 364404 618054 365004 653498
rect 364404 617818 364586 618054
rect 364822 617818 365004 618054
rect 364404 617734 365004 617818
rect 364404 617498 364586 617734
rect 364822 617498 365004 617734
rect 364404 614247 365004 617498
rect 368004 693654 368604 708042
rect 368004 693418 368186 693654
rect 368422 693418 368604 693654
rect 368004 693334 368604 693418
rect 368004 693098 368186 693334
rect 368422 693098 368604 693334
rect 368004 657654 368604 693098
rect 368004 657418 368186 657654
rect 368422 657418 368604 657654
rect 368004 657334 368604 657418
rect 368004 657098 368186 657334
rect 368422 657098 368604 657334
rect 368004 621654 368604 657098
rect 368004 621418 368186 621654
rect 368422 621418 368604 621654
rect 368004 621334 368604 621418
rect 368004 621098 368186 621334
rect 368422 621098 368604 621334
rect 368004 614247 368604 621098
rect 371604 697254 372204 709922
rect 389604 711418 390204 711440
rect 389604 711182 389786 711418
rect 390022 711182 390204 711418
rect 389604 711098 390204 711182
rect 389604 710862 389786 711098
rect 390022 710862 390204 711098
rect 386004 709538 386604 709560
rect 386004 709302 386186 709538
rect 386422 709302 386604 709538
rect 386004 709218 386604 709302
rect 386004 708982 386186 709218
rect 386422 708982 386604 709218
rect 382404 707658 383004 707680
rect 382404 707422 382586 707658
rect 382822 707422 383004 707658
rect 382404 707338 383004 707422
rect 382404 707102 382586 707338
rect 382822 707102 383004 707338
rect 371604 697018 371786 697254
rect 372022 697018 372204 697254
rect 371604 696934 372204 697018
rect 371604 696698 371786 696934
rect 372022 696698 372204 696934
rect 371604 661254 372204 696698
rect 371604 661018 371786 661254
rect 372022 661018 372204 661254
rect 371604 660934 372204 661018
rect 371604 660698 371786 660934
rect 372022 660698 372204 660934
rect 371604 625254 372204 660698
rect 371604 625018 371786 625254
rect 372022 625018 372204 625254
rect 371604 624934 372204 625018
rect 371604 624698 371786 624934
rect 372022 624698 372204 624934
rect 371604 614247 372204 624698
rect 378804 705778 379404 705800
rect 378804 705542 378986 705778
rect 379222 705542 379404 705778
rect 378804 705458 379404 705542
rect 378804 705222 378986 705458
rect 379222 705222 379404 705458
rect 378804 668454 379404 705222
rect 378804 668218 378986 668454
rect 379222 668218 379404 668454
rect 378804 668134 379404 668218
rect 378804 667898 378986 668134
rect 379222 667898 379404 668134
rect 378804 632454 379404 667898
rect 378804 632218 378986 632454
rect 379222 632218 379404 632454
rect 378804 632134 379404 632218
rect 378804 631898 378986 632134
rect 379222 631898 379404 632134
rect 378804 614247 379404 631898
rect 382404 672054 383004 707102
rect 382404 671818 382586 672054
rect 382822 671818 383004 672054
rect 382404 671734 383004 671818
rect 382404 671498 382586 671734
rect 382822 671498 383004 671734
rect 382404 636054 383004 671498
rect 382404 635818 382586 636054
rect 382822 635818 383004 636054
rect 382404 635734 383004 635818
rect 382404 635498 382586 635734
rect 382822 635498 383004 635734
rect 373579 612780 373645 612781
rect 373579 612716 373580 612780
rect 373644 612716 373645 612780
rect 373579 612715 373645 612716
rect 369163 611012 369229 611013
rect 369163 611010 369164 611012
rect 368608 610950 369164 611010
rect 369163 610948 369164 610950
rect 369228 610948 369229 611012
rect 369163 610947 369229 610948
rect 373027 611012 373093 611013
rect 373027 610948 373028 611012
rect 373092 611010 373093 611012
rect 373582 611010 373642 612715
rect 373092 610950 373642 611010
rect 373092 610948 373093 610950
rect 373027 610947 373093 610948
rect 382404 600054 383004 635498
rect 382404 599818 382586 600054
rect 382822 599818 383004 600054
rect 382404 599734 383004 599818
rect 382404 599498 382586 599734
rect 382822 599498 383004 599734
rect 376938 596454 377262 596476
rect 376938 596218 376982 596454
rect 377218 596218 377262 596454
rect 376938 596134 377262 596218
rect 376938 595898 376982 596134
rect 377218 595898 377262 596134
rect 376938 595876 377262 595898
rect 296004 585418 296186 585654
rect 296422 585418 296604 585654
rect 296004 585334 296604 585418
rect 296004 585098 296186 585334
rect 296422 585098 296604 585334
rect 296004 549654 296604 585098
rect 376494 578454 376814 578476
rect 376494 578218 376536 578454
rect 376772 578218 376814 578454
rect 376494 578134 376814 578218
rect 376494 577898 376536 578134
rect 376772 577898 376814 578134
rect 376494 577876 376814 577898
rect 382404 564054 383004 599498
rect 382404 563818 382586 564054
rect 382822 563818 383004 564054
rect 382404 563734 383004 563818
rect 382404 563498 382586 563734
rect 382822 563498 383004 563734
rect 376938 560454 377262 560476
rect 376938 560218 376982 560454
rect 377218 560218 377262 560454
rect 376938 560134 377262 560218
rect 376938 559898 376982 560134
rect 377218 559898 377262 560134
rect 376938 559876 377262 559898
rect 296004 549418 296186 549654
rect 296422 549418 296604 549654
rect 296004 549334 296604 549418
rect 296004 549098 296186 549334
rect 296422 549098 296604 549334
rect 296004 513654 296604 549098
rect 376494 542454 376814 542476
rect 376494 542218 376536 542454
rect 376772 542218 376814 542454
rect 376494 542134 376814 542218
rect 376494 541898 376536 542134
rect 376772 541898 376814 542134
rect 376494 541876 376814 541898
rect 382404 528054 383004 563498
rect 382404 527818 382586 528054
rect 382822 527818 383004 528054
rect 382404 527734 383004 527818
rect 382404 527498 382586 527734
rect 382822 527498 383004 527734
rect 376938 524454 377262 524476
rect 376938 524218 376982 524454
rect 377218 524218 377262 524454
rect 376938 524134 377262 524218
rect 376938 523898 376982 524134
rect 377218 523898 377262 524134
rect 376938 523876 377262 523898
rect 314702 520510 315008 520570
rect 316300 520510 316602 520570
rect 319804 520510 320098 520570
rect 303662 520170 303833 520230
rect 306832 520170 307402 520230
rect 308000 520170 308690 520230
rect 309168 520170 309794 520230
rect 303662 518261 303722 520170
rect 303659 518260 303725 518261
rect 303659 518196 303660 518260
rect 303724 518196 303725 518260
rect 303659 518195 303725 518196
rect 307342 517581 307402 520170
rect 308630 517581 308690 520170
rect 309734 517717 309794 520170
rect 309731 517716 309797 517717
rect 309731 517652 309732 517716
rect 309796 517652 309797 517716
rect 309731 517651 309797 517652
rect 310286 517581 310346 520230
rect 311504 520170 311818 520230
rect 311758 517581 311818 520170
rect 312494 520170 312672 520230
rect 312494 518669 312554 520170
rect 312766 519890 312826 520200
rect 312678 519830 312826 519890
rect 312491 518668 312557 518669
rect 312491 518604 312492 518668
rect 312556 518604 312557 518668
rect 312491 518603 312557 518604
rect 312678 517853 312738 519830
rect 313782 518805 313842 520230
rect 313964 520170 314026 520230
rect 313779 518804 313845 518805
rect 313779 518740 313780 518804
rect 313844 518740 313845 518804
rect 313779 518739 313845 518740
rect 313966 518397 314026 520170
rect 313963 518396 314029 518397
rect 313963 518332 313964 518396
rect 314028 518332 314029 518396
rect 313963 518331 314029 518332
rect 314702 518125 314762 520510
rect 315102 519890 315162 520200
rect 315070 519830 315162 519890
rect 316146 519890 316206 520200
rect 316146 519830 316234 519890
rect 315070 518533 315130 519830
rect 316174 518669 316234 519830
rect 316171 518668 316237 518669
rect 316171 518604 316172 518668
rect 316236 518604 316237 518668
rect 316171 518603 316237 518604
rect 316542 518533 316602 520510
rect 317278 520170 317344 520230
rect 317278 518533 317338 520170
rect 315067 518532 315133 518533
rect 315067 518468 315068 518532
rect 315132 518468 315133 518532
rect 315067 518467 315133 518468
rect 316539 518532 316605 518533
rect 316539 518468 316540 518532
rect 316604 518468 316605 518532
rect 316539 518467 316605 518468
rect 317275 518532 317341 518533
rect 317275 518468 317276 518532
rect 317340 518468 317341 518532
rect 317275 518467 317341 518468
rect 314699 518124 314765 518125
rect 314699 518060 314700 518124
rect 314764 518060 314765 518124
rect 314699 518059 314765 518060
rect 317462 517989 317522 520230
rect 318482 519890 318542 520200
rect 318636 520170 318810 520230
rect 318482 519830 318626 519890
rect 318566 518669 318626 519830
rect 318563 518668 318629 518669
rect 318563 518604 318564 518668
rect 318628 518604 318629 518668
rect 318563 518603 318629 518604
rect 318563 518532 318629 518533
rect 318563 518468 318564 518532
rect 318628 518530 318629 518532
rect 318750 518530 318810 520170
rect 319650 519890 319710 520200
rect 319650 519830 319730 519890
rect 319670 518805 319730 519830
rect 319667 518804 319733 518805
rect 319667 518740 319668 518804
rect 319732 518740 319733 518804
rect 319667 518739 319733 518740
rect 318628 518470 318810 518530
rect 318628 518468 318629 518470
rect 318563 518467 318629 518468
rect 320038 518125 320098 520510
rect 321694 520510 322016 520570
rect 323308 520510 323594 520570
rect 320774 520170 320848 520230
rect 320774 518669 320834 520170
rect 320771 518668 320837 518669
rect 320771 518604 320772 518668
rect 320836 518604 320837 518668
rect 320771 518603 320837 518604
rect 320958 518397 321018 520230
rect 321694 518533 321754 520510
rect 322110 519890 322170 520200
rect 322062 519830 322170 519890
rect 323154 519890 323214 520200
rect 323154 519830 323226 519890
rect 321691 518532 321757 518533
rect 321691 518468 321692 518532
rect 321756 518468 321757 518532
rect 321691 518467 321757 518468
rect 320955 518396 321021 518397
rect 320955 518332 320956 518396
rect 321020 518332 321021 518396
rect 320955 518331 321021 518332
rect 322062 518261 322122 519830
rect 323166 518669 323226 519830
rect 323534 518805 323594 520510
rect 325190 520510 325520 520570
rect 334574 520510 334864 520570
rect 338070 520510 338368 520570
rect 339660 520510 339970 520570
rect 324270 520170 324352 520230
rect 324270 518805 324330 520170
rect 323531 518804 323597 518805
rect 323531 518740 323532 518804
rect 323596 518740 323597 518804
rect 323531 518739 323597 518740
rect 324267 518804 324333 518805
rect 324267 518740 324268 518804
rect 324332 518740 324333 518804
rect 324267 518739 324333 518740
rect 323163 518668 323229 518669
rect 323163 518604 323164 518668
rect 323228 518604 323229 518668
rect 323163 518603 323229 518604
rect 322059 518260 322125 518261
rect 322059 518196 322060 518260
rect 322124 518196 322125 518260
rect 322059 518195 322125 518196
rect 320035 518124 320101 518125
rect 320035 518060 320036 518124
rect 320100 518060 320101 518124
rect 320035 518059 320101 518060
rect 317459 517988 317525 517989
rect 317459 517924 317460 517988
rect 317524 517924 317525 517988
rect 317459 517923 317525 517924
rect 312675 517852 312741 517853
rect 312675 517788 312676 517852
rect 312740 517788 312741 517852
rect 312675 517787 312741 517788
rect 324454 517717 324514 520230
rect 325190 518805 325250 520510
rect 325614 519890 325674 520200
rect 325558 519830 325674 519890
rect 326478 520170 326688 520230
rect 325187 518804 325253 518805
rect 325187 518740 325188 518804
rect 325252 518740 325253 518804
rect 325187 518739 325253 518740
rect 324451 517716 324517 517717
rect 324451 517652 324452 517716
rect 324516 517652 324517 517716
rect 324451 517651 324517 517652
rect 325558 517581 325618 519830
rect 326478 518805 326538 520170
rect 326782 519890 326842 520200
rect 326662 519830 326842 519890
rect 327398 520170 327856 520230
rect 326475 518804 326541 518805
rect 326475 518740 326476 518804
rect 326540 518740 326541 518804
rect 326475 518739 326541 518740
rect 326662 517717 326722 519830
rect 327398 518805 327458 520170
rect 327395 518804 327461 518805
rect 327395 518740 327396 518804
rect 327460 518740 327461 518804
rect 327395 518739 327461 518740
rect 327950 517717 328010 520200
rect 328870 520170 329024 520230
rect 328870 518805 328930 520170
rect 329118 519890 329178 520200
rect 329054 519830 329178 519890
rect 328867 518804 328933 518805
rect 328867 518740 328868 518804
rect 328932 518740 328933 518804
rect 328867 518739 328933 518740
rect 329054 517717 329114 519830
rect 330158 518805 330218 520230
rect 330316 520170 330402 520230
rect 330155 518804 330221 518805
rect 330155 518740 330156 518804
rect 330220 518740 330221 518804
rect 330155 518739 330221 518740
rect 330342 518533 330402 520170
rect 331330 519890 331390 520200
rect 331484 520170 331690 520230
rect 331262 519830 331390 519890
rect 331262 518669 331322 519830
rect 331630 518805 331690 520170
rect 332366 520170 332528 520230
rect 332366 518805 332426 520170
rect 332622 519890 332682 520200
rect 332550 519830 332682 519890
rect 331627 518804 331693 518805
rect 331627 518740 331628 518804
rect 331692 518740 331693 518804
rect 331627 518739 331693 518740
rect 332363 518804 332429 518805
rect 332363 518740 332364 518804
rect 332428 518740 332429 518804
rect 332363 518739 332429 518740
rect 331259 518668 331325 518669
rect 331259 518604 331260 518668
rect 331324 518604 331325 518668
rect 331259 518603 331325 518604
rect 330339 518532 330405 518533
rect 330339 518468 330340 518532
rect 330404 518468 330405 518532
rect 330339 518467 330405 518468
rect 332550 517717 332610 519830
rect 333654 518805 333714 520230
rect 333820 520170 333898 520230
rect 333651 518804 333717 518805
rect 333651 518740 333652 518804
rect 333716 518740 333717 518804
rect 333651 518739 333717 518740
rect 333838 518261 333898 520170
rect 334574 518805 334634 520510
rect 334958 519890 335018 520200
rect 334942 519830 335018 519890
rect 335862 520170 336032 520230
rect 334571 518804 334637 518805
rect 334571 518740 334572 518804
rect 334636 518740 334637 518804
rect 334571 518739 334637 518740
rect 333835 518260 333901 518261
rect 333835 518196 333836 518260
rect 333900 518196 333901 518260
rect 333835 518195 333901 518196
rect 334942 517853 335002 519830
rect 335862 518805 335922 520170
rect 336126 519890 336186 520200
rect 336046 519830 336186 519890
rect 336966 520170 337200 520230
rect 337324 520170 337394 520230
rect 335859 518804 335925 518805
rect 335859 518740 335860 518804
rect 335924 518740 335925 518804
rect 335859 518739 335925 518740
rect 334939 517852 335005 517853
rect 334939 517788 334940 517852
rect 335004 517788 335005 517852
rect 334939 517787 335005 517788
rect 336046 517717 336106 519830
rect 336966 518805 337026 520170
rect 336963 518804 337029 518805
rect 336963 518740 336964 518804
rect 337028 518740 337029 518804
rect 336963 518739 337029 518740
rect 337334 518397 337394 520170
rect 338070 518805 338130 520510
rect 338462 519890 338522 520200
rect 338438 519830 338522 519890
rect 339506 519890 339566 520200
rect 339506 519830 339602 519890
rect 338067 518804 338133 518805
rect 338067 518740 338068 518804
rect 338132 518740 338133 518804
rect 338067 518739 338133 518740
rect 338438 518397 338498 519830
rect 339542 518805 339602 519830
rect 339539 518804 339605 518805
rect 339539 518740 339540 518804
rect 339604 518740 339605 518804
rect 339539 518739 339605 518740
rect 339910 518397 339970 520510
rect 341566 520510 341872 520570
rect 343164 520510 343466 520570
rect 340462 520170 340704 520230
rect 340462 518805 340522 520170
rect 340798 519890 340858 520200
rect 340646 519830 340858 519890
rect 340459 518804 340525 518805
rect 340459 518740 340460 518804
rect 340524 518740 340525 518804
rect 340459 518739 340525 518740
rect 340646 518669 340706 519830
rect 341566 518805 341626 520510
rect 341966 519890 342026 520200
rect 341934 519830 342026 519890
rect 343010 519890 343070 520200
rect 343010 519830 343098 519890
rect 341563 518804 341629 518805
rect 341563 518740 341564 518804
rect 341628 518740 341629 518804
rect 341563 518739 341629 518740
rect 340643 518668 340709 518669
rect 340643 518604 340644 518668
rect 340708 518604 340709 518668
rect 340643 518603 340709 518604
rect 337331 518396 337397 518397
rect 337331 518332 337332 518396
rect 337396 518332 337397 518396
rect 337331 518331 337397 518332
rect 338435 518396 338501 518397
rect 338435 518332 338436 518396
rect 338500 518332 338501 518396
rect 338435 518331 338501 518332
rect 339907 518396 339973 518397
rect 339907 518332 339908 518396
rect 339972 518332 339973 518396
rect 339907 518331 339973 518332
rect 341934 518261 341994 519830
rect 343038 518533 343098 519830
rect 343035 518532 343101 518533
rect 343035 518468 343036 518532
rect 343100 518468 343101 518532
rect 343035 518467 343101 518468
rect 341931 518260 341997 518261
rect 341931 518196 341932 518260
rect 341996 518196 341997 518260
rect 341931 518195 341997 518196
rect 343406 517853 343466 520510
rect 343774 520170 344208 520230
rect 343774 518397 343834 520170
rect 343771 518396 343837 518397
rect 343771 518332 343772 518396
rect 343836 518332 343837 518396
rect 343771 518331 343837 518332
rect 343403 517852 343469 517853
rect 343403 517788 343404 517852
rect 343468 517788 343469 517852
rect 343403 517787 343469 517788
rect 344326 517717 344386 520230
rect 345062 520170 345376 520230
rect 345062 518805 345122 520170
rect 345470 519890 345530 520200
rect 345430 519830 345530 519890
rect 345059 518804 345125 518805
rect 345059 518740 345060 518804
rect 345124 518740 345125 518804
rect 345059 518739 345125 518740
rect 345430 517717 345490 519830
rect 346514 519210 346574 520200
rect 346638 519890 346698 520200
rect 347638 520170 347712 520230
rect 346638 519830 346778 519890
rect 346514 519150 346594 519210
rect 346534 518805 346594 519150
rect 346531 518804 346597 518805
rect 346531 518740 346532 518804
rect 346596 518740 346597 518804
rect 346531 518739 346597 518740
rect 346718 517717 346778 519830
rect 347638 518669 347698 520170
rect 347635 518668 347701 518669
rect 347635 518604 347636 518668
rect 347700 518604 347701 518668
rect 347635 518603 347701 518604
rect 347822 517853 347882 520230
rect 348850 519890 348910 520200
rect 349004 520170 349170 520230
rect 348850 519830 348986 519890
rect 348926 518805 348986 519830
rect 348923 518804 348989 518805
rect 348923 518740 348924 518804
rect 348988 518740 348989 518804
rect 348923 518739 348989 518740
rect 348923 518532 348989 518533
rect 348923 518468 348924 518532
rect 348988 518530 348989 518532
rect 349110 518530 349170 520170
rect 348988 518470 349170 518530
rect 348988 518468 348989 518470
rect 348923 518467 348989 518468
rect 347819 517852 347885 517853
rect 347819 517788 347820 517852
rect 347884 517788 347885 517852
rect 347819 517787 347885 517788
rect 326659 517716 326725 517717
rect 326659 517652 326660 517716
rect 326724 517652 326725 517716
rect 326659 517651 326725 517652
rect 327947 517716 328013 517717
rect 327947 517652 327948 517716
rect 328012 517652 328013 517716
rect 327947 517651 328013 517652
rect 329051 517716 329117 517717
rect 329051 517652 329052 517716
rect 329116 517652 329117 517716
rect 329051 517651 329117 517652
rect 332547 517716 332613 517717
rect 332547 517652 332548 517716
rect 332612 517652 332613 517716
rect 332547 517651 332613 517652
rect 336043 517716 336109 517717
rect 336043 517652 336044 517716
rect 336108 517652 336109 517716
rect 336043 517651 336109 517652
rect 344323 517716 344389 517717
rect 344323 517652 344324 517716
rect 344388 517652 344389 517716
rect 344323 517651 344389 517652
rect 345427 517716 345493 517717
rect 345427 517652 345428 517716
rect 345492 517652 345493 517716
rect 345427 517651 345493 517652
rect 346715 517716 346781 517717
rect 346715 517652 346716 517716
rect 346780 517652 346781 517716
rect 346715 517651 346781 517652
rect 307339 517580 307405 517581
rect 307339 517516 307340 517580
rect 307404 517516 307405 517580
rect 307339 517515 307405 517516
rect 308627 517580 308693 517581
rect 308627 517516 308628 517580
rect 308692 517516 308693 517580
rect 308627 517515 308693 517516
rect 310283 517580 310349 517581
rect 310283 517516 310284 517580
rect 310348 517516 310349 517580
rect 310283 517515 310349 517516
rect 311755 517580 311821 517581
rect 311755 517516 311756 517580
rect 311820 517516 311821 517580
rect 311755 517515 311821 517516
rect 325555 517580 325621 517581
rect 325555 517516 325556 517580
rect 325620 517516 325621 517580
rect 325555 517515 325621 517516
rect 296004 513418 296186 513654
rect 296422 513418 296604 513654
rect 296004 513334 296604 513418
rect 296004 513098 296186 513334
rect 296422 513098 296604 513334
rect 296004 483000 296604 513098
rect 299604 483000 300204 517000
rect 306804 488454 307404 517000
rect 306804 488218 306986 488454
rect 307222 488218 307404 488454
rect 306804 488134 307404 488218
rect 306804 487898 306986 488134
rect 307222 487898 307404 488134
rect 306804 483000 307404 487898
rect 310404 492054 311004 517000
rect 310404 491818 310586 492054
rect 310822 491818 311004 492054
rect 310404 491734 311004 491818
rect 310404 491498 310586 491734
rect 310822 491498 311004 491734
rect 310404 483000 311004 491498
rect 314004 495654 314604 517000
rect 314004 495418 314186 495654
rect 314422 495418 314604 495654
rect 314004 495334 314604 495418
rect 314004 495098 314186 495334
rect 314422 495098 314604 495334
rect 314004 483000 314604 495098
rect 317604 499254 318204 517000
rect 317604 499018 317786 499254
rect 318022 499018 318204 499254
rect 317604 498934 318204 499018
rect 317604 498698 317786 498934
rect 318022 498698 318204 498934
rect 317604 483000 318204 498698
rect 324804 506454 325404 517000
rect 324804 506218 324986 506454
rect 325222 506218 325404 506454
rect 324804 506134 325404 506218
rect 324804 505898 324986 506134
rect 325222 505898 325404 506134
rect 324804 483000 325404 505898
rect 328404 510054 329004 517000
rect 328404 509818 328586 510054
rect 328822 509818 329004 510054
rect 328404 509734 329004 509818
rect 328404 509498 328586 509734
rect 328822 509498 329004 509734
rect 328404 483000 329004 509498
rect 332004 513654 332604 517000
rect 332004 513418 332186 513654
rect 332422 513418 332604 513654
rect 332004 513334 332604 513418
rect 332004 513098 332186 513334
rect 332422 513098 332604 513334
rect 332004 483000 332604 513098
rect 335604 483000 336204 517000
rect 342804 488454 343404 517000
rect 342804 488218 342986 488454
rect 343222 488218 343404 488454
rect 342804 488134 343404 488218
rect 342804 487898 342986 488134
rect 343222 487898 343404 488134
rect 342804 483000 343404 487898
rect 346404 492054 347004 517000
rect 346404 491818 346586 492054
rect 346822 491818 347004 492054
rect 346404 491734 347004 491818
rect 346404 491498 346586 491734
rect 346822 491498 347004 491734
rect 346404 483000 347004 491498
rect 350004 495654 350604 517000
rect 350004 495418 350186 495654
rect 350422 495418 350604 495654
rect 350004 495334 350604 495418
rect 350004 495098 350186 495334
rect 350422 495098 350604 495334
rect 350004 483000 350604 495098
rect 353604 499254 354204 517000
rect 353604 499018 353786 499254
rect 354022 499018 354204 499254
rect 353604 498934 354204 499018
rect 353604 498698 353786 498934
rect 354022 498698 354204 498934
rect 353604 483000 354204 498698
rect 360804 506454 361404 517000
rect 360804 506218 360986 506454
rect 361222 506218 361404 506454
rect 360804 506134 361404 506218
rect 360804 505898 360986 506134
rect 361222 505898 361404 506134
rect 360804 483000 361404 505898
rect 364404 510054 365004 517000
rect 364404 509818 364586 510054
rect 364822 509818 365004 510054
rect 364404 509734 365004 509818
rect 364404 509498 364586 509734
rect 364822 509498 365004 509734
rect 364404 483000 365004 509498
rect 368004 513654 368604 517000
rect 368004 513418 368186 513654
rect 368422 513418 368604 513654
rect 368004 513334 368604 513418
rect 368004 513098 368186 513334
rect 368422 513098 368604 513334
rect 368004 483000 368604 513098
rect 371604 483000 372204 517000
rect 378804 488454 379404 517000
rect 378804 488218 378986 488454
rect 379222 488218 379404 488454
rect 378804 488134 379404 488218
rect 378804 487898 378986 488134
rect 379222 487898 379404 488134
rect 378804 483000 379404 487898
rect 382404 492054 383004 527498
rect 382404 491818 382586 492054
rect 382822 491818 383004 492054
rect 382404 491734 383004 491818
rect 382404 491498 382586 491734
rect 382822 491498 383004 491734
rect 382404 483000 383004 491498
rect 386004 675654 386604 708982
rect 386004 675418 386186 675654
rect 386422 675418 386604 675654
rect 386004 675334 386604 675418
rect 386004 675098 386186 675334
rect 386422 675098 386604 675334
rect 386004 639654 386604 675098
rect 386004 639418 386186 639654
rect 386422 639418 386604 639654
rect 386004 639334 386604 639418
rect 386004 639098 386186 639334
rect 386422 639098 386604 639334
rect 386004 603654 386604 639098
rect 386004 603418 386186 603654
rect 386422 603418 386604 603654
rect 386004 603334 386604 603418
rect 386004 603098 386186 603334
rect 386422 603098 386604 603334
rect 386004 567654 386604 603098
rect 386004 567418 386186 567654
rect 386422 567418 386604 567654
rect 386004 567334 386604 567418
rect 386004 567098 386186 567334
rect 386422 567098 386604 567334
rect 386004 531654 386604 567098
rect 386004 531418 386186 531654
rect 386422 531418 386604 531654
rect 386004 531334 386604 531418
rect 386004 531098 386186 531334
rect 386422 531098 386604 531334
rect 386004 495654 386604 531098
rect 386004 495418 386186 495654
rect 386422 495418 386604 495654
rect 386004 495334 386604 495418
rect 386004 495098 386186 495334
rect 386422 495098 386604 495334
rect 386004 483000 386604 495098
rect 389604 679254 390204 710862
rect 407604 710478 408204 711440
rect 407604 710242 407786 710478
rect 408022 710242 408204 710478
rect 407604 710158 408204 710242
rect 407604 709922 407786 710158
rect 408022 709922 408204 710158
rect 404004 708598 404604 709560
rect 404004 708362 404186 708598
rect 404422 708362 404604 708598
rect 404004 708278 404604 708362
rect 404004 708042 404186 708278
rect 404422 708042 404604 708278
rect 400404 706718 401004 707680
rect 400404 706482 400586 706718
rect 400822 706482 401004 706718
rect 400404 706398 401004 706482
rect 400404 706162 400586 706398
rect 400822 706162 401004 706398
rect 389604 679018 389786 679254
rect 390022 679018 390204 679254
rect 389604 678934 390204 679018
rect 389604 678698 389786 678934
rect 390022 678698 390204 678934
rect 389604 643254 390204 678698
rect 389604 643018 389786 643254
rect 390022 643018 390204 643254
rect 389604 642934 390204 643018
rect 389604 642698 389786 642934
rect 390022 642698 390204 642934
rect 389604 607254 390204 642698
rect 389604 607018 389786 607254
rect 390022 607018 390204 607254
rect 389604 606934 390204 607018
rect 389604 606698 389786 606934
rect 390022 606698 390204 606934
rect 389604 571254 390204 606698
rect 389604 571018 389786 571254
rect 390022 571018 390204 571254
rect 389604 570934 390204 571018
rect 389604 570698 389786 570934
rect 390022 570698 390204 570934
rect 389604 535254 390204 570698
rect 389604 535018 389786 535254
rect 390022 535018 390204 535254
rect 389604 534934 390204 535018
rect 389604 534698 389786 534934
rect 390022 534698 390204 534934
rect 389604 499254 390204 534698
rect 389604 499018 389786 499254
rect 390022 499018 390204 499254
rect 389604 498934 390204 499018
rect 389604 498698 389786 498934
rect 390022 498698 390204 498934
rect 389604 483000 390204 498698
rect 396804 704838 397404 705800
rect 396804 704602 396986 704838
rect 397222 704602 397404 704838
rect 396804 704518 397404 704602
rect 396804 704282 396986 704518
rect 397222 704282 397404 704518
rect 396804 686454 397404 704282
rect 396804 686218 396986 686454
rect 397222 686218 397404 686454
rect 396804 686134 397404 686218
rect 396804 685898 396986 686134
rect 397222 685898 397404 686134
rect 396804 650454 397404 685898
rect 396804 650218 396986 650454
rect 397222 650218 397404 650454
rect 396804 650134 397404 650218
rect 396804 649898 396986 650134
rect 397222 649898 397404 650134
rect 396804 614454 397404 649898
rect 396804 614218 396986 614454
rect 397222 614218 397404 614454
rect 396804 614134 397404 614218
rect 396804 613898 396986 614134
rect 397222 613898 397404 614134
rect 396804 578454 397404 613898
rect 396804 578218 396986 578454
rect 397222 578218 397404 578454
rect 396804 578134 397404 578218
rect 396804 577898 396986 578134
rect 397222 577898 397404 578134
rect 396804 542454 397404 577898
rect 396804 542218 396986 542454
rect 397222 542218 397404 542454
rect 396804 542134 397404 542218
rect 396804 541898 396986 542134
rect 397222 541898 397404 542134
rect 396804 506454 397404 541898
rect 396804 506218 396986 506454
rect 397222 506218 397404 506454
rect 396804 506134 397404 506218
rect 396804 505898 396986 506134
rect 397222 505898 397404 506134
rect 396804 483000 397404 505898
rect 400404 690054 401004 706162
rect 400404 689818 400586 690054
rect 400822 689818 401004 690054
rect 400404 689734 401004 689818
rect 400404 689498 400586 689734
rect 400822 689498 401004 689734
rect 400404 654054 401004 689498
rect 400404 653818 400586 654054
rect 400822 653818 401004 654054
rect 400404 653734 401004 653818
rect 400404 653498 400586 653734
rect 400822 653498 401004 653734
rect 400404 618054 401004 653498
rect 400404 617818 400586 618054
rect 400822 617818 401004 618054
rect 400404 617734 401004 617818
rect 400404 617498 400586 617734
rect 400822 617498 401004 617734
rect 400404 582054 401004 617498
rect 400404 581818 400586 582054
rect 400822 581818 401004 582054
rect 400404 581734 401004 581818
rect 400404 581498 400586 581734
rect 400822 581498 401004 581734
rect 400404 546054 401004 581498
rect 400404 545818 400586 546054
rect 400822 545818 401004 546054
rect 400404 545734 401004 545818
rect 400404 545498 400586 545734
rect 400822 545498 401004 545734
rect 400404 510054 401004 545498
rect 400404 509818 400586 510054
rect 400822 509818 401004 510054
rect 400404 509734 401004 509818
rect 400404 509498 400586 509734
rect 400822 509498 401004 509734
rect 400404 483000 401004 509498
rect 404004 693654 404604 708042
rect 404004 693418 404186 693654
rect 404422 693418 404604 693654
rect 404004 693334 404604 693418
rect 404004 693098 404186 693334
rect 404422 693098 404604 693334
rect 404004 657654 404604 693098
rect 404004 657418 404186 657654
rect 404422 657418 404604 657654
rect 404004 657334 404604 657418
rect 404004 657098 404186 657334
rect 404422 657098 404604 657334
rect 404004 621654 404604 657098
rect 404004 621418 404186 621654
rect 404422 621418 404604 621654
rect 404004 621334 404604 621418
rect 404004 621098 404186 621334
rect 404422 621098 404604 621334
rect 404004 585654 404604 621098
rect 404004 585418 404186 585654
rect 404422 585418 404604 585654
rect 404004 585334 404604 585418
rect 404004 585098 404186 585334
rect 404422 585098 404604 585334
rect 404004 549654 404604 585098
rect 404004 549418 404186 549654
rect 404422 549418 404604 549654
rect 404004 549334 404604 549418
rect 404004 549098 404186 549334
rect 404422 549098 404604 549334
rect 404004 513654 404604 549098
rect 404004 513418 404186 513654
rect 404422 513418 404604 513654
rect 404004 513334 404604 513418
rect 404004 513098 404186 513334
rect 404422 513098 404604 513334
rect 404004 483000 404604 513098
rect 407604 697254 408204 709922
rect 425604 711418 426204 711440
rect 425604 711182 425786 711418
rect 426022 711182 426204 711418
rect 425604 711098 426204 711182
rect 425604 710862 425786 711098
rect 426022 710862 426204 711098
rect 422004 709538 422604 709560
rect 422004 709302 422186 709538
rect 422422 709302 422604 709538
rect 422004 709218 422604 709302
rect 422004 708982 422186 709218
rect 422422 708982 422604 709218
rect 418404 707658 419004 707680
rect 418404 707422 418586 707658
rect 418822 707422 419004 707658
rect 418404 707338 419004 707422
rect 418404 707102 418586 707338
rect 418822 707102 419004 707338
rect 407604 697018 407786 697254
rect 408022 697018 408204 697254
rect 407604 696934 408204 697018
rect 407604 696698 407786 696934
rect 408022 696698 408204 696934
rect 407604 661254 408204 696698
rect 407604 661018 407786 661254
rect 408022 661018 408204 661254
rect 407604 660934 408204 661018
rect 407604 660698 407786 660934
rect 408022 660698 408204 660934
rect 407604 625254 408204 660698
rect 407604 625018 407786 625254
rect 408022 625018 408204 625254
rect 407604 624934 408204 625018
rect 407604 624698 407786 624934
rect 408022 624698 408204 624934
rect 407604 589254 408204 624698
rect 407604 589018 407786 589254
rect 408022 589018 408204 589254
rect 407604 588934 408204 589018
rect 407604 588698 407786 588934
rect 408022 588698 408204 588934
rect 407604 553254 408204 588698
rect 407604 553018 407786 553254
rect 408022 553018 408204 553254
rect 407604 552934 408204 553018
rect 407604 552698 407786 552934
rect 408022 552698 408204 552934
rect 407604 517254 408204 552698
rect 407604 517018 407786 517254
rect 408022 517018 408204 517254
rect 407604 516934 408204 517018
rect 407604 516698 407786 516934
rect 408022 516698 408204 516934
rect 407604 483000 408204 516698
rect 414804 705778 415404 705800
rect 414804 705542 414986 705778
rect 415222 705542 415404 705778
rect 414804 705458 415404 705542
rect 414804 705222 414986 705458
rect 415222 705222 415404 705458
rect 414804 668454 415404 705222
rect 414804 668218 414986 668454
rect 415222 668218 415404 668454
rect 414804 668134 415404 668218
rect 414804 667898 414986 668134
rect 415222 667898 415404 668134
rect 414804 632454 415404 667898
rect 414804 632218 414986 632454
rect 415222 632218 415404 632454
rect 414804 632134 415404 632218
rect 414804 631898 414986 632134
rect 415222 631898 415404 632134
rect 414804 596454 415404 631898
rect 418404 672054 419004 707102
rect 418404 671818 418586 672054
rect 418822 671818 419004 672054
rect 418404 671734 419004 671818
rect 418404 671498 418586 671734
rect 418822 671498 419004 671734
rect 418404 636054 419004 671498
rect 418404 635818 418586 636054
rect 418822 635818 419004 636054
rect 418404 635734 419004 635818
rect 418404 635498 418586 635734
rect 418822 635498 419004 635734
rect 418404 614247 419004 635498
rect 422004 675654 422604 708982
rect 422004 675418 422186 675654
rect 422422 675418 422604 675654
rect 422004 675334 422604 675418
rect 422004 675098 422186 675334
rect 422422 675098 422604 675334
rect 422004 639654 422604 675098
rect 422004 639418 422186 639654
rect 422422 639418 422604 639654
rect 422004 639334 422604 639418
rect 422004 639098 422186 639334
rect 422422 639098 422604 639334
rect 422004 614247 422604 639098
rect 425604 679254 426204 710862
rect 443604 710478 444204 711440
rect 443604 710242 443786 710478
rect 444022 710242 444204 710478
rect 443604 710158 444204 710242
rect 443604 709922 443786 710158
rect 444022 709922 444204 710158
rect 440004 708598 440604 709560
rect 440004 708362 440186 708598
rect 440422 708362 440604 708598
rect 440004 708278 440604 708362
rect 440004 708042 440186 708278
rect 440422 708042 440604 708278
rect 436404 706718 437004 707680
rect 436404 706482 436586 706718
rect 436822 706482 437004 706718
rect 436404 706398 437004 706482
rect 436404 706162 436586 706398
rect 436822 706162 437004 706398
rect 425604 679018 425786 679254
rect 426022 679018 426204 679254
rect 425604 678934 426204 679018
rect 425604 678698 425786 678934
rect 426022 678698 426204 678934
rect 425604 643254 426204 678698
rect 425604 643018 425786 643254
rect 426022 643018 426204 643254
rect 425604 642934 426204 643018
rect 425604 642698 425786 642934
rect 426022 642698 426204 642934
rect 425604 614247 426204 642698
rect 432804 704838 433404 705800
rect 432804 704602 432986 704838
rect 433222 704602 433404 704838
rect 432804 704518 433404 704602
rect 432804 704282 432986 704518
rect 433222 704282 433404 704518
rect 432804 686454 433404 704282
rect 432804 686218 432986 686454
rect 433222 686218 433404 686454
rect 432804 686134 433404 686218
rect 432804 685898 432986 686134
rect 433222 685898 433404 686134
rect 432804 650454 433404 685898
rect 432804 650218 432986 650454
rect 433222 650218 433404 650454
rect 432804 650134 433404 650218
rect 432804 649898 432986 650134
rect 433222 649898 433404 650134
rect 432804 614247 433404 649898
rect 436404 690054 437004 706162
rect 436404 689818 436586 690054
rect 436822 689818 437004 690054
rect 436404 689734 437004 689818
rect 436404 689498 436586 689734
rect 436822 689498 437004 689734
rect 436404 654054 437004 689498
rect 436404 653818 436586 654054
rect 436822 653818 437004 654054
rect 436404 653734 437004 653818
rect 436404 653498 436586 653734
rect 436822 653498 437004 653734
rect 436404 618054 437004 653498
rect 436404 617818 436586 618054
rect 436822 617818 437004 618054
rect 436404 617734 437004 617818
rect 436404 617498 436586 617734
rect 436822 617498 437004 617734
rect 436404 614247 437004 617498
rect 440004 693654 440604 708042
rect 440004 693418 440186 693654
rect 440422 693418 440604 693654
rect 440004 693334 440604 693418
rect 440004 693098 440186 693334
rect 440422 693098 440604 693334
rect 440004 657654 440604 693098
rect 440004 657418 440186 657654
rect 440422 657418 440604 657654
rect 440004 657334 440604 657418
rect 440004 657098 440186 657334
rect 440422 657098 440604 657334
rect 440004 621654 440604 657098
rect 440004 621418 440186 621654
rect 440422 621418 440604 621654
rect 440004 621334 440604 621418
rect 440004 621098 440186 621334
rect 440422 621098 440604 621334
rect 440004 614247 440604 621098
rect 443604 697254 444204 709922
rect 461604 711418 462204 711440
rect 461604 711182 461786 711418
rect 462022 711182 462204 711418
rect 461604 711098 462204 711182
rect 461604 710862 461786 711098
rect 462022 710862 462204 711098
rect 458004 709538 458604 709560
rect 458004 709302 458186 709538
rect 458422 709302 458604 709538
rect 458004 709218 458604 709302
rect 458004 708982 458186 709218
rect 458422 708982 458604 709218
rect 454404 707658 455004 707680
rect 454404 707422 454586 707658
rect 454822 707422 455004 707658
rect 454404 707338 455004 707422
rect 454404 707102 454586 707338
rect 454822 707102 455004 707338
rect 443604 697018 443786 697254
rect 444022 697018 444204 697254
rect 443604 696934 444204 697018
rect 443604 696698 443786 696934
rect 444022 696698 444204 696934
rect 443604 661254 444204 696698
rect 443604 661018 443786 661254
rect 444022 661018 444204 661254
rect 443604 660934 444204 661018
rect 443604 660698 443786 660934
rect 444022 660698 444204 660934
rect 443604 625254 444204 660698
rect 443604 625018 443786 625254
rect 444022 625018 444204 625254
rect 443604 624934 444204 625018
rect 443604 624698 443786 624934
rect 444022 624698 444204 624934
rect 443604 614247 444204 624698
rect 450804 705778 451404 705800
rect 450804 705542 450986 705778
rect 451222 705542 451404 705778
rect 450804 705458 451404 705542
rect 450804 705222 450986 705458
rect 451222 705222 451404 705458
rect 450804 668454 451404 705222
rect 450804 668218 450986 668454
rect 451222 668218 451404 668454
rect 450804 668134 451404 668218
rect 450804 667898 450986 668134
rect 451222 667898 451404 668134
rect 450804 632454 451404 667898
rect 450804 632218 450986 632454
rect 451222 632218 451404 632454
rect 450804 632134 451404 632218
rect 450804 631898 450986 632134
rect 451222 631898 451404 632134
rect 450804 614247 451404 631898
rect 454404 672054 455004 707102
rect 454404 671818 454586 672054
rect 454822 671818 455004 672054
rect 454404 671734 455004 671818
rect 454404 671498 454586 671734
rect 454822 671498 455004 671734
rect 454404 636054 455004 671498
rect 454404 635818 454586 636054
rect 454822 635818 455004 636054
rect 454404 635734 455004 635818
rect 454404 635498 454586 635734
rect 454822 635498 455004 635734
rect 454404 614247 455004 635498
rect 458004 675654 458604 708982
rect 458004 675418 458186 675654
rect 458422 675418 458604 675654
rect 458004 675334 458604 675418
rect 458004 675098 458186 675334
rect 458422 675098 458604 675334
rect 458004 639654 458604 675098
rect 458004 639418 458186 639654
rect 458422 639418 458604 639654
rect 458004 639334 458604 639418
rect 458004 639098 458186 639334
rect 458422 639098 458604 639334
rect 458004 614247 458604 639098
rect 461604 679254 462204 710862
rect 479604 710478 480204 711440
rect 479604 710242 479786 710478
rect 480022 710242 480204 710478
rect 479604 710158 480204 710242
rect 479604 709922 479786 710158
rect 480022 709922 480204 710158
rect 476004 708598 476604 709560
rect 476004 708362 476186 708598
rect 476422 708362 476604 708598
rect 476004 708278 476604 708362
rect 476004 708042 476186 708278
rect 476422 708042 476604 708278
rect 472404 706718 473004 707680
rect 472404 706482 472586 706718
rect 472822 706482 473004 706718
rect 472404 706398 473004 706482
rect 472404 706162 472586 706398
rect 472822 706162 473004 706398
rect 461604 679018 461786 679254
rect 462022 679018 462204 679254
rect 461604 678934 462204 679018
rect 461604 678698 461786 678934
rect 462022 678698 462204 678934
rect 461604 643254 462204 678698
rect 461604 643018 461786 643254
rect 462022 643018 462204 643254
rect 461604 642934 462204 643018
rect 461604 642698 461786 642934
rect 462022 642698 462204 642934
rect 461604 614247 462204 642698
rect 468804 704838 469404 705800
rect 468804 704602 468986 704838
rect 469222 704602 469404 704838
rect 468804 704518 469404 704602
rect 468804 704282 468986 704518
rect 469222 704282 469404 704518
rect 468804 686454 469404 704282
rect 468804 686218 468986 686454
rect 469222 686218 469404 686454
rect 468804 686134 469404 686218
rect 468804 685898 468986 686134
rect 469222 685898 469404 686134
rect 468804 650454 469404 685898
rect 468804 650218 468986 650454
rect 469222 650218 469404 650454
rect 468804 650134 469404 650218
rect 468804 649898 468986 650134
rect 469222 649898 469404 650134
rect 468804 614247 469404 649898
rect 472404 690054 473004 706162
rect 472404 689818 472586 690054
rect 472822 689818 473004 690054
rect 472404 689734 473004 689818
rect 472404 689498 472586 689734
rect 472822 689498 473004 689734
rect 472404 654054 473004 689498
rect 472404 653818 472586 654054
rect 472822 653818 473004 654054
rect 472404 653734 473004 653818
rect 472404 653498 472586 653734
rect 472822 653498 473004 653734
rect 472404 618054 473004 653498
rect 472404 617818 472586 618054
rect 472822 617818 473004 618054
rect 472404 617734 473004 617818
rect 472404 617498 472586 617734
rect 472822 617498 473004 617734
rect 472404 614247 473004 617498
rect 476004 693654 476604 708042
rect 476004 693418 476186 693654
rect 476422 693418 476604 693654
rect 476004 693334 476604 693418
rect 476004 693098 476186 693334
rect 476422 693098 476604 693334
rect 476004 657654 476604 693098
rect 476004 657418 476186 657654
rect 476422 657418 476604 657654
rect 476004 657334 476604 657418
rect 476004 657098 476186 657334
rect 476422 657098 476604 657334
rect 476004 621654 476604 657098
rect 476004 621418 476186 621654
rect 476422 621418 476604 621654
rect 476004 621334 476604 621418
rect 476004 621098 476186 621334
rect 476422 621098 476604 621334
rect 476004 614247 476604 621098
rect 479604 697254 480204 709922
rect 497604 711418 498204 711440
rect 497604 711182 497786 711418
rect 498022 711182 498204 711418
rect 497604 711098 498204 711182
rect 497604 710862 497786 711098
rect 498022 710862 498204 711098
rect 494004 709538 494604 709560
rect 494004 709302 494186 709538
rect 494422 709302 494604 709538
rect 494004 709218 494604 709302
rect 494004 708982 494186 709218
rect 494422 708982 494604 709218
rect 490404 707658 491004 707680
rect 490404 707422 490586 707658
rect 490822 707422 491004 707658
rect 490404 707338 491004 707422
rect 490404 707102 490586 707338
rect 490822 707102 491004 707338
rect 479604 697018 479786 697254
rect 480022 697018 480204 697254
rect 479604 696934 480204 697018
rect 479604 696698 479786 696934
rect 480022 696698 480204 696934
rect 479604 661254 480204 696698
rect 479604 661018 479786 661254
rect 480022 661018 480204 661254
rect 479604 660934 480204 661018
rect 479604 660698 479786 660934
rect 480022 660698 480204 660934
rect 479604 625254 480204 660698
rect 479604 625018 479786 625254
rect 480022 625018 480204 625254
rect 479604 624934 480204 625018
rect 479604 624698 479786 624934
rect 480022 624698 480204 624934
rect 479604 614247 480204 624698
rect 486804 705778 487404 705800
rect 486804 705542 486986 705778
rect 487222 705542 487404 705778
rect 486804 705458 487404 705542
rect 486804 705222 486986 705458
rect 487222 705222 487404 705458
rect 486804 668454 487404 705222
rect 486804 668218 486986 668454
rect 487222 668218 487404 668454
rect 486804 668134 487404 668218
rect 486804 667898 486986 668134
rect 487222 667898 487404 668134
rect 486804 632454 487404 667898
rect 486804 632218 486986 632454
rect 487222 632218 487404 632454
rect 486804 632134 487404 632218
rect 486804 631898 486986 632134
rect 487222 631898 487404 632134
rect 486804 614247 487404 631898
rect 490404 672054 491004 707102
rect 490404 671818 490586 672054
rect 490822 671818 491004 672054
rect 490404 671734 491004 671818
rect 490404 671498 490586 671734
rect 490822 671498 491004 671734
rect 490404 636054 491004 671498
rect 490404 635818 490586 636054
rect 490822 635818 491004 636054
rect 490404 635734 491004 635818
rect 490404 635498 490586 635734
rect 490822 635498 491004 635734
rect 490404 614247 491004 635498
rect 494004 675654 494604 708982
rect 494004 675418 494186 675654
rect 494422 675418 494604 675654
rect 494004 675334 494604 675418
rect 494004 675098 494186 675334
rect 494422 675098 494604 675334
rect 494004 639654 494604 675098
rect 494004 639418 494186 639654
rect 494422 639418 494604 639654
rect 494004 639334 494604 639418
rect 494004 639098 494186 639334
rect 494422 639098 494604 639334
rect 494004 614247 494604 639098
rect 497604 679254 498204 710862
rect 515604 710478 516204 711440
rect 515604 710242 515786 710478
rect 516022 710242 516204 710478
rect 515604 710158 516204 710242
rect 515604 709922 515786 710158
rect 516022 709922 516204 710158
rect 512004 708598 512604 709560
rect 512004 708362 512186 708598
rect 512422 708362 512604 708598
rect 512004 708278 512604 708362
rect 512004 708042 512186 708278
rect 512422 708042 512604 708278
rect 508404 706718 509004 707680
rect 508404 706482 508586 706718
rect 508822 706482 509004 706718
rect 508404 706398 509004 706482
rect 508404 706162 508586 706398
rect 508822 706162 509004 706398
rect 497604 679018 497786 679254
rect 498022 679018 498204 679254
rect 497604 678934 498204 679018
rect 497604 678698 497786 678934
rect 498022 678698 498204 678934
rect 497604 643254 498204 678698
rect 497604 643018 497786 643254
rect 498022 643018 498204 643254
rect 497604 642934 498204 643018
rect 497604 642698 497786 642934
rect 498022 642698 498204 642934
rect 497604 614247 498204 642698
rect 504804 704838 505404 705800
rect 504804 704602 504986 704838
rect 505222 704602 505404 704838
rect 504804 704518 505404 704602
rect 504804 704282 504986 704518
rect 505222 704282 505404 704518
rect 504804 686454 505404 704282
rect 504804 686218 504986 686454
rect 505222 686218 505404 686454
rect 504804 686134 505404 686218
rect 504804 685898 504986 686134
rect 505222 685898 505404 686134
rect 504804 650454 505404 685898
rect 504804 650218 504986 650454
rect 505222 650218 505404 650454
rect 504804 650134 505404 650218
rect 504804 649898 504986 650134
rect 505222 649898 505404 650134
rect 504804 614454 505404 649898
rect 504804 614218 504986 614454
rect 505222 614218 505404 614454
rect 504804 614134 505404 614218
rect 504804 613898 504986 614134
rect 505222 613898 505404 614134
rect 488579 612780 488645 612781
rect 488579 612716 488580 612780
rect 488644 612716 488645 612780
rect 488579 612715 488645 612716
rect 493915 612780 493981 612781
rect 493915 612716 493916 612780
rect 493980 612716 493981 612780
rect 493915 612715 493981 612716
rect 488582 610950 488642 612715
rect 493918 611010 493978 612715
rect 493603 610950 493978 611010
rect 414804 596218 414986 596454
rect 415222 596218 415404 596454
rect 414804 596134 415404 596218
rect 414804 595898 414986 596134
rect 415222 595898 415404 596134
rect 414804 560454 415404 595898
rect 496938 596454 497262 596476
rect 496938 596218 496982 596454
rect 497218 596218 497262 596454
rect 496938 596134 497262 596218
rect 496938 595898 496982 596134
rect 497218 595898 497262 596134
rect 496938 595876 497262 595898
rect 496494 578454 496814 578476
rect 496494 578218 496536 578454
rect 496772 578218 496814 578454
rect 496494 578134 496814 578218
rect 496494 577898 496536 578134
rect 496772 577898 496814 578134
rect 496494 577876 496814 577898
rect 504804 578454 505404 613898
rect 504804 578218 504986 578454
rect 505222 578218 505404 578454
rect 504804 578134 505404 578218
rect 504804 577898 504986 578134
rect 505222 577898 505404 578134
rect 414804 560218 414986 560454
rect 415222 560218 415404 560454
rect 414804 560134 415404 560218
rect 414804 559898 414986 560134
rect 415222 559898 415404 560134
rect 414804 524454 415404 559898
rect 496938 560454 497262 560476
rect 496938 560218 496982 560454
rect 497218 560218 497262 560454
rect 496938 560134 497262 560218
rect 496938 559898 496982 560134
rect 497218 559898 497262 560134
rect 496938 559876 497262 559898
rect 496494 542454 496814 542476
rect 496494 542218 496536 542454
rect 496772 542218 496814 542454
rect 496494 542134 496814 542218
rect 496494 541898 496536 542134
rect 496772 541898 496814 542134
rect 496494 541876 496814 541898
rect 504804 542454 505404 577898
rect 504804 542218 504986 542454
rect 505222 542218 505404 542454
rect 504804 542134 505404 542218
rect 504804 541898 504986 542134
rect 505222 541898 505404 542134
rect 414804 524218 414986 524454
rect 415222 524218 415404 524454
rect 414804 524134 415404 524218
rect 414804 523898 414986 524134
rect 415222 523898 415404 524134
rect 414804 488454 415404 523898
rect 496938 524454 497262 524476
rect 496938 524218 496982 524454
rect 497218 524218 497262 524454
rect 496938 524134 497262 524218
rect 496938 523898 496982 524134
rect 497218 523898 497262 524134
rect 496938 523876 497262 523898
rect 423814 518261 423874 520230
rect 426574 520170 426832 520230
rect 426574 518533 426634 520170
rect 427970 519757 428030 520200
rect 427967 519756 428033 519757
rect 427967 519692 427968 519756
rect 428032 519692 428033 519756
rect 427967 519691 428033 519692
rect 426571 518532 426637 518533
rect 426571 518468 426572 518532
rect 426636 518468 426637 518532
rect 426571 518467 426637 518468
rect 429150 518261 429210 520230
rect 429702 520170 430336 520230
rect 430806 520170 431504 520230
rect 429702 518669 429762 520170
rect 429699 518668 429765 518669
rect 429699 518604 429700 518668
rect 429764 518604 429765 518668
rect 429699 518603 429765 518604
rect 430806 518397 430866 520170
rect 432642 519890 432702 520200
rect 432796 520170 433074 520230
rect 432642 519830 432706 519890
rect 430803 518396 430869 518397
rect 430803 518332 430804 518396
rect 430868 518332 430869 518396
rect 430803 518331 430869 518332
rect 423811 518260 423877 518261
rect 423811 518196 423812 518260
rect 423876 518196 423877 518260
rect 423811 518195 423877 518196
rect 429147 518260 429213 518261
rect 429147 518196 429148 518260
rect 429212 518196 429213 518260
rect 429147 518195 429213 518196
rect 432646 517853 432706 519830
rect 432643 517852 432709 517853
rect 432643 517788 432644 517852
rect 432708 517788 432709 517852
rect 432643 517787 432709 517788
rect 433014 517717 433074 520170
rect 433810 519757 433870 520200
rect 433807 519756 433873 519757
rect 433807 519692 433808 519756
rect 433872 519692 433873 519756
rect 433807 519691 433873 519692
rect 433934 517717 433994 520200
rect 434978 519890 435038 520200
rect 435132 520170 435834 520230
rect 434978 519830 435098 519890
rect 435038 518397 435098 519830
rect 435035 518396 435101 518397
rect 435035 518332 435036 518396
rect 435100 518332 435101 518396
rect 435035 518331 435101 518332
rect 435774 517717 435834 520170
rect 436142 518261 436202 520230
rect 436300 520170 436938 520230
rect 436139 518260 436205 518261
rect 436139 518196 436140 518260
rect 436204 518196 436205 518260
rect 436139 518195 436205 518196
rect 436878 517717 436938 520170
rect 437314 519890 437374 520200
rect 437468 520170 438042 520230
rect 437246 519830 437374 519890
rect 437246 517853 437306 519830
rect 437243 517852 437309 517853
rect 437243 517788 437244 517852
rect 437308 517788 437309 517852
rect 437243 517787 437309 517788
rect 437982 517717 438042 520170
rect 438350 520170 438512 520230
rect 433011 517716 433077 517717
rect 433011 517652 433012 517716
rect 433076 517652 433077 517716
rect 433011 517651 433077 517652
rect 433931 517716 433997 517717
rect 433931 517652 433932 517716
rect 433996 517652 433997 517716
rect 433931 517651 433997 517652
rect 435771 517716 435837 517717
rect 435771 517652 435772 517716
rect 435836 517652 435837 517716
rect 435771 517651 435837 517652
rect 436875 517716 436941 517717
rect 436875 517652 436876 517716
rect 436940 517652 436941 517716
rect 436875 517651 436941 517652
rect 437979 517716 438045 517717
rect 437979 517652 437980 517716
rect 438044 517652 438045 517716
rect 437979 517651 438045 517652
rect 438350 517581 438410 520170
rect 438606 519890 438666 520200
rect 438606 519830 438778 519890
rect 438718 517581 438778 519830
rect 439638 517581 439698 520230
rect 439804 520170 440066 520230
rect 440006 517581 440066 520170
rect 440818 519890 440878 520200
rect 440972 520170 441538 520230
rect 440742 519830 440878 519890
rect 440742 518261 440802 519830
rect 440739 518260 440805 518261
rect 440739 518196 440740 518260
rect 440804 518196 440805 518260
rect 440739 518195 440805 518196
rect 441478 517581 441538 520170
rect 441662 520170 442016 520230
rect 442140 520170 442826 520230
rect 441662 518669 441722 520170
rect 441659 518668 441725 518669
rect 441659 518604 441660 518668
rect 441724 518604 441725 518668
rect 441659 518603 441725 518604
rect 442766 517581 442826 520170
rect 443134 518805 443194 520230
rect 443308 520170 443930 520230
rect 443131 518804 443197 518805
rect 443131 518740 443132 518804
rect 443196 518740 443197 518804
rect 443131 518739 443197 518740
rect 443870 518533 443930 520170
rect 444054 520170 444352 520230
rect 444476 520170 445034 520230
rect 444054 518669 444114 520170
rect 444051 518668 444117 518669
rect 444051 518604 444052 518668
rect 444116 518604 444117 518668
rect 444051 518603 444117 518604
rect 444974 518533 445034 520170
rect 445342 520170 445520 520230
rect 445342 518669 445402 520170
rect 445614 519890 445674 520200
rect 445526 519830 445674 519890
rect 445339 518668 445405 518669
rect 445339 518604 445340 518668
rect 445404 518604 445405 518668
rect 445339 518603 445405 518604
rect 443867 518532 443933 518533
rect 443867 518468 443868 518532
rect 443932 518468 443933 518532
rect 443867 518467 443933 518468
rect 444971 518532 445037 518533
rect 444971 518468 444972 518532
rect 445036 518468 445037 518532
rect 444971 518467 445037 518468
rect 445526 518397 445586 519830
rect 446630 518669 446690 520230
rect 446812 520170 447058 520230
rect 446627 518668 446693 518669
rect 446627 518604 446628 518668
rect 446692 518604 446693 518668
rect 446627 518603 446693 518604
rect 446998 518397 447058 520170
rect 447826 519890 447886 520200
rect 447980 520170 448346 520230
rect 447734 519830 447886 519890
rect 447734 518533 447794 519830
rect 447731 518532 447797 518533
rect 447731 518468 447732 518532
rect 447796 518468 447797 518532
rect 447731 518467 447797 518468
rect 445523 518396 445589 518397
rect 445523 518332 445524 518396
rect 445588 518332 445589 518396
rect 445523 518331 445589 518332
rect 446995 518396 447061 518397
rect 446995 518332 446996 518396
rect 447060 518332 447061 518396
rect 446995 518331 447061 518332
rect 448286 518261 448346 520170
rect 448838 520170 449024 520230
rect 449148 520170 449818 520230
rect 448838 518533 448898 520170
rect 448835 518532 448901 518533
rect 448835 518468 448836 518532
rect 448900 518468 448901 518532
rect 448835 518467 448901 518468
rect 448283 518260 448349 518261
rect 448283 518196 448284 518260
rect 448348 518196 448349 518260
rect 448283 518195 448349 518196
rect 449758 517581 449818 520170
rect 450126 520170 450192 520230
rect 450316 520170 450922 520230
rect 450126 518397 450186 520170
rect 450123 518396 450189 518397
rect 450123 518332 450124 518396
rect 450188 518332 450189 518396
rect 450123 518331 450189 518332
rect 450862 517581 450922 520170
rect 451330 519890 451390 520200
rect 451484 520170 452026 520230
rect 451230 519830 451390 519890
rect 451230 518805 451290 519830
rect 451227 518804 451293 518805
rect 451227 518740 451228 518804
rect 451292 518740 451293 518804
rect 451227 518739 451293 518740
rect 451966 517581 452026 520170
rect 452498 519890 452558 520200
rect 452652 520170 453314 520230
rect 452498 519830 452578 519890
rect 452518 518805 452578 519830
rect 452515 518804 452581 518805
rect 452515 518740 452516 518804
rect 452580 518740 452581 518804
rect 452515 518739 452581 518740
rect 453254 517717 453314 520170
rect 453622 520170 453696 520230
rect 453622 518533 453682 520170
rect 453619 518532 453685 518533
rect 453619 518468 453620 518532
rect 453684 518468 453685 518532
rect 453619 518467 453685 518468
rect 453251 517716 453317 517717
rect 453251 517652 453252 517716
rect 453316 517652 453317 517716
rect 453251 517651 453317 517652
rect 453806 517581 453866 520230
rect 454834 519890 454894 520200
rect 454988 520170 455338 520230
rect 454726 519830 454894 519890
rect 454726 518533 454786 519830
rect 454723 518532 454789 518533
rect 454723 518468 454724 518532
rect 454788 518468 454789 518532
rect 454723 518467 454789 518468
rect 455278 517581 455338 520170
rect 456002 519890 456062 520200
rect 456156 520170 456442 520230
rect 456002 519830 456074 519890
rect 456014 518533 456074 519830
rect 456011 518532 456077 518533
rect 456011 518468 456012 518532
rect 456076 518468 456077 518532
rect 456011 518467 456077 518468
rect 456382 517581 456442 520170
rect 457118 520170 457200 520230
rect 457324 520170 457914 520230
rect 457118 518669 457178 520170
rect 457115 518668 457181 518669
rect 457115 518604 457116 518668
rect 457180 518604 457181 518668
rect 457115 518603 457181 518604
rect 457854 517581 457914 520170
rect 458338 519890 458398 520200
rect 458492 520170 459202 520230
rect 458338 519830 458466 519890
rect 458406 518805 458466 519830
rect 458403 518804 458469 518805
rect 458403 518740 458404 518804
rect 458468 518740 458469 518804
rect 458403 518739 458469 518740
rect 459142 517581 459202 520170
rect 459506 519890 459566 520200
rect 459660 520170 460306 520230
rect 459506 519830 459570 519890
rect 459510 518397 459570 519830
rect 459507 518396 459573 518397
rect 459507 518332 459508 518396
rect 459572 518332 459573 518396
rect 459507 518331 459573 518332
rect 460246 517717 460306 520170
rect 460430 520170 460704 520230
rect 460430 518805 460490 520170
rect 460427 518804 460493 518805
rect 460427 518740 460428 518804
rect 460492 518740 460493 518804
rect 460427 518739 460493 518740
rect 460243 517716 460309 517717
rect 460243 517652 460244 517716
rect 460308 517652 460309 517716
rect 460243 517651 460309 517652
rect 460798 517581 460858 520200
rect 461166 520170 461872 520230
rect 461996 520170 462146 520230
rect 461166 518669 461226 520170
rect 461163 518668 461229 518669
rect 461163 518604 461164 518668
rect 461228 518604 461229 518668
rect 461163 518603 461229 518604
rect 462086 517581 462146 520170
rect 462454 520170 463040 520230
rect 463164 520170 463618 520230
rect 462454 518533 462514 520170
rect 462451 518532 462517 518533
rect 462451 518468 462452 518532
rect 462516 518468 462517 518532
rect 462451 518467 462517 518468
rect 463558 517581 463618 520170
rect 463926 520170 464208 520230
rect 464332 520170 464906 520230
rect 463926 518533 463986 520170
rect 463923 518532 463989 518533
rect 463923 518468 463924 518532
rect 463988 518468 463989 518532
rect 463923 518467 463989 518468
rect 464846 517581 464906 520170
rect 465214 520170 465376 520230
rect 465500 520170 466194 520230
rect 465214 518397 465274 520170
rect 465211 518396 465277 518397
rect 465211 518332 465212 518396
rect 465276 518332 465277 518396
rect 465211 518331 465277 518332
rect 466134 517581 466194 520170
rect 466502 518805 466562 520230
rect 466668 520170 467298 520230
rect 466499 518804 466565 518805
rect 466499 518740 466500 518804
rect 466564 518740 466565 518804
rect 466499 518739 466565 518740
rect 467238 517581 467298 520170
rect 467422 520170 467712 520230
rect 467836 520170 468402 520230
rect 467422 518533 467482 520170
rect 467419 518532 467485 518533
rect 467419 518468 467420 518532
rect 467484 518468 467485 518532
rect 467419 518467 467485 518468
rect 468342 517717 468402 520170
rect 468526 520170 468880 520230
rect 468526 518261 468586 520170
rect 468974 519890 469034 520200
rect 468974 519830 469138 519890
rect 468523 518260 468589 518261
rect 468523 518196 468524 518260
rect 468588 518196 468589 518260
rect 468523 518195 468589 518196
rect 468339 517716 468405 517717
rect 468339 517652 468340 517716
rect 468404 517652 468405 517716
rect 468339 517651 468405 517652
rect 469078 517581 469138 519830
rect 438347 517580 438413 517581
rect 438347 517516 438348 517580
rect 438412 517516 438413 517580
rect 438347 517515 438413 517516
rect 438715 517580 438781 517581
rect 438715 517516 438716 517580
rect 438780 517516 438781 517580
rect 438715 517515 438781 517516
rect 439635 517580 439701 517581
rect 439635 517516 439636 517580
rect 439700 517516 439701 517580
rect 439635 517515 439701 517516
rect 440003 517580 440069 517581
rect 440003 517516 440004 517580
rect 440068 517516 440069 517580
rect 440003 517515 440069 517516
rect 441475 517580 441541 517581
rect 441475 517516 441476 517580
rect 441540 517516 441541 517580
rect 441475 517515 441541 517516
rect 442763 517580 442829 517581
rect 442763 517516 442764 517580
rect 442828 517516 442829 517580
rect 442763 517515 442829 517516
rect 449755 517580 449821 517581
rect 449755 517516 449756 517580
rect 449820 517516 449821 517580
rect 449755 517515 449821 517516
rect 450859 517580 450925 517581
rect 450859 517516 450860 517580
rect 450924 517516 450925 517580
rect 450859 517515 450925 517516
rect 451963 517580 452029 517581
rect 451963 517516 451964 517580
rect 452028 517516 452029 517580
rect 451963 517515 452029 517516
rect 453803 517580 453869 517581
rect 453803 517516 453804 517580
rect 453868 517516 453869 517580
rect 453803 517515 453869 517516
rect 455275 517580 455341 517581
rect 455275 517516 455276 517580
rect 455340 517516 455341 517580
rect 455275 517515 455341 517516
rect 456379 517580 456445 517581
rect 456379 517516 456380 517580
rect 456444 517516 456445 517580
rect 456379 517515 456445 517516
rect 457851 517580 457917 517581
rect 457851 517516 457852 517580
rect 457916 517516 457917 517580
rect 457851 517515 457917 517516
rect 459139 517580 459205 517581
rect 459139 517516 459140 517580
rect 459204 517516 459205 517580
rect 459139 517515 459205 517516
rect 460795 517580 460861 517581
rect 460795 517516 460796 517580
rect 460860 517516 460861 517580
rect 460795 517515 460861 517516
rect 462083 517580 462149 517581
rect 462083 517516 462084 517580
rect 462148 517516 462149 517580
rect 462083 517515 462149 517516
rect 463555 517580 463621 517581
rect 463555 517516 463556 517580
rect 463620 517516 463621 517580
rect 463555 517515 463621 517516
rect 464843 517580 464909 517581
rect 464843 517516 464844 517580
rect 464908 517516 464909 517580
rect 464843 517515 464909 517516
rect 466131 517580 466197 517581
rect 466131 517516 466132 517580
rect 466196 517516 466197 517580
rect 466131 517515 466197 517516
rect 467235 517580 467301 517581
rect 467235 517516 467236 517580
rect 467300 517516 467301 517580
rect 467235 517515 467301 517516
rect 469075 517580 469141 517581
rect 469075 517516 469076 517580
rect 469140 517516 469141 517580
rect 469075 517515 469141 517516
rect 414804 488218 414986 488454
rect 415222 488218 415404 488454
rect 414804 488134 415404 488218
rect 414804 487898 414986 488134
rect 415222 487898 415404 488134
rect 414804 483000 415404 487898
rect 418404 492054 419004 517000
rect 418404 491818 418586 492054
rect 418822 491818 419004 492054
rect 418404 491734 419004 491818
rect 418404 491498 418586 491734
rect 418822 491498 419004 491734
rect 418404 483000 419004 491498
rect 422004 495654 422604 517000
rect 422004 495418 422186 495654
rect 422422 495418 422604 495654
rect 422004 495334 422604 495418
rect 422004 495098 422186 495334
rect 422422 495098 422604 495334
rect 422004 483000 422604 495098
rect 425604 499254 426204 517000
rect 425604 499018 425786 499254
rect 426022 499018 426204 499254
rect 425604 498934 426204 499018
rect 425604 498698 425786 498934
rect 426022 498698 426204 498934
rect 425604 483000 426204 498698
rect 432804 506454 433404 517000
rect 432804 506218 432986 506454
rect 433222 506218 433404 506454
rect 432804 506134 433404 506218
rect 432804 505898 432986 506134
rect 433222 505898 433404 506134
rect 432804 483000 433404 505898
rect 436404 510054 437004 517000
rect 436404 509818 436586 510054
rect 436822 509818 437004 510054
rect 436404 509734 437004 509818
rect 436404 509498 436586 509734
rect 436822 509498 437004 509734
rect 433931 495548 433997 495549
rect 433931 495484 433932 495548
rect 433996 495484 433997 495548
rect 433931 495483 433997 495484
rect 433934 492693 433994 495483
rect 433931 492692 433997 492693
rect 433931 492628 433932 492692
rect 433996 492628 433997 492692
rect 433931 492627 433997 492628
rect 436404 483000 437004 509498
rect 440004 513654 440604 517000
rect 440004 513418 440186 513654
rect 440422 513418 440604 513654
rect 440004 513334 440604 513418
rect 440004 513098 440186 513334
rect 440422 513098 440604 513334
rect 440004 483000 440604 513098
rect 443604 483000 444204 517000
rect 450804 488454 451404 517000
rect 450804 488218 450986 488454
rect 451222 488218 451404 488454
rect 450804 488134 451404 488218
rect 450804 487898 450986 488134
rect 451222 487898 451404 488134
rect 450804 483000 451404 487898
rect 454404 492054 455004 517000
rect 454404 491818 454586 492054
rect 454822 491818 455004 492054
rect 454404 491734 455004 491818
rect 454404 491498 454586 491734
rect 454822 491498 455004 491734
rect 454404 483000 455004 491498
rect 458004 495654 458604 517000
rect 458004 495418 458186 495654
rect 458422 495418 458604 495654
rect 458004 495334 458604 495418
rect 458004 495098 458186 495334
rect 458422 495098 458604 495334
rect 458004 483000 458604 495098
rect 461604 499254 462204 517000
rect 461604 499018 461786 499254
rect 462022 499018 462204 499254
rect 461604 498934 462204 499018
rect 461604 498698 461786 498934
rect 462022 498698 462204 498934
rect 461604 483000 462204 498698
rect 468804 506454 469404 517000
rect 468804 506218 468986 506454
rect 469222 506218 469404 506454
rect 468804 506134 469404 506218
rect 468804 505898 468986 506134
rect 469222 505898 469404 506134
rect 468804 483000 469404 505898
rect 472404 510054 473004 517000
rect 472404 509818 472586 510054
rect 472822 509818 473004 510054
rect 472404 509734 473004 509818
rect 472404 509498 472586 509734
rect 472822 509498 473004 509734
rect 472404 483000 473004 509498
rect 476004 513654 476604 517000
rect 476004 513418 476186 513654
rect 476422 513418 476604 513654
rect 476004 513334 476604 513418
rect 476004 513098 476186 513334
rect 476422 513098 476604 513334
rect 476004 483000 476604 513098
rect 479604 483000 480204 517000
rect 486804 488454 487404 517000
rect 486804 488218 486986 488454
rect 487222 488218 487404 488454
rect 486804 488134 487404 488218
rect 486804 487898 486986 488134
rect 487222 487898 487404 488134
rect 486804 483000 487404 487898
rect 490404 492054 491004 517000
rect 490404 491818 490586 492054
rect 490822 491818 491004 492054
rect 490404 491734 491004 491818
rect 490404 491498 490586 491734
rect 490822 491498 491004 491734
rect 490404 483000 491004 491498
rect 494004 495654 494604 517000
rect 494004 495418 494186 495654
rect 494422 495418 494604 495654
rect 494004 495334 494604 495418
rect 494004 495098 494186 495334
rect 494422 495098 494604 495334
rect 494004 483000 494604 495098
rect 497604 499254 498204 517000
rect 497604 499018 497786 499254
rect 498022 499018 498204 499254
rect 497604 498934 498204 499018
rect 497604 498698 497786 498934
rect 498022 498698 498204 498934
rect 497604 483000 498204 498698
rect 504804 506454 505404 541898
rect 504804 506218 504986 506454
rect 505222 506218 505404 506454
rect 504804 506134 505404 506218
rect 504804 505898 504986 506134
rect 505222 505898 505404 506134
rect 504804 483000 505404 505898
rect 508404 690054 509004 706162
rect 508404 689818 508586 690054
rect 508822 689818 509004 690054
rect 508404 689734 509004 689818
rect 508404 689498 508586 689734
rect 508822 689498 509004 689734
rect 508404 654054 509004 689498
rect 508404 653818 508586 654054
rect 508822 653818 509004 654054
rect 508404 653734 509004 653818
rect 508404 653498 508586 653734
rect 508822 653498 509004 653734
rect 508404 618054 509004 653498
rect 508404 617818 508586 618054
rect 508822 617818 509004 618054
rect 508404 617734 509004 617818
rect 508404 617498 508586 617734
rect 508822 617498 509004 617734
rect 508404 582054 509004 617498
rect 508404 581818 508586 582054
rect 508822 581818 509004 582054
rect 508404 581734 509004 581818
rect 508404 581498 508586 581734
rect 508822 581498 509004 581734
rect 508404 546054 509004 581498
rect 508404 545818 508586 546054
rect 508822 545818 509004 546054
rect 508404 545734 509004 545818
rect 508404 545498 508586 545734
rect 508822 545498 509004 545734
rect 508404 510054 509004 545498
rect 508404 509818 508586 510054
rect 508822 509818 509004 510054
rect 508404 509734 509004 509818
rect 508404 509498 508586 509734
rect 508822 509498 509004 509734
rect 508404 483000 509004 509498
rect 512004 693654 512604 708042
rect 512004 693418 512186 693654
rect 512422 693418 512604 693654
rect 512004 693334 512604 693418
rect 512004 693098 512186 693334
rect 512422 693098 512604 693334
rect 512004 657654 512604 693098
rect 512004 657418 512186 657654
rect 512422 657418 512604 657654
rect 512004 657334 512604 657418
rect 512004 657098 512186 657334
rect 512422 657098 512604 657334
rect 512004 621654 512604 657098
rect 512004 621418 512186 621654
rect 512422 621418 512604 621654
rect 512004 621334 512604 621418
rect 512004 621098 512186 621334
rect 512422 621098 512604 621334
rect 512004 585654 512604 621098
rect 512004 585418 512186 585654
rect 512422 585418 512604 585654
rect 512004 585334 512604 585418
rect 512004 585098 512186 585334
rect 512422 585098 512604 585334
rect 512004 549654 512604 585098
rect 512004 549418 512186 549654
rect 512422 549418 512604 549654
rect 512004 549334 512604 549418
rect 512004 549098 512186 549334
rect 512422 549098 512604 549334
rect 512004 513654 512604 549098
rect 512004 513418 512186 513654
rect 512422 513418 512604 513654
rect 512004 513334 512604 513418
rect 512004 513098 512186 513334
rect 512422 513098 512604 513334
rect 512004 483000 512604 513098
rect 515604 697254 516204 709922
rect 533604 711418 534204 711440
rect 533604 711182 533786 711418
rect 534022 711182 534204 711418
rect 533604 711098 534204 711182
rect 533604 710862 533786 711098
rect 534022 710862 534204 711098
rect 530004 709538 530604 709560
rect 530004 709302 530186 709538
rect 530422 709302 530604 709538
rect 530004 709218 530604 709302
rect 530004 708982 530186 709218
rect 530422 708982 530604 709218
rect 526404 707658 527004 707680
rect 526404 707422 526586 707658
rect 526822 707422 527004 707658
rect 526404 707338 527004 707422
rect 526404 707102 526586 707338
rect 526822 707102 527004 707338
rect 515604 697018 515786 697254
rect 516022 697018 516204 697254
rect 515604 696934 516204 697018
rect 515604 696698 515786 696934
rect 516022 696698 516204 696934
rect 515604 661254 516204 696698
rect 515604 661018 515786 661254
rect 516022 661018 516204 661254
rect 515604 660934 516204 661018
rect 515604 660698 515786 660934
rect 516022 660698 516204 660934
rect 515604 625254 516204 660698
rect 515604 625018 515786 625254
rect 516022 625018 516204 625254
rect 515604 624934 516204 625018
rect 515604 624698 515786 624934
rect 516022 624698 516204 624934
rect 515604 589254 516204 624698
rect 515604 589018 515786 589254
rect 516022 589018 516204 589254
rect 515604 588934 516204 589018
rect 515604 588698 515786 588934
rect 516022 588698 516204 588934
rect 515604 553254 516204 588698
rect 515604 553018 515786 553254
rect 516022 553018 516204 553254
rect 515604 552934 516204 553018
rect 515604 552698 515786 552934
rect 516022 552698 516204 552934
rect 515604 517254 516204 552698
rect 515604 517018 515786 517254
rect 516022 517018 516204 517254
rect 515604 516934 516204 517018
rect 515604 516698 515786 516934
rect 516022 516698 516204 516934
rect 515604 483000 516204 516698
rect 522804 705778 523404 705800
rect 522804 705542 522986 705778
rect 523222 705542 523404 705778
rect 522804 705458 523404 705542
rect 522804 705222 522986 705458
rect 523222 705222 523404 705458
rect 522804 668454 523404 705222
rect 522804 668218 522986 668454
rect 523222 668218 523404 668454
rect 522804 668134 523404 668218
rect 522804 667898 522986 668134
rect 523222 667898 523404 668134
rect 522804 632454 523404 667898
rect 522804 632218 522986 632454
rect 523222 632218 523404 632454
rect 522804 632134 523404 632218
rect 522804 631898 522986 632134
rect 523222 631898 523404 632134
rect 522804 596454 523404 631898
rect 522804 596218 522986 596454
rect 523222 596218 523404 596454
rect 522804 596134 523404 596218
rect 522804 595898 522986 596134
rect 523222 595898 523404 596134
rect 522804 560454 523404 595898
rect 522804 560218 522986 560454
rect 523222 560218 523404 560454
rect 522804 560134 523404 560218
rect 522804 559898 522986 560134
rect 523222 559898 523404 560134
rect 522804 524454 523404 559898
rect 522804 524218 522986 524454
rect 523222 524218 523404 524454
rect 522804 524134 523404 524218
rect 522804 523898 522986 524134
rect 523222 523898 523404 524134
rect 522804 488454 523404 523898
rect 522804 488218 522986 488454
rect 523222 488218 523404 488454
rect 522804 488134 523404 488218
rect 522804 487898 522986 488134
rect 523222 487898 523404 488134
rect 522804 483000 523404 487898
rect 526404 672054 527004 707102
rect 526404 671818 526586 672054
rect 526822 671818 527004 672054
rect 526404 671734 527004 671818
rect 526404 671498 526586 671734
rect 526822 671498 527004 671734
rect 526404 636054 527004 671498
rect 526404 635818 526586 636054
rect 526822 635818 527004 636054
rect 526404 635734 527004 635818
rect 526404 635498 526586 635734
rect 526822 635498 527004 635734
rect 526404 600054 527004 635498
rect 526404 599818 526586 600054
rect 526822 599818 527004 600054
rect 526404 599734 527004 599818
rect 526404 599498 526586 599734
rect 526822 599498 527004 599734
rect 526404 564054 527004 599498
rect 526404 563818 526586 564054
rect 526822 563818 527004 564054
rect 526404 563734 527004 563818
rect 526404 563498 526586 563734
rect 526822 563498 527004 563734
rect 526404 528054 527004 563498
rect 526404 527818 526586 528054
rect 526822 527818 527004 528054
rect 526404 527734 527004 527818
rect 526404 527498 526586 527734
rect 526822 527498 527004 527734
rect 526404 492054 527004 527498
rect 526404 491818 526586 492054
rect 526822 491818 527004 492054
rect 526404 491734 527004 491818
rect 526404 491498 526586 491734
rect 526822 491498 527004 491734
rect 526404 483000 527004 491498
rect 530004 675654 530604 708982
rect 530004 675418 530186 675654
rect 530422 675418 530604 675654
rect 530004 675334 530604 675418
rect 530004 675098 530186 675334
rect 530422 675098 530604 675334
rect 530004 639654 530604 675098
rect 530004 639418 530186 639654
rect 530422 639418 530604 639654
rect 530004 639334 530604 639418
rect 530004 639098 530186 639334
rect 530422 639098 530604 639334
rect 530004 603654 530604 639098
rect 530004 603418 530186 603654
rect 530422 603418 530604 603654
rect 530004 603334 530604 603418
rect 530004 603098 530186 603334
rect 530422 603098 530604 603334
rect 530004 567654 530604 603098
rect 530004 567418 530186 567654
rect 530422 567418 530604 567654
rect 530004 567334 530604 567418
rect 530004 567098 530186 567334
rect 530422 567098 530604 567334
rect 530004 531654 530604 567098
rect 530004 531418 530186 531654
rect 530422 531418 530604 531654
rect 530004 531334 530604 531418
rect 530004 531098 530186 531334
rect 530422 531098 530604 531334
rect 530004 495654 530604 531098
rect 530004 495418 530186 495654
rect 530422 495418 530604 495654
rect 530004 495334 530604 495418
rect 530004 495098 530186 495334
rect 530422 495098 530604 495334
rect 530004 483000 530604 495098
rect 533604 679254 534204 710862
rect 551604 710478 552204 711440
rect 551604 710242 551786 710478
rect 552022 710242 552204 710478
rect 551604 710158 552204 710242
rect 551604 709922 551786 710158
rect 552022 709922 552204 710158
rect 548004 708598 548604 709560
rect 548004 708362 548186 708598
rect 548422 708362 548604 708598
rect 548004 708278 548604 708362
rect 548004 708042 548186 708278
rect 548422 708042 548604 708278
rect 544404 706718 545004 707680
rect 544404 706482 544586 706718
rect 544822 706482 545004 706718
rect 544404 706398 545004 706482
rect 544404 706162 544586 706398
rect 544822 706162 545004 706398
rect 540804 704838 541404 705800
rect 540804 704602 540986 704838
rect 541222 704602 541404 704838
rect 540804 704518 541404 704602
rect 540804 704282 540986 704518
rect 541222 704282 541404 704518
rect 538259 700772 538325 700773
rect 538259 700708 538260 700772
rect 538324 700708 538325 700772
rect 538259 700707 538325 700708
rect 533604 679018 533786 679254
rect 534022 679018 534204 679254
rect 533604 678934 534204 679018
rect 533604 678698 533786 678934
rect 534022 678698 534204 678934
rect 533604 643254 534204 678698
rect 533604 643018 533786 643254
rect 534022 643018 534204 643254
rect 533604 642934 534204 643018
rect 533604 642698 533786 642934
rect 534022 642698 534204 642934
rect 533604 607254 534204 642698
rect 533604 607018 533786 607254
rect 534022 607018 534204 607254
rect 533604 606934 534204 607018
rect 533604 606698 533786 606934
rect 534022 606698 534204 606934
rect 533604 571254 534204 606698
rect 533604 571018 533786 571254
rect 534022 571018 534204 571254
rect 533604 570934 534204 571018
rect 533604 570698 533786 570934
rect 534022 570698 534204 570934
rect 533604 535254 534204 570698
rect 533604 535018 533786 535254
rect 534022 535018 534204 535254
rect 533604 534934 534204 535018
rect 533604 534698 533786 534934
rect 534022 534698 534204 534934
rect 533604 499254 534204 534698
rect 533604 499018 533786 499254
rect 534022 499018 534204 499254
rect 533604 498934 534204 499018
rect 533604 498698 533786 498934
rect 534022 498698 534204 498934
rect 533604 483000 534204 498698
rect 252804 470218 252986 470454
rect 253222 470218 253404 470454
rect 252804 470134 253404 470218
rect 252804 469898 252986 470134
rect 253222 469898 253404 470134
rect 252804 434454 253404 469898
rect 264208 470454 264528 470476
rect 264208 470218 264250 470454
rect 264486 470218 264528 470454
rect 264208 470134 264528 470218
rect 264208 469898 264250 470134
rect 264486 469898 264528 470134
rect 264208 469876 264528 469898
rect 279568 452454 279888 452476
rect 279568 452218 279610 452454
rect 279846 452218 279888 452454
rect 279568 452134 279888 452218
rect 279568 451898 279610 452134
rect 279846 451898 279888 452134
rect 279568 451876 279888 451898
rect 252804 434218 252986 434454
rect 253222 434218 253404 434454
rect 252804 434134 253404 434218
rect 252804 433898 252986 434134
rect 253222 433898 253404 434134
rect 252804 398454 253404 433898
rect 264208 434454 264528 434476
rect 264208 434218 264250 434454
rect 264486 434218 264528 434454
rect 264208 434134 264528 434218
rect 264208 433898 264250 434134
rect 264486 433898 264528 434134
rect 264208 433876 264528 433898
rect 538262 427410 538322 700707
rect 538443 700636 538509 700637
rect 538443 700572 538444 700636
rect 538508 700572 538509 700636
rect 538443 700571 538509 700572
rect 538078 427350 538322 427410
rect 538078 426050 538138 427350
rect 538078 425990 538322 426050
rect 279568 416454 279888 416476
rect 279568 416218 279610 416454
rect 279846 416218 279888 416454
rect 279568 416134 279888 416218
rect 279568 415898 279610 416134
rect 279846 415898 279888 416134
rect 279568 415876 279888 415898
rect 538262 399530 538322 425990
rect 538078 399470 538322 399530
rect 538446 399530 538506 700571
rect 540099 700500 540165 700501
rect 540099 700436 540100 700500
rect 540164 700436 540165 700500
rect 540099 700435 540165 700436
rect 539915 700364 539981 700365
rect 539915 700300 539916 700364
rect 539980 700300 539981 700364
rect 539915 700299 539981 700300
rect 538811 623796 538877 623797
rect 538811 623732 538812 623796
rect 538876 623732 538877 623796
rect 538811 623731 538877 623732
rect 538814 437610 538874 623731
rect 539547 469980 539613 469981
rect 539547 469916 539548 469980
rect 539612 469916 539613 469980
rect 539547 469915 539613 469916
rect 539363 455292 539429 455293
rect 539363 455290 539364 455292
rect 539182 455230 539364 455290
rect 539182 451210 539242 455230
rect 539363 455228 539364 455230
rect 539428 455228 539429 455292
rect 539363 455227 539429 455228
rect 539363 451212 539429 451213
rect 539363 451210 539364 451212
rect 539182 451150 539364 451210
rect 539363 451148 539364 451150
rect 539428 451148 539429 451212
rect 539363 451147 539429 451148
rect 539363 442644 539429 442645
rect 539363 442580 539364 442644
rect 539428 442580 539429 442644
rect 539363 442579 539429 442580
rect 539366 442370 539426 442579
rect 538630 437550 538874 437610
rect 538998 442310 539426 442370
rect 538630 436250 538690 437550
rect 538630 436190 538874 436250
rect 538814 416530 538874 436190
rect 538998 428770 539058 442310
rect 539363 442236 539429 442237
rect 539363 442172 539364 442236
rect 539428 442172 539429 442236
rect 539363 442171 539429 442172
rect 538998 428710 539242 428770
rect 539182 417346 539242 428710
rect 539366 417890 539426 442171
rect 539550 418437 539610 469915
rect 539731 463724 539797 463725
rect 539731 463660 539732 463724
rect 539796 463660 539797 463724
rect 539731 463659 539797 463660
rect 539734 452029 539794 463659
rect 539731 452028 539797 452029
rect 539731 451964 539732 452028
rect 539796 451964 539797 452028
rect 539731 451963 539797 451964
rect 539731 451212 539797 451213
rect 539731 451148 539732 451212
rect 539796 451148 539797 451212
rect 539731 451147 539797 451148
rect 539734 442509 539794 451147
rect 539731 442508 539797 442509
rect 539731 442444 539732 442508
rect 539796 442444 539797 442508
rect 539731 442443 539797 442444
rect 539731 442372 539797 442373
rect 539731 442308 539732 442372
rect 539796 442308 539797 442372
rect 539731 442307 539797 442308
rect 539734 432717 539794 442307
rect 539731 432716 539797 432717
rect 539731 432652 539732 432716
rect 539796 432652 539797 432716
rect 539731 432651 539797 432652
rect 539547 418436 539613 418437
rect 539547 418372 539548 418436
rect 539612 418372 539613 418436
rect 539547 418371 539613 418372
rect 539366 417830 539794 417890
rect 539182 417286 539610 417346
rect 538814 416470 539242 416530
rect 539182 415034 539242 416470
rect 539363 415036 539429 415037
rect 539363 415034 539364 415036
rect 539182 414974 539364 415034
rect 539363 414972 539364 414974
rect 539428 414972 539429 415036
rect 539363 414971 539429 414972
rect 539363 414492 539429 414493
rect 539363 414490 539364 414492
rect 538630 414430 539364 414490
rect 538630 401570 538690 414430
rect 539363 414428 539364 414430
rect 539428 414428 539429 414492
rect 539363 414427 539429 414428
rect 539363 413812 539429 413813
rect 539363 413810 539364 413812
rect 539182 413750 539364 413810
rect 539182 413130 539242 413750
rect 539363 413748 539364 413750
rect 539428 413748 539429 413812
rect 539363 413747 539429 413748
rect 538814 413070 539242 413130
rect 538814 403746 538874 413070
rect 539550 406469 539610 417286
rect 539734 414493 539794 417830
rect 539731 414492 539797 414493
rect 539731 414428 539732 414492
rect 539796 414428 539797 414492
rect 539731 414427 539797 414428
rect 539731 413404 539797 413405
rect 539731 413340 539732 413404
rect 539796 413340 539797 413404
rect 539731 413339 539797 413340
rect 539547 406468 539613 406469
rect 539547 406404 539548 406468
rect 539612 406404 539613 406468
rect 539547 406403 539613 406404
rect 539363 405788 539429 405789
rect 539363 405724 539364 405788
rect 539428 405724 539429 405788
rect 539363 405723 539429 405724
rect 538814 403686 539058 403746
rect 538630 401510 538874 401570
rect 538446 399470 538690 399530
rect 538078 398850 538138 399470
rect 538630 398850 538690 399470
rect 538078 398790 538322 398850
rect 252804 398218 252986 398454
rect 253222 398218 253404 398454
rect 252804 398134 253404 398218
rect 252804 397898 252986 398134
rect 253222 397898 253404 398134
rect 252804 362454 253404 397898
rect 264208 398454 264528 398476
rect 264208 398218 264250 398454
rect 264486 398218 264528 398454
rect 264208 398134 264528 398218
rect 264208 397898 264250 398134
rect 264486 397898 264528 398134
rect 264208 397876 264528 397898
rect 279568 380454 279888 380476
rect 279568 380218 279610 380454
rect 279846 380218 279888 380454
rect 279568 380134 279888 380218
rect 279568 379898 279610 380134
rect 279846 379898 279888 380134
rect 279568 379876 279888 379898
rect 538262 377770 538322 398790
rect 538446 398790 538690 398850
rect 538814 398850 538874 401510
rect 538998 399530 539058 403686
rect 539366 402253 539426 405723
rect 539734 403749 539794 413339
rect 539731 403748 539797 403749
rect 539731 403684 539732 403748
rect 539796 403684 539797 403748
rect 539731 403683 539797 403684
rect 539363 402252 539429 402253
rect 539363 402188 539364 402252
rect 539428 402188 539429 402252
rect 539363 402187 539429 402188
rect 539363 399532 539429 399533
rect 539363 399530 539364 399532
rect 538998 399470 539364 399530
rect 539363 399468 539364 399470
rect 539428 399468 539429 399532
rect 539363 399467 539429 399468
rect 539547 399124 539613 399125
rect 539547 399060 539548 399124
rect 539612 399060 539613 399124
rect 539547 399059 539613 399060
rect 539550 398850 539610 399059
rect 538814 398790 539610 398850
rect 538446 384570 538506 398790
rect 539547 398580 539613 398581
rect 539547 398516 539548 398580
rect 539612 398516 539613 398580
rect 539547 398515 539613 398516
rect 539363 395452 539429 395453
rect 539363 395450 539364 395452
rect 538814 395390 539364 395450
rect 538814 388514 538874 395390
rect 539363 395388 539364 395390
rect 539428 395388 539429 395452
rect 539363 395387 539429 395388
rect 539363 391372 539429 391373
rect 539363 391370 539364 391372
rect 539182 391310 539364 391370
rect 539182 388650 539242 391310
rect 539363 391308 539364 391310
rect 539428 391308 539429 391372
rect 539363 391307 539429 391308
rect 539363 388652 539429 388653
rect 539363 388650 539364 388652
rect 539182 388590 539364 388650
rect 539363 388588 539364 388590
rect 539428 388588 539429 388652
rect 539363 388587 539429 388588
rect 539363 388516 539429 388517
rect 539363 388514 539364 388516
rect 538814 388454 539364 388514
rect 539363 388452 539364 388454
rect 539428 388452 539429 388516
rect 539363 388451 539429 388452
rect 539363 384572 539429 384573
rect 539363 384570 539364 384572
rect 538446 384510 539364 384570
rect 539363 384508 539364 384510
rect 539428 384508 539429 384572
rect 539363 384507 539429 384508
rect 539363 383484 539429 383485
rect 539363 383420 539364 383484
rect 539428 383420 539429 383484
rect 539363 383419 539429 383420
rect 538262 377710 538506 377770
rect 538446 376274 538506 377710
rect 539366 376413 539426 383419
rect 539363 376412 539429 376413
rect 539363 376348 539364 376412
rect 539428 376348 539429 376412
rect 539363 376347 539429 376348
rect 539363 376276 539429 376277
rect 539363 376274 539364 376276
rect 538446 376214 539364 376274
rect 539363 376212 539364 376214
rect 539428 376212 539429 376276
rect 539363 376211 539429 376212
rect 539363 374644 539429 374645
rect 539363 374580 539364 374644
rect 539428 374580 539429 374644
rect 539363 374579 539429 374580
rect 539366 372330 539426 374579
rect 538814 372270 539426 372330
rect 538814 369746 538874 372270
rect 538630 369686 538874 369746
rect 252804 362218 252986 362454
rect 253222 362218 253404 362454
rect 252804 362134 253404 362218
rect 252804 361898 252986 362134
rect 253222 361898 253404 362134
rect 252804 326454 253404 361898
rect 264208 362454 264528 362476
rect 264208 362218 264250 362454
rect 264486 362218 264528 362454
rect 264208 362134 264528 362218
rect 264208 361898 264250 362134
rect 264486 361898 264528 362134
rect 264208 361876 264528 361898
rect 538630 352610 538690 369686
rect 539363 364172 539429 364173
rect 539363 364170 539364 364172
rect 539182 364110 539364 364170
rect 538630 352550 538874 352610
rect 279568 344454 279888 344476
rect 279568 344218 279610 344454
rect 279846 344218 279888 344454
rect 279568 344134 279888 344218
rect 279568 343898 279610 344134
rect 279846 343898 279888 344134
rect 279568 343876 279888 343898
rect 538814 342410 538874 352550
rect 538446 342350 538874 342410
rect 538446 341730 538506 342350
rect 538262 341670 538506 341730
rect 538262 327450 538322 341670
rect 539182 330170 539242 364110
rect 539363 364108 539364 364110
rect 539428 364108 539429 364172
rect 539363 364107 539429 364108
rect 539550 359549 539610 398515
rect 539918 388517 539978 700299
rect 540102 390557 540162 700435
rect 540804 686454 541404 704282
rect 540804 686218 540986 686454
rect 541222 686218 541404 686454
rect 540804 686134 541404 686218
rect 540804 685898 540986 686134
rect 541222 685898 541404 686134
rect 540804 650454 541404 685898
rect 540804 650218 540986 650454
rect 541222 650218 541404 650454
rect 540804 650134 541404 650218
rect 540804 649898 540986 650134
rect 541222 649898 541404 650134
rect 540804 614454 541404 649898
rect 540804 614218 540986 614454
rect 541222 614218 541404 614454
rect 540804 614134 541404 614218
rect 540804 613898 540986 614134
rect 541222 613898 541404 614134
rect 540804 578454 541404 613898
rect 540804 578218 540986 578454
rect 541222 578218 541404 578454
rect 540804 578134 541404 578218
rect 540804 577898 540986 578134
rect 541222 577898 541404 578134
rect 540804 542454 541404 577898
rect 540804 542218 540986 542454
rect 541222 542218 541404 542454
rect 540804 542134 541404 542218
rect 540804 541898 540986 542134
rect 541222 541898 541404 542134
rect 540804 506454 541404 541898
rect 540804 506218 540986 506454
rect 541222 506218 541404 506454
rect 540804 506134 541404 506218
rect 540804 505898 540986 506134
rect 541222 505898 541404 506134
rect 540804 483000 541404 505898
rect 544404 690054 545004 706162
rect 544404 689818 544586 690054
rect 544822 689818 545004 690054
rect 544404 689734 545004 689818
rect 544404 689498 544586 689734
rect 544822 689498 545004 689734
rect 544404 654054 545004 689498
rect 544404 653818 544586 654054
rect 544822 653818 545004 654054
rect 544404 653734 545004 653818
rect 544404 653498 544586 653734
rect 544822 653498 545004 653734
rect 544404 618054 545004 653498
rect 544404 617818 544586 618054
rect 544822 617818 545004 618054
rect 544404 617734 545004 617818
rect 544404 617498 544586 617734
rect 544822 617498 545004 617734
rect 544404 582054 545004 617498
rect 544404 581818 544586 582054
rect 544822 581818 545004 582054
rect 544404 581734 545004 581818
rect 544404 581498 544586 581734
rect 544822 581498 545004 581734
rect 544404 546054 545004 581498
rect 544404 545818 544586 546054
rect 544822 545818 545004 546054
rect 544404 545734 545004 545818
rect 544404 545498 544586 545734
rect 544822 545498 545004 545734
rect 544404 510054 545004 545498
rect 544404 509818 544586 510054
rect 544822 509818 545004 510054
rect 544404 509734 545004 509818
rect 544404 509498 544586 509734
rect 544822 509498 545004 509734
rect 542491 478956 542557 478957
rect 542491 478892 542492 478956
rect 542556 478892 542557 478956
rect 542491 478891 542557 478892
rect 542307 476916 542373 476917
rect 542307 476852 542308 476916
rect 542372 476852 542373 476916
rect 542307 476851 542373 476852
rect 541571 472700 541637 472701
rect 541571 472636 541572 472700
rect 541636 472636 541637 472700
rect 541571 472635 541637 472636
rect 540283 462092 540349 462093
rect 540283 462028 540284 462092
rect 540348 462028 540349 462092
rect 540283 462027 540349 462028
rect 540099 390556 540165 390557
rect 540099 390492 540100 390556
rect 540164 390492 540165 390556
rect 540099 390491 540165 390492
rect 539731 388516 539797 388517
rect 539731 388452 539732 388516
rect 539796 388452 539797 388516
rect 539731 388451 539797 388452
rect 539915 388516 539981 388517
rect 539915 388452 539916 388516
rect 539980 388452 539981 388516
rect 539915 388451 539981 388452
rect 539734 383485 539794 388451
rect 539731 383484 539797 383485
rect 539731 383420 539732 383484
rect 539796 383420 539797 383484
rect 539731 383419 539797 383420
rect 539731 381036 539797 381037
rect 539731 380972 539732 381036
rect 539796 380972 539797 381036
rect 539731 380971 539797 380972
rect 539734 379130 539794 380971
rect 539734 379070 539978 379130
rect 539731 376412 539797 376413
rect 539731 376348 539732 376412
rect 539796 376348 539797 376412
rect 539731 376347 539797 376348
rect 539734 374645 539794 376347
rect 539731 374644 539797 374645
rect 539731 374580 539732 374644
rect 539796 374580 539797 374644
rect 539731 374579 539797 374580
rect 539731 373284 539797 373285
rect 539731 373220 539732 373284
rect 539796 373220 539797 373284
rect 539731 373219 539797 373220
rect 539734 364173 539794 373219
rect 539731 364172 539797 364173
rect 539731 364108 539732 364172
rect 539796 364108 539797 364172
rect 539731 364107 539797 364108
rect 539918 363490 539978 379070
rect 539734 363430 539978 363490
rect 539547 359548 539613 359549
rect 539547 359484 539548 359548
rect 539612 359484 539613 359548
rect 539547 359483 539613 359484
rect 539547 359412 539613 359413
rect 539547 359348 539548 359412
rect 539612 359348 539613 359412
rect 539547 359347 539613 359348
rect 538998 330110 539242 330170
rect 538262 327390 538690 327450
rect 252804 326218 252986 326454
rect 253222 326218 253404 326454
rect 252804 326134 253404 326218
rect 252804 325898 252986 326134
rect 253222 325898 253404 326134
rect 252804 290454 253404 325898
rect 264208 326454 264528 326476
rect 264208 326218 264250 326454
rect 264486 326218 264528 326454
rect 264208 326134 264528 326218
rect 264208 325898 264250 326134
rect 264486 325898 264528 326134
rect 264208 325876 264528 325898
rect 538630 322690 538690 327390
rect 538262 322630 538690 322690
rect 538262 321330 538322 322630
rect 538998 322010 539058 330110
rect 538998 321950 539242 322010
rect 539182 321330 539242 321950
rect 538262 321270 538506 321330
rect 538446 317386 538506 321270
rect 538078 317326 538506 317386
rect 538814 321270 539242 321330
rect 279568 308454 279888 308476
rect 279568 308218 279610 308454
rect 279846 308218 279888 308454
rect 279568 308134 279888 308218
rect 279568 307898 279610 308134
rect 279846 307898 279888 308134
rect 279568 307876 279888 307898
rect 538078 300250 538138 317326
rect 538814 313170 538874 321270
rect 538814 313110 539058 313170
rect 538998 300930 539058 313110
rect 537894 300190 538138 300250
rect 538814 300870 539058 300930
rect 537894 291410 537954 300190
rect 538814 298210 538874 300870
rect 538814 298150 539242 298210
rect 539182 292770 539242 298150
rect 539363 292772 539429 292773
rect 539363 292770 539364 292772
rect 539182 292710 539364 292770
rect 539363 292708 539364 292710
rect 539428 292708 539429 292772
rect 539363 292707 539429 292708
rect 539363 292092 539429 292093
rect 539363 292090 539364 292092
rect 538998 292030 539364 292090
rect 537894 291350 538322 291410
rect 252804 290218 252986 290454
rect 253222 290218 253404 290454
rect 252804 290134 253404 290218
rect 252804 289898 252986 290134
rect 253222 289898 253404 290134
rect 252804 254454 253404 289898
rect 264208 290454 264528 290476
rect 264208 290218 264250 290454
rect 264486 290218 264528 290454
rect 264208 290134 264528 290218
rect 264208 289898 264250 290134
rect 264486 289898 264528 290134
rect 264208 289876 264528 289898
rect 538262 281890 538322 291350
rect 538998 286650 539058 292030
rect 539363 292028 539364 292030
rect 539428 292028 539429 292092
rect 539363 292027 539429 292028
rect 539363 286652 539429 286653
rect 539363 286650 539364 286652
rect 538998 286590 539364 286650
rect 539363 286588 539364 286590
rect 539428 286588 539429 286652
rect 539363 286587 539429 286588
rect 538262 281830 538874 281890
rect 279568 272454 279888 272476
rect 279568 272218 279610 272454
rect 279846 272218 279888 272454
rect 279568 272134 279888 272218
rect 279568 271898 279610 272134
rect 279846 271898 279888 272134
rect 279568 271876 279888 271898
rect 538814 265570 538874 281830
rect 538814 265510 539058 265570
rect 538998 256730 539058 265510
rect 539363 265028 539429 265029
rect 539363 264964 539364 265028
rect 539428 264964 539429 265028
rect 539363 264963 539429 264964
rect 539366 256869 539426 264963
rect 539363 256868 539429 256869
rect 539363 256804 539364 256868
rect 539428 256804 539429 256868
rect 539363 256803 539429 256804
rect 539363 256732 539429 256733
rect 539363 256730 539364 256732
rect 538814 256670 539058 256730
rect 539182 256670 539364 256730
rect 538814 254690 538874 256670
rect 538814 254630 539058 254690
rect 252804 254218 252986 254454
rect 253222 254218 253404 254454
rect 252804 254134 253404 254218
rect 252804 253898 252986 254134
rect 253222 253898 253404 254134
rect 252804 218454 253404 253898
rect 264208 254454 264528 254476
rect 264208 254218 264250 254454
rect 264486 254218 264528 254454
rect 264208 254134 264528 254218
rect 264208 253898 264250 254134
rect 264486 253898 264528 254134
rect 264208 253876 264528 253898
rect 538998 251290 539058 254630
rect 538446 251230 539058 251290
rect 538446 246530 538506 251230
rect 539182 250610 539242 256670
rect 539363 256668 539364 256670
rect 539428 256668 539429 256732
rect 539363 256667 539429 256668
rect 538998 250550 539242 250610
rect 538446 246470 538874 246530
rect 538814 242450 538874 246470
rect 538446 242390 538874 242450
rect 252804 218218 252986 218454
rect 253222 218218 253404 218454
rect 252804 218134 253404 218218
rect 252804 217898 252986 218134
rect 253222 217898 253404 218134
rect 252804 182454 253404 217898
rect 252804 182218 252986 182454
rect 253222 182218 253404 182454
rect 252804 182134 253404 182218
rect 252804 181898 252986 182134
rect 253222 181898 253404 182134
rect 252804 146454 253404 181898
rect 252804 146218 252986 146454
rect 253222 146218 253404 146454
rect 252804 146134 253404 146218
rect 252804 145898 252986 146134
rect 253222 145898 253404 146134
rect 252804 110454 253404 145898
rect 252804 110218 252986 110454
rect 253222 110218 253404 110454
rect 252804 110134 253404 110218
rect 252804 109898 252986 110134
rect 253222 109898 253404 110134
rect 252804 74454 253404 109898
rect 252804 74218 252986 74454
rect 253222 74218 253404 74454
rect 252804 74134 253404 74218
rect 252804 73898 252986 74134
rect 253222 73898 253404 74134
rect 252804 38454 253404 73898
rect 252804 38218 252986 38454
rect 253222 38218 253404 38454
rect 252804 38134 253404 38218
rect 252804 37898 252986 38134
rect 253222 37898 253404 38134
rect 252804 2454 253404 37898
rect 252804 2218 252986 2454
rect 253222 2218 253404 2454
rect 252804 2134 253404 2218
rect 252804 1898 252986 2134
rect 253222 1898 253404 2134
rect 252804 -346 253404 1898
rect 252804 -582 252986 -346
rect 253222 -582 253404 -346
rect 252804 -666 253404 -582
rect 252804 -902 252986 -666
rect 253222 -902 253404 -666
rect 252804 -1864 253404 -902
rect 256404 222054 257004 237000
rect 256404 221818 256586 222054
rect 256822 221818 257004 222054
rect 256404 221734 257004 221818
rect 256404 221498 256586 221734
rect 256822 221498 257004 221734
rect 256404 186054 257004 221498
rect 256404 185818 256586 186054
rect 256822 185818 257004 186054
rect 256404 185734 257004 185818
rect 256404 185498 256586 185734
rect 256822 185498 257004 185734
rect 256404 150054 257004 185498
rect 256404 149818 256586 150054
rect 256822 149818 257004 150054
rect 256404 149734 257004 149818
rect 256404 149498 256586 149734
rect 256822 149498 257004 149734
rect 256404 114054 257004 149498
rect 256404 113818 256586 114054
rect 256822 113818 257004 114054
rect 256404 113734 257004 113818
rect 256404 113498 256586 113734
rect 256822 113498 257004 113734
rect 256404 78054 257004 113498
rect 256404 77818 256586 78054
rect 256822 77818 257004 78054
rect 256404 77734 257004 77818
rect 256404 77498 256586 77734
rect 256822 77498 257004 77734
rect 256404 42054 257004 77498
rect 256404 41818 256586 42054
rect 256822 41818 257004 42054
rect 256404 41734 257004 41818
rect 256404 41498 256586 41734
rect 256822 41498 257004 41734
rect 256404 6054 257004 41498
rect 256404 5818 256586 6054
rect 256822 5818 257004 6054
rect 256404 5734 257004 5818
rect 256404 5498 256586 5734
rect 256822 5498 257004 5734
rect 256404 -2226 257004 5498
rect 256404 -2462 256586 -2226
rect 256822 -2462 257004 -2226
rect 256404 -2546 257004 -2462
rect 256404 -2782 256586 -2546
rect 256822 -2782 257004 -2546
rect 256404 -3744 257004 -2782
rect 260004 225654 260604 237000
rect 260004 225418 260186 225654
rect 260422 225418 260604 225654
rect 260004 225334 260604 225418
rect 260004 225098 260186 225334
rect 260422 225098 260604 225334
rect 260004 189654 260604 225098
rect 260004 189418 260186 189654
rect 260422 189418 260604 189654
rect 260004 189334 260604 189418
rect 260004 189098 260186 189334
rect 260422 189098 260604 189334
rect 260004 153654 260604 189098
rect 260004 153418 260186 153654
rect 260422 153418 260604 153654
rect 260004 153334 260604 153418
rect 260004 153098 260186 153334
rect 260422 153098 260604 153334
rect 260004 117654 260604 153098
rect 260004 117418 260186 117654
rect 260422 117418 260604 117654
rect 260004 117334 260604 117418
rect 260004 117098 260186 117334
rect 260422 117098 260604 117334
rect 260004 81654 260604 117098
rect 260004 81418 260186 81654
rect 260422 81418 260604 81654
rect 260004 81334 260604 81418
rect 260004 81098 260186 81334
rect 260422 81098 260604 81334
rect 260004 45654 260604 81098
rect 260004 45418 260186 45654
rect 260422 45418 260604 45654
rect 260004 45334 260604 45418
rect 260004 45098 260186 45334
rect 260422 45098 260604 45334
rect 260004 9654 260604 45098
rect 260004 9418 260186 9654
rect 260422 9418 260604 9654
rect 260004 9334 260604 9418
rect 260004 9098 260186 9334
rect 260422 9098 260604 9334
rect 260004 -4106 260604 9098
rect 260004 -4342 260186 -4106
rect 260422 -4342 260604 -4106
rect 260004 -4426 260604 -4342
rect 260004 -4662 260186 -4426
rect 260422 -4662 260604 -4426
rect 260004 -5624 260604 -4662
rect 263604 229254 264204 237000
rect 263604 229018 263786 229254
rect 264022 229018 264204 229254
rect 263604 228934 264204 229018
rect 263604 228698 263786 228934
rect 264022 228698 264204 228934
rect 263604 193254 264204 228698
rect 263604 193018 263786 193254
rect 264022 193018 264204 193254
rect 263604 192934 264204 193018
rect 263604 192698 263786 192934
rect 264022 192698 264204 192934
rect 263604 157254 264204 192698
rect 263604 157018 263786 157254
rect 264022 157018 264204 157254
rect 263604 156934 264204 157018
rect 263604 156698 263786 156934
rect 264022 156698 264204 156934
rect 263604 121254 264204 156698
rect 263604 121018 263786 121254
rect 264022 121018 264204 121254
rect 263604 120934 264204 121018
rect 263604 120698 263786 120934
rect 264022 120698 264204 120934
rect 263604 85254 264204 120698
rect 263604 85018 263786 85254
rect 264022 85018 264204 85254
rect 263604 84934 264204 85018
rect 263604 84698 263786 84934
rect 264022 84698 264204 84934
rect 263604 49254 264204 84698
rect 263604 49018 263786 49254
rect 264022 49018 264204 49254
rect 263604 48934 264204 49018
rect 263604 48698 263786 48934
rect 264022 48698 264204 48934
rect 263604 13254 264204 48698
rect 263604 13018 263786 13254
rect 264022 13018 264204 13254
rect 263604 12934 264204 13018
rect 263604 12698 263786 12934
rect 264022 12698 264204 12934
rect 245604 -7162 245786 -6926
rect 246022 -7162 246204 -6926
rect 245604 -7246 246204 -7162
rect 245604 -7482 245786 -7246
rect 246022 -7482 246204 -7246
rect 245604 -7504 246204 -7482
rect 263604 -5986 264204 12698
rect 270804 236454 271404 237000
rect 270804 236218 270986 236454
rect 271222 236218 271404 236454
rect 270804 236134 271404 236218
rect 270804 235898 270986 236134
rect 271222 235898 271404 236134
rect 270804 200454 271404 235898
rect 270804 200218 270986 200454
rect 271222 200218 271404 200454
rect 270804 200134 271404 200218
rect 270804 199898 270986 200134
rect 271222 199898 271404 200134
rect 270804 164454 271404 199898
rect 270804 164218 270986 164454
rect 271222 164218 271404 164454
rect 270804 164134 271404 164218
rect 270804 163898 270986 164134
rect 271222 163898 271404 164134
rect 270804 128454 271404 163898
rect 270804 128218 270986 128454
rect 271222 128218 271404 128454
rect 270804 128134 271404 128218
rect 270804 127898 270986 128134
rect 271222 127898 271404 128134
rect 270804 92454 271404 127898
rect 270804 92218 270986 92454
rect 271222 92218 271404 92454
rect 270804 92134 271404 92218
rect 270804 91898 270986 92134
rect 271222 91898 271404 92134
rect 270804 56454 271404 91898
rect 270804 56218 270986 56454
rect 271222 56218 271404 56454
rect 270804 56134 271404 56218
rect 270804 55898 270986 56134
rect 271222 55898 271404 56134
rect 270804 20454 271404 55898
rect 270804 20218 270986 20454
rect 271222 20218 271404 20454
rect 270804 20134 271404 20218
rect 270804 19898 270986 20134
rect 271222 19898 271404 20134
rect 270804 -1286 271404 19898
rect 270804 -1522 270986 -1286
rect 271222 -1522 271404 -1286
rect 270804 -1606 271404 -1522
rect 270804 -1842 270986 -1606
rect 271222 -1842 271404 -1606
rect 270804 -1864 271404 -1842
rect 274404 204054 275004 237000
rect 274404 203818 274586 204054
rect 274822 203818 275004 204054
rect 274404 203734 275004 203818
rect 274404 203498 274586 203734
rect 274822 203498 275004 203734
rect 274404 168054 275004 203498
rect 274404 167818 274586 168054
rect 274822 167818 275004 168054
rect 274404 167734 275004 167818
rect 274404 167498 274586 167734
rect 274822 167498 275004 167734
rect 274404 132054 275004 167498
rect 274404 131818 274586 132054
rect 274822 131818 275004 132054
rect 274404 131734 275004 131818
rect 274404 131498 274586 131734
rect 274822 131498 275004 131734
rect 274404 96054 275004 131498
rect 274404 95818 274586 96054
rect 274822 95818 275004 96054
rect 274404 95734 275004 95818
rect 274404 95498 274586 95734
rect 274822 95498 275004 95734
rect 274404 60054 275004 95498
rect 274404 59818 274586 60054
rect 274822 59818 275004 60054
rect 274404 59734 275004 59818
rect 274404 59498 274586 59734
rect 274822 59498 275004 59734
rect 274404 24054 275004 59498
rect 274404 23818 274586 24054
rect 274822 23818 275004 24054
rect 274404 23734 275004 23818
rect 274404 23498 274586 23734
rect 274822 23498 275004 23734
rect 274404 -3166 275004 23498
rect 274404 -3402 274586 -3166
rect 274822 -3402 275004 -3166
rect 274404 -3486 275004 -3402
rect 274404 -3722 274586 -3486
rect 274822 -3722 275004 -3486
rect 274404 -3744 275004 -3722
rect 278004 207654 278604 237000
rect 278004 207418 278186 207654
rect 278422 207418 278604 207654
rect 278004 207334 278604 207418
rect 278004 207098 278186 207334
rect 278422 207098 278604 207334
rect 278004 171654 278604 207098
rect 278004 171418 278186 171654
rect 278422 171418 278604 171654
rect 278004 171334 278604 171418
rect 278004 171098 278186 171334
rect 278422 171098 278604 171334
rect 278004 135654 278604 171098
rect 278004 135418 278186 135654
rect 278422 135418 278604 135654
rect 278004 135334 278604 135418
rect 278004 135098 278186 135334
rect 278422 135098 278604 135334
rect 278004 99654 278604 135098
rect 278004 99418 278186 99654
rect 278422 99418 278604 99654
rect 278004 99334 278604 99418
rect 278004 99098 278186 99334
rect 278422 99098 278604 99334
rect 278004 63654 278604 99098
rect 278004 63418 278186 63654
rect 278422 63418 278604 63654
rect 278004 63334 278604 63418
rect 278004 63098 278186 63334
rect 278422 63098 278604 63334
rect 278004 27654 278604 63098
rect 278004 27418 278186 27654
rect 278422 27418 278604 27654
rect 278004 27334 278604 27418
rect 278004 27098 278186 27334
rect 278422 27098 278604 27334
rect 278004 -5046 278604 27098
rect 278004 -5282 278186 -5046
rect 278422 -5282 278604 -5046
rect 278004 -5366 278604 -5282
rect 278004 -5602 278186 -5366
rect 278422 -5602 278604 -5366
rect 278004 -5624 278604 -5602
rect 281604 211254 282204 237000
rect 281604 211018 281786 211254
rect 282022 211018 282204 211254
rect 281604 210934 282204 211018
rect 281604 210698 281786 210934
rect 282022 210698 282204 210934
rect 281604 175254 282204 210698
rect 281604 175018 281786 175254
rect 282022 175018 282204 175254
rect 281604 174934 282204 175018
rect 281604 174698 281786 174934
rect 282022 174698 282204 174934
rect 281604 139254 282204 174698
rect 281604 139018 281786 139254
rect 282022 139018 282204 139254
rect 281604 138934 282204 139018
rect 281604 138698 281786 138934
rect 282022 138698 282204 138934
rect 281604 103254 282204 138698
rect 281604 103018 281786 103254
rect 282022 103018 282204 103254
rect 281604 102934 282204 103018
rect 281604 102698 281786 102934
rect 282022 102698 282204 102934
rect 281604 67254 282204 102698
rect 281604 67018 281786 67254
rect 282022 67018 282204 67254
rect 281604 66934 282204 67018
rect 281604 66698 281786 66934
rect 282022 66698 282204 66934
rect 281604 31254 282204 66698
rect 281604 31018 281786 31254
rect 282022 31018 282204 31254
rect 281604 30934 282204 31018
rect 281604 30698 281786 30934
rect 282022 30698 282204 30934
rect 263604 -6222 263786 -5986
rect 264022 -6222 264204 -5986
rect 263604 -6306 264204 -6222
rect 263604 -6542 263786 -6306
rect 264022 -6542 264204 -6306
rect 263604 -7504 264204 -6542
rect 281604 -6926 282204 30698
rect 288804 218454 289404 237000
rect 288804 218218 288986 218454
rect 289222 218218 289404 218454
rect 288804 218134 289404 218218
rect 288804 217898 288986 218134
rect 289222 217898 289404 218134
rect 288804 182454 289404 217898
rect 288804 182218 288986 182454
rect 289222 182218 289404 182454
rect 288804 182134 289404 182218
rect 288804 181898 288986 182134
rect 289222 181898 289404 182134
rect 288804 146454 289404 181898
rect 288804 146218 288986 146454
rect 289222 146218 289404 146454
rect 288804 146134 289404 146218
rect 288804 145898 288986 146134
rect 289222 145898 289404 146134
rect 288804 110454 289404 145898
rect 288804 110218 288986 110454
rect 289222 110218 289404 110454
rect 288804 110134 289404 110218
rect 288804 109898 288986 110134
rect 289222 109898 289404 110134
rect 288804 74454 289404 109898
rect 288804 74218 288986 74454
rect 289222 74218 289404 74454
rect 288804 74134 289404 74218
rect 288804 73898 288986 74134
rect 289222 73898 289404 74134
rect 288804 38454 289404 73898
rect 288804 38218 288986 38454
rect 289222 38218 289404 38454
rect 288804 38134 289404 38218
rect 288804 37898 288986 38134
rect 289222 37898 289404 38134
rect 288804 2454 289404 37898
rect 288804 2218 288986 2454
rect 289222 2218 289404 2454
rect 288804 2134 289404 2218
rect 288804 1898 288986 2134
rect 289222 1898 289404 2134
rect 288804 -346 289404 1898
rect 288804 -582 288986 -346
rect 289222 -582 289404 -346
rect 288804 -666 289404 -582
rect 288804 -902 288986 -666
rect 289222 -902 289404 -666
rect 288804 -1864 289404 -902
rect 292404 222054 293004 237000
rect 292404 221818 292586 222054
rect 292822 221818 293004 222054
rect 292404 221734 293004 221818
rect 292404 221498 292586 221734
rect 292822 221498 293004 221734
rect 292404 186054 293004 221498
rect 292404 185818 292586 186054
rect 292822 185818 293004 186054
rect 292404 185734 293004 185818
rect 292404 185498 292586 185734
rect 292822 185498 293004 185734
rect 292404 150054 293004 185498
rect 292404 149818 292586 150054
rect 292822 149818 293004 150054
rect 292404 149734 293004 149818
rect 292404 149498 292586 149734
rect 292822 149498 293004 149734
rect 292404 114054 293004 149498
rect 292404 113818 292586 114054
rect 292822 113818 293004 114054
rect 292404 113734 293004 113818
rect 292404 113498 292586 113734
rect 292822 113498 293004 113734
rect 292404 78054 293004 113498
rect 292404 77818 292586 78054
rect 292822 77818 293004 78054
rect 292404 77734 293004 77818
rect 292404 77498 292586 77734
rect 292822 77498 293004 77734
rect 292404 42054 293004 77498
rect 292404 41818 292586 42054
rect 292822 41818 293004 42054
rect 292404 41734 293004 41818
rect 292404 41498 292586 41734
rect 292822 41498 293004 41734
rect 292404 6054 293004 41498
rect 292404 5818 292586 6054
rect 292822 5818 293004 6054
rect 292404 5734 293004 5818
rect 292404 5498 292586 5734
rect 292822 5498 293004 5734
rect 292404 -2226 293004 5498
rect 292404 -2462 292586 -2226
rect 292822 -2462 293004 -2226
rect 292404 -2546 293004 -2462
rect 292404 -2782 292586 -2546
rect 292822 -2782 293004 -2546
rect 292404 -3744 293004 -2782
rect 296004 225654 296604 237000
rect 296004 225418 296186 225654
rect 296422 225418 296604 225654
rect 296004 225334 296604 225418
rect 296004 225098 296186 225334
rect 296422 225098 296604 225334
rect 296004 189654 296604 225098
rect 299604 229254 300204 237000
rect 299604 229018 299786 229254
rect 300022 229018 300204 229254
rect 299604 228934 300204 229018
rect 299604 228698 299786 228934
rect 300022 228698 300204 228934
rect 299604 204247 300204 228698
rect 306804 236454 307404 237000
rect 306804 236218 306986 236454
rect 307222 236218 307404 236454
rect 306804 236134 307404 236218
rect 306804 235898 306986 236134
rect 307222 235898 307404 236134
rect 306804 204247 307404 235898
rect 310404 204247 311004 237000
rect 314004 207654 314604 237000
rect 314004 207418 314186 207654
rect 314422 207418 314604 207654
rect 314004 207334 314604 207418
rect 314004 207098 314186 207334
rect 314422 207098 314604 207334
rect 314004 204247 314604 207098
rect 317604 211254 318204 237000
rect 317604 211018 317786 211254
rect 318022 211018 318204 211254
rect 317604 210934 318204 211018
rect 317604 210698 317786 210934
rect 318022 210698 318204 210934
rect 317604 204247 318204 210698
rect 324804 218454 325404 237000
rect 324804 218218 324986 218454
rect 325222 218218 325404 218454
rect 324804 218134 325404 218218
rect 324804 217898 324986 218134
rect 325222 217898 325404 218134
rect 324804 204247 325404 217898
rect 328404 222054 329004 237000
rect 328404 221818 328586 222054
rect 328822 221818 329004 222054
rect 328404 221734 329004 221818
rect 328404 221498 328586 221734
rect 328822 221498 329004 221734
rect 328404 204247 329004 221498
rect 332004 225654 332604 237000
rect 332004 225418 332186 225654
rect 332422 225418 332604 225654
rect 332004 225334 332604 225418
rect 332004 225098 332186 225334
rect 332422 225098 332604 225334
rect 332004 204247 332604 225098
rect 335604 229254 336204 237000
rect 335604 229018 335786 229254
rect 336022 229018 336204 229254
rect 335604 228934 336204 229018
rect 335604 228698 335786 228934
rect 336022 228698 336204 228934
rect 335604 204247 336204 228698
rect 342804 236454 343404 237000
rect 342804 236218 342986 236454
rect 343222 236218 343404 236454
rect 342804 236134 343404 236218
rect 342804 235898 342986 236134
rect 343222 235898 343404 236134
rect 342804 204247 343404 235898
rect 346404 204247 347004 237000
rect 350004 207654 350604 237000
rect 350004 207418 350186 207654
rect 350422 207418 350604 207654
rect 350004 207334 350604 207418
rect 350004 207098 350186 207334
rect 350422 207098 350604 207334
rect 350004 204247 350604 207098
rect 353604 211254 354204 237000
rect 353604 211018 353786 211254
rect 354022 211018 354204 211254
rect 353604 210934 354204 211018
rect 353604 210698 353786 210934
rect 354022 210698 354204 210934
rect 353604 204247 354204 210698
rect 360804 218454 361404 237000
rect 360804 218218 360986 218454
rect 361222 218218 361404 218454
rect 360804 218134 361404 218218
rect 360804 217898 360986 218134
rect 361222 217898 361404 218134
rect 360804 204247 361404 217898
rect 364404 222054 365004 237000
rect 364404 221818 364586 222054
rect 364822 221818 365004 222054
rect 364404 221734 365004 221818
rect 364404 221498 364586 221734
rect 364822 221498 365004 221734
rect 364404 204247 365004 221498
rect 368004 225654 368604 237000
rect 368004 225418 368186 225654
rect 368422 225418 368604 225654
rect 368004 225334 368604 225418
rect 368004 225098 368186 225334
rect 368422 225098 368604 225334
rect 368004 204247 368604 225098
rect 371604 229254 372204 237000
rect 371604 229018 371786 229254
rect 372022 229018 372204 229254
rect 371604 228934 372204 229018
rect 371604 228698 371786 228934
rect 372022 228698 372204 228934
rect 371604 204247 372204 228698
rect 378804 236454 379404 237000
rect 378804 236218 378986 236454
rect 379222 236218 379404 236454
rect 378804 236134 379404 236218
rect 378804 235898 378986 236134
rect 379222 235898 379404 236134
rect 378804 204247 379404 235898
rect 359227 204236 359293 204237
rect 359227 204172 359228 204236
rect 359292 204172 359293 204236
rect 359227 204171 359293 204172
rect 366035 204236 366101 204237
rect 366035 204172 366036 204236
rect 366100 204172 366101 204236
rect 366035 204171 366101 204172
rect 371003 204236 371069 204237
rect 371003 204172 371004 204236
rect 371068 204172 371069 204236
rect 371003 204171 371069 204172
rect 328131 203692 328197 203693
rect 328131 203628 328132 203692
rect 328196 203628 328197 203692
rect 328131 203627 328197 203628
rect 329419 203692 329485 203693
rect 329419 203628 329420 203692
rect 329484 203628 329485 203692
rect 329419 203627 329485 203628
rect 330707 203692 330773 203693
rect 330707 203628 330708 203692
rect 330772 203628 330773 203692
rect 330707 203627 330773 203628
rect 334939 203692 335005 203693
rect 334939 203628 334940 203692
rect 335004 203628 335005 203692
rect 334939 203627 335005 203628
rect 342851 203692 342917 203693
rect 342851 203628 342852 203692
rect 342916 203628 342917 203692
rect 342851 203627 342917 203628
rect 343955 203692 344021 203693
rect 343955 203628 343956 203692
rect 344020 203628 344021 203692
rect 343955 203627 344021 203628
rect 349107 203692 349173 203693
rect 349107 203628 349108 203692
rect 349172 203628 349173 203692
rect 349107 203627 349173 203628
rect 351131 203692 351197 203693
rect 351131 203628 351132 203692
rect 351196 203628 351197 203692
rect 351131 203627 351197 203628
rect 328134 200970 328194 203627
rect 328315 203420 328381 203421
rect 328315 203356 328316 203420
rect 328380 203356 328381 203420
rect 328315 203355 328381 203356
rect 328318 201650 328378 203355
rect 328318 201590 328446 201650
rect 328134 200910 328292 200970
rect 328386 200940 328446 201590
rect 329422 200910 329482 203627
rect 329603 203148 329669 203149
rect 329603 203084 329604 203148
rect 329668 203084 329669 203148
rect 329603 203083 329669 203084
rect 329606 200970 329666 203083
rect 330710 201650 330770 203627
rect 332363 203420 332429 203421
rect 332363 203356 332364 203420
rect 332428 203356 332429 203420
rect 332363 203355 332429 203356
rect 332915 203420 332981 203421
rect 332915 203356 332916 203420
rect 332980 203356 332981 203420
rect 332915 203355 332981 203356
rect 331075 203284 331141 203285
rect 331075 203220 331076 203284
rect 331140 203220 331141 203284
rect 331075 203219 331141 203220
rect 331627 203284 331693 203285
rect 331627 203220 331628 203284
rect 331692 203220 331693 203284
rect 331627 203219 331693 203220
rect 329584 200910 329666 200970
rect 330598 201590 330770 201650
rect 330598 200940 330658 201590
rect 331078 200970 331138 203219
rect 330752 200910 331138 200970
rect 331630 200970 331690 203219
rect 332366 200970 332426 203355
rect 331630 200910 331796 200970
rect 331920 200910 332426 200970
rect 332918 200910 332978 203355
rect 334019 203284 334085 203285
rect 334019 203220 334020 203284
rect 334084 203220 334085 203284
rect 334019 203219 334085 203220
rect 333651 203148 333717 203149
rect 333651 203084 333652 203148
rect 333716 203084 333717 203148
rect 333651 203083 333717 203084
rect 333654 200970 333714 203083
rect 334022 201650 334082 203219
rect 334755 203148 334821 203149
rect 334755 203084 334756 203148
rect 334820 203084 334821 203148
rect 334755 203083 334821 203084
rect 334022 201590 334162 201650
rect 333088 200910 333714 200970
rect 334102 200940 334162 201590
rect 334758 200970 334818 203083
rect 334256 200910 334818 200970
rect 334942 200970 335002 203627
rect 340091 203556 340157 203557
rect 340091 203492 340092 203556
rect 340156 203492 340157 203556
rect 340091 203491 340157 203492
rect 340827 203556 340893 203557
rect 340827 203492 340828 203556
rect 340892 203492 340893 203556
rect 340827 203491 340893 203492
rect 336595 203420 336661 203421
rect 336595 203356 336596 203420
rect 336660 203356 336661 203420
rect 336595 203355 336661 203356
rect 338251 203420 338317 203421
rect 338251 203356 338252 203420
rect 338316 203356 338317 203420
rect 338251 203355 338317 203356
rect 336227 203284 336293 203285
rect 336227 203220 336228 203284
rect 336292 203220 336293 203284
rect 336227 203219 336293 203220
rect 336043 203012 336109 203013
rect 336043 202948 336044 203012
rect 336108 202948 336109 203012
rect 336043 202947 336109 202948
rect 336046 200970 336106 202947
rect 334942 200910 335300 200970
rect 335424 200910 336106 200970
rect 336230 200970 336290 203219
rect 336598 200970 336658 203355
rect 336963 203284 337029 203285
rect 336963 203220 336964 203284
rect 337028 203220 337029 203284
rect 336963 203219 337029 203220
rect 336230 200910 336468 200970
rect 336592 200910 336658 200970
rect 336966 200970 337026 203219
rect 337883 203012 337949 203013
rect 337883 202948 337884 203012
rect 337948 202948 337949 203012
rect 337883 202947 337949 202948
rect 337886 200970 337946 202947
rect 336966 200910 337636 200970
rect 337760 200910 337946 200970
rect 338254 200970 338314 203355
rect 339539 203284 339605 203285
rect 339539 203220 339540 203284
rect 339604 203220 339605 203284
rect 339539 203219 339605 203220
rect 339171 203012 339237 203013
rect 339171 202948 339172 203012
rect 339236 202948 339237 203012
rect 339171 202947 339237 202948
rect 338254 200910 338804 200970
rect 339174 200817 339234 202947
rect 339542 200970 339602 203219
rect 339542 200910 339972 200970
rect 340094 200910 340154 203491
rect 338928 200757 339234 200817
rect 340830 200817 340890 203491
rect 341747 203148 341813 203149
rect 341747 203084 341748 203148
rect 341812 203084 341813 203148
rect 341747 203083 341813 203084
rect 341750 200970 341810 203083
rect 342299 203012 342365 203013
rect 342299 202948 342300 203012
rect 342364 202948 342365 203012
rect 342299 202947 342365 202948
rect 342483 203012 342549 203013
rect 342483 202948 342484 203012
rect 342548 202948 342549 203012
rect 342483 202947 342549 202948
rect 342302 201789 342362 202947
rect 342299 201788 342365 201789
rect 342299 201724 342300 201788
rect 342364 201724 342365 201788
rect 342299 201723 342365 201724
rect 342486 201650 342546 202947
rect 342402 201590 342546 201650
rect 342275 201516 342341 201517
rect 342275 201452 342276 201516
rect 342340 201452 342341 201516
rect 342275 201451 342341 201452
rect 341264 200910 341810 200970
rect 342278 200940 342338 201451
rect 342402 200940 342462 201590
rect 342854 200970 342914 203627
rect 343587 203012 343653 203013
rect 343587 202948 343588 203012
rect 343652 202948 343653 203012
rect 343587 202947 343653 202948
rect 342854 200910 343476 200970
rect 343590 200910 343650 202947
rect 343958 200970 344018 203627
rect 345243 203284 345309 203285
rect 345243 203220 345244 203284
rect 345308 203220 345309 203284
rect 345243 203219 345309 203220
rect 344875 203012 344941 203013
rect 344875 202948 344876 203012
rect 344940 202948 344941 203012
rect 344875 202947 344941 202948
rect 344878 200970 344938 202947
rect 343958 200910 344644 200970
rect 344768 200910 344938 200970
rect 345246 200970 345306 203219
rect 346531 203148 346597 203149
rect 346531 203084 346532 203148
rect 346596 203084 346597 203148
rect 346531 203083 346597 203084
rect 347819 203148 347885 203149
rect 347819 203084 347820 203148
rect 347884 203084 347885 203148
rect 347819 203083 347885 203084
rect 345979 203012 346045 203013
rect 345979 202948 345980 203012
rect 346044 202948 346045 203012
rect 345979 202947 346045 202948
rect 345982 201650 346042 202947
rect 345906 201590 346042 201650
rect 345246 200910 345812 200970
rect 345906 200940 345966 201590
rect 346534 200970 346594 203083
rect 347083 203012 347149 203013
rect 347083 202948 347084 203012
rect 347148 202948 347149 203012
rect 347083 202947 347149 202948
rect 346534 200910 346980 200970
rect 347086 200910 347146 202947
rect 347822 200970 347882 203083
rect 348371 203012 348437 203013
rect 348371 202948 348372 203012
rect 348436 202948 348437 203012
rect 348371 202947 348437 202948
rect 348374 200970 348434 202947
rect 347822 200910 348148 200970
rect 348272 200910 348434 200970
rect 349110 200970 349170 203627
rect 349843 203284 349909 203285
rect 349843 203220 349844 203284
rect 349908 203220 349909 203284
rect 349843 203219 349909 203220
rect 349659 203012 349725 203013
rect 349659 202948 349660 203012
rect 349724 202948 349725 203012
rect 349659 202947 349725 202948
rect 349110 200910 349316 200970
rect 349662 200817 349722 202947
rect 349846 200970 349906 203219
rect 350947 203012 351013 203013
rect 350947 202948 350948 203012
rect 351012 202948 351013 203012
rect 350947 202947 351013 202948
rect 350950 200970 351010 202947
rect 349846 200910 350484 200970
rect 350608 200910 351010 200970
rect 351134 200970 351194 203627
rect 357387 203420 357453 203421
rect 357387 203356 357388 203420
rect 357452 203356 357453 203420
rect 357387 203355 357453 203356
rect 352787 203148 352853 203149
rect 352787 203084 352788 203148
rect 352852 203084 352853 203148
rect 352787 203083 352853 203084
rect 353155 203148 353221 203149
rect 353155 203084 353156 203148
rect 353220 203084 353221 203148
rect 353155 203083 353221 203084
rect 354811 203148 354877 203149
rect 354811 203084 354812 203148
rect 354876 203084 354877 203148
rect 354811 203083 354877 203084
rect 356099 203148 356165 203149
rect 356099 203084 356100 203148
rect 356164 203084 356165 203148
rect 356099 203083 356165 203084
rect 351683 203012 351749 203013
rect 351683 202948 351684 203012
rect 351748 202948 351749 203012
rect 351683 202947 351749 202948
rect 351686 201650 351746 202947
rect 351686 201590 351806 201650
rect 351134 200910 351652 200970
rect 351746 200940 351806 201590
rect 352790 200940 352850 203083
rect 353158 200970 353218 203083
rect 353339 203012 353405 203013
rect 353339 202948 353340 203012
rect 353404 202948 353405 203012
rect 353339 202947 353405 202948
rect 354259 203012 354325 203013
rect 354259 202948 354260 203012
rect 354324 202948 354325 203012
rect 354259 202947 354325 202948
rect 352944 200910 353218 200970
rect 353342 200970 353402 202947
rect 354262 200970 354322 202947
rect 353342 200910 353988 200970
rect 354112 200910 354322 200970
rect 354814 200970 354874 203083
rect 355547 203012 355613 203013
rect 355547 202948 355548 203012
rect 355612 202948 355613 203012
rect 355547 202947 355613 202948
rect 354814 200910 355156 200970
rect 355550 200817 355610 202947
rect 356102 200970 356162 203083
rect 356467 203012 356533 203013
rect 356467 202948 356468 203012
rect 356532 202948 356533 203012
rect 356467 202947 356533 202948
rect 356470 200970 356530 202947
rect 357390 201650 357450 203355
rect 357755 203148 357821 203149
rect 357755 203084 357756 203148
rect 357820 203084 357821 203148
rect 357755 203083 357821 203084
rect 357390 201590 357522 201650
rect 356102 200910 356324 200970
rect 356448 200910 356530 200970
rect 357462 200940 357522 201590
rect 357758 200970 357818 203083
rect 357939 203012 358005 203013
rect 357939 202948 357940 203012
rect 358004 202948 358005 203012
rect 357939 202947 358005 202948
rect 358675 203012 358741 203013
rect 358675 202948 358676 203012
rect 358740 202948 358741 203012
rect 358675 202947 358741 202948
rect 357616 200910 357818 200970
rect 357942 200970 358002 202947
rect 358678 201650 358738 202947
rect 358678 201590 358814 201650
rect 357942 200910 358660 200970
rect 358754 200940 358814 201590
rect 359230 200970 359290 204171
rect 360331 204100 360397 204101
rect 360331 204036 360332 204100
rect 360396 204036 360397 204100
rect 360331 204035 360397 204036
rect 359963 203012 360029 203013
rect 359963 202948 359964 203012
rect 360028 202948 360029 203012
rect 359963 202947 360029 202948
rect 359966 200970 360026 202947
rect 359230 200910 359828 200970
rect 359952 200910 360026 200970
rect 360334 200970 360394 204035
rect 361619 203964 361685 203965
rect 361619 203900 361620 203964
rect 361684 203900 361685 203964
rect 361619 203899 361685 203900
rect 361251 203012 361317 203013
rect 361251 202948 361252 203012
rect 361316 202948 361317 203012
rect 361251 202947 361317 202948
rect 361254 200970 361314 202947
rect 360334 200910 360996 200970
rect 361120 200910 361314 200970
rect 361622 200970 361682 203899
rect 362907 203828 362973 203829
rect 362907 203764 362908 203828
rect 362972 203764 362973 203828
rect 362907 203763 362973 203764
rect 364379 203828 364445 203829
rect 364379 203764 364380 203828
rect 364444 203764 364445 203828
rect 364379 203763 364445 203764
rect 362539 203012 362605 203013
rect 362539 202948 362540 203012
rect 362604 202948 362605 203012
rect 362539 202947 362605 202948
rect 361622 200910 362164 200970
rect 362542 200817 362602 202947
rect 362910 200970 362970 203763
rect 363459 203012 363525 203013
rect 363459 202948 363460 203012
rect 363524 202948 363525 203012
rect 363459 202947 363525 202948
rect 363462 200970 363522 202947
rect 364382 201650 364442 203763
rect 364747 203012 364813 203013
rect 364747 202948 364748 203012
rect 364812 202948 364813 203012
rect 364747 202947 364813 202948
rect 364382 201590 364530 201650
rect 362910 200910 363332 200970
rect 363456 200910 363522 200970
rect 364470 200940 364530 201590
rect 364750 200970 364810 202947
rect 366038 200970 366098 204171
rect 367507 204100 367573 204101
rect 367507 204036 367508 204100
rect 367572 204036 367573 204100
rect 367507 204035 367573 204036
rect 366403 203964 366469 203965
rect 366403 203900 366404 203964
rect 366468 203900 366469 203964
rect 366403 203899 366469 203900
rect 364624 200910 364810 200970
rect 365792 200910 366098 200970
rect 366406 200970 366466 203899
rect 367510 200970 367570 204035
rect 368611 203284 368677 203285
rect 368611 203220 368612 203284
rect 368676 203220 368677 203284
rect 368611 203219 368677 203220
rect 368614 200970 368674 203219
rect 371006 200970 371066 204171
rect 382404 204054 383004 237000
rect 382404 203818 382586 204054
rect 382822 203818 383004 204054
rect 382404 203734 383004 203818
rect 382404 203498 382586 203734
rect 382822 203498 383004 203734
rect 373395 203148 373461 203149
rect 373395 203084 373396 203148
rect 373460 203084 373461 203148
rect 373395 203083 373461 203084
rect 366406 200910 366960 200970
rect 367510 200910 368128 200970
rect 368614 200910 369296 200970
rect 370464 200910 371066 200970
rect 373398 200970 373458 203083
rect 373398 200910 373463 200970
rect 340830 200757 341140 200817
rect 349440 200757 349722 200817
rect 355280 200757 355610 200817
rect 362288 200757 362602 200817
rect 296004 189418 296186 189654
rect 296422 189418 296604 189654
rect 296004 189334 296604 189418
rect 296004 189098 296186 189334
rect 296422 189098 296604 189334
rect 296004 153654 296604 189098
rect 300482 182454 300802 182476
rect 300482 182218 300524 182454
rect 300760 182218 300802 182454
rect 300482 182134 300802 182218
rect 300482 181898 300524 182134
rect 300760 181898 300802 182134
rect 300482 181876 300802 181898
rect 382404 168054 383004 203498
rect 382404 167818 382586 168054
rect 382822 167818 383004 168054
rect 382404 167734 383004 167818
rect 382404 167498 382586 167734
rect 382822 167498 383004 167734
rect 300034 164454 300358 164476
rect 300034 164218 300078 164454
rect 300314 164218 300358 164454
rect 300034 164134 300358 164218
rect 300034 163898 300078 164134
rect 300314 163898 300358 164134
rect 300034 163876 300358 163898
rect 296004 153418 296186 153654
rect 296422 153418 296604 153654
rect 296004 153334 296604 153418
rect 296004 153098 296186 153334
rect 296422 153098 296604 153334
rect 296004 117654 296604 153098
rect 300482 146454 300802 146476
rect 300482 146218 300524 146454
rect 300760 146218 300802 146454
rect 300482 146134 300802 146218
rect 300482 145898 300524 146134
rect 300760 145898 300802 146134
rect 300482 145876 300802 145898
rect 382404 132054 383004 167498
rect 382404 131818 382586 132054
rect 382822 131818 383004 132054
rect 382404 131734 383004 131818
rect 382404 131498 382586 131734
rect 382822 131498 383004 131734
rect 300034 128454 300358 128476
rect 300034 128218 300078 128454
rect 300314 128218 300358 128454
rect 300034 128134 300358 128218
rect 300034 127898 300078 128134
rect 300314 127898 300358 128134
rect 300034 127876 300358 127898
rect 296004 117418 296186 117654
rect 296422 117418 296604 117654
rect 296004 117334 296604 117418
rect 296004 117098 296186 117334
rect 296422 117098 296604 117334
rect 296004 81654 296604 117098
rect 303662 109037 303722 110190
rect 308078 110130 308688 110190
rect 308078 109037 308138 110130
rect 303659 109036 303725 109037
rect 303659 108972 303660 109036
rect 303724 108972 303725 109036
rect 303659 108971 303725 108972
rect 308075 109036 308141 109037
rect 308075 108972 308076 109036
rect 308140 108972 308141 109036
rect 308075 108971 308141 108972
rect 296004 81418 296186 81654
rect 296422 81418 296604 81654
rect 296004 81334 296604 81418
rect 296004 81098 296186 81334
rect 296422 81098 296604 81334
rect 296004 45654 296604 81098
rect 296004 45418 296186 45654
rect 296422 45418 296604 45654
rect 296004 45334 296604 45418
rect 296004 45098 296186 45334
rect 296422 45098 296604 45334
rect 296004 9654 296604 45098
rect 296004 9418 296186 9654
rect 296422 9418 296604 9654
rect 296004 9334 296604 9418
rect 296004 9098 296186 9334
rect 296422 9098 296604 9334
rect 296004 -4106 296604 9098
rect 296004 -4342 296186 -4106
rect 296422 -4342 296604 -4106
rect 296004 -4426 296604 -4342
rect 296004 -4662 296186 -4426
rect 296422 -4662 296604 -4426
rect 296004 -5624 296604 -4662
rect 299604 85254 300204 107000
rect 299604 85018 299786 85254
rect 300022 85018 300204 85254
rect 299604 84934 300204 85018
rect 299604 84698 299786 84934
rect 300022 84698 300204 84934
rect 299604 49254 300204 84698
rect 299604 49018 299786 49254
rect 300022 49018 300204 49254
rect 299604 48934 300204 49018
rect 299604 48698 299786 48934
rect 300022 48698 300204 48934
rect 299604 13254 300204 48698
rect 299604 13018 299786 13254
rect 300022 13018 300204 13254
rect 299604 12934 300204 13018
rect 299604 12698 299786 12934
rect 300022 12698 300204 12934
rect 281604 -7162 281786 -6926
rect 282022 -7162 282204 -6926
rect 281604 -7246 282204 -7162
rect 281604 -7482 281786 -7246
rect 282022 -7482 282204 -7246
rect 281604 -7504 282204 -7482
rect 299604 -5986 300204 12698
rect 306804 92454 307404 107000
rect 306804 92218 306986 92454
rect 307222 92218 307404 92454
rect 306804 92134 307404 92218
rect 306804 91898 306986 92134
rect 307222 91898 307404 92134
rect 306804 56454 307404 91898
rect 306804 56218 306986 56454
rect 307222 56218 307404 56454
rect 306804 56134 307404 56218
rect 306804 55898 306986 56134
rect 307222 55898 307404 56134
rect 306804 20454 307404 55898
rect 306804 20218 306986 20454
rect 307222 20218 307404 20454
rect 306804 20134 307404 20218
rect 306804 19898 306986 20134
rect 307222 19898 307404 20134
rect 306804 -1286 307404 19898
rect 306804 -1522 306986 -1286
rect 307222 -1522 307404 -1286
rect 306804 -1606 307404 -1522
rect 306804 -1842 306986 -1606
rect 307222 -1842 307404 -1606
rect 306804 -1864 307404 -1842
rect 310404 96054 311004 107000
rect 310404 95818 310586 96054
rect 310822 95818 311004 96054
rect 310404 95734 311004 95818
rect 310404 95498 310586 95734
rect 310822 95498 311004 95734
rect 310404 60054 311004 95498
rect 310404 59818 310586 60054
rect 310822 59818 311004 60054
rect 310404 59734 311004 59818
rect 310404 59498 310586 59734
rect 310822 59498 311004 59734
rect 310404 24054 311004 59498
rect 310404 23818 310586 24054
rect 310822 23818 311004 24054
rect 310404 23734 311004 23818
rect 310404 23498 310586 23734
rect 310822 23498 311004 23734
rect 310404 -3166 311004 23498
rect 310404 -3402 310586 -3166
rect 310822 -3402 311004 -3166
rect 310404 -3486 311004 -3402
rect 310404 -3722 310586 -3486
rect 310822 -3722 311004 -3486
rect 310404 -3744 311004 -3722
rect 314004 99654 314604 107000
rect 314004 99418 314186 99654
rect 314422 99418 314604 99654
rect 314004 99334 314604 99418
rect 314004 99098 314186 99334
rect 314422 99098 314604 99334
rect 314004 63654 314604 99098
rect 314004 63418 314186 63654
rect 314422 63418 314604 63654
rect 314004 63334 314604 63418
rect 314004 63098 314186 63334
rect 314422 63098 314604 63334
rect 314004 27654 314604 63098
rect 314004 27418 314186 27654
rect 314422 27418 314604 27654
rect 314004 27334 314604 27418
rect 314004 27098 314186 27334
rect 314422 27098 314604 27334
rect 314004 -5046 314604 27098
rect 314004 -5282 314186 -5046
rect 314422 -5282 314604 -5046
rect 314004 -5366 314604 -5282
rect 314004 -5602 314186 -5366
rect 314422 -5602 314604 -5366
rect 314004 -5624 314604 -5602
rect 317604 103254 318204 107000
rect 317604 103018 317786 103254
rect 318022 103018 318204 103254
rect 317604 102934 318204 103018
rect 317604 102698 317786 102934
rect 318022 102698 318204 102934
rect 317604 67254 318204 102698
rect 317604 67018 317786 67254
rect 318022 67018 318204 67254
rect 317604 66934 318204 67018
rect 317604 66698 317786 66934
rect 318022 66698 318204 66934
rect 317604 31254 318204 66698
rect 317604 31018 317786 31254
rect 318022 31018 318204 31254
rect 317604 30934 318204 31018
rect 317604 30698 317786 30934
rect 318022 30698 318204 30934
rect 299604 -6222 299786 -5986
rect 300022 -6222 300204 -5986
rect 299604 -6306 300204 -6222
rect 299604 -6542 299786 -6306
rect 300022 -6542 300204 -6306
rect 299604 -7504 300204 -6542
rect 317604 -6926 318204 30698
rect 324804 74454 325404 107000
rect 324804 74218 324986 74454
rect 325222 74218 325404 74454
rect 324804 74134 325404 74218
rect 324804 73898 324986 74134
rect 325222 73898 325404 74134
rect 324804 38454 325404 73898
rect 324804 38218 324986 38454
rect 325222 38218 325404 38454
rect 324804 38134 325404 38218
rect 324804 37898 324986 38134
rect 325222 37898 325404 38134
rect 324804 2454 325404 37898
rect 324804 2218 324986 2454
rect 325222 2218 325404 2454
rect 324804 2134 325404 2218
rect 324804 1898 324986 2134
rect 325222 1898 325404 2134
rect 324804 -346 325404 1898
rect 324804 -582 324986 -346
rect 325222 -582 325404 -346
rect 324804 -666 325404 -582
rect 324804 -902 324986 -666
rect 325222 -902 325404 -666
rect 324804 -1864 325404 -902
rect 328404 78054 329004 107000
rect 328404 77818 328586 78054
rect 328822 77818 329004 78054
rect 328404 77734 329004 77818
rect 328404 77498 328586 77734
rect 328822 77498 329004 77734
rect 328404 42054 329004 77498
rect 328404 41818 328586 42054
rect 328822 41818 329004 42054
rect 328404 41734 329004 41818
rect 328404 41498 328586 41734
rect 328822 41498 329004 41734
rect 328404 6054 329004 41498
rect 328404 5818 328586 6054
rect 328822 5818 329004 6054
rect 328404 5734 329004 5818
rect 328404 5498 328586 5734
rect 328822 5498 329004 5734
rect 328404 -2226 329004 5498
rect 328404 -2462 328586 -2226
rect 328822 -2462 329004 -2226
rect 328404 -2546 329004 -2462
rect 328404 -2782 328586 -2546
rect 328822 -2782 329004 -2546
rect 328404 -3744 329004 -2782
rect 332004 81654 332604 107000
rect 332004 81418 332186 81654
rect 332422 81418 332604 81654
rect 332004 81334 332604 81418
rect 332004 81098 332186 81334
rect 332422 81098 332604 81334
rect 332004 45654 332604 81098
rect 332004 45418 332186 45654
rect 332422 45418 332604 45654
rect 332004 45334 332604 45418
rect 332004 45098 332186 45334
rect 332422 45098 332604 45334
rect 332004 9654 332604 45098
rect 332004 9418 332186 9654
rect 332422 9418 332604 9654
rect 332004 9334 332604 9418
rect 332004 9098 332186 9334
rect 332422 9098 332604 9334
rect 332004 -4106 332604 9098
rect 332004 -4342 332186 -4106
rect 332422 -4342 332604 -4106
rect 332004 -4426 332604 -4342
rect 332004 -4662 332186 -4426
rect 332422 -4662 332604 -4426
rect 332004 -5624 332604 -4662
rect 335604 85254 336204 107000
rect 335604 85018 335786 85254
rect 336022 85018 336204 85254
rect 335604 84934 336204 85018
rect 335604 84698 335786 84934
rect 336022 84698 336204 84934
rect 335604 49254 336204 84698
rect 335604 49018 335786 49254
rect 336022 49018 336204 49254
rect 335604 48934 336204 49018
rect 335604 48698 335786 48934
rect 336022 48698 336204 48934
rect 335604 13254 336204 48698
rect 335604 13018 335786 13254
rect 336022 13018 336204 13254
rect 335604 12934 336204 13018
rect 335604 12698 335786 12934
rect 336022 12698 336204 12934
rect 317604 -7162 317786 -6926
rect 318022 -7162 318204 -6926
rect 317604 -7246 318204 -7162
rect 317604 -7482 317786 -7246
rect 318022 -7482 318204 -7246
rect 317604 -7504 318204 -7482
rect 335604 -5986 336204 12698
rect 342804 92454 343404 107000
rect 342804 92218 342986 92454
rect 343222 92218 343404 92454
rect 342804 92134 343404 92218
rect 342804 91898 342986 92134
rect 343222 91898 343404 92134
rect 342804 56454 343404 91898
rect 342804 56218 342986 56454
rect 343222 56218 343404 56454
rect 342804 56134 343404 56218
rect 342804 55898 342986 56134
rect 343222 55898 343404 56134
rect 342804 20454 343404 55898
rect 342804 20218 342986 20454
rect 343222 20218 343404 20454
rect 342804 20134 343404 20218
rect 342804 19898 342986 20134
rect 343222 19898 343404 20134
rect 342804 -1286 343404 19898
rect 342804 -1522 342986 -1286
rect 343222 -1522 343404 -1286
rect 342804 -1606 343404 -1522
rect 342804 -1842 342986 -1606
rect 343222 -1842 343404 -1606
rect 342804 -1864 343404 -1842
rect 346404 96054 347004 107000
rect 346404 95818 346586 96054
rect 346822 95818 347004 96054
rect 346404 95734 347004 95818
rect 346404 95498 346586 95734
rect 346822 95498 347004 95734
rect 346404 60054 347004 95498
rect 346404 59818 346586 60054
rect 346822 59818 347004 60054
rect 346404 59734 347004 59818
rect 346404 59498 346586 59734
rect 346822 59498 347004 59734
rect 346404 24054 347004 59498
rect 346404 23818 346586 24054
rect 346822 23818 347004 24054
rect 346404 23734 347004 23818
rect 346404 23498 346586 23734
rect 346822 23498 347004 23734
rect 346404 -3166 347004 23498
rect 346404 -3402 346586 -3166
rect 346822 -3402 347004 -3166
rect 346404 -3486 347004 -3402
rect 346404 -3722 346586 -3486
rect 346822 -3722 347004 -3486
rect 346404 -3744 347004 -3722
rect 350004 99654 350604 107000
rect 350004 99418 350186 99654
rect 350422 99418 350604 99654
rect 350004 99334 350604 99418
rect 350004 99098 350186 99334
rect 350422 99098 350604 99334
rect 350004 63654 350604 99098
rect 350004 63418 350186 63654
rect 350422 63418 350604 63654
rect 350004 63334 350604 63418
rect 350004 63098 350186 63334
rect 350422 63098 350604 63334
rect 350004 27654 350604 63098
rect 350004 27418 350186 27654
rect 350422 27418 350604 27654
rect 350004 27334 350604 27418
rect 350004 27098 350186 27334
rect 350422 27098 350604 27334
rect 350004 -5046 350604 27098
rect 350004 -5282 350186 -5046
rect 350422 -5282 350604 -5046
rect 350004 -5366 350604 -5282
rect 350004 -5602 350186 -5366
rect 350422 -5602 350604 -5366
rect 350004 -5624 350604 -5602
rect 353604 103254 354204 107000
rect 353604 103018 353786 103254
rect 354022 103018 354204 103254
rect 353604 102934 354204 103018
rect 353604 102698 353786 102934
rect 354022 102698 354204 102934
rect 353604 67254 354204 102698
rect 353604 67018 353786 67254
rect 354022 67018 354204 67254
rect 353604 66934 354204 67018
rect 353604 66698 353786 66934
rect 354022 66698 354204 66934
rect 353604 31254 354204 66698
rect 353604 31018 353786 31254
rect 354022 31018 354204 31254
rect 353604 30934 354204 31018
rect 353604 30698 353786 30934
rect 354022 30698 354204 30934
rect 335604 -6222 335786 -5986
rect 336022 -6222 336204 -5986
rect 335604 -6306 336204 -6222
rect 335604 -6542 335786 -6306
rect 336022 -6542 336204 -6306
rect 335604 -7504 336204 -6542
rect 353604 -6926 354204 30698
rect 360804 74454 361404 107000
rect 360804 74218 360986 74454
rect 361222 74218 361404 74454
rect 360804 74134 361404 74218
rect 360804 73898 360986 74134
rect 361222 73898 361404 74134
rect 360804 38454 361404 73898
rect 360804 38218 360986 38454
rect 361222 38218 361404 38454
rect 360804 38134 361404 38218
rect 360804 37898 360986 38134
rect 361222 37898 361404 38134
rect 360804 2454 361404 37898
rect 360804 2218 360986 2454
rect 361222 2218 361404 2454
rect 360804 2134 361404 2218
rect 360804 1898 360986 2134
rect 361222 1898 361404 2134
rect 360804 -346 361404 1898
rect 360804 -582 360986 -346
rect 361222 -582 361404 -346
rect 360804 -666 361404 -582
rect 360804 -902 360986 -666
rect 361222 -902 361404 -666
rect 360804 -1864 361404 -902
rect 364404 78054 365004 107000
rect 364404 77818 364586 78054
rect 364822 77818 365004 78054
rect 364404 77734 365004 77818
rect 364404 77498 364586 77734
rect 364822 77498 365004 77734
rect 364404 42054 365004 77498
rect 364404 41818 364586 42054
rect 364822 41818 365004 42054
rect 364404 41734 365004 41818
rect 364404 41498 364586 41734
rect 364822 41498 365004 41734
rect 364404 6054 365004 41498
rect 364404 5818 364586 6054
rect 364822 5818 365004 6054
rect 364404 5734 365004 5818
rect 364404 5498 364586 5734
rect 364822 5498 365004 5734
rect 364404 -2226 365004 5498
rect 364404 -2462 364586 -2226
rect 364822 -2462 365004 -2226
rect 364404 -2546 365004 -2462
rect 364404 -2782 364586 -2546
rect 364822 -2782 365004 -2546
rect 364404 -3744 365004 -2782
rect 368004 81654 368604 107000
rect 368004 81418 368186 81654
rect 368422 81418 368604 81654
rect 368004 81334 368604 81418
rect 368004 81098 368186 81334
rect 368422 81098 368604 81334
rect 368004 45654 368604 81098
rect 368004 45418 368186 45654
rect 368422 45418 368604 45654
rect 368004 45334 368604 45418
rect 368004 45098 368186 45334
rect 368422 45098 368604 45334
rect 368004 9654 368604 45098
rect 368004 9418 368186 9654
rect 368422 9418 368604 9654
rect 368004 9334 368604 9418
rect 368004 9098 368186 9334
rect 368422 9098 368604 9334
rect 368004 -4106 368604 9098
rect 368004 -4342 368186 -4106
rect 368422 -4342 368604 -4106
rect 368004 -4426 368604 -4342
rect 368004 -4662 368186 -4426
rect 368422 -4662 368604 -4426
rect 368004 -5624 368604 -4662
rect 371604 85254 372204 107000
rect 371604 85018 371786 85254
rect 372022 85018 372204 85254
rect 371604 84934 372204 85018
rect 371604 84698 371786 84934
rect 372022 84698 372204 84934
rect 371604 49254 372204 84698
rect 371604 49018 371786 49254
rect 372022 49018 372204 49254
rect 371604 48934 372204 49018
rect 371604 48698 371786 48934
rect 372022 48698 372204 48934
rect 371604 13254 372204 48698
rect 371604 13018 371786 13254
rect 372022 13018 372204 13254
rect 371604 12934 372204 13018
rect 371604 12698 371786 12934
rect 372022 12698 372204 12934
rect 353604 -7162 353786 -6926
rect 354022 -7162 354204 -6926
rect 353604 -7246 354204 -7162
rect 353604 -7482 353786 -7246
rect 354022 -7482 354204 -7246
rect 353604 -7504 354204 -7482
rect 371604 -5986 372204 12698
rect 378804 92454 379404 107000
rect 378804 92218 378986 92454
rect 379222 92218 379404 92454
rect 378804 92134 379404 92218
rect 378804 91898 378986 92134
rect 379222 91898 379404 92134
rect 378804 56454 379404 91898
rect 378804 56218 378986 56454
rect 379222 56218 379404 56454
rect 378804 56134 379404 56218
rect 378804 55898 378986 56134
rect 379222 55898 379404 56134
rect 378804 20454 379404 55898
rect 378804 20218 378986 20454
rect 379222 20218 379404 20454
rect 378804 20134 379404 20218
rect 378804 19898 378986 20134
rect 379222 19898 379404 20134
rect 378804 -1286 379404 19898
rect 378804 -1522 378986 -1286
rect 379222 -1522 379404 -1286
rect 378804 -1606 379404 -1522
rect 378804 -1842 378986 -1606
rect 379222 -1842 379404 -1606
rect 378804 -1864 379404 -1842
rect 382404 96054 383004 131498
rect 382404 95818 382586 96054
rect 382822 95818 383004 96054
rect 382404 95734 383004 95818
rect 382404 95498 382586 95734
rect 382822 95498 383004 95734
rect 382404 60054 383004 95498
rect 382404 59818 382586 60054
rect 382822 59818 383004 60054
rect 382404 59734 383004 59818
rect 382404 59498 382586 59734
rect 382822 59498 383004 59734
rect 382404 24054 383004 59498
rect 382404 23818 382586 24054
rect 382822 23818 383004 24054
rect 382404 23734 383004 23818
rect 382404 23498 382586 23734
rect 382822 23498 383004 23734
rect 382404 -3166 383004 23498
rect 382404 -3402 382586 -3166
rect 382822 -3402 383004 -3166
rect 382404 -3486 383004 -3402
rect 382404 -3722 382586 -3486
rect 382822 -3722 383004 -3486
rect 382404 -3744 383004 -3722
rect 386004 207654 386604 237000
rect 386004 207418 386186 207654
rect 386422 207418 386604 207654
rect 386004 207334 386604 207418
rect 386004 207098 386186 207334
rect 386422 207098 386604 207334
rect 386004 171654 386604 207098
rect 386004 171418 386186 171654
rect 386422 171418 386604 171654
rect 386004 171334 386604 171418
rect 386004 171098 386186 171334
rect 386422 171098 386604 171334
rect 386004 135654 386604 171098
rect 386004 135418 386186 135654
rect 386422 135418 386604 135654
rect 386004 135334 386604 135418
rect 386004 135098 386186 135334
rect 386422 135098 386604 135334
rect 386004 99654 386604 135098
rect 386004 99418 386186 99654
rect 386422 99418 386604 99654
rect 386004 99334 386604 99418
rect 386004 99098 386186 99334
rect 386422 99098 386604 99334
rect 386004 63654 386604 99098
rect 386004 63418 386186 63654
rect 386422 63418 386604 63654
rect 386004 63334 386604 63418
rect 386004 63098 386186 63334
rect 386422 63098 386604 63334
rect 386004 27654 386604 63098
rect 386004 27418 386186 27654
rect 386422 27418 386604 27654
rect 386004 27334 386604 27418
rect 386004 27098 386186 27334
rect 386422 27098 386604 27334
rect 386004 -5046 386604 27098
rect 386004 -5282 386186 -5046
rect 386422 -5282 386604 -5046
rect 386004 -5366 386604 -5282
rect 386004 -5602 386186 -5366
rect 386422 -5602 386604 -5366
rect 386004 -5624 386604 -5602
rect 389604 211254 390204 237000
rect 389604 211018 389786 211254
rect 390022 211018 390204 211254
rect 389604 210934 390204 211018
rect 389604 210698 389786 210934
rect 390022 210698 390204 210934
rect 389604 175254 390204 210698
rect 389604 175018 389786 175254
rect 390022 175018 390204 175254
rect 389604 174934 390204 175018
rect 389604 174698 389786 174934
rect 390022 174698 390204 174934
rect 389604 139254 390204 174698
rect 389604 139018 389786 139254
rect 390022 139018 390204 139254
rect 389604 138934 390204 139018
rect 389604 138698 389786 138934
rect 390022 138698 390204 138934
rect 389604 103254 390204 138698
rect 389604 103018 389786 103254
rect 390022 103018 390204 103254
rect 389604 102934 390204 103018
rect 389604 102698 389786 102934
rect 390022 102698 390204 102934
rect 389604 67254 390204 102698
rect 389604 67018 389786 67254
rect 390022 67018 390204 67254
rect 389604 66934 390204 67018
rect 389604 66698 389786 66934
rect 390022 66698 390204 66934
rect 389604 31254 390204 66698
rect 389604 31018 389786 31254
rect 390022 31018 390204 31254
rect 389604 30934 390204 31018
rect 389604 30698 389786 30934
rect 390022 30698 390204 30934
rect 371604 -6222 371786 -5986
rect 372022 -6222 372204 -5986
rect 371604 -6306 372204 -6222
rect 371604 -6542 371786 -6306
rect 372022 -6542 372204 -6306
rect 371604 -7504 372204 -6542
rect 389604 -6926 390204 30698
rect 396804 218454 397404 237000
rect 396804 218218 396986 218454
rect 397222 218218 397404 218454
rect 396804 218134 397404 218218
rect 396804 217898 396986 218134
rect 397222 217898 397404 218134
rect 396804 182454 397404 217898
rect 396804 182218 396986 182454
rect 397222 182218 397404 182454
rect 396804 182134 397404 182218
rect 396804 181898 396986 182134
rect 397222 181898 397404 182134
rect 396804 146454 397404 181898
rect 396804 146218 396986 146454
rect 397222 146218 397404 146454
rect 396804 146134 397404 146218
rect 396804 145898 396986 146134
rect 397222 145898 397404 146134
rect 396804 110454 397404 145898
rect 396804 110218 396986 110454
rect 397222 110218 397404 110454
rect 396804 110134 397404 110218
rect 396804 109898 396986 110134
rect 397222 109898 397404 110134
rect 396804 74454 397404 109898
rect 396804 74218 396986 74454
rect 397222 74218 397404 74454
rect 396804 74134 397404 74218
rect 396804 73898 396986 74134
rect 397222 73898 397404 74134
rect 396804 38454 397404 73898
rect 396804 38218 396986 38454
rect 397222 38218 397404 38454
rect 396804 38134 397404 38218
rect 396804 37898 396986 38134
rect 397222 37898 397404 38134
rect 396804 2454 397404 37898
rect 396804 2218 396986 2454
rect 397222 2218 397404 2454
rect 396804 2134 397404 2218
rect 396804 1898 396986 2134
rect 397222 1898 397404 2134
rect 396804 -346 397404 1898
rect 396804 -582 396986 -346
rect 397222 -582 397404 -346
rect 396804 -666 397404 -582
rect 396804 -902 396986 -666
rect 397222 -902 397404 -666
rect 396804 -1864 397404 -902
rect 400404 222054 401004 237000
rect 400404 221818 400586 222054
rect 400822 221818 401004 222054
rect 400404 221734 401004 221818
rect 400404 221498 400586 221734
rect 400822 221498 401004 221734
rect 400404 186054 401004 221498
rect 400404 185818 400586 186054
rect 400822 185818 401004 186054
rect 400404 185734 401004 185818
rect 400404 185498 400586 185734
rect 400822 185498 401004 185734
rect 400404 150054 401004 185498
rect 400404 149818 400586 150054
rect 400822 149818 401004 150054
rect 400404 149734 401004 149818
rect 400404 149498 400586 149734
rect 400822 149498 401004 149734
rect 400404 114054 401004 149498
rect 400404 113818 400586 114054
rect 400822 113818 401004 114054
rect 400404 113734 401004 113818
rect 400404 113498 400586 113734
rect 400822 113498 401004 113734
rect 400404 78054 401004 113498
rect 400404 77818 400586 78054
rect 400822 77818 401004 78054
rect 400404 77734 401004 77818
rect 400404 77498 400586 77734
rect 400822 77498 401004 77734
rect 400404 42054 401004 77498
rect 400404 41818 400586 42054
rect 400822 41818 401004 42054
rect 400404 41734 401004 41818
rect 400404 41498 400586 41734
rect 400822 41498 401004 41734
rect 400404 6054 401004 41498
rect 400404 5818 400586 6054
rect 400822 5818 401004 6054
rect 400404 5734 401004 5818
rect 400404 5498 400586 5734
rect 400822 5498 401004 5734
rect 400404 -2226 401004 5498
rect 400404 -2462 400586 -2226
rect 400822 -2462 401004 -2226
rect 400404 -2546 401004 -2462
rect 400404 -2782 400586 -2546
rect 400822 -2782 401004 -2546
rect 400404 -3744 401004 -2782
rect 404004 225654 404604 237000
rect 404004 225418 404186 225654
rect 404422 225418 404604 225654
rect 404004 225334 404604 225418
rect 404004 225098 404186 225334
rect 404422 225098 404604 225334
rect 404004 189654 404604 225098
rect 404004 189418 404186 189654
rect 404422 189418 404604 189654
rect 404004 189334 404604 189418
rect 404004 189098 404186 189334
rect 404422 189098 404604 189334
rect 404004 153654 404604 189098
rect 404004 153418 404186 153654
rect 404422 153418 404604 153654
rect 404004 153334 404604 153418
rect 404004 153098 404186 153334
rect 404422 153098 404604 153334
rect 404004 117654 404604 153098
rect 404004 117418 404186 117654
rect 404422 117418 404604 117654
rect 404004 117334 404604 117418
rect 404004 117098 404186 117334
rect 404422 117098 404604 117334
rect 404004 81654 404604 117098
rect 404004 81418 404186 81654
rect 404422 81418 404604 81654
rect 404004 81334 404604 81418
rect 404004 81098 404186 81334
rect 404422 81098 404604 81334
rect 404004 45654 404604 81098
rect 404004 45418 404186 45654
rect 404422 45418 404604 45654
rect 404004 45334 404604 45418
rect 404004 45098 404186 45334
rect 404422 45098 404604 45334
rect 404004 9654 404604 45098
rect 404004 9418 404186 9654
rect 404422 9418 404604 9654
rect 404004 9334 404604 9418
rect 404004 9098 404186 9334
rect 404422 9098 404604 9334
rect 404004 -4106 404604 9098
rect 404004 -4342 404186 -4106
rect 404422 -4342 404604 -4106
rect 404004 -4426 404604 -4342
rect 404004 -4662 404186 -4426
rect 404422 -4662 404604 -4426
rect 404004 -5624 404604 -4662
rect 407604 229254 408204 237000
rect 407604 229018 407786 229254
rect 408022 229018 408204 229254
rect 407604 228934 408204 229018
rect 407604 228698 407786 228934
rect 408022 228698 408204 228934
rect 407604 193254 408204 228698
rect 407604 193018 407786 193254
rect 408022 193018 408204 193254
rect 407604 192934 408204 193018
rect 407604 192698 407786 192934
rect 408022 192698 408204 192934
rect 407604 157254 408204 192698
rect 407604 157018 407786 157254
rect 408022 157018 408204 157254
rect 407604 156934 408204 157018
rect 407604 156698 407786 156934
rect 408022 156698 408204 156934
rect 407604 121254 408204 156698
rect 407604 121018 407786 121254
rect 408022 121018 408204 121254
rect 407604 120934 408204 121018
rect 407604 120698 407786 120934
rect 408022 120698 408204 120934
rect 407604 85254 408204 120698
rect 407604 85018 407786 85254
rect 408022 85018 408204 85254
rect 407604 84934 408204 85018
rect 407604 84698 407786 84934
rect 408022 84698 408204 84934
rect 407604 49254 408204 84698
rect 407604 49018 407786 49254
rect 408022 49018 408204 49254
rect 407604 48934 408204 49018
rect 407604 48698 407786 48934
rect 408022 48698 408204 48934
rect 407604 13254 408204 48698
rect 407604 13018 407786 13254
rect 408022 13018 408204 13254
rect 407604 12934 408204 13018
rect 407604 12698 407786 12934
rect 408022 12698 408204 12934
rect 389604 -7162 389786 -6926
rect 390022 -7162 390204 -6926
rect 389604 -7246 390204 -7162
rect 389604 -7482 389786 -7246
rect 390022 -7482 390204 -7246
rect 389604 -7504 390204 -7482
rect 407604 -5986 408204 12698
rect 414804 236454 415404 237000
rect 414804 236218 414986 236454
rect 415222 236218 415404 236454
rect 414804 236134 415404 236218
rect 414804 235898 414986 236134
rect 415222 235898 415404 236134
rect 414804 200454 415404 235898
rect 418404 204247 419004 237000
rect 422004 207654 422604 237000
rect 422004 207418 422186 207654
rect 422422 207418 422604 207654
rect 422004 207334 422604 207418
rect 422004 207098 422186 207334
rect 422422 207098 422604 207334
rect 422004 204247 422604 207098
rect 425604 211254 426204 237000
rect 425604 211018 425786 211254
rect 426022 211018 426204 211254
rect 425604 210934 426204 211018
rect 425604 210698 425786 210934
rect 426022 210698 426204 210934
rect 425604 204247 426204 210698
rect 432804 218454 433404 237000
rect 432804 218218 432986 218454
rect 433222 218218 433404 218454
rect 432804 218134 433404 218218
rect 432804 217898 432986 218134
rect 433222 217898 433404 218134
rect 432804 204247 433404 217898
rect 436404 222054 437004 237000
rect 436404 221818 436586 222054
rect 436822 221818 437004 222054
rect 436404 221734 437004 221818
rect 436404 221498 436586 221734
rect 436822 221498 437004 221734
rect 436404 204247 437004 221498
rect 440004 225654 440604 237000
rect 440004 225418 440186 225654
rect 440422 225418 440604 225654
rect 440004 225334 440604 225418
rect 440004 225098 440186 225334
rect 440422 225098 440604 225334
rect 440004 204247 440604 225098
rect 443604 229254 444204 237000
rect 443604 229018 443786 229254
rect 444022 229018 444204 229254
rect 443604 228934 444204 229018
rect 443604 228698 443786 228934
rect 444022 228698 444204 228934
rect 443604 204247 444204 228698
rect 450804 236454 451404 237000
rect 450804 236218 450986 236454
rect 451222 236218 451404 236454
rect 450804 236134 451404 236218
rect 450804 235898 450986 236134
rect 451222 235898 451404 236134
rect 450804 204247 451404 235898
rect 454404 204247 455004 237000
rect 458004 207654 458604 237000
rect 458004 207418 458186 207654
rect 458422 207418 458604 207654
rect 458004 207334 458604 207418
rect 458004 207098 458186 207334
rect 458422 207098 458604 207334
rect 458004 204247 458604 207098
rect 461604 211254 462204 237000
rect 461604 211018 461786 211254
rect 462022 211018 462204 211254
rect 461604 210934 462204 211018
rect 461604 210698 461786 210934
rect 462022 210698 462204 210934
rect 461604 204247 462204 210698
rect 468804 218454 469404 237000
rect 468804 218218 468986 218454
rect 469222 218218 469404 218454
rect 468804 218134 469404 218218
rect 468804 217898 468986 218134
rect 469222 217898 469404 218134
rect 468804 204247 469404 217898
rect 472404 222054 473004 237000
rect 472404 221818 472586 222054
rect 472822 221818 473004 222054
rect 472404 221734 473004 221818
rect 472404 221498 472586 221734
rect 472822 221498 473004 221734
rect 472404 204247 473004 221498
rect 476004 225654 476604 237000
rect 476004 225418 476186 225654
rect 476422 225418 476604 225654
rect 476004 225334 476604 225418
rect 476004 225098 476186 225334
rect 476422 225098 476604 225334
rect 474043 207772 474109 207773
rect 474043 207708 474044 207772
rect 474108 207708 474109 207772
rect 474043 207707 474109 207708
rect 456563 204236 456629 204237
rect 456563 204172 456564 204236
rect 456628 204172 456629 204236
rect 456563 204171 456629 204172
rect 468155 204236 468221 204237
rect 468155 204172 468156 204236
rect 468220 204172 468221 204236
rect 468155 204171 468221 204172
rect 470363 204236 470429 204237
rect 470363 204172 470364 204236
rect 470428 204172 470429 204236
rect 470363 204171 470429 204172
rect 449387 204100 449453 204101
rect 449387 204036 449388 204100
rect 449452 204036 449453 204100
rect 449387 204035 449453 204036
rect 448283 203828 448349 203829
rect 448283 203764 448284 203828
rect 448348 203764 448349 203828
rect 448283 203763 448349 203764
rect 448286 201650 448346 203763
rect 448262 201590 448346 201650
rect 448262 200940 448322 201590
rect 448383 201516 448449 201517
rect 448383 201452 448384 201516
rect 448448 201452 448449 201516
rect 448383 201451 448449 201452
rect 448386 200940 448446 201451
rect 449390 200970 449450 204035
rect 449571 203420 449637 203421
rect 449571 203356 449572 203420
rect 449636 203356 449637 203420
rect 449571 203355 449637 203356
rect 450859 203420 450925 203421
rect 450859 203356 450860 203420
rect 450924 203356 450925 203420
rect 450859 203355 450925 203356
rect 452147 203420 452213 203421
rect 452147 203356 452148 203420
rect 452212 203356 452213 203420
rect 452147 203355 452213 203356
rect 453251 203420 453317 203421
rect 453251 203356 453252 203420
rect 453316 203356 453317 203420
rect 453251 203355 453317 203356
rect 456011 203420 456077 203421
rect 456011 203356 456012 203420
rect 456076 203356 456077 203420
rect 456011 203355 456077 203356
rect 449390 200910 449460 200970
rect 449574 200910 449634 203355
rect 450675 203284 450741 203285
rect 450675 203220 450676 203284
rect 450740 203220 450741 203284
rect 450675 203219 450741 203220
rect 450678 201650 450738 203219
rect 450598 201590 450738 201650
rect 450598 200940 450658 201590
rect 450862 200970 450922 203355
rect 451779 203012 451845 203013
rect 451779 202948 451780 203012
rect 451844 202948 451845 203012
rect 451779 202947 451845 202948
rect 451782 201650 451842 202947
rect 450752 200910 450922 200970
rect 451766 201590 451842 201650
rect 451766 200940 451826 201590
rect 452150 200817 452210 203355
rect 452883 203284 452949 203285
rect 452883 203220 452884 203284
rect 452948 203220 452949 203284
rect 452883 203219 452949 203220
rect 452886 200970 452946 203219
rect 453254 200970 453314 203355
rect 454907 203284 454973 203285
rect 454907 203220 454908 203284
rect 454972 203220 454973 203284
rect 454907 203219 454973 203220
rect 455275 203284 455341 203285
rect 455275 203220 455276 203284
rect 455340 203220 455341 203284
rect 455275 203219 455341 203220
rect 454171 203012 454237 203013
rect 454171 202948 454172 203012
rect 454236 202948 454237 203012
rect 454171 202947 454237 202948
rect 454174 201650 454234 202947
rect 452886 200910 452964 200970
rect 453088 200910 453314 200970
rect 454102 201590 454234 201650
rect 454102 200940 454162 201590
rect 454910 200970 454970 203219
rect 455278 201650 455338 203219
rect 454256 200910 454970 200970
rect 455270 201590 455338 201650
rect 455270 200940 455330 201590
rect 456014 200970 456074 203355
rect 456379 203012 456445 203013
rect 456379 202948 456380 203012
rect 456444 202948 456445 203012
rect 456379 202947 456445 202948
rect 455424 200910 456074 200970
rect 456382 200970 456442 202947
rect 456382 200910 456468 200970
rect 456566 200910 456626 204171
rect 467051 204100 467117 204101
rect 467051 204036 467052 204100
rect 467116 204036 467117 204100
rect 467051 204035 467117 204036
rect 458771 203420 458837 203421
rect 458771 203356 458772 203420
rect 458836 203356 458837 203420
rect 458771 203355 458837 203356
rect 460979 203420 461045 203421
rect 460979 203356 460980 203420
rect 461044 203356 461045 203420
rect 460979 203355 461045 203356
rect 462267 203420 462333 203421
rect 462267 203356 462268 203420
rect 462332 203356 462333 203420
rect 462267 203355 462333 203356
rect 457483 203284 457549 203285
rect 457483 203220 457484 203284
rect 457548 203220 457549 203284
rect 457483 203219 457549 203220
rect 457486 200970 457546 203219
rect 457851 203012 457917 203013
rect 457851 202948 457852 203012
rect 457916 202948 457917 203012
rect 457851 202947 457917 202948
rect 457854 200970 457914 202947
rect 457486 200910 457636 200970
rect 457760 200910 457914 200970
rect 458774 200940 458834 203355
rect 460059 203284 460125 203285
rect 460059 203220 460060 203284
rect 460124 203220 460125 203284
rect 460059 203219 460125 203220
rect 458955 203012 459021 203013
rect 458955 202948 458956 203012
rect 459020 202948 459021 203012
rect 458955 202947 459021 202948
rect 458958 200970 459018 202947
rect 460062 201650 460122 203219
rect 460427 203012 460493 203013
rect 460427 202948 460428 203012
rect 460492 202948 460493 203012
rect 460427 202947 460493 202948
rect 458928 200910 459018 200970
rect 459942 201590 460122 201650
rect 459942 200940 460002 201590
rect 460430 200970 460490 202947
rect 460096 200910 460490 200970
rect 460982 200970 461042 203355
rect 461531 203012 461597 203013
rect 461531 202948 461532 203012
rect 461596 202948 461597 203012
rect 461531 202947 461597 202948
rect 460982 200910 461140 200970
rect 461534 200817 461594 202947
rect 462270 200910 462330 203355
rect 463187 203284 463253 203285
rect 463187 203220 463188 203284
rect 463252 203220 463253 203284
rect 463187 203219 463253 203220
rect 464659 203284 464725 203285
rect 464659 203220 464660 203284
rect 464724 203220 464725 203284
rect 464659 203219 464725 203220
rect 465947 203284 466013 203285
rect 465947 203220 465948 203284
rect 466012 203220 466013 203284
rect 465947 203219 466013 203220
rect 462451 203012 462517 203013
rect 462451 202948 462452 203012
rect 462516 202948 462517 203012
rect 462451 202947 462517 202948
rect 462454 200970 462514 202947
rect 462432 200910 462514 200970
rect 451920 200757 452210 200817
rect 461264 200757 461594 200817
rect 463190 200817 463250 203219
rect 463555 203012 463621 203013
rect 463555 202948 463556 203012
rect 463620 202948 463621 203012
rect 463555 202947 463621 202948
rect 464475 203012 464541 203013
rect 464475 202948 464476 203012
rect 464540 202948 464541 203012
rect 464475 202947 464541 202948
rect 463558 201650 463618 202947
rect 463558 201590 463630 201650
rect 463570 200940 463630 201590
rect 464478 200970 464538 202947
rect 464662 201650 464722 203219
rect 465763 203012 465829 203013
rect 465763 202948 465764 203012
rect 465828 202948 465829 203012
rect 465763 202947 465829 202948
rect 464662 201590 464798 201650
rect 464478 200910 464644 200970
rect 464738 200940 464798 201590
rect 465766 200910 465826 202947
rect 465950 200970 466010 203219
rect 467054 201650 467114 204035
rect 467235 203012 467301 203013
rect 467235 202948 467236 203012
rect 467300 202948 467301 203012
rect 467235 202947 467301 202948
rect 465936 200910 466010 200970
rect 466950 201590 467114 201650
rect 466950 200940 467010 201590
rect 467238 200970 467298 202947
rect 468158 201650 468218 204171
rect 469259 204100 469325 204101
rect 469259 204036 469260 204100
rect 469324 204036 469325 204100
rect 469259 204035 469325 204036
rect 468523 203012 468589 203013
rect 468523 202948 468524 203012
rect 468588 202948 468589 203012
rect 468523 202947 468589 202948
rect 467104 200910 467298 200970
rect 468118 201590 468218 201650
rect 468118 200940 468178 201590
rect 468526 200817 468586 202947
rect 469262 200910 469322 204035
rect 469443 203012 469509 203013
rect 469443 202948 469444 203012
rect 469508 202948 469509 203012
rect 469443 202947 469509 202948
rect 469446 200970 469506 202947
rect 470366 201650 470426 204171
rect 471651 203284 471717 203285
rect 471651 203220 471652 203284
rect 471716 203220 471717 203284
rect 471651 203219 471717 203220
rect 472755 203284 472821 203285
rect 472755 203220 472756 203284
rect 472820 203220 472821 203284
rect 472755 203219 472821 203220
rect 470731 203012 470797 203013
rect 470731 202948 470732 203012
rect 470796 202948 470797 203012
rect 470731 202947 470797 202948
rect 470366 201590 470514 201650
rect 469440 200910 469506 200970
rect 470454 200940 470514 201590
rect 470734 200970 470794 202947
rect 471654 201650 471714 203219
rect 471835 203012 471901 203013
rect 471835 202948 471836 203012
rect 471900 202948 471901 203012
rect 471835 202947 471901 202948
rect 470608 200910 470794 200970
rect 471622 201590 471714 201650
rect 471838 201650 471898 202947
rect 471838 201590 472082 201650
rect 471622 200940 471682 201590
rect 472022 200817 472082 201590
rect 472758 200970 472818 203219
rect 472939 203012 473005 203013
rect 472939 202948 472940 203012
rect 473004 202948 473005 203012
rect 472939 202947 473005 202948
rect 472758 200910 472820 200970
rect 472942 200910 473002 202947
rect 474046 201650 474106 207707
rect 476004 204247 476604 225098
rect 479604 229254 480204 237000
rect 479604 229018 479786 229254
rect 480022 229018 480204 229254
rect 479604 228934 480204 229018
rect 479604 228698 479786 228934
rect 480022 228698 480204 228934
rect 479604 204247 480204 228698
rect 486804 236454 487404 237000
rect 486804 236218 486986 236454
rect 487222 236218 487404 236454
rect 486804 236134 487404 236218
rect 486804 235898 486986 236134
rect 487222 235898 487404 236134
rect 486804 204247 487404 235898
rect 490404 204247 491004 237000
rect 494004 207654 494604 237000
rect 494004 207418 494186 207654
rect 494422 207418 494604 207654
rect 494004 207334 494604 207418
rect 494004 207098 494186 207334
rect 494422 207098 494604 207334
rect 494004 204247 494604 207098
rect 497604 211254 498204 237000
rect 497604 211018 497786 211254
rect 498022 211018 498204 211254
rect 497604 210934 498204 211018
rect 497604 210698 497786 210934
rect 498022 210698 498204 210934
rect 497604 204247 498204 210698
rect 504804 218454 505404 237000
rect 504804 218218 504986 218454
rect 505222 218218 505404 218454
rect 504804 218134 505404 218218
rect 504804 217898 504986 218134
rect 505222 217898 505404 218134
rect 477539 204236 477605 204237
rect 477539 204172 477540 204236
rect 477604 204172 477605 204236
rect 477539 204171 477605 204172
rect 479195 204236 479261 204237
rect 479195 204172 479196 204236
rect 479260 204172 479261 204236
rect 479195 204171 479261 204172
rect 481771 204236 481837 204237
rect 481771 204172 481772 204236
rect 481836 204172 481837 204236
rect 481771 204171 481837 204172
rect 490235 204236 490301 204237
rect 490235 204172 490236 204236
rect 490300 204172 490301 204236
rect 490235 204171 490301 204172
rect 476251 204100 476317 204101
rect 476251 204036 476252 204100
rect 476316 204036 476317 204100
rect 476251 204035 476317 204036
rect 475147 203284 475213 203285
rect 475147 203220 475148 203284
rect 475212 203220 475213 203284
rect 475147 203219 475213 203220
rect 474227 203012 474293 203013
rect 474227 202948 474228 203012
rect 474292 202948 474293 203012
rect 474227 202947 474293 202948
rect 473958 201590 474106 201650
rect 473958 200940 474018 201590
rect 474230 200970 474290 202947
rect 475150 201650 475210 203219
rect 475515 203012 475581 203013
rect 475515 202948 475516 203012
rect 475580 202948 475581 203012
rect 475515 202947 475581 202948
rect 474112 200910 474290 200970
rect 475126 201590 475210 201650
rect 475126 200940 475186 201590
rect 475518 200817 475578 202947
rect 476254 200970 476314 204035
rect 476435 203012 476501 203013
rect 476435 202948 476436 203012
rect 476500 202948 476501 203012
rect 476435 202947 476501 202948
rect 476254 200910 476324 200970
rect 476438 200910 476498 202947
rect 477542 201514 477602 204171
rect 478091 204100 478157 204101
rect 478091 204036 478092 204100
rect 478156 204036 478157 204100
rect 478091 204035 478157 204036
rect 477723 203284 477789 203285
rect 477723 203220 477724 203284
rect 477788 203220 477789 203284
rect 477723 203219 477789 203220
rect 477462 201454 477602 201514
rect 477462 200940 477522 201454
rect 477726 200970 477786 203219
rect 477616 200910 477786 200970
rect 478094 200970 478154 204035
rect 478643 203420 478709 203421
rect 478643 203356 478644 203420
rect 478708 203356 478709 203420
rect 478643 203355 478709 203356
rect 478646 201514 478706 203355
rect 478646 201454 478814 201514
rect 478094 200910 478660 200970
rect 478754 200940 478814 201454
rect 479198 200970 479258 204171
rect 480483 203964 480549 203965
rect 480483 203900 480484 203964
rect 480548 203900 480549 203964
rect 480483 203899 480549 203900
rect 479931 203012 479997 203013
rect 479931 202948 479932 203012
rect 479996 202948 479997 203012
rect 479931 202947 479997 202948
rect 479198 200910 479828 200970
rect 479934 200910 479994 202947
rect 480486 200970 480546 203899
rect 481219 203012 481285 203013
rect 481219 202948 481220 203012
rect 481284 202948 481285 203012
rect 481219 202947 481285 202948
rect 481222 200970 481282 202947
rect 480486 200910 480996 200970
rect 481120 200910 481282 200970
rect 481774 200970 481834 204171
rect 485819 204100 485885 204101
rect 485819 204036 485820 204100
rect 485884 204036 485885 204100
rect 485819 204035 485885 204036
rect 483059 203692 483125 203693
rect 483059 203628 483060 203692
rect 483124 203628 483125 203692
rect 483059 203627 483125 203628
rect 482139 203012 482205 203013
rect 482139 202948 482140 203012
rect 482204 202948 482205 203012
rect 482139 202947 482205 202948
rect 482142 201650 482202 202947
rect 482142 201590 482318 201650
rect 481774 200910 482164 200970
rect 482258 200940 482318 201590
rect 483062 200970 483122 203627
rect 484347 203556 484413 203557
rect 484347 203492 484348 203556
rect 484412 203492 484413 203556
rect 484347 203491 484413 203492
rect 483427 203012 483493 203013
rect 483427 202948 483428 203012
rect 483492 202948 483493 203012
rect 483427 202947 483493 202948
rect 483062 200910 483332 200970
rect 483430 200910 483490 202947
rect 484350 200970 484410 203491
rect 484715 203012 484781 203013
rect 484715 202948 484716 203012
rect 484780 202948 484781 203012
rect 484715 202947 484781 202948
rect 484718 200970 484778 202947
rect 485822 200970 485882 204035
rect 487475 203692 487541 203693
rect 487475 203628 487476 203692
rect 487540 203628 487541 203692
rect 487475 203627 487541 203628
rect 486371 203284 486437 203285
rect 486371 203220 486372 203284
rect 486436 203220 486437 203284
rect 486371 203219 486437 203220
rect 484350 200910 484500 200970
rect 484624 200910 484778 200970
rect 485792 200910 485882 200970
rect 486374 200970 486434 203219
rect 487478 200970 487538 203627
rect 488579 203556 488645 203557
rect 488579 203492 488580 203556
rect 488644 203492 488645 203556
rect 488579 203491 488645 203492
rect 488582 200970 488642 203491
rect 490238 200970 490298 204171
rect 492811 203148 492877 203149
rect 492811 203084 492812 203148
rect 492876 203084 492877 203148
rect 492811 203083 492877 203084
rect 492814 200970 492874 203083
rect 486374 200910 486960 200970
rect 487478 200910 488128 200970
rect 488582 200910 489296 200970
rect 490238 200910 490464 200970
rect 492814 200910 493463 200970
rect 463190 200757 463476 200817
rect 468272 200757 468586 200817
rect 471776 200757 472082 200817
rect 475280 200757 475578 200817
rect 414804 200218 414986 200454
rect 415222 200218 415404 200454
rect 414804 200134 415404 200218
rect 414804 199898 414986 200134
rect 415222 199898 415404 200134
rect 414804 164454 415404 199898
rect 420482 182454 420802 182476
rect 420482 182218 420524 182454
rect 420760 182218 420802 182454
rect 420482 182134 420802 182218
rect 420482 181898 420524 182134
rect 420760 181898 420802 182134
rect 420482 181876 420802 181898
rect 504804 182454 505404 217898
rect 504804 182218 504986 182454
rect 505222 182218 505404 182454
rect 504804 182134 505404 182218
rect 504804 181898 504986 182134
rect 505222 181898 505404 182134
rect 414804 164218 414986 164454
rect 415222 164218 415404 164454
rect 414804 164134 415404 164218
rect 414804 163898 414986 164134
rect 415222 163898 415404 164134
rect 414804 128454 415404 163898
rect 420034 164454 420358 164476
rect 420034 164218 420078 164454
rect 420314 164218 420358 164454
rect 420034 164134 420358 164218
rect 420034 163898 420078 164134
rect 420314 163898 420358 164134
rect 420034 163876 420358 163898
rect 420482 146454 420802 146476
rect 420482 146218 420524 146454
rect 420760 146218 420802 146454
rect 420482 146134 420802 146218
rect 420482 145898 420524 146134
rect 420760 145898 420802 146134
rect 420482 145876 420802 145898
rect 504804 146454 505404 181898
rect 504804 146218 504986 146454
rect 505222 146218 505404 146454
rect 504804 146134 505404 146218
rect 504804 145898 504986 146134
rect 505222 145898 505404 146134
rect 414804 128218 414986 128454
rect 415222 128218 415404 128454
rect 414804 128134 415404 128218
rect 414804 127898 414986 128134
rect 415222 127898 415404 128134
rect 414804 92454 415404 127898
rect 420034 128454 420358 128476
rect 420034 128218 420078 128454
rect 420314 128218 420358 128454
rect 420034 128134 420358 128218
rect 420034 127898 420078 128134
rect 420314 127898 420358 128134
rect 420034 127876 420358 127898
rect 504804 110454 505404 145898
rect 504804 110218 504986 110454
rect 505222 110218 505404 110454
rect 423693 110130 424242 110190
rect 424182 109037 424242 110130
rect 428046 110130 428688 110190
rect 504804 110134 505404 110218
rect 428046 109037 428106 110130
rect 504804 109898 504986 110134
rect 505222 109898 505404 110134
rect 424179 109036 424245 109037
rect 424179 108972 424180 109036
rect 424244 108972 424245 109036
rect 424179 108971 424245 108972
rect 428043 109036 428109 109037
rect 428043 108972 428044 109036
rect 428108 108972 428109 109036
rect 428043 108971 428109 108972
rect 414804 92218 414986 92454
rect 415222 92218 415404 92454
rect 414804 92134 415404 92218
rect 414804 91898 414986 92134
rect 415222 91898 415404 92134
rect 414804 56454 415404 91898
rect 414804 56218 414986 56454
rect 415222 56218 415404 56454
rect 414804 56134 415404 56218
rect 414804 55898 414986 56134
rect 415222 55898 415404 56134
rect 414804 20454 415404 55898
rect 414804 20218 414986 20454
rect 415222 20218 415404 20454
rect 414804 20134 415404 20218
rect 414804 19898 414986 20134
rect 415222 19898 415404 20134
rect 414804 -1286 415404 19898
rect 414804 -1522 414986 -1286
rect 415222 -1522 415404 -1286
rect 414804 -1606 415404 -1522
rect 414804 -1842 414986 -1606
rect 415222 -1842 415404 -1606
rect 414804 -1864 415404 -1842
rect 418404 96054 419004 107000
rect 418404 95818 418586 96054
rect 418822 95818 419004 96054
rect 418404 95734 419004 95818
rect 418404 95498 418586 95734
rect 418822 95498 419004 95734
rect 418404 60054 419004 95498
rect 418404 59818 418586 60054
rect 418822 59818 419004 60054
rect 418404 59734 419004 59818
rect 418404 59498 418586 59734
rect 418822 59498 419004 59734
rect 418404 24054 419004 59498
rect 418404 23818 418586 24054
rect 418822 23818 419004 24054
rect 418404 23734 419004 23818
rect 418404 23498 418586 23734
rect 418822 23498 419004 23734
rect 418404 -3166 419004 23498
rect 418404 -3402 418586 -3166
rect 418822 -3402 419004 -3166
rect 418404 -3486 419004 -3402
rect 418404 -3722 418586 -3486
rect 418822 -3722 419004 -3486
rect 418404 -3744 419004 -3722
rect 422004 99654 422604 107000
rect 422004 99418 422186 99654
rect 422422 99418 422604 99654
rect 422004 99334 422604 99418
rect 422004 99098 422186 99334
rect 422422 99098 422604 99334
rect 422004 63654 422604 99098
rect 422004 63418 422186 63654
rect 422422 63418 422604 63654
rect 422004 63334 422604 63418
rect 422004 63098 422186 63334
rect 422422 63098 422604 63334
rect 422004 27654 422604 63098
rect 422004 27418 422186 27654
rect 422422 27418 422604 27654
rect 422004 27334 422604 27418
rect 422004 27098 422186 27334
rect 422422 27098 422604 27334
rect 422004 -5046 422604 27098
rect 422004 -5282 422186 -5046
rect 422422 -5282 422604 -5046
rect 422004 -5366 422604 -5282
rect 422004 -5602 422186 -5366
rect 422422 -5602 422604 -5366
rect 422004 -5624 422604 -5602
rect 425604 103254 426204 107000
rect 425604 103018 425786 103254
rect 426022 103018 426204 103254
rect 425604 102934 426204 103018
rect 425604 102698 425786 102934
rect 426022 102698 426204 102934
rect 425604 67254 426204 102698
rect 425604 67018 425786 67254
rect 426022 67018 426204 67254
rect 425604 66934 426204 67018
rect 425604 66698 425786 66934
rect 426022 66698 426204 66934
rect 425604 31254 426204 66698
rect 425604 31018 425786 31254
rect 426022 31018 426204 31254
rect 425604 30934 426204 31018
rect 425604 30698 425786 30934
rect 426022 30698 426204 30934
rect 407604 -6222 407786 -5986
rect 408022 -6222 408204 -5986
rect 407604 -6306 408204 -6222
rect 407604 -6542 407786 -6306
rect 408022 -6542 408204 -6306
rect 407604 -7504 408204 -6542
rect 425604 -6926 426204 30698
rect 432804 74454 433404 107000
rect 432804 74218 432986 74454
rect 433222 74218 433404 74454
rect 432804 74134 433404 74218
rect 432804 73898 432986 74134
rect 433222 73898 433404 74134
rect 432804 38454 433404 73898
rect 432804 38218 432986 38454
rect 433222 38218 433404 38454
rect 432804 38134 433404 38218
rect 432804 37898 432986 38134
rect 433222 37898 433404 38134
rect 432804 2454 433404 37898
rect 432804 2218 432986 2454
rect 433222 2218 433404 2454
rect 432804 2134 433404 2218
rect 432804 1898 432986 2134
rect 433222 1898 433404 2134
rect 432804 -346 433404 1898
rect 432804 -582 432986 -346
rect 433222 -582 433404 -346
rect 432804 -666 433404 -582
rect 432804 -902 432986 -666
rect 433222 -902 433404 -666
rect 432804 -1864 433404 -902
rect 436404 78054 437004 107000
rect 436404 77818 436586 78054
rect 436822 77818 437004 78054
rect 436404 77734 437004 77818
rect 436404 77498 436586 77734
rect 436822 77498 437004 77734
rect 436404 42054 437004 77498
rect 436404 41818 436586 42054
rect 436822 41818 437004 42054
rect 436404 41734 437004 41818
rect 436404 41498 436586 41734
rect 436822 41498 437004 41734
rect 436404 6054 437004 41498
rect 436404 5818 436586 6054
rect 436822 5818 437004 6054
rect 436404 5734 437004 5818
rect 436404 5498 436586 5734
rect 436822 5498 437004 5734
rect 436404 -2226 437004 5498
rect 436404 -2462 436586 -2226
rect 436822 -2462 437004 -2226
rect 436404 -2546 437004 -2462
rect 436404 -2782 436586 -2546
rect 436822 -2782 437004 -2546
rect 436404 -3744 437004 -2782
rect 440004 81654 440604 107000
rect 440004 81418 440186 81654
rect 440422 81418 440604 81654
rect 440004 81334 440604 81418
rect 440004 81098 440186 81334
rect 440422 81098 440604 81334
rect 440004 45654 440604 81098
rect 440004 45418 440186 45654
rect 440422 45418 440604 45654
rect 440004 45334 440604 45418
rect 440004 45098 440186 45334
rect 440422 45098 440604 45334
rect 440004 9654 440604 45098
rect 440004 9418 440186 9654
rect 440422 9418 440604 9654
rect 440004 9334 440604 9418
rect 440004 9098 440186 9334
rect 440422 9098 440604 9334
rect 440004 -4106 440604 9098
rect 440004 -4342 440186 -4106
rect 440422 -4342 440604 -4106
rect 440004 -4426 440604 -4342
rect 440004 -4662 440186 -4426
rect 440422 -4662 440604 -4426
rect 440004 -5624 440604 -4662
rect 443604 85254 444204 107000
rect 443604 85018 443786 85254
rect 444022 85018 444204 85254
rect 443604 84934 444204 85018
rect 443604 84698 443786 84934
rect 444022 84698 444204 84934
rect 443604 49254 444204 84698
rect 443604 49018 443786 49254
rect 444022 49018 444204 49254
rect 443604 48934 444204 49018
rect 443604 48698 443786 48934
rect 444022 48698 444204 48934
rect 443604 13254 444204 48698
rect 443604 13018 443786 13254
rect 444022 13018 444204 13254
rect 443604 12934 444204 13018
rect 443604 12698 443786 12934
rect 444022 12698 444204 12934
rect 425604 -7162 425786 -6926
rect 426022 -7162 426204 -6926
rect 425604 -7246 426204 -7162
rect 425604 -7482 425786 -7246
rect 426022 -7482 426204 -7246
rect 425604 -7504 426204 -7482
rect 443604 -5986 444204 12698
rect 450804 92454 451404 107000
rect 450804 92218 450986 92454
rect 451222 92218 451404 92454
rect 450804 92134 451404 92218
rect 450804 91898 450986 92134
rect 451222 91898 451404 92134
rect 450804 56454 451404 91898
rect 450804 56218 450986 56454
rect 451222 56218 451404 56454
rect 450804 56134 451404 56218
rect 450804 55898 450986 56134
rect 451222 55898 451404 56134
rect 450804 20454 451404 55898
rect 450804 20218 450986 20454
rect 451222 20218 451404 20454
rect 450804 20134 451404 20218
rect 450804 19898 450986 20134
rect 451222 19898 451404 20134
rect 450804 -1286 451404 19898
rect 450804 -1522 450986 -1286
rect 451222 -1522 451404 -1286
rect 450804 -1606 451404 -1522
rect 450804 -1842 450986 -1606
rect 451222 -1842 451404 -1606
rect 450804 -1864 451404 -1842
rect 454404 96054 455004 107000
rect 454404 95818 454586 96054
rect 454822 95818 455004 96054
rect 454404 95734 455004 95818
rect 454404 95498 454586 95734
rect 454822 95498 455004 95734
rect 454404 60054 455004 95498
rect 454404 59818 454586 60054
rect 454822 59818 455004 60054
rect 454404 59734 455004 59818
rect 454404 59498 454586 59734
rect 454822 59498 455004 59734
rect 454404 24054 455004 59498
rect 454404 23818 454586 24054
rect 454822 23818 455004 24054
rect 454404 23734 455004 23818
rect 454404 23498 454586 23734
rect 454822 23498 455004 23734
rect 454404 -3166 455004 23498
rect 454404 -3402 454586 -3166
rect 454822 -3402 455004 -3166
rect 454404 -3486 455004 -3402
rect 454404 -3722 454586 -3486
rect 454822 -3722 455004 -3486
rect 454404 -3744 455004 -3722
rect 458004 99654 458604 107000
rect 458004 99418 458186 99654
rect 458422 99418 458604 99654
rect 458004 99334 458604 99418
rect 458004 99098 458186 99334
rect 458422 99098 458604 99334
rect 458004 63654 458604 99098
rect 458004 63418 458186 63654
rect 458422 63418 458604 63654
rect 458004 63334 458604 63418
rect 458004 63098 458186 63334
rect 458422 63098 458604 63334
rect 458004 27654 458604 63098
rect 458004 27418 458186 27654
rect 458422 27418 458604 27654
rect 458004 27334 458604 27418
rect 458004 27098 458186 27334
rect 458422 27098 458604 27334
rect 458004 -5046 458604 27098
rect 458004 -5282 458186 -5046
rect 458422 -5282 458604 -5046
rect 458004 -5366 458604 -5282
rect 458004 -5602 458186 -5366
rect 458422 -5602 458604 -5366
rect 458004 -5624 458604 -5602
rect 461604 103254 462204 107000
rect 461604 103018 461786 103254
rect 462022 103018 462204 103254
rect 461604 102934 462204 103018
rect 461604 102698 461786 102934
rect 462022 102698 462204 102934
rect 461604 67254 462204 102698
rect 461604 67018 461786 67254
rect 462022 67018 462204 67254
rect 461604 66934 462204 67018
rect 461604 66698 461786 66934
rect 462022 66698 462204 66934
rect 461604 31254 462204 66698
rect 461604 31018 461786 31254
rect 462022 31018 462204 31254
rect 461604 30934 462204 31018
rect 461604 30698 461786 30934
rect 462022 30698 462204 30934
rect 443604 -6222 443786 -5986
rect 444022 -6222 444204 -5986
rect 443604 -6306 444204 -6222
rect 443604 -6542 443786 -6306
rect 444022 -6542 444204 -6306
rect 443604 -7504 444204 -6542
rect 461604 -6926 462204 30698
rect 468804 74454 469404 107000
rect 468804 74218 468986 74454
rect 469222 74218 469404 74454
rect 468804 74134 469404 74218
rect 468804 73898 468986 74134
rect 469222 73898 469404 74134
rect 468804 38454 469404 73898
rect 468804 38218 468986 38454
rect 469222 38218 469404 38454
rect 468804 38134 469404 38218
rect 468804 37898 468986 38134
rect 469222 37898 469404 38134
rect 468804 2454 469404 37898
rect 468804 2218 468986 2454
rect 469222 2218 469404 2454
rect 468804 2134 469404 2218
rect 468804 1898 468986 2134
rect 469222 1898 469404 2134
rect 468804 -346 469404 1898
rect 468804 -582 468986 -346
rect 469222 -582 469404 -346
rect 468804 -666 469404 -582
rect 468804 -902 468986 -666
rect 469222 -902 469404 -666
rect 468804 -1864 469404 -902
rect 472404 78054 473004 107000
rect 472404 77818 472586 78054
rect 472822 77818 473004 78054
rect 472404 77734 473004 77818
rect 472404 77498 472586 77734
rect 472822 77498 473004 77734
rect 472404 42054 473004 77498
rect 472404 41818 472586 42054
rect 472822 41818 473004 42054
rect 472404 41734 473004 41818
rect 472404 41498 472586 41734
rect 472822 41498 473004 41734
rect 472404 6054 473004 41498
rect 472404 5818 472586 6054
rect 472822 5818 473004 6054
rect 472404 5734 473004 5818
rect 472404 5498 472586 5734
rect 472822 5498 473004 5734
rect 472404 -2226 473004 5498
rect 472404 -2462 472586 -2226
rect 472822 -2462 473004 -2226
rect 472404 -2546 473004 -2462
rect 472404 -2782 472586 -2546
rect 472822 -2782 473004 -2546
rect 472404 -3744 473004 -2782
rect 476004 81654 476604 107000
rect 476004 81418 476186 81654
rect 476422 81418 476604 81654
rect 476004 81334 476604 81418
rect 476004 81098 476186 81334
rect 476422 81098 476604 81334
rect 476004 45654 476604 81098
rect 476004 45418 476186 45654
rect 476422 45418 476604 45654
rect 476004 45334 476604 45418
rect 476004 45098 476186 45334
rect 476422 45098 476604 45334
rect 476004 9654 476604 45098
rect 476004 9418 476186 9654
rect 476422 9418 476604 9654
rect 476004 9334 476604 9418
rect 476004 9098 476186 9334
rect 476422 9098 476604 9334
rect 476004 -4106 476604 9098
rect 476004 -4342 476186 -4106
rect 476422 -4342 476604 -4106
rect 476004 -4426 476604 -4342
rect 476004 -4662 476186 -4426
rect 476422 -4662 476604 -4426
rect 476004 -5624 476604 -4662
rect 479604 85254 480204 107000
rect 479604 85018 479786 85254
rect 480022 85018 480204 85254
rect 479604 84934 480204 85018
rect 479604 84698 479786 84934
rect 480022 84698 480204 84934
rect 479604 49254 480204 84698
rect 479604 49018 479786 49254
rect 480022 49018 480204 49254
rect 479604 48934 480204 49018
rect 479604 48698 479786 48934
rect 480022 48698 480204 48934
rect 479604 13254 480204 48698
rect 479604 13018 479786 13254
rect 480022 13018 480204 13254
rect 479604 12934 480204 13018
rect 479604 12698 479786 12934
rect 480022 12698 480204 12934
rect 461604 -7162 461786 -6926
rect 462022 -7162 462204 -6926
rect 461604 -7246 462204 -7162
rect 461604 -7482 461786 -7246
rect 462022 -7482 462204 -7246
rect 461604 -7504 462204 -7482
rect 479604 -5986 480204 12698
rect 486804 92454 487404 107000
rect 486804 92218 486986 92454
rect 487222 92218 487404 92454
rect 486804 92134 487404 92218
rect 486804 91898 486986 92134
rect 487222 91898 487404 92134
rect 486804 56454 487404 91898
rect 486804 56218 486986 56454
rect 487222 56218 487404 56454
rect 486804 56134 487404 56218
rect 486804 55898 486986 56134
rect 487222 55898 487404 56134
rect 486804 20454 487404 55898
rect 486804 20218 486986 20454
rect 487222 20218 487404 20454
rect 486804 20134 487404 20218
rect 486804 19898 486986 20134
rect 487222 19898 487404 20134
rect 486804 -1286 487404 19898
rect 486804 -1522 486986 -1286
rect 487222 -1522 487404 -1286
rect 486804 -1606 487404 -1522
rect 486804 -1842 486986 -1606
rect 487222 -1842 487404 -1606
rect 486804 -1864 487404 -1842
rect 490404 96054 491004 107000
rect 490404 95818 490586 96054
rect 490822 95818 491004 96054
rect 490404 95734 491004 95818
rect 490404 95498 490586 95734
rect 490822 95498 491004 95734
rect 490404 60054 491004 95498
rect 490404 59818 490586 60054
rect 490822 59818 491004 60054
rect 490404 59734 491004 59818
rect 490404 59498 490586 59734
rect 490822 59498 491004 59734
rect 490404 24054 491004 59498
rect 490404 23818 490586 24054
rect 490822 23818 491004 24054
rect 490404 23734 491004 23818
rect 490404 23498 490586 23734
rect 490822 23498 491004 23734
rect 490404 -3166 491004 23498
rect 490404 -3402 490586 -3166
rect 490822 -3402 491004 -3166
rect 490404 -3486 491004 -3402
rect 490404 -3722 490586 -3486
rect 490822 -3722 491004 -3486
rect 490404 -3744 491004 -3722
rect 494004 99654 494604 107000
rect 494004 99418 494186 99654
rect 494422 99418 494604 99654
rect 494004 99334 494604 99418
rect 494004 99098 494186 99334
rect 494422 99098 494604 99334
rect 494004 63654 494604 99098
rect 494004 63418 494186 63654
rect 494422 63418 494604 63654
rect 494004 63334 494604 63418
rect 494004 63098 494186 63334
rect 494422 63098 494604 63334
rect 494004 27654 494604 63098
rect 494004 27418 494186 27654
rect 494422 27418 494604 27654
rect 494004 27334 494604 27418
rect 494004 27098 494186 27334
rect 494422 27098 494604 27334
rect 494004 -5046 494604 27098
rect 494004 -5282 494186 -5046
rect 494422 -5282 494604 -5046
rect 494004 -5366 494604 -5282
rect 494004 -5602 494186 -5366
rect 494422 -5602 494604 -5366
rect 494004 -5624 494604 -5602
rect 497604 103254 498204 107000
rect 497604 103018 497786 103254
rect 498022 103018 498204 103254
rect 497604 102934 498204 103018
rect 497604 102698 497786 102934
rect 498022 102698 498204 102934
rect 497604 67254 498204 102698
rect 497604 67018 497786 67254
rect 498022 67018 498204 67254
rect 497604 66934 498204 67018
rect 497604 66698 497786 66934
rect 498022 66698 498204 66934
rect 497604 31254 498204 66698
rect 497604 31018 497786 31254
rect 498022 31018 498204 31254
rect 497604 30934 498204 31018
rect 497604 30698 497786 30934
rect 498022 30698 498204 30934
rect 479604 -6222 479786 -5986
rect 480022 -6222 480204 -5986
rect 479604 -6306 480204 -6222
rect 479604 -6542 479786 -6306
rect 480022 -6542 480204 -6306
rect 479604 -7504 480204 -6542
rect 497604 -6926 498204 30698
rect 504804 74454 505404 109898
rect 504804 74218 504986 74454
rect 505222 74218 505404 74454
rect 504804 74134 505404 74218
rect 504804 73898 504986 74134
rect 505222 73898 505404 74134
rect 504804 38454 505404 73898
rect 504804 38218 504986 38454
rect 505222 38218 505404 38454
rect 504804 38134 505404 38218
rect 504804 37898 504986 38134
rect 505222 37898 505404 38134
rect 504804 2454 505404 37898
rect 504804 2218 504986 2454
rect 505222 2218 505404 2454
rect 504804 2134 505404 2218
rect 504804 1898 504986 2134
rect 505222 1898 505404 2134
rect 504804 -346 505404 1898
rect 504804 -582 504986 -346
rect 505222 -582 505404 -346
rect 504804 -666 505404 -582
rect 504804 -902 504986 -666
rect 505222 -902 505404 -666
rect 504804 -1864 505404 -902
rect 508404 222054 509004 237000
rect 508404 221818 508586 222054
rect 508822 221818 509004 222054
rect 508404 221734 509004 221818
rect 508404 221498 508586 221734
rect 508822 221498 509004 221734
rect 508404 186054 509004 221498
rect 508404 185818 508586 186054
rect 508822 185818 509004 186054
rect 508404 185734 509004 185818
rect 508404 185498 508586 185734
rect 508822 185498 509004 185734
rect 508404 150054 509004 185498
rect 508404 149818 508586 150054
rect 508822 149818 509004 150054
rect 508404 149734 509004 149818
rect 508404 149498 508586 149734
rect 508822 149498 509004 149734
rect 508404 114054 509004 149498
rect 508404 113818 508586 114054
rect 508822 113818 509004 114054
rect 508404 113734 509004 113818
rect 508404 113498 508586 113734
rect 508822 113498 509004 113734
rect 508404 78054 509004 113498
rect 508404 77818 508586 78054
rect 508822 77818 509004 78054
rect 508404 77734 509004 77818
rect 508404 77498 508586 77734
rect 508822 77498 509004 77734
rect 508404 42054 509004 77498
rect 508404 41818 508586 42054
rect 508822 41818 509004 42054
rect 508404 41734 509004 41818
rect 508404 41498 508586 41734
rect 508822 41498 509004 41734
rect 508404 6054 509004 41498
rect 508404 5818 508586 6054
rect 508822 5818 509004 6054
rect 508404 5734 509004 5818
rect 508404 5498 508586 5734
rect 508822 5498 509004 5734
rect 508404 -2226 509004 5498
rect 508404 -2462 508586 -2226
rect 508822 -2462 509004 -2226
rect 508404 -2546 509004 -2462
rect 508404 -2782 508586 -2546
rect 508822 -2782 509004 -2546
rect 508404 -3744 509004 -2782
rect 512004 225654 512604 237000
rect 512004 225418 512186 225654
rect 512422 225418 512604 225654
rect 512004 225334 512604 225418
rect 512004 225098 512186 225334
rect 512422 225098 512604 225334
rect 512004 189654 512604 225098
rect 512004 189418 512186 189654
rect 512422 189418 512604 189654
rect 512004 189334 512604 189418
rect 512004 189098 512186 189334
rect 512422 189098 512604 189334
rect 512004 153654 512604 189098
rect 512004 153418 512186 153654
rect 512422 153418 512604 153654
rect 512004 153334 512604 153418
rect 512004 153098 512186 153334
rect 512422 153098 512604 153334
rect 512004 117654 512604 153098
rect 512004 117418 512186 117654
rect 512422 117418 512604 117654
rect 512004 117334 512604 117418
rect 512004 117098 512186 117334
rect 512422 117098 512604 117334
rect 512004 81654 512604 117098
rect 512004 81418 512186 81654
rect 512422 81418 512604 81654
rect 512004 81334 512604 81418
rect 512004 81098 512186 81334
rect 512422 81098 512604 81334
rect 512004 45654 512604 81098
rect 512004 45418 512186 45654
rect 512422 45418 512604 45654
rect 512004 45334 512604 45418
rect 512004 45098 512186 45334
rect 512422 45098 512604 45334
rect 512004 9654 512604 45098
rect 512004 9418 512186 9654
rect 512422 9418 512604 9654
rect 512004 9334 512604 9418
rect 512004 9098 512186 9334
rect 512422 9098 512604 9334
rect 512004 -4106 512604 9098
rect 512004 -4342 512186 -4106
rect 512422 -4342 512604 -4106
rect 512004 -4426 512604 -4342
rect 512004 -4662 512186 -4426
rect 512422 -4662 512604 -4426
rect 512004 -5624 512604 -4662
rect 515604 229254 516204 237000
rect 515604 229018 515786 229254
rect 516022 229018 516204 229254
rect 515604 228934 516204 229018
rect 515604 228698 515786 228934
rect 516022 228698 516204 228934
rect 515604 193254 516204 228698
rect 515604 193018 515786 193254
rect 516022 193018 516204 193254
rect 515604 192934 516204 193018
rect 515604 192698 515786 192934
rect 516022 192698 516204 192934
rect 515604 157254 516204 192698
rect 515604 157018 515786 157254
rect 516022 157018 516204 157254
rect 515604 156934 516204 157018
rect 515604 156698 515786 156934
rect 516022 156698 516204 156934
rect 515604 121254 516204 156698
rect 515604 121018 515786 121254
rect 516022 121018 516204 121254
rect 515604 120934 516204 121018
rect 515604 120698 515786 120934
rect 516022 120698 516204 120934
rect 515604 85254 516204 120698
rect 515604 85018 515786 85254
rect 516022 85018 516204 85254
rect 515604 84934 516204 85018
rect 515604 84698 515786 84934
rect 516022 84698 516204 84934
rect 515604 49254 516204 84698
rect 515604 49018 515786 49254
rect 516022 49018 516204 49254
rect 515604 48934 516204 49018
rect 515604 48698 515786 48934
rect 516022 48698 516204 48934
rect 515604 13254 516204 48698
rect 515604 13018 515786 13254
rect 516022 13018 516204 13254
rect 515604 12934 516204 13018
rect 515604 12698 515786 12934
rect 516022 12698 516204 12934
rect 497604 -7162 497786 -6926
rect 498022 -7162 498204 -6926
rect 497604 -7246 498204 -7162
rect 497604 -7482 497786 -7246
rect 498022 -7482 498204 -7246
rect 497604 -7504 498204 -7482
rect 515604 -5986 516204 12698
rect 522804 236454 523404 237000
rect 522804 236218 522986 236454
rect 523222 236218 523404 236454
rect 522804 236134 523404 236218
rect 522804 235898 522986 236134
rect 523222 235898 523404 236134
rect 522804 200454 523404 235898
rect 522804 200218 522986 200454
rect 523222 200218 523404 200454
rect 522804 200134 523404 200218
rect 522804 199898 522986 200134
rect 523222 199898 523404 200134
rect 522804 164454 523404 199898
rect 522804 164218 522986 164454
rect 523222 164218 523404 164454
rect 522804 164134 523404 164218
rect 522804 163898 522986 164134
rect 523222 163898 523404 164134
rect 522804 128454 523404 163898
rect 522804 128218 522986 128454
rect 523222 128218 523404 128454
rect 522804 128134 523404 128218
rect 522804 127898 522986 128134
rect 523222 127898 523404 128134
rect 522804 92454 523404 127898
rect 522804 92218 522986 92454
rect 523222 92218 523404 92454
rect 522804 92134 523404 92218
rect 522804 91898 522986 92134
rect 523222 91898 523404 92134
rect 522804 56454 523404 91898
rect 522804 56218 522986 56454
rect 523222 56218 523404 56454
rect 522804 56134 523404 56218
rect 522804 55898 522986 56134
rect 523222 55898 523404 56134
rect 522804 20454 523404 55898
rect 522804 20218 522986 20454
rect 523222 20218 523404 20454
rect 522804 20134 523404 20218
rect 522804 19898 522986 20134
rect 523222 19898 523404 20134
rect 522804 -1286 523404 19898
rect 522804 -1522 522986 -1286
rect 523222 -1522 523404 -1286
rect 522804 -1606 523404 -1522
rect 522804 -1842 522986 -1606
rect 523222 -1842 523404 -1606
rect 522804 -1864 523404 -1842
rect 526404 204054 527004 237000
rect 526404 203818 526586 204054
rect 526822 203818 527004 204054
rect 526404 203734 527004 203818
rect 526404 203498 526586 203734
rect 526822 203498 527004 203734
rect 526404 168054 527004 203498
rect 526404 167818 526586 168054
rect 526822 167818 527004 168054
rect 526404 167734 527004 167818
rect 526404 167498 526586 167734
rect 526822 167498 527004 167734
rect 526404 132054 527004 167498
rect 526404 131818 526586 132054
rect 526822 131818 527004 132054
rect 526404 131734 527004 131818
rect 526404 131498 526586 131734
rect 526822 131498 527004 131734
rect 526404 96054 527004 131498
rect 526404 95818 526586 96054
rect 526822 95818 527004 96054
rect 526404 95734 527004 95818
rect 526404 95498 526586 95734
rect 526822 95498 527004 95734
rect 526404 60054 527004 95498
rect 526404 59818 526586 60054
rect 526822 59818 527004 60054
rect 526404 59734 527004 59818
rect 526404 59498 526586 59734
rect 526822 59498 527004 59734
rect 526404 24054 527004 59498
rect 526404 23818 526586 24054
rect 526822 23818 527004 24054
rect 526404 23734 527004 23818
rect 526404 23498 526586 23734
rect 526822 23498 527004 23734
rect 526404 -3166 527004 23498
rect 526404 -3402 526586 -3166
rect 526822 -3402 527004 -3166
rect 526404 -3486 527004 -3402
rect 526404 -3722 526586 -3486
rect 526822 -3722 527004 -3486
rect 526404 -3744 527004 -3722
rect 530004 207654 530604 237000
rect 530004 207418 530186 207654
rect 530422 207418 530604 207654
rect 530004 207334 530604 207418
rect 530004 207098 530186 207334
rect 530422 207098 530604 207334
rect 530004 171654 530604 207098
rect 530004 171418 530186 171654
rect 530422 171418 530604 171654
rect 530004 171334 530604 171418
rect 530004 171098 530186 171334
rect 530422 171098 530604 171334
rect 530004 135654 530604 171098
rect 530004 135418 530186 135654
rect 530422 135418 530604 135654
rect 530004 135334 530604 135418
rect 530004 135098 530186 135334
rect 530422 135098 530604 135334
rect 530004 99654 530604 135098
rect 530004 99418 530186 99654
rect 530422 99418 530604 99654
rect 530004 99334 530604 99418
rect 530004 99098 530186 99334
rect 530422 99098 530604 99334
rect 530004 63654 530604 99098
rect 530004 63418 530186 63654
rect 530422 63418 530604 63654
rect 530004 63334 530604 63418
rect 530004 63098 530186 63334
rect 530422 63098 530604 63334
rect 530004 27654 530604 63098
rect 530004 27418 530186 27654
rect 530422 27418 530604 27654
rect 530004 27334 530604 27418
rect 530004 27098 530186 27334
rect 530422 27098 530604 27334
rect 530004 -5046 530604 27098
rect 530004 -5282 530186 -5046
rect 530422 -5282 530604 -5046
rect 530004 -5366 530604 -5282
rect 530004 -5602 530186 -5366
rect 530422 -5602 530604 -5366
rect 530004 -5624 530604 -5602
rect 533604 211254 534204 237000
rect 538446 227765 538506 242390
rect 538998 240821 539058 250550
rect 538995 240820 539061 240821
rect 538995 240756 538996 240820
rect 539060 240756 539061 240820
rect 538995 240755 539061 240756
rect 538443 227764 538509 227765
rect 538443 227700 538444 227764
rect 538508 227700 538509 227764
rect 538443 227699 538509 227700
rect 538627 227764 538693 227765
rect 538627 227700 538628 227764
rect 538692 227700 538693 227764
rect 538627 227699 538693 227700
rect 538630 222869 538690 227699
rect 538627 222868 538693 222869
rect 538627 222804 538628 222868
rect 538692 222804 538693 222868
rect 538627 222803 538693 222804
rect 533604 211018 533786 211254
rect 534022 211018 534204 211254
rect 533604 210934 534204 211018
rect 533604 210698 533786 210934
rect 534022 210698 534204 210934
rect 533604 175254 534204 210698
rect 538259 205460 538325 205461
rect 538259 205396 538260 205460
rect 538324 205396 538325 205460
rect 538259 205395 538325 205396
rect 538262 201109 538322 205395
rect 538259 201108 538325 201109
rect 538259 201044 538260 201108
rect 538324 201044 538325 201108
rect 538259 201043 538325 201044
rect 533604 175018 533786 175254
rect 534022 175018 534204 175254
rect 533604 174934 534204 175018
rect 533604 174698 533786 174934
rect 534022 174698 534204 174934
rect 533604 139254 534204 174698
rect 533604 139018 533786 139254
rect 534022 139018 534204 139254
rect 533604 138934 534204 139018
rect 533604 138698 533786 138934
rect 534022 138698 534204 138934
rect 533604 103254 534204 138698
rect 533604 103018 533786 103254
rect 534022 103018 534204 103254
rect 533604 102934 534204 103018
rect 533604 102698 533786 102934
rect 534022 102698 534204 102934
rect 533604 67254 534204 102698
rect 533604 67018 533786 67254
rect 534022 67018 534204 67254
rect 533604 66934 534204 67018
rect 533604 66698 533786 66934
rect 534022 66698 534204 66934
rect 533604 31254 534204 66698
rect 539550 50965 539610 359347
rect 539734 349077 539794 363430
rect 539731 349076 539797 349077
rect 539731 349012 539732 349076
rect 539796 349012 539797 349076
rect 539731 349011 539797 349012
rect 539915 331260 539981 331261
rect 539915 331196 539916 331260
rect 539980 331196 539981 331260
rect 539915 331195 539981 331196
rect 539918 320650 539978 331195
rect 539918 320590 540162 320650
rect 540102 314530 540162 320590
rect 539918 314470 540162 314530
rect 539918 302429 539978 314470
rect 539915 302428 539981 302429
rect 539915 302364 539916 302428
rect 539980 302364 539981 302428
rect 539915 302363 539981 302364
rect 540099 302156 540165 302157
rect 540099 302092 540100 302156
rect 540164 302092 540165 302156
rect 540099 302091 540165 302092
rect 540102 291957 540162 302091
rect 540099 291956 540165 291957
rect 540099 291892 540100 291956
rect 540164 291892 540165 291956
rect 540099 291891 540165 291892
rect 540099 279172 540165 279173
rect 540099 279108 540100 279172
rect 540164 279108 540165 279172
rect 540099 279107 540165 279108
rect 540102 273461 540162 279107
rect 540099 273460 540165 273461
rect 540099 273396 540100 273460
rect 540164 273396 540165 273460
rect 540099 273395 540165 273396
rect 539731 265028 539797 265029
rect 539731 264964 539732 265028
rect 539796 264964 539797 265028
rect 539731 264963 539797 264964
rect 539734 263669 539794 264963
rect 539731 263668 539797 263669
rect 539731 263604 539732 263668
rect 539796 263604 539797 263668
rect 539731 263603 539797 263604
rect 539915 263532 539981 263533
rect 539915 263468 539916 263532
rect 539980 263468 539981 263532
rect 539915 263467 539981 263468
rect 539918 256730 539978 263467
rect 539918 256670 540162 256730
rect 540102 216069 540162 256670
rect 540099 216068 540165 216069
rect 540099 216004 540100 216068
rect 540164 216004 540165 216068
rect 540099 216003 540165 216004
rect 539915 203012 539981 203013
rect 539915 202948 539916 203012
rect 539980 202948 539981 203012
rect 539915 202947 539981 202948
rect 539918 196077 539978 202947
rect 540286 200973 540346 462027
rect 540467 452028 540533 452029
rect 540467 451964 540468 452028
rect 540532 451964 540533 452028
rect 540467 451963 540533 451964
rect 540470 442373 540530 451963
rect 540467 442372 540533 442373
rect 540467 442308 540468 442372
rect 540532 442308 540533 442372
rect 540467 442307 540533 442308
rect 540467 432716 540533 432717
rect 540467 432652 540468 432716
rect 540532 432652 540533 432716
rect 540467 432651 540533 432652
rect 540470 413405 540530 432651
rect 540467 413404 540533 413405
rect 540467 413340 540468 413404
rect 540532 413340 540533 413404
rect 540467 413339 540533 413340
rect 540467 403748 540533 403749
rect 540467 403684 540468 403748
rect 540532 403684 540533 403748
rect 540467 403683 540533 403684
rect 540470 381037 540530 403683
rect 540467 381036 540533 381037
rect 540467 380972 540468 381036
rect 540532 380972 540533 381036
rect 540467 380971 540533 380972
rect 540804 218454 541404 237000
rect 540804 218218 540986 218454
rect 541222 218218 541404 218454
rect 540804 218134 541404 218218
rect 540804 217898 540986 218134
rect 541222 217898 541404 218134
rect 540283 200972 540349 200973
rect 540283 200908 540284 200972
rect 540348 200908 540349 200972
rect 540283 200907 540349 200908
rect 539915 196076 539981 196077
rect 539915 196012 539916 196076
rect 539980 196012 539981 196076
rect 539915 196011 539981 196012
rect 540099 195804 540165 195805
rect 540099 195740 540100 195804
rect 540164 195740 540165 195804
rect 540099 195739 540165 195740
rect 540102 193221 540162 195739
rect 540099 193220 540165 193221
rect 540099 193156 540100 193220
rect 540164 193156 540165 193220
rect 540099 193155 540165 193156
rect 539915 183700 539981 183701
rect 539915 183636 539916 183700
rect 539980 183636 539981 183700
rect 539915 183635 539981 183636
rect 539918 176765 539978 183635
rect 540804 182454 541404 217898
rect 540804 182218 540986 182454
rect 541222 182218 541404 182454
rect 540804 182134 541404 182218
rect 540804 181898 540986 182134
rect 541222 181898 541404 182134
rect 539915 176764 539981 176765
rect 539915 176700 539916 176764
rect 539980 176700 539981 176764
rect 539915 176699 539981 176700
rect 540099 176492 540165 176493
rect 540099 176428 540100 176492
rect 540164 176428 540165 176492
rect 540099 176427 540165 176428
rect 540102 167109 540162 176427
rect 540099 167108 540165 167109
rect 540099 167044 540100 167108
rect 540164 167044 540165 167108
rect 540099 167043 540165 167044
rect 540099 164252 540165 164253
rect 540099 164250 540100 164252
rect 539918 164190 540100 164250
rect 539918 162757 539978 164190
rect 540099 164188 540100 164190
rect 540164 164188 540165 164252
rect 540099 164187 540165 164188
rect 539915 162756 539981 162757
rect 539915 162692 539916 162756
rect 539980 162692 539981 162756
rect 539915 162691 539981 162692
rect 540099 153236 540165 153237
rect 540099 153172 540100 153236
rect 540164 153172 540165 153236
rect 540099 153171 540165 153172
rect 540102 147797 540162 153171
rect 540099 147796 540165 147797
rect 540099 147732 540100 147796
rect 540164 147732 540165 147796
rect 540099 147731 540165 147732
rect 540804 146454 541404 181898
rect 540804 146218 540986 146454
rect 541222 146218 541404 146454
rect 540804 146134 541404 146218
rect 540804 145898 540986 146134
rect 541222 145898 541404 146134
rect 539731 144940 539797 144941
rect 539731 144876 539732 144940
rect 539796 144876 539797 144940
rect 539731 144875 539797 144876
rect 539734 137730 539794 144875
rect 539734 137670 540162 137730
rect 540102 128210 540162 137670
rect 539918 128150 540162 128210
rect 539918 120733 539978 128150
rect 539915 120732 539981 120733
rect 539915 120668 539916 120732
rect 539980 120668 539981 120732
rect 539915 120667 539981 120668
rect 540099 115972 540165 115973
rect 540099 115908 540100 115972
rect 540164 115908 540165 115972
rect 540099 115907 540165 115908
rect 540102 93533 540162 115907
rect 540804 110454 541404 145898
rect 540804 110218 540986 110454
rect 541222 110218 541404 110454
rect 540804 110134 541404 110218
rect 540804 109898 540986 110134
rect 541222 109898 541404 110134
rect 540099 93532 540165 93533
rect 540099 93468 540100 93532
rect 540164 93468 540165 93532
rect 540099 93467 540165 93468
rect 540804 74454 541404 109898
rect 540804 74218 540986 74454
rect 541222 74218 541404 74454
rect 540804 74134 541404 74218
rect 540804 73898 540986 74134
rect 541222 73898 541404 74134
rect 539547 50964 539613 50965
rect 539547 50900 539548 50964
rect 539612 50900 539613 50964
rect 539547 50899 539613 50900
rect 533604 31018 533786 31254
rect 534022 31018 534204 31254
rect 533604 30934 534204 31018
rect 533604 30698 533786 30934
rect 534022 30698 534204 30934
rect 515604 -6222 515786 -5986
rect 516022 -6222 516204 -5986
rect 515604 -6306 516204 -6222
rect 515604 -6542 515786 -6306
rect 516022 -6542 516204 -6306
rect 515604 -7504 516204 -6542
rect 533604 -6926 534204 30698
rect 540804 38454 541404 73898
rect 541574 64837 541634 472635
rect 541571 64836 541637 64837
rect 541571 64772 541572 64836
rect 541636 64772 541637 64836
rect 541571 64771 541637 64772
rect 540804 38218 540986 38454
rect 541222 38218 541404 38454
rect 540804 38134 541404 38218
rect 540804 37898 540986 38134
rect 541222 37898 541404 38134
rect 540804 2454 541404 37898
rect 542310 8261 542370 476851
rect 542494 21997 542554 478891
rect 542675 474740 542741 474741
rect 542675 474676 542676 474740
rect 542740 474676 542741 474740
rect 542675 474675 542741 474676
rect 542678 35869 542738 474675
rect 544404 474054 545004 509498
rect 544404 473818 544586 474054
rect 544822 473818 545004 474054
rect 544404 473734 545004 473818
rect 544404 473498 544586 473734
rect 544822 473498 545004 473734
rect 542859 468484 542925 468485
rect 542859 468420 542860 468484
rect 542924 468420 542925 468484
rect 542859 468419 542925 468420
rect 542862 80069 542922 468419
rect 543043 460052 543109 460053
rect 543043 459988 543044 460052
rect 543108 459988 543109 460052
rect 543043 459987 543109 459988
rect 543046 200837 543106 459987
rect 543227 457876 543293 457877
rect 543227 457812 543228 457876
rect 543292 457812 543293 457876
rect 543227 457811 543293 457812
rect 543043 200836 543109 200837
rect 543043 200772 543044 200836
rect 543108 200772 543109 200836
rect 543043 200771 543109 200772
rect 543230 200701 543290 457811
rect 544404 438054 545004 473498
rect 544404 437818 544586 438054
rect 544822 437818 545004 438054
rect 544404 437734 545004 437818
rect 544404 437498 544586 437734
rect 544822 437498 545004 437734
rect 544404 402054 545004 437498
rect 544404 401818 544586 402054
rect 544822 401818 545004 402054
rect 544404 401734 545004 401818
rect 544404 401498 544586 401734
rect 544822 401498 545004 401734
rect 543411 399532 543477 399533
rect 543411 399468 543412 399532
rect 543476 399468 543477 399532
rect 543411 399467 543477 399468
rect 543414 389061 543474 399467
rect 543411 389060 543477 389061
rect 543411 388996 543412 389060
rect 543476 388996 543477 389060
rect 543411 388995 543477 388996
rect 543411 376684 543477 376685
rect 543411 376620 543412 376684
rect 543476 376620 543477 376684
rect 543411 376619 543477 376620
rect 543414 369749 543474 376619
rect 543411 369748 543477 369749
rect 543411 369684 543412 369748
rect 543476 369684 543477 369748
rect 543411 369683 543477 369684
rect 544404 366054 545004 401498
rect 544404 365818 544586 366054
rect 544822 365818 545004 366054
rect 544404 365734 545004 365818
rect 544404 365498 544586 365734
rect 544822 365498 545004 365734
rect 543411 357372 543477 357373
rect 543411 357308 543412 357372
rect 543476 357308 543477 357372
rect 543411 357307 543477 357308
rect 543414 350437 543474 357307
rect 543411 350436 543477 350437
rect 543411 350372 543412 350436
rect 543476 350372 543477 350436
rect 543411 350371 543477 350372
rect 544404 330054 545004 365498
rect 544404 329818 544586 330054
rect 544822 329818 545004 330054
rect 544404 329734 545004 329818
rect 544404 329498 544586 329734
rect 544822 329498 545004 329734
rect 544404 294054 545004 329498
rect 544404 293818 544586 294054
rect 544822 293818 545004 294054
rect 544404 293734 545004 293818
rect 544404 293498 544586 293734
rect 544822 293498 545004 293734
rect 544404 258054 545004 293498
rect 544404 257818 544586 258054
rect 544822 257818 545004 258054
rect 544404 257734 545004 257818
rect 544404 257498 544586 257734
rect 544822 257498 545004 257734
rect 544404 222054 545004 257498
rect 544404 221818 544586 222054
rect 544822 221818 545004 222054
rect 544404 221734 545004 221818
rect 544404 221498 544586 221734
rect 544822 221498 545004 221734
rect 543227 200700 543293 200701
rect 543227 200636 543228 200700
rect 543292 200636 543293 200700
rect 543227 200635 543293 200636
rect 544404 186054 545004 221498
rect 544404 185818 544586 186054
rect 544822 185818 545004 186054
rect 544404 185734 545004 185818
rect 544404 185498 544586 185734
rect 544822 185498 545004 185734
rect 543043 173908 543109 173909
rect 543043 173844 543044 173908
rect 543108 173844 543109 173908
rect 543043 173843 543109 173844
rect 543046 164253 543106 173843
rect 543043 164252 543109 164253
rect 543043 164188 543044 164252
rect 543108 164188 543109 164252
rect 543043 164187 543109 164188
rect 544404 150054 545004 185498
rect 544404 149818 544586 150054
rect 544822 149818 545004 150054
rect 544404 149734 545004 149818
rect 544404 149498 544586 149734
rect 544822 149498 545004 149734
rect 544404 114054 545004 149498
rect 544404 113818 544586 114054
rect 544822 113818 545004 114054
rect 544404 113734 545004 113818
rect 544404 113498 544586 113734
rect 544822 113498 545004 113734
rect 542859 80068 542925 80069
rect 542859 80004 542860 80068
rect 542924 80004 542925 80068
rect 542859 80003 542925 80004
rect 544404 78054 545004 113498
rect 544404 77818 544586 78054
rect 544822 77818 545004 78054
rect 544404 77734 545004 77818
rect 544404 77498 544586 77734
rect 544822 77498 545004 77734
rect 544404 42054 545004 77498
rect 544404 41818 544586 42054
rect 544822 41818 545004 42054
rect 544404 41734 545004 41818
rect 544404 41498 544586 41734
rect 544822 41498 545004 41734
rect 542675 35868 542741 35869
rect 542675 35804 542676 35868
rect 542740 35804 542741 35868
rect 542675 35803 542741 35804
rect 542491 21996 542557 21997
rect 542491 21932 542492 21996
rect 542556 21932 542557 21996
rect 542491 21931 542557 21932
rect 542307 8260 542373 8261
rect 542307 8196 542308 8260
rect 542372 8196 542373 8260
rect 542307 8195 542373 8196
rect 540804 2218 540986 2454
rect 541222 2218 541404 2454
rect 540804 2134 541404 2218
rect 540804 1898 540986 2134
rect 541222 1898 541404 2134
rect 540804 -346 541404 1898
rect 540804 -582 540986 -346
rect 541222 -582 541404 -346
rect 540804 -666 541404 -582
rect 540804 -902 540986 -666
rect 541222 -902 541404 -666
rect 540804 -1864 541404 -902
rect 544404 6054 545004 41498
rect 544404 5818 544586 6054
rect 544822 5818 545004 6054
rect 544404 5734 545004 5818
rect 544404 5498 544586 5734
rect 544822 5498 545004 5734
rect 544404 -2226 545004 5498
rect 544404 -2462 544586 -2226
rect 544822 -2462 545004 -2226
rect 544404 -2546 545004 -2462
rect 544404 -2782 544586 -2546
rect 544822 -2782 545004 -2546
rect 544404 -3744 545004 -2782
rect 548004 693654 548604 708042
rect 548004 693418 548186 693654
rect 548422 693418 548604 693654
rect 548004 693334 548604 693418
rect 548004 693098 548186 693334
rect 548422 693098 548604 693334
rect 548004 657654 548604 693098
rect 548004 657418 548186 657654
rect 548422 657418 548604 657654
rect 548004 657334 548604 657418
rect 548004 657098 548186 657334
rect 548422 657098 548604 657334
rect 548004 621654 548604 657098
rect 548004 621418 548186 621654
rect 548422 621418 548604 621654
rect 548004 621334 548604 621418
rect 548004 621098 548186 621334
rect 548422 621098 548604 621334
rect 548004 585654 548604 621098
rect 548004 585418 548186 585654
rect 548422 585418 548604 585654
rect 548004 585334 548604 585418
rect 548004 585098 548186 585334
rect 548422 585098 548604 585334
rect 548004 549654 548604 585098
rect 548004 549418 548186 549654
rect 548422 549418 548604 549654
rect 548004 549334 548604 549418
rect 548004 549098 548186 549334
rect 548422 549098 548604 549334
rect 548004 513654 548604 549098
rect 548004 513418 548186 513654
rect 548422 513418 548604 513654
rect 548004 513334 548604 513418
rect 548004 513098 548186 513334
rect 548422 513098 548604 513334
rect 548004 477654 548604 513098
rect 548004 477418 548186 477654
rect 548422 477418 548604 477654
rect 548004 477334 548604 477418
rect 548004 477098 548186 477334
rect 548422 477098 548604 477334
rect 548004 441654 548604 477098
rect 548004 441418 548186 441654
rect 548422 441418 548604 441654
rect 548004 441334 548604 441418
rect 548004 441098 548186 441334
rect 548422 441098 548604 441334
rect 548004 405654 548604 441098
rect 548004 405418 548186 405654
rect 548422 405418 548604 405654
rect 548004 405334 548604 405418
rect 548004 405098 548186 405334
rect 548422 405098 548604 405334
rect 548004 369654 548604 405098
rect 548004 369418 548186 369654
rect 548422 369418 548604 369654
rect 548004 369334 548604 369418
rect 548004 369098 548186 369334
rect 548422 369098 548604 369334
rect 548004 333654 548604 369098
rect 548004 333418 548186 333654
rect 548422 333418 548604 333654
rect 548004 333334 548604 333418
rect 548004 333098 548186 333334
rect 548422 333098 548604 333334
rect 548004 297654 548604 333098
rect 548004 297418 548186 297654
rect 548422 297418 548604 297654
rect 548004 297334 548604 297418
rect 548004 297098 548186 297334
rect 548422 297098 548604 297334
rect 548004 261654 548604 297098
rect 548004 261418 548186 261654
rect 548422 261418 548604 261654
rect 548004 261334 548604 261418
rect 548004 261098 548186 261334
rect 548422 261098 548604 261334
rect 548004 225654 548604 261098
rect 548004 225418 548186 225654
rect 548422 225418 548604 225654
rect 548004 225334 548604 225418
rect 548004 225098 548186 225334
rect 548422 225098 548604 225334
rect 548004 189654 548604 225098
rect 548004 189418 548186 189654
rect 548422 189418 548604 189654
rect 548004 189334 548604 189418
rect 548004 189098 548186 189334
rect 548422 189098 548604 189334
rect 548004 153654 548604 189098
rect 548004 153418 548186 153654
rect 548422 153418 548604 153654
rect 548004 153334 548604 153418
rect 548004 153098 548186 153334
rect 548422 153098 548604 153334
rect 548004 117654 548604 153098
rect 548004 117418 548186 117654
rect 548422 117418 548604 117654
rect 548004 117334 548604 117418
rect 548004 117098 548186 117334
rect 548422 117098 548604 117334
rect 548004 81654 548604 117098
rect 548004 81418 548186 81654
rect 548422 81418 548604 81654
rect 548004 81334 548604 81418
rect 548004 81098 548186 81334
rect 548422 81098 548604 81334
rect 548004 45654 548604 81098
rect 548004 45418 548186 45654
rect 548422 45418 548604 45654
rect 548004 45334 548604 45418
rect 548004 45098 548186 45334
rect 548422 45098 548604 45334
rect 548004 9654 548604 45098
rect 548004 9418 548186 9654
rect 548422 9418 548604 9654
rect 548004 9334 548604 9418
rect 548004 9098 548186 9334
rect 548422 9098 548604 9334
rect 548004 -4106 548604 9098
rect 548004 -4342 548186 -4106
rect 548422 -4342 548604 -4106
rect 548004 -4426 548604 -4342
rect 548004 -4662 548186 -4426
rect 548422 -4662 548604 -4426
rect 548004 -5624 548604 -4662
rect 551604 697254 552204 709922
rect 569604 711418 570204 711440
rect 569604 711182 569786 711418
rect 570022 711182 570204 711418
rect 569604 711098 570204 711182
rect 569604 710862 569786 711098
rect 570022 710862 570204 711098
rect 566004 709538 566604 709560
rect 566004 709302 566186 709538
rect 566422 709302 566604 709538
rect 566004 709218 566604 709302
rect 566004 708982 566186 709218
rect 566422 708982 566604 709218
rect 562404 707658 563004 707680
rect 562404 707422 562586 707658
rect 562822 707422 563004 707658
rect 562404 707338 563004 707422
rect 562404 707102 562586 707338
rect 562822 707102 563004 707338
rect 551604 697018 551786 697254
rect 552022 697018 552204 697254
rect 551604 696934 552204 697018
rect 551604 696698 551786 696934
rect 552022 696698 552204 696934
rect 551604 661254 552204 696698
rect 551604 661018 551786 661254
rect 552022 661018 552204 661254
rect 551604 660934 552204 661018
rect 551604 660698 551786 660934
rect 552022 660698 552204 660934
rect 551604 625254 552204 660698
rect 551604 625018 551786 625254
rect 552022 625018 552204 625254
rect 551604 624934 552204 625018
rect 551604 624698 551786 624934
rect 552022 624698 552204 624934
rect 551604 589254 552204 624698
rect 551604 589018 551786 589254
rect 552022 589018 552204 589254
rect 551604 588934 552204 589018
rect 551604 588698 551786 588934
rect 552022 588698 552204 588934
rect 551604 553254 552204 588698
rect 551604 553018 551786 553254
rect 552022 553018 552204 553254
rect 551604 552934 552204 553018
rect 551604 552698 551786 552934
rect 552022 552698 552204 552934
rect 551604 517254 552204 552698
rect 551604 517018 551786 517254
rect 552022 517018 552204 517254
rect 551604 516934 552204 517018
rect 551604 516698 551786 516934
rect 552022 516698 552204 516934
rect 551604 481254 552204 516698
rect 551604 481018 551786 481254
rect 552022 481018 552204 481254
rect 551604 480934 552204 481018
rect 551604 480698 551786 480934
rect 552022 480698 552204 480934
rect 551604 445254 552204 480698
rect 551604 445018 551786 445254
rect 552022 445018 552204 445254
rect 551604 444934 552204 445018
rect 551604 444698 551786 444934
rect 552022 444698 552204 444934
rect 551604 409254 552204 444698
rect 551604 409018 551786 409254
rect 552022 409018 552204 409254
rect 551604 408934 552204 409018
rect 551604 408698 551786 408934
rect 552022 408698 552204 408934
rect 551604 373254 552204 408698
rect 551604 373018 551786 373254
rect 552022 373018 552204 373254
rect 551604 372934 552204 373018
rect 551604 372698 551786 372934
rect 552022 372698 552204 372934
rect 551604 337254 552204 372698
rect 551604 337018 551786 337254
rect 552022 337018 552204 337254
rect 551604 336934 552204 337018
rect 551604 336698 551786 336934
rect 552022 336698 552204 336934
rect 551604 301254 552204 336698
rect 551604 301018 551786 301254
rect 552022 301018 552204 301254
rect 551604 300934 552204 301018
rect 551604 300698 551786 300934
rect 552022 300698 552204 300934
rect 551604 265254 552204 300698
rect 551604 265018 551786 265254
rect 552022 265018 552204 265254
rect 551604 264934 552204 265018
rect 551604 264698 551786 264934
rect 552022 264698 552204 264934
rect 551604 229254 552204 264698
rect 551604 229018 551786 229254
rect 552022 229018 552204 229254
rect 551604 228934 552204 229018
rect 551604 228698 551786 228934
rect 552022 228698 552204 228934
rect 551604 193254 552204 228698
rect 551604 193018 551786 193254
rect 552022 193018 552204 193254
rect 551604 192934 552204 193018
rect 551604 192698 551786 192934
rect 552022 192698 552204 192934
rect 551604 157254 552204 192698
rect 551604 157018 551786 157254
rect 552022 157018 552204 157254
rect 551604 156934 552204 157018
rect 551604 156698 551786 156934
rect 552022 156698 552204 156934
rect 551604 121254 552204 156698
rect 551604 121018 551786 121254
rect 552022 121018 552204 121254
rect 551604 120934 552204 121018
rect 551604 120698 551786 120934
rect 552022 120698 552204 120934
rect 551604 85254 552204 120698
rect 551604 85018 551786 85254
rect 552022 85018 552204 85254
rect 551604 84934 552204 85018
rect 551604 84698 551786 84934
rect 552022 84698 552204 84934
rect 551604 49254 552204 84698
rect 551604 49018 551786 49254
rect 552022 49018 552204 49254
rect 551604 48934 552204 49018
rect 551604 48698 551786 48934
rect 552022 48698 552204 48934
rect 551604 13254 552204 48698
rect 551604 13018 551786 13254
rect 552022 13018 552204 13254
rect 551604 12934 552204 13018
rect 551604 12698 551786 12934
rect 552022 12698 552204 12934
rect 533604 -7162 533786 -6926
rect 534022 -7162 534204 -6926
rect 533604 -7246 534204 -7162
rect 533604 -7482 533786 -7246
rect 534022 -7482 534204 -7246
rect 533604 -7504 534204 -7482
rect 551604 -5986 552204 12698
rect 558804 705778 559404 705800
rect 558804 705542 558986 705778
rect 559222 705542 559404 705778
rect 558804 705458 559404 705542
rect 558804 705222 558986 705458
rect 559222 705222 559404 705458
rect 558804 668454 559404 705222
rect 558804 668218 558986 668454
rect 559222 668218 559404 668454
rect 558804 668134 559404 668218
rect 558804 667898 558986 668134
rect 559222 667898 559404 668134
rect 558804 632454 559404 667898
rect 558804 632218 558986 632454
rect 559222 632218 559404 632454
rect 558804 632134 559404 632218
rect 558804 631898 558986 632134
rect 559222 631898 559404 632134
rect 558804 596454 559404 631898
rect 558804 596218 558986 596454
rect 559222 596218 559404 596454
rect 558804 596134 559404 596218
rect 558804 595898 558986 596134
rect 559222 595898 559404 596134
rect 558804 560454 559404 595898
rect 558804 560218 558986 560454
rect 559222 560218 559404 560454
rect 558804 560134 559404 560218
rect 558804 559898 558986 560134
rect 559222 559898 559404 560134
rect 558804 524454 559404 559898
rect 558804 524218 558986 524454
rect 559222 524218 559404 524454
rect 558804 524134 559404 524218
rect 558804 523898 558986 524134
rect 559222 523898 559404 524134
rect 558804 488454 559404 523898
rect 558804 488218 558986 488454
rect 559222 488218 559404 488454
rect 558804 488134 559404 488218
rect 558804 487898 558986 488134
rect 559222 487898 559404 488134
rect 558804 452454 559404 487898
rect 558804 452218 558986 452454
rect 559222 452218 559404 452454
rect 558804 452134 559404 452218
rect 558804 451898 558986 452134
rect 559222 451898 559404 452134
rect 558804 416454 559404 451898
rect 558804 416218 558986 416454
rect 559222 416218 559404 416454
rect 558804 416134 559404 416218
rect 558804 415898 558986 416134
rect 559222 415898 559404 416134
rect 558804 380454 559404 415898
rect 558804 380218 558986 380454
rect 559222 380218 559404 380454
rect 558804 380134 559404 380218
rect 558804 379898 558986 380134
rect 559222 379898 559404 380134
rect 558804 344454 559404 379898
rect 558804 344218 558986 344454
rect 559222 344218 559404 344454
rect 558804 344134 559404 344218
rect 558804 343898 558986 344134
rect 559222 343898 559404 344134
rect 558804 308454 559404 343898
rect 558804 308218 558986 308454
rect 559222 308218 559404 308454
rect 558804 308134 559404 308218
rect 558804 307898 558986 308134
rect 559222 307898 559404 308134
rect 558804 272454 559404 307898
rect 558804 272218 558986 272454
rect 559222 272218 559404 272454
rect 558804 272134 559404 272218
rect 558804 271898 558986 272134
rect 559222 271898 559404 272134
rect 558804 236454 559404 271898
rect 558804 236218 558986 236454
rect 559222 236218 559404 236454
rect 558804 236134 559404 236218
rect 558804 235898 558986 236134
rect 559222 235898 559404 236134
rect 558804 200454 559404 235898
rect 558804 200218 558986 200454
rect 559222 200218 559404 200454
rect 558804 200134 559404 200218
rect 558804 199898 558986 200134
rect 559222 199898 559404 200134
rect 558804 164454 559404 199898
rect 558804 164218 558986 164454
rect 559222 164218 559404 164454
rect 558804 164134 559404 164218
rect 558804 163898 558986 164134
rect 559222 163898 559404 164134
rect 558804 128454 559404 163898
rect 558804 128218 558986 128454
rect 559222 128218 559404 128454
rect 558804 128134 559404 128218
rect 558804 127898 558986 128134
rect 559222 127898 559404 128134
rect 558804 92454 559404 127898
rect 558804 92218 558986 92454
rect 559222 92218 559404 92454
rect 558804 92134 559404 92218
rect 558804 91898 558986 92134
rect 559222 91898 559404 92134
rect 558804 56454 559404 91898
rect 558804 56218 558986 56454
rect 559222 56218 559404 56454
rect 558804 56134 559404 56218
rect 558804 55898 558986 56134
rect 559222 55898 559404 56134
rect 558804 20454 559404 55898
rect 558804 20218 558986 20454
rect 559222 20218 559404 20454
rect 558804 20134 559404 20218
rect 558804 19898 558986 20134
rect 559222 19898 559404 20134
rect 558804 -1286 559404 19898
rect 558804 -1522 558986 -1286
rect 559222 -1522 559404 -1286
rect 558804 -1606 559404 -1522
rect 558804 -1842 558986 -1606
rect 559222 -1842 559404 -1606
rect 558804 -1864 559404 -1842
rect 562404 672054 563004 707102
rect 562404 671818 562586 672054
rect 562822 671818 563004 672054
rect 562404 671734 563004 671818
rect 562404 671498 562586 671734
rect 562822 671498 563004 671734
rect 562404 636054 563004 671498
rect 562404 635818 562586 636054
rect 562822 635818 563004 636054
rect 562404 635734 563004 635818
rect 562404 635498 562586 635734
rect 562822 635498 563004 635734
rect 562404 600054 563004 635498
rect 562404 599818 562586 600054
rect 562822 599818 563004 600054
rect 562404 599734 563004 599818
rect 562404 599498 562586 599734
rect 562822 599498 563004 599734
rect 562404 564054 563004 599498
rect 562404 563818 562586 564054
rect 562822 563818 563004 564054
rect 562404 563734 563004 563818
rect 562404 563498 562586 563734
rect 562822 563498 563004 563734
rect 562404 528054 563004 563498
rect 562404 527818 562586 528054
rect 562822 527818 563004 528054
rect 562404 527734 563004 527818
rect 562404 527498 562586 527734
rect 562822 527498 563004 527734
rect 562404 492054 563004 527498
rect 562404 491818 562586 492054
rect 562822 491818 563004 492054
rect 562404 491734 563004 491818
rect 562404 491498 562586 491734
rect 562822 491498 563004 491734
rect 562404 456054 563004 491498
rect 562404 455818 562586 456054
rect 562822 455818 563004 456054
rect 562404 455734 563004 455818
rect 562404 455498 562586 455734
rect 562822 455498 563004 455734
rect 562404 420054 563004 455498
rect 562404 419818 562586 420054
rect 562822 419818 563004 420054
rect 562404 419734 563004 419818
rect 562404 419498 562586 419734
rect 562822 419498 563004 419734
rect 562404 384054 563004 419498
rect 562404 383818 562586 384054
rect 562822 383818 563004 384054
rect 562404 383734 563004 383818
rect 562404 383498 562586 383734
rect 562822 383498 563004 383734
rect 562404 348054 563004 383498
rect 562404 347818 562586 348054
rect 562822 347818 563004 348054
rect 562404 347734 563004 347818
rect 562404 347498 562586 347734
rect 562822 347498 563004 347734
rect 562404 312054 563004 347498
rect 562404 311818 562586 312054
rect 562822 311818 563004 312054
rect 562404 311734 563004 311818
rect 562404 311498 562586 311734
rect 562822 311498 563004 311734
rect 562404 276054 563004 311498
rect 562404 275818 562586 276054
rect 562822 275818 563004 276054
rect 562404 275734 563004 275818
rect 562404 275498 562586 275734
rect 562822 275498 563004 275734
rect 562404 240054 563004 275498
rect 562404 239818 562586 240054
rect 562822 239818 563004 240054
rect 562404 239734 563004 239818
rect 562404 239498 562586 239734
rect 562822 239498 563004 239734
rect 562404 204054 563004 239498
rect 562404 203818 562586 204054
rect 562822 203818 563004 204054
rect 562404 203734 563004 203818
rect 562404 203498 562586 203734
rect 562822 203498 563004 203734
rect 562404 168054 563004 203498
rect 562404 167818 562586 168054
rect 562822 167818 563004 168054
rect 562404 167734 563004 167818
rect 562404 167498 562586 167734
rect 562822 167498 563004 167734
rect 562404 132054 563004 167498
rect 562404 131818 562586 132054
rect 562822 131818 563004 132054
rect 562404 131734 563004 131818
rect 562404 131498 562586 131734
rect 562822 131498 563004 131734
rect 562404 96054 563004 131498
rect 562404 95818 562586 96054
rect 562822 95818 563004 96054
rect 562404 95734 563004 95818
rect 562404 95498 562586 95734
rect 562822 95498 563004 95734
rect 562404 60054 563004 95498
rect 562404 59818 562586 60054
rect 562822 59818 563004 60054
rect 562404 59734 563004 59818
rect 562404 59498 562586 59734
rect 562822 59498 563004 59734
rect 562404 24054 563004 59498
rect 562404 23818 562586 24054
rect 562822 23818 563004 24054
rect 562404 23734 563004 23818
rect 562404 23498 562586 23734
rect 562822 23498 563004 23734
rect 562404 -3166 563004 23498
rect 562404 -3402 562586 -3166
rect 562822 -3402 563004 -3166
rect 562404 -3486 563004 -3402
rect 562404 -3722 562586 -3486
rect 562822 -3722 563004 -3486
rect 562404 -3744 563004 -3722
rect 566004 675654 566604 708982
rect 566004 675418 566186 675654
rect 566422 675418 566604 675654
rect 566004 675334 566604 675418
rect 566004 675098 566186 675334
rect 566422 675098 566604 675334
rect 566004 639654 566604 675098
rect 566004 639418 566186 639654
rect 566422 639418 566604 639654
rect 566004 639334 566604 639418
rect 566004 639098 566186 639334
rect 566422 639098 566604 639334
rect 566004 603654 566604 639098
rect 566004 603418 566186 603654
rect 566422 603418 566604 603654
rect 566004 603334 566604 603418
rect 566004 603098 566186 603334
rect 566422 603098 566604 603334
rect 566004 567654 566604 603098
rect 566004 567418 566186 567654
rect 566422 567418 566604 567654
rect 566004 567334 566604 567418
rect 566004 567098 566186 567334
rect 566422 567098 566604 567334
rect 566004 531654 566604 567098
rect 566004 531418 566186 531654
rect 566422 531418 566604 531654
rect 566004 531334 566604 531418
rect 566004 531098 566186 531334
rect 566422 531098 566604 531334
rect 566004 495654 566604 531098
rect 566004 495418 566186 495654
rect 566422 495418 566604 495654
rect 566004 495334 566604 495418
rect 566004 495098 566186 495334
rect 566422 495098 566604 495334
rect 566004 459654 566604 495098
rect 566004 459418 566186 459654
rect 566422 459418 566604 459654
rect 566004 459334 566604 459418
rect 566004 459098 566186 459334
rect 566422 459098 566604 459334
rect 566004 423654 566604 459098
rect 566004 423418 566186 423654
rect 566422 423418 566604 423654
rect 566004 423334 566604 423418
rect 566004 423098 566186 423334
rect 566422 423098 566604 423334
rect 566004 387654 566604 423098
rect 566004 387418 566186 387654
rect 566422 387418 566604 387654
rect 566004 387334 566604 387418
rect 566004 387098 566186 387334
rect 566422 387098 566604 387334
rect 566004 351654 566604 387098
rect 566004 351418 566186 351654
rect 566422 351418 566604 351654
rect 566004 351334 566604 351418
rect 566004 351098 566186 351334
rect 566422 351098 566604 351334
rect 566004 315654 566604 351098
rect 566004 315418 566186 315654
rect 566422 315418 566604 315654
rect 566004 315334 566604 315418
rect 566004 315098 566186 315334
rect 566422 315098 566604 315334
rect 566004 279654 566604 315098
rect 566004 279418 566186 279654
rect 566422 279418 566604 279654
rect 566004 279334 566604 279418
rect 566004 279098 566186 279334
rect 566422 279098 566604 279334
rect 566004 243654 566604 279098
rect 566004 243418 566186 243654
rect 566422 243418 566604 243654
rect 566004 243334 566604 243418
rect 566004 243098 566186 243334
rect 566422 243098 566604 243334
rect 566004 207654 566604 243098
rect 566004 207418 566186 207654
rect 566422 207418 566604 207654
rect 566004 207334 566604 207418
rect 566004 207098 566186 207334
rect 566422 207098 566604 207334
rect 566004 171654 566604 207098
rect 566004 171418 566186 171654
rect 566422 171418 566604 171654
rect 566004 171334 566604 171418
rect 566004 171098 566186 171334
rect 566422 171098 566604 171334
rect 566004 135654 566604 171098
rect 566004 135418 566186 135654
rect 566422 135418 566604 135654
rect 566004 135334 566604 135418
rect 566004 135098 566186 135334
rect 566422 135098 566604 135334
rect 566004 99654 566604 135098
rect 566004 99418 566186 99654
rect 566422 99418 566604 99654
rect 566004 99334 566604 99418
rect 566004 99098 566186 99334
rect 566422 99098 566604 99334
rect 566004 63654 566604 99098
rect 566004 63418 566186 63654
rect 566422 63418 566604 63654
rect 566004 63334 566604 63418
rect 566004 63098 566186 63334
rect 566422 63098 566604 63334
rect 566004 27654 566604 63098
rect 566004 27418 566186 27654
rect 566422 27418 566604 27654
rect 566004 27334 566604 27418
rect 566004 27098 566186 27334
rect 566422 27098 566604 27334
rect 566004 -5046 566604 27098
rect 566004 -5282 566186 -5046
rect 566422 -5282 566604 -5046
rect 566004 -5366 566604 -5282
rect 566004 -5602 566186 -5366
rect 566422 -5602 566604 -5366
rect 566004 -5624 566604 -5602
rect 569604 679254 570204 710862
rect 591900 711418 592500 711440
rect 591900 711182 592082 711418
rect 592318 711182 592500 711418
rect 591900 711098 592500 711182
rect 591900 710862 592082 711098
rect 592318 710862 592500 711098
rect 590960 710478 591560 710500
rect 590960 710242 591142 710478
rect 591378 710242 591560 710478
rect 590960 710158 591560 710242
rect 590960 709922 591142 710158
rect 591378 709922 591560 710158
rect 590020 709538 590620 709560
rect 590020 709302 590202 709538
rect 590438 709302 590620 709538
rect 590020 709218 590620 709302
rect 590020 708982 590202 709218
rect 590438 708982 590620 709218
rect 589080 708598 589680 708620
rect 589080 708362 589262 708598
rect 589498 708362 589680 708598
rect 589080 708278 589680 708362
rect 589080 708042 589262 708278
rect 589498 708042 589680 708278
rect 580404 706718 581004 707680
rect 588140 707658 588740 707680
rect 588140 707422 588322 707658
rect 588558 707422 588740 707658
rect 588140 707338 588740 707422
rect 588140 707102 588322 707338
rect 588558 707102 588740 707338
rect 580404 706482 580586 706718
rect 580822 706482 581004 706718
rect 580404 706398 581004 706482
rect 580404 706162 580586 706398
rect 580822 706162 581004 706398
rect 569604 679018 569786 679254
rect 570022 679018 570204 679254
rect 569604 678934 570204 679018
rect 569604 678698 569786 678934
rect 570022 678698 570204 678934
rect 569604 643254 570204 678698
rect 569604 643018 569786 643254
rect 570022 643018 570204 643254
rect 569604 642934 570204 643018
rect 569604 642698 569786 642934
rect 570022 642698 570204 642934
rect 569604 607254 570204 642698
rect 569604 607018 569786 607254
rect 570022 607018 570204 607254
rect 569604 606934 570204 607018
rect 569604 606698 569786 606934
rect 570022 606698 570204 606934
rect 569604 571254 570204 606698
rect 569604 571018 569786 571254
rect 570022 571018 570204 571254
rect 569604 570934 570204 571018
rect 569604 570698 569786 570934
rect 570022 570698 570204 570934
rect 569604 535254 570204 570698
rect 569604 535018 569786 535254
rect 570022 535018 570204 535254
rect 569604 534934 570204 535018
rect 569604 534698 569786 534934
rect 570022 534698 570204 534934
rect 569604 499254 570204 534698
rect 569604 499018 569786 499254
rect 570022 499018 570204 499254
rect 569604 498934 570204 499018
rect 569604 498698 569786 498934
rect 570022 498698 570204 498934
rect 569604 463254 570204 498698
rect 569604 463018 569786 463254
rect 570022 463018 570204 463254
rect 569604 462934 570204 463018
rect 569604 462698 569786 462934
rect 570022 462698 570204 462934
rect 569604 427254 570204 462698
rect 569604 427018 569786 427254
rect 570022 427018 570204 427254
rect 569604 426934 570204 427018
rect 569604 426698 569786 426934
rect 570022 426698 570204 426934
rect 569604 391254 570204 426698
rect 569604 391018 569786 391254
rect 570022 391018 570204 391254
rect 569604 390934 570204 391018
rect 569604 390698 569786 390934
rect 570022 390698 570204 390934
rect 569604 355254 570204 390698
rect 569604 355018 569786 355254
rect 570022 355018 570204 355254
rect 569604 354934 570204 355018
rect 569604 354698 569786 354934
rect 570022 354698 570204 354934
rect 569604 319254 570204 354698
rect 569604 319018 569786 319254
rect 570022 319018 570204 319254
rect 569604 318934 570204 319018
rect 569604 318698 569786 318934
rect 570022 318698 570204 318934
rect 569604 283254 570204 318698
rect 569604 283018 569786 283254
rect 570022 283018 570204 283254
rect 569604 282934 570204 283018
rect 569604 282698 569786 282934
rect 570022 282698 570204 282934
rect 569604 247254 570204 282698
rect 569604 247018 569786 247254
rect 570022 247018 570204 247254
rect 569604 246934 570204 247018
rect 569604 246698 569786 246934
rect 570022 246698 570204 246934
rect 569604 211254 570204 246698
rect 569604 211018 569786 211254
rect 570022 211018 570204 211254
rect 569604 210934 570204 211018
rect 569604 210698 569786 210934
rect 570022 210698 570204 210934
rect 569604 175254 570204 210698
rect 569604 175018 569786 175254
rect 570022 175018 570204 175254
rect 569604 174934 570204 175018
rect 569604 174698 569786 174934
rect 570022 174698 570204 174934
rect 569604 139254 570204 174698
rect 569604 139018 569786 139254
rect 570022 139018 570204 139254
rect 569604 138934 570204 139018
rect 569604 138698 569786 138934
rect 570022 138698 570204 138934
rect 569604 103254 570204 138698
rect 569604 103018 569786 103254
rect 570022 103018 570204 103254
rect 569604 102934 570204 103018
rect 569604 102698 569786 102934
rect 570022 102698 570204 102934
rect 569604 67254 570204 102698
rect 569604 67018 569786 67254
rect 570022 67018 570204 67254
rect 569604 66934 570204 67018
rect 569604 66698 569786 66934
rect 570022 66698 570204 66934
rect 569604 31254 570204 66698
rect 569604 31018 569786 31254
rect 570022 31018 570204 31254
rect 569604 30934 570204 31018
rect 569604 30698 569786 30934
rect 570022 30698 570204 30934
rect 551604 -6222 551786 -5986
rect 552022 -6222 552204 -5986
rect 551604 -6306 552204 -6222
rect 551604 -6542 551786 -6306
rect 552022 -6542 552204 -6306
rect 551604 -7504 552204 -6542
rect 569604 -6926 570204 30698
rect 576804 704838 577404 705800
rect 576804 704602 576986 704838
rect 577222 704602 577404 704838
rect 576804 704518 577404 704602
rect 576804 704282 576986 704518
rect 577222 704282 577404 704518
rect 576804 686454 577404 704282
rect 576804 686218 576986 686454
rect 577222 686218 577404 686454
rect 576804 686134 577404 686218
rect 576804 685898 576986 686134
rect 577222 685898 577404 686134
rect 576804 650454 577404 685898
rect 576804 650218 576986 650454
rect 577222 650218 577404 650454
rect 576804 650134 577404 650218
rect 576804 649898 576986 650134
rect 577222 649898 577404 650134
rect 576804 614454 577404 649898
rect 576804 614218 576986 614454
rect 577222 614218 577404 614454
rect 576804 614134 577404 614218
rect 576804 613898 576986 614134
rect 577222 613898 577404 614134
rect 576804 578454 577404 613898
rect 576804 578218 576986 578454
rect 577222 578218 577404 578454
rect 576804 578134 577404 578218
rect 576804 577898 576986 578134
rect 577222 577898 577404 578134
rect 576804 542454 577404 577898
rect 576804 542218 576986 542454
rect 577222 542218 577404 542454
rect 576804 542134 577404 542218
rect 576804 541898 576986 542134
rect 577222 541898 577404 542134
rect 576804 506454 577404 541898
rect 576804 506218 576986 506454
rect 577222 506218 577404 506454
rect 576804 506134 577404 506218
rect 576804 505898 576986 506134
rect 577222 505898 577404 506134
rect 576804 470454 577404 505898
rect 576804 470218 576986 470454
rect 577222 470218 577404 470454
rect 576804 470134 577404 470218
rect 576804 469898 576986 470134
rect 577222 469898 577404 470134
rect 576804 434454 577404 469898
rect 576804 434218 576986 434454
rect 577222 434218 577404 434454
rect 576804 434134 577404 434218
rect 576804 433898 576986 434134
rect 577222 433898 577404 434134
rect 576804 398454 577404 433898
rect 576804 398218 576986 398454
rect 577222 398218 577404 398454
rect 576804 398134 577404 398218
rect 576804 397898 576986 398134
rect 577222 397898 577404 398134
rect 576804 362454 577404 397898
rect 576804 362218 576986 362454
rect 577222 362218 577404 362454
rect 576804 362134 577404 362218
rect 576804 361898 576986 362134
rect 577222 361898 577404 362134
rect 576804 326454 577404 361898
rect 576804 326218 576986 326454
rect 577222 326218 577404 326454
rect 576804 326134 577404 326218
rect 576804 325898 576986 326134
rect 577222 325898 577404 326134
rect 576804 290454 577404 325898
rect 576804 290218 576986 290454
rect 577222 290218 577404 290454
rect 576804 290134 577404 290218
rect 576804 289898 576986 290134
rect 577222 289898 577404 290134
rect 576804 254454 577404 289898
rect 576804 254218 576986 254454
rect 577222 254218 577404 254454
rect 576804 254134 577404 254218
rect 576804 253898 576986 254134
rect 577222 253898 577404 254134
rect 576804 218454 577404 253898
rect 576804 218218 576986 218454
rect 577222 218218 577404 218454
rect 576804 218134 577404 218218
rect 576804 217898 576986 218134
rect 577222 217898 577404 218134
rect 576804 182454 577404 217898
rect 576804 182218 576986 182454
rect 577222 182218 577404 182454
rect 576804 182134 577404 182218
rect 576804 181898 576986 182134
rect 577222 181898 577404 182134
rect 576804 146454 577404 181898
rect 576804 146218 576986 146454
rect 577222 146218 577404 146454
rect 576804 146134 577404 146218
rect 576804 145898 576986 146134
rect 577222 145898 577404 146134
rect 576804 110454 577404 145898
rect 576804 110218 576986 110454
rect 577222 110218 577404 110454
rect 576804 110134 577404 110218
rect 576804 109898 576986 110134
rect 577222 109898 577404 110134
rect 576804 74454 577404 109898
rect 576804 74218 576986 74454
rect 577222 74218 577404 74454
rect 576804 74134 577404 74218
rect 576804 73898 576986 74134
rect 577222 73898 577404 74134
rect 576804 38454 577404 73898
rect 576804 38218 576986 38454
rect 577222 38218 577404 38454
rect 576804 38134 577404 38218
rect 576804 37898 576986 38134
rect 577222 37898 577404 38134
rect 576804 2454 577404 37898
rect 576804 2218 576986 2454
rect 577222 2218 577404 2454
rect 576804 2134 577404 2218
rect 576804 1898 576986 2134
rect 577222 1898 577404 2134
rect 576804 -346 577404 1898
rect 576804 -582 576986 -346
rect 577222 -582 577404 -346
rect 576804 -666 577404 -582
rect 576804 -902 576986 -666
rect 577222 -902 577404 -666
rect 576804 -1864 577404 -902
rect 580404 690054 581004 706162
rect 587200 706718 587800 706740
rect 587200 706482 587382 706718
rect 587618 706482 587800 706718
rect 587200 706398 587800 706482
rect 587200 706162 587382 706398
rect 587618 706162 587800 706398
rect 586260 705778 586860 705800
rect 586260 705542 586442 705778
rect 586678 705542 586860 705778
rect 586260 705458 586860 705542
rect 586260 705222 586442 705458
rect 586678 705222 586860 705458
rect 580404 689818 580586 690054
rect 580822 689818 581004 690054
rect 580404 689734 581004 689818
rect 580404 689498 580586 689734
rect 580822 689498 581004 689734
rect 580404 654054 581004 689498
rect 580404 653818 580586 654054
rect 580822 653818 581004 654054
rect 580404 653734 581004 653818
rect 580404 653498 580586 653734
rect 580822 653498 581004 653734
rect 580404 618054 581004 653498
rect 580404 617818 580586 618054
rect 580822 617818 581004 618054
rect 580404 617734 581004 617818
rect 580404 617498 580586 617734
rect 580822 617498 581004 617734
rect 580404 582054 581004 617498
rect 580404 581818 580586 582054
rect 580822 581818 581004 582054
rect 580404 581734 581004 581818
rect 580404 581498 580586 581734
rect 580822 581498 581004 581734
rect 580404 546054 581004 581498
rect 580404 545818 580586 546054
rect 580822 545818 581004 546054
rect 580404 545734 581004 545818
rect 580404 545498 580586 545734
rect 580822 545498 581004 545734
rect 580404 510054 581004 545498
rect 580404 509818 580586 510054
rect 580822 509818 581004 510054
rect 580404 509734 581004 509818
rect 580404 509498 580586 509734
rect 580822 509498 581004 509734
rect 580404 474054 581004 509498
rect 580404 473818 580586 474054
rect 580822 473818 581004 474054
rect 580404 473734 581004 473818
rect 580404 473498 580586 473734
rect 580822 473498 581004 473734
rect 580404 438054 581004 473498
rect 580404 437818 580586 438054
rect 580822 437818 581004 438054
rect 580404 437734 581004 437818
rect 580404 437498 580586 437734
rect 580822 437498 581004 437734
rect 580404 402054 581004 437498
rect 580404 401818 580586 402054
rect 580822 401818 581004 402054
rect 580404 401734 581004 401818
rect 580404 401498 580586 401734
rect 580822 401498 581004 401734
rect 580404 366054 581004 401498
rect 580404 365818 580586 366054
rect 580822 365818 581004 366054
rect 580404 365734 581004 365818
rect 580404 365498 580586 365734
rect 580822 365498 581004 365734
rect 580404 330054 581004 365498
rect 580404 329818 580586 330054
rect 580822 329818 581004 330054
rect 580404 329734 581004 329818
rect 580404 329498 580586 329734
rect 580822 329498 581004 329734
rect 580404 294054 581004 329498
rect 580404 293818 580586 294054
rect 580822 293818 581004 294054
rect 580404 293734 581004 293818
rect 580404 293498 580586 293734
rect 580822 293498 581004 293734
rect 580404 258054 581004 293498
rect 580404 257818 580586 258054
rect 580822 257818 581004 258054
rect 580404 257734 581004 257818
rect 580404 257498 580586 257734
rect 580822 257498 581004 257734
rect 580404 222054 581004 257498
rect 580404 221818 580586 222054
rect 580822 221818 581004 222054
rect 580404 221734 581004 221818
rect 580404 221498 580586 221734
rect 580822 221498 581004 221734
rect 580404 186054 581004 221498
rect 580404 185818 580586 186054
rect 580822 185818 581004 186054
rect 580404 185734 581004 185818
rect 580404 185498 580586 185734
rect 580822 185498 581004 185734
rect 580404 150054 581004 185498
rect 580404 149818 580586 150054
rect 580822 149818 581004 150054
rect 580404 149734 581004 149818
rect 580404 149498 580586 149734
rect 580822 149498 581004 149734
rect 580404 114054 581004 149498
rect 580404 113818 580586 114054
rect 580822 113818 581004 114054
rect 580404 113734 581004 113818
rect 580404 113498 580586 113734
rect 580822 113498 581004 113734
rect 580404 78054 581004 113498
rect 580404 77818 580586 78054
rect 580822 77818 581004 78054
rect 580404 77734 581004 77818
rect 580404 77498 580586 77734
rect 580822 77498 581004 77734
rect 580404 42054 581004 77498
rect 580404 41818 580586 42054
rect 580822 41818 581004 42054
rect 580404 41734 581004 41818
rect 580404 41498 580586 41734
rect 580822 41498 581004 41734
rect 580404 6054 581004 41498
rect 580404 5818 580586 6054
rect 580822 5818 581004 6054
rect 580404 5734 581004 5818
rect 580404 5498 580586 5734
rect 580822 5498 581004 5734
rect 580404 -2226 581004 5498
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 585320 686454 585920 704282
rect 585320 686218 585502 686454
rect 585738 686218 585920 686454
rect 585320 686134 585920 686218
rect 585320 685898 585502 686134
rect 585738 685898 585920 686134
rect 585320 650454 585920 685898
rect 585320 650218 585502 650454
rect 585738 650218 585920 650454
rect 585320 650134 585920 650218
rect 585320 649898 585502 650134
rect 585738 649898 585920 650134
rect 585320 614454 585920 649898
rect 585320 614218 585502 614454
rect 585738 614218 585920 614454
rect 585320 614134 585920 614218
rect 585320 613898 585502 614134
rect 585738 613898 585920 614134
rect 585320 578454 585920 613898
rect 585320 578218 585502 578454
rect 585738 578218 585920 578454
rect 585320 578134 585920 578218
rect 585320 577898 585502 578134
rect 585738 577898 585920 578134
rect 585320 542454 585920 577898
rect 585320 542218 585502 542454
rect 585738 542218 585920 542454
rect 585320 542134 585920 542218
rect 585320 541898 585502 542134
rect 585738 541898 585920 542134
rect 585320 506454 585920 541898
rect 585320 506218 585502 506454
rect 585738 506218 585920 506454
rect 585320 506134 585920 506218
rect 585320 505898 585502 506134
rect 585738 505898 585920 506134
rect 585320 470454 585920 505898
rect 585320 470218 585502 470454
rect 585738 470218 585920 470454
rect 585320 470134 585920 470218
rect 585320 469898 585502 470134
rect 585738 469898 585920 470134
rect 585320 434454 585920 469898
rect 585320 434218 585502 434454
rect 585738 434218 585920 434454
rect 585320 434134 585920 434218
rect 585320 433898 585502 434134
rect 585738 433898 585920 434134
rect 585320 398454 585920 433898
rect 585320 398218 585502 398454
rect 585738 398218 585920 398454
rect 585320 398134 585920 398218
rect 585320 397898 585502 398134
rect 585738 397898 585920 398134
rect 585320 362454 585920 397898
rect 585320 362218 585502 362454
rect 585738 362218 585920 362454
rect 585320 362134 585920 362218
rect 585320 361898 585502 362134
rect 585738 361898 585920 362134
rect 585320 326454 585920 361898
rect 585320 326218 585502 326454
rect 585738 326218 585920 326454
rect 585320 326134 585920 326218
rect 585320 325898 585502 326134
rect 585738 325898 585920 326134
rect 585320 290454 585920 325898
rect 585320 290218 585502 290454
rect 585738 290218 585920 290454
rect 585320 290134 585920 290218
rect 585320 289898 585502 290134
rect 585738 289898 585920 290134
rect 585320 254454 585920 289898
rect 585320 254218 585502 254454
rect 585738 254218 585920 254454
rect 585320 254134 585920 254218
rect 585320 253898 585502 254134
rect 585738 253898 585920 254134
rect 585320 218454 585920 253898
rect 585320 218218 585502 218454
rect 585738 218218 585920 218454
rect 585320 218134 585920 218218
rect 585320 217898 585502 218134
rect 585738 217898 585920 218134
rect 585320 182454 585920 217898
rect 585320 182218 585502 182454
rect 585738 182218 585920 182454
rect 585320 182134 585920 182218
rect 585320 181898 585502 182134
rect 585738 181898 585920 182134
rect 585320 146454 585920 181898
rect 585320 146218 585502 146454
rect 585738 146218 585920 146454
rect 585320 146134 585920 146218
rect 585320 145898 585502 146134
rect 585738 145898 585920 146134
rect 585320 110454 585920 145898
rect 585320 110218 585502 110454
rect 585738 110218 585920 110454
rect 585320 110134 585920 110218
rect 585320 109898 585502 110134
rect 585738 109898 585920 110134
rect 585320 74454 585920 109898
rect 585320 74218 585502 74454
rect 585738 74218 585920 74454
rect 585320 74134 585920 74218
rect 585320 73898 585502 74134
rect 585738 73898 585920 74134
rect 585320 38454 585920 73898
rect 585320 38218 585502 38454
rect 585738 38218 585920 38454
rect 585320 38134 585920 38218
rect 585320 37898 585502 38134
rect 585738 37898 585920 38134
rect 585320 2454 585920 37898
rect 585320 2218 585502 2454
rect 585738 2218 585920 2454
rect 585320 2134 585920 2218
rect 585320 1898 585502 2134
rect 585738 1898 585920 2134
rect 585320 -346 585920 1898
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586260 668454 586860 705222
rect 586260 668218 586442 668454
rect 586678 668218 586860 668454
rect 586260 668134 586860 668218
rect 586260 667898 586442 668134
rect 586678 667898 586860 668134
rect 586260 632454 586860 667898
rect 586260 632218 586442 632454
rect 586678 632218 586860 632454
rect 586260 632134 586860 632218
rect 586260 631898 586442 632134
rect 586678 631898 586860 632134
rect 586260 596454 586860 631898
rect 586260 596218 586442 596454
rect 586678 596218 586860 596454
rect 586260 596134 586860 596218
rect 586260 595898 586442 596134
rect 586678 595898 586860 596134
rect 586260 560454 586860 595898
rect 586260 560218 586442 560454
rect 586678 560218 586860 560454
rect 586260 560134 586860 560218
rect 586260 559898 586442 560134
rect 586678 559898 586860 560134
rect 586260 524454 586860 559898
rect 586260 524218 586442 524454
rect 586678 524218 586860 524454
rect 586260 524134 586860 524218
rect 586260 523898 586442 524134
rect 586678 523898 586860 524134
rect 586260 488454 586860 523898
rect 586260 488218 586442 488454
rect 586678 488218 586860 488454
rect 586260 488134 586860 488218
rect 586260 487898 586442 488134
rect 586678 487898 586860 488134
rect 586260 452454 586860 487898
rect 586260 452218 586442 452454
rect 586678 452218 586860 452454
rect 586260 452134 586860 452218
rect 586260 451898 586442 452134
rect 586678 451898 586860 452134
rect 586260 416454 586860 451898
rect 586260 416218 586442 416454
rect 586678 416218 586860 416454
rect 586260 416134 586860 416218
rect 586260 415898 586442 416134
rect 586678 415898 586860 416134
rect 586260 380454 586860 415898
rect 586260 380218 586442 380454
rect 586678 380218 586860 380454
rect 586260 380134 586860 380218
rect 586260 379898 586442 380134
rect 586678 379898 586860 380134
rect 586260 344454 586860 379898
rect 586260 344218 586442 344454
rect 586678 344218 586860 344454
rect 586260 344134 586860 344218
rect 586260 343898 586442 344134
rect 586678 343898 586860 344134
rect 586260 308454 586860 343898
rect 586260 308218 586442 308454
rect 586678 308218 586860 308454
rect 586260 308134 586860 308218
rect 586260 307898 586442 308134
rect 586678 307898 586860 308134
rect 586260 272454 586860 307898
rect 586260 272218 586442 272454
rect 586678 272218 586860 272454
rect 586260 272134 586860 272218
rect 586260 271898 586442 272134
rect 586678 271898 586860 272134
rect 586260 236454 586860 271898
rect 586260 236218 586442 236454
rect 586678 236218 586860 236454
rect 586260 236134 586860 236218
rect 586260 235898 586442 236134
rect 586678 235898 586860 236134
rect 586260 200454 586860 235898
rect 586260 200218 586442 200454
rect 586678 200218 586860 200454
rect 586260 200134 586860 200218
rect 586260 199898 586442 200134
rect 586678 199898 586860 200134
rect 586260 164454 586860 199898
rect 586260 164218 586442 164454
rect 586678 164218 586860 164454
rect 586260 164134 586860 164218
rect 586260 163898 586442 164134
rect 586678 163898 586860 164134
rect 586260 128454 586860 163898
rect 586260 128218 586442 128454
rect 586678 128218 586860 128454
rect 586260 128134 586860 128218
rect 586260 127898 586442 128134
rect 586678 127898 586860 128134
rect 586260 92454 586860 127898
rect 586260 92218 586442 92454
rect 586678 92218 586860 92454
rect 586260 92134 586860 92218
rect 586260 91898 586442 92134
rect 586678 91898 586860 92134
rect 586260 56454 586860 91898
rect 586260 56218 586442 56454
rect 586678 56218 586860 56454
rect 586260 56134 586860 56218
rect 586260 55898 586442 56134
rect 586678 55898 586860 56134
rect 586260 20454 586860 55898
rect 586260 20218 586442 20454
rect 586678 20218 586860 20454
rect 586260 20134 586860 20218
rect 586260 19898 586442 20134
rect 586678 19898 586860 20134
rect 586260 -1286 586860 19898
rect 586260 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect 586260 -1606 586860 -1522
rect 586260 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect 586260 -1864 586860 -1842
rect 587200 690054 587800 706162
rect 587200 689818 587382 690054
rect 587618 689818 587800 690054
rect 587200 689734 587800 689818
rect 587200 689498 587382 689734
rect 587618 689498 587800 689734
rect 587200 654054 587800 689498
rect 587200 653818 587382 654054
rect 587618 653818 587800 654054
rect 587200 653734 587800 653818
rect 587200 653498 587382 653734
rect 587618 653498 587800 653734
rect 587200 618054 587800 653498
rect 587200 617818 587382 618054
rect 587618 617818 587800 618054
rect 587200 617734 587800 617818
rect 587200 617498 587382 617734
rect 587618 617498 587800 617734
rect 587200 582054 587800 617498
rect 587200 581818 587382 582054
rect 587618 581818 587800 582054
rect 587200 581734 587800 581818
rect 587200 581498 587382 581734
rect 587618 581498 587800 581734
rect 587200 546054 587800 581498
rect 587200 545818 587382 546054
rect 587618 545818 587800 546054
rect 587200 545734 587800 545818
rect 587200 545498 587382 545734
rect 587618 545498 587800 545734
rect 587200 510054 587800 545498
rect 587200 509818 587382 510054
rect 587618 509818 587800 510054
rect 587200 509734 587800 509818
rect 587200 509498 587382 509734
rect 587618 509498 587800 509734
rect 587200 474054 587800 509498
rect 587200 473818 587382 474054
rect 587618 473818 587800 474054
rect 587200 473734 587800 473818
rect 587200 473498 587382 473734
rect 587618 473498 587800 473734
rect 587200 438054 587800 473498
rect 587200 437818 587382 438054
rect 587618 437818 587800 438054
rect 587200 437734 587800 437818
rect 587200 437498 587382 437734
rect 587618 437498 587800 437734
rect 587200 402054 587800 437498
rect 587200 401818 587382 402054
rect 587618 401818 587800 402054
rect 587200 401734 587800 401818
rect 587200 401498 587382 401734
rect 587618 401498 587800 401734
rect 587200 366054 587800 401498
rect 587200 365818 587382 366054
rect 587618 365818 587800 366054
rect 587200 365734 587800 365818
rect 587200 365498 587382 365734
rect 587618 365498 587800 365734
rect 587200 330054 587800 365498
rect 587200 329818 587382 330054
rect 587618 329818 587800 330054
rect 587200 329734 587800 329818
rect 587200 329498 587382 329734
rect 587618 329498 587800 329734
rect 587200 294054 587800 329498
rect 587200 293818 587382 294054
rect 587618 293818 587800 294054
rect 587200 293734 587800 293818
rect 587200 293498 587382 293734
rect 587618 293498 587800 293734
rect 587200 258054 587800 293498
rect 587200 257818 587382 258054
rect 587618 257818 587800 258054
rect 587200 257734 587800 257818
rect 587200 257498 587382 257734
rect 587618 257498 587800 257734
rect 587200 222054 587800 257498
rect 587200 221818 587382 222054
rect 587618 221818 587800 222054
rect 587200 221734 587800 221818
rect 587200 221498 587382 221734
rect 587618 221498 587800 221734
rect 587200 186054 587800 221498
rect 587200 185818 587382 186054
rect 587618 185818 587800 186054
rect 587200 185734 587800 185818
rect 587200 185498 587382 185734
rect 587618 185498 587800 185734
rect 587200 150054 587800 185498
rect 587200 149818 587382 150054
rect 587618 149818 587800 150054
rect 587200 149734 587800 149818
rect 587200 149498 587382 149734
rect 587618 149498 587800 149734
rect 587200 114054 587800 149498
rect 587200 113818 587382 114054
rect 587618 113818 587800 114054
rect 587200 113734 587800 113818
rect 587200 113498 587382 113734
rect 587618 113498 587800 113734
rect 587200 78054 587800 113498
rect 587200 77818 587382 78054
rect 587618 77818 587800 78054
rect 587200 77734 587800 77818
rect 587200 77498 587382 77734
rect 587618 77498 587800 77734
rect 587200 42054 587800 77498
rect 587200 41818 587382 42054
rect 587618 41818 587800 42054
rect 587200 41734 587800 41818
rect 587200 41498 587382 41734
rect 587618 41498 587800 41734
rect 587200 6054 587800 41498
rect 587200 5818 587382 6054
rect 587618 5818 587800 6054
rect 587200 5734 587800 5818
rect 587200 5498 587382 5734
rect 587618 5498 587800 5734
rect 580404 -2462 580586 -2226
rect 580822 -2462 581004 -2226
rect 580404 -2546 581004 -2462
rect 580404 -2782 580586 -2546
rect 580822 -2782 581004 -2546
rect 580404 -3744 581004 -2782
rect 587200 -2226 587800 5498
rect 587200 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect 587200 -2546 587800 -2462
rect 587200 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect 587200 -2804 587800 -2782
rect 588140 672054 588740 707102
rect 588140 671818 588322 672054
rect 588558 671818 588740 672054
rect 588140 671734 588740 671818
rect 588140 671498 588322 671734
rect 588558 671498 588740 671734
rect 588140 636054 588740 671498
rect 588140 635818 588322 636054
rect 588558 635818 588740 636054
rect 588140 635734 588740 635818
rect 588140 635498 588322 635734
rect 588558 635498 588740 635734
rect 588140 600054 588740 635498
rect 588140 599818 588322 600054
rect 588558 599818 588740 600054
rect 588140 599734 588740 599818
rect 588140 599498 588322 599734
rect 588558 599498 588740 599734
rect 588140 564054 588740 599498
rect 588140 563818 588322 564054
rect 588558 563818 588740 564054
rect 588140 563734 588740 563818
rect 588140 563498 588322 563734
rect 588558 563498 588740 563734
rect 588140 528054 588740 563498
rect 588140 527818 588322 528054
rect 588558 527818 588740 528054
rect 588140 527734 588740 527818
rect 588140 527498 588322 527734
rect 588558 527498 588740 527734
rect 588140 492054 588740 527498
rect 588140 491818 588322 492054
rect 588558 491818 588740 492054
rect 588140 491734 588740 491818
rect 588140 491498 588322 491734
rect 588558 491498 588740 491734
rect 588140 456054 588740 491498
rect 588140 455818 588322 456054
rect 588558 455818 588740 456054
rect 588140 455734 588740 455818
rect 588140 455498 588322 455734
rect 588558 455498 588740 455734
rect 588140 420054 588740 455498
rect 588140 419818 588322 420054
rect 588558 419818 588740 420054
rect 588140 419734 588740 419818
rect 588140 419498 588322 419734
rect 588558 419498 588740 419734
rect 588140 384054 588740 419498
rect 588140 383818 588322 384054
rect 588558 383818 588740 384054
rect 588140 383734 588740 383818
rect 588140 383498 588322 383734
rect 588558 383498 588740 383734
rect 588140 348054 588740 383498
rect 588140 347818 588322 348054
rect 588558 347818 588740 348054
rect 588140 347734 588740 347818
rect 588140 347498 588322 347734
rect 588558 347498 588740 347734
rect 588140 312054 588740 347498
rect 588140 311818 588322 312054
rect 588558 311818 588740 312054
rect 588140 311734 588740 311818
rect 588140 311498 588322 311734
rect 588558 311498 588740 311734
rect 588140 276054 588740 311498
rect 588140 275818 588322 276054
rect 588558 275818 588740 276054
rect 588140 275734 588740 275818
rect 588140 275498 588322 275734
rect 588558 275498 588740 275734
rect 588140 240054 588740 275498
rect 588140 239818 588322 240054
rect 588558 239818 588740 240054
rect 588140 239734 588740 239818
rect 588140 239498 588322 239734
rect 588558 239498 588740 239734
rect 588140 204054 588740 239498
rect 588140 203818 588322 204054
rect 588558 203818 588740 204054
rect 588140 203734 588740 203818
rect 588140 203498 588322 203734
rect 588558 203498 588740 203734
rect 588140 168054 588740 203498
rect 588140 167818 588322 168054
rect 588558 167818 588740 168054
rect 588140 167734 588740 167818
rect 588140 167498 588322 167734
rect 588558 167498 588740 167734
rect 588140 132054 588740 167498
rect 588140 131818 588322 132054
rect 588558 131818 588740 132054
rect 588140 131734 588740 131818
rect 588140 131498 588322 131734
rect 588558 131498 588740 131734
rect 588140 96054 588740 131498
rect 588140 95818 588322 96054
rect 588558 95818 588740 96054
rect 588140 95734 588740 95818
rect 588140 95498 588322 95734
rect 588558 95498 588740 95734
rect 588140 60054 588740 95498
rect 588140 59818 588322 60054
rect 588558 59818 588740 60054
rect 588140 59734 588740 59818
rect 588140 59498 588322 59734
rect 588558 59498 588740 59734
rect 588140 24054 588740 59498
rect 588140 23818 588322 24054
rect 588558 23818 588740 24054
rect 588140 23734 588740 23818
rect 588140 23498 588322 23734
rect 588558 23498 588740 23734
rect 588140 -3166 588740 23498
rect 588140 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect 588140 -3486 588740 -3402
rect 588140 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect 588140 -3744 588740 -3722
rect 589080 693654 589680 708042
rect 589080 693418 589262 693654
rect 589498 693418 589680 693654
rect 589080 693334 589680 693418
rect 589080 693098 589262 693334
rect 589498 693098 589680 693334
rect 589080 657654 589680 693098
rect 589080 657418 589262 657654
rect 589498 657418 589680 657654
rect 589080 657334 589680 657418
rect 589080 657098 589262 657334
rect 589498 657098 589680 657334
rect 589080 621654 589680 657098
rect 589080 621418 589262 621654
rect 589498 621418 589680 621654
rect 589080 621334 589680 621418
rect 589080 621098 589262 621334
rect 589498 621098 589680 621334
rect 589080 585654 589680 621098
rect 589080 585418 589262 585654
rect 589498 585418 589680 585654
rect 589080 585334 589680 585418
rect 589080 585098 589262 585334
rect 589498 585098 589680 585334
rect 589080 549654 589680 585098
rect 589080 549418 589262 549654
rect 589498 549418 589680 549654
rect 589080 549334 589680 549418
rect 589080 549098 589262 549334
rect 589498 549098 589680 549334
rect 589080 513654 589680 549098
rect 589080 513418 589262 513654
rect 589498 513418 589680 513654
rect 589080 513334 589680 513418
rect 589080 513098 589262 513334
rect 589498 513098 589680 513334
rect 589080 477654 589680 513098
rect 589080 477418 589262 477654
rect 589498 477418 589680 477654
rect 589080 477334 589680 477418
rect 589080 477098 589262 477334
rect 589498 477098 589680 477334
rect 589080 441654 589680 477098
rect 589080 441418 589262 441654
rect 589498 441418 589680 441654
rect 589080 441334 589680 441418
rect 589080 441098 589262 441334
rect 589498 441098 589680 441334
rect 589080 405654 589680 441098
rect 589080 405418 589262 405654
rect 589498 405418 589680 405654
rect 589080 405334 589680 405418
rect 589080 405098 589262 405334
rect 589498 405098 589680 405334
rect 589080 369654 589680 405098
rect 589080 369418 589262 369654
rect 589498 369418 589680 369654
rect 589080 369334 589680 369418
rect 589080 369098 589262 369334
rect 589498 369098 589680 369334
rect 589080 333654 589680 369098
rect 589080 333418 589262 333654
rect 589498 333418 589680 333654
rect 589080 333334 589680 333418
rect 589080 333098 589262 333334
rect 589498 333098 589680 333334
rect 589080 297654 589680 333098
rect 589080 297418 589262 297654
rect 589498 297418 589680 297654
rect 589080 297334 589680 297418
rect 589080 297098 589262 297334
rect 589498 297098 589680 297334
rect 589080 261654 589680 297098
rect 589080 261418 589262 261654
rect 589498 261418 589680 261654
rect 589080 261334 589680 261418
rect 589080 261098 589262 261334
rect 589498 261098 589680 261334
rect 589080 225654 589680 261098
rect 589080 225418 589262 225654
rect 589498 225418 589680 225654
rect 589080 225334 589680 225418
rect 589080 225098 589262 225334
rect 589498 225098 589680 225334
rect 589080 189654 589680 225098
rect 589080 189418 589262 189654
rect 589498 189418 589680 189654
rect 589080 189334 589680 189418
rect 589080 189098 589262 189334
rect 589498 189098 589680 189334
rect 589080 153654 589680 189098
rect 589080 153418 589262 153654
rect 589498 153418 589680 153654
rect 589080 153334 589680 153418
rect 589080 153098 589262 153334
rect 589498 153098 589680 153334
rect 589080 117654 589680 153098
rect 589080 117418 589262 117654
rect 589498 117418 589680 117654
rect 589080 117334 589680 117418
rect 589080 117098 589262 117334
rect 589498 117098 589680 117334
rect 589080 81654 589680 117098
rect 589080 81418 589262 81654
rect 589498 81418 589680 81654
rect 589080 81334 589680 81418
rect 589080 81098 589262 81334
rect 589498 81098 589680 81334
rect 589080 45654 589680 81098
rect 589080 45418 589262 45654
rect 589498 45418 589680 45654
rect 589080 45334 589680 45418
rect 589080 45098 589262 45334
rect 589498 45098 589680 45334
rect 589080 9654 589680 45098
rect 589080 9418 589262 9654
rect 589498 9418 589680 9654
rect 589080 9334 589680 9418
rect 589080 9098 589262 9334
rect 589498 9098 589680 9334
rect 589080 -4106 589680 9098
rect 589080 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect 589080 -4426 589680 -4342
rect 589080 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect 589080 -4684 589680 -4662
rect 590020 675654 590620 708982
rect 590020 675418 590202 675654
rect 590438 675418 590620 675654
rect 590020 675334 590620 675418
rect 590020 675098 590202 675334
rect 590438 675098 590620 675334
rect 590020 639654 590620 675098
rect 590020 639418 590202 639654
rect 590438 639418 590620 639654
rect 590020 639334 590620 639418
rect 590020 639098 590202 639334
rect 590438 639098 590620 639334
rect 590020 603654 590620 639098
rect 590020 603418 590202 603654
rect 590438 603418 590620 603654
rect 590020 603334 590620 603418
rect 590020 603098 590202 603334
rect 590438 603098 590620 603334
rect 590020 567654 590620 603098
rect 590020 567418 590202 567654
rect 590438 567418 590620 567654
rect 590020 567334 590620 567418
rect 590020 567098 590202 567334
rect 590438 567098 590620 567334
rect 590020 531654 590620 567098
rect 590020 531418 590202 531654
rect 590438 531418 590620 531654
rect 590020 531334 590620 531418
rect 590020 531098 590202 531334
rect 590438 531098 590620 531334
rect 590020 495654 590620 531098
rect 590020 495418 590202 495654
rect 590438 495418 590620 495654
rect 590020 495334 590620 495418
rect 590020 495098 590202 495334
rect 590438 495098 590620 495334
rect 590020 459654 590620 495098
rect 590020 459418 590202 459654
rect 590438 459418 590620 459654
rect 590020 459334 590620 459418
rect 590020 459098 590202 459334
rect 590438 459098 590620 459334
rect 590020 423654 590620 459098
rect 590020 423418 590202 423654
rect 590438 423418 590620 423654
rect 590020 423334 590620 423418
rect 590020 423098 590202 423334
rect 590438 423098 590620 423334
rect 590020 387654 590620 423098
rect 590020 387418 590202 387654
rect 590438 387418 590620 387654
rect 590020 387334 590620 387418
rect 590020 387098 590202 387334
rect 590438 387098 590620 387334
rect 590020 351654 590620 387098
rect 590020 351418 590202 351654
rect 590438 351418 590620 351654
rect 590020 351334 590620 351418
rect 590020 351098 590202 351334
rect 590438 351098 590620 351334
rect 590020 315654 590620 351098
rect 590020 315418 590202 315654
rect 590438 315418 590620 315654
rect 590020 315334 590620 315418
rect 590020 315098 590202 315334
rect 590438 315098 590620 315334
rect 590020 279654 590620 315098
rect 590020 279418 590202 279654
rect 590438 279418 590620 279654
rect 590020 279334 590620 279418
rect 590020 279098 590202 279334
rect 590438 279098 590620 279334
rect 590020 243654 590620 279098
rect 590020 243418 590202 243654
rect 590438 243418 590620 243654
rect 590020 243334 590620 243418
rect 590020 243098 590202 243334
rect 590438 243098 590620 243334
rect 590020 207654 590620 243098
rect 590020 207418 590202 207654
rect 590438 207418 590620 207654
rect 590020 207334 590620 207418
rect 590020 207098 590202 207334
rect 590438 207098 590620 207334
rect 590020 171654 590620 207098
rect 590020 171418 590202 171654
rect 590438 171418 590620 171654
rect 590020 171334 590620 171418
rect 590020 171098 590202 171334
rect 590438 171098 590620 171334
rect 590020 135654 590620 171098
rect 590020 135418 590202 135654
rect 590438 135418 590620 135654
rect 590020 135334 590620 135418
rect 590020 135098 590202 135334
rect 590438 135098 590620 135334
rect 590020 99654 590620 135098
rect 590020 99418 590202 99654
rect 590438 99418 590620 99654
rect 590020 99334 590620 99418
rect 590020 99098 590202 99334
rect 590438 99098 590620 99334
rect 590020 63654 590620 99098
rect 590020 63418 590202 63654
rect 590438 63418 590620 63654
rect 590020 63334 590620 63418
rect 590020 63098 590202 63334
rect 590438 63098 590620 63334
rect 590020 27654 590620 63098
rect 590020 27418 590202 27654
rect 590438 27418 590620 27654
rect 590020 27334 590620 27418
rect 590020 27098 590202 27334
rect 590438 27098 590620 27334
rect 590020 -5046 590620 27098
rect 590020 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect 590020 -5366 590620 -5282
rect 590020 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect 590020 -5624 590620 -5602
rect 590960 697254 591560 709922
rect 590960 697018 591142 697254
rect 591378 697018 591560 697254
rect 590960 696934 591560 697018
rect 590960 696698 591142 696934
rect 591378 696698 591560 696934
rect 590960 661254 591560 696698
rect 590960 661018 591142 661254
rect 591378 661018 591560 661254
rect 590960 660934 591560 661018
rect 590960 660698 591142 660934
rect 591378 660698 591560 660934
rect 590960 625254 591560 660698
rect 590960 625018 591142 625254
rect 591378 625018 591560 625254
rect 590960 624934 591560 625018
rect 590960 624698 591142 624934
rect 591378 624698 591560 624934
rect 590960 589254 591560 624698
rect 590960 589018 591142 589254
rect 591378 589018 591560 589254
rect 590960 588934 591560 589018
rect 590960 588698 591142 588934
rect 591378 588698 591560 588934
rect 590960 553254 591560 588698
rect 590960 553018 591142 553254
rect 591378 553018 591560 553254
rect 590960 552934 591560 553018
rect 590960 552698 591142 552934
rect 591378 552698 591560 552934
rect 590960 517254 591560 552698
rect 590960 517018 591142 517254
rect 591378 517018 591560 517254
rect 590960 516934 591560 517018
rect 590960 516698 591142 516934
rect 591378 516698 591560 516934
rect 590960 481254 591560 516698
rect 590960 481018 591142 481254
rect 591378 481018 591560 481254
rect 590960 480934 591560 481018
rect 590960 480698 591142 480934
rect 591378 480698 591560 480934
rect 590960 445254 591560 480698
rect 590960 445018 591142 445254
rect 591378 445018 591560 445254
rect 590960 444934 591560 445018
rect 590960 444698 591142 444934
rect 591378 444698 591560 444934
rect 590960 409254 591560 444698
rect 590960 409018 591142 409254
rect 591378 409018 591560 409254
rect 590960 408934 591560 409018
rect 590960 408698 591142 408934
rect 591378 408698 591560 408934
rect 590960 373254 591560 408698
rect 590960 373018 591142 373254
rect 591378 373018 591560 373254
rect 590960 372934 591560 373018
rect 590960 372698 591142 372934
rect 591378 372698 591560 372934
rect 590960 337254 591560 372698
rect 590960 337018 591142 337254
rect 591378 337018 591560 337254
rect 590960 336934 591560 337018
rect 590960 336698 591142 336934
rect 591378 336698 591560 336934
rect 590960 301254 591560 336698
rect 590960 301018 591142 301254
rect 591378 301018 591560 301254
rect 590960 300934 591560 301018
rect 590960 300698 591142 300934
rect 591378 300698 591560 300934
rect 590960 265254 591560 300698
rect 590960 265018 591142 265254
rect 591378 265018 591560 265254
rect 590960 264934 591560 265018
rect 590960 264698 591142 264934
rect 591378 264698 591560 264934
rect 590960 229254 591560 264698
rect 590960 229018 591142 229254
rect 591378 229018 591560 229254
rect 590960 228934 591560 229018
rect 590960 228698 591142 228934
rect 591378 228698 591560 228934
rect 590960 193254 591560 228698
rect 590960 193018 591142 193254
rect 591378 193018 591560 193254
rect 590960 192934 591560 193018
rect 590960 192698 591142 192934
rect 591378 192698 591560 192934
rect 590960 157254 591560 192698
rect 590960 157018 591142 157254
rect 591378 157018 591560 157254
rect 590960 156934 591560 157018
rect 590960 156698 591142 156934
rect 591378 156698 591560 156934
rect 590960 121254 591560 156698
rect 590960 121018 591142 121254
rect 591378 121018 591560 121254
rect 590960 120934 591560 121018
rect 590960 120698 591142 120934
rect 591378 120698 591560 120934
rect 590960 85254 591560 120698
rect 590960 85018 591142 85254
rect 591378 85018 591560 85254
rect 590960 84934 591560 85018
rect 590960 84698 591142 84934
rect 591378 84698 591560 84934
rect 590960 49254 591560 84698
rect 590960 49018 591142 49254
rect 591378 49018 591560 49254
rect 590960 48934 591560 49018
rect 590960 48698 591142 48934
rect 591378 48698 591560 48934
rect 590960 13254 591560 48698
rect 590960 13018 591142 13254
rect 591378 13018 591560 13254
rect 590960 12934 591560 13018
rect 590960 12698 591142 12934
rect 591378 12698 591560 12934
rect 590960 -5986 591560 12698
rect 590960 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect 590960 -6306 591560 -6222
rect 590960 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect 590960 -6564 591560 -6542
rect 591900 679254 592500 710862
rect 591900 679018 592082 679254
rect 592318 679018 592500 679254
rect 591900 678934 592500 679018
rect 591900 678698 592082 678934
rect 592318 678698 592500 678934
rect 591900 643254 592500 678698
rect 591900 643018 592082 643254
rect 592318 643018 592500 643254
rect 591900 642934 592500 643018
rect 591900 642698 592082 642934
rect 592318 642698 592500 642934
rect 591900 607254 592500 642698
rect 591900 607018 592082 607254
rect 592318 607018 592500 607254
rect 591900 606934 592500 607018
rect 591900 606698 592082 606934
rect 592318 606698 592500 606934
rect 591900 571254 592500 606698
rect 591900 571018 592082 571254
rect 592318 571018 592500 571254
rect 591900 570934 592500 571018
rect 591900 570698 592082 570934
rect 592318 570698 592500 570934
rect 591900 535254 592500 570698
rect 591900 535018 592082 535254
rect 592318 535018 592500 535254
rect 591900 534934 592500 535018
rect 591900 534698 592082 534934
rect 592318 534698 592500 534934
rect 591900 499254 592500 534698
rect 591900 499018 592082 499254
rect 592318 499018 592500 499254
rect 591900 498934 592500 499018
rect 591900 498698 592082 498934
rect 592318 498698 592500 498934
rect 591900 463254 592500 498698
rect 591900 463018 592082 463254
rect 592318 463018 592500 463254
rect 591900 462934 592500 463018
rect 591900 462698 592082 462934
rect 592318 462698 592500 462934
rect 591900 427254 592500 462698
rect 591900 427018 592082 427254
rect 592318 427018 592500 427254
rect 591900 426934 592500 427018
rect 591900 426698 592082 426934
rect 592318 426698 592500 426934
rect 591900 391254 592500 426698
rect 591900 391018 592082 391254
rect 592318 391018 592500 391254
rect 591900 390934 592500 391018
rect 591900 390698 592082 390934
rect 592318 390698 592500 390934
rect 591900 355254 592500 390698
rect 591900 355018 592082 355254
rect 592318 355018 592500 355254
rect 591900 354934 592500 355018
rect 591900 354698 592082 354934
rect 592318 354698 592500 354934
rect 591900 319254 592500 354698
rect 591900 319018 592082 319254
rect 592318 319018 592500 319254
rect 591900 318934 592500 319018
rect 591900 318698 592082 318934
rect 592318 318698 592500 318934
rect 591900 283254 592500 318698
rect 591900 283018 592082 283254
rect 592318 283018 592500 283254
rect 591900 282934 592500 283018
rect 591900 282698 592082 282934
rect 592318 282698 592500 282934
rect 591900 247254 592500 282698
rect 591900 247018 592082 247254
rect 592318 247018 592500 247254
rect 591900 246934 592500 247018
rect 591900 246698 592082 246934
rect 592318 246698 592500 246934
rect 591900 211254 592500 246698
rect 591900 211018 592082 211254
rect 592318 211018 592500 211254
rect 591900 210934 592500 211018
rect 591900 210698 592082 210934
rect 592318 210698 592500 210934
rect 591900 175254 592500 210698
rect 591900 175018 592082 175254
rect 592318 175018 592500 175254
rect 591900 174934 592500 175018
rect 591900 174698 592082 174934
rect 592318 174698 592500 174934
rect 591900 139254 592500 174698
rect 591900 139018 592082 139254
rect 592318 139018 592500 139254
rect 591900 138934 592500 139018
rect 591900 138698 592082 138934
rect 592318 138698 592500 138934
rect 591900 103254 592500 138698
rect 591900 103018 592082 103254
rect 592318 103018 592500 103254
rect 591900 102934 592500 103018
rect 591900 102698 592082 102934
rect 592318 102698 592500 102934
rect 591900 67254 592500 102698
rect 591900 67018 592082 67254
rect 592318 67018 592500 67254
rect 591900 66934 592500 67018
rect 591900 66698 592082 66934
rect 592318 66698 592500 66934
rect 591900 31254 592500 66698
rect 591900 31018 592082 31254
rect 592318 31018 592500 31254
rect 591900 30934 592500 31018
rect 591900 30698 592082 30934
rect 592318 30698 592500 30934
rect 569604 -7162 569786 -6926
rect 570022 -7162 570204 -6926
rect 569604 -7246 570204 -7162
rect 569604 -7482 569786 -7246
rect 570022 -7482 570204 -7246
rect 569604 -7504 570204 -7482
rect 591900 -6926 592500 30698
rect 591900 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect 591900 -7246 592500 -7162
rect 591900 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect 591900 -7504 592500 -7482
<< via4 >>
rect -8394 711182 -8158 711418
rect -8394 710862 -8158 711098
rect -8394 679018 -8158 679254
rect -8394 678698 -8158 678934
rect -8394 643018 -8158 643254
rect -8394 642698 -8158 642934
rect -8394 607018 -8158 607254
rect -8394 606698 -8158 606934
rect -8394 571018 -8158 571254
rect -8394 570698 -8158 570934
rect -8394 535018 -8158 535254
rect -8394 534698 -8158 534934
rect -8394 499018 -8158 499254
rect -8394 498698 -8158 498934
rect -8394 463018 -8158 463254
rect -8394 462698 -8158 462934
rect -8394 427018 -8158 427254
rect -8394 426698 -8158 426934
rect -8394 391018 -8158 391254
rect -8394 390698 -8158 390934
rect -8394 355018 -8158 355254
rect -8394 354698 -8158 354934
rect -8394 319018 -8158 319254
rect -8394 318698 -8158 318934
rect -8394 283018 -8158 283254
rect -8394 282698 -8158 282934
rect -8394 247018 -8158 247254
rect -8394 246698 -8158 246934
rect -8394 211018 -8158 211254
rect -8394 210698 -8158 210934
rect -8394 175018 -8158 175254
rect -8394 174698 -8158 174934
rect -8394 139018 -8158 139254
rect -8394 138698 -8158 138934
rect -8394 103018 -8158 103254
rect -8394 102698 -8158 102934
rect -8394 67018 -8158 67254
rect -8394 66698 -8158 66934
rect -8394 31018 -8158 31254
rect -8394 30698 -8158 30934
rect -7454 710242 -7218 710478
rect -7454 709922 -7218 710158
rect 11786 710242 12022 710478
rect 11786 709922 12022 710158
rect -7454 697018 -7218 697254
rect -7454 696698 -7218 696934
rect -7454 661018 -7218 661254
rect -7454 660698 -7218 660934
rect -7454 625018 -7218 625254
rect -7454 624698 -7218 624934
rect -7454 589018 -7218 589254
rect -7454 588698 -7218 588934
rect -7454 553018 -7218 553254
rect -7454 552698 -7218 552934
rect -7454 517018 -7218 517254
rect -7454 516698 -7218 516934
rect -7454 481018 -7218 481254
rect -7454 480698 -7218 480934
rect -7454 445018 -7218 445254
rect -7454 444698 -7218 444934
rect -7454 409018 -7218 409254
rect -7454 408698 -7218 408934
rect -7454 373018 -7218 373254
rect -7454 372698 -7218 372934
rect -7454 337018 -7218 337254
rect -7454 336698 -7218 336934
rect -7454 301018 -7218 301254
rect -7454 300698 -7218 300934
rect -7454 265018 -7218 265254
rect -7454 264698 -7218 264934
rect -7454 229018 -7218 229254
rect -7454 228698 -7218 228934
rect -7454 193018 -7218 193254
rect -7454 192698 -7218 192934
rect -7454 157018 -7218 157254
rect -7454 156698 -7218 156934
rect -7454 121018 -7218 121254
rect -7454 120698 -7218 120934
rect -7454 85018 -7218 85254
rect -7454 84698 -7218 84934
rect -7454 49018 -7218 49254
rect -7454 48698 -7218 48934
rect -7454 13018 -7218 13254
rect -7454 12698 -7218 12934
rect -6514 709302 -6278 709538
rect -6514 708982 -6278 709218
rect -6514 675418 -6278 675654
rect -6514 675098 -6278 675334
rect -6514 639418 -6278 639654
rect -6514 639098 -6278 639334
rect -6514 603418 -6278 603654
rect -6514 603098 -6278 603334
rect -6514 567418 -6278 567654
rect -6514 567098 -6278 567334
rect -6514 531418 -6278 531654
rect -6514 531098 -6278 531334
rect -6514 495418 -6278 495654
rect -6514 495098 -6278 495334
rect -6514 459418 -6278 459654
rect -6514 459098 -6278 459334
rect -6514 423418 -6278 423654
rect -6514 423098 -6278 423334
rect -6514 387418 -6278 387654
rect -6514 387098 -6278 387334
rect -6514 351418 -6278 351654
rect -6514 351098 -6278 351334
rect -6514 315418 -6278 315654
rect -6514 315098 -6278 315334
rect -6514 279418 -6278 279654
rect -6514 279098 -6278 279334
rect -6514 243418 -6278 243654
rect -6514 243098 -6278 243334
rect -6514 207418 -6278 207654
rect -6514 207098 -6278 207334
rect -6514 171418 -6278 171654
rect -6514 171098 -6278 171334
rect -6514 135418 -6278 135654
rect -6514 135098 -6278 135334
rect -6514 99418 -6278 99654
rect -6514 99098 -6278 99334
rect -6514 63418 -6278 63654
rect -6514 63098 -6278 63334
rect -6514 27418 -6278 27654
rect -6514 27098 -6278 27334
rect -5574 708362 -5338 708598
rect -5574 708042 -5338 708278
rect 8186 708362 8422 708598
rect 8186 708042 8422 708278
rect -5574 693418 -5338 693654
rect -5574 693098 -5338 693334
rect -5574 657418 -5338 657654
rect -5574 657098 -5338 657334
rect -5574 621418 -5338 621654
rect -5574 621098 -5338 621334
rect -5574 585418 -5338 585654
rect -5574 585098 -5338 585334
rect -5574 549418 -5338 549654
rect -5574 549098 -5338 549334
rect -5574 513418 -5338 513654
rect -5574 513098 -5338 513334
rect -5574 477418 -5338 477654
rect -5574 477098 -5338 477334
rect -5574 441418 -5338 441654
rect -5574 441098 -5338 441334
rect -5574 405418 -5338 405654
rect -5574 405098 -5338 405334
rect -5574 369418 -5338 369654
rect -5574 369098 -5338 369334
rect -5574 333418 -5338 333654
rect -5574 333098 -5338 333334
rect -5574 297418 -5338 297654
rect -5574 297098 -5338 297334
rect -5574 261418 -5338 261654
rect -5574 261098 -5338 261334
rect -5574 225418 -5338 225654
rect -5574 225098 -5338 225334
rect -5574 189418 -5338 189654
rect -5574 189098 -5338 189334
rect -5574 153418 -5338 153654
rect -5574 153098 -5338 153334
rect -5574 117418 -5338 117654
rect -5574 117098 -5338 117334
rect -5574 81418 -5338 81654
rect -5574 81098 -5338 81334
rect -5574 45418 -5338 45654
rect -5574 45098 -5338 45334
rect -5574 9418 -5338 9654
rect -5574 9098 -5338 9334
rect -4634 707422 -4398 707658
rect -4634 707102 -4398 707338
rect -4634 671818 -4398 672054
rect -4634 671498 -4398 671734
rect -4634 635818 -4398 636054
rect -4634 635498 -4398 635734
rect -4634 599818 -4398 600054
rect -4634 599498 -4398 599734
rect -4634 563818 -4398 564054
rect -4634 563498 -4398 563734
rect -4634 527818 -4398 528054
rect -4634 527498 -4398 527734
rect -4634 491818 -4398 492054
rect -4634 491498 -4398 491734
rect -4634 455818 -4398 456054
rect -4634 455498 -4398 455734
rect -4634 419818 -4398 420054
rect -4634 419498 -4398 419734
rect -4634 383818 -4398 384054
rect -4634 383498 -4398 383734
rect -4634 347818 -4398 348054
rect -4634 347498 -4398 347734
rect -4634 311818 -4398 312054
rect -4634 311498 -4398 311734
rect -4634 275818 -4398 276054
rect -4634 275498 -4398 275734
rect -4634 239818 -4398 240054
rect -4634 239498 -4398 239734
rect -4634 203818 -4398 204054
rect -4634 203498 -4398 203734
rect -4634 167818 -4398 168054
rect -4634 167498 -4398 167734
rect -4634 131818 -4398 132054
rect -4634 131498 -4398 131734
rect -4634 95818 -4398 96054
rect -4634 95498 -4398 95734
rect -4634 59818 -4398 60054
rect -4634 59498 -4398 59734
rect -4634 23818 -4398 24054
rect -4634 23498 -4398 23734
rect -3694 706482 -3458 706718
rect -3694 706162 -3458 706398
rect 4586 706482 4822 706718
rect 4586 706162 4822 706398
rect -3694 689818 -3458 690054
rect -3694 689498 -3458 689734
rect -3694 653818 -3458 654054
rect -3694 653498 -3458 653734
rect -3694 617818 -3458 618054
rect -3694 617498 -3458 617734
rect -3694 581818 -3458 582054
rect -3694 581498 -3458 581734
rect -3694 545818 -3458 546054
rect -3694 545498 -3458 545734
rect -3694 509818 -3458 510054
rect -3694 509498 -3458 509734
rect -3694 473818 -3458 474054
rect -3694 473498 -3458 473734
rect -3694 437818 -3458 438054
rect -3694 437498 -3458 437734
rect -3694 401818 -3458 402054
rect -3694 401498 -3458 401734
rect -3694 365818 -3458 366054
rect -3694 365498 -3458 365734
rect -3694 329818 -3458 330054
rect -3694 329498 -3458 329734
rect -3694 293818 -3458 294054
rect -3694 293498 -3458 293734
rect -3694 257818 -3458 258054
rect -3694 257498 -3458 257734
rect -3694 221818 -3458 222054
rect -3694 221498 -3458 221734
rect -3694 185818 -3458 186054
rect -3694 185498 -3458 185734
rect -3694 149818 -3458 150054
rect -3694 149498 -3458 149734
rect -3694 113818 -3458 114054
rect -3694 113498 -3458 113734
rect -3694 77818 -3458 78054
rect -3694 77498 -3458 77734
rect -3694 41818 -3458 42054
rect -3694 41498 -3458 41734
rect -3694 5818 -3458 6054
rect -3694 5498 -3458 5734
rect -2754 705542 -2518 705778
rect -2754 705222 -2518 705458
rect -2754 668218 -2518 668454
rect -2754 667898 -2518 668134
rect -2754 632218 -2518 632454
rect -2754 631898 -2518 632134
rect -2754 596218 -2518 596454
rect -2754 595898 -2518 596134
rect -2754 560218 -2518 560454
rect -2754 559898 -2518 560134
rect -2754 524218 -2518 524454
rect -2754 523898 -2518 524134
rect -2754 488218 -2518 488454
rect -2754 487898 -2518 488134
rect -2754 452218 -2518 452454
rect -2754 451898 -2518 452134
rect -2754 416218 -2518 416454
rect -2754 415898 -2518 416134
rect -2754 380218 -2518 380454
rect -2754 379898 -2518 380134
rect -2754 344218 -2518 344454
rect -2754 343898 -2518 344134
rect -2754 308218 -2518 308454
rect -2754 307898 -2518 308134
rect -2754 272218 -2518 272454
rect -2754 271898 -2518 272134
rect -2754 236218 -2518 236454
rect -2754 235898 -2518 236134
rect -2754 200218 -2518 200454
rect -2754 199898 -2518 200134
rect -2754 164218 -2518 164454
rect -2754 163898 -2518 164134
rect -2754 128218 -2518 128454
rect -2754 127898 -2518 128134
rect -2754 92218 -2518 92454
rect -2754 91898 -2518 92134
rect -2754 56218 -2518 56454
rect -2754 55898 -2518 56134
rect -2754 20218 -2518 20454
rect -2754 19898 -2518 20134
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect -1814 686218 -1578 686454
rect -1814 685898 -1578 686134
rect -1814 650218 -1578 650454
rect -1814 649898 -1578 650134
rect -1814 614218 -1578 614454
rect -1814 613898 -1578 614134
rect -1814 578218 -1578 578454
rect -1814 577898 -1578 578134
rect -1814 542218 -1578 542454
rect -1814 541898 -1578 542134
rect -1814 506218 -1578 506454
rect -1814 505898 -1578 506134
rect -1814 470218 -1578 470454
rect -1814 469898 -1578 470134
rect -1814 434218 -1578 434454
rect -1814 433898 -1578 434134
rect -1814 398218 -1578 398454
rect -1814 397898 -1578 398134
rect -1814 362218 -1578 362454
rect -1814 361898 -1578 362134
rect -1814 326218 -1578 326454
rect -1814 325898 -1578 326134
rect -1814 290218 -1578 290454
rect -1814 289898 -1578 290134
rect -1814 254218 -1578 254454
rect -1814 253898 -1578 254134
rect -1814 218218 -1578 218454
rect -1814 217898 -1578 218134
rect -1814 182218 -1578 182454
rect -1814 181898 -1578 182134
rect -1814 146218 -1578 146454
rect -1814 145898 -1578 146134
rect -1814 110218 -1578 110454
rect -1814 109898 -1578 110134
rect -1814 74218 -1578 74454
rect -1814 73898 -1578 74134
rect -1814 38218 -1578 38454
rect -1814 37898 -1578 38134
rect -1814 2218 -1578 2454
rect -1814 1898 -1578 2134
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 986 704602 1222 704838
rect 986 704282 1222 704518
rect 986 686218 1222 686454
rect 986 685898 1222 686134
rect 986 650218 1222 650454
rect 986 649898 1222 650134
rect 986 614218 1222 614454
rect 986 613898 1222 614134
rect 986 578218 1222 578454
rect 986 577898 1222 578134
rect 986 542218 1222 542454
rect 986 541898 1222 542134
rect 986 506218 1222 506454
rect 986 505898 1222 506134
rect 986 470218 1222 470454
rect 986 469898 1222 470134
rect 986 434218 1222 434454
rect 986 433898 1222 434134
rect 986 398218 1222 398454
rect 986 397898 1222 398134
rect 986 362218 1222 362454
rect 986 361898 1222 362134
rect 986 326218 1222 326454
rect 986 325898 1222 326134
rect 986 290218 1222 290454
rect 986 289898 1222 290134
rect 986 254218 1222 254454
rect 986 253898 1222 254134
rect 986 218218 1222 218454
rect 986 217898 1222 218134
rect 986 182218 1222 182454
rect 986 181898 1222 182134
rect 986 146218 1222 146454
rect 986 145898 1222 146134
rect 986 110218 1222 110454
rect 986 109898 1222 110134
rect 986 74218 1222 74454
rect 986 73898 1222 74134
rect 986 38218 1222 38454
rect 986 37898 1222 38134
rect 986 2218 1222 2454
rect 986 1898 1222 2134
rect 986 -582 1222 -346
rect 986 -902 1222 -666
rect -2754 -1522 -2518 -1286
rect -2754 -1842 -2518 -1606
rect 4586 689818 4822 690054
rect 4586 689498 4822 689734
rect 4586 653818 4822 654054
rect 4586 653498 4822 653734
rect 4586 617818 4822 618054
rect 4586 617498 4822 617734
rect 4586 581818 4822 582054
rect 4586 581498 4822 581734
rect 4586 545818 4822 546054
rect 4586 545498 4822 545734
rect 4586 509818 4822 510054
rect 4586 509498 4822 509734
rect 4586 473818 4822 474054
rect 4586 473498 4822 473734
rect 4586 437818 4822 438054
rect 4586 437498 4822 437734
rect 4586 401818 4822 402054
rect 4586 401498 4822 401734
rect 4586 365818 4822 366054
rect 4586 365498 4822 365734
rect 4586 329818 4822 330054
rect 4586 329498 4822 329734
rect 4586 293818 4822 294054
rect 4586 293498 4822 293734
rect 4586 257818 4822 258054
rect 4586 257498 4822 257734
rect 4586 221818 4822 222054
rect 4586 221498 4822 221734
rect 4586 185818 4822 186054
rect 4586 185498 4822 185734
rect 4586 149818 4822 150054
rect 4586 149498 4822 149734
rect 4586 113818 4822 114054
rect 4586 113498 4822 113734
rect 4586 77818 4822 78054
rect 4586 77498 4822 77734
rect 4586 41818 4822 42054
rect 4586 41498 4822 41734
rect 4586 5818 4822 6054
rect 4586 5498 4822 5734
rect -3694 -2462 -3458 -2226
rect -3694 -2782 -3458 -2546
rect 4586 -2462 4822 -2226
rect 4586 -2782 4822 -2546
rect -4634 -3402 -4398 -3166
rect -4634 -3722 -4398 -3486
rect 8186 693418 8422 693654
rect 8186 693098 8422 693334
rect 8186 657418 8422 657654
rect 8186 657098 8422 657334
rect 8186 621418 8422 621654
rect 8186 621098 8422 621334
rect 8186 585418 8422 585654
rect 8186 585098 8422 585334
rect 8186 549418 8422 549654
rect 8186 549098 8422 549334
rect 8186 513418 8422 513654
rect 8186 513098 8422 513334
rect 8186 477418 8422 477654
rect 8186 477098 8422 477334
rect 8186 441418 8422 441654
rect 8186 441098 8422 441334
rect 8186 405418 8422 405654
rect 8186 405098 8422 405334
rect 8186 369418 8422 369654
rect 8186 369098 8422 369334
rect 8186 333418 8422 333654
rect 8186 333098 8422 333334
rect 8186 297418 8422 297654
rect 8186 297098 8422 297334
rect 8186 261418 8422 261654
rect 8186 261098 8422 261334
rect 8186 225418 8422 225654
rect 8186 225098 8422 225334
rect 8186 189418 8422 189654
rect 8186 189098 8422 189334
rect 8186 153418 8422 153654
rect 8186 153098 8422 153334
rect 8186 117418 8422 117654
rect 8186 117098 8422 117334
rect 29786 711182 30022 711418
rect 29786 710862 30022 711098
rect 26186 709302 26422 709538
rect 26186 708982 26422 709218
rect 22586 707422 22822 707658
rect 22586 707102 22822 707338
rect 11786 697018 12022 697254
rect 11786 696698 12022 696934
rect 11786 661018 12022 661254
rect 11786 660698 12022 660934
rect 11786 625018 12022 625254
rect 11786 624698 12022 624934
rect 11786 589018 12022 589254
rect 11786 588698 12022 588934
rect 11786 553018 12022 553254
rect 11786 552698 12022 552934
rect 11786 517018 12022 517254
rect 11786 516698 12022 516934
rect 11786 481018 12022 481254
rect 11786 480698 12022 480934
rect 11786 445018 12022 445254
rect 11786 444698 12022 444934
rect 11786 409018 12022 409254
rect 11786 408698 12022 408934
rect 11786 373018 12022 373254
rect 11786 372698 12022 372934
rect 11786 337018 12022 337254
rect 11786 336698 12022 336934
rect 11786 301018 12022 301254
rect 11786 300698 12022 300934
rect 11786 265018 12022 265254
rect 11786 264698 12022 264934
rect 11786 229018 12022 229254
rect 11786 228698 12022 228934
rect 11786 193018 12022 193254
rect 11786 192698 12022 192934
rect 11786 157018 12022 157254
rect 11786 156698 12022 156934
rect 11786 121018 12022 121254
rect 11786 120698 12022 120934
rect 8186 81418 8422 81654
rect 8186 81098 8422 81334
rect 8186 45418 8422 45654
rect 8186 45098 8422 45334
rect 8186 9418 8422 9654
rect 8186 9098 8422 9334
rect -5574 -4342 -5338 -4106
rect -5574 -4662 -5338 -4426
rect 8186 -4342 8422 -4106
rect 8186 -4662 8422 -4426
rect -6514 -5282 -6278 -5046
rect -6514 -5602 -6278 -5366
rect 11786 85018 12022 85254
rect 11786 84698 12022 84934
rect 11786 49018 12022 49254
rect 11786 48698 12022 48934
rect 11786 13018 12022 13254
rect 11786 12698 12022 12934
rect -7454 -6222 -7218 -5986
rect -7454 -6542 -7218 -6306
rect 18986 705542 19222 705778
rect 18986 705222 19222 705458
rect 18986 668218 19222 668454
rect 18986 667898 19222 668134
rect 18986 632218 19222 632454
rect 18986 631898 19222 632134
rect 18986 596218 19222 596454
rect 18986 595898 19222 596134
rect 18986 560218 19222 560454
rect 18986 559898 19222 560134
rect 18986 524218 19222 524454
rect 18986 523898 19222 524134
rect 18986 488218 19222 488454
rect 18986 487898 19222 488134
rect 18986 452218 19222 452454
rect 18986 451898 19222 452134
rect 18986 416218 19222 416454
rect 18986 415898 19222 416134
rect 18986 380218 19222 380454
rect 18986 379898 19222 380134
rect 18986 344218 19222 344454
rect 18986 343898 19222 344134
rect 18986 308218 19222 308454
rect 18986 307898 19222 308134
rect 18986 272218 19222 272454
rect 18986 271898 19222 272134
rect 18986 236218 19222 236454
rect 18986 235898 19222 236134
rect 18986 200218 19222 200454
rect 18986 199898 19222 200134
rect 18986 164218 19222 164454
rect 18986 163898 19222 164134
rect 18986 128218 19222 128454
rect 18986 127898 19222 128134
rect 18986 92218 19222 92454
rect 18986 91898 19222 92134
rect 18986 56218 19222 56454
rect 18986 55898 19222 56134
rect 18986 20218 19222 20454
rect 18986 19898 19222 20134
rect 18986 -1522 19222 -1286
rect 18986 -1842 19222 -1606
rect 22586 671818 22822 672054
rect 22586 671498 22822 671734
rect 22586 635818 22822 636054
rect 22586 635498 22822 635734
rect 22586 599818 22822 600054
rect 22586 599498 22822 599734
rect 22586 563818 22822 564054
rect 22586 563498 22822 563734
rect 22586 527818 22822 528054
rect 22586 527498 22822 527734
rect 22586 491818 22822 492054
rect 22586 491498 22822 491734
rect 22586 455818 22822 456054
rect 22586 455498 22822 455734
rect 22586 419818 22822 420054
rect 22586 419498 22822 419734
rect 22586 383818 22822 384054
rect 22586 383498 22822 383734
rect 22586 347818 22822 348054
rect 22586 347498 22822 347734
rect 22586 311818 22822 312054
rect 22586 311498 22822 311734
rect 22586 275818 22822 276054
rect 22586 275498 22822 275734
rect 22586 239818 22822 240054
rect 22586 239498 22822 239734
rect 22586 203818 22822 204054
rect 22586 203498 22822 203734
rect 22586 167818 22822 168054
rect 22586 167498 22822 167734
rect 22586 131818 22822 132054
rect 22586 131498 22822 131734
rect 22586 95818 22822 96054
rect 22586 95498 22822 95734
rect 22586 59818 22822 60054
rect 22586 59498 22822 59734
rect 22586 23818 22822 24054
rect 22586 23498 22822 23734
rect 22586 -3402 22822 -3166
rect 22586 -3722 22822 -3486
rect 26186 675418 26422 675654
rect 26186 675098 26422 675334
rect 26186 639418 26422 639654
rect 26186 639098 26422 639334
rect 26186 603418 26422 603654
rect 26186 603098 26422 603334
rect 26186 567418 26422 567654
rect 26186 567098 26422 567334
rect 26186 531418 26422 531654
rect 26186 531098 26422 531334
rect 26186 495418 26422 495654
rect 26186 495098 26422 495334
rect 26186 459418 26422 459654
rect 26186 459098 26422 459334
rect 26186 423418 26422 423654
rect 26186 423098 26422 423334
rect 26186 387418 26422 387654
rect 26186 387098 26422 387334
rect 26186 351418 26422 351654
rect 26186 351098 26422 351334
rect 26186 315418 26422 315654
rect 26186 315098 26422 315334
rect 26186 279418 26422 279654
rect 26186 279098 26422 279334
rect 26186 243418 26422 243654
rect 26186 243098 26422 243334
rect 26186 207418 26422 207654
rect 26186 207098 26422 207334
rect 26186 171418 26422 171654
rect 26186 171098 26422 171334
rect 26186 135418 26422 135654
rect 26186 135098 26422 135334
rect 26186 99418 26422 99654
rect 26186 99098 26422 99334
rect 47786 710242 48022 710478
rect 47786 709922 48022 710158
rect 44186 708362 44422 708598
rect 44186 708042 44422 708278
rect 40586 706482 40822 706718
rect 40586 706162 40822 706398
rect 29786 679018 30022 679254
rect 29786 678698 30022 678934
rect 29786 643018 30022 643254
rect 29786 642698 30022 642934
rect 29786 607018 30022 607254
rect 29786 606698 30022 606934
rect 29786 571018 30022 571254
rect 29786 570698 30022 570934
rect 29786 535018 30022 535254
rect 29786 534698 30022 534934
rect 29786 499018 30022 499254
rect 29786 498698 30022 498934
rect 29786 463018 30022 463254
rect 29786 462698 30022 462934
rect 29786 427018 30022 427254
rect 29786 426698 30022 426934
rect 29786 391018 30022 391254
rect 29786 390698 30022 390934
rect 29786 355018 30022 355254
rect 29786 354698 30022 354934
rect 29786 319018 30022 319254
rect 29786 318698 30022 318934
rect 29786 283018 30022 283254
rect 29786 282698 30022 282934
rect 29786 247018 30022 247254
rect 29786 246698 30022 246934
rect 29786 211018 30022 211254
rect 29786 210698 30022 210934
rect 29786 175018 30022 175254
rect 29786 174698 30022 174934
rect 29786 139018 30022 139254
rect 29786 138698 30022 138934
rect 29786 103018 30022 103254
rect 29786 102698 30022 102934
rect 26186 63418 26422 63654
rect 26186 63098 26422 63334
rect 26186 27418 26422 27654
rect 26186 27098 26422 27334
rect 26186 -5282 26422 -5046
rect 26186 -5602 26422 -5366
rect 29786 67018 30022 67254
rect 29786 66698 30022 66934
rect 29786 31018 30022 31254
rect 29786 30698 30022 30934
rect 11786 -6222 12022 -5986
rect 11786 -6542 12022 -6306
rect -8394 -7162 -8158 -6926
rect -8394 -7482 -8158 -7246
rect 36986 704602 37222 704838
rect 36986 704282 37222 704518
rect 36986 686218 37222 686454
rect 36986 685898 37222 686134
rect 36986 650218 37222 650454
rect 36986 649898 37222 650134
rect 36986 614218 37222 614454
rect 36986 613898 37222 614134
rect 36986 578218 37222 578454
rect 36986 577898 37222 578134
rect 36986 542218 37222 542454
rect 36986 541898 37222 542134
rect 36986 506218 37222 506454
rect 36986 505898 37222 506134
rect 36986 470218 37222 470454
rect 36986 469898 37222 470134
rect 36986 434218 37222 434454
rect 36986 433898 37222 434134
rect 36986 398218 37222 398454
rect 36986 397898 37222 398134
rect 36986 362218 37222 362454
rect 36986 361898 37222 362134
rect 36986 326218 37222 326454
rect 36986 325898 37222 326134
rect 36986 290218 37222 290454
rect 36986 289898 37222 290134
rect 36986 254218 37222 254454
rect 36986 253898 37222 254134
rect 36986 218218 37222 218454
rect 36986 217898 37222 218134
rect 36986 182218 37222 182454
rect 36986 181898 37222 182134
rect 36986 146218 37222 146454
rect 36986 145898 37222 146134
rect 36986 110218 37222 110454
rect 36986 109898 37222 110134
rect 36986 74218 37222 74454
rect 36986 73898 37222 74134
rect 36986 38218 37222 38454
rect 36986 37898 37222 38134
rect 36986 2218 37222 2454
rect 36986 1898 37222 2134
rect 36986 -582 37222 -346
rect 36986 -902 37222 -666
rect 40586 689818 40822 690054
rect 40586 689498 40822 689734
rect 40586 653818 40822 654054
rect 40586 653498 40822 653734
rect 40586 617818 40822 618054
rect 40586 617498 40822 617734
rect 40586 581818 40822 582054
rect 40586 581498 40822 581734
rect 40586 545818 40822 546054
rect 40586 545498 40822 545734
rect 40586 509818 40822 510054
rect 40586 509498 40822 509734
rect 40586 473818 40822 474054
rect 40586 473498 40822 473734
rect 40586 437818 40822 438054
rect 40586 437498 40822 437734
rect 40586 401818 40822 402054
rect 40586 401498 40822 401734
rect 40586 365818 40822 366054
rect 40586 365498 40822 365734
rect 40586 329818 40822 330054
rect 40586 329498 40822 329734
rect 40586 293818 40822 294054
rect 40586 293498 40822 293734
rect 40586 257818 40822 258054
rect 40586 257498 40822 257734
rect 40586 221818 40822 222054
rect 40586 221498 40822 221734
rect 40586 185818 40822 186054
rect 40586 185498 40822 185734
rect 40586 149818 40822 150054
rect 40586 149498 40822 149734
rect 40586 113818 40822 114054
rect 40586 113498 40822 113734
rect 40586 77818 40822 78054
rect 40586 77498 40822 77734
rect 40586 41818 40822 42054
rect 40586 41498 40822 41734
rect 40586 5818 40822 6054
rect 40586 5498 40822 5734
rect 40586 -2462 40822 -2226
rect 40586 -2782 40822 -2546
rect 44186 693418 44422 693654
rect 44186 693098 44422 693334
rect 44186 657418 44422 657654
rect 44186 657098 44422 657334
rect 44186 621418 44422 621654
rect 44186 621098 44422 621334
rect 44186 585418 44422 585654
rect 44186 585098 44422 585334
rect 44186 549418 44422 549654
rect 44186 549098 44422 549334
rect 44186 513418 44422 513654
rect 44186 513098 44422 513334
rect 44186 477418 44422 477654
rect 44186 477098 44422 477334
rect 44186 441418 44422 441654
rect 44186 441098 44422 441334
rect 44186 405418 44422 405654
rect 44186 405098 44422 405334
rect 44186 369418 44422 369654
rect 44186 369098 44422 369334
rect 44186 333418 44422 333654
rect 44186 333098 44422 333334
rect 44186 297418 44422 297654
rect 44186 297098 44422 297334
rect 44186 261418 44422 261654
rect 44186 261098 44422 261334
rect 44186 225418 44422 225654
rect 44186 225098 44422 225334
rect 44186 189418 44422 189654
rect 44186 189098 44422 189334
rect 44186 153418 44422 153654
rect 44186 153098 44422 153334
rect 44186 117418 44422 117654
rect 44186 117098 44422 117334
rect 44186 81418 44422 81654
rect 44186 81098 44422 81334
rect 44186 45418 44422 45654
rect 44186 45098 44422 45334
rect 44186 9418 44422 9654
rect 44186 9098 44422 9334
rect 44186 -4342 44422 -4106
rect 44186 -4662 44422 -4426
rect 65786 711182 66022 711418
rect 65786 710862 66022 711098
rect 62186 709302 62422 709538
rect 62186 708982 62422 709218
rect 58586 707422 58822 707658
rect 58586 707102 58822 707338
rect 47786 697018 48022 697254
rect 47786 696698 48022 696934
rect 47786 661018 48022 661254
rect 47786 660698 48022 660934
rect 47786 625018 48022 625254
rect 47786 624698 48022 624934
rect 47786 589018 48022 589254
rect 47786 588698 48022 588934
rect 47786 553018 48022 553254
rect 47786 552698 48022 552934
rect 47786 517018 48022 517254
rect 47786 516698 48022 516934
rect 47786 481018 48022 481254
rect 47786 480698 48022 480934
rect 47786 445018 48022 445254
rect 47786 444698 48022 444934
rect 47786 409018 48022 409254
rect 47786 408698 48022 408934
rect 47786 373018 48022 373254
rect 47786 372698 48022 372934
rect 47786 337018 48022 337254
rect 47786 336698 48022 336934
rect 47786 301018 48022 301254
rect 47786 300698 48022 300934
rect 47786 265018 48022 265254
rect 47786 264698 48022 264934
rect 47786 229018 48022 229254
rect 47786 228698 48022 228934
rect 47786 193018 48022 193254
rect 47786 192698 48022 192934
rect 47786 157018 48022 157254
rect 47786 156698 48022 156934
rect 47786 121018 48022 121254
rect 47786 120698 48022 120934
rect 54986 705542 55222 705778
rect 54986 705222 55222 705458
rect 54986 668218 55222 668454
rect 54986 667898 55222 668134
rect 54986 632218 55222 632454
rect 54986 631898 55222 632134
rect 54986 596218 55222 596454
rect 54986 595898 55222 596134
rect 54986 560218 55222 560454
rect 54986 559898 55222 560134
rect 54986 524218 55222 524454
rect 54986 523898 55222 524134
rect 54986 488218 55222 488454
rect 54986 487898 55222 488134
rect 54986 452218 55222 452454
rect 54986 451898 55222 452134
rect 54986 416218 55222 416454
rect 54986 415898 55222 416134
rect 54986 380218 55222 380454
rect 54986 379898 55222 380134
rect 54986 344218 55222 344454
rect 54986 343898 55222 344134
rect 54986 308218 55222 308454
rect 54986 307898 55222 308134
rect 54986 272218 55222 272454
rect 54986 271898 55222 272134
rect 54986 236218 55222 236454
rect 54986 235898 55222 236134
rect 54986 200218 55222 200454
rect 54986 199898 55222 200134
rect 54986 164218 55222 164454
rect 54986 163898 55222 164134
rect 54986 128218 55222 128454
rect 54986 127898 55222 128134
rect 47786 85018 48022 85254
rect 47786 84698 48022 84934
rect 47786 49018 48022 49254
rect 47786 48698 48022 48934
rect 47786 13018 48022 13254
rect 47786 12698 48022 12934
rect 29786 -7162 30022 -6926
rect 29786 -7482 30022 -7246
rect 58586 671818 58822 672054
rect 58586 671498 58822 671734
rect 58586 635818 58822 636054
rect 58586 635498 58822 635734
rect 58586 599818 58822 600054
rect 58586 599498 58822 599734
rect 58586 563818 58822 564054
rect 58586 563498 58822 563734
rect 58586 527818 58822 528054
rect 58586 527498 58822 527734
rect 58586 491818 58822 492054
rect 58586 491498 58822 491734
rect 58586 455818 58822 456054
rect 58586 455498 58822 455734
rect 58586 419818 58822 420054
rect 58586 419498 58822 419734
rect 58586 383818 58822 384054
rect 58586 383498 58822 383734
rect 58586 347818 58822 348054
rect 58586 347498 58822 347734
rect 58586 311818 58822 312054
rect 58586 311498 58822 311734
rect 58586 275818 58822 276054
rect 58586 275498 58822 275734
rect 58586 239818 58822 240054
rect 58586 239498 58822 239734
rect 58586 203818 58822 204054
rect 58586 203498 58822 203734
rect 58586 167818 58822 168054
rect 58586 167498 58822 167734
rect 58586 131818 58822 132054
rect 58586 131498 58822 131734
rect 58586 95818 58822 96054
rect 58586 95498 58822 95734
rect 54986 92218 55222 92454
rect 54986 91898 55222 92134
rect 54986 56218 55222 56454
rect 54986 55898 55222 56134
rect 54986 20218 55222 20454
rect 54986 19898 55222 20134
rect 54986 -1522 55222 -1286
rect 54986 -1842 55222 -1606
rect 58586 59818 58822 60054
rect 58586 59498 58822 59734
rect 58586 23818 58822 24054
rect 58586 23498 58822 23734
rect 58586 -3402 58822 -3166
rect 58586 -3722 58822 -3486
rect 62186 675418 62422 675654
rect 62186 675098 62422 675334
rect 62186 639418 62422 639654
rect 62186 639098 62422 639334
rect 62186 603418 62422 603654
rect 62186 603098 62422 603334
rect 62186 567418 62422 567654
rect 62186 567098 62422 567334
rect 62186 531418 62422 531654
rect 62186 531098 62422 531334
rect 62186 495418 62422 495654
rect 62186 495098 62422 495334
rect 62186 459418 62422 459654
rect 62186 459098 62422 459334
rect 62186 423418 62422 423654
rect 62186 423098 62422 423334
rect 62186 387418 62422 387654
rect 62186 387098 62422 387334
rect 62186 351418 62422 351654
rect 62186 351098 62422 351334
rect 62186 315418 62422 315654
rect 62186 315098 62422 315334
rect 62186 279418 62422 279654
rect 62186 279098 62422 279334
rect 62186 243418 62422 243654
rect 62186 243098 62422 243334
rect 62186 207418 62422 207654
rect 62186 207098 62422 207334
rect 62186 171418 62422 171654
rect 62186 171098 62422 171334
rect 62186 135418 62422 135654
rect 62186 135098 62422 135334
rect 62186 99418 62422 99654
rect 62186 99098 62422 99334
rect 62186 63418 62422 63654
rect 62186 63098 62422 63334
rect 62186 27418 62422 27654
rect 62186 27098 62422 27334
rect 62186 -5282 62422 -5046
rect 62186 -5602 62422 -5366
rect 83786 710242 84022 710478
rect 83786 709922 84022 710158
rect 80186 708362 80422 708598
rect 80186 708042 80422 708278
rect 76586 706482 76822 706718
rect 76586 706162 76822 706398
rect 65786 679018 66022 679254
rect 65786 678698 66022 678934
rect 65786 643018 66022 643254
rect 65786 642698 66022 642934
rect 65786 607018 66022 607254
rect 65786 606698 66022 606934
rect 65786 571018 66022 571254
rect 65786 570698 66022 570934
rect 65786 535018 66022 535254
rect 65786 534698 66022 534934
rect 65786 499018 66022 499254
rect 65786 498698 66022 498934
rect 65786 463018 66022 463254
rect 65786 462698 66022 462934
rect 65786 427018 66022 427254
rect 65786 426698 66022 426934
rect 65786 391018 66022 391254
rect 65786 390698 66022 390934
rect 65786 355018 66022 355254
rect 65786 354698 66022 354934
rect 65786 319018 66022 319254
rect 65786 318698 66022 318934
rect 65786 283018 66022 283254
rect 65786 282698 66022 282934
rect 65786 247018 66022 247254
rect 65786 246698 66022 246934
rect 65786 211018 66022 211254
rect 65786 210698 66022 210934
rect 65786 175018 66022 175254
rect 65786 174698 66022 174934
rect 65786 139018 66022 139254
rect 65786 138698 66022 138934
rect 65786 103018 66022 103254
rect 65786 102698 66022 102934
rect 72986 704602 73222 704838
rect 72986 704282 73222 704518
rect 72986 686218 73222 686454
rect 72986 685898 73222 686134
rect 72986 650218 73222 650454
rect 72986 649898 73222 650134
rect 72986 614218 73222 614454
rect 72986 613898 73222 614134
rect 72986 578218 73222 578454
rect 72986 577898 73222 578134
rect 72986 542218 73222 542454
rect 72986 541898 73222 542134
rect 72986 506218 73222 506454
rect 72986 505898 73222 506134
rect 72986 470218 73222 470454
rect 72986 469898 73222 470134
rect 72986 434218 73222 434454
rect 72986 433898 73222 434134
rect 72986 398218 73222 398454
rect 72986 397898 73222 398134
rect 72986 362218 73222 362454
rect 72986 361898 73222 362134
rect 72986 326218 73222 326454
rect 72986 325898 73222 326134
rect 72986 290218 73222 290454
rect 72986 289898 73222 290134
rect 72986 254218 73222 254454
rect 72986 253898 73222 254134
rect 72986 218218 73222 218454
rect 72986 217898 73222 218134
rect 72986 182218 73222 182454
rect 72986 181898 73222 182134
rect 72986 146218 73222 146454
rect 72986 145898 73222 146134
rect 72986 110218 73222 110454
rect 72986 109898 73222 110134
rect 65786 67018 66022 67254
rect 65786 66698 66022 66934
rect 65786 31018 66022 31254
rect 65786 30698 66022 30934
rect 47786 -6222 48022 -5986
rect 47786 -6542 48022 -6306
rect 72986 74218 73222 74454
rect 72986 73898 73222 74134
rect 72986 38218 73222 38454
rect 72986 37898 73222 38134
rect 72986 2218 73222 2454
rect 72986 1898 73222 2134
rect 72986 -582 73222 -346
rect 72986 -902 73222 -666
rect 76586 689818 76822 690054
rect 76586 689498 76822 689734
rect 76586 653818 76822 654054
rect 76586 653498 76822 653734
rect 76586 617818 76822 618054
rect 76586 617498 76822 617734
rect 76586 581818 76822 582054
rect 76586 581498 76822 581734
rect 76586 545818 76822 546054
rect 76586 545498 76822 545734
rect 76586 509818 76822 510054
rect 76586 509498 76822 509734
rect 76586 473818 76822 474054
rect 76586 473498 76822 473734
rect 76586 437818 76822 438054
rect 76586 437498 76822 437734
rect 76586 401818 76822 402054
rect 76586 401498 76822 401734
rect 76586 365818 76822 366054
rect 76586 365498 76822 365734
rect 76586 329818 76822 330054
rect 76586 329498 76822 329734
rect 76586 293818 76822 294054
rect 76586 293498 76822 293734
rect 76586 257818 76822 258054
rect 76586 257498 76822 257734
rect 76586 221818 76822 222054
rect 76586 221498 76822 221734
rect 76586 185818 76822 186054
rect 76586 185498 76822 185734
rect 76586 149818 76822 150054
rect 76586 149498 76822 149734
rect 76586 113818 76822 114054
rect 76586 113498 76822 113734
rect 76586 77818 76822 78054
rect 76586 77498 76822 77734
rect 76586 41818 76822 42054
rect 76586 41498 76822 41734
rect 76586 5818 76822 6054
rect 76586 5498 76822 5734
rect 76586 -2462 76822 -2226
rect 76586 -2782 76822 -2546
rect 80186 693418 80422 693654
rect 80186 693098 80422 693334
rect 80186 657418 80422 657654
rect 80186 657098 80422 657334
rect 80186 621418 80422 621654
rect 80186 621098 80422 621334
rect 80186 585418 80422 585654
rect 80186 585098 80422 585334
rect 80186 549418 80422 549654
rect 80186 549098 80422 549334
rect 80186 513418 80422 513654
rect 80186 513098 80422 513334
rect 80186 477418 80422 477654
rect 80186 477098 80422 477334
rect 80186 441418 80422 441654
rect 80186 441098 80422 441334
rect 80186 405418 80422 405654
rect 80186 405098 80422 405334
rect 80186 369418 80422 369654
rect 80186 369098 80422 369334
rect 80186 333418 80422 333654
rect 80186 333098 80422 333334
rect 80186 297418 80422 297654
rect 80186 297098 80422 297334
rect 80186 261418 80422 261654
rect 80186 261098 80422 261334
rect 80186 225418 80422 225654
rect 80186 225098 80422 225334
rect 80186 189418 80422 189654
rect 80186 189098 80422 189334
rect 80186 153418 80422 153654
rect 80186 153098 80422 153334
rect 80186 117418 80422 117654
rect 80186 117098 80422 117334
rect 80186 81418 80422 81654
rect 80186 81098 80422 81334
rect 80186 45418 80422 45654
rect 80186 45098 80422 45334
rect 80186 9418 80422 9654
rect 80186 9098 80422 9334
rect 80186 -4342 80422 -4106
rect 80186 -4662 80422 -4426
rect 101786 711182 102022 711418
rect 101786 710862 102022 711098
rect 98186 709302 98422 709538
rect 98186 708982 98422 709218
rect 94586 707422 94822 707658
rect 94586 707102 94822 707338
rect 83786 697018 84022 697254
rect 83786 696698 84022 696934
rect 83786 661018 84022 661254
rect 83786 660698 84022 660934
rect 83786 625018 84022 625254
rect 83786 624698 84022 624934
rect 83786 589018 84022 589254
rect 83786 588698 84022 588934
rect 83786 553018 84022 553254
rect 83786 552698 84022 552934
rect 83786 517018 84022 517254
rect 83786 516698 84022 516934
rect 83786 481018 84022 481254
rect 83786 480698 84022 480934
rect 83786 445018 84022 445254
rect 83786 444698 84022 444934
rect 83786 409018 84022 409254
rect 83786 408698 84022 408934
rect 83786 373018 84022 373254
rect 83786 372698 84022 372934
rect 83786 337018 84022 337254
rect 83786 336698 84022 336934
rect 83786 301018 84022 301254
rect 83786 300698 84022 300934
rect 83786 265018 84022 265254
rect 83786 264698 84022 264934
rect 83786 229018 84022 229254
rect 83786 228698 84022 228934
rect 83786 193018 84022 193254
rect 83786 192698 84022 192934
rect 83786 157018 84022 157254
rect 83786 156698 84022 156934
rect 83786 121018 84022 121254
rect 83786 120698 84022 120934
rect 90986 705542 91222 705778
rect 90986 705222 91222 705458
rect 90986 668218 91222 668454
rect 90986 667898 91222 668134
rect 90986 632218 91222 632454
rect 90986 631898 91222 632134
rect 90986 596218 91222 596454
rect 90986 595898 91222 596134
rect 90986 560218 91222 560454
rect 90986 559898 91222 560134
rect 90986 524218 91222 524454
rect 90986 523898 91222 524134
rect 90986 488218 91222 488454
rect 90986 487898 91222 488134
rect 90986 452218 91222 452454
rect 90986 451898 91222 452134
rect 90986 416218 91222 416454
rect 90986 415898 91222 416134
rect 90986 380218 91222 380454
rect 90986 379898 91222 380134
rect 90986 344218 91222 344454
rect 90986 343898 91222 344134
rect 90986 308218 91222 308454
rect 90986 307898 91222 308134
rect 90986 272218 91222 272454
rect 90986 271898 91222 272134
rect 90986 236218 91222 236454
rect 90986 235898 91222 236134
rect 90986 200218 91222 200454
rect 90986 199898 91222 200134
rect 90986 164218 91222 164454
rect 90986 163898 91222 164134
rect 90986 128218 91222 128454
rect 90986 127898 91222 128134
rect 83786 85018 84022 85254
rect 83786 84698 84022 84934
rect 83786 49018 84022 49254
rect 83786 48698 84022 48934
rect 83786 13018 84022 13254
rect 83786 12698 84022 12934
rect 65786 -7162 66022 -6926
rect 65786 -7482 66022 -7246
rect 90986 92218 91222 92454
rect 90986 91898 91222 92134
rect 90986 56218 91222 56454
rect 90986 55898 91222 56134
rect 90986 20218 91222 20454
rect 90986 19898 91222 20134
rect 90986 -1522 91222 -1286
rect 90986 -1842 91222 -1606
rect 94586 671818 94822 672054
rect 94586 671498 94822 671734
rect 94586 635818 94822 636054
rect 94586 635498 94822 635734
rect 94586 599818 94822 600054
rect 94586 599498 94822 599734
rect 94586 563818 94822 564054
rect 94586 563498 94822 563734
rect 94586 527818 94822 528054
rect 94586 527498 94822 527734
rect 94586 491818 94822 492054
rect 94586 491498 94822 491734
rect 94586 455818 94822 456054
rect 94586 455498 94822 455734
rect 94586 419818 94822 420054
rect 94586 419498 94822 419734
rect 94586 383818 94822 384054
rect 94586 383498 94822 383734
rect 94586 347818 94822 348054
rect 94586 347498 94822 347734
rect 94586 311818 94822 312054
rect 94586 311498 94822 311734
rect 94586 275818 94822 276054
rect 94586 275498 94822 275734
rect 94586 239818 94822 240054
rect 94586 239498 94822 239734
rect 94586 203818 94822 204054
rect 94586 203498 94822 203734
rect 94586 167818 94822 168054
rect 94586 167498 94822 167734
rect 94586 131818 94822 132054
rect 94586 131498 94822 131734
rect 94586 95818 94822 96054
rect 94586 95498 94822 95734
rect 94586 59818 94822 60054
rect 94586 59498 94822 59734
rect 94586 23818 94822 24054
rect 94586 23498 94822 23734
rect 94586 -3402 94822 -3166
rect 94586 -3722 94822 -3486
rect 98186 675418 98422 675654
rect 98186 675098 98422 675334
rect 98186 639418 98422 639654
rect 98186 639098 98422 639334
rect 98186 603418 98422 603654
rect 98186 603098 98422 603334
rect 98186 567418 98422 567654
rect 98186 567098 98422 567334
rect 98186 531418 98422 531654
rect 98186 531098 98422 531334
rect 98186 495418 98422 495654
rect 98186 495098 98422 495334
rect 98186 459418 98422 459654
rect 98186 459098 98422 459334
rect 98186 423418 98422 423654
rect 98186 423098 98422 423334
rect 98186 387418 98422 387654
rect 98186 387098 98422 387334
rect 98186 351418 98422 351654
rect 98186 351098 98422 351334
rect 98186 315418 98422 315654
rect 98186 315098 98422 315334
rect 98186 279418 98422 279654
rect 98186 279098 98422 279334
rect 98186 243418 98422 243654
rect 98186 243098 98422 243334
rect 98186 207418 98422 207654
rect 98186 207098 98422 207334
rect 98186 171418 98422 171654
rect 98186 171098 98422 171334
rect 98186 135418 98422 135654
rect 98186 135098 98422 135334
rect 98186 99418 98422 99654
rect 98186 99098 98422 99334
rect 98186 63418 98422 63654
rect 98186 63098 98422 63334
rect 98186 27418 98422 27654
rect 98186 27098 98422 27334
rect 98186 -5282 98422 -5046
rect 98186 -5602 98422 -5366
rect 119786 710242 120022 710478
rect 119786 709922 120022 710158
rect 116186 708362 116422 708598
rect 116186 708042 116422 708278
rect 112586 706482 112822 706718
rect 112586 706162 112822 706398
rect 101786 679018 102022 679254
rect 101786 678698 102022 678934
rect 101786 643018 102022 643254
rect 101786 642698 102022 642934
rect 101786 607018 102022 607254
rect 101786 606698 102022 606934
rect 101786 571018 102022 571254
rect 101786 570698 102022 570934
rect 101786 535018 102022 535254
rect 101786 534698 102022 534934
rect 101786 499018 102022 499254
rect 101786 498698 102022 498934
rect 101786 463018 102022 463254
rect 101786 462698 102022 462934
rect 101786 427018 102022 427254
rect 101786 426698 102022 426934
rect 101786 391018 102022 391254
rect 101786 390698 102022 390934
rect 101786 355018 102022 355254
rect 101786 354698 102022 354934
rect 101786 319018 102022 319254
rect 101786 318698 102022 318934
rect 101786 283018 102022 283254
rect 101786 282698 102022 282934
rect 101786 247018 102022 247254
rect 101786 246698 102022 246934
rect 101786 211018 102022 211254
rect 101786 210698 102022 210934
rect 101786 175018 102022 175254
rect 101786 174698 102022 174934
rect 101786 139018 102022 139254
rect 101786 138698 102022 138934
rect 101786 103018 102022 103254
rect 101786 102698 102022 102934
rect 108986 704602 109222 704838
rect 108986 704282 109222 704518
rect 108986 686218 109222 686454
rect 108986 685898 109222 686134
rect 108986 650218 109222 650454
rect 108986 649898 109222 650134
rect 108986 614218 109222 614454
rect 108986 613898 109222 614134
rect 108986 578218 109222 578454
rect 108986 577898 109222 578134
rect 108986 542218 109222 542454
rect 108986 541898 109222 542134
rect 108986 506218 109222 506454
rect 108986 505898 109222 506134
rect 108986 470218 109222 470454
rect 108986 469898 109222 470134
rect 108986 434218 109222 434454
rect 108986 433898 109222 434134
rect 108986 398218 109222 398454
rect 108986 397898 109222 398134
rect 108986 362218 109222 362454
rect 108986 361898 109222 362134
rect 108986 326218 109222 326454
rect 108986 325898 109222 326134
rect 108986 290218 109222 290454
rect 108986 289898 109222 290134
rect 108986 254218 109222 254454
rect 108986 253898 109222 254134
rect 108986 218218 109222 218454
rect 108986 217898 109222 218134
rect 108986 182218 109222 182454
rect 108986 181898 109222 182134
rect 108986 146218 109222 146454
rect 108986 145898 109222 146134
rect 108986 110218 109222 110454
rect 108986 109898 109222 110134
rect 101786 67018 102022 67254
rect 101786 66698 102022 66934
rect 101786 31018 102022 31254
rect 101786 30698 102022 30934
rect 83786 -6222 84022 -5986
rect 83786 -6542 84022 -6306
rect 108986 74218 109222 74454
rect 108986 73898 109222 74134
rect 108986 38218 109222 38454
rect 108986 37898 109222 38134
rect 108986 2218 109222 2454
rect 108986 1898 109222 2134
rect 108986 -582 109222 -346
rect 108986 -902 109222 -666
rect 112586 689818 112822 690054
rect 112586 689498 112822 689734
rect 112586 653818 112822 654054
rect 112586 653498 112822 653734
rect 112586 617818 112822 618054
rect 112586 617498 112822 617734
rect 112586 581818 112822 582054
rect 112586 581498 112822 581734
rect 112586 545818 112822 546054
rect 112586 545498 112822 545734
rect 112586 509818 112822 510054
rect 112586 509498 112822 509734
rect 112586 473818 112822 474054
rect 112586 473498 112822 473734
rect 112586 437818 112822 438054
rect 112586 437498 112822 437734
rect 112586 401818 112822 402054
rect 112586 401498 112822 401734
rect 112586 365818 112822 366054
rect 112586 365498 112822 365734
rect 112586 329818 112822 330054
rect 112586 329498 112822 329734
rect 112586 293818 112822 294054
rect 112586 293498 112822 293734
rect 112586 257818 112822 258054
rect 112586 257498 112822 257734
rect 112586 221818 112822 222054
rect 112586 221498 112822 221734
rect 112586 185818 112822 186054
rect 112586 185498 112822 185734
rect 112586 149818 112822 150054
rect 112586 149498 112822 149734
rect 112586 113818 112822 114054
rect 112586 113498 112822 113734
rect 112586 77818 112822 78054
rect 112586 77498 112822 77734
rect 112586 41818 112822 42054
rect 112586 41498 112822 41734
rect 112586 5818 112822 6054
rect 112586 5498 112822 5734
rect 112586 -2462 112822 -2226
rect 112586 -2782 112822 -2546
rect 116186 693418 116422 693654
rect 116186 693098 116422 693334
rect 116186 657418 116422 657654
rect 116186 657098 116422 657334
rect 116186 621418 116422 621654
rect 116186 621098 116422 621334
rect 116186 585418 116422 585654
rect 116186 585098 116422 585334
rect 116186 549418 116422 549654
rect 116186 549098 116422 549334
rect 116186 513418 116422 513654
rect 116186 513098 116422 513334
rect 116186 477418 116422 477654
rect 116186 477098 116422 477334
rect 116186 441418 116422 441654
rect 116186 441098 116422 441334
rect 116186 405418 116422 405654
rect 116186 405098 116422 405334
rect 116186 369418 116422 369654
rect 116186 369098 116422 369334
rect 116186 333418 116422 333654
rect 116186 333098 116422 333334
rect 116186 297418 116422 297654
rect 116186 297098 116422 297334
rect 116186 261418 116422 261654
rect 116186 261098 116422 261334
rect 116186 225418 116422 225654
rect 116186 225098 116422 225334
rect 116186 189418 116422 189654
rect 116186 189098 116422 189334
rect 116186 153418 116422 153654
rect 116186 153098 116422 153334
rect 116186 117418 116422 117654
rect 116186 117098 116422 117334
rect 116186 81418 116422 81654
rect 116186 81098 116422 81334
rect 116186 45418 116422 45654
rect 116186 45098 116422 45334
rect 116186 9418 116422 9654
rect 116186 9098 116422 9334
rect 116186 -4342 116422 -4106
rect 116186 -4662 116422 -4426
rect 137786 711182 138022 711418
rect 137786 710862 138022 711098
rect 134186 709302 134422 709538
rect 134186 708982 134422 709218
rect 130586 707422 130822 707658
rect 130586 707102 130822 707338
rect 119786 697018 120022 697254
rect 119786 696698 120022 696934
rect 119786 661018 120022 661254
rect 119786 660698 120022 660934
rect 119786 625018 120022 625254
rect 119786 624698 120022 624934
rect 119786 589018 120022 589254
rect 119786 588698 120022 588934
rect 119786 553018 120022 553254
rect 119786 552698 120022 552934
rect 119786 517018 120022 517254
rect 119786 516698 120022 516934
rect 119786 481018 120022 481254
rect 119786 480698 120022 480934
rect 119786 445018 120022 445254
rect 119786 444698 120022 444934
rect 119786 409018 120022 409254
rect 119786 408698 120022 408934
rect 119786 373018 120022 373254
rect 119786 372698 120022 372934
rect 119786 337018 120022 337254
rect 119786 336698 120022 336934
rect 119786 301018 120022 301254
rect 119786 300698 120022 300934
rect 119786 265018 120022 265254
rect 119786 264698 120022 264934
rect 119786 229018 120022 229254
rect 119786 228698 120022 228934
rect 119786 193018 120022 193254
rect 119786 192698 120022 192934
rect 119786 157018 120022 157254
rect 119786 156698 120022 156934
rect 119786 121018 120022 121254
rect 119786 120698 120022 120934
rect 126986 705542 127222 705778
rect 126986 705222 127222 705458
rect 126986 668218 127222 668454
rect 126986 667898 127222 668134
rect 126986 632218 127222 632454
rect 126986 631898 127222 632134
rect 126986 596218 127222 596454
rect 126986 595898 127222 596134
rect 126986 560218 127222 560454
rect 126986 559898 127222 560134
rect 126986 524218 127222 524454
rect 126986 523898 127222 524134
rect 126986 488218 127222 488454
rect 126986 487898 127222 488134
rect 126986 452218 127222 452454
rect 126986 451898 127222 452134
rect 126986 416218 127222 416454
rect 126986 415898 127222 416134
rect 126986 380218 127222 380454
rect 126986 379898 127222 380134
rect 126986 344218 127222 344454
rect 126986 343898 127222 344134
rect 126986 308218 127222 308454
rect 126986 307898 127222 308134
rect 126986 272218 127222 272454
rect 126986 271898 127222 272134
rect 126986 236218 127222 236454
rect 126986 235898 127222 236134
rect 126986 200218 127222 200454
rect 126986 199898 127222 200134
rect 126986 164218 127222 164454
rect 126986 163898 127222 164134
rect 126986 128218 127222 128454
rect 126986 127898 127222 128134
rect 119786 85018 120022 85254
rect 119786 84698 120022 84934
rect 119786 49018 120022 49254
rect 119786 48698 120022 48934
rect 119786 13018 120022 13254
rect 119786 12698 120022 12934
rect 101786 -7162 102022 -6926
rect 101786 -7482 102022 -7246
rect 126986 92218 127222 92454
rect 126986 91898 127222 92134
rect 126986 56218 127222 56454
rect 126986 55898 127222 56134
rect 126986 20218 127222 20454
rect 126986 19898 127222 20134
rect 126986 -1522 127222 -1286
rect 126986 -1842 127222 -1606
rect 130586 671818 130822 672054
rect 130586 671498 130822 671734
rect 130586 635818 130822 636054
rect 130586 635498 130822 635734
rect 130586 599818 130822 600054
rect 130586 599498 130822 599734
rect 130586 563818 130822 564054
rect 130586 563498 130822 563734
rect 130586 527818 130822 528054
rect 130586 527498 130822 527734
rect 130586 491818 130822 492054
rect 130586 491498 130822 491734
rect 130586 455818 130822 456054
rect 130586 455498 130822 455734
rect 130586 419818 130822 420054
rect 130586 419498 130822 419734
rect 130586 383818 130822 384054
rect 130586 383498 130822 383734
rect 130586 347818 130822 348054
rect 130586 347498 130822 347734
rect 130586 311818 130822 312054
rect 130586 311498 130822 311734
rect 130586 275818 130822 276054
rect 130586 275498 130822 275734
rect 130586 239818 130822 240054
rect 130586 239498 130822 239734
rect 130586 203818 130822 204054
rect 130586 203498 130822 203734
rect 130586 167818 130822 168054
rect 130586 167498 130822 167734
rect 130586 131818 130822 132054
rect 130586 131498 130822 131734
rect 130586 95818 130822 96054
rect 130586 95498 130822 95734
rect 130586 59818 130822 60054
rect 130586 59498 130822 59734
rect 130586 23818 130822 24054
rect 130586 23498 130822 23734
rect 130586 -3402 130822 -3166
rect 130586 -3722 130822 -3486
rect 134186 675418 134422 675654
rect 134186 675098 134422 675334
rect 134186 639418 134422 639654
rect 134186 639098 134422 639334
rect 134186 603418 134422 603654
rect 134186 603098 134422 603334
rect 134186 567418 134422 567654
rect 134186 567098 134422 567334
rect 134186 531418 134422 531654
rect 134186 531098 134422 531334
rect 134186 495418 134422 495654
rect 134186 495098 134422 495334
rect 134186 459418 134422 459654
rect 134186 459098 134422 459334
rect 134186 423418 134422 423654
rect 134186 423098 134422 423334
rect 134186 387418 134422 387654
rect 134186 387098 134422 387334
rect 134186 351418 134422 351654
rect 134186 351098 134422 351334
rect 134186 315418 134422 315654
rect 134186 315098 134422 315334
rect 134186 279418 134422 279654
rect 134186 279098 134422 279334
rect 134186 243418 134422 243654
rect 134186 243098 134422 243334
rect 134186 207418 134422 207654
rect 134186 207098 134422 207334
rect 134186 171418 134422 171654
rect 134186 171098 134422 171334
rect 134186 135418 134422 135654
rect 134186 135098 134422 135334
rect 134186 99418 134422 99654
rect 134186 99098 134422 99334
rect 134186 63418 134422 63654
rect 134186 63098 134422 63334
rect 134186 27418 134422 27654
rect 134186 27098 134422 27334
rect 134186 -5282 134422 -5046
rect 134186 -5602 134422 -5366
rect 155786 710242 156022 710478
rect 155786 709922 156022 710158
rect 152186 708362 152422 708598
rect 152186 708042 152422 708278
rect 148586 706482 148822 706718
rect 148586 706162 148822 706398
rect 137786 679018 138022 679254
rect 137786 678698 138022 678934
rect 137786 643018 138022 643254
rect 137786 642698 138022 642934
rect 137786 607018 138022 607254
rect 137786 606698 138022 606934
rect 137786 571018 138022 571254
rect 137786 570698 138022 570934
rect 137786 535018 138022 535254
rect 137786 534698 138022 534934
rect 137786 499018 138022 499254
rect 137786 498698 138022 498934
rect 137786 463018 138022 463254
rect 137786 462698 138022 462934
rect 137786 427018 138022 427254
rect 137786 426698 138022 426934
rect 137786 391018 138022 391254
rect 137786 390698 138022 390934
rect 137786 355018 138022 355254
rect 137786 354698 138022 354934
rect 137786 319018 138022 319254
rect 137786 318698 138022 318934
rect 137786 283018 138022 283254
rect 137786 282698 138022 282934
rect 137786 247018 138022 247254
rect 137786 246698 138022 246934
rect 137786 211018 138022 211254
rect 137786 210698 138022 210934
rect 137786 175018 138022 175254
rect 137786 174698 138022 174934
rect 137786 139018 138022 139254
rect 137786 138698 138022 138934
rect 137786 103018 138022 103254
rect 137786 102698 138022 102934
rect 137786 67018 138022 67254
rect 137786 66698 138022 66934
rect 137786 31018 138022 31254
rect 137786 30698 138022 30934
rect 119786 -6222 120022 -5986
rect 119786 -6542 120022 -6306
rect 144986 704602 145222 704838
rect 144986 704282 145222 704518
rect 144986 686218 145222 686454
rect 144986 685898 145222 686134
rect 144986 650218 145222 650454
rect 144986 649898 145222 650134
rect 144986 614218 145222 614454
rect 144986 613898 145222 614134
rect 144986 578218 145222 578454
rect 144986 577898 145222 578134
rect 144986 542218 145222 542454
rect 144986 541898 145222 542134
rect 144986 506218 145222 506454
rect 144986 505898 145222 506134
rect 144986 470218 145222 470454
rect 144986 469898 145222 470134
rect 144986 434218 145222 434454
rect 144986 433898 145222 434134
rect 144986 398218 145222 398454
rect 144986 397898 145222 398134
rect 144986 362218 145222 362454
rect 144986 361898 145222 362134
rect 144986 326218 145222 326454
rect 144986 325898 145222 326134
rect 144986 290218 145222 290454
rect 144986 289898 145222 290134
rect 144986 254218 145222 254454
rect 144986 253898 145222 254134
rect 144986 218218 145222 218454
rect 144986 217898 145222 218134
rect 144986 182218 145222 182454
rect 144986 181898 145222 182134
rect 144986 146218 145222 146454
rect 144986 145898 145222 146134
rect 144986 110218 145222 110454
rect 144986 109898 145222 110134
rect 144986 74218 145222 74454
rect 144986 73898 145222 74134
rect 144986 38218 145222 38454
rect 144986 37898 145222 38134
rect 144986 2218 145222 2454
rect 144986 1898 145222 2134
rect 144986 -582 145222 -346
rect 144986 -902 145222 -666
rect 148586 689818 148822 690054
rect 148586 689498 148822 689734
rect 148586 653818 148822 654054
rect 148586 653498 148822 653734
rect 148586 617818 148822 618054
rect 148586 617498 148822 617734
rect 148586 581818 148822 582054
rect 148586 581498 148822 581734
rect 148586 545818 148822 546054
rect 148586 545498 148822 545734
rect 148586 509818 148822 510054
rect 148586 509498 148822 509734
rect 148586 473818 148822 474054
rect 148586 473498 148822 473734
rect 148586 437818 148822 438054
rect 148586 437498 148822 437734
rect 148586 401818 148822 402054
rect 148586 401498 148822 401734
rect 148586 365818 148822 366054
rect 148586 365498 148822 365734
rect 148586 329818 148822 330054
rect 148586 329498 148822 329734
rect 148586 293818 148822 294054
rect 148586 293498 148822 293734
rect 148586 257818 148822 258054
rect 148586 257498 148822 257734
rect 148586 221818 148822 222054
rect 148586 221498 148822 221734
rect 148586 185818 148822 186054
rect 148586 185498 148822 185734
rect 148586 149818 148822 150054
rect 148586 149498 148822 149734
rect 148586 113818 148822 114054
rect 148586 113498 148822 113734
rect 148586 77818 148822 78054
rect 148586 77498 148822 77734
rect 148586 41818 148822 42054
rect 148586 41498 148822 41734
rect 148586 5818 148822 6054
rect 148586 5498 148822 5734
rect 148586 -2462 148822 -2226
rect 148586 -2782 148822 -2546
rect 152186 693418 152422 693654
rect 152186 693098 152422 693334
rect 152186 657418 152422 657654
rect 152186 657098 152422 657334
rect 152186 621418 152422 621654
rect 152186 621098 152422 621334
rect 152186 585418 152422 585654
rect 152186 585098 152422 585334
rect 152186 549418 152422 549654
rect 152186 549098 152422 549334
rect 152186 513418 152422 513654
rect 152186 513098 152422 513334
rect 152186 477418 152422 477654
rect 152186 477098 152422 477334
rect 152186 441418 152422 441654
rect 152186 441098 152422 441334
rect 152186 405418 152422 405654
rect 152186 405098 152422 405334
rect 152186 369418 152422 369654
rect 152186 369098 152422 369334
rect 152186 333418 152422 333654
rect 152186 333098 152422 333334
rect 152186 297418 152422 297654
rect 152186 297098 152422 297334
rect 152186 261418 152422 261654
rect 152186 261098 152422 261334
rect 152186 225418 152422 225654
rect 152186 225098 152422 225334
rect 152186 189418 152422 189654
rect 152186 189098 152422 189334
rect 152186 153418 152422 153654
rect 152186 153098 152422 153334
rect 152186 117418 152422 117654
rect 152186 117098 152422 117334
rect 152186 81418 152422 81654
rect 152186 81098 152422 81334
rect 152186 45418 152422 45654
rect 152186 45098 152422 45334
rect 152186 9418 152422 9654
rect 152186 9098 152422 9334
rect 152186 -4342 152422 -4106
rect 152186 -4662 152422 -4426
rect 173786 711182 174022 711418
rect 173786 710862 174022 711098
rect 170186 709302 170422 709538
rect 170186 708982 170422 709218
rect 166586 707422 166822 707658
rect 166586 707102 166822 707338
rect 155786 697018 156022 697254
rect 155786 696698 156022 696934
rect 155786 661018 156022 661254
rect 155786 660698 156022 660934
rect 155786 625018 156022 625254
rect 155786 624698 156022 624934
rect 155786 589018 156022 589254
rect 155786 588698 156022 588934
rect 155786 553018 156022 553254
rect 155786 552698 156022 552934
rect 155786 517018 156022 517254
rect 155786 516698 156022 516934
rect 155786 481018 156022 481254
rect 155786 480698 156022 480934
rect 155786 445018 156022 445254
rect 155786 444698 156022 444934
rect 155786 409018 156022 409254
rect 155786 408698 156022 408934
rect 155786 373018 156022 373254
rect 155786 372698 156022 372934
rect 155786 337018 156022 337254
rect 155786 336698 156022 336934
rect 155786 301018 156022 301254
rect 155786 300698 156022 300934
rect 155786 265018 156022 265254
rect 155786 264698 156022 264934
rect 155786 229018 156022 229254
rect 155786 228698 156022 228934
rect 155786 193018 156022 193254
rect 155786 192698 156022 192934
rect 155786 157018 156022 157254
rect 155786 156698 156022 156934
rect 155786 121018 156022 121254
rect 155786 120698 156022 120934
rect 155786 85018 156022 85254
rect 155786 84698 156022 84934
rect 155786 49018 156022 49254
rect 155786 48698 156022 48934
rect 155786 13018 156022 13254
rect 155786 12698 156022 12934
rect 137786 -7162 138022 -6926
rect 137786 -7482 138022 -7246
rect 162986 705542 163222 705778
rect 162986 705222 163222 705458
rect 162986 668218 163222 668454
rect 162986 667898 163222 668134
rect 162986 632218 163222 632454
rect 162986 631898 163222 632134
rect 162986 596218 163222 596454
rect 162986 595898 163222 596134
rect 162986 560218 163222 560454
rect 162986 559898 163222 560134
rect 162986 524218 163222 524454
rect 162986 523898 163222 524134
rect 162986 488218 163222 488454
rect 162986 487898 163222 488134
rect 162986 452218 163222 452454
rect 162986 451898 163222 452134
rect 162986 416218 163222 416454
rect 162986 415898 163222 416134
rect 162986 380218 163222 380454
rect 162986 379898 163222 380134
rect 162986 344218 163222 344454
rect 162986 343898 163222 344134
rect 162986 308218 163222 308454
rect 162986 307898 163222 308134
rect 162986 272218 163222 272454
rect 162986 271898 163222 272134
rect 162986 236218 163222 236454
rect 162986 235898 163222 236134
rect 162986 200218 163222 200454
rect 162986 199898 163222 200134
rect 162986 164218 163222 164454
rect 162986 163898 163222 164134
rect 162986 128218 163222 128454
rect 162986 127898 163222 128134
rect 162986 92218 163222 92454
rect 162986 91898 163222 92134
rect 162986 56218 163222 56454
rect 162986 55898 163222 56134
rect 162986 20218 163222 20454
rect 162986 19898 163222 20134
rect 162986 -1522 163222 -1286
rect 162986 -1842 163222 -1606
rect 166586 671818 166822 672054
rect 166586 671498 166822 671734
rect 166586 635818 166822 636054
rect 166586 635498 166822 635734
rect 166586 599818 166822 600054
rect 166586 599498 166822 599734
rect 166586 563818 166822 564054
rect 166586 563498 166822 563734
rect 166586 527818 166822 528054
rect 166586 527498 166822 527734
rect 166586 491818 166822 492054
rect 166586 491498 166822 491734
rect 166586 455818 166822 456054
rect 166586 455498 166822 455734
rect 166586 419818 166822 420054
rect 166586 419498 166822 419734
rect 166586 383818 166822 384054
rect 166586 383498 166822 383734
rect 166586 347818 166822 348054
rect 166586 347498 166822 347734
rect 166586 311818 166822 312054
rect 166586 311498 166822 311734
rect 166586 275818 166822 276054
rect 166586 275498 166822 275734
rect 166586 239818 166822 240054
rect 166586 239498 166822 239734
rect 166586 203818 166822 204054
rect 166586 203498 166822 203734
rect 166586 167818 166822 168054
rect 166586 167498 166822 167734
rect 166586 131818 166822 132054
rect 166586 131498 166822 131734
rect 166586 95818 166822 96054
rect 166586 95498 166822 95734
rect 166586 59818 166822 60054
rect 166586 59498 166822 59734
rect 166586 23818 166822 24054
rect 166586 23498 166822 23734
rect 166586 -3402 166822 -3166
rect 166586 -3722 166822 -3486
rect 170186 675418 170422 675654
rect 170186 675098 170422 675334
rect 170186 639418 170422 639654
rect 170186 639098 170422 639334
rect 170186 603418 170422 603654
rect 170186 603098 170422 603334
rect 170186 567418 170422 567654
rect 170186 567098 170422 567334
rect 170186 531418 170422 531654
rect 170186 531098 170422 531334
rect 170186 495418 170422 495654
rect 170186 495098 170422 495334
rect 170186 459418 170422 459654
rect 170186 459098 170422 459334
rect 170186 423418 170422 423654
rect 170186 423098 170422 423334
rect 170186 387418 170422 387654
rect 170186 387098 170422 387334
rect 170186 351418 170422 351654
rect 170186 351098 170422 351334
rect 170186 315418 170422 315654
rect 170186 315098 170422 315334
rect 170186 279418 170422 279654
rect 170186 279098 170422 279334
rect 170186 243418 170422 243654
rect 170186 243098 170422 243334
rect 170186 207418 170422 207654
rect 170186 207098 170422 207334
rect 170186 171418 170422 171654
rect 170186 171098 170422 171334
rect 170186 135418 170422 135654
rect 170186 135098 170422 135334
rect 170186 99418 170422 99654
rect 170186 99098 170422 99334
rect 170186 63418 170422 63654
rect 170186 63098 170422 63334
rect 170186 27418 170422 27654
rect 170186 27098 170422 27334
rect 170186 -5282 170422 -5046
rect 170186 -5602 170422 -5366
rect 191786 710242 192022 710478
rect 191786 709922 192022 710158
rect 188186 708362 188422 708598
rect 188186 708042 188422 708278
rect 184586 706482 184822 706718
rect 184586 706162 184822 706398
rect 173786 679018 174022 679254
rect 173786 678698 174022 678934
rect 173786 643018 174022 643254
rect 173786 642698 174022 642934
rect 173786 607018 174022 607254
rect 173786 606698 174022 606934
rect 173786 571018 174022 571254
rect 173786 570698 174022 570934
rect 173786 535018 174022 535254
rect 173786 534698 174022 534934
rect 173786 499018 174022 499254
rect 173786 498698 174022 498934
rect 173786 463018 174022 463254
rect 173786 462698 174022 462934
rect 173786 427018 174022 427254
rect 173786 426698 174022 426934
rect 173786 391018 174022 391254
rect 173786 390698 174022 390934
rect 173786 355018 174022 355254
rect 173786 354698 174022 354934
rect 173786 319018 174022 319254
rect 173786 318698 174022 318934
rect 173786 283018 174022 283254
rect 173786 282698 174022 282934
rect 173786 247018 174022 247254
rect 173786 246698 174022 246934
rect 173786 211018 174022 211254
rect 173786 210698 174022 210934
rect 173786 175018 174022 175254
rect 173786 174698 174022 174934
rect 173786 139018 174022 139254
rect 173786 138698 174022 138934
rect 173786 103018 174022 103254
rect 173786 102698 174022 102934
rect 173786 67018 174022 67254
rect 173786 66698 174022 66934
rect 173786 31018 174022 31254
rect 173786 30698 174022 30934
rect 155786 -6222 156022 -5986
rect 155786 -6542 156022 -6306
rect 180986 704602 181222 704838
rect 180986 704282 181222 704518
rect 180986 686218 181222 686454
rect 180986 685898 181222 686134
rect 180986 650218 181222 650454
rect 180986 649898 181222 650134
rect 180986 614218 181222 614454
rect 180986 613898 181222 614134
rect 180986 578218 181222 578454
rect 180986 577898 181222 578134
rect 180986 542218 181222 542454
rect 180986 541898 181222 542134
rect 180986 506218 181222 506454
rect 180986 505898 181222 506134
rect 180986 470218 181222 470454
rect 180986 469898 181222 470134
rect 180986 434218 181222 434454
rect 180986 433898 181222 434134
rect 180986 398218 181222 398454
rect 180986 397898 181222 398134
rect 180986 362218 181222 362454
rect 180986 361898 181222 362134
rect 180986 326218 181222 326454
rect 180986 325898 181222 326134
rect 180986 290218 181222 290454
rect 180986 289898 181222 290134
rect 180986 254218 181222 254454
rect 180986 253898 181222 254134
rect 180986 218218 181222 218454
rect 180986 217898 181222 218134
rect 180986 182218 181222 182454
rect 180986 181898 181222 182134
rect 180986 146218 181222 146454
rect 180986 145898 181222 146134
rect 180986 110218 181222 110454
rect 180986 109898 181222 110134
rect 180986 74218 181222 74454
rect 180986 73898 181222 74134
rect 180986 38218 181222 38454
rect 180986 37898 181222 38134
rect 180986 2218 181222 2454
rect 180986 1898 181222 2134
rect 180986 -582 181222 -346
rect 180986 -902 181222 -666
rect 184586 689818 184822 690054
rect 184586 689498 184822 689734
rect 184586 653818 184822 654054
rect 184586 653498 184822 653734
rect 184586 617818 184822 618054
rect 184586 617498 184822 617734
rect 184586 581818 184822 582054
rect 184586 581498 184822 581734
rect 184586 545818 184822 546054
rect 184586 545498 184822 545734
rect 184586 509818 184822 510054
rect 184586 509498 184822 509734
rect 184586 473818 184822 474054
rect 184586 473498 184822 473734
rect 184586 437818 184822 438054
rect 184586 437498 184822 437734
rect 184586 401818 184822 402054
rect 184586 401498 184822 401734
rect 184586 365818 184822 366054
rect 184586 365498 184822 365734
rect 184586 329818 184822 330054
rect 184586 329498 184822 329734
rect 184586 293818 184822 294054
rect 184586 293498 184822 293734
rect 184586 257818 184822 258054
rect 184586 257498 184822 257734
rect 184586 221818 184822 222054
rect 184586 221498 184822 221734
rect 184586 185818 184822 186054
rect 184586 185498 184822 185734
rect 184586 149818 184822 150054
rect 184586 149498 184822 149734
rect 184586 113818 184822 114054
rect 184586 113498 184822 113734
rect 184586 77818 184822 78054
rect 184586 77498 184822 77734
rect 184586 41818 184822 42054
rect 184586 41498 184822 41734
rect 184586 5818 184822 6054
rect 184586 5498 184822 5734
rect 184586 -2462 184822 -2226
rect 184586 -2782 184822 -2546
rect 188186 693418 188422 693654
rect 188186 693098 188422 693334
rect 188186 657418 188422 657654
rect 188186 657098 188422 657334
rect 188186 621418 188422 621654
rect 188186 621098 188422 621334
rect 188186 585418 188422 585654
rect 188186 585098 188422 585334
rect 188186 549418 188422 549654
rect 188186 549098 188422 549334
rect 188186 513418 188422 513654
rect 188186 513098 188422 513334
rect 188186 477418 188422 477654
rect 188186 477098 188422 477334
rect 188186 441418 188422 441654
rect 188186 441098 188422 441334
rect 188186 405418 188422 405654
rect 188186 405098 188422 405334
rect 188186 369418 188422 369654
rect 188186 369098 188422 369334
rect 188186 333418 188422 333654
rect 188186 333098 188422 333334
rect 188186 297418 188422 297654
rect 188186 297098 188422 297334
rect 188186 261418 188422 261654
rect 188186 261098 188422 261334
rect 188186 225418 188422 225654
rect 188186 225098 188422 225334
rect 188186 189418 188422 189654
rect 188186 189098 188422 189334
rect 188186 153418 188422 153654
rect 188186 153098 188422 153334
rect 188186 117418 188422 117654
rect 188186 117098 188422 117334
rect 188186 81418 188422 81654
rect 188186 81098 188422 81334
rect 188186 45418 188422 45654
rect 188186 45098 188422 45334
rect 188186 9418 188422 9654
rect 188186 9098 188422 9334
rect 188186 -4342 188422 -4106
rect 188186 -4662 188422 -4426
rect 209786 711182 210022 711418
rect 209786 710862 210022 711098
rect 206186 709302 206422 709538
rect 206186 708982 206422 709218
rect 202586 707422 202822 707658
rect 202586 707102 202822 707338
rect 191786 697018 192022 697254
rect 191786 696698 192022 696934
rect 191786 661018 192022 661254
rect 191786 660698 192022 660934
rect 191786 625018 192022 625254
rect 191786 624698 192022 624934
rect 191786 589018 192022 589254
rect 191786 588698 192022 588934
rect 191786 553018 192022 553254
rect 191786 552698 192022 552934
rect 191786 517018 192022 517254
rect 191786 516698 192022 516934
rect 191786 481018 192022 481254
rect 191786 480698 192022 480934
rect 191786 445018 192022 445254
rect 191786 444698 192022 444934
rect 191786 409018 192022 409254
rect 191786 408698 192022 408934
rect 191786 373018 192022 373254
rect 191786 372698 192022 372934
rect 191786 337018 192022 337254
rect 191786 336698 192022 336934
rect 191786 301018 192022 301254
rect 191786 300698 192022 300934
rect 191786 265018 192022 265254
rect 191786 264698 192022 264934
rect 191786 229018 192022 229254
rect 191786 228698 192022 228934
rect 191786 193018 192022 193254
rect 191786 192698 192022 192934
rect 191786 157018 192022 157254
rect 191786 156698 192022 156934
rect 191786 121018 192022 121254
rect 191786 120698 192022 120934
rect 191786 85018 192022 85254
rect 191786 84698 192022 84934
rect 191786 49018 192022 49254
rect 191786 48698 192022 48934
rect 191786 13018 192022 13254
rect 191786 12698 192022 12934
rect 173786 -7162 174022 -6926
rect 173786 -7482 174022 -7246
rect 198986 705542 199222 705778
rect 198986 705222 199222 705458
rect 198986 668218 199222 668454
rect 198986 667898 199222 668134
rect 198986 632218 199222 632454
rect 198986 631898 199222 632134
rect 198986 596218 199222 596454
rect 198986 595898 199222 596134
rect 198986 560218 199222 560454
rect 198986 559898 199222 560134
rect 198986 524218 199222 524454
rect 198986 523898 199222 524134
rect 198986 488218 199222 488454
rect 198986 487898 199222 488134
rect 198986 452218 199222 452454
rect 198986 451898 199222 452134
rect 198986 416218 199222 416454
rect 198986 415898 199222 416134
rect 198986 380218 199222 380454
rect 198986 379898 199222 380134
rect 198986 344218 199222 344454
rect 198986 343898 199222 344134
rect 198986 308218 199222 308454
rect 198986 307898 199222 308134
rect 198986 272218 199222 272454
rect 198986 271898 199222 272134
rect 198986 236218 199222 236454
rect 198986 235898 199222 236134
rect 198986 200218 199222 200454
rect 198986 199898 199222 200134
rect 198986 164218 199222 164454
rect 198986 163898 199222 164134
rect 198986 128218 199222 128454
rect 198986 127898 199222 128134
rect 198986 92218 199222 92454
rect 198986 91898 199222 92134
rect 198986 56218 199222 56454
rect 198986 55898 199222 56134
rect 198986 20218 199222 20454
rect 198986 19898 199222 20134
rect 198986 -1522 199222 -1286
rect 198986 -1842 199222 -1606
rect 202586 671818 202822 672054
rect 202586 671498 202822 671734
rect 202586 635818 202822 636054
rect 202586 635498 202822 635734
rect 202586 599818 202822 600054
rect 202586 599498 202822 599734
rect 202586 563818 202822 564054
rect 202586 563498 202822 563734
rect 202586 527818 202822 528054
rect 202586 527498 202822 527734
rect 202586 491818 202822 492054
rect 202586 491498 202822 491734
rect 202586 455818 202822 456054
rect 202586 455498 202822 455734
rect 202586 419818 202822 420054
rect 202586 419498 202822 419734
rect 202586 383818 202822 384054
rect 202586 383498 202822 383734
rect 202586 347818 202822 348054
rect 202586 347498 202822 347734
rect 202586 311818 202822 312054
rect 202586 311498 202822 311734
rect 202586 275818 202822 276054
rect 202586 275498 202822 275734
rect 202586 239818 202822 240054
rect 202586 239498 202822 239734
rect 202586 203818 202822 204054
rect 202586 203498 202822 203734
rect 202586 167818 202822 168054
rect 202586 167498 202822 167734
rect 202586 131818 202822 132054
rect 202586 131498 202822 131734
rect 202586 95818 202822 96054
rect 202586 95498 202822 95734
rect 202586 59818 202822 60054
rect 202586 59498 202822 59734
rect 202586 23818 202822 24054
rect 202586 23498 202822 23734
rect 202586 -3402 202822 -3166
rect 202586 -3722 202822 -3486
rect 206186 675418 206422 675654
rect 206186 675098 206422 675334
rect 206186 639418 206422 639654
rect 206186 639098 206422 639334
rect 206186 603418 206422 603654
rect 206186 603098 206422 603334
rect 206186 567418 206422 567654
rect 206186 567098 206422 567334
rect 206186 531418 206422 531654
rect 206186 531098 206422 531334
rect 206186 495418 206422 495654
rect 206186 495098 206422 495334
rect 206186 459418 206422 459654
rect 206186 459098 206422 459334
rect 206186 423418 206422 423654
rect 206186 423098 206422 423334
rect 206186 387418 206422 387654
rect 206186 387098 206422 387334
rect 206186 351418 206422 351654
rect 206186 351098 206422 351334
rect 206186 315418 206422 315654
rect 206186 315098 206422 315334
rect 206186 279418 206422 279654
rect 206186 279098 206422 279334
rect 206186 243418 206422 243654
rect 206186 243098 206422 243334
rect 206186 207418 206422 207654
rect 206186 207098 206422 207334
rect 206186 171418 206422 171654
rect 206186 171098 206422 171334
rect 206186 135418 206422 135654
rect 206186 135098 206422 135334
rect 206186 99418 206422 99654
rect 206186 99098 206422 99334
rect 206186 63418 206422 63654
rect 206186 63098 206422 63334
rect 206186 27418 206422 27654
rect 206186 27098 206422 27334
rect 206186 -5282 206422 -5046
rect 206186 -5602 206422 -5366
rect 227786 710242 228022 710478
rect 227786 709922 228022 710158
rect 224186 708362 224422 708598
rect 224186 708042 224422 708278
rect 220586 706482 220822 706718
rect 220586 706162 220822 706398
rect 209786 679018 210022 679254
rect 209786 678698 210022 678934
rect 209786 643018 210022 643254
rect 209786 642698 210022 642934
rect 209786 607018 210022 607254
rect 209786 606698 210022 606934
rect 209786 571018 210022 571254
rect 209786 570698 210022 570934
rect 209786 535018 210022 535254
rect 209786 534698 210022 534934
rect 209786 499018 210022 499254
rect 209786 498698 210022 498934
rect 209786 463018 210022 463254
rect 209786 462698 210022 462934
rect 209786 427018 210022 427254
rect 209786 426698 210022 426934
rect 209786 391018 210022 391254
rect 209786 390698 210022 390934
rect 209786 355018 210022 355254
rect 209786 354698 210022 354934
rect 209786 319018 210022 319254
rect 209786 318698 210022 318934
rect 209786 283018 210022 283254
rect 209786 282698 210022 282934
rect 209786 247018 210022 247254
rect 209786 246698 210022 246934
rect 209786 211018 210022 211254
rect 209786 210698 210022 210934
rect 209786 175018 210022 175254
rect 209786 174698 210022 174934
rect 209786 139018 210022 139254
rect 209786 138698 210022 138934
rect 209786 103018 210022 103254
rect 209786 102698 210022 102934
rect 209786 67018 210022 67254
rect 209786 66698 210022 66934
rect 209786 31018 210022 31254
rect 209786 30698 210022 30934
rect 191786 -6222 192022 -5986
rect 191786 -6542 192022 -6306
rect 216986 704602 217222 704838
rect 216986 704282 217222 704518
rect 216986 686218 217222 686454
rect 216986 685898 217222 686134
rect 216986 650218 217222 650454
rect 216986 649898 217222 650134
rect 216986 614218 217222 614454
rect 216986 613898 217222 614134
rect 216986 578218 217222 578454
rect 216986 577898 217222 578134
rect 216986 542218 217222 542454
rect 216986 541898 217222 542134
rect 216986 506218 217222 506454
rect 216986 505898 217222 506134
rect 216986 470218 217222 470454
rect 216986 469898 217222 470134
rect 216986 434218 217222 434454
rect 216986 433898 217222 434134
rect 216986 398218 217222 398454
rect 216986 397898 217222 398134
rect 216986 362218 217222 362454
rect 216986 361898 217222 362134
rect 216986 326218 217222 326454
rect 216986 325898 217222 326134
rect 216986 290218 217222 290454
rect 216986 289898 217222 290134
rect 216986 254218 217222 254454
rect 216986 253898 217222 254134
rect 216986 218218 217222 218454
rect 216986 217898 217222 218134
rect 216986 182218 217222 182454
rect 216986 181898 217222 182134
rect 216986 146218 217222 146454
rect 216986 145898 217222 146134
rect 216986 110218 217222 110454
rect 216986 109898 217222 110134
rect 216986 74218 217222 74454
rect 216986 73898 217222 74134
rect 216986 38218 217222 38454
rect 216986 37898 217222 38134
rect 216986 2218 217222 2454
rect 216986 1898 217222 2134
rect 216986 -582 217222 -346
rect 216986 -902 217222 -666
rect 220586 689818 220822 690054
rect 220586 689498 220822 689734
rect 220586 653818 220822 654054
rect 220586 653498 220822 653734
rect 220586 617818 220822 618054
rect 220586 617498 220822 617734
rect 220586 581818 220822 582054
rect 220586 581498 220822 581734
rect 220586 545818 220822 546054
rect 220586 545498 220822 545734
rect 220586 509818 220822 510054
rect 220586 509498 220822 509734
rect 220586 473818 220822 474054
rect 220586 473498 220822 473734
rect 220586 437818 220822 438054
rect 220586 437498 220822 437734
rect 220586 401818 220822 402054
rect 220586 401498 220822 401734
rect 220586 365818 220822 366054
rect 220586 365498 220822 365734
rect 220586 329818 220822 330054
rect 220586 329498 220822 329734
rect 220586 293818 220822 294054
rect 220586 293498 220822 293734
rect 220586 257818 220822 258054
rect 220586 257498 220822 257734
rect 220586 221818 220822 222054
rect 220586 221498 220822 221734
rect 220586 185818 220822 186054
rect 220586 185498 220822 185734
rect 220586 149818 220822 150054
rect 220586 149498 220822 149734
rect 220586 113818 220822 114054
rect 220586 113498 220822 113734
rect 220586 77818 220822 78054
rect 220586 77498 220822 77734
rect 220586 41818 220822 42054
rect 220586 41498 220822 41734
rect 220586 5818 220822 6054
rect 220586 5498 220822 5734
rect 220586 -2462 220822 -2226
rect 220586 -2782 220822 -2546
rect 224186 693418 224422 693654
rect 224186 693098 224422 693334
rect 224186 657418 224422 657654
rect 224186 657098 224422 657334
rect 224186 621418 224422 621654
rect 224186 621098 224422 621334
rect 224186 585418 224422 585654
rect 224186 585098 224422 585334
rect 224186 549418 224422 549654
rect 224186 549098 224422 549334
rect 224186 513418 224422 513654
rect 224186 513098 224422 513334
rect 224186 477418 224422 477654
rect 224186 477098 224422 477334
rect 224186 441418 224422 441654
rect 224186 441098 224422 441334
rect 224186 405418 224422 405654
rect 224186 405098 224422 405334
rect 224186 369418 224422 369654
rect 224186 369098 224422 369334
rect 224186 333418 224422 333654
rect 224186 333098 224422 333334
rect 224186 297418 224422 297654
rect 224186 297098 224422 297334
rect 224186 261418 224422 261654
rect 224186 261098 224422 261334
rect 224186 225418 224422 225654
rect 224186 225098 224422 225334
rect 224186 189418 224422 189654
rect 224186 189098 224422 189334
rect 224186 153418 224422 153654
rect 224186 153098 224422 153334
rect 224186 117418 224422 117654
rect 224186 117098 224422 117334
rect 224186 81418 224422 81654
rect 224186 81098 224422 81334
rect 224186 45418 224422 45654
rect 224186 45098 224422 45334
rect 224186 9418 224422 9654
rect 224186 9098 224422 9334
rect 224186 -4342 224422 -4106
rect 224186 -4662 224422 -4426
rect 245786 711182 246022 711418
rect 245786 710862 246022 711098
rect 242186 709302 242422 709538
rect 242186 708982 242422 709218
rect 238586 707422 238822 707658
rect 238586 707102 238822 707338
rect 227786 697018 228022 697254
rect 227786 696698 228022 696934
rect 227786 661018 228022 661254
rect 227786 660698 228022 660934
rect 227786 625018 228022 625254
rect 227786 624698 228022 624934
rect 227786 589018 228022 589254
rect 227786 588698 228022 588934
rect 227786 553018 228022 553254
rect 227786 552698 228022 552934
rect 227786 517018 228022 517254
rect 227786 516698 228022 516934
rect 227786 481018 228022 481254
rect 227786 480698 228022 480934
rect 227786 445018 228022 445254
rect 227786 444698 228022 444934
rect 227786 409018 228022 409254
rect 227786 408698 228022 408934
rect 227786 373018 228022 373254
rect 227786 372698 228022 372934
rect 227786 337018 228022 337254
rect 227786 336698 228022 336934
rect 227786 301018 228022 301254
rect 227786 300698 228022 300934
rect 227786 265018 228022 265254
rect 227786 264698 228022 264934
rect 227786 229018 228022 229254
rect 227786 228698 228022 228934
rect 227786 193018 228022 193254
rect 227786 192698 228022 192934
rect 227786 157018 228022 157254
rect 227786 156698 228022 156934
rect 227786 121018 228022 121254
rect 227786 120698 228022 120934
rect 227786 85018 228022 85254
rect 227786 84698 228022 84934
rect 227786 49018 228022 49254
rect 227786 48698 228022 48934
rect 227786 13018 228022 13254
rect 227786 12698 228022 12934
rect 209786 -7162 210022 -6926
rect 209786 -7482 210022 -7246
rect 234986 705542 235222 705778
rect 234986 705222 235222 705458
rect 234986 668218 235222 668454
rect 234986 667898 235222 668134
rect 234986 632218 235222 632454
rect 234986 631898 235222 632134
rect 234986 596218 235222 596454
rect 234986 595898 235222 596134
rect 234986 560218 235222 560454
rect 234986 559898 235222 560134
rect 234986 524218 235222 524454
rect 234986 523898 235222 524134
rect 234986 488218 235222 488454
rect 234986 487898 235222 488134
rect 234986 452218 235222 452454
rect 234986 451898 235222 452134
rect 234986 416218 235222 416454
rect 234986 415898 235222 416134
rect 234986 380218 235222 380454
rect 234986 379898 235222 380134
rect 234986 344218 235222 344454
rect 234986 343898 235222 344134
rect 234986 308218 235222 308454
rect 234986 307898 235222 308134
rect 234986 272218 235222 272454
rect 234986 271898 235222 272134
rect 234986 236218 235222 236454
rect 234986 235898 235222 236134
rect 234986 200218 235222 200454
rect 234986 199898 235222 200134
rect 234986 164218 235222 164454
rect 234986 163898 235222 164134
rect 234986 128218 235222 128454
rect 234986 127898 235222 128134
rect 234986 92218 235222 92454
rect 234986 91898 235222 92134
rect 234986 56218 235222 56454
rect 234986 55898 235222 56134
rect 234986 20218 235222 20454
rect 234986 19898 235222 20134
rect 234986 -1522 235222 -1286
rect 234986 -1842 235222 -1606
rect 238586 671818 238822 672054
rect 238586 671498 238822 671734
rect 238586 635818 238822 636054
rect 238586 635498 238822 635734
rect 238586 599818 238822 600054
rect 238586 599498 238822 599734
rect 238586 563818 238822 564054
rect 238586 563498 238822 563734
rect 238586 527818 238822 528054
rect 238586 527498 238822 527734
rect 238586 491818 238822 492054
rect 238586 491498 238822 491734
rect 238586 455818 238822 456054
rect 238586 455498 238822 455734
rect 238586 419818 238822 420054
rect 238586 419498 238822 419734
rect 238586 383818 238822 384054
rect 238586 383498 238822 383734
rect 238586 347818 238822 348054
rect 238586 347498 238822 347734
rect 238586 311818 238822 312054
rect 238586 311498 238822 311734
rect 238586 275818 238822 276054
rect 238586 275498 238822 275734
rect 238586 239818 238822 240054
rect 238586 239498 238822 239734
rect 238586 203818 238822 204054
rect 238586 203498 238822 203734
rect 238586 167818 238822 168054
rect 238586 167498 238822 167734
rect 238586 131818 238822 132054
rect 238586 131498 238822 131734
rect 238586 95818 238822 96054
rect 238586 95498 238822 95734
rect 238586 59818 238822 60054
rect 238586 59498 238822 59734
rect 238586 23818 238822 24054
rect 238586 23498 238822 23734
rect 238586 -3402 238822 -3166
rect 238586 -3722 238822 -3486
rect 242186 675418 242422 675654
rect 242186 675098 242422 675334
rect 242186 639418 242422 639654
rect 242186 639098 242422 639334
rect 242186 603418 242422 603654
rect 242186 603098 242422 603334
rect 242186 567418 242422 567654
rect 242186 567098 242422 567334
rect 242186 531418 242422 531654
rect 242186 531098 242422 531334
rect 242186 495418 242422 495654
rect 242186 495098 242422 495334
rect 242186 459418 242422 459654
rect 242186 459098 242422 459334
rect 242186 423418 242422 423654
rect 242186 423098 242422 423334
rect 242186 387418 242422 387654
rect 242186 387098 242422 387334
rect 242186 351418 242422 351654
rect 242186 351098 242422 351334
rect 242186 315418 242422 315654
rect 242186 315098 242422 315334
rect 242186 279418 242422 279654
rect 242186 279098 242422 279334
rect 242186 243418 242422 243654
rect 242186 243098 242422 243334
rect 242186 207418 242422 207654
rect 242186 207098 242422 207334
rect 242186 171418 242422 171654
rect 242186 171098 242422 171334
rect 242186 135418 242422 135654
rect 242186 135098 242422 135334
rect 242186 99418 242422 99654
rect 242186 99098 242422 99334
rect 242186 63418 242422 63654
rect 242186 63098 242422 63334
rect 242186 27418 242422 27654
rect 242186 27098 242422 27334
rect 242186 -5282 242422 -5046
rect 242186 -5602 242422 -5366
rect 263786 710242 264022 710478
rect 263786 709922 264022 710158
rect 260186 708362 260422 708598
rect 260186 708042 260422 708278
rect 256586 706482 256822 706718
rect 256586 706162 256822 706398
rect 245786 679018 246022 679254
rect 245786 678698 246022 678934
rect 245786 643018 246022 643254
rect 245786 642698 246022 642934
rect 245786 607018 246022 607254
rect 245786 606698 246022 606934
rect 245786 571018 246022 571254
rect 245786 570698 246022 570934
rect 245786 535018 246022 535254
rect 245786 534698 246022 534934
rect 245786 499018 246022 499254
rect 245786 498698 246022 498934
rect 245786 463018 246022 463254
rect 245786 462698 246022 462934
rect 245786 427018 246022 427254
rect 245786 426698 246022 426934
rect 245786 391018 246022 391254
rect 245786 390698 246022 390934
rect 245786 355018 246022 355254
rect 245786 354698 246022 354934
rect 245786 319018 246022 319254
rect 245786 318698 246022 318934
rect 245786 283018 246022 283254
rect 245786 282698 246022 282934
rect 245786 247018 246022 247254
rect 245786 246698 246022 246934
rect 245786 211018 246022 211254
rect 245786 210698 246022 210934
rect 245786 175018 246022 175254
rect 245786 174698 246022 174934
rect 245786 139018 246022 139254
rect 245786 138698 246022 138934
rect 245786 103018 246022 103254
rect 245786 102698 246022 102934
rect 245786 67018 246022 67254
rect 245786 66698 246022 66934
rect 245786 31018 246022 31254
rect 245786 30698 246022 30934
rect 227786 -6222 228022 -5986
rect 227786 -6542 228022 -6306
rect 252986 704602 253222 704838
rect 252986 704282 253222 704518
rect 252986 686218 253222 686454
rect 252986 685898 253222 686134
rect 252986 650218 253222 650454
rect 252986 649898 253222 650134
rect 252986 614218 253222 614454
rect 252986 613898 253222 614134
rect 252986 578218 253222 578454
rect 252986 577898 253222 578134
rect 252986 542218 253222 542454
rect 252986 541898 253222 542134
rect 252986 506218 253222 506454
rect 252986 505898 253222 506134
rect 256586 689818 256822 690054
rect 256586 689498 256822 689734
rect 256586 653818 256822 654054
rect 256586 653498 256822 653734
rect 256586 617818 256822 618054
rect 256586 617498 256822 617734
rect 256586 581818 256822 582054
rect 256586 581498 256822 581734
rect 256586 545818 256822 546054
rect 256586 545498 256822 545734
rect 256586 509818 256822 510054
rect 256586 509498 256822 509734
rect 260186 693418 260422 693654
rect 260186 693098 260422 693334
rect 260186 657418 260422 657654
rect 260186 657098 260422 657334
rect 260186 621418 260422 621654
rect 260186 621098 260422 621334
rect 260186 585418 260422 585654
rect 260186 585098 260422 585334
rect 260186 549418 260422 549654
rect 260186 549098 260422 549334
rect 260186 513418 260422 513654
rect 260186 513098 260422 513334
rect 281786 711182 282022 711418
rect 281786 710862 282022 711098
rect 278186 709302 278422 709538
rect 278186 708982 278422 709218
rect 274586 707422 274822 707658
rect 274586 707102 274822 707338
rect 263786 697018 264022 697254
rect 263786 696698 264022 696934
rect 263786 661018 264022 661254
rect 263786 660698 264022 660934
rect 263786 625018 264022 625254
rect 263786 624698 264022 624934
rect 263786 589018 264022 589254
rect 263786 588698 264022 588934
rect 263786 553018 264022 553254
rect 263786 552698 264022 552934
rect 263786 517018 264022 517254
rect 263786 516698 264022 516934
rect 270986 705542 271222 705778
rect 270986 705222 271222 705458
rect 270986 668218 271222 668454
rect 270986 667898 271222 668134
rect 270986 632218 271222 632454
rect 270986 631898 271222 632134
rect 270986 596218 271222 596454
rect 270986 595898 271222 596134
rect 270986 560218 271222 560454
rect 270986 559898 271222 560134
rect 270986 524218 271222 524454
rect 270986 523898 271222 524134
rect 270986 488218 271222 488454
rect 270986 487898 271222 488134
rect 274586 671818 274822 672054
rect 274586 671498 274822 671734
rect 274586 635818 274822 636054
rect 274586 635498 274822 635734
rect 274586 599818 274822 600054
rect 274586 599498 274822 599734
rect 274586 563818 274822 564054
rect 274586 563498 274822 563734
rect 274586 527818 274822 528054
rect 274586 527498 274822 527734
rect 274586 491818 274822 492054
rect 274586 491498 274822 491734
rect 278186 675418 278422 675654
rect 278186 675098 278422 675334
rect 278186 639418 278422 639654
rect 278186 639098 278422 639334
rect 278186 603418 278422 603654
rect 278186 603098 278422 603334
rect 278186 567418 278422 567654
rect 278186 567098 278422 567334
rect 278186 531418 278422 531654
rect 278186 531098 278422 531334
rect 278186 495418 278422 495654
rect 278186 495098 278422 495334
rect 299786 710242 300022 710478
rect 299786 709922 300022 710158
rect 296186 708362 296422 708598
rect 296186 708042 296422 708278
rect 292586 706482 292822 706718
rect 292586 706162 292822 706398
rect 281786 679018 282022 679254
rect 281786 678698 282022 678934
rect 281786 643018 282022 643254
rect 281786 642698 282022 642934
rect 281786 607018 282022 607254
rect 281786 606698 282022 606934
rect 281786 571018 282022 571254
rect 281786 570698 282022 570934
rect 281786 535018 282022 535254
rect 281786 534698 282022 534934
rect 281786 499018 282022 499254
rect 281786 498698 282022 498934
rect 288986 704602 289222 704838
rect 288986 704282 289222 704518
rect 288986 686218 289222 686454
rect 288986 685898 289222 686134
rect 288986 650218 289222 650454
rect 288986 649898 289222 650134
rect 288986 614218 289222 614454
rect 288986 613898 289222 614134
rect 288986 578218 289222 578454
rect 288986 577898 289222 578134
rect 288986 542218 289222 542454
rect 288986 541898 289222 542134
rect 288986 506218 289222 506454
rect 288986 505898 289222 506134
rect 292586 689818 292822 690054
rect 292586 689498 292822 689734
rect 292586 653818 292822 654054
rect 292586 653498 292822 653734
rect 292586 617818 292822 618054
rect 292586 617498 292822 617734
rect 292586 581818 292822 582054
rect 292586 581498 292822 581734
rect 292586 545818 292822 546054
rect 292586 545498 292822 545734
rect 292586 509818 292822 510054
rect 292586 509498 292822 509734
rect 296186 693418 296422 693654
rect 296186 693098 296422 693334
rect 296186 657418 296422 657654
rect 296186 657098 296422 657334
rect 296186 621418 296422 621654
rect 296186 621098 296422 621334
rect 317786 711182 318022 711418
rect 317786 710862 318022 711098
rect 314186 709302 314422 709538
rect 314186 708982 314422 709218
rect 310586 707422 310822 707658
rect 310586 707102 310822 707338
rect 299786 697018 300022 697254
rect 299786 696698 300022 696934
rect 299786 661018 300022 661254
rect 299786 660698 300022 660934
rect 299786 625018 300022 625254
rect 299786 624698 300022 624934
rect 306986 705542 307222 705778
rect 306986 705222 307222 705458
rect 306986 668218 307222 668454
rect 306986 667898 307222 668134
rect 306986 632218 307222 632454
rect 306986 631898 307222 632134
rect 310586 671818 310822 672054
rect 310586 671498 310822 671734
rect 310586 635818 310822 636054
rect 310586 635498 310822 635734
rect 314186 675418 314422 675654
rect 314186 675098 314422 675334
rect 314186 639418 314422 639654
rect 314186 639098 314422 639334
rect 335786 710242 336022 710478
rect 335786 709922 336022 710158
rect 332186 708362 332422 708598
rect 332186 708042 332422 708278
rect 328586 706482 328822 706718
rect 328586 706162 328822 706398
rect 317786 679018 318022 679254
rect 317786 678698 318022 678934
rect 317786 643018 318022 643254
rect 317786 642698 318022 642934
rect 324986 704602 325222 704838
rect 324986 704282 325222 704518
rect 324986 686218 325222 686454
rect 324986 685898 325222 686134
rect 324986 650218 325222 650454
rect 324986 649898 325222 650134
rect 328586 689818 328822 690054
rect 328586 689498 328822 689734
rect 328586 653818 328822 654054
rect 328586 653498 328822 653734
rect 328586 617818 328822 618054
rect 328586 617498 328822 617734
rect 332186 693418 332422 693654
rect 332186 693098 332422 693334
rect 332186 657418 332422 657654
rect 332186 657098 332422 657334
rect 332186 621418 332422 621654
rect 332186 621098 332422 621334
rect 353786 711182 354022 711418
rect 353786 710862 354022 711098
rect 350186 709302 350422 709538
rect 350186 708982 350422 709218
rect 346586 707422 346822 707658
rect 346586 707102 346822 707338
rect 335786 697018 336022 697254
rect 335786 696698 336022 696934
rect 335786 661018 336022 661254
rect 335786 660698 336022 660934
rect 335786 625018 336022 625254
rect 335786 624698 336022 624934
rect 342986 705542 343222 705778
rect 342986 705222 343222 705458
rect 342986 668218 343222 668454
rect 342986 667898 343222 668134
rect 342986 632218 343222 632454
rect 342986 631898 343222 632134
rect 346586 671818 346822 672054
rect 346586 671498 346822 671734
rect 346586 635818 346822 636054
rect 346586 635498 346822 635734
rect 350186 675418 350422 675654
rect 350186 675098 350422 675334
rect 350186 639418 350422 639654
rect 350186 639098 350422 639334
rect 371786 710242 372022 710478
rect 371786 709922 372022 710158
rect 368186 708362 368422 708598
rect 368186 708042 368422 708278
rect 364586 706482 364822 706718
rect 364586 706162 364822 706398
rect 353786 679018 354022 679254
rect 353786 678698 354022 678934
rect 353786 643018 354022 643254
rect 353786 642698 354022 642934
rect 360986 704602 361222 704838
rect 360986 704282 361222 704518
rect 360986 686218 361222 686454
rect 360986 685898 361222 686134
rect 360986 650218 361222 650454
rect 360986 649898 361222 650134
rect 364586 689818 364822 690054
rect 364586 689498 364822 689734
rect 364586 653818 364822 654054
rect 364586 653498 364822 653734
rect 364586 617818 364822 618054
rect 364586 617498 364822 617734
rect 368186 693418 368422 693654
rect 368186 693098 368422 693334
rect 368186 657418 368422 657654
rect 368186 657098 368422 657334
rect 368186 621418 368422 621654
rect 368186 621098 368422 621334
rect 389786 711182 390022 711418
rect 389786 710862 390022 711098
rect 386186 709302 386422 709538
rect 386186 708982 386422 709218
rect 382586 707422 382822 707658
rect 382586 707102 382822 707338
rect 371786 697018 372022 697254
rect 371786 696698 372022 696934
rect 371786 661018 372022 661254
rect 371786 660698 372022 660934
rect 371786 625018 372022 625254
rect 371786 624698 372022 624934
rect 378986 705542 379222 705778
rect 378986 705222 379222 705458
rect 378986 668218 379222 668454
rect 378986 667898 379222 668134
rect 378986 632218 379222 632454
rect 378986 631898 379222 632134
rect 382586 671818 382822 672054
rect 382586 671498 382822 671734
rect 382586 635818 382822 636054
rect 382586 635498 382822 635734
rect 382586 599818 382822 600054
rect 382586 599498 382822 599734
rect 376982 596218 377218 596454
rect 376982 595898 377218 596134
rect 296186 585418 296422 585654
rect 296186 585098 296422 585334
rect 376536 578218 376772 578454
rect 376536 577898 376772 578134
rect 382586 563818 382822 564054
rect 382586 563498 382822 563734
rect 376982 560218 377218 560454
rect 376982 559898 377218 560134
rect 296186 549418 296422 549654
rect 296186 549098 296422 549334
rect 376536 542218 376772 542454
rect 376536 541898 376772 542134
rect 382586 527818 382822 528054
rect 382586 527498 382822 527734
rect 376982 524218 377218 524454
rect 376982 523898 377218 524134
rect 296186 513418 296422 513654
rect 296186 513098 296422 513334
rect 306986 488218 307222 488454
rect 306986 487898 307222 488134
rect 310586 491818 310822 492054
rect 310586 491498 310822 491734
rect 314186 495418 314422 495654
rect 314186 495098 314422 495334
rect 317786 499018 318022 499254
rect 317786 498698 318022 498934
rect 324986 506218 325222 506454
rect 324986 505898 325222 506134
rect 328586 509818 328822 510054
rect 328586 509498 328822 509734
rect 332186 513418 332422 513654
rect 332186 513098 332422 513334
rect 342986 488218 343222 488454
rect 342986 487898 343222 488134
rect 346586 491818 346822 492054
rect 346586 491498 346822 491734
rect 350186 495418 350422 495654
rect 350186 495098 350422 495334
rect 353786 499018 354022 499254
rect 353786 498698 354022 498934
rect 360986 506218 361222 506454
rect 360986 505898 361222 506134
rect 364586 509818 364822 510054
rect 364586 509498 364822 509734
rect 368186 513418 368422 513654
rect 368186 513098 368422 513334
rect 378986 488218 379222 488454
rect 378986 487898 379222 488134
rect 382586 491818 382822 492054
rect 382586 491498 382822 491734
rect 386186 675418 386422 675654
rect 386186 675098 386422 675334
rect 386186 639418 386422 639654
rect 386186 639098 386422 639334
rect 386186 603418 386422 603654
rect 386186 603098 386422 603334
rect 386186 567418 386422 567654
rect 386186 567098 386422 567334
rect 386186 531418 386422 531654
rect 386186 531098 386422 531334
rect 386186 495418 386422 495654
rect 386186 495098 386422 495334
rect 407786 710242 408022 710478
rect 407786 709922 408022 710158
rect 404186 708362 404422 708598
rect 404186 708042 404422 708278
rect 400586 706482 400822 706718
rect 400586 706162 400822 706398
rect 389786 679018 390022 679254
rect 389786 678698 390022 678934
rect 389786 643018 390022 643254
rect 389786 642698 390022 642934
rect 389786 607018 390022 607254
rect 389786 606698 390022 606934
rect 389786 571018 390022 571254
rect 389786 570698 390022 570934
rect 389786 535018 390022 535254
rect 389786 534698 390022 534934
rect 389786 499018 390022 499254
rect 389786 498698 390022 498934
rect 396986 704602 397222 704838
rect 396986 704282 397222 704518
rect 396986 686218 397222 686454
rect 396986 685898 397222 686134
rect 396986 650218 397222 650454
rect 396986 649898 397222 650134
rect 396986 614218 397222 614454
rect 396986 613898 397222 614134
rect 396986 578218 397222 578454
rect 396986 577898 397222 578134
rect 396986 542218 397222 542454
rect 396986 541898 397222 542134
rect 396986 506218 397222 506454
rect 396986 505898 397222 506134
rect 400586 689818 400822 690054
rect 400586 689498 400822 689734
rect 400586 653818 400822 654054
rect 400586 653498 400822 653734
rect 400586 617818 400822 618054
rect 400586 617498 400822 617734
rect 400586 581818 400822 582054
rect 400586 581498 400822 581734
rect 400586 545818 400822 546054
rect 400586 545498 400822 545734
rect 400586 509818 400822 510054
rect 400586 509498 400822 509734
rect 404186 693418 404422 693654
rect 404186 693098 404422 693334
rect 404186 657418 404422 657654
rect 404186 657098 404422 657334
rect 404186 621418 404422 621654
rect 404186 621098 404422 621334
rect 404186 585418 404422 585654
rect 404186 585098 404422 585334
rect 404186 549418 404422 549654
rect 404186 549098 404422 549334
rect 404186 513418 404422 513654
rect 404186 513098 404422 513334
rect 425786 711182 426022 711418
rect 425786 710862 426022 711098
rect 422186 709302 422422 709538
rect 422186 708982 422422 709218
rect 418586 707422 418822 707658
rect 418586 707102 418822 707338
rect 407786 697018 408022 697254
rect 407786 696698 408022 696934
rect 407786 661018 408022 661254
rect 407786 660698 408022 660934
rect 407786 625018 408022 625254
rect 407786 624698 408022 624934
rect 407786 589018 408022 589254
rect 407786 588698 408022 588934
rect 407786 553018 408022 553254
rect 407786 552698 408022 552934
rect 407786 517018 408022 517254
rect 407786 516698 408022 516934
rect 414986 705542 415222 705778
rect 414986 705222 415222 705458
rect 414986 668218 415222 668454
rect 414986 667898 415222 668134
rect 414986 632218 415222 632454
rect 414986 631898 415222 632134
rect 418586 671818 418822 672054
rect 418586 671498 418822 671734
rect 418586 635818 418822 636054
rect 418586 635498 418822 635734
rect 422186 675418 422422 675654
rect 422186 675098 422422 675334
rect 422186 639418 422422 639654
rect 422186 639098 422422 639334
rect 443786 710242 444022 710478
rect 443786 709922 444022 710158
rect 440186 708362 440422 708598
rect 440186 708042 440422 708278
rect 436586 706482 436822 706718
rect 436586 706162 436822 706398
rect 425786 679018 426022 679254
rect 425786 678698 426022 678934
rect 425786 643018 426022 643254
rect 425786 642698 426022 642934
rect 432986 704602 433222 704838
rect 432986 704282 433222 704518
rect 432986 686218 433222 686454
rect 432986 685898 433222 686134
rect 432986 650218 433222 650454
rect 432986 649898 433222 650134
rect 436586 689818 436822 690054
rect 436586 689498 436822 689734
rect 436586 653818 436822 654054
rect 436586 653498 436822 653734
rect 436586 617818 436822 618054
rect 436586 617498 436822 617734
rect 440186 693418 440422 693654
rect 440186 693098 440422 693334
rect 440186 657418 440422 657654
rect 440186 657098 440422 657334
rect 440186 621418 440422 621654
rect 440186 621098 440422 621334
rect 461786 711182 462022 711418
rect 461786 710862 462022 711098
rect 458186 709302 458422 709538
rect 458186 708982 458422 709218
rect 454586 707422 454822 707658
rect 454586 707102 454822 707338
rect 443786 697018 444022 697254
rect 443786 696698 444022 696934
rect 443786 661018 444022 661254
rect 443786 660698 444022 660934
rect 443786 625018 444022 625254
rect 443786 624698 444022 624934
rect 450986 705542 451222 705778
rect 450986 705222 451222 705458
rect 450986 668218 451222 668454
rect 450986 667898 451222 668134
rect 450986 632218 451222 632454
rect 450986 631898 451222 632134
rect 454586 671818 454822 672054
rect 454586 671498 454822 671734
rect 454586 635818 454822 636054
rect 454586 635498 454822 635734
rect 458186 675418 458422 675654
rect 458186 675098 458422 675334
rect 458186 639418 458422 639654
rect 458186 639098 458422 639334
rect 479786 710242 480022 710478
rect 479786 709922 480022 710158
rect 476186 708362 476422 708598
rect 476186 708042 476422 708278
rect 472586 706482 472822 706718
rect 472586 706162 472822 706398
rect 461786 679018 462022 679254
rect 461786 678698 462022 678934
rect 461786 643018 462022 643254
rect 461786 642698 462022 642934
rect 468986 704602 469222 704838
rect 468986 704282 469222 704518
rect 468986 686218 469222 686454
rect 468986 685898 469222 686134
rect 468986 650218 469222 650454
rect 468986 649898 469222 650134
rect 472586 689818 472822 690054
rect 472586 689498 472822 689734
rect 472586 653818 472822 654054
rect 472586 653498 472822 653734
rect 472586 617818 472822 618054
rect 472586 617498 472822 617734
rect 476186 693418 476422 693654
rect 476186 693098 476422 693334
rect 476186 657418 476422 657654
rect 476186 657098 476422 657334
rect 476186 621418 476422 621654
rect 476186 621098 476422 621334
rect 497786 711182 498022 711418
rect 497786 710862 498022 711098
rect 494186 709302 494422 709538
rect 494186 708982 494422 709218
rect 490586 707422 490822 707658
rect 490586 707102 490822 707338
rect 479786 697018 480022 697254
rect 479786 696698 480022 696934
rect 479786 661018 480022 661254
rect 479786 660698 480022 660934
rect 479786 625018 480022 625254
rect 479786 624698 480022 624934
rect 486986 705542 487222 705778
rect 486986 705222 487222 705458
rect 486986 668218 487222 668454
rect 486986 667898 487222 668134
rect 486986 632218 487222 632454
rect 486986 631898 487222 632134
rect 490586 671818 490822 672054
rect 490586 671498 490822 671734
rect 490586 635818 490822 636054
rect 490586 635498 490822 635734
rect 494186 675418 494422 675654
rect 494186 675098 494422 675334
rect 494186 639418 494422 639654
rect 494186 639098 494422 639334
rect 515786 710242 516022 710478
rect 515786 709922 516022 710158
rect 512186 708362 512422 708598
rect 512186 708042 512422 708278
rect 508586 706482 508822 706718
rect 508586 706162 508822 706398
rect 497786 679018 498022 679254
rect 497786 678698 498022 678934
rect 497786 643018 498022 643254
rect 497786 642698 498022 642934
rect 504986 704602 505222 704838
rect 504986 704282 505222 704518
rect 504986 686218 505222 686454
rect 504986 685898 505222 686134
rect 504986 650218 505222 650454
rect 504986 649898 505222 650134
rect 504986 614218 505222 614454
rect 504986 613898 505222 614134
rect 414986 596218 415222 596454
rect 414986 595898 415222 596134
rect 496982 596218 497218 596454
rect 496982 595898 497218 596134
rect 496536 578218 496772 578454
rect 496536 577898 496772 578134
rect 504986 578218 505222 578454
rect 504986 577898 505222 578134
rect 414986 560218 415222 560454
rect 414986 559898 415222 560134
rect 496982 560218 497218 560454
rect 496982 559898 497218 560134
rect 496536 542218 496772 542454
rect 496536 541898 496772 542134
rect 504986 542218 505222 542454
rect 504986 541898 505222 542134
rect 414986 524218 415222 524454
rect 414986 523898 415222 524134
rect 496982 524218 497218 524454
rect 496982 523898 497218 524134
rect 414986 488218 415222 488454
rect 414986 487898 415222 488134
rect 418586 491818 418822 492054
rect 418586 491498 418822 491734
rect 422186 495418 422422 495654
rect 422186 495098 422422 495334
rect 425786 499018 426022 499254
rect 425786 498698 426022 498934
rect 432986 506218 433222 506454
rect 432986 505898 433222 506134
rect 436586 509818 436822 510054
rect 436586 509498 436822 509734
rect 440186 513418 440422 513654
rect 440186 513098 440422 513334
rect 450986 488218 451222 488454
rect 450986 487898 451222 488134
rect 454586 491818 454822 492054
rect 454586 491498 454822 491734
rect 458186 495418 458422 495654
rect 458186 495098 458422 495334
rect 461786 499018 462022 499254
rect 461786 498698 462022 498934
rect 468986 506218 469222 506454
rect 468986 505898 469222 506134
rect 472586 509818 472822 510054
rect 472586 509498 472822 509734
rect 476186 513418 476422 513654
rect 476186 513098 476422 513334
rect 486986 488218 487222 488454
rect 486986 487898 487222 488134
rect 490586 491818 490822 492054
rect 490586 491498 490822 491734
rect 494186 495418 494422 495654
rect 494186 495098 494422 495334
rect 497786 499018 498022 499254
rect 497786 498698 498022 498934
rect 504986 506218 505222 506454
rect 504986 505898 505222 506134
rect 508586 689818 508822 690054
rect 508586 689498 508822 689734
rect 508586 653818 508822 654054
rect 508586 653498 508822 653734
rect 508586 617818 508822 618054
rect 508586 617498 508822 617734
rect 508586 581818 508822 582054
rect 508586 581498 508822 581734
rect 508586 545818 508822 546054
rect 508586 545498 508822 545734
rect 508586 509818 508822 510054
rect 508586 509498 508822 509734
rect 512186 693418 512422 693654
rect 512186 693098 512422 693334
rect 512186 657418 512422 657654
rect 512186 657098 512422 657334
rect 512186 621418 512422 621654
rect 512186 621098 512422 621334
rect 512186 585418 512422 585654
rect 512186 585098 512422 585334
rect 512186 549418 512422 549654
rect 512186 549098 512422 549334
rect 512186 513418 512422 513654
rect 512186 513098 512422 513334
rect 533786 711182 534022 711418
rect 533786 710862 534022 711098
rect 530186 709302 530422 709538
rect 530186 708982 530422 709218
rect 526586 707422 526822 707658
rect 526586 707102 526822 707338
rect 515786 697018 516022 697254
rect 515786 696698 516022 696934
rect 515786 661018 516022 661254
rect 515786 660698 516022 660934
rect 515786 625018 516022 625254
rect 515786 624698 516022 624934
rect 515786 589018 516022 589254
rect 515786 588698 516022 588934
rect 515786 553018 516022 553254
rect 515786 552698 516022 552934
rect 515786 517018 516022 517254
rect 515786 516698 516022 516934
rect 522986 705542 523222 705778
rect 522986 705222 523222 705458
rect 522986 668218 523222 668454
rect 522986 667898 523222 668134
rect 522986 632218 523222 632454
rect 522986 631898 523222 632134
rect 522986 596218 523222 596454
rect 522986 595898 523222 596134
rect 522986 560218 523222 560454
rect 522986 559898 523222 560134
rect 522986 524218 523222 524454
rect 522986 523898 523222 524134
rect 522986 488218 523222 488454
rect 522986 487898 523222 488134
rect 526586 671818 526822 672054
rect 526586 671498 526822 671734
rect 526586 635818 526822 636054
rect 526586 635498 526822 635734
rect 526586 599818 526822 600054
rect 526586 599498 526822 599734
rect 526586 563818 526822 564054
rect 526586 563498 526822 563734
rect 526586 527818 526822 528054
rect 526586 527498 526822 527734
rect 526586 491818 526822 492054
rect 526586 491498 526822 491734
rect 530186 675418 530422 675654
rect 530186 675098 530422 675334
rect 530186 639418 530422 639654
rect 530186 639098 530422 639334
rect 530186 603418 530422 603654
rect 530186 603098 530422 603334
rect 530186 567418 530422 567654
rect 530186 567098 530422 567334
rect 530186 531418 530422 531654
rect 530186 531098 530422 531334
rect 530186 495418 530422 495654
rect 530186 495098 530422 495334
rect 551786 710242 552022 710478
rect 551786 709922 552022 710158
rect 548186 708362 548422 708598
rect 548186 708042 548422 708278
rect 544586 706482 544822 706718
rect 544586 706162 544822 706398
rect 540986 704602 541222 704838
rect 540986 704282 541222 704518
rect 533786 679018 534022 679254
rect 533786 678698 534022 678934
rect 533786 643018 534022 643254
rect 533786 642698 534022 642934
rect 533786 607018 534022 607254
rect 533786 606698 534022 606934
rect 533786 571018 534022 571254
rect 533786 570698 534022 570934
rect 533786 535018 534022 535254
rect 533786 534698 534022 534934
rect 533786 499018 534022 499254
rect 533786 498698 534022 498934
rect 252986 470218 253222 470454
rect 252986 469898 253222 470134
rect 264250 470218 264486 470454
rect 264250 469898 264486 470134
rect 279610 452218 279846 452454
rect 279610 451898 279846 452134
rect 252986 434218 253222 434454
rect 252986 433898 253222 434134
rect 264250 434218 264486 434454
rect 264250 433898 264486 434134
rect 279610 416218 279846 416454
rect 279610 415898 279846 416134
rect 252986 398218 253222 398454
rect 252986 397898 253222 398134
rect 264250 398218 264486 398454
rect 264250 397898 264486 398134
rect 279610 380218 279846 380454
rect 279610 379898 279846 380134
rect 252986 362218 253222 362454
rect 252986 361898 253222 362134
rect 264250 362218 264486 362454
rect 264250 361898 264486 362134
rect 279610 344218 279846 344454
rect 279610 343898 279846 344134
rect 540986 686218 541222 686454
rect 540986 685898 541222 686134
rect 540986 650218 541222 650454
rect 540986 649898 541222 650134
rect 540986 614218 541222 614454
rect 540986 613898 541222 614134
rect 540986 578218 541222 578454
rect 540986 577898 541222 578134
rect 540986 542218 541222 542454
rect 540986 541898 541222 542134
rect 540986 506218 541222 506454
rect 540986 505898 541222 506134
rect 544586 689818 544822 690054
rect 544586 689498 544822 689734
rect 544586 653818 544822 654054
rect 544586 653498 544822 653734
rect 544586 617818 544822 618054
rect 544586 617498 544822 617734
rect 544586 581818 544822 582054
rect 544586 581498 544822 581734
rect 544586 545818 544822 546054
rect 544586 545498 544822 545734
rect 544586 509818 544822 510054
rect 544586 509498 544822 509734
rect 252986 326218 253222 326454
rect 252986 325898 253222 326134
rect 264250 326218 264486 326454
rect 264250 325898 264486 326134
rect 279610 308218 279846 308454
rect 279610 307898 279846 308134
rect 252986 290218 253222 290454
rect 252986 289898 253222 290134
rect 264250 290218 264486 290454
rect 264250 289898 264486 290134
rect 279610 272218 279846 272454
rect 279610 271898 279846 272134
rect 252986 254218 253222 254454
rect 252986 253898 253222 254134
rect 264250 254218 264486 254454
rect 264250 253898 264486 254134
rect 252986 218218 253222 218454
rect 252986 217898 253222 218134
rect 252986 182218 253222 182454
rect 252986 181898 253222 182134
rect 252986 146218 253222 146454
rect 252986 145898 253222 146134
rect 252986 110218 253222 110454
rect 252986 109898 253222 110134
rect 252986 74218 253222 74454
rect 252986 73898 253222 74134
rect 252986 38218 253222 38454
rect 252986 37898 253222 38134
rect 252986 2218 253222 2454
rect 252986 1898 253222 2134
rect 252986 -582 253222 -346
rect 252986 -902 253222 -666
rect 256586 221818 256822 222054
rect 256586 221498 256822 221734
rect 256586 185818 256822 186054
rect 256586 185498 256822 185734
rect 256586 149818 256822 150054
rect 256586 149498 256822 149734
rect 256586 113818 256822 114054
rect 256586 113498 256822 113734
rect 256586 77818 256822 78054
rect 256586 77498 256822 77734
rect 256586 41818 256822 42054
rect 256586 41498 256822 41734
rect 256586 5818 256822 6054
rect 256586 5498 256822 5734
rect 256586 -2462 256822 -2226
rect 256586 -2782 256822 -2546
rect 260186 225418 260422 225654
rect 260186 225098 260422 225334
rect 260186 189418 260422 189654
rect 260186 189098 260422 189334
rect 260186 153418 260422 153654
rect 260186 153098 260422 153334
rect 260186 117418 260422 117654
rect 260186 117098 260422 117334
rect 260186 81418 260422 81654
rect 260186 81098 260422 81334
rect 260186 45418 260422 45654
rect 260186 45098 260422 45334
rect 260186 9418 260422 9654
rect 260186 9098 260422 9334
rect 260186 -4342 260422 -4106
rect 260186 -4662 260422 -4426
rect 263786 229018 264022 229254
rect 263786 228698 264022 228934
rect 263786 193018 264022 193254
rect 263786 192698 264022 192934
rect 263786 157018 264022 157254
rect 263786 156698 264022 156934
rect 263786 121018 264022 121254
rect 263786 120698 264022 120934
rect 263786 85018 264022 85254
rect 263786 84698 264022 84934
rect 263786 49018 264022 49254
rect 263786 48698 264022 48934
rect 263786 13018 264022 13254
rect 263786 12698 264022 12934
rect 245786 -7162 246022 -6926
rect 245786 -7482 246022 -7246
rect 270986 236218 271222 236454
rect 270986 235898 271222 236134
rect 270986 200218 271222 200454
rect 270986 199898 271222 200134
rect 270986 164218 271222 164454
rect 270986 163898 271222 164134
rect 270986 128218 271222 128454
rect 270986 127898 271222 128134
rect 270986 92218 271222 92454
rect 270986 91898 271222 92134
rect 270986 56218 271222 56454
rect 270986 55898 271222 56134
rect 270986 20218 271222 20454
rect 270986 19898 271222 20134
rect 270986 -1522 271222 -1286
rect 270986 -1842 271222 -1606
rect 274586 203818 274822 204054
rect 274586 203498 274822 203734
rect 274586 167818 274822 168054
rect 274586 167498 274822 167734
rect 274586 131818 274822 132054
rect 274586 131498 274822 131734
rect 274586 95818 274822 96054
rect 274586 95498 274822 95734
rect 274586 59818 274822 60054
rect 274586 59498 274822 59734
rect 274586 23818 274822 24054
rect 274586 23498 274822 23734
rect 274586 -3402 274822 -3166
rect 274586 -3722 274822 -3486
rect 278186 207418 278422 207654
rect 278186 207098 278422 207334
rect 278186 171418 278422 171654
rect 278186 171098 278422 171334
rect 278186 135418 278422 135654
rect 278186 135098 278422 135334
rect 278186 99418 278422 99654
rect 278186 99098 278422 99334
rect 278186 63418 278422 63654
rect 278186 63098 278422 63334
rect 278186 27418 278422 27654
rect 278186 27098 278422 27334
rect 278186 -5282 278422 -5046
rect 278186 -5602 278422 -5366
rect 281786 211018 282022 211254
rect 281786 210698 282022 210934
rect 281786 175018 282022 175254
rect 281786 174698 282022 174934
rect 281786 139018 282022 139254
rect 281786 138698 282022 138934
rect 281786 103018 282022 103254
rect 281786 102698 282022 102934
rect 281786 67018 282022 67254
rect 281786 66698 282022 66934
rect 281786 31018 282022 31254
rect 281786 30698 282022 30934
rect 263786 -6222 264022 -5986
rect 263786 -6542 264022 -6306
rect 288986 218218 289222 218454
rect 288986 217898 289222 218134
rect 288986 182218 289222 182454
rect 288986 181898 289222 182134
rect 288986 146218 289222 146454
rect 288986 145898 289222 146134
rect 288986 110218 289222 110454
rect 288986 109898 289222 110134
rect 288986 74218 289222 74454
rect 288986 73898 289222 74134
rect 288986 38218 289222 38454
rect 288986 37898 289222 38134
rect 288986 2218 289222 2454
rect 288986 1898 289222 2134
rect 288986 -582 289222 -346
rect 288986 -902 289222 -666
rect 292586 221818 292822 222054
rect 292586 221498 292822 221734
rect 292586 185818 292822 186054
rect 292586 185498 292822 185734
rect 292586 149818 292822 150054
rect 292586 149498 292822 149734
rect 292586 113818 292822 114054
rect 292586 113498 292822 113734
rect 292586 77818 292822 78054
rect 292586 77498 292822 77734
rect 292586 41818 292822 42054
rect 292586 41498 292822 41734
rect 292586 5818 292822 6054
rect 292586 5498 292822 5734
rect 292586 -2462 292822 -2226
rect 292586 -2782 292822 -2546
rect 296186 225418 296422 225654
rect 296186 225098 296422 225334
rect 299786 229018 300022 229254
rect 299786 228698 300022 228934
rect 306986 236218 307222 236454
rect 306986 235898 307222 236134
rect 314186 207418 314422 207654
rect 314186 207098 314422 207334
rect 317786 211018 318022 211254
rect 317786 210698 318022 210934
rect 324986 218218 325222 218454
rect 324986 217898 325222 218134
rect 328586 221818 328822 222054
rect 328586 221498 328822 221734
rect 332186 225418 332422 225654
rect 332186 225098 332422 225334
rect 335786 229018 336022 229254
rect 335786 228698 336022 228934
rect 342986 236218 343222 236454
rect 342986 235898 343222 236134
rect 350186 207418 350422 207654
rect 350186 207098 350422 207334
rect 353786 211018 354022 211254
rect 353786 210698 354022 210934
rect 360986 218218 361222 218454
rect 360986 217898 361222 218134
rect 364586 221818 364822 222054
rect 364586 221498 364822 221734
rect 368186 225418 368422 225654
rect 368186 225098 368422 225334
rect 371786 229018 372022 229254
rect 371786 228698 372022 228934
rect 378986 236218 379222 236454
rect 378986 235898 379222 236134
rect 382586 203818 382822 204054
rect 382586 203498 382822 203734
rect 296186 189418 296422 189654
rect 296186 189098 296422 189334
rect 300524 182218 300760 182454
rect 300524 181898 300760 182134
rect 382586 167818 382822 168054
rect 382586 167498 382822 167734
rect 300078 164218 300314 164454
rect 300078 163898 300314 164134
rect 296186 153418 296422 153654
rect 296186 153098 296422 153334
rect 300524 146218 300760 146454
rect 300524 145898 300760 146134
rect 382586 131818 382822 132054
rect 382586 131498 382822 131734
rect 300078 128218 300314 128454
rect 300078 127898 300314 128134
rect 296186 117418 296422 117654
rect 296186 117098 296422 117334
rect 296186 81418 296422 81654
rect 296186 81098 296422 81334
rect 296186 45418 296422 45654
rect 296186 45098 296422 45334
rect 296186 9418 296422 9654
rect 296186 9098 296422 9334
rect 296186 -4342 296422 -4106
rect 296186 -4662 296422 -4426
rect 299786 85018 300022 85254
rect 299786 84698 300022 84934
rect 299786 49018 300022 49254
rect 299786 48698 300022 48934
rect 299786 13018 300022 13254
rect 299786 12698 300022 12934
rect 281786 -7162 282022 -6926
rect 281786 -7482 282022 -7246
rect 306986 92218 307222 92454
rect 306986 91898 307222 92134
rect 306986 56218 307222 56454
rect 306986 55898 307222 56134
rect 306986 20218 307222 20454
rect 306986 19898 307222 20134
rect 306986 -1522 307222 -1286
rect 306986 -1842 307222 -1606
rect 310586 95818 310822 96054
rect 310586 95498 310822 95734
rect 310586 59818 310822 60054
rect 310586 59498 310822 59734
rect 310586 23818 310822 24054
rect 310586 23498 310822 23734
rect 310586 -3402 310822 -3166
rect 310586 -3722 310822 -3486
rect 314186 99418 314422 99654
rect 314186 99098 314422 99334
rect 314186 63418 314422 63654
rect 314186 63098 314422 63334
rect 314186 27418 314422 27654
rect 314186 27098 314422 27334
rect 314186 -5282 314422 -5046
rect 314186 -5602 314422 -5366
rect 317786 103018 318022 103254
rect 317786 102698 318022 102934
rect 317786 67018 318022 67254
rect 317786 66698 318022 66934
rect 317786 31018 318022 31254
rect 317786 30698 318022 30934
rect 299786 -6222 300022 -5986
rect 299786 -6542 300022 -6306
rect 324986 74218 325222 74454
rect 324986 73898 325222 74134
rect 324986 38218 325222 38454
rect 324986 37898 325222 38134
rect 324986 2218 325222 2454
rect 324986 1898 325222 2134
rect 324986 -582 325222 -346
rect 324986 -902 325222 -666
rect 328586 77818 328822 78054
rect 328586 77498 328822 77734
rect 328586 41818 328822 42054
rect 328586 41498 328822 41734
rect 328586 5818 328822 6054
rect 328586 5498 328822 5734
rect 328586 -2462 328822 -2226
rect 328586 -2782 328822 -2546
rect 332186 81418 332422 81654
rect 332186 81098 332422 81334
rect 332186 45418 332422 45654
rect 332186 45098 332422 45334
rect 332186 9418 332422 9654
rect 332186 9098 332422 9334
rect 332186 -4342 332422 -4106
rect 332186 -4662 332422 -4426
rect 335786 85018 336022 85254
rect 335786 84698 336022 84934
rect 335786 49018 336022 49254
rect 335786 48698 336022 48934
rect 335786 13018 336022 13254
rect 335786 12698 336022 12934
rect 317786 -7162 318022 -6926
rect 317786 -7482 318022 -7246
rect 342986 92218 343222 92454
rect 342986 91898 343222 92134
rect 342986 56218 343222 56454
rect 342986 55898 343222 56134
rect 342986 20218 343222 20454
rect 342986 19898 343222 20134
rect 342986 -1522 343222 -1286
rect 342986 -1842 343222 -1606
rect 346586 95818 346822 96054
rect 346586 95498 346822 95734
rect 346586 59818 346822 60054
rect 346586 59498 346822 59734
rect 346586 23818 346822 24054
rect 346586 23498 346822 23734
rect 346586 -3402 346822 -3166
rect 346586 -3722 346822 -3486
rect 350186 99418 350422 99654
rect 350186 99098 350422 99334
rect 350186 63418 350422 63654
rect 350186 63098 350422 63334
rect 350186 27418 350422 27654
rect 350186 27098 350422 27334
rect 350186 -5282 350422 -5046
rect 350186 -5602 350422 -5366
rect 353786 103018 354022 103254
rect 353786 102698 354022 102934
rect 353786 67018 354022 67254
rect 353786 66698 354022 66934
rect 353786 31018 354022 31254
rect 353786 30698 354022 30934
rect 335786 -6222 336022 -5986
rect 335786 -6542 336022 -6306
rect 360986 74218 361222 74454
rect 360986 73898 361222 74134
rect 360986 38218 361222 38454
rect 360986 37898 361222 38134
rect 360986 2218 361222 2454
rect 360986 1898 361222 2134
rect 360986 -582 361222 -346
rect 360986 -902 361222 -666
rect 364586 77818 364822 78054
rect 364586 77498 364822 77734
rect 364586 41818 364822 42054
rect 364586 41498 364822 41734
rect 364586 5818 364822 6054
rect 364586 5498 364822 5734
rect 364586 -2462 364822 -2226
rect 364586 -2782 364822 -2546
rect 368186 81418 368422 81654
rect 368186 81098 368422 81334
rect 368186 45418 368422 45654
rect 368186 45098 368422 45334
rect 368186 9418 368422 9654
rect 368186 9098 368422 9334
rect 368186 -4342 368422 -4106
rect 368186 -4662 368422 -4426
rect 371786 85018 372022 85254
rect 371786 84698 372022 84934
rect 371786 49018 372022 49254
rect 371786 48698 372022 48934
rect 371786 13018 372022 13254
rect 371786 12698 372022 12934
rect 353786 -7162 354022 -6926
rect 353786 -7482 354022 -7246
rect 378986 92218 379222 92454
rect 378986 91898 379222 92134
rect 378986 56218 379222 56454
rect 378986 55898 379222 56134
rect 378986 20218 379222 20454
rect 378986 19898 379222 20134
rect 378986 -1522 379222 -1286
rect 378986 -1842 379222 -1606
rect 382586 95818 382822 96054
rect 382586 95498 382822 95734
rect 382586 59818 382822 60054
rect 382586 59498 382822 59734
rect 382586 23818 382822 24054
rect 382586 23498 382822 23734
rect 382586 -3402 382822 -3166
rect 382586 -3722 382822 -3486
rect 386186 207418 386422 207654
rect 386186 207098 386422 207334
rect 386186 171418 386422 171654
rect 386186 171098 386422 171334
rect 386186 135418 386422 135654
rect 386186 135098 386422 135334
rect 386186 99418 386422 99654
rect 386186 99098 386422 99334
rect 386186 63418 386422 63654
rect 386186 63098 386422 63334
rect 386186 27418 386422 27654
rect 386186 27098 386422 27334
rect 386186 -5282 386422 -5046
rect 386186 -5602 386422 -5366
rect 389786 211018 390022 211254
rect 389786 210698 390022 210934
rect 389786 175018 390022 175254
rect 389786 174698 390022 174934
rect 389786 139018 390022 139254
rect 389786 138698 390022 138934
rect 389786 103018 390022 103254
rect 389786 102698 390022 102934
rect 389786 67018 390022 67254
rect 389786 66698 390022 66934
rect 389786 31018 390022 31254
rect 389786 30698 390022 30934
rect 371786 -6222 372022 -5986
rect 371786 -6542 372022 -6306
rect 396986 218218 397222 218454
rect 396986 217898 397222 218134
rect 396986 182218 397222 182454
rect 396986 181898 397222 182134
rect 396986 146218 397222 146454
rect 396986 145898 397222 146134
rect 396986 110218 397222 110454
rect 396986 109898 397222 110134
rect 396986 74218 397222 74454
rect 396986 73898 397222 74134
rect 396986 38218 397222 38454
rect 396986 37898 397222 38134
rect 396986 2218 397222 2454
rect 396986 1898 397222 2134
rect 396986 -582 397222 -346
rect 396986 -902 397222 -666
rect 400586 221818 400822 222054
rect 400586 221498 400822 221734
rect 400586 185818 400822 186054
rect 400586 185498 400822 185734
rect 400586 149818 400822 150054
rect 400586 149498 400822 149734
rect 400586 113818 400822 114054
rect 400586 113498 400822 113734
rect 400586 77818 400822 78054
rect 400586 77498 400822 77734
rect 400586 41818 400822 42054
rect 400586 41498 400822 41734
rect 400586 5818 400822 6054
rect 400586 5498 400822 5734
rect 400586 -2462 400822 -2226
rect 400586 -2782 400822 -2546
rect 404186 225418 404422 225654
rect 404186 225098 404422 225334
rect 404186 189418 404422 189654
rect 404186 189098 404422 189334
rect 404186 153418 404422 153654
rect 404186 153098 404422 153334
rect 404186 117418 404422 117654
rect 404186 117098 404422 117334
rect 404186 81418 404422 81654
rect 404186 81098 404422 81334
rect 404186 45418 404422 45654
rect 404186 45098 404422 45334
rect 404186 9418 404422 9654
rect 404186 9098 404422 9334
rect 404186 -4342 404422 -4106
rect 404186 -4662 404422 -4426
rect 407786 229018 408022 229254
rect 407786 228698 408022 228934
rect 407786 193018 408022 193254
rect 407786 192698 408022 192934
rect 407786 157018 408022 157254
rect 407786 156698 408022 156934
rect 407786 121018 408022 121254
rect 407786 120698 408022 120934
rect 407786 85018 408022 85254
rect 407786 84698 408022 84934
rect 407786 49018 408022 49254
rect 407786 48698 408022 48934
rect 407786 13018 408022 13254
rect 407786 12698 408022 12934
rect 389786 -7162 390022 -6926
rect 389786 -7482 390022 -7246
rect 414986 236218 415222 236454
rect 414986 235898 415222 236134
rect 422186 207418 422422 207654
rect 422186 207098 422422 207334
rect 425786 211018 426022 211254
rect 425786 210698 426022 210934
rect 432986 218218 433222 218454
rect 432986 217898 433222 218134
rect 436586 221818 436822 222054
rect 436586 221498 436822 221734
rect 440186 225418 440422 225654
rect 440186 225098 440422 225334
rect 443786 229018 444022 229254
rect 443786 228698 444022 228934
rect 450986 236218 451222 236454
rect 450986 235898 451222 236134
rect 458186 207418 458422 207654
rect 458186 207098 458422 207334
rect 461786 211018 462022 211254
rect 461786 210698 462022 210934
rect 468986 218218 469222 218454
rect 468986 217898 469222 218134
rect 472586 221818 472822 222054
rect 472586 221498 472822 221734
rect 476186 225418 476422 225654
rect 476186 225098 476422 225334
rect 479786 229018 480022 229254
rect 479786 228698 480022 228934
rect 486986 236218 487222 236454
rect 486986 235898 487222 236134
rect 494186 207418 494422 207654
rect 494186 207098 494422 207334
rect 497786 211018 498022 211254
rect 497786 210698 498022 210934
rect 504986 218218 505222 218454
rect 504986 217898 505222 218134
rect 414986 200218 415222 200454
rect 414986 199898 415222 200134
rect 420524 182218 420760 182454
rect 420524 181898 420760 182134
rect 504986 182218 505222 182454
rect 504986 181898 505222 182134
rect 414986 164218 415222 164454
rect 414986 163898 415222 164134
rect 420078 164218 420314 164454
rect 420078 163898 420314 164134
rect 420524 146218 420760 146454
rect 420524 145898 420760 146134
rect 504986 146218 505222 146454
rect 504986 145898 505222 146134
rect 414986 128218 415222 128454
rect 414986 127898 415222 128134
rect 420078 128218 420314 128454
rect 420078 127898 420314 128134
rect 504986 110218 505222 110454
rect 504986 109898 505222 110134
rect 414986 92218 415222 92454
rect 414986 91898 415222 92134
rect 414986 56218 415222 56454
rect 414986 55898 415222 56134
rect 414986 20218 415222 20454
rect 414986 19898 415222 20134
rect 414986 -1522 415222 -1286
rect 414986 -1842 415222 -1606
rect 418586 95818 418822 96054
rect 418586 95498 418822 95734
rect 418586 59818 418822 60054
rect 418586 59498 418822 59734
rect 418586 23818 418822 24054
rect 418586 23498 418822 23734
rect 418586 -3402 418822 -3166
rect 418586 -3722 418822 -3486
rect 422186 99418 422422 99654
rect 422186 99098 422422 99334
rect 422186 63418 422422 63654
rect 422186 63098 422422 63334
rect 422186 27418 422422 27654
rect 422186 27098 422422 27334
rect 422186 -5282 422422 -5046
rect 422186 -5602 422422 -5366
rect 425786 103018 426022 103254
rect 425786 102698 426022 102934
rect 425786 67018 426022 67254
rect 425786 66698 426022 66934
rect 425786 31018 426022 31254
rect 425786 30698 426022 30934
rect 407786 -6222 408022 -5986
rect 407786 -6542 408022 -6306
rect 432986 74218 433222 74454
rect 432986 73898 433222 74134
rect 432986 38218 433222 38454
rect 432986 37898 433222 38134
rect 432986 2218 433222 2454
rect 432986 1898 433222 2134
rect 432986 -582 433222 -346
rect 432986 -902 433222 -666
rect 436586 77818 436822 78054
rect 436586 77498 436822 77734
rect 436586 41818 436822 42054
rect 436586 41498 436822 41734
rect 436586 5818 436822 6054
rect 436586 5498 436822 5734
rect 436586 -2462 436822 -2226
rect 436586 -2782 436822 -2546
rect 440186 81418 440422 81654
rect 440186 81098 440422 81334
rect 440186 45418 440422 45654
rect 440186 45098 440422 45334
rect 440186 9418 440422 9654
rect 440186 9098 440422 9334
rect 440186 -4342 440422 -4106
rect 440186 -4662 440422 -4426
rect 443786 85018 444022 85254
rect 443786 84698 444022 84934
rect 443786 49018 444022 49254
rect 443786 48698 444022 48934
rect 443786 13018 444022 13254
rect 443786 12698 444022 12934
rect 425786 -7162 426022 -6926
rect 425786 -7482 426022 -7246
rect 450986 92218 451222 92454
rect 450986 91898 451222 92134
rect 450986 56218 451222 56454
rect 450986 55898 451222 56134
rect 450986 20218 451222 20454
rect 450986 19898 451222 20134
rect 450986 -1522 451222 -1286
rect 450986 -1842 451222 -1606
rect 454586 95818 454822 96054
rect 454586 95498 454822 95734
rect 454586 59818 454822 60054
rect 454586 59498 454822 59734
rect 454586 23818 454822 24054
rect 454586 23498 454822 23734
rect 454586 -3402 454822 -3166
rect 454586 -3722 454822 -3486
rect 458186 99418 458422 99654
rect 458186 99098 458422 99334
rect 458186 63418 458422 63654
rect 458186 63098 458422 63334
rect 458186 27418 458422 27654
rect 458186 27098 458422 27334
rect 458186 -5282 458422 -5046
rect 458186 -5602 458422 -5366
rect 461786 103018 462022 103254
rect 461786 102698 462022 102934
rect 461786 67018 462022 67254
rect 461786 66698 462022 66934
rect 461786 31018 462022 31254
rect 461786 30698 462022 30934
rect 443786 -6222 444022 -5986
rect 443786 -6542 444022 -6306
rect 468986 74218 469222 74454
rect 468986 73898 469222 74134
rect 468986 38218 469222 38454
rect 468986 37898 469222 38134
rect 468986 2218 469222 2454
rect 468986 1898 469222 2134
rect 468986 -582 469222 -346
rect 468986 -902 469222 -666
rect 472586 77818 472822 78054
rect 472586 77498 472822 77734
rect 472586 41818 472822 42054
rect 472586 41498 472822 41734
rect 472586 5818 472822 6054
rect 472586 5498 472822 5734
rect 472586 -2462 472822 -2226
rect 472586 -2782 472822 -2546
rect 476186 81418 476422 81654
rect 476186 81098 476422 81334
rect 476186 45418 476422 45654
rect 476186 45098 476422 45334
rect 476186 9418 476422 9654
rect 476186 9098 476422 9334
rect 476186 -4342 476422 -4106
rect 476186 -4662 476422 -4426
rect 479786 85018 480022 85254
rect 479786 84698 480022 84934
rect 479786 49018 480022 49254
rect 479786 48698 480022 48934
rect 479786 13018 480022 13254
rect 479786 12698 480022 12934
rect 461786 -7162 462022 -6926
rect 461786 -7482 462022 -7246
rect 486986 92218 487222 92454
rect 486986 91898 487222 92134
rect 486986 56218 487222 56454
rect 486986 55898 487222 56134
rect 486986 20218 487222 20454
rect 486986 19898 487222 20134
rect 486986 -1522 487222 -1286
rect 486986 -1842 487222 -1606
rect 490586 95818 490822 96054
rect 490586 95498 490822 95734
rect 490586 59818 490822 60054
rect 490586 59498 490822 59734
rect 490586 23818 490822 24054
rect 490586 23498 490822 23734
rect 490586 -3402 490822 -3166
rect 490586 -3722 490822 -3486
rect 494186 99418 494422 99654
rect 494186 99098 494422 99334
rect 494186 63418 494422 63654
rect 494186 63098 494422 63334
rect 494186 27418 494422 27654
rect 494186 27098 494422 27334
rect 494186 -5282 494422 -5046
rect 494186 -5602 494422 -5366
rect 497786 103018 498022 103254
rect 497786 102698 498022 102934
rect 497786 67018 498022 67254
rect 497786 66698 498022 66934
rect 497786 31018 498022 31254
rect 497786 30698 498022 30934
rect 479786 -6222 480022 -5986
rect 479786 -6542 480022 -6306
rect 504986 74218 505222 74454
rect 504986 73898 505222 74134
rect 504986 38218 505222 38454
rect 504986 37898 505222 38134
rect 504986 2218 505222 2454
rect 504986 1898 505222 2134
rect 504986 -582 505222 -346
rect 504986 -902 505222 -666
rect 508586 221818 508822 222054
rect 508586 221498 508822 221734
rect 508586 185818 508822 186054
rect 508586 185498 508822 185734
rect 508586 149818 508822 150054
rect 508586 149498 508822 149734
rect 508586 113818 508822 114054
rect 508586 113498 508822 113734
rect 508586 77818 508822 78054
rect 508586 77498 508822 77734
rect 508586 41818 508822 42054
rect 508586 41498 508822 41734
rect 508586 5818 508822 6054
rect 508586 5498 508822 5734
rect 508586 -2462 508822 -2226
rect 508586 -2782 508822 -2546
rect 512186 225418 512422 225654
rect 512186 225098 512422 225334
rect 512186 189418 512422 189654
rect 512186 189098 512422 189334
rect 512186 153418 512422 153654
rect 512186 153098 512422 153334
rect 512186 117418 512422 117654
rect 512186 117098 512422 117334
rect 512186 81418 512422 81654
rect 512186 81098 512422 81334
rect 512186 45418 512422 45654
rect 512186 45098 512422 45334
rect 512186 9418 512422 9654
rect 512186 9098 512422 9334
rect 512186 -4342 512422 -4106
rect 512186 -4662 512422 -4426
rect 515786 229018 516022 229254
rect 515786 228698 516022 228934
rect 515786 193018 516022 193254
rect 515786 192698 516022 192934
rect 515786 157018 516022 157254
rect 515786 156698 516022 156934
rect 515786 121018 516022 121254
rect 515786 120698 516022 120934
rect 515786 85018 516022 85254
rect 515786 84698 516022 84934
rect 515786 49018 516022 49254
rect 515786 48698 516022 48934
rect 515786 13018 516022 13254
rect 515786 12698 516022 12934
rect 497786 -7162 498022 -6926
rect 497786 -7482 498022 -7246
rect 522986 236218 523222 236454
rect 522986 235898 523222 236134
rect 522986 200218 523222 200454
rect 522986 199898 523222 200134
rect 522986 164218 523222 164454
rect 522986 163898 523222 164134
rect 522986 128218 523222 128454
rect 522986 127898 523222 128134
rect 522986 92218 523222 92454
rect 522986 91898 523222 92134
rect 522986 56218 523222 56454
rect 522986 55898 523222 56134
rect 522986 20218 523222 20454
rect 522986 19898 523222 20134
rect 522986 -1522 523222 -1286
rect 522986 -1842 523222 -1606
rect 526586 203818 526822 204054
rect 526586 203498 526822 203734
rect 526586 167818 526822 168054
rect 526586 167498 526822 167734
rect 526586 131818 526822 132054
rect 526586 131498 526822 131734
rect 526586 95818 526822 96054
rect 526586 95498 526822 95734
rect 526586 59818 526822 60054
rect 526586 59498 526822 59734
rect 526586 23818 526822 24054
rect 526586 23498 526822 23734
rect 526586 -3402 526822 -3166
rect 526586 -3722 526822 -3486
rect 530186 207418 530422 207654
rect 530186 207098 530422 207334
rect 530186 171418 530422 171654
rect 530186 171098 530422 171334
rect 530186 135418 530422 135654
rect 530186 135098 530422 135334
rect 530186 99418 530422 99654
rect 530186 99098 530422 99334
rect 530186 63418 530422 63654
rect 530186 63098 530422 63334
rect 530186 27418 530422 27654
rect 530186 27098 530422 27334
rect 530186 -5282 530422 -5046
rect 530186 -5602 530422 -5366
rect 533786 211018 534022 211254
rect 533786 210698 534022 210934
rect 533786 175018 534022 175254
rect 533786 174698 534022 174934
rect 533786 139018 534022 139254
rect 533786 138698 534022 138934
rect 533786 103018 534022 103254
rect 533786 102698 534022 102934
rect 533786 67018 534022 67254
rect 533786 66698 534022 66934
rect 540986 218218 541222 218454
rect 540986 217898 541222 218134
rect 540986 182218 541222 182454
rect 540986 181898 541222 182134
rect 540986 146218 541222 146454
rect 540986 145898 541222 146134
rect 540986 110218 541222 110454
rect 540986 109898 541222 110134
rect 540986 74218 541222 74454
rect 540986 73898 541222 74134
rect 533786 31018 534022 31254
rect 533786 30698 534022 30934
rect 515786 -6222 516022 -5986
rect 515786 -6542 516022 -6306
rect 540986 38218 541222 38454
rect 540986 37898 541222 38134
rect 544586 473818 544822 474054
rect 544586 473498 544822 473734
rect 544586 437818 544822 438054
rect 544586 437498 544822 437734
rect 544586 401818 544822 402054
rect 544586 401498 544822 401734
rect 544586 365818 544822 366054
rect 544586 365498 544822 365734
rect 544586 329818 544822 330054
rect 544586 329498 544822 329734
rect 544586 293818 544822 294054
rect 544586 293498 544822 293734
rect 544586 257818 544822 258054
rect 544586 257498 544822 257734
rect 544586 221818 544822 222054
rect 544586 221498 544822 221734
rect 544586 185818 544822 186054
rect 544586 185498 544822 185734
rect 544586 149818 544822 150054
rect 544586 149498 544822 149734
rect 544586 113818 544822 114054
rect 544586 113498 544822 113734
rect 544586 77818 544822 78054
rect 544586 77498 544822 77734
rect 544586 41818 544822 42054
rect 544586 41498 544822 41734
rect 540986 2218 541222 2454
rect 540986 1898 541222 2134
rect 540986 -582 541222 -346
rect 540986 -902 541222 -666
rect 544586 5818 544822 6054
rect 544586 5498 544822 5734
rect 544586 -2462 544822 -2226
rect 544586 -2782 544822 -2546
rect 548186 693418 548422 693654
rect 548186 693098 548422 693334
rect 548186 657418 548422 657654
rect 548186 657098 548422 657334
rect 548186 621418 548422 621654
rect 548186 621098 548422 621334
rect 548186 585418 548422 585654
rect 548186 585098 548422 585334
rect 548186 549418 548422 549654
rect 548186 549098 548422 549334
rect 548186 513418 548422 513654
rect 548186 513098 548422 513334
rect 548186 477418 548422 477654
rect 548186 477098 548422 477334
rect 548186 441418 548422 441654
rect 548186 441098 548422 441334
rect 548186 405418 548422 405654
rect 548186 405098 548422 405334
rect 548186 369418 548422 369654
rect 548186 369098 548422 369334
rect 548186 333418 548422 333654
rect 548186 333098 548422 333334
rect 548186 297418 548422 297654
rect 548186 297098 548422 297334
rect 548186 261418 548422 261654
rect 548186 261098 548422 261334
rect 548186 225418 548422 225654
rect 548186 225098 548422 225334
rect 548186 189418 548422 189654
rect 548186 189098 548422 189334
rect 548186 153418 548422 153654
rect 548186 153098 548422 153334
rect 548186 117418 548422 117654
rect 548186 117098 548422 117334
rect 548186 81418 548422 81654
rect 548186 81098 548422 81334
rect 548186 45418 548422 45654
rect 548186 45098 548422 45334
rect 548186 9418 548422 9654
rect 548186 9098 548422 9334
rect 548186 -4342 548422 -4106
rect 548186 -4662 548422 -4426
rect 569786 711182 570022 711418
rect 569786 710862 570022 711098
rect 566186 709302 566422 709538
rect 566186 708982 566422 709218
rect 562586 707422 562822 707658
rect 562586 707102 562822 707338
rect 551786 697018 552022 697254
rect 551786 696698 552022 696934
rect 551786 661018 552022 661254
rect 551786 660698 552022 660934
rect 551786 625018 552022 625254
rect 551786 624698 552022 624934
rect 551786 589018 552022 589254
rect 551786 588698 552022 588934
rect 551786 553018 552022 553254
rect 551786 552698 552022 552934
rect 551786 517018 552022 517254
rect 551786 516698 552022 516934
rect 551786 481018 552022 481254
rect 551786 480698 552022 480934
rect 551786 445018 552022 445254
rect 551786 444698 552022 444934
rect 551786 409018 552022 409254
rect 551786 408698 552022 408934
rect 551786 373018 552022 373254
rect 551786 372698 552022 372934
rect 551786 337018 552022 337254
rect 551786 336698 552022 336934
rect 551786 301018 552022 301254
rect 551786 300698 552022 300934
rect 551786 265018 552022 265254
rect 551786 264698 552022 264934
rect 551786 229018 552022 229254
rect 551786 228698 552022 228934
rect 551786 193018 552022 193254
rect 551786 192698 552022 192934
rect 551786 157018 552022 157254
rect 551786 156698 552022 156934
rect 551786 121018 552022 121254
rect 551786 120698 552022 120934
rect 551786 85018 552022 85254
rect 551786 84698 552022 84934
rect 551786 49018 552022 49254
rect 551786 48698 552022 48934
rect 551786 13018 552022 13254
rect 551786 12698 552022 12934
rect 533786 -7162 534022 -6926
rect 533786 -7482 534022 -7246
rect 558986 705542 559222 705778
rect 558986 705222 559222 705458
rect 558986 668218 559222 668454
rect 558986 667898 559222 668134
rect 558986 632218 559222 632454
rect 558986 631898 559222 632134
rect 558986 596218 559222 596454
rect 558986 595898 559222 596134
rect 558986 560218 559222 560454
rect 558986 559898 559222 560134
rect 558986 524218 559222 524454
rect 558986 523898 559222 524134
rect 558986 488218 559222 488454
rect 558986 487898 559222 488134
rect 558986 452218 559222 452454
rect 558986 451898 559222 452134
rect 558986 416218 559222 416454
rect 558986 415898 559222 416134
rect 558986 380218 559222 380454
rect 558986 379898 559222 380134
rect 558986 344218 559222 344454
rect 558986 343898 559222 344134
rect 558986 308218 559222 308454
rect 558986 307898 559222 308134
rect 558986 272218 559222 272454
rect 558986 271898 559222 272134
rect 558986 236218 559222 236454
rect 558986 235898 559222 236134
rect 558986 200218 559222 200454
rect 558986 199898 559222 200134
rect 558986 164218 559222 164454
rect 558986 163898 559222 164134
rect 558986 128218 559222 128454
rect 558986 127898 559222 128134
rect 558986 92218 559222 92454
rect 558986 91898 559222 92134
rect 558986 56218 559222 56454
rect 558986 55898 559222 56134
rect 558986 20218 559222 20454
rect 558986 19898 559222 20134
rect 558986 -1522 559222 -1286
rect 558986 -1842 559222 -1606
rect 562586 671818 562822 672054
rect 562586 671498 562822 671734
rect 562586 635818 562822 636054
rect 562586 635498 562822 635734
rect 562586 599818 562822 600054
rect 562586 599498 562822 599734
rect 562586 563818 562822 564054
rect 562586 563498 562822 563734
rect 562586 527818 562822 528054
rect 562586 527498 562822 527734
rect 562586 491818 562822 492054
rect 562586 491498 562822 491734
rect 562586 455818 562822 456054
rect 562586 455498 562822 455734
rect 562586 419818 562822 420054
rect 562586 419498 562822 419734
rect 562586 383818 562822 384054
rect 562586 383498 562822 383734
rect 562586 347818 562822 348054
rect 562586 347498 562822 347734
rect 562586 311818 562822 312054
rect 562586 311498 562822 311734
rect 562586 275818 562822 276054
rect 562586 275498 562822 275734
rect 562586 239818 562822 240054
rect 562586 239498 562822 239734
rect 562586 203818 562822 204054
rect 562586 203498 562822 203734
rect 562586 167818 562822 168054
rect 562586 167498 562822 167734
rect 562586 131818 562822 132054
rect 562586 131498 562822 131734
rect 562586 95818 562822 96054
rect 562586 95498 562822 95734
rect 562586 59818 562822 60054
rect 562586 59498 562822 59734
rect 562586 23818 562822 24054
rect 562586 23498 562822 23734
rect 562586 -3402 562822 -3166
rect 562586 -3722 562822 -3486
rect 566186 675418 566422 675654
rect 566186 675098 566422 675334
rect 566186 639418 566422 639654
rect 566186 639098 566422 639334
rect 566186 603418 566422 603654
rect 566186 603098 566422 603334
rect 566186 567418 566422 567654
rect 566186 567098 566422 567334
rect 566186 531418 566422 531654
rect 566186 531098 566422 531334
rect 566186 495418 566422 495654
rect 566186 495098 566422 495334
rect 566186 459418 566422 459654
rect 566186 459098 566422 459334
rect 566186 423418 566422 423654
rect 566186 423098 566422 423334
rect 566186 387418 566422 387654
rect 566186 387098 566422 387334
rect 566186 351418 566422 351654
rect 566186 351098 566422 351334
rect 566186 315418 566422 315654
rect 566186 315098 566422 315334
rect 566186 279418 566422 279654
rect 566186 279098 566422 279334
rect 566186 243418 566422 243654
rect 566186 243098 566422 243334
rect 566186 207418 566422 207654
rect 566186 207098 566422 207334
rect 566186 171418 566422 171654
rect 566186 171098 566422 171334
rect 566186 135418 566422 135654
rect 566186 135098 566422 135334
rect 566186 99418 566422 99654
rect 566186 99098 566422 99334
rect 566186 63418 566422 63654
rect 566186 63098 566422 63334
rect 566186 27418 566422 27654
rect 566186 27098 566422 27334
rect 566186 -5282 566422 -5046
rect 566186 -5602 566422 -5366
rect 592082 711182 592318 711418
rect 592082 710862 592318 711098
rect 591142 710242 591378 710478
rect 591142 709922 591378 710158
rect 590202 709302 590438 709538
rect 590202 708982 590438 709218
rect 589262 708362 589498 708598
rect 589262 708042 589498 708278
rect 588322 707422 588558 707658
rect 588322 707102 588558 707338
rect 580586 706482 580822 706718
rect 580586 706162 580822 706398
rect 569786 679018 570022 679254
rect 569786 678698 570022 678934
rect 569786 643018 570022 643254
rect 569786 642698 570022 642934
rect 569786 607018 570022 607254
rect 569786 606698 570022 606934
rect 569786 571018 570022 571254
rect 569786 570698 570022 570934
rect 569786 535018 570022 535254
rect 569786 534698 570022 534934
rect 569786 499018 570022 499254
rect 569786 498698 570022 498934
rect 569786 463018 570022 463254
rect 569786 462698 570022 462934
rect 569786 427018 570022 427254
rect 569786 426698 570022 426934
rect 569786 391018 570022 391254
rect 569786 390698 570022 390934
rect 569786 355018 570022 355254
rect 569786 354698 570022 354934
rect 569786 319018 570022 319254
rect 569786 318698 570022 318934
rect 569786 283018 570022 283254
rect 569786 282698 570022 282934
rect 569786 247018 570022 247254
rect 569786 246698 570022 246934
rect 569786 211018 570022 211254
rect 569786 210698 570022 210934
rect 569786 175018 570022 175254
rect 569786 174698 570022 174934
rect 569786 139018 570022 139254
rect 569786 138698 570022 138934
rect 569786 103018 570022 103254
rect 569786 102698 570022 102934
rect 569786 67018 570022 67254
rect 569786 66698 570022 66934
rect 569786 31018 570022 31254
rect 569786 30698 570022 30934
rect 551786 -6222 552022 -5986
rect 551786 -6542 552022 -6306
rect 576986 704602 577222 704838
rect 576986 704282 577222 704518
rect 576986 686218 577222 686454
rect 576986 685898 577222 686134
rect 576986 650218 577222 650454
rect 576986 649898 577222 650134
rect 576986 614218 577222 614454
rect 576986 613898 577222 614134
rect 576986 578218 577222 578454
rect 576986 577898 577222 578134
rect 576986 542218 577222 542454
rect 576986 541898 577222 542134
rect 576986 506218 577222 506454
rect 576986 505898 577222 506134
rect 576986 470218 577222 470454
rect 576986 469898 577222 470134
rect 576986 434218 577222 434454
rect 576986 433898 577222 434134
rect 576986 398218 577222 398454
rect 576986 397898 577222 398134
rect 576986 362218 577222 362454
rect 576986 361898 577222 362134
rect 576986 326218 577222 326454
rect 576986 325898 577222 326134
rect 576986 290218 577222 290454
rect 576986 289898 577222 290134
rect 576986 254218 577222 254454
rect 576986 253898 577222 254134
rect 576986 218218 577222 218454
rect 576986 217898 577222 218134
rect 576986 182218 577222 182454
rect 576986 181898 577222 182134
rect 576986 146218 577222 146454
rect 576986 145898 577222 146134
rect 576986 110218 577222 110454
rect 576986 109898 577222 110134
rect 576986 74218 577222 74454
rect 576986 73898 577222 74134
rect 576986 38218 577222 38454
rect 576986 37898 577222 38134
rect 576986 2218 577222 2454
rect 576986 1898 577222 2134
rect 576986 -582 577222 -346
rect 576986 -902 577222 -666
rect 587382 706482 587618 706718
rect 587382 706162 587618 706398
rect 586442 705542 586678 705778
rect 586442 705222 586678 705458
rect 580586 689818 580822 690054
rect 580586 689498 580822 689734
rect 580586 653818 580822 654054
rect 580586 653498 580822 653734
rect 580586 617818 580822 618054
rect 580586 617498 580822 617734
rect 580586 581818 580822 582054
rect 580586 581498 580822 581734
rect 580586 545818 580822 546054
rect 580586 545498 580822 545734
rect 580586 509818 580822 510054
rect 580586 509498 580822 509734
rect 580586 473818 580822 474054
rect 580586 473498 580822 473734
rect 580586 437818 580822 438054
rect 580586 437498 580822 437734
rect 580586 401818 580822 402054
rect 580586 401498 580822 401734
rect 580586 365818 580822 366054
rect 580586 365498 580822 365734
rect 580586 329818 580822 330054
rect 580586 329498 580822 329734
rect 580586 293818 580822 294054
rect 580586 293498 580822 293734
rect 580586 257818 580822 258054
rect 580586 257498 580822 257734
rect 580586 221818 580822 222054
rect 580586 221498 580822 221734
rect 580586 185818 580822 186054
rect 580586 185498 580822 185734
rect 580586 149818 580822 150054
rect 580586 149498 580822 149734
rect 580586 113818 580822 114054
rect 580586 113498 580822 113734
rect 580586 77818 580822 78054
rect 580586 77498 580822 77734
rect 580586 41818 580822 42054
rect 580586 41498 580822 41734
rect 580586 5818 580822 6054
rect 580586 5498 580822 5734
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 686218 585738 686454
rect 585502 685898 585738 686134
rect 585502 650218 585738 650454
rect 585502 649898 585738 650134
rect 585502 614218 585738 614454
rect 585502 613898 585738 614134
rect 585502 578218 585738 578454
rect 585502 577898 585738 578134
rect 585502 542218 585738 542454
rect 585502 541898 585738 542134
rect 585502 506218 585738 506454
rect 585502 505898 585738 506134
rect 585502 470218 585738 470454
rect 585502 469898 585738 470134
rect 585502 434218 585738 434454
rect 585502 433898 585738 434134
rect 585502 398218 585738 398454
rect 585502 397898 585738 398134
rect 585502 362218 585738 362454
rect 585502 361898 585738 362134
rect 585502 326218 585738 326454
rect 585502 325898 585738 326134
rect 585502 290218 585738 290454
rect 585502 289898 585738 290134
rect 585502 254218 585738 254454
rect 585502 253898 585738 254134
rect 585502 218218 585738 218454
rect 585502 217898 585738 218134
rect 585502 182218 585738 182454
rect 585502 181898 585738 182134
rect 585502 146218 585738 146454
rect 585502 145898 585738 146134
rect 585502 110218 585738 110454
rect 585502 109898 585738 110134
rect 585502 74218 585738 74454
rect 585502 73898 585738 74134
rect 585502 38218 585738 38454
rect 585502 37898 585738 38134
rect 585502 2218 585738 2454
rect 585502 1898 585738 2134
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586442 668218 586678 668454
rect 586442 667898 586678 668134
rect 586442 632218 586678 632454
rect 586442 631898 586678 632134
rect 586442 596218 586678 596454
rect 586442 595898 586678 596134
rect 586442 560218 586678 560454
rect 586442 559898 586678 560134
rect 586442 524218 586678 524454
rect 586442 523898 586678 524134
rect 586442 488218 586678 488454
rect 586442 487898 586678 488134
rect 586442 452218 586678 452454
rect 586442 451898 586678 452134
rect 586442 416218 586678 416454
rect 586442 415898 586678 416134
rect 586442 380218 586678 380454
rect 586442 379898 586678 380134
rect 586442 344218 586678 344454
rect 586442 343898 586678 344134
rect 586442 308218 586678 308454
rect 586442 307898 586678 308134
rect 586442 272218 586678 272454
rect 586442 271898 586678 272134
rect 586442 236218 586678 236454
rect 586442 235898 586678 236134
rect 586442 200218 586678 200454
rect 586442 199898 586678 200134
rect 586442 164218 586678 164454
rect 586442 163898 586678 164134
rect 586442 128218 586678 128454
rect 586442 127898 586678 128134
rect 586442 92218 586678 92454
rect 586442 91898 586678 92134
rect 586442 56218 586678 56454
rect 586442 55898 586678 56134
rect 586442 20218 586678 20454
rect 586442 19898 586678 20134
rect 586442 -1522 586678 -1286
rect 586442 -1842 586678 -1606
rect 587382 689818 587618 690054
rect 587382 689498 587618 689734
rect 587382 653818 587618 654054
rect 587382 653498 587618 653734
rect 587382 617818 587618 618054
rect 587382 617498 587618 617734
rect 587382 581818 587618 582054
rect 587382 581498 587618 581734
rect 587382 545818 587618 546054
rect 587382 545498 587618 545734
rect 587382 509818 587618 510054
rect 587382 509498 587618 509734
rect 587382 473818 587618 474054
rect 587382 473498 587618 473734
rect 587382 437818 587618 438054
rect 587382 437498 587618 437734
rect 587382 401818 587618 402054
rect 587382 401498 587618 401734
rect 587382 365818 587618 366054
rect 587382 365498 587618 365734
rect 587382 329818 587618 330054
rect 587382 329498 587618 329734
rect 587382 293818 587618 294054
rect 587382 293498 587618 293734
rect 587382 257818 587618 258054
rect 587382 257498 587618 257734
rect 587382 221818 587618 222054
rect 587382 221498 587618 221734
rect 587382 185818 587618 186054
rect 587382 185498 587618 185734
rect 587382 149818 587618 150054
rect 587382 149498 587618 149734
rect 587382 113818 587618 114054
rect 587382 113498 587618 113734
rect 587382 77818 587618 78054
rect 587382 77498 587618 77734
rect 587382 41818 587618 42054
rect 587382 41498 587618 41734
rect 587382 5818 587618 6054
rect 587382 5498 587618 5734
rect 580586 -2462 580822 -2226
rect 580586 -2782 580822 -2546
rect 587382 -2462 587618 -2226
rect 587382 -2782 587618 -2546
rect 588322 671818 588558 672054
rect 588322 671498 588558 671734
rect 588322 635818 588558 636054
rect 588322 635498 588558 635734
rect 588322 599818 588558 600054
rect 588322 599498 588558 599734
rect 588322 563818 588558 564054
rect 588322 563498 588558 563734
rect 588322 527818 588558 528054
rect 588322 527498 588558 527734
rect 588322 491818 588558 492054
rect 588322 491498 588558 491734
rect 588322 455818 588558 456054
rect 588322 455498 588558 455734
rect 588322 419818 588558 420054
rect 588322 419498 588558 419734
rect 588322 383818 588558 384054
rect 588322 383498 588558 383734
rect 588322 347818 588558 348054
rect 588322 347498 588558 347734
rect 588322 311818 588558 312054
rect 588322 311498 588558 311734
rect 588322 275818 588558 276054
rect 588322 275498 588558 275734
rect 588322 239818 588558 240054
rect 588322 239498 588558 239734
rect 588322 203818 588558 204054
rect 588322 203498 588558 203734
rect 588322 167818 588558 168054
rect 588322 167498 588558 167734
rect 588322 131818 588558 132054
rect 588322 131498 588558 131734
rect 588322 95818 588558 96054
rect 588322 95498 588558 95734
rect 588322 59818 588558 60054
rect 588322 59498 588558 59734
rect 588322 23818 588558 24054
rect 588322 23498 588558 23734
rect 588322 -3402 588558 -3166
rect 588322 -3722 588558 -3486
rect 589262 693418 589498 693654
rect 589262 693098 589498 693334
rect 589262 657418 589498 657654
rect 589262 657098 589498 657334
rect 589262 621418 589498 621654
rect 589262 621098 589498 621334
rect 589262 585418 589498 585654
rect 589262 585098 589498 585334
rect 589262 549418 589498 549654
rect 589262 549098 589498 549334
rect 589262 513418 589498 513654
rect 589262 513098 589498 513334
rect 589262 477418 589498 477654
rect 589262 477098 589498 477334
rect 589262 441418 589498 441654
rect 589262 441098 589498 441334
rect 589262 405418 589498 405654
rect 589262 405098 589498 405334
rect 589262 369418 589498 369654
rect 589262 369098 589498 369334
rect 589262 333418 589498 333654
rect 589262 333098 589498 333334
rect 589262 297418 589498 297654
rect 589262 297098 589498 297334
rect 589262 261418 589498 261654
rect 589262 261098 589498 261334
rect 589262 225418 589498 225654
rect 589262 225098 589498 225334
rect 589262 189418 589498 189654
rect 589262 189098 589498 189334
rect 589262 153418 589498 153654
rect 589262 153098 589498 153334
rect 589262 117418 589498 117654
rect 589262 117098 589498 117334
rect 589262 81418 589498 81654
rect 589262 81098 589498 81334
rect 589262 45418 589498 45654
rect 589262 45098 589498 45334
rect 589262 9418 589498 9654
rect 589262 9098 589498 9334
rect 589262 -4342 589498 -4106
rect 589262 -4662 589498 -4426
rect 590202 675418 590438 675654
rect 590202 675098 590438 675334
rect 590202 639418 590438 639654
rect 590202 639098 590438 639334
rect 590202 603418 590438 603654
rect 590202 603098 590438 603334
rect 590202 567418 590438 567654
rect 590202 567098 590438 567334
rect 590202 531418 590438 531654
rect 590202 531098 590438 531334
rect 590202 495418 590438 495654
rect 590202 495098 590438 495334
rect 590202 459418 590438 459654
rect 590202 459098 590438 459334
rect 590202 423418 590438 423654
rect 590202 423098 590438 423334
rect 590202 387418 590438 387654
rect 590202 387098 590438 387334
rect 590202 351418 590438 351654
rect 590202 351098 590438 351334
rect 590202 315418 590438 315654
rect 590202 315098 590438 315334
rect 590202 279418 590438 279654
rect 590202 279098 590438 279334
rect 590202 243418 590438 243654
rect 590202 243098 590438 243334
rect 590202 207418 590438 207654
rect 590202 207098 590438 207334
rect 590202 171418 590438 171654
rect 590202 171098 590438 171334
rect 590202 135418 590438 135654
rect 590202 135098 590438 135334
rect 590202 99418 590438 99654
rect 590202 99098 590438 99334
rect 590202 63418 590438 63654
rect 590202 63098 590438 63334
rect 590202 27418 590438 27654
rect 590202 27098 590438 27334
rect 590202 -5282 590438 -5046
rect 590202 -5602 590438 -5366
rect 591142 697018 591378 697254
rect 591142 696698 591378 696934
rect 591142 661018 591378 661254
rect 591142 660698 591378 660934
rect 591142 625018 591378 625254
rect 591142 624698 591378 624934
rect 591142 589018 591378 589254
rect 591142 588698 591378 588934
rect 591142 553018 591378 553254
rect 591142 552698 591378 552934
rect 591142 517018 591378 517254
rect 591142 516698 591378 516934
rect 591142 481018 591378 481254
rect 591142 480698 591378 480934
rect 591142 445018 591378 445254
rect 591142 444698 591378 444934
rect 591142 409018 591378 409254
rect 591142 408698 591378 408934
rect 591142 373018 591378 373254
rect 591142 372698 591378 372934
rect 591142 337018 591378 337254
rect 591142 336698 591378 336934
rect 591142 301018 591378 301254
rect 591142 300698 591378 300934
rect 591142 265018 591378 265254
rect 591142 264698 591378 264934
rect 591142 229018 591378 229254
rect 591142 228698 591378 228934
rect 591142 193018 591378 193254
rect 591142 192698 591378 192934
rect 591142 157018 591378 157254
rect 591142 156698 591378 156934
rect 591142 121018 591378 121254
rect 591142 120698 591378 120934
rect 591142 85018 591378 85254
rect 591142 84698 591378 84934
rect 591142 49018 591378 49254
rect 591142 48698 591378 48934
rect 591142 13018 591378 13254
rect 591142 12698 591378 12934
rect 591142 -6222 591378 -5986
rect 591142 -6542 591378 -6306
rect 592082 679018 592318 679254
rect 592082 678698 592318 678934
rect 592082 643018 592318 643254
rect 592082 642698 592318 642934
rect 592082 607018 592318 607254
rect 592082 606698 592318 606934
rect 592082 571018 592318 571254
rect 592082 570698 592318 570934
rect 592082 535018 592318 535254
rect 592082 534698 592318 534934
rect 592082 499018 592318 499254
rect 592082 498698 592318 498934
rect 592082 463018 592318 463254
rect 592082 462698 592318 462934
rect 592082 427018 592318 427254
rect 592082 426698 592318 426934
rect 592082 391018 592318 391254
rect 592082 390698 592318 390934
rect 592082 355018 592318 355254
rect 592082 354698 592318 354934
rect 592082 319018 592318 319254
rect 592082 318698 592318 318934
rect 592082 283018 592318 283254
rect 592082 282698 592318 282934
rect 592082 247018 592318 247254
rect 592082 246698 592318 246934
rect 592082 211018 592318 211254
rect 592082 210698 592318 210934
rect 592082 175018 592318 175254
rect 592082 174698 592318 174934
rect 592082 139018 592318 139254
rect 592082 138698 592318 138934
rect 592082 103018 592318 103254
rect 592082 102698 592318 102934
rect 592082 67018 592318 67254
rect 592082 66698 592318 66934
rect 592082 31018 592318 31254
rect 592082 30698 592318 30934
rect 569786 -7162 570022 -6926
rect 569786 -7482 570022 -7246
rect 592082 -7162 592318 -6926
rect 592082 -7482 592318 -7246
<< metal5 >>
rect -8576 711440 -7976 711442
rect 29604 711440 30204 711442
rect 65604 711440 66204 711442
rect 101604 711440 102204 711442
rect 137604 711440 138204 711442
rect 173604 711440 174204 711442
rect 209604 711440 210204 711442
rect 245604 711440 246204 711442
rect 281604 711440 282204 711442
rect 317604 711440 318204 711442
rect 353604 711440 354204 711442
rect 389604 711440 390204 711442
rect 425604 711440 426204 711442
rect 461604 711440 462204 711442
rect 497604 711440 498204 711442
rect 533604 711440 534204 711442
rect 569604 711440 570204 711442
rect 591900 711440 592500 711442
rect -8576 711418 592500 711440
rect -8576 711182 -8394 711418
rect -8158 711182 29786 711418
rect 30022 711182 65786 711418
rect 66022 711182 101786 711418
rect 102022 711182 137786 711418
rect 138022 711182 173786 711418
rect 174022 711182 209786 711418
rect 210022 711182 245786 711418
rect 246022 711182 281786 711418
rect 282022 711182 317786 711418
rect 318022 711182 353786 711418
rect 354022 711182 389786 711418
rect 390022 711182 425786 711418
rect 426022 711182 461786 711418
rect 462022 711182 497786 711418
rect 498022 711182 533786 711418
rect 534022 711182 569786 711418
rect 570022 711182 592082 711418
rect 592318 711182 592500 711418
rect -8576 711098 592500 711182
rect -8576 710862 -8394 711098
rect -8158 710862 29786 711098
rect 30022 710862 65786 711098
rect 66022 710862 101786 711098
rect 102022 710862 137786 711098
rect 138022 710862 173786 711098
rect 174022 710862 209786 711098
rect 210022 710862 245786 711098
rect 246022 710862 281786 711098
rect 282022 710862 317786 711098
rect 318022 710862 353786 711098
rect 354022 710862 389786 711098
rect 390022 710862 425786 711098
rect 426022 710862 461786 711098
rect 462022 710862 497786 711098
rect 498022 710862 533786 711098
rect 534022 710862 569786 711098
rect 570022 710862 592082 711098
rect 592318 710862 592500 711098
rect -8576 710840 592500 710862
rect -8576 710838 -7976 710840
rect 29604 710838 30204 710840
rect 65604 710838 66204 710840
rect 101604 710838 102204 710840
rect 137604 710838 138204 710840
rect 173604 710838 174204 710840
rect 209604 710838 210204 710840
rect 245604 710838 246204 710840
rect 281604 710838 282204 710840
rect 317604 710838 318204 710840
rect 353604 710838 354204 710840
rect 389604 710838 390204 710840
rect 425604 710838 426204 710840
rect 461604 710838 462204 710840
rect 497604 710838 498204 710840
rect 533604 710838 534204 710840
rect 569604 710838 570204 710840
rect 591900 710838 592500 710840
rect -7636 710500 -7036 710502
rect 11604 710500 12204 710502
rect 47604 710500 48204 710502
rect 83604 710500 84204 710502
rect 119604 710500 120204 710502
rect 155604 710500 156204 710502
rect 191604 710500 192204 710502
rect 227604 710500 228204 710502
rect 263604 710500 264204 710502
rect 299604 710500 300204 710502
rect 335604 710500 336204 710502
rect 371604 710500 372204 710502
rect 407604 710500 408204 710502
rect 443604 710500 444204 710502
rect 479604 710500 480204 710502
rect 515604 710500 516204 710502
rect 551604 710500 552204 710502
rect 590960 710500 591560 710502
rect -7636 710478 591560 710500
rect -7636 710242 -7454 710478
rect -7218 710242 11786 710478
rect 12022 710242 47786 710478
rect 48022 710242 83786 710478
rect 84022 710242 119786 710478
rect 120022 710242 155786 710478
rect 156022 710242 191786 710478
rect 192022 710242 227786 710478
rect 228022 710242 263786 710478
rect 264022 710242 299786 710478
rect 300022 710242 335786 710478
rect 336022 710242 371786 710478
rect 372022 710242 407786 710478
rect 408022 710242 443786 710478
rect 444022 710242 479786 710478
rect 480022 710242 515786 710478
rect 516022 710242 551786 710478
rect 552022 710242 591142 710478
rect 591378 710242 591560 710478
rect -7636 710158 591560 710242
rect -7636 709922 -7454 710158
rect -7218 709922 11786 710158
rect 12022 709922 47786 710158
rect 48022 709922 83786 710158
rect 84022 709922 119786 710158
rect 120022 709922 155786 710158
rect 156022 709922 191786 710158
rect 192022 709922 227786 710158
rect 228022 709922 263786 710158
rect 264022 709922 299786 710158
rect 300022 709922 335786 710158
rect 336022 709922 371786 710158
rect 372022 709922 407786 710158
rect 408022 709922 443786 710158
rect 444022 709922 479786 710158
rect 480022 709922 515786 710158
rect 516022 709922 551786 710158
rect 552022 709922 591142 710158
rect 591378 709922 591560 710158
rect -7636 709900 591560 709922
rect -7636 709898 -7036 709900
rect 11604 709898 12204 709900
rect 47604 709898 48204 709900
rect 83604 709898 84204 709900
rect 119604 709898 120204 709900
rect 155604 709898 156204 709900
rect 191604 709898 192204 709900
rect 227604 709898 228204 709900
rect 263604 709898 264204 709900
rect 299604 709898 300204 709900
rect 335604 709898 336204 709900
rect 371604 709898 372204 709900
rect 407604 709898 408204 709900
rect 443604 709898 444204 709900
rect 479604 709898 480204 709900
rect 515604 709898 516204 709900
rect 551604 709898 552204 709900
rect 590960 709898 591560 709900
rect -6696 709560 -6096 709562
rect 26004 709560 26604 709562
rect 62004 709560 62604 709562
rect 98004 709560 98604 709562
rect 134004 709560 134604 709562
rect 170004 709560 170604 709562
rect 206004 709560 206604 709562
rect 242004 709560 242604 709562
rect 278004 709560 278604 709562
rect 314004 709560 314604 709562
rect 350004 709560 350604 709562
rect 386004 709560 386604 709562
rect 422004 709560 422604 709562
rect 458004 709560 458604 709562
rect 494004 709560 494604 709562
rect 530004 709560 530604 709562
rect 566004 709560 566604 709562
rect 590020 709560 590620 709562
rect -6696 709538 590620 709560
rect -6696 709302 -6514 709538
rect -6278 709302 26186 709538
rect 26422 709302 62186 709538
rect 62422 709302 98186 709538
rect 98422 709302 134186 709538
rect 134422 709302 170186 709538
rect 170422 709302 206186 709538
rect 206422 709302 242186 709538
rect 242422 709302 278186 709538
rect 278422 709302 314186 709538
rect 314422 709302 350186 709538
rect 350422 709302 386186 709538
rect 386422 709302 422186 709538
rect 422422 709302 458186 709538
rect 458422 709302 494186 709538
rect 494422 709302 530186 709538
rect 530422 709302 566186 709538
rect 566422 709302 590202 709538
rect 590438 709302 590620 709538
rect -6696 709218 590620 709302
rect -6696 708982 -6514 709218
rect -6278 708982 26186 709218
rect 26422 708982 62186 709218
rect 62422 708982 98186 709218
rect 98422 708982 134186 709218
rect 134422 708982 170186 709218
rect 170422 708982 206186 709218
rect 206422 708982 242186 709218
rect 242422 708982 278186 709218
rect 278422 708982 314186 709218
rect 314422 708982 350186 709218
rect 350422 708982 386186 709218
rect 386422 708982 422186 709218
rect 422422 708982 458186 709218
rect 458422 708982 494186 709218
rect 494422 708982 530186 709218
rect 530422 708982 566186 709218
rect 566422 708982 590202 709218
rect 590438 708982 590620 709218
rect -6696 708960 590620 708982
rect -6696 708958 -6096 708960
rect 26004 708958 26604 708960
rect 62004 708958 62604 708960
rect 98004 708958 98604 708960
rect 134004 708958 134604 708960
rect 170004 708958 170604 708960
rect 206004 708958 206604 708960
rect 242004 708958 242604 708960
rect 278004 708958 278604 708960
rect 314004 708958 314604 708960
rect 350004 708958 350604 708960
rect 386004 708958 386604 708960
rect 422004 708958 422604 708960
rect 458004 708958 458604 708960
rect 494004 708958 494604 708960
rect 530004 708958 530604 708960
rect 566004 708958 566604 708960
rect 590020 708958 590620 708960
rect -5756 708620 -5156 708622
rect 8004 708620 8604 708622
rect 44004 708620 44604 708622
rect 80004 708620 80604 708622
rect 116004 708620 116604 708622
rect 152004 708620 152604 708622
rect 188004 708620 188604 708622
rect 224004 708620 224604 708622
rect 260004 708620 260604 708622
rect 296004 708620 296604 708622
rect 332004 708620 332604 708622
rect 368004 708620 368604 708622
rect 404004 708620 404604 708622
rect 440004 708620 440604 708622
rect 476004 708620 476604 708622
rect 512004 708620 512604 708622
rect 548004 708620 548604 708622
rect 589080 708620 589680 708622
rect -5756 708598 589680 708620
rect -5756 708362 -5574 708598
rect -5338 708362 8186 708598
rect 8422 708362 44186 708598
rect 44422 708362 80186 708598
rect 80422 708362 116186 708598
rect 116422 708362 152186 708598
rect 152422 708362 188186 708598
rect 188422 708362 224186 708598
rect 224422 708362 260186 708598
rect 260422 708362 296186 708598
rect 296422 708362 332186 708598
rect 332422 708362 368186 708598
rect 368422 708362 404186 708598
rect 404422 708362 440186 708598
rect 440422 708362 476186 708598
rect 476422 708362 512186 708598
rect 512422 708362 548186 708598
rect 548422 708362 589262 708598
rect 589498 708362 589680 708598
rect -5756 708278 589680 708362
rect -5756 708042 -5574 708278
rect -5338 708042 8186 708278
rect 8422 708042 44186 708278
rect 44422 708042 80186 708278
rect 80422 708042 116186 708278
rect 116422 708042 152186 708278
rect 152422 708042 188186 708278
rect 188422 708042 224186 708278
rect 224422 708042 260186 708278
rect 260422 708042 296186 708278
rect 296422 708042 332186 708278
rect 332422 708042 368186 708278
rect 368422 708042 404186 708278
rect 404422 708042 440186 708278
rect 440422 708042 476186 708278
rect 476422 708042 512186 708278
rect 512422 708042 548186 708278
rect 548422 708042 589262 708278
rect 589498 708042 589680 708278
rect -5756 708020 589680 708042
rect -5756 708018 -5156 708020
rect 8004 708018 8604 708020
rect 44004 708018 44604 708020
rect 80004 708018 80604 708020
rect 116004 708018 116604 708020
rect 152004 708018 152604 708020
rect 188004 708018 188604 708020
rect 224004 708018 224604 708020
rect 260004 708018 260604 708020
rect 296004 708018 296604 708020
rect 332004 708018 332604 708020
rect 368004 708018 368604 708020
rect 404004 708018 404604 708020
rect 440004 708018 440604 708020
rect 476004 708018 476604 708020
rect 512004 708018 512604 708020
rect 548004 708018 548604 708020
rect 589080 708018 589680 708020
rect -4816 707680 -4216 707682
rect 22404 707680 23004 707682
rect 58404 707680 59004 707682
rect 94404 707680 95004 707682
rect 130404 707680 131004 707682
rect 166404 707680 167004 707682
rect 202404 707680 203004 707682
rect 238404 707680 239004 707682
rect 274404 707680 275004 707682
rect 310404 707680 311004 707682
rect 346404 707680 347004 707682
rect 382404 707680 383004 707682
rect 418404 707680 419004 707682
rect 454404 707680 455004 707682
rect 490404 707680 491004 707682
rect 526404 707680 527004 707682
rect 562404 707680 563004 707682
rect 588140 707680 588740 707682
rect -4816 707658 588740 707680
rect -4816 707422 -4634 707658
rect -4398 707422 22586 707658
rect 22822 707422 58586 707658
rect 58822 707422 94586 707658
rect 94822 707422 130586 707658
rect 130822 707422 166586 707658
rect 166822 707422 202586 707658
rect 202822 707422 238586 707658
rect 238822 707422 274586 707658
rect 274822 707422 310586 707658
rect 310822 707422 346586 707658
rect 346822 707422 382586 707658
rect 382822 707422 418586 707658
rect 418822 707422 454586 707658
rect 454822 707422 490586 707658
rect 490822 707422 526586 707658
rect 526822 707422 562586 707658
rect 562822 707422 588322 707658
rect 588558 707422 588740 707658
rect -4816 707338 588740 707422
rect -4816 707102 -4634 707338
rect -4398 707102 22586 707338
rect 22822 707102 58586 707338
rect 58822 707102 94586 707338
rect 94822 707102 130586 707338
rect 130822 707102 166586 707338
rect 166822 707102 202586 707338
rect 202822 707102 238586 707338
rect 238822 707102 274586 707338
rect 274822 707102 310586 707338
rect 310822 707102 346586 707338
rect 346822 707102 382586 707338
rect 382822 707102 418586 707338
rect 418822 707102 454586 707338
rect 454822 707102 490586 707338
rect 490822 707102 526586 707338
rect 526822 707102 562586 707338
rect 562822 707102 588322 707338
rect 588558 707102 588740 707338
rect -4816 707080 588740 707102
rect -4816 707078 -4216 707080
rect 22404 707078 23004 707080
rect 58404 707078 59004 707080
rect 94404 707078 95004 707080
rect 130404 707078 131004 707080
rect 166404 707078 167004 707080
rect 202404 707078 203004 707080
rect 238404 707078 239004 707080
rect 274404 707078 275004 707080
rect 310404 707078 311004 707080
rect 346404 707078 347004 707080
rect 382404 707078 383004 707080
rect 418404 707078 419004 707080
rect 454404 707078 455004 707080
rect 490404 707078 491004 707080
rect 526404 707078 527004 707080
rect 562404 707078 563004 707080
rect 588140 707078 588740 707080
rect -3876 706740 -3276 706742
rect 4404 706740 5004 706742
rect 40404 706740 41004 706742
rect 76404 706740 77004 706742
rect 112404 706740 113004 706742
rect 148404 706740 149004 706742
rect 184404 706740 185004 706742
rect 220404 706740 221004 706742
rect 256404 706740 257004 706742
rect 292404 706740 293004 706742
rect 328404 706740 329004 706742
rect 364404 706740 365004 706742
rect 400404 706740 401004 706742
rect 436404 706740 437004 706742
rect 472404 706740 473004 706742
rect 508404 706740 509004 706742
rect 544404 706740 545004 706742
rect 580404 706740 581004 706742
rect 587200 706740 587800 706742
rect -3876 706718 587800 706740
rect -3876 706482 -3694 706718
rect -3458 706482 4586 706718
rect 4822 706482 40586 706718
rect 40822 706482 76586 706718
rect 76822 706482 112586 706718
rect 112822 706482 148586 706718
rect 148822 706482 184586 706718
rect 184822 706482 220586 706718
rect 220822 706482 256586 706718
rect 256822 706482 292586 706718
rect 292822 706482 328586 706718
rect 328822 706482 364586 706718
rect 364822 706482 400586 706718
rect 400822 706482 436586 706718
rect 436822 706482 472586 706718
rect 472822 706482 508586 706718
rect 508822 706482 544586 706718
rect 544822 706482 580586 706718
rect 580822 706482 587382 706718
rect 587618 706482 587800 706718
rect -3876 706398 587800 706482
rect -3876 706162 -3694 706398
rect -3458 706162 4586 706398
rect 4822 706162 40586 706398
rect 40822 706162 76586 706398
rect 76822 706162 112586 706398
rect 112822 706162 148586 706398
rect 148822 706162 184586 706398
rect 184822 706162 220586 706398
rect 220822 706162 256586 706398
rect 256822 706162 292586 706398
rect 292822 706162 328586 706398
rect 328822 706162 364586 706398
rect 364822 706162 400586 706398
rect 400822 706162 436586 706398
rect 436822 706162 472586 706398
rect 472822 706162 508586 706398
rect 508822 706162 544586 706398
rect 544822 706162 580586 706398
rect 580822 706162 587382 706398
rect 587618 706162 587800 706398
rect -3876 706140 587800 706162
rect -3876 706138 -3276 706140
rect 4404 706138 5004 706140
rect 40404 706138 41004 706140
rect 76404 706138 77004 706140
rect 112404 706138 113004 706140
rect 148404 706138 149004 706140
rect 184404 706138 185004 706140
rect 220404 706138 221004 706140
rect 256404 706138 257004 706140
rect 292404 706138 293004 706140
rect 328404 706138 329004 706140
rect 364404 706138 365004 706140
rect 400404 706138 401004 706140
rect 436404 706138 437004 706140
rect 472404 706138 473004 706140
rect 508404 706138 509004 706140
rect 544404 706138 545004 706140
rect 580404 706138 581004 706140
rect 587200 706138 587800 706140
rect -2936 705800 -2336 705802
rect 18804 705800 19404 705802
rect 54804 705800 55404 705802
rect 90804 705800 91404 705802
rect 126804 705800 127404 705802
rect 162804 705800 163404 705802
rect 198804 705800 199404 705802
rect 234804 705800 235404 705802
rect 270804 705800 271404 705802
rect 306804 705800 307404 705802
rect 342804 705800 343404 705802
rect 378804 705800 379404 705802
rect 414804 705800 415404 705802
rect 450804 705800 451404 705802
rect 486804 705800 487404 705802
rect 522804 705800 523404 705802
rect 558804 705800 559404 705802
rect 586260 705800 586860 705802
rect -2936 705778 586860 705800
rect -2936 705542 -2754 705778
rect -2518 705542 18986 705778
rect 19222 705542 54986 705778
rect 55222 705542 90986 705778
rect 91222 705542 126986 705778
rect 127222 705542 162986 705778
rect 163222 705542 198986 705778
rect 199222 705542 234986 705778
rect 235222 705542 270986 705778
rect 271222 705542 306986 705778
rect 307222 705542 342986 705778
rect 343222 705542 378986 705778
rect 379222 705542 414986 705778
rect 415222 705542 450986 705778
rect 451222 705542 486986 705778
rect 487222 705542 522986 705778
rect 523222 705542 558986 705778
rect 559222 705542 586442 705778
rect 586678 705542 586860 705778
rect -2936 705458 586860 705542
rect -2936 705222 -2754 705458
rect -2518 705222 18986 705458
rect 19222 705222 54986 705458
rect 55222 705222 90986 705458
rect 91222 705222 126986 705458
rect 127222 705222 162986 705458
rect 163222 705222 198986 705458
rect 199222 705222 234986 705458
rect 235222 705222 270986 705458
rect 271222 705222 306986 705458
rect 307222 705222 342986 705458
rect 343222 705222 378986 705458
rect 379222 705222 414986 705458
rect 415222 705222 450986 705458
rect 451222 705222 486986 705458
rect 487222 705222 522986 705458
rect 523222 705222 558986 705458
rect 559222 705222 586442 705458
rect 586678 705222 586860 705458
rect -2936 705200 586860 705222
rect -2936 705198 -2336 705200
rect 18804 705198 19404 705200
rect 54804 705198 55404 705200
rect 90804 705198 91404 705200
rect 126804 705198 127404 705200
rect 162804 705198 163404 705200
rect 198804 705198 199404 705200
rect 234804 705198 235404 705200
rect 270804 705198 271404 705200
rect 306804 705198 307404 705200
rect 342804 705198 343404 705200
rect 378804 705198 379404 705200
rect 414804 705198 415404 705200
rect 450804 705198 451404 705200
rect 486804 705198 487404 705200
rect 522804 705198 523404 705200
rect 558804 705198 559404 705200
rect 586260 705198 586860 705200
rect -1996 704860 -1396 704862
rect 804 704860 1404 704862
rect 36804 704860 37404 704862
rect 72804 704860 73404 704862
rect 108804 704860 109404 704862
rect 144804 704860 145404 704862
rect 180804 704860 181404 704862
rect 216804 704860 217404 704862
rect 252804 704860 253404 704862
rect 288804 704860 289404 704862
rect 324804 704860 325404 704862
rect 360804 704860 361404 704862
rect 396804 704860 397404 704862
rect 432804 704860 433404 704862
rect 468804 704860 469404 704862
rect 504804 704860 505404 704862
rect 540804 704860 541404 704862
rect 576804 704860 577404 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 986 704838
rect 1222 704602 36986 704838
rect 37222 704602 72986 704838
rect 73222 704602 108986 704838
rect 109222 704602 144986 704838
rect 145222 704602 180986 704838
rect 181222 704602 216986 704838
rect 217222 704602 252986 704838
rect 253222 704602 288986 704838
rect 289222 704602 324986 704838
rect 325222 704602 360986 704838
rect 361222 704602 396986 704838
rect 397222 704602 432986 704838
rect 433222 704602 468986 704838
rect 469222 704602 504986 704838
rect 505222 704602 540986 704838
rect 541222 704602 576986 704838
rect 577222 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 986 704518
rect 1222 704282 36986 704518
rect 37222 704282 72986 704518
rect 73222 704282 108986 704518
rect 109222 704282 144986 704518
rect 145222 704282 180986 704518
rect 181222 704282 216986 704518
rect 217222 704282 252986 704518
rect 253222 704282 288986 704518
rect 289222 704282 324986 704518
rect 325222 704282 360986 704518
rect 361222 704282 396986 704518
rect 397222 704282 432986 704518
rect 433222 704282 468986 704518
rect 469222 704282 504986 704518
rect 505222 704282 540986 704518
rect 541222 704282 576986 704518
rect 577222 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 804 704258 1404 704260
rect 36804 704258 37404 704260
rect 72804 704258 73404 704260
rect 108804 704258 109404 704260
rect 144804 704258 145404 704260
rect 180804 704258 181404 704260
rect 216804 704258 217404 704260
rect 252804 704258 253404 704260
rect 288804 704258 289404 704260
rect 324804 704258 325404 704260
rect 360804 704258 361404 704260
rect 396804 704258 397404 704260
rect 432804 704258 433404 704260
rect 468804 704258 469404 704260
rect 504804 704258 505404 704260
rect 540804 704258 541404 704260
rect 576804 704258 577404 704260
rect 585320 704258 585920 704260
rect -7636 697276 -7036 697278
rect 11604 697276 12204 697278
rect 47604 697276 48204 697278
rect 83604 697276 84204 697278
rect 119604 697276 120204 697278
rect 155604 697276 156204 697278
rect 191604 697276 192204 697278
rect 227604 697276 228204 697278
rect 263604 697276 264204 697278
rect 299604 697276 300204 697278
rect 335604 697276 336204 697278
rect 371604 697276 372204 697278
rect 407604 697276 408204 697278
rect 443604 697276 444204 697278
rect 479604 697276 480204 697278
rect 515604 697276 516204 697278
rect 551604 697276 552204 697278
rect 590960 697276 591560 697278
rect -8576 697254 592500 697276
rect -8576 697018 -7454 697254
rect -7218 697018 11786 697254
rect 12022 697018 47786 697254
rect 48022 697018 83786 697254
rect 84022 697018 119786 697254
rect 120022 697018 155786 697254
rect 156022 697018 191786 697254
rect 192022 697018 227786 697254
rect 228022 697018 263786 697254
rect 264022 697018 299786 697254
rect 300022 697018 335786 697254
rect 336022 697018 371786 697254
rect 372022 697018 407786 697254
rect 408022 697018 443786 697254
rect 444022 697018 479786 697254
rect 480022 697018 515786 697254
rect 516022 697018 551786 697254
rect 552022 697018 591142 697254
rect 591378 697018 592500 697254
rect -8576 696934 592500 697018
rect -8576 696698 -7454 696934
rect -7218 696698 11786 696934
rect 12022 696698 47786 696934
rect 48022 696698 83786 696934
rect 84022 696698 119786 696934
rect 120022 696698 155786 696934
rect 156022 696698 191786 696934
rect 192022 696698 227786 696934
rect 228022 696698 263786 696934
rect 264022 696698 299786 696934
rect 300022 696698 335786 696934
rect 336022 696698 371786 696934
rect 372022 696698 407786 696934
rect 408022 696698 443786 696934
rect 444022 696698 479786 696934
rect 480022 696698 515786 696934
rect 516022 696698 551786 696934
rect 552022 696698 591142 696934
rect 591378 696698 592500 696934
rect -8576 696676 592500 696698
rect -7636 696674 -7036 696676
rect 11604 696674 12204 696676
rect 47604 696674 48204 696676
rect 83604 696674 84204 696676
rect 119604 696674 120204 696676
rect 155604 696674 156204 696676
rect 191604 696674 192204 696676
rect 227604 696674 228204 696676
rect 263604 696674 264204 696676
rect 299604 696674 300204 696676
rect 335604 696674 336204 696676
rect 371604 696674 372204 696676
rect 407604 696674 408204 696676
rect 443604 696674 444204 696676
rect 479604 696674 480204 696676
rect 515604 696674 516204 696676
rect 551604 696674 552204 696676
rect 590960 696674 591560 696676
rect -5756 693676 -5156 693678
rect 8004 693676 8604 693678
rect 44004 693676 44604 693678
rect 80004 693676 80604 693678
rect 116004 693676 116604 693678
rect 152004 693676 152604 693678
rect 188004 693676 188604 693678
rect 224004 693676 224604 693678
rect 260004 693676 260604 693678
rect 296004 693676 296604 693678
rect 332004 693676 332604 693678
rect 368004 693676 368604 693678
rect 404004 693676 404604 693678
rect 440004 693676 440604 693678
rect 476004 693676 476604 693678
rect 512004 693676 512604 693678
rect 548004 693676 548604 693678
rect 589080 693676 589680 693678
rect -6696 693654 590620 693676
rect -6696 693418 -5574 693654
rect -5338 693418 8186 693654
rect 8422 693418 44186 693654
rect 44422 693418 80186 693654
rect 80422 693418 116186 693654
rect 116422 693418 152186 693654
rect 152422 693418 188186 693654
rect 188422 693418 224186 693654
rect 224422 693418 260186 693654
rect 260422 693418 296186 693654
rect 296422 693418 332186 693654
rect 332422 693418 368186 693654
rect 368422 693418 404186 693654
rect 404422 693418 440186 693654
rect 440422 693418 476186 693654
rect 476422 693418 512186 693654
rect 512422 693418 548186 693654
rect 548422 693418 589262 693654
rect 589498 693418 590620 693654
rect -6696 693334 590620 693418
rect -6696 693098 -5574 693334
rect -5338 693098 8186 693334
rect 8422 693098 44186 693334
rect 44422 693098 80186 693334
rect 80422 693098 116186 693334
rect 116422 693098 152186 693334
rect 152422 693098 188186 693334
rect 188422 693098 224186 693334
rect 224422 693098 260186 693334
rect 260422 693098 296186 693334
rect 296422 693098 332186 693334
rect 332422 693098 368186 693334
rect 368422 693098 404186 693334
rect 404422 693098 440186 693334
rect 440422 693098 476186 693334
rect 476422 693098 512186 693334
rect 512422 693098 548186 693334
rect 548422 693098 589262 693334
rect 589498 693098 590620 693334
rect -6696 693076 590620 693098
rect -5756 693074 -5156 693076
rect 8004 693074 8604 693076
rect 44004 693074 44604 693076
rect 80004 693074 80604 693076
rect 116004 693074 116604 693076
rect 152004 693074 152604 693076
rect 188004 693074 188604 693076
rect 224004 693074 224604 693076
rect 260004 693074 260604 693076
rect 296004 693074 296604 693076
rect 332004 693074 332604 693076
rect 368004 693074 368604 693076
rect 404004 693074 404604 693076
rect 440004 693074 440604 693076
rect 476004 693074 476604 693076
rect 512004 693074 512604 693076
rect 548004 693074 548604 693076
rect 589080 693074 589680 693076
rect -3876 690076 -3276 690078
rect 4404 690076 5004 690078
rect 40404 690076 41004 690078
rect 76404 690076 77004 690078
rect 112404 690076 113004 690078
rect 148404 690076 149004 690078
rect 184404 690076 185004 690078
rect 220404 690076 221004 690078
rect 256404 690076 257004 690078
rect 292404 690076 293004 690078
rect 328404 690076 329004 690078
rect 364404 690076 365004 690078
rect 400404 690076 401004 690078
rect 436404 690076 437004 690078
rect 472404 690076 473004 690078
rect 508404 690076 509004 690078
rect 544404 690076 545004 690078
rect 580404 690076 581004 690078
rect 587200 690076 587800 690078
rect -4816 690054 588740 690076
rect -4816 689818 -3694 690054
rect -3458 689818 4586 690054
rect 4822 689818 40586 690054
rect 40822 689818 76586 690054
rect 76822 689818 112586 690054
rect 112822 689818 148586 690054
rect 148822 689818 184586 690054
rect 184822 689818 220586 690054
rect 220822 689818 256586 690054
rect 256822 689818 292586 690054
rect 292822 689818 328586 690054
rect 328822 689818 364586 690054
rect 364822 689818 400586 690054
rect 400822 689818 436586 690054
rect 436822 689818 472586 690054
rect 472822 689818 508586 690054
rect 508822 689818 544586 690054
rect 544822 689818 580586 690054
rect 580822 689818 587382 690054
rect 587618 689818 588740 690054
rect -4816 689734 588740 689818
rect -4816 689498 -3694 689734
rect -3458 689498 4586 689734
rect 4822 689498 40586 689734
rect 40822 689498 76586 689734
rect 76822 689498 112586 689734
rect 112822 689498 148586 689734
rect 148822 689498 184586 689734
rect 184822 689498 220586 689734
rect 220822 689498 256586 689734
rect 256822 689498 292586 689734
rect 292822 689498 328586 689734
rect 328822 689498 364586 689734
rect 364822 689498 400586 689734
rect 400822 689498 436586 689734
rect 436822 689498 472586 689734
rect 472822 689498 508586 689734
rect 508822 689498 544586 689734
rect 544822 689498 580586 689734
rect 580822 689498 587382 689734
rect 587618 689498 588740 689734
rect -4816 689476 588740 689498
rect -3876 689474 -3276 689476
rect 4404 689474 5004 689476
rect 40404 689474 41004 689476
rect 76404 689474 77004 689476
rect 112404 689474 113004 689476
rect 148404 689474 149004 689476
rect 184404 689474 185004 689476
rect 220404 689474 221004 689476
rect 256404 689474 257004 689476
rect 292404 689474 293004 689476
rect 328404 689474 329004 689476
rect 364404 689474 365004 689476
rect 400404 689474 401004 689476
rect 436404 689474 437004 689476
rect 472404 689474 473004 689476
rect 508404 689474 509004 689476
rect 544404 689474 545004 689476
rect 580404 689474 581004 689476
rect 587200 689474 587800 689476
rect -1996 686476 -1396 686478
rect 804 686476 1404 686478
rect 36804 686476 37404 686478
rect 72804 686476 73404 686478
rect 108804 686476 109404 686478
rect 144804 686476 145404 686478
rect 180804 686476 181404 686478
rect 216804 686476 217404 686478
rect 252804 686476 253404 686478
rect 288804 686476 289404 686478
rect 324804 686476 325404 686478
rect 360804 686476 361404 686478
rect 396804 686476 397404 686478
rect 432804 686476 433404 686478
rect 468804 686476 469404 686478
rect 504804 686476 505404 686478
rect 540804 686476 541404 686478
rect 576804 686476 577404 686478
rect 585320 686476 585920 686478
rect -2936 686454 586860 686476
rect -2936 686218 -1814 686454
rect -1578 686218 986 686454
rect 1222 686218 36986 686454
rect 37222 686218 72986 686454
rect 73222 686218 108986 686454
rect 109222 686218 144986 686454
rect 145222 686218 180986 686454
rect 181222 686218 216986 686454
rect 217222 686218 252986 686454
rect 253222 686218 288986 686454
rect 289222 686218 324986 686454
rect 325222 686218 360986 686454
rect 361222 686218 396986 686454
rect 397222 686218 432986 686454
rect 433222 686218 468986 686454
rect 469222 686218 504986 686454
rect 505222 686218 540986 686454
rect 541222 686218 576986 686454
rect 577222 686218 585502 686454
rect 585738 686218 586860 686454
rect -2936 686134 586860 686218
rect -2936 685898 -1814 686134
rect -1578 685898 986 686134
rect 1222 685898 36986 686134
rect 37222 685898 72986 686134
rect 73222 685898 108986 686134
rect 109222 685898 144986 686134
rect 145222 685898 180986 686134
rect 181222 685898 216986 686134
rect 217222 685898 252986 686134
rect 253222 685898 288986 686134
rect 289222 685898 324986 686134
rect 325222 685898 360986 686134
rect 361222 685898 396986 686134
rect 397222 685898 432986 686134
rect 433222 685898 468986 686134
rect 469222 685898 504986 686134
rect 505222 685898 540986 686134
rect 541222 685898 576986 686134
rect 577222 685898 585502 686134
rect 585738 685898 586860 686134
rect -2936 685876 586860 685898
rect -1996 685874 -1396 685876
rect 804 685874 1404 685876
rect 36804 685874 37404 685876
rect 72804 685874 73404 685876
rect 108804 685874 109404 685876
rect 144804 685874 145404 685876
rect 180804 685874 181404 685876
rect 216804 685874 217404 685876
rect 252804 685874 253404 685876
rect 288804 685874 289404 685876
rect 324804 685874 325404 685876
rect 360804 685874 361404 685876
rect 396804 685874 397404 685876
rect 432804 685874 433404 685876
rect 468804 685874 469404 685876
rect 504804 685874 505404 685876
rect 540804 685874 541404 685876
rect 576804 685874 577404 685876
rect 585320 685874 585920 685876
rect -8576 679276 -7976 679278
rect 29604 679276 30204 679278
rect 65604 679276 66204 679278
rect 101604 679276 102204 679278
rect 137604 679276 138204 679278
rect 173604 679276 174204 679278
rect 209604 679276 210204 679278
rect 245604 679276 246204 679278
rect 281604 679276 282204 679278
rect 317604 679276 318204 679278
rect 353604 679276 354204 679278
rect 389604 679276 390204 679278
rect 425604 679276 426204 679278
rect 461604 679276 462204 679278
rect 497604 679276 498204 679278
rect 533604 679276 534204 679278
rect 569604 679276 570204 679278
rect 591900 679276 592500 679278
rect -8576 679254 592500 679276
rect -8576 679018 -8394 679254
rect -8158 679018 29786 679254
rect 30022 679018 65786 679254
rect 66022 679018 101786 679254
rect 102022 679018 137786 679254
rect 138022 679018 173786 679254
rect 174022 679018 209786 679254
rect 210022 679018 245786 679254
rect 246022 679018 281786 679254
rect 282022 679018 317786 679254
rect 318022 679018 353786 679254
rect 354022 679018 389786 679254
rect 390022 679018 425786 679254
rect 426022 679018 461786 679254
rect 462022 679018 497786 679254
rect 498022 679018 533786 679254
rect 534022 679018 569786 679254
rect 570022 679018 592082 679254
rect 592318 679018 592500 679254
rect -8576 678934 592500 679018
rect -8576 678698 -8394 678934
rect -8158 678698 29786 678934
rect 30022 678698 65786 678934
rect 66022 678698 101786 678934
rect 102022 678698 137786 678934
rect 138022 678698 173786 678934
rect 174022 678698 209786 678934
rect 210022 678698 245786 678934
rect 246022 678698 281786 678934
rect 282022 678698 317786 678934
rect 318022 678698 353786 678934
rect 354022 678698 389786 678934
rect 390022 678698 425786 678934
rect 426022 678698 461786 678934
rect 462022 678698 497786 678934
rect 498022 678698 533786 678934
rect 534022 678698 569786 678934
rect 570022 678698 592082 678934
rect 592318 678698 592500 678934
rect -8576 678676 592500 678698
rect -8576 678674 -7976 678676
rect 29604 678674 30204 678676
rect 65604 678674 66204 678676
rect 101604 678674 102204 678676
rect 137604 678674 138204 678676
rect 173604 678674 174204 678676
rect 209604 678674 210204 678676
rect 245604 678674 246204 678676
rect 281604 678674 282204 678676
rect 317604 678674 318204 678676
rect 353604 678674 354204 678676
rect 389604 678674 390204 678676
rect 425604 678674 426204 678676
rect 461604 678674 462204 678676
rect 497604 678674 498204 678676
rect 533604 678674 534204 678676
rect 569604 678674 570204 678676
rect 591900 678674 592500 678676
rect -6696 675676 -6096 675678
rect 26004 675676 26604 675678
rect 62004 675676 62604 675678
rect 98004 675676 98604 675678
rect 134004 675676 134604 675678
rect 170004 675676 170604 675678
rect 206004 675676 206604 675678
rect 242004 675676 242604 675678
rect 278004 675676 278604 675678
rect 314004 675676 314604 675678
rect 350004 675676 350604 675678
rect 386004 675676 386604 675678
rect 422004 675676 422604 675678
rect 458004 675676 458604 675678
rect 494004 675676 494604 675678
rect 530004 675676 530604 675678
rect 566004 675676 566604 675678
rect 590020 675676 590620 675678
rect -6696 675654 590620 675676
rect -6696 675418 -6514 675654
rect -6278 675418 26186 675654
rect 26422 675418 62186 675654
rect 62422 675418 98186 675654
rect 98422 675418 134186 675654
rect 134422 675418 170186 675654
rect 170422 675418 206186 675654
rect 206422 675418 242186 675654
rect 242422 675418 278186 675654
rect 278422 675418 314186 675654
rect 314422 675418 350186 675654
rect 350422 675418 386186 675654
rect 386422 675418 422186 675654
rect 422422 675418 458186 675654
rect 458422 675418 494186 675654
rect 494422 675418 530186 675654
rect 530422 675418 566186 675654
rect 566422 675418 590202 675654
rect 590438 675418 590620 675654
rect -6696 675334 590620 675418
rect -6696 675098 -6514 675334
rect -6278 675098 26186 675334
rect 26422 675098 62186 675334
rect 62422 675098 98186 675334
rect 98422 675098 134186 675334
rect 134422 675098 170186 675334
rect 170422 675098 206186 675334
rect 206422 675098 242186 675334
rect 242422 675098 278186 675334
rect 278422 675098 314186 675334
rect 314422 675098 350186 675334
rect 350422 675098 386186 675334
rect 386422 675098 422186 675334
rect 422422 675098 458186 675334
rect 458422 675098 494186 675334
rect 494422 675098 530186 675334
rect 530422 675098 566186 675334
rect 566422 675098 590202 675334
rect 590438 675098 590620 675334
rect -6696 675076 590620 675098
rect -6696 675074 -6096 675076
rect 26004 675074 26604 675076
rect 62004 675074 62604 675076
rect 98004 675074 98604 675076
rect 134004 675074 134604 675076
rect 170004 675074 170604 675076
rect 206004 675074 206604 675076
rect 242004 675074 242604 675076
rect 278004 675074 278604 675076
rect 314004 675074 314604 675076
rect 350004 675074 350604 675076
rect 386004 675074 386604 675076
rect 422004 675074 422604 675076
rect 458004 675074 458604 675076
rect 494004 675074 494604 675076
rect 530004 675074 530604 675076
rect 566004 675074 566604 675076
rect 590020 675074 590620 675076
rect -4816 672076 -4216 672078
rect 22404 672076 23004 672078
rect 58404 672076 59004 672078
rect 94404 672076 95004 672078
rect 130404 672076 131004 672078
rect 166404 672076 167004 672078
rect 202404 672076 203004 672078
rect 238404 672076 239004 672078
rect 274404 672076 275004 672078
rect 310404 672076 311004 672078
rect 346404 672076 347004 672078
rect 382404 672076 383004 672078
rect 418404 672076 419004 672078
rect 454404 672076 455004 672078
rect 490404 672076 491004 672078
rect 526404 672076 527004 672078
rect 562404 672076 563004 672078
rect 588140 672076 588740 672078
rect -4816 672054 588740 672076
rect -4816 671818 -4634 672054
rect -4398 671818 22586 672054
rect 22822 671818 58586 672054
rect 58822 671818 94586 672054
rect 94822 671818 130586 672054
rect 130822 671818 166586 672054
rect 166822 671818 202586 672054
rect 202822 671818 238586 672054
rect 238822 671818 274586 672054
rect 274822 671818 310586 672054
rect 310822 671818 346586 672054
rect 346822 671818 382586 672054
rect 382822 671818 418586 672054
rect 418822 671818 454586 672054
rect 454822 671818 490586 672054
rect 490822 671818 526586 672054
rect 526822 671818 562586 672054
rect 562822 671818 588322 672054
rect 588558 671818 588740 672054
rect -4816 671734 588740 671818
rect -4816 671498 -4634 671734
rect -4398 671498 22586 671734
rect 22822 671498 58586 671734
rect 58822 671498 94586 671734
rect 94822 671498 130586 671734
rect 130822 671498 166586 671734
rect 166822 671498 202586 671734
rect 202822 671498 238586 671734
rect 238822 671498 274586 671734
rect 274822 671498 310586 671734
rect 310822 671498 346586 671734
rect 346822 671498 382586 671734
rect 382822 671498 418586 671734
rect 418822 671498 454586 671734
rect 454822 671498 490586 671734
rect 490822 671498 526586 671734
rect 526822 671498 562586 671734
rect 562822 671498 588322 671734
rect 588558 671498 588740 671734
rect -4816 671476 588740 671498
rect -4816 671474 -4216 671476
rect 22404 671474 23004 671476
rect 58404 671474 59004 671476
rect 94404 671474 95004 671476
rect 130404 671474 131004 671476
rect 166404 671474 167004 671476
rect 202404 671474 203004 671476
rect 238404 671474 239004 671476
rect 274404 671474 275004 671476
rect 310404 671474 311004 671476
rect 346404 671474 347004 671476
rect 382404 671474 383004 671476
rect 418404 671474 419004 671476
rect 454404 671474 455004 671476
rect 490404 671474 491004 671476
rect 526404 671474 527004 671476
rect 562404 671474 563004 671476
rect 588140 671474 588740 671476
rect -2936 668476 -2336 668478
rect 18804 668476 19404 668478
rect 54804 668476 55404 668478
rect 90804 668476 91404 668478
rect 126804 668476 127404 668478
rect 162804 668476 163404 668478
rect 198804 668476 199404 668478
rect 234804 668476 235404 668478
rect 270804 668476 271404 668478
rect 306804 668476 307404 668478
rect 342804 668476 343404 668478
rect 378804 668476 379404 668478
rect 414804 668476 415404 668478
rect 450804 668476 451404 668478
rect 486804 668476 487404 668478
rect 522804 668476 523404 668478
rect 558804 668476 559404 668478
rect 586260 668476 586860 668478
rect -2936 668454 586860 668476
rect -2936 668218 -2754 668454
rect -2518 668218 18986 668454
rect 19222 668218 54986 668454
rect 55222 668218 90986 668454
rect 91222 668218 126986 668454
rect 127222 668218 162986 668454
rect 163222 668218 198986 668454
rect 199222 668218 234986 668454
rect 235222 668218 270986 668454
rect 271222 668218 306986 668454
rect 307222 668218 342986 668454
rect 343222 668218 378986 668454
rect 379222 668218 414986 668454
rect 415222 668218 450986 668454
rect 451222 668218 486986 668454
rect 487222 668218 522986 668454
rect 523222 668218 558986 668454
rect 559222 668218 586442 668454
rect 586678 668218 586860 668454
rect -2936 668134 586860 668218
rect -2936 667898 -2754 668134
rect -2518 667898 18986 668134
rect 19222 667898 54986 668134
rect 55222 667898 90986 668134
rect 91222 667898 126986 668134
rect 127222 667898 162986 668134
rect 163222 667898 198986 668134
rect 199222 667898 234986 668134
rect 235222 667898 270986 668134
rect 271222 667898 306986 668134
rect 307222 667898 342986 668134
rect 343222 667898 378986 668134
rect 379222 667898 414986 668134
rect 415222 667898 450986 668134
rect 451222 667898 486986 668134
rect 487222 667898 522986 668134
rect 523222 667898 558986 668134
rect 559222 667898 586442 668134
rect 586678 667898 586860 668134
rect -2936 667876 586860 667898
rect -2936 667874 -2336 667876
rect 18804 667874 19404 667876
rect 54804 667874 55404 667876
rect 90804 667874 91404 667876
rect 126804 667874 127404 667876
rect 162804 667874 163404 667876
rect 198804 667874 199404 667876
rect 234804 667874 235404 667876
rect 270804 667874 271404 667876
rect 306804 667874 307404 667876
rect 342804 667874 343404 667876
rect 378804 667874 379404 667876
rect 414804 667874 415404 667876
rect 450804 667874 451404 667876
rect 486804 667874 487404 667876
rect 522804 667874 523404 667876
rect 558804 667874 559404 667876
rect 586260 667874 586860 667876
rect -7636 661276 -7036 661278
rect 11604 661276 12204 661278
rect 47604 661276 48204 661278
rect 83604 661276 84204 661278
rect 119604 661276 120204 661278
rect 155604 661276 156204 661278
rect 191604 661276 192204 661278
rect 227604 661276 228204 661278
rect 263604 661276 264204 661278
rect 299604 661276 300204 661278
rect 335604 661276 336204 661278
rect 371604 661276 372204 661278
rect 407604 661276 408204 661278
rect 443604 661276 444204 661278
rect 479604 661276 480204 661278
rect 515604 661276 516204 661278
rect 551604 661276 552204 661278
rect 590960 661276 591560 661278
rect -8576 661254 592500 661276
rect -8576 661018 -7454 661254
rect -7218 661018 11786 661254
rect 12022 661018 47786 661254
rect 48022 661018 83786 661254
rect 84022 661018 119786 661254
rect 120022 661018 155786 661254
rect 156022 661018 191786 661254
rect 192022 661018 227786 661254
rect 228022 661018 263786 661254
rect 264022 661018 299786 661254
rect 300022 661018 335786 661254
rect 336022 661018 371786 661254
rect 372022 661018 407786 661254
rect 408022 661018 443786 661254
rect 444022 661018 479786 661254
rect 480022 661018 515786 661254
rect 516022 661018 551786 661254
rect 552022 661018 591142 661254
rect 591378 661018 592500 661254
rect -8576 660934 592500 661018
rect -8576 660698 -7454 660934
rect -7218 660698 11786 660934
rect 12022 660698 47786 660934
rect 48022 660698 83786 660934
rect 84022 660698 119786 660934
rect 120022 660698 155786 660934
rect 156022 660698 191786 660934
rect 192022 660698 227786 660934
rect 228022 660698 263786 660934
rect 264022 660698 299786 660934
rect 300022 660698 335786 660934
rect 336022 660698 371786 660934
rect 372022 660698 407786 660934
rect 408022 660698 443786 660934
rect 444022 660698 479786 660934
rect 480022 660698 515786 660934
rect 516022 660698 551786 660934
rect 552022 660698 591142 660934
rect 591378 660698 592500 660934
rect -8576 660676 592500 660698
rect -7636 660674 -7036 660676
rect 11604 660674 12204 660676
rect 47604 660674 48204 660676
rect 83604 660674 84204 660676
rect 119604 660674 120204 660676
rect 155604 660674 156204 660676
rect 191604 660674 192204 660676
rect 227604 660674 228204 660676
rect 263604 660674 264204 660676
rect 299604 660674 300204 660676
rect 335604 660674 336204 660676
rect 371604 660674 372204 660676
rect 407604 660674 408204 660676
rect 443604 660674 444204 660676
rect 479604 660674 480204 660676
rect 515604 660674 516204 660676
rect 551604 660674 552204 660676
rect 590960 660674 591560 660676
rect -5756 657676 -5156 657678
rect 8004 657676 8604 657678
rect 44004 657676 44604 657678
rect 80004 657676 80604 657678
rect 116004 657676 116604 657678
rect 152004 657676 152604 657678
rect 188004 657676 188604 657678
rect 224004 657676 224604 657678
rect 260004 657676 260604 657678
rect 296004 657676 296604 657678
rect 332004 657676 332604 657678
rect 368004 657676 368604 657678
rect 404004 657676 404604 657678
rect 440004 657676 440604 657678
rect 476004 657676 476604 657678
rect 512004 657676 512604 657678
rect 548004 657676 548604 657678
rect 589080 657676 589680 657678
rect -6696 657654 590620 657676
rect -6696 657418 -5574 657654
rect -5338 657418 8186 657654
rect 8422 657418 44186 657654
rect 44422 657418 80186 657654
rect 80422 657418 116186 657654
rect 116422 657418 152186 657654
rect 152422 657418 188186 657654
rect 188422 657418 224186 657654
rect 224422 657418 260186 657654
rect 260422 657418 296186 657654
rect 296422 657418 332186 657654
rect 332422 657418 368186 657654
rect 368422 657418 404186 657654
rect 404422 657418 440186 657654
rect 440422 657418 476186 657654
rect 476422 657418 512186 657654
rect 512422 657418 548186 657654
rect 548422 657418 589262 657654
rect 589498 657418 590620 657654
rect -6696 657334 590620 657418
rect -6696 657098 -5574 657334
rect -5338 657098 8186 657334
rect 8422 657098 44186 657334
rect 44422 657098 80186 657334
rect 80422 657098 116186 657334
rect 116422 657098 152186 657334
rect 152422 657098 188186 657334
rect 188422 657098 224186 657334
rect 224422 657098 260186 657334
rect 260422 657098 296186 657334
rect 296422 657098 332186 657334
rect 332422 657098 368186 657334
rect 368422 657098 404186 657334
rect 404422 657098 440186 657334
rect 440422 657098 476186 657334
rect 476422 657098 512186 657334
rect 512422 657098 548186 657334
rect 548422 657098 589262 657334
rect 589498 657098 590620 657334
rect -6696 657076 590620 657098
rect -5756 657074 -5156 657076
rect 8004 657074 8604 657076
rect 44004 657074 44604 657076
rect 80004 657074 80604 657076
rect 116004 657074 116604 657076
rect 152004 657074 152604 657076
rect 188004 657074 188604 657076
rect 224004 657074 224604 657076
rect 260004 657074 260604 657076
rect 296004 657074 296604 657076
rect 332004 657074 332604 657076
rect 368004 657074 368604 657076
rect 404004 657074 404604 657076
rect 440004 657074 440604 657076
rect 476004 657074 476604 657076
rect 512004 657074 512604 657076
rect 548004 657074 548604 657076
rect 589080 657074 589680 657076
rect -3876 654076 -3276 654078
rect 4404 654076 5004 654078
rect 40404 654076 41004 654078
rect 76404 654076 77004 654078
rect 112404 654076 113004 654078
rect 148404 654076 149004 654078
rect 184404 654076 185004 654078
rect 220404 654076 221004 654078
rect 256404 654076 257004 654078
rect 292404 654076 293004 654078
rect 328404 654076 329004 654078
rect 364404 654076 365004 654078
rect 400404 654076 401004 654078
rect 436404 654076 437004 654078
rect 472404 654076 473004 654078
rect 508404 654076 509004 654078
rect 544404 654076 545004 654078
rect 580404 654076 581004 654078
rect 587200 654076 587800 654078
rect -4816 654054 588740 654076
rect -4816 653818 -3694 654054
rect -3458 653818 4586 654054
rect 4822 653818 40586 654054
rect 40822 653818 76586 654054
rect 76822 653818 112586 654054
rect 112822 653818 148586 654054
rect 148822 653818 184586 654054
rect 184822 653818 220586 654054
rect 220822 653818 256586 654054
rect 256822 653818 292586 654054
rect 292822 653818 328586 654054
rect 328822 653818 364586 654054
rect 364822 653818 400586 654054
rect 400822 653818 436586 654054
rect 436822 653818 472586 654054
rect 472822 653818 508586 654054
rect 508822 653818 544586 654054
rect 544822 653818 580586 654054
rect 580822 653818 587382 654054
rect 587618 653818 588740 654054
rect -4816 653734 588740 653818
rect -4816 653498 -3694 653734
rect -3458 653498 4586 653734
rect 4822 653498 40586 653734
rect 40822 653498 76586 653734
rect 76822 653498 112586 653734
rect 112822 653498 148586 653734
rect 148822 653498 184586 653734
rect 184822 653498 220586 653734
rect 220822 653498 256586 653734
rect 256822 653498 292586 653734
rect 292822 653498 328586 653734
rect 328822 653498 364586 653734
rect 364822 653498 400586 653734
rect 400822 653498 436586 653734
rect 436822 653498 472586 653734
rect 472822 653498 508586 653734
rect 508822 653498 544586 653734
rect 544822 653498 580586 653734
rect 580822 653498 587382 653734
rect 587618 653498 588740 653734
rect -4816 653476 588740 653498
rect -3876 653474 -3276 653476
rect 4404 653474 5004 653476
rect 40404 653474 41004 653476
rect 76404 653474 77004 653476
rect 112404 653474 113004 653476
rect 148404 653474 149004 653476
rect 184404 653474 185004 653476
rect 220404 653474 221004 653476
rect 256404 653474 257004 653476
rect 292404 653474 293004 653476
rect 328404 653474 329004 653476
rect 364404 653474 365004 653476
rect 400404 653474 401004 653476
rect 436404 653474 437004 653476
rect 472404 653474 473004 653476
rect 508404 653474 509004 653476
rect 544404 653474 545004 653476
rect 580404 653474 581004 653476
rect 587200 653474 587800 653476
rect -1996 650476 -1396 650478
rect 804 650476 1404 650478
rect 36804 650476 37404 650478
rect 72804 650476 73404 650478
rect 108804 650476 109404 650478
rect 144804 650476 145404 650478
rect 180804 650476 181404 650478
rect 216804 650476 217404 650478
rect 252804 650476 253404 650478
rect 288804 650476 289404 650478
rect 324804 650476 325404 650478
rect 360804 650476 361404 650478
rect 396804 650476 397404 650478
rect 432804 650476 433404 650478
rect 468804 650476 469404 650478
rect 504804 650476 505404 650478
rect 540804 650476 541404 650478
rect 576804 650476 577404 650478
rect 585320 650476 585920 650478
rect -2936 650454 586860 650476
rect -2936 650218 -1814 650454
rect -1578 650218 986 650454
rect 1222 650218 36986 650454
rect 37222 650218 72986 650454
rect 73222 650218 108986 650454
rect 109222 650218 144986 650454
rect 145222 650218 180986 650454
rect 181222 650218 216986 650454
rect 217222 650218 252986 650454
rect 253222 650218 288986 650454
rect 289222 650218 324986 650454
rect 325222 650218 360986 650454
rect 361222 650218 396986 650454
rect 397222 650218 432986 650454
rect 433222 650218 468986 650454
rect 469222 650218 504986 650454
rect 505222 650218 540986 650454
rect 541222 650218 576986 650454
rect 577222 650218 585502 650454
rect 585738 650218 586860 650454
rect -2936 650134 586860 650218
rect -2936 649898 -1814 650134
rect -1578 649898 986 650134
rect 1222 649898 36986 650134
rect 37222 649898 72986 650134
rect 73222 649898 108986 650134
rect 109222 649898 144986 650134
rect 145222 649898 180986 650134
rect 181222 649898 216986 650134
rect 217222 649898 252986 650134
rect 253222 649898 288986 650134
rect 289222 649898 324986 650134
rect 325222 649898 360986 650134
rect 361222 649898 396986 650134
rect 397222 649898 432986 650134
rect 433222 649898 468986 650134
rect 469222 649898 504986 650134
rect 505222 649898 540986 650134
rect 541222 649898 576986 650134
rect 577222 649898 585502 650134
rect 585738 649898 586860 650134
rect -2936 649876 586860 649898
rect -1996 649874 -1396 649876
rect 804 649874 1404 649876
rect 36804 649874 37404 649876
rect 72804 649874 73404 649876
rect 108804 649874 109404 649876
rect 144804 649874 145404 649876
rect 180804 649874 181404 649876
rect 216804 649874 217404 649876
rect 252804 649874 253404 649876
rect 288804 649874 289404 649876
rect 324804 649874 325404 649876
rect 360804 649874 361404 649876
rect 396804 649874 397404 649876
rect 432804 649874 433404 649876
rect 468804 649874 469404 649876
rect 504804 649874 505404 649876
rect 540804 649874 541404 649876
rect 576804 649874 577404 649876
rect 585320 649874 585920 649876
rect -8576 643276 -7976 643278
rect 29604 643276 30204 643278
rect 65604 643276 66204 643278
rect 101604 643276 102204 643278
rect 137604 643276 138204 643278
rect 173604 643276 174204 643278
rect 209604 643276 210204 643278
rect 245604 643276 246204 643278
rect 281604 643276 282204 643278
rect 317604 643276 318204 643278
rect 353604 643276 354204 643278
rect 389604 643276 390204 643278
rect 425604 643276 426204 643278
rect 461604 643276 462204 643278
rect 497604 643276 498204 643278
rect 533604 643276 534204 643278
rect 569604 643276 570204 643278
rect 591900 643276 592500 643278
rect -8576 643254 592500 643276
rect -8576 643018 -8394 643254
rect -8158 643018 29786 643254
rect 30022 643018 65786 643254
rect 66022 643018 101786 643254
rect 102022 643018 137786 643254
rect 138022 643018 173786 643254
rect 174022 643018 209786 643254
rect 210022 643018 245786 643254
rect 246022 643018 281786 643254
rect 282022 643018 317786 643254
rect 318022 643018 353786 643254
rect 354022 643018 389786 643254
rect 390022 643018 425786 643254
rect 426022 643018 461786 643254
rect 462022 643018 497786 643254
rect 498022 643018 533786 643254
rect 534022 643018 569786 643254
rect 570022 643018 592082 643254
rect 592318 643018 592500 643254
rect -8576 642934 592500 643018
rect -8576 642698 -8394 642934
rect -8158 642698 29786 642934
rect 30022 642698 65786 642934
rect 66022 642698 101786 642934
rect 102022 642698 137786 642934
rect 138022 642698 173786 642934
rect 174022 642698 209786 642934
rect 210022 642698 245786 642934
rect 246022 642698 281786 642934
rect 282022 642698 317786 642934
rect 318022 642698 353786 642934
rect 354022 642698 389786 642934
rect 390022 642698 425786 642934
rect 426022 642698 461786 642934
rect 462022 642698 497786 642934
rect 498022 642698 533786 642934
rect 534022 642698 569786 642934
rect 570022 642698 592082 642934
rect 592318 642698 592500 642934
rect -8576 642676 592500 642698
rect -8576 642674 -7976 642676
rect 29604 642674 30204 642676
rect 65604 642674 66204 642676
rect 101604 642674 102204 642676
rect 137604 642674 138204 642676
rect 173604 642674 174204 642676
rect 209604 642674 210204 642676
rect 245604 642674 246204 642676
rect 281604 642674 282204 642676
rect 317604 642674 318204 642676
rect 353604 642674 354204 642676
rect 389604 642674 390204 642676
rect 425604 642674 426204 642676
rect 461604 642674 462204 642676
rect 497604 642674 498204 642676
rect 533604 642674 534204 642676
rect 569604 642674 570204 642676
rect 591900 642674 592500 642676
rect -6696 639676 -6096 639678
rect 26004 639676 26604 639678
rect 62004 639676 62604 639678
rect 98004 639676 98604 639678
rect 134004 639676 134604 639678
rect 170004 639676 170604 639678
rect 206004 639676 206604 639678
rect 242004 639676 242604 639678
rect 278004 639676 278604 639678
rect 314004 639676 314604 639678
rect 350004 639676 350604 639678
rect 386004 639676 386604 639678
rect 422004 639676 422604 639678
rect 458004 639676 458604 639678
rect 494004 639676 494604 639678
rect 530004 639676 530604 639678
rect 566004 639676 566604 639678
rect 590020 639676 590620 639678
rect -6696 639654 590620 639676
rect -6696 639418 -6514 639654
rect -6278 639418 26186 639654
rect 26422 639418 62186 639654
rect 62422 639418 98186 639654
rect 98422 639418 134186 639654
rect 134422 639418 170186 639654
rect 170422 639418 206186 639654
rect 206422 639418 242186 639654
rect 242422 639418 278186 639654
rect 278422 639418 314186 639654
rect 314422 639418 350186 639654
rect 350422 639418 386186 639654
rect 386422 639418 422186 639654
rect 422422 639418 458186 639654
rect 458422 639418 494186 639654
rect 494422 639418 530186 639654
rect 530422 639418 566186 639654
rect 566422 639418 590202 639654
rect 590438 639418 590620 639654
rect -6696 639334 590620 639418
rect -6696 639098 -6514 639334
rect -6278 639098 26186 639334
rect 26422 639098 62186 639334
rect 62422 639098 98186 639334
rect 98422 639098 134186 639334
rect 134422 639098 170186 639334
rect 170422 639098 206186 639334
rect 206422 639098 242186 639334
rect 242422 639098 278186 639334
rect 278422 639098 314186 639334
rect 314422 639098 350186 639334
rect 350422 639098 386186 639334
rect 386422 639098 422186 639334
rect 422422 639098 458186 639334
rect 458422 639098 494186 639334
rect 494422 639098 530186 639334
rect 530422 639098 566186 639334
rect 566422 639098 590202 639334
rect 590438 639098 590620 639334
rect -6696 639076 590620 639098
rect -6696 639074 -6096 639076
rect 26004 639074 26604 639076
rect 62004 639074 62604 639076
rect 98004 639074 98604 639076
rect 134004 639074 134604 639076
rect 170004 639074 170604 639076
rect 206004 639074 206604 639076
rect 242004 639074 242604 639076
rect 278004 639074 278604 639076
rect 314004 639074 314604 639076
rect 350004 639074 350604 639076
rect 386004 639074 386604 639076
rect 422004 639074 422604 639076
rect 458004 639074 458604 639076
rect 494004 639074 494604 639076
rect 530004 639074 530604 639076
rect 566004 639074 566604 639076
rect 590020 639074 590620 639076
rect -4816 636076 -4216 636078
rect 22404 636076 23004 636078
rect 58404 636076 59004 636078
rect 94404 636076 95004 636078
rect 130404 636076 131004 636078
rect 166404 636076 167004 636078
rect 202404 636076 203004 636078
rect 238404 636076 239004 636078
rect 274404 636076 275004 636078
rect 310404 636076 311004 636078
rect 346404 636076 347004 636078
rect 382404 636076 383004 636078
rect 418404 636076 419004 636078
rect 454404 636076 455004 636078
rect 490404 636076 491004 636078
rect 526404 636076 527004 636078
rect 562404 636076 563004 636078
rect 588140 636076 588740 636078
rect -4816 636054 588740 636076
rect -4816 635818 -4634 636054
rect -4398 635818 22586 636054
rect 22822 635818 58586 636054
rect 58822 635818 94586 636054
rect 94822 635818 130586 636054
rect 130822 635818 166586 636054
rect 166822 635818 202586 636054
rect 202822 635818 238586 636054
rect 238822 635818 274586 636054
rect 274822 635818 310586 636054
rect 310822 635818 346586 636054
rect 346822 635818 382586 636054
rect 382822 635818 418586 636054
rect 418822 635818 454586 636054
rect 454822 635818 490586 636054
rect 490822 635818 526586 636054
rect 526822 635818 562586 636054
rect 562822 635818 588322 636054
rect 588558 635818 588740 636054
rect -4816 635734 588740 635818
rect -4816 635498 -4634 635734
rect -4398 635498 22586 635734
rect 22822 635498 58586 635734
rect 58822 635498 94586 635734
rect 94822 635498 130586 635734
rect 130822 635498 166586 635734
rect 166822 635498 202586 635734
rect 202822 635498 238586 635734
rect 238822 635498 274586 635734
rect 274822 635498 310586 635734
rect 310822 635498 346586 635734
rect 346822 635498 382586 635734
rect 382822 635498 418586 635734
rect 418822 635498 454586 635734
rect 454822 635498 490586 635734
rect 490822 635498 526586 635734
rect 526822 635498 562586 635734
rect 562822 635498 588322 635734
rect 588558 635498 588740 635734
rect -4816 635476 588740 635498
rect -4816 635474 -4216 635476
rect 22404 635474 23004 635476
rect 58404 635474 59004 635476
rect 94404 635474 95004 635476
rect 130404 635474 131004 635476
rect 166404 635474 167004 635476
rect 202404 635474 203004 635476
rect 238404 635474 239004 635476
rect 274404 635474 275004 635476
rect 310404 635474 311004 635476
rect 346404 635474 347004 635476
rect 382404 635474 383004 635476
rect 418404 635474 419004 635476
rect 454404 635474 455004 635476
rect 490404 635474 491004 635476
rect 526404 635474 527004 635476
rect 562404 635474 563004 635476
rect 588140 635474 588740 635476
rect -2936 632476 -2336 632478
rect 18804 632476 19404 632478
rect 54804 632476 55404 632478
rect 90804 632476 91404 632478
rect 126804 632476 127404 632478
rect 162804 632476 163404 632478
rect 198804 632476 199404 632478
rect 234804 632476 235404 632478
rect 270804 632476 271404 632478
rect 306804 632476 307404 632478
rect 342804 632476 343404 632478
rect 378804 632476 379404 632478
rect 414804 632476 415404 632478
rect 450804 632476 451404 632478
rect 486804 632476 487404 632478
rect 522804 632476 523404 632478
rect 558804 632476 559404 632478
rect 586260 632476 586860 632478
rect -2936 632454 586860 632476
rect -2936 632218 -2754 632454
rect -2518 632218 18986 632454
rect 19222 632218 54986 632454
rect 55222 632218 90986 632454
rect 91222 632218 126986 632454
rect 127222 632218 162986 632454
rect 163222 632218 198986 632454
rect 199222 632218 234986 632454
rect 235222 632218 270986 632454
rect 271222 632218 306986 632454
rect 307222 632218 342986 632454
rect 343222 632218 378986 632454
rect 379222 632218 414986 632454
rect 415222 632218 450986 632454
rect 451222 632218 486986 632454
rect 487222 632218 522986 632454
rect 523222 632218 558986 632454
rect 559222 632218 586442 632454
rect 586678 632218 586860 632454
rect -2936 632134 586860 632218
rect -2936 631898 -2754 632134
rect -2518 631898 18986 632134
rect 19222 631898 54986 632134
rect 55222 631898 90986 632134
rect 91222 631898 126986 632134
rect 127222 631898 162986 632134
rect 163222 631898 198986 632134
rect 199222 631898 234986 632134
rect 235222 631898 270986 632134
rect 271222 631898 306986 632134
rect 307222 631898 342986 632134
rect 343222 631898 378986 632134
rect 379222 631898 414986 632134
rect 415222 631898 450986 632134
rect 451222 631898 486986 632134
rect 487222 631898 522986 632134
rect 523222 631898 558986 632134
rect 559222 631898 586442 632134
rect 586678 631898 586860 632134
rect -2936 631876 586860 631898
rect -2936 631874 -2336 631876
rect 18804 631874 19404 631876
rect 54804 631874 55404 631876
rect 90804 631874 91404 631876
rect 126804 631874 127404 631876
rect 162804 631874 163404 631876
rect 198804 631874 199404 631876
rect 234804 631874 235404 631876
rect 270804 631874 271404 631876
rect 306804 631874 307404 631876
rect 342804 631874 343404 631876
rect 378804 631874 379404 631876
rect 414804 631874 415404 631876
rect 450804 631874 451404 631876
rect 486804 631874 487404 631876
rect 522804 631874 523404 631876
rect 558804 631874 559404 631876
rect 586260 631874 586860 631876
rect -7636 625276 -7036 625278
rect 11604 625276 12204 625278
rect 47604 625276 48204 625278
rect 83604 625276 84204 625278
rect 119604 625276 120204 625278
rect 155604 625276 156204 625278
rect 191604 625276 192204 625278
rect 227604 625276 228204 625278
rect 263604 625276 264204 625278
rect 299604 625276 300204 625278
rect 335604 625276 336204 625278
rect 371604 625276 372204 625278
rect 407604 625276 408204 625278
rect 443604 625276 444204 625278
rect 479604 625276 480204 625278
rect 515604 625276 516204 625278
rect 551604 625276 552204 625278
rect 590960 625276 591560 625278
rect -8576 625254 592500 625276
rect -8576 625018 -7454 625254
rect -7218 625018 11786 625254
rect 12022 625018 47786 625254
rect 48022 625018 83786 625254
rect 84022 625018 119786 625254
rect 120022 625018 155786 625254
rect 156022 625018 191786 625254
rect 192022 625018 227786 625254
rect 228022 625018 263786 625254
rect 264022 625018 299786 625254
rect 300022 625018 335786 625254
rect 336022 625018 371786 625254
rect 372022 625018 407786 625254
rect 408022 625018 443786 625254
rect 444022 625018 479786 625254
rect 480022 625018 515786 625254
rect 516022 625018 551786 625254
rect 552022 625018 591142 625254
rect 591378 625018 592500 625254
rect -8576 624934 592500 625018
rect -8576 624698 -7454 624934
rect -7218 624698 11786 624934
rect 12022 624698 47786 624934
rect 48022 624698 83786 624934
rect 84022 624698 119786 624934
rect 120022 624698 155786 624934
rect 156022 624698 191786 624934
rect 192022 624698 227786 624934
rect 228022 624698 263786 624934
rect 264022 624698 299786 624934
rect 300022 624698 335786 624934
rect 336022 624698 371786 624934
rect 372022 624698 407786 624934
rect 408022 624698 443786 624934
rect 444022 624698 479786 624934
rect 480022 624698 515786 624934
rect 516022 624698 551786 624934
rect 552022 624698 591142 624934
rect 591378 624698 592500 624934
rect -8576 624676 592500 624698
rect -7636 624674 -7036 624676
rect 11604 624674 12204 624676
rect 47604 624674 48204 624676
rect 83604 624674 84204 624676
rect 119604 624674 120204 624676
rect 155604 624674 156204 624676
rect 191604 624674 192204 624676
rect 227604 624674 228204 624676
rect 263604 624674 264204 624676
rect 299604 624674 300204 624676
rect 335604 624674 336204 624676
rect 371604 624674 372204 624676
rect 407604 624674 408204 624676
rect 443604 624674 444204 624676
rect 479604 624674 480204 624676
rect 515604 624674 516204 624676
rect 551604 624674 552204 624676
rect 590960 624674 591560 624676
rect -5756 621676 -5156 621678
rect 8004 621676 8604 621678
rect 44004 621676 44604 621678
rect 80004 621676 80604 621678
rect 116004 621676 116604 621678
rect 152004 621676 152604 621678
rect 188004 621676 188604 621678
rect 224004 621676 224604 621678
rect 260004 621676 260604 621678
rect 296004 621676 296604 621678
rect 332004 621676 332604 621678
rect 368004 621676 368604 621678
rect 404004 621676 404604 621678
rect 440004 621676 440604 621678
rect 476004 621676 476604 621678
rect 512004 621676 512604 621678
rect 548004 621676 548604 621678
rect 589080 621676 589680 621678
rect -6696 621654 590620 621676
rect -6696 621418 -5574 621654
rect -5338 621418 8186 621654
rect 8422 621418 44186 621654
rect 44422 621418 80186 621654
rect 80422 621418 116186 621654
rect 116422 621418 152186 621654
rect 152422 621418 188186 621654
rect 188422 621418 224186 621654
rect 224422 621418 260186 621654
rect 260422 621418 296186 621654
rect 296422 621418 332186 621654
rect 332422 621418 368186 621654
rect 368422 621418 404186 621654
rect 404422 621418 440186 621654
rect 440422 621418 476186 621654
rect 476422 621418 512186 621654
rect 512422 621418 548186 621654
rect 548422 621418 589262 621654
rect 589498 621418 590620 621654
rect -6696 621334 590620 621418
rect -6696 621098 -5574 621334
rect -5338 621098 8186 621334
rect 8422 621098 44186 621334
rect 44422 621098 80186 621334
rect 80422 621098 116186 621334
rect 116422 621098 152186 621334
rect 152422 621098 188186 621334
rect 188422 621098 224186 621334
rect 224422 621098 260186 621334
rect 260422 621098 296186 621334
rect 296422 621098 332186 621334
rect 332422 621098 368186 621334
rect 368422 621098 404186 621334
rect 404422 621098 440186 621334
rect 440422 621098 476186 621334
rect 476422 621098 512186 621334
rect 512422 621098 548186 621334
rect 548422 621098 589262 621334
rect 589498 621098 590620 621334
rect -6696 621076 590620 621098
rect -5756 621074 -5156 621076
rect 8004 621074 8604 621076
rect 44004 621074 44604 621076
rect 80004 621074 80604 621076
rect 116004 621074 116604 621076
rect 152004 621074 152604 621076
rect 188004 621074 188604 621076
rect 224004 621074 224604 621076
rect 260004 621074 260604 621076
rect 296004 621074 296604 621076
rect 332004 621074 332604 621076
rect 368004 621074 368604 621076
rect 404004 621074 404604 621076
rect 440004 621074 440604 621076
rect 476004 621074 476604 621076
rect 512004 621074 512604 621076
rect 548004 621074 548604 621076
rect 589080 621074 589680 621076
rect -3876 618076 -3276 618078
rect 4404 618076 5004 618078
rect 40404 618076 41004 618078
rect 76404 618076 77004 618078
rect 112404 618076 113004 618078
rect 148404 618076 149004 618078
rect 184404 618076 185004 618078
rect 220404 618076 221004 618078
rect 256404 618076 257004 618078
rect 292404 618076 293004 618078
rect 328404 618076 329004 618078
rect 364404 618076 365004 618078
rect 400404 618076 401004 618078
rect 436404 618076 437004 618078
rect 472404 618076 473004 618078
rect 508404 618076 509004 618078
rect 544404 618076 545004 618078
rect 580404 618076 581004 618078
rect 587200 618076 587800 618078
rect -4816 618054 588740 618076
rect -4816 617818 -3694 618054
rect -3458 617818 4586 618054
rect 4822 617818 40586 618054
rect 40822 617818 76586 618054
rect 76822 617818 112586 618054
rect 112822 617818 148586 618054
rect 148822 617818 184586 618054
rect 184822 617818 220586 618054
rect 220822 617818 256586 618054
rect 256822 617818 292586 618054
rect 292822 617818 328586 618054
rect 328822 617818 364586 618054
rect 364822 617818 400586 618054
rect 400822 617818 436586 618054
rect 436822 617818 472586 618054
rect 472822 617818 508586 618054
rect 508822 617818 544586 618054
rect 544822 617818 580586 618054
rect 580822 617818 587382 618054
rect 587618 617818 588740 618054
rect -4816 617734 588740 617818
rect -4816 617498 -3694 617734
rect -3458 617498 4586 617734
rect 4822 617498 40586 617734
rect 40822 617498 76586 617734
rect 76822 617498 112586 617734
rect 112822 617498 148586 617734
rect 148822 617498 184586 617734
rect 184822 617498 220586 617734
rect 220822 617498 256586 617734
rect 256822 617498 292586 617734
rect 292822 617498 328586 617734
rect 328822 617498 364586 617734
rect 364822 617498 400586 617734
rect 400822 617498 436586 617734
rect 436822 617498 472586 617734
rect 472822 617498 508586 617734
rect 508822 617498 544586 617734
rect 544822 617498 580586 617734
rect 580822 617498 587382 617734
rect 587618 617498 588740 617734
rect -4816 617476 588740 617498
rect -3876 617474 -3276 617476
rect 4404 617474 5004 617476
rect 40404 617474 41004 617476
rect 76404 617474 77004 617476
rect 112404 617474 113004 617476
rect 148404 617474 149004 617476
rect 184404 617474 185004 617476
rect 220404 617474 221004 617476
rect 256404 617474 257004 617476
rect 292404 617474 293004 617476
rect 328404 617474 329004 617476
rect 364404 617474 365004 617476
rect 400404 617474 401004 617476
rect 436404 617474 437004 617476
rect 472404 617474 473004 617476
rect 508404 617474 509004 617476
rect 544404 617474 545004 617476
rect 580404 617474 581004 617476
rect 587200 617474 587800 617476
rect -1996 614476 -1396 614478
rect 804 614476 1404 614478
rect 36804 614476 37404 614478
rect 72804 614476 73404 614478
rect 108804 614476 109404 614478
rect 144804 614476 145404 614478
rect 180804 614476 181404 614478
rect 216804 614476 217404 614478
rect 252804 614476 253404 614478
rect 288804 614476 289404 614478
rect 396804 614476 397404 614478
rect 504804 614476 505404 614478
rect 540804 614476 541404 614478
rect 576804 614476 577404 614478
rect 585320 614476 585920 614478
rect -2936 614454 586860 614476
rect -2936 614218 -1814 614454
rect -1578 614218 986 614454
rect 1222 614218 36986 614454
rect 37222 614218 72986 614454
rect 73222 614218 108986 614454
rect 109222 614218 144986 614454
rect 145222 614218 180986 614454
rect 181222 614218 216986 614454
rect 217222 614218 252986 614454
rect 253222 614218 288986 614454
rect 289222 614218 396986 614454
rect 397222 614218 504986 614454
rect 505222 614218 540986 614454
rect 541222 614218 576986 614454
rect 577222 614218 585502 614454
rect 585738 614218 586860 614454
rect -2936 614134 586860 614218
rect -2936 613898 -1814 614134
rect -1578 613898 986 614134
rect 1222 613898 36986 614134
rect 37222 613898 72986 614134
rect 73222 613898 108986 614134
rect 109222 613898 144986 614134
rect 145222 613898 180986 614134
rect 181222 613898 216986 614134
rect 217222 613898 252986 614134
rect 253222 613898 288986 614134
rect 289222 613898 396986 614134
rect 397222 613898 504986 614134
rect 505222 613898 540986 614134
rect 541222 613898 576986 614134
rect 577222 613898 585502 614134
rect 585738 613898 586860 614134
rect -2936 613876 586860 613898
rect -1996 613874 -1396 613876
rect 804 613874 1404 613876
rect 36804 613874 37404 613876
rect 72804 613874 73404 613876
rect 108804 613874 109404 613876
rect 144804 613874 145404 613876
rect 180804 613874 181404 613876
rect 216804 613874 217404 613876
rect 252804 613874 253404 613876
rect 288804 613874 289404 613876
rect 396804 613874 397404 613876
rect 504804 613874 505404 613876
rect 540804 613874 541404 613876
rect 576804 613874 577404 613876
rect 585320 613874 585920 613876
rect -8576 607276 -7976 607278
rect 29604 607276 30204 607278
rect 65604 607276 66204 607278
rect 101604 607276 102204 607278
rect 137604 607276 138204 607278
rect 173604 607276 174204 607278
rect 209604 607276 210204 607278
rect 245604 607276 246204 607278
rect 281604 607276 282204 607278
rect 389604 607276 390204 607278
rect 533604 607276 534204 607278
rect 569604 607276 570204 607278
rect 591900 607276 592500 607278
rect -8576 607254 592500 607276
rect -8576 607018 -8394 607254
rect -8158 607018 29786 607254
rect 30022 607018 65786 607254
rect 66022 607018 101786 607254
rect 102022 607018 137786 607254
rect 138022 607018 173786 607254
rect 174022 607018 209786 607254
rect 210022 607018 245786 607254
rect 246022 607018 281786 607254
rect 282022 607018 389786 607254
rect 390022 607018 533786 607254
rect 534022 607018 569786 607254
rect 570022 607018 592082 607254
rect 592318 607018 592500 607254
rect -8576 606934 592500 607018
rect -8576 606698 -8394 606934
rect -8158 606698 29786 606934
rect 30022 606698 65786 606934
rect 66022 606698 101786 606934
rect 102022 606698 137786 606934
rect 138022 606698 173786 606934
rect 174022 606698 209786 606934
rect 210022 606698 245786 606934
rect 246022 606698 281786 606934
rect 282022 606698 389786 606934
rect 390022 606698 533786 606934
rect 534022 606698 569786 606934
rect 570022 606698 592082 606934
rect 592318 606698 592500 606934
rect -8576 606676 592500 606698
rect -8576 606674 -7976 606676
rect 29604 606674 30204 606676
rect 65604 606674 66204 606676
rect 101604 606674 102204 606676
rect 137604 606674 138204 606676
rect 173604 606674 174204 606676
rect 209604 606674 210204 606676
rect 245604 606674 246204 606676
rect 281604 606674 282204 606676
rect 389604 606674 390204 606676
rect 533604 606674 534204 606676
rect 569604 606674 570204 606676
rect 591900 606674 592500 606676
rect -6696 603676 -6096 603678
rect 26004 603676 26604 603678
rect 62004 603676 62604 603678
rect 98004 603676 98604 603678
rect 134004 603676 134604 603678
rect 170004 603676 170604 603678
rect 206004 603676 206604 603678
rect 242004 603676 242604 603678
rect 278004 603676 278604 603678
rect 386004 603676 386604 603678
rect 530004 603676 530604 603678
rect 566004 603676 566604 603678
rect 590020 603676 590620 603678
rect -6696 603654 590620 603676
rect -6696 603418 -6514 603654
rect -6278 603418 26186 603654
rect 26422 603418 62186 603654
rect 62422 603418 98186 603654
rect 98422 603418 134186 603654
rect 134422 603418 170186 603654
rect 170422 603418 206186 603654
rect 206422 603418 242186 603654
rect 242422 603418 278186 603654
rect 278422 603418 386186 603654
rect 386422 603418 530186 603654
rect 530422 603418 566186 603654
rect 566422 603418 590202 603654
rect 590438 603418 590620 603654
rect -6696 603334 590620 603418
rect -6696 603098 -6514 603334
rect -6278 603098 26186 603334
rect 26422 603098 62186 603334
rect 62422 603098 98186 603334
rect 98422 603098 134186 603334
rect 134422 603098 170186 603334
rect 170422 603098 206186 603334
rect 206422 603098 242186 603334
rect 242422 603098 278186 603334
rect 278422 603098 386186 603334
rect 386422 603098 530186 603334
rect 530422 603098 566186 603334
rect 566422 603098 590202 603334
rect 590438 603098 590620 603334
rect -6696 603076 590620 603098
rect -6696 603074 -6096 603076
rect 26004 603074 26604 603076
rect 62004 603074 62604 603076
rect 98004 603074 98604 603076
rect 134004 603074 134604 603076
rect 170004 603074 170604 603076
rect 206004 603074 206604 603076
rect 242004 603074 242604 603076
rect 278004 603074 278604 603076
rect 386004 603074 386604 603076
rect 530004 603074 530604 603076
rect 566004 603074 566604 603076
rect 590020 603074 590620 603076
rect -4816 600076 -4216 600078
rect 22404 600076 23004 600078
rect 58404 600076 59004 600078
rect 94404 600076 95004 600078
rect 130404 600076 131004 600078
rect 166404 600076 167004 600078
rect 202404 600076 203004 600078
rect 238404 600076 239004 600078
rect 274404 600076 275004 600078
rect 382404 600076 383004 600078
rect 526404 600076 527004 600078
rect 562404 600076 563004 600078
rect 588140 600076 588740 600078
rect -4816 600054 588740 600076
rect -4816 599818 -4634 600054
rect -4398 599818 22586 600054
rect 22822 599818 58586 600054
rect 58822 599818 94586 600054
rect 94822 599818 130586 600054
rect 130822 599818 166586 600054
rect 166822 599818 202586 600054
rect 202822 599818 238586 600054
rect 238822 599818 274586 600054
rect 274822 599818 382586 600054
rect 382822 599818 526586 600054
rect 526822 599818 562586 600054
rect 562822 599818 588322 600054
rect 588558 599818 588740 600054
rect -4816 599734 588740 599818
rect -4816 599498 -4634 599734
rect -4398 599498 22586 599734
rect 22822 599498 58586 599734
rect 58822 599498 94586 599734
rect 94822 599498 130586 599734
rect 130822 599498 166586 599734
rect 166822 599498 202586 599734
rect 202822 599498 238586 599734
rect 238822 599498 274586 599734
rect 274822 599498 382586 599734
rect 382822 599498 526586 599734
rect 526822 599498 562586 599734
rect 562822 599498 588322 599734
rect 588558 599498 588740 599734
rect -4816 599476 588740 599498
rect -4816 599474 -4216 599476
rect 22404 599474 23004 599476
rect 58404 599474 59004 599476
rect 94404 599474 95004 599476
rect 130404 599474 131004 599476
rect 166404 599474 167004 599476
rect 202404 599474 203004 599476
rect 238404 599474 239004 599476
rect 274404 599474 275004 599476
rect 382404 599474 383004 599476
rect 526404 599474 527004 599476
rect 562404 599474 563004 599476
rect 588140 599474 588740 599476
rect -2936 596476 -2336 596478
rect 18804 596476 19404 596478
rect 54804 596476 55404 596478
rect 90804 596476 91404 596478
rect 126804 596476 127404 596478
rect 162804 596476 163404 596478
rect 198804 596476 199404 596478
rect 234804 596476 235404 596478
rect 270804 596476 271404 596478
rect 376938 596476 377262 596478
rect 414804 596476 415404 596478
rect 496938 596476 497262 596478
rect 522804 596476 523404 596478
rect 558804 596476 559404 596478
rect 586260 596476 586860 596478
rect -2936 596454 586860 596476
rect -2936 596218 -2754 596454
rect -2518 596218 18986 596454
rect 19222 596218 54986 596454
rect 55222 596218 90986 596454
rect 91222 596218 126986 596454
rect 127222 596218 162986 596454
rect 163222 596218 198986 596454
rect 199222 596218 234986 596454
rect 235222 596218 270986 596454
rect 271222 596218 376982 596454
rect 377218 596218 414986 596454
rect 415222 596218 496982 596454
rect 497218 596218 522986 596454
rect 523222 596218 558986 596454
rect 559222 596218 586442 596454
rect 586678 596218 586860 596454
rect -2936 596134 586860 596218
rect -2936 595898 -2754 596134
rect -2518 595898 18986 596134
rect 19222 595898 54986 596134
rect 55222 595898 90986 596134
rect 91222 595898 126986 596134
rect 127222 595898 162986 596134
rect 163222 595898 198986 596134
rect 199222 595898 234986 596134
rect 235222 595898 270986 596134
rect 271222 595898 376982 596134
rect 377218 595898 414986 596134
rect 415222 595898 496982 596134
rect 497218 595898 522986 596134
rect 523222 595898 558986 596134
rect 559222 595898 586442 596134
rect 586678 595898 586860 596134
rect -2936 595876 586860 595898
rect -2936 595874 -2336 595876
rect 18804 595874 19404 595876
rect 54804 595874 55404 595876
rect 90804 595874 91404 595876
rect 126804 595874 127404 595876
rect 162804 595874 163404 595876
rect 198804 595874 199404 595876
rect 234804 595874 235404 595876
rect 270804 595874 271404 595876
rect 376938 595874 377262 595876
rect 414804 595874 415404 595876
rect 496938 595874 497262 595876
rect 522804 595874 523404 595876
rect 558804 595874 559404 595876
rect 586260 595874 586860 595876
rect -7636 589276 -7036 589278
rect 11604 589276 12204 589278
rect 47604 589276 48204 589278
rect 83604 589276 84204 589278
rect 119604 589276 120204 589278
rect 155604 589276 156204 589278
rect 191604 589276 192204 589278
rect 227604 589276 228204 589278
rect 263604 589276 264204 589278
rect 407604 589276 408204 589278
rect 515604 589276 516204 589278
rect 551604 589276 552204 589278
rect 590960 589276 591560 589278
rect -8576 589254 592500 589276
rect -8576 589018 -7454 589254
rect -7218 589018 11786 589254
rect 12022 589018 47786 589254
rect 48022 589018 83786 589254
rect 84022 589018 119786 589254
rect 120022 589018 155786 589254
rect 156022 589018 191786 589254
rect 192022 589018 227786 589254
rect 228022 589018 263786 589254
rect 264022 589018 407786 589254
rect 408022 589018 515786 589254
rect 516022 589018 551786 589254
rect 552022 589018 591142 589254
rect 591378 589018 592500 589254
rect -8576 588934 592500 589018
rect -8576 588698 -7454 588934
rect -7218 588698 11786 588934
rect 12022 588698 47786 588934
rect 48022 588698 83786 588934
rect 84022 588698 119786 588934
rect 120022 588698 155786 588934
rect 156022 588698 191786 588934
rect 192022 588698 227786 588934
rect 228022 588698 263786 588934
rect 264022 588698 407786 588934
rect 408022 588698 515786 588934
rect 516022 588698 551786 588934
rect 552022 588698 591142 588934
rect 591378 588698 592500 588934
rect -8576 588676 592500 588698
rect -7636 588674 -7036 588676
rect 11604 588674 12204 588676
rect 47604 588674 48204 588676
rect 83604 588674 84204 588676
rect 119604 588674 120204 588676
rect 155604 588674 156204 588676
rect 191604 588674 192204 588676
rect 227604 588674 228204 588676
rect 263604 588674 264204 588676
rect 407604 588674 408204 588676
rect 515604 588674 516204 588676
rect 551604 588674 552204 588676
rect 590960 588674 591560 588676
rect -5756 585676 -5156 585678
rect 8004 585676 8604 585678
rect 44004 585676 44604 585678
rect 80004 585676 80604 585678
rect 116004 585676 116604 585678
rect 152004 585676 152604 585678
rect 188004 585676 188604 585678
rect 224004 585676 224604 585678
rect 260004 585676 260604 585678
rect 296004 585676 296604 585678
rect 404004 585676 404604 585678
rect 512004 585676 512604 585678
rect 548004 585676 548604 585678
rect 589080 585676 589680 585678
rect -6696 585654 590620 585676
rect -6696 585418 -5574 585654
rect -5338 585418 8186 585654
rect 8422 585418 44186 585654
rect 44422 585418 80186 585654
rect 80422 585418 116186 585654
rect 116422 585418 152186 585654
rect 152422 585418 188186 585654
rect 188422 585418 224186 585654
rect 224422 585418 260186 585654
rect 260422 585418 296186 585654
rect 296422 585418 404186 585654
rect 404422 585418 512186 585654
rect 512422 585418 548186 585654
rect 548422 585418 589262 585654
rect 589498 585418 590620 585654
rect -6696 585334 590620 585418
rect -6696 585098 -5574 585334
rect -5338 585098 8186 585334
rect 8422 585098 44186 585334
rect 44422 585098 80186 585334
rect 80422 585098 116186 585334
rect 116422 585098 152186 585334
rect 152422 585098 188186 585334
rect 188422 585098 224186 585334
rect 224422 585098 260186 585334
rect 260422 585098 296186 585334
rect 296422 585098 404186 585334
rect 404422 585098 512186 585334
rect 512422 585098 548186 585334
rect 548422 585098 589262 585334
rect 589498 585098 590620 585334
rect -6696 585076 590620 585098
rect -5756 585074 -5156 585076
rect 8004 585074 8604 585076
rect 44004 585074 44604 585076
rect 80004 585074 80604 585076
rect 116004 585074 116604 585076
rect 152004 585074 152604 585076
rect 188004 585074 188604 585076
rect 224004 585074 224604 585076
rect 260004 585074 260604 585076
rect 296004 585074 296604 585076
rect 404004 585074 404604 585076
rect 512004 585074 512604 585076
rect 548004 585074 548604 585076
rect 589080 585074 589680 585076
rect -3876 582076 -3276 582078
rect 4404 582076 5004 582078
rect 40404 582076 41004 582078
rect 76404 582076 77004 582078
rect 112404 582076 113004 582078
rect 148404 582076 149004 582078
rect 184404 582076 185004 582078
rect 220404 582076 221004 582078
rect 256404 582076 257004 582078
rect 292404 582076 293004 582078
rect 400404 582076 401004 582078
rect 508404 582076 509004 582078
rect 544404 582076 545004 582078
rect 580404 582076 581004 582078
rect 587200 582076 587800 582078
rect -4816 582054 588740 582076
rect -4816 581818 -3694 582054
rect -3458 581818 4586 582054
rect 4822 581818 40586 582054
rect 40822 581818 76586 582054
rect 76822 581818 112586 582054
rect 112822 581818 148586 582054
rect 148822 581818 184586 582054
rect 184822 581818 220586 582054
rect 220822 581818 256586 582054
rect 256822 581818 292586 582054
rect 292822 581818 400586 582054
rect 400822 581818 508586 582054
rect 508822 581818 544586 582054
rect 544822 581818 580586 582054
rect 580822 581818 587382 582054
rect 587618 581818 588740 582054
rect -4816 581734 588740 581818
rect -4816 581498 -3694 581734
rect -3458 581498 4586 581734
rect 4822 581498 40586 581734
rect 40822 581498 76586 581734
rect 76822 581498 112586 581734
rect 112822 581498 148586 581734
rect 148822 581498 184586 581734
rect 184822 581498 220586 581734
rect 220822 581498 256586 581734
rect 256822 581498 292586 581734
rect 292822 581498 400586 581734
rect 400822 581498 508586 581734
rect 508822 581498 544586 581734
rect 544822 581498 580586 581734
rect 580822 581498 587382 581734
rect 587618 581498 588740 581734
rect -4816 581476 588740 581498
rect -3876 581474 -3276 581476
rect 4404 581474 5004 581476
rect 40404 581474 41004 581476
rect 76404 581474 77004 581476
rect 112404 581474 113004 581476
rect 148404 581474 149004 581476
rect 184404 581474 185004 581476
rect 220404 581474 221004 581476
rect 256404 581474 257004 581476
rect 292404 581474 293004 581476
rect 400404 581474 401004 581476
rect 508404 581474 509004 581476
rect 544404 581474 545004 581476
rect 580404 581474 581004 581476
rect 587200 581474 587800 581476
rect -1996 578476 -1396 578478
rect 804 578476 1404 578478
rect 36804 578476 37404 578478
rect 72804 578476 73404 578478
rect 108804 578476 109404 578478
rect 144804 578476 145404 578478
rect 180804 578476 181404 578478
rect 216804 578476 217404 578478
rect 252804 578476 253404 578478
rect 288804 578476 289404 578478
rect 376494 578476 376814 578478
rect 396804 578476 397404 578478
rect 496494 578476 496814 578478
rect 504804 578476 505404 578478
rect 540804 578476 541404 578478
rect 576804 578476 577404 578478
rect 585320 578476 585920 578478
rect -2936 578454 586860 578476
rect -2936 578218 -1814 578454
rect -1578 578218 986 578454
rect 1222 578218 36986 578454
rect 37222 578218 72986 578454
rect 73222 578218 108986 578454
rect 109222 578218 144986 578454
rect 145222 578218 180986 578454
rect 181222 578218 216986 578454
rect 217222 578218 252986 578454
rect 253222 578218 288986 578454
rect 289222 578218 376536 578454
rect 376772 578218 396986 578454
rect 397222 578218 496536 578454
rect 496772 578218 504986 578454
rect 505222 578218 540986 578454
rect 541222 578218 576986 578454
rect 577222 578218 585502 578454
rect 585738 578218 586860 578454
rect -2936 578134 586860 578218
rect -2936 577898 -1814 578134
rect -1578 577898 986 578134
rect 1222 577898 36986 578134
rect 37222 577898 72986 578134
rect 73222 577898 108986 578134
rect 109222 577898 144986 578134
rect 145222 577898 180986 578134
rect 181222 577898 216986 578134
rect 217222 577898 252986 578134
rect 253222 577898 288986 578134
rect 289222 577898 376536 578134
rect 376772 577898 396986 578134
rect 397222 577898 496536 578134
rect 496772 577898 504986 578134
rect 505222 577898 540986 578134
rect 541222 577898 576986 578134
rect 577222 577898 585502 578134
rect 585738 577898 586860 578134
rect -2936 577876 586860 577898
rect -1996 577874 -1396 577876
rect 804 577874 1404 577876
rect 36804 577874 37404 577876
rect 72804 577874 73404 577876
rect 108804 577874 109404 577876
rect 144804 577874 145404 577876
rect 180804 577874 181404 577876
rect 216804 577874 217404 577876
rect 252804 577874 253404 577876
rect 288804 577874 289404 577876
rect 376494 577874 376814 577876
rect 396804 577874 397404 577876
rect 496494 577874 496814 577876
rect 504804 577874 505404 577876
rect 540804 577874 541404 577876
rect 576804 577874 577404 577876
rect 585320 577874 585920 577876
rect -8576 571276 -7976 571278
rect 29604 571276 30204 571278
rect 65604 571276 66204 571278
rect 101604 571276 102204 571278
rect 137604 571276 138204 571278
rect 173604 571276 174204 571278
rect 209604 571276 210204 571278
rect 245604 571276 246204 571278
rect 281604 571276 282204 571278
rect 389604 571276 390204 571278
rect 533604 571276 534204 571278
rect 569604 571276 570204 571278
rect 591900 571276 592500 571278
rect -8576 571254 592500 571276
rect -8576 571018 -8394 571254
rect -8158 571018 29786 571254
rect 30022 571018 65786 571254
rect 66022 571018 101786 571254
rect 102022 571018 137786 571254
rect 138022 571018 173786 571254
rect 174022 571018 209786 571254
rect 210022 571018 245786 571254
rect 246022 571018 281786 571254
rect 282022 571018 389786 571254
rect 390022 571018 533786 571254
rect 534022 571018 569786 571254
rect 570022 571018 592082 571254
rect 592318 571018 592500 571254
rect -8576 570934 592500 571018
rect -8576 570698 -8394 570934
rect -8158 570698 29786 570934
rect 30022 570698 65786 570934
rect 66022 570698 101786 570934
rect 102022 570698 137786 570934
rect 138022 570698 173786 570934
rect 174022 570698 209786 570934
rect 210022 570698 245786 570934
rect 246022 570698 281786 570934
rect 282022 570698 389786 570934
rect 390022 570698 533786 570934
rect 534022 570698 569786 570934
rect 570022 570698 592082 570934
rect 592318 570698 592500 570934
rect -8576 570676 592500 570698
rect -8576 570674 -7976 570676
rect 29604 570674 30204 570676
rect 65604 570674 66204 570676
rect 101604 570674 102204 570676
rect 137604 570674 138204 570676
rect 173604 570674 174204 570676
rect 209604 570674 210204 570676
rect 245604 570674 246204 570676
rect 281604 570674 282204 570676
rect 389604 570674 390204 570676
rect 533604 570674 534204 570676
rect 569604 570674 570204 570676
rect 591900 570674 592500 570676
rect -6696 567676 -6096 567678
rect 26004 567676 26604 567678
rect 62004 567676 62604 567678
rect 98004 567676 98604 567678
rect 134004 567676 134604 567678
rect 170004 567676 170604 567678
rect 206004 567676 206604 567678
rect 242004 567676 242604 567678
rect 278004 567676 278604 567678
rect 386004 567676 386604 567678
rect 530004 567676 530604 567678
rect 566004 567676 566604 567678
rect 590020 567676 590620 567678
rect -6696 567654 590620 567676
rect -6696 567418 -6514 567654
rect -6278 567418 26186 567654
rect 26422 567418 62186 567654
rect 62422 567418 98186 567654
rect 98422 567418 134186 567654
rect 134422 567418 170186 567654
rect 170422 567418 206186 567654
rect 206422 567418 242186 567654
rect 242422 567418 278186 567654
rect 278422 567418 386186 567654
rect 386422 567418 530186 567654
rect 530422 567418 566186 567654
rect 566422 567418 590202 567654
rect 590438 567418 590620 567654
rect -6696 567334 590620 567418
rect -6696 567098 -6514 567334
rect -6278 567098 26186 567334
rect 26422 567098 62186 567334
rect 62422 567098 98186 567334
rect 98422 567098 134186 567334
rect 134422 567098 170186 567334
rect 170422 567098 206186 567334
rect 206422 567098 242186 567334
rect 242422 567098 278186 567334
rect 278422 567098 386186 567334
rect 386422 567098 530186 567334
rect 530422 567098 566186 567334
rect 566422 567098 590202 567334
rect 590438 567098 590620 567334
rect -6696 567076 590620 567098
rect -6696 567074 -6096 567076
rect 26004 567074 26604 567076
rect 62004 567074 62604 567076
rect 98004 567074 98604 567076
rect 134004 567074 134604 567076
rect 170004 567074 170604 567076
rect 206004 567074 206604 567076
rect 242004 567074 242604 567076
rect 278004 567074 278604 567076
rect 386004 567074 386604 567076
rect 530004 567074 530604 567076
rect 566004 567074 566604 567076
rect 590020 567074 590620 567076
rect -4816 564076 -4216 564078
rect 22404 564076 23004 564078
rect 58404 564076 59004 564078
rect 94404 564076 95004 564078
rect 130404 564076 131004 564078
rect 166404 564076 167004 564078
rect 202404 564076 203004 564078
rect 238404 564076 239004 564078
rect 274404 564076 275004 564078
rect 382404 564076 383004 564078
rect 526404 564076 527004 564078
rect 562404 564076 563004 564078
rect 588140 564076 588740 564078
rect -4816 564054 588740 564076
rect -4816 563818 -4634 564054
rect -4398 563818 22586 564054
rect 22822 563818 58586 564054
rect 58822 563818 94586 564054
rect 94822 563818 130586 564054
rect 130822 563818 166586 564054
rect 166822 563818 202586 564054
rect 202822 563818 238586 564054
rect 238822 563818 274586 564054
rect 274822 563818 382586 564054
rect 382822 563818 526586 564054
rect 526822 563818 562586 564054
rect 562822 563818 588322 564054
rect 588558 563818 588740 564054
rect -4816 563734 588740 563818
rect -4816 563498 -4634 563734
rect -4398 563498 22586 563734
rect 22822 563498 58586 563734
rect 58822 563498 94586 563734
rect 94822 563498 130586 563734
rect 130822 563498 166586 563734
rect 166822 563498 202586 563734
rect 202822 563498 238586 563734
rect 238822 563498 274586 563734
rect 274822 563498 382586 563734
rect 382822 563498 526586 563734
rect 526822 563498 562586 563734
rect 562822 563498 588322 563734
rect 588558 563498 588740 563734
rect -4816 563476 588740 563498
rect -4816 563474 -4216 563476
rect 22404 563474 23004 563476
rect 58404 563474 59004 563476
rect 94404 563474 95004 563476
rect 130404 563474 131004 563476
rect 166404 563474 167004 563476
rect 202404 563474 203004 563476
rect 238404 563474 239004 563476
rect 274404 563474 275004 563476
rect 382404 563474 383004 563476
rect 526404 563474 527004 563476
rect 562404 563474 563004 563476
rect 588140 563474 588740 563476
rect -2936 560476 -2336 560478
rect 18804 560476 19404 560478
rect 54804 560476 55404 560478
rect 90804 560476 91404 560478
rect 126804 560476 127404 560478
rect 162804 560476 163404 560478
rect 198804 560476 199404 560478
rect 234804 560476 235404 560478
rect 270804 560476 271404 560478
rect 376938 560476 377262 560478
rect 414804 560476 415404 560478
rect 496938 560476 497262 560478
rect 522804 560476 523404 560478
rect 558804 560476 559404 560478
rect 586260 560476 586860 560478
rect -2936 560454 586860 560476
rect -2936 560218 -2754 560454
rect -2518 560218 18986 560454
rect 19222 560218 54986 560454
rect 55222 560218 90986 560454
rect 91222 560218 126986 560454
rect 127222 560218 162986 560454
rect 163222 560218 198986 560454
rect 199222 560218 234986 560454
rect 235222 560218 270986 560454
rect 271222 560218 376982 560454
rect 377218 560218 414986 560454
rect 415222 560218 496982 560454
rect 497218 560218 522986 560454
rect 523222 560218 558986 560454
rect 559222 560218 586442 560454
rect 586678 560218 586860 560454
rect -2936 560134 586860 560218
rect -2936 559898 -2754 560134
rect -2518 559898 18986 560134
rect 19222 559898 54986 560134
rect 55222 559898 90986 560134
rect 91222 559898 126986 560134
rect 127222 559898 162986 560134
rect 163222 559898 198986 560134
rect 199222 559898 234986 560134
rect 235222 559898 270986 560134
rect 271222 559898 376982 560134
rect 377218 559898 414986 560134
rect 415222 559898 496982 560134
rect 497218 559898 522986 560134
rect 523222 559898 558986 560134
rect 559222 559898 586442 560134
rect 586678 559898 586860 560134
rect -2936 559876 586860 559898
rect -2936 559874 -2336 559876
rect 18804 559874 19404 559876
rect 54804 559874 55404 559876
rect 90804 559874 91404 559876
rect 126804 559874 127404 559876
rect 162804 559874 163404 559876
rect 198804 559874 199404 559876
rect 234804 559874 235404 559876
rect 270804 559874 271404 559876
rect 376938 559874 377262 559876
rect 414804 559874 415404 559876
rect 496938 559874 497262 559876
rect 522804 559874 523404 559876
rect 558804 559874 559404 559876
rect 586260 559874 586860 559876
rect -7636 553276 -7036 553278
rect 11604 553276 12204 553278
rect 47604 553276 48204 553278
rect 83604 553276 84204 553278
rect 119604 553276 120204 553278
rect 155604 553276 156204 553278
rect 191604 553276 192204 553278
rect 227604 553276 228204 553278
rect 263604 553276 264204 553278
rect 407604 553276 408204 553278
rect 515604 553276 516204 553278
rect 551604 553276 552204 553278
rect 590960 553276 591560 553278
rect -8576 553254 592500 553276
rect -8576 553018 -7454 553254
rect -7218 553018 11786 553254
rect 12022 553018 47786 553254
rect 48022 553018 83786 553254
rect 84022 553018 119786 553254
rect 120022 553018 155786 553254
rect 156022 553018 191786 553254
rect 192022 553018 227786 553254
rect 228022 553018 263786 553254
rect 264022 553018 407786 553254
rect 408022 553018 515786 553254
rect 516022 553018 551786 553254
rect 552022 553018 591142 553254
rect 591378 553018 592500 553254
rect -8576 552934 592500 553018
rect -8576 552698 -7454 552934
rect -7218 552698 11786 552934
rect 12022 552698 47786 552934
rect 48022 552698 83786 552934
rect 84022 552698 119786 552934
rect 120022 552698 155786 552934
rect 156022 552698 191786 552934
rect 192022 552698 227786 552934
rect 228022 552698 263786 552934
rect 264022 552698 407786 552934
rect 408022 552698 515786 552934
rect 516022 552698 551786 552934
rect 552022 552698 591142 552934
rect 591378 552698 592500 552934
rect -8576 552676 592500 552698
rect -7636 552674 -7036 552676
rect 11604 552674 12204 552676
rect 47604 552674 48204 552676
rect 83604 552674 84204 552676
rect 119604 552674 120204 552676
rect 155604 552674 156204 552676
rect 191604 552674 192204 552676
rect 227604 552674 228204 552676
rect 263604 552674 264204 552676
rect 407604 552674 408204 552676
rect 515604 552674 516204 552676
rect 551604 552674 552204 552676
rect 590960 552674 591560 552676
rect -5756 549676 -5156 549678
rect 8004 549676 8604 549678
rect 44004 549676 44604 549678
rect 80004 549676 80604 549678
rect 116004 549676 116604 549678
rect 152004 549676 152604 549678
rect 188004 549676 188604 549678
rect 224004 549676 224604 549678
rect 260004 549676 260604 549678
rect 296004 549676 296604 549678
rect 404004 549676 404604 549678
rect 512004 549676 512604 549678
rect 548004 549676 548604 549678
rect 589080 549676 589680 549678
rect -6696 549654 590620 549676
rect -6696 549418 -5574 549654
rect -5338 549418 8186 549654
rect 8422 549418 44186 549654
rect 44422 549418 80186 549654
rect 80422 549418 116186 549654
rect 116422 549418 152186 549654
rect 152422 549418 188186 549654
rect 188422 549418 224186 549654
rect 224422 549418 260186 549654
rect 260422 549418 296186 549654
rect 296422 549418 404186 549654
rect 404422 549418 512186 549654
rect 512422 549418 548186 549654
rect 548422 549418 589262 549654
rect 589498 549418 590620 549654
rect -6696 549334 590620 549418
rect -6696 549098 -5574 549334
rect -5338 549098 8186 549334
rect 8422 549098 44186 549334
rect 44422 549098 80186 549334
rect 80422 549098 116186 549334
rect 116422 549098 152186 549334
rect 152422 549098 188186 549334
rect 188422 549098 224186 549334
rect 224422 549098 260186 549334
rect 260422 549098 296186 549334
rect 296422 549098 404186 549334
rect 404422 549098 512186 549334
rect 512422 549098 548186 549334
rect 548422 549098 589262 549334
rect 589498 549098 590620 549334
rect -6696 549076 590620 549098
rect -5756 549074 -5156 549076
rect 8004 549074 8604 549076
rect 44004 549074 44604 549076
rect 80004 549074 80604 549076
rect 116004 549074 116604 549076
rect 152004 549074 152604 549076
rect 188004 549074 188604 549076
rect 224004 549074 224604 549076
rect 260004 549074 260604 549076
rect 296004 549074 296604 549076
rect 404004 549074 404604 549076
rect 512004 549074 512604 549076
rect 548004 549074 548604 549076
rect 589080 549074 589680 549076
rect -3876 546076 -3276 546078
rect 4404 546076 5004 546078
rect 40404 546076 41004 546078
rect 76404 546076 77004 546078
rect 112404 546076 113004 546078
rect 148404 546076 149004 546078
rect 184404 546076 185004 546078
rect 220404 546076 221004 546078
rect 256404 546076 257004 546078
rect 292404 546076 293004 546078
rect 400404 546076 401004 546078
rect 508404 546076 509004 546078
rect 544404 546076 545004 546078
rect 580404 546076 581004 546078
rect 587200 546076 587800 546078
rect -4816 546054 588740 546076
rect -4816 545818 -3694 546054
rect -3458 545818 4586 546054
rect 4822 545818 40586 546054
rect 40822 545818 76586 546054
rect 76822 545818 112586 546054
rect 112822 545818 148586 546054
rect 148822 545818 184586 546054
rect 184822 545818 220586 546054
rect 220822 545818 256586 546054
rect 256822 545818 292586 546054
rect 292822 545818 400586 546054
rect 400822 545818 508586 546054
rect 508822 545818 544586 546054
rect 544822 545818 580586 546054
rect 580822 545818 587382 546054
rect 587618 545818 588740 546054
rect -4816 545734 588740 545818
rect -4816 545498 -3694 545734
rect -3458 545498 4586 545734
rect 4822 545498 40586 545734
rect 40822 545498 76586 545734
rect 76822 545498 112586 545734
rect 112822 545498 148586 545734
rect 148822 545498 184586 545734
rect 184822 545498 220586 545734
rect 220822 545498 256586 545734
rect 256822 545498 292586 545734
rect 292822 545498 400586 545734
rect 400822 545498 508586 545734
rect 508822 545498 544586 545734
rect 544822 545498 580586 545734
rect 580822 545498 587382 545734
rect 587618 545498 588740 545734
rect -4816 545476 588740 545498
rect -3876 545474 -3276 545476
rect 4404 545474 5004 545476
rect 40404 545474 41004 545476
rect 76404 545474 77004 545476
rect 112404 545474 113004 545476
rect 148404 545474 149004 545476
rect 184404 545474 185004 545476
rect 220404 545474 221004 545476
rect 256404 545474 257004 545476
rect 292404 545474 293004 545476
rect 400404 545474 401004 545476
rect 508404 545474 509004 545476
rect 544404 545474 545004 545476
rect 580404 545474 581004 545476
rect 587200 545474 587800 545476
rect -1996 542476 -1396 542478
rect 804 542476 1404 542478
rect 36804 542476 37404 542478
rect 72804 542476 73404 542478
rect 108804 542476 109404 542478
rect 144804 542476 145404 542478
rect 180804 542476 181404 542478
rect 216804 542476 217404 542478
rect 252804 542476 253404 542478
rect 288804 542476 289404 542478
rect 376494 542476 376814 542478
rect 396804 542476 397404 542478
rect 496494 542476 496814 542478
rect 504804 542476 505404 542478
rect 540804 542476 541404 542478
rect 576804 542476 577404 542478
rect 585320 542476 585920 542478
rect -2936 542454 586860 542476
rect -2936 542218 -1814 542454
rect -1578 542218 986 542454
rect 1222 542218 36986 542454
rect 37222 542218 72986 542454
rect 73222 542218 108986 542454
rect 109222 542218 144986 542454
rect 145222 542218 180986 542454
rect 181222 542218 216986 542454
rect 217222 542218 252986 542454
rect 253222 542218 288986 542454
rect 289222 542218 376536 542454
rect 376772 542218 396986 542454
rect 397222 542218 496536 542454
rect 496772 542218 504986 542454
rect 505222 542218 540986 542454
rect 541222 542218 576986 542454
rect 577222 542218 585502 542454
rect 585738 542218 586860 542454
rect -2936 542134 586860 542218
rect -2936 541898 -1814 542134
rect -1578 541898 986 542134
rect 1222 541898 36986 542134
rect 37222 541898 72986 542134
rect 73222 541898 108986 542134
rect 109222 541898 144986 542134
rect 145222 541898 180986 542134
rect 181222 541898 216986 542134
rect 217222 541898 252986 542134
rect 253222 541898 288986 542134
rect 289222 541898 376536 542134
rect 376772 541898 396986 542134
rect 397222 541898 496536 542134
rect 496772 541898 504986 542134
rect 505222 541898 540986 542134
rect 541222 541898 576986 542134
rect 577222 541898 585502 542134
rect 585738 541898 586860 542134
rect -2936 541876 586860 541898
rect -1996 541874 -1396 541876
rect 804 541874 1404 541876
rect 36804 541874 37404 541876
rect 72804 541874 73404 541876
rect 108804 541874 109404 541876
rect 144804 541874 145404 541876
rect 180804 541874 181404 541876
rect 216804 541874 217404 541876
rect 252804 541874 253404 541876
rect 288804 541874 289404 541876
rect 376494 541874 376814 541876
rect 396804 541874 397404 541876
rect 496494 541874 496814 541876
rect 504804 541874 505404 541876
rect 540804 541874 541404 541876
rect 576804 541874 577404 541876
rect 585320 541874 585920 541876
rect -8576 535276 -7976 535278
rect 29604 535276 30204 535278
rect 65604 535276 66204 535278
rect 101604 535276 102204 535278
rect 137604 535276 138204 535278
rect 173604 535276 174204 535278
rect 209604 535276 210204 535278
rect 245604 535276 246204 535278
rect 281604 535276 282204 535278
rect 389604 535276 390204 535278
rect 533604 535276 534204 535278
rect 569604 535276 570204 535278
rect 591900 535276 592500 535278
rect -8576 535254 592500 535276
rect -8576 535018 -8394 535254
rect -8158 535018 29786 535254
rect 30022 535018 65786 535254
rect 66022 535018 101786 535254
rect 102022 535018 137786 535254
rect 138022 535018 173786 535254
rect 174022 535018 209786 535254
rect 210022 535018 245786 535254
rect 246022 535018 281786 535254
rect 282022 535018 389786 535254
rect 390022 535018 533786 535254
rect 534022 535018 569786 535254
rect 570022 535018 592082 535254
rect 592318 535018 592500 535254
rect -8576 534934 592500 535018
rect -8576 534698 -8394 534934
rect -8158 534698 29786 534934
rect 30022 534698 65786 534934
rect 66022 534698 101786 534934
rect 102022 534698 137786 534934
rect 138022 534698 173786 534934
rect 174022 534698 209786 534934
rect 210022 534698 245786 534934
rect 246022 534698 281786 534934
rect 282022 534698 389786 534934
rect 390022 534698 533786 534934
rect 534022 534698 569786 534934
rect 570022 534698 592082 534934
rect 592318 534698 592500 534934
rect -8576 534676 592500 534698
rect -8576 534674 -7976 534676
rect 29604 534674 30204 534676
rect 65604 534674 66204 534676
rect 101604 534674 102204 534676
rect 137604 534674 138204 534676
rect 173604 534674 174204 534676
rect 209604 534674 210204 534676
rect 245604 534674 246204 534676
rect 281604 534674 282204 534676
rect 389604 534674 390204 534676
rect 533604 534674 534204 534676
rect 569604 534674 570204 534676
rect 591900 534674 592500 534676
rect -6696 531676 -6096 531678
rect 26004 531676 26604 531678
rect 62004 531676 62604 531678
rect 98004 531676 98604 531678
rect 134004 531676 134604 531678
rect 170004 531676 170604 531678
rect 206004 531676 206604 531678
rect 242004 531676 242604 531678
rect 278004 531676 278604 531678
rect 386004 531676 386604 531678
rect 530004 531676 530604 531678
rect 566004 531676 566604 531678
rect 590020 531676 590620 531678
rect -6696 531654 590620 531676
rect -6696 531418 -6514 531654
rect -6278 531418 26186 531654
rect 26422 531418 62186 531654
rect 62422 531418 98186 531654
rect 98422 531418 134186 531654
rect 134422 531418 170186 531654
rect 170422 531418 206186 531654
rect 206422 531418 242186 531654
rect 242422 531418 278186 531654
rect 278422 531418 386186 531654
rect 386422 531418 530186 531654
rect 530422 531418 566186 531654
rect 566422 531418 590202 531654
rect 590438 531418 590620 531654
rect -6696 531334 590620 531418
rect -6696 531098 -6514 531334
rect -6278 531098 26186 531334
rect 26422 531098 62186 531334
rect 62422 531098 98186 531334
rect 98422 531098 134186 531334
rect 134422 531098 170186 531334
rect 170422 531098 206186 531334
rect 206422 531098 242186 531334
rect 242422 531098 278186 531334
rect 278422 531098 386186 531334
rect 386422 531098 530186 531334
rect 530422 531098 566186 531334
rect 566422 531098 590202 531334
rect 590438 531098 590620 531334
rect -6696 531076 590620 531098
rect -6696 531074 -6096 531076
rect 26004 531074 26604 531076
rect 62004 531074 62604 531076
rect 98004 531074 98604 531076
rect 134004 531074 134604 531076
rect 170004 531074 170604 531076
rect 206004 531074 206604 531076
rect 242004 531074 242604 531076
rect 278004 531074 278604 531076
rect 386004 531074 386604 531076
rect 530004 531074 530604 531076
rect 566004 531074 566604 531076
rect 590020 531074 590620 531076
rect -4816 528076 -4216 528078
rect 22404 528076 23004 528078
rect 58404 528076 59004 528078
rect 94404 528076 95004 528078
rect 130404 528076 131004 528078
rect 166404 528076 167004 528078
rect 202404 528076 203004 528078
rect 238404 528076 239004 528078
rect 274404 528076 275004 528078
rect 382404 528076 383004 528078
rect 526404 528076 527004 528078
rect 562404 528076 563004 528078
rect 588140 528076 588740 528078
rect -4816 528054 588740 528076
rect -4816 527818 -4634 528054
rect -4398 527818 22586 528054
rect 22822 527818 58586 528054
rect 58822 527818 94586 528054
rect 94822 527818 130586 528054
rect 130822 527818 166586 528054
rect 166822 527818 202586 528054
rect 202822 527818 238586 528054
rect 238822 527818 274586 528054
rect 274822 527818 382586 528054
rect 382822 527818 526586 528054
rect 526822 527818 562586 528054
rect 562822 527818 588322 528054
rect 588558 527818 588740 528054
rect -4816 527734 588740 527818
rect -4816 527498 -4634 527734
rect -4398 527498 22586 527734
rect 22822 527498 58586 527734
rect 58822 527498 94586 527734
rect 94822 527498 130586 527734
rect 130822 527498 166586 527734
rect 166822 527498 202586 527734
rect 202822 527498 238586 527734
rect 238822 527498 274586 527734
rect 274822 527498 382586 527734
rect 382822 527498 526586 527734
rect 526822 527498 562586 527734
rect 562822 527498 588322 527734
rect 588558 527498 588740 527734
rect -4816 527476 588740 527498
rect -4816 527474 -4216 527476
rect 22404 527474 23004 527476
rect 58404 527474 59004 527476
rect 94404 527474 95004 527476
rect 130404 527474 131004 527476
rect 166404 527474 167004 527476
rect 202404 527474 203004 527476
rect 238404 527474 239004 527476
rect 274404 527474 275004 527476
rect 382404 527474 383004 527476
rect 526404 527474 527004 527476
rect 562404 527474 563004 527476
rect 588140 527474 588740 527476
rect -2936 524476 -2336 524478
rect 18804 524476 19404 524478
rect 54804 524476 55404 524478
rect 90804 524476 91404 524478
rect 126804 524476 127404 524478
rect 162804 524476 163404 524478
rect 198804 524476 199404 524478
rect 234804 524476 235404 524478
rect 270804 524476 271404 524478
rect 376938 524476 377262 524478
rect 414804 524476 415404 524478
rect 496938 524476 497262 524478
rect 522804 524476 523404 524478
rect 558804 524476 559404 524478
rect 586260 524476 586860 524478
rect -2936 524454 586860 524476
rect -2936 524218 -2754 524454
rect -2518 524218 18986 524454
rect 19222 524218 54986 524454
rect 55222 524218 90986 524454
rect 91222 524218 126986 524454
rect 127222 524218 162986 524454
rect 163222 524218 198986 524454
rect 199222 524218 234986 524454
rect 235222 524218 270986 524454
rect 271222 524218 376982 524454
rect 377218 524218 414986 524454
rect 415222 524218 496982 524454
rect 497218 524218 522986 524454
rect 523222 524218 558986 524454
rect 559222 524218 586442 524454
rect 586678 524218 586860 524454
rect -2936 524134 586860 524218
rect -2936 523898 -2754 524134
rect -2518 523898 18986 524134
rect 19222 523898 54986 524134
rect 55222 523898 90986 524134
rect 91222 523898 126986 524134
rect 127222 523898 162986 524134
rect 163222 523898 198986 524134
rect 199222 523898 234986 524134
rect 235222 523898 270986 524134
rect 271222 523898 376982 524134
rect 377218 523898 414986 524134
rect 415222 523898 496982 524134
rect 497218 523898 522986 524134
rect 523222 523898 558986 524134
rect 559222 523898 586442 524134
rect 586678 523898 586860 524134
rect -2936 523876 586860 523898
rect -2936 523874 -2336 523876
rect 18804 523874 19404 523876
rect 54804 523874 55404 523876
rect 90804 523874 91404 523876
rect 126804 523874 127404 523876
rect 162804 523874 163404 523876
rect 198804 523874 199404 523876
rect 234804 523874 235404 523876
rect 270804 523874 271404 523876
rect 376938 523874 377262 523876
rect 414804 523874 415404 523876
rect 496938 523874 497262 523876
rect 522804 523874 523404 523876
rect 558804 523874 559404 523876
rect 586260 523874 586860 523876
rect -7636 517276 -7036 517278
rect 11604 517276 12204 517278
rect 47604 517276 48204 517278
rect 83604 517276 84204 517278
rect 119604 517276 120204 517278
rect 155604 517276 156204 517278
rect 191604 517276 192204 517278
rect 227604 517276 228204 517278
rect 263604 517276 264204 517278
rect 407604 517276 408204 517278
rect 515604 517276 516204 517278
rect 551604 517276 552204 517278
rect 590960 517276 591560 517278
rect -8576 517254 592500 517276
rect -8576 517018 -7454 517254
rect -7218 517018 11786 517254
rect 12022 517018 47786 517254
rect 48022 517018 83786 517254
rect 84022 517018 119786 517254
rect 120022 517018 155786 517254
rect 156022 517018 191786 517254
rect 192022 517018 227786 517254
rect 228022 517018 263786 517254
rect 264022 517018 407786 517254
rect 408022 517018 515786 517254
rect 516022 517018 551786 517254
rect 552022 517018 591142 517254
rect 591378 517018 592500 517254
rect -8576 516934 592500 517018
rect -8576 516698 -7454 516934
rect -7218 516698 11786 516934
rect 12022 516698 47786 516934
rect 48022 516698 83786 516934
rect 84022 516698 119786 516934
rect 120022 516698 155786 516934
rect 156022 516698 191786 516934
rect 192022 516698 227786 516934
rect 228022 516698 263786 516934
rect 264022 516698 407786 516934
rect 408022 516698 515786 516934
rect 516022 516698 551786 516934
rect 552022 516698 591142 516934
rect 591378 516698 592500 516934
rect -8576 516676 592500 516698
rect -7636 516674 -7036 516676
rect 11604 516674 12204 516676
rect 47604 516674 48204 516676
rect 83604 516674 84204 516676
rect 119604 516674 120204 516676
rect 155604 516674 156204 516676
rect 191604 516674 192204 516676
rect 227604 516674 228204 516676
rect 263604 516674 264204 516676
rect 407604 516674 408204 516676
rect 515604 516674 516204 516676
rect 551604 516674 552204 516676
rect 590960 516674 591560 516676
rect -5756 513676 -5156 513678
rect 8004 513676 8604 513678
rect 44004 513676 44604 513678
rect 80004 513676 80604 513678
rect 116004 513676 116604 513678
rect 152004 513676 152604 513678
rect 188004 513676 188604 513678
rect 224004 513676 224604 513678
rect 260004 513676 260604 513678
rect 296004 513676 296604 513678
rect 332004 513676 332604 513678
rect 368004 513676 368604 513678
rect 404004 513676 404604 513678
rect 440004 513676 440604 513678
rect 476004 513676 476604 513678
rect 512004 513676 512604 513678
rect 548004 513676 548604 513678
rect 589080 513676 589680 513678
rect -6696 513654 590620 513676
rect -6696 513418 -5574 513654
rect -5338 513418 8186 513654
rect 8422 513418 44186 513654
rect 44422 513418 80186 513654
rect 80422 513418 116186 513654
rect 116422 513418 152186 513654
rect 152422 513418 188186 513654
rect 188422 513418 224186 513654
rect 224422 513418 260186 513654
rect 260422 513418 296186 513654
rect 296422 513418 332186 513654
rect 332422 513418 368186 513654
rect 368422 513418 404186 513654
rect 404422 513418 440186 513654
rect 440422 513418 476186 513654
rect 476422 513418 512186 513654
rect 512422 513418 548186 513654
rect 548422 513418 589262 513654
rect 589498 513418 590620 513654
rect -6696 513334 590620 513418
rect -6696 513098 -5574 513334
rect -5338 513098 8186 513334
rect 8422 513098 44186 513334
rect 44422 513098 80186 513334
rect 80422 513098 116186 513334
rect 116422 513098 152186 513334
rect 152422 513098 188186 513334
rect 188422 513098 224186 513334
rect 224422 513098 260186 513334
rect 260422 513098 296186 513334
rect 296422 513098 332186 513334
rect 332422 513098 368186 513334
rect 368422 513098 404186 513334
rect 404422 513098 440186 513334
rect 440422 513098 476186 513334
rect 476422 513098 512186 513334
rect 512422 513098 548186 513334
rect 548422 513098 589262 513334
rect 589498 513098 590620 513334
rect -6696 513076 590620 513098
rect -5756 513074 -5156 513076
rect 8004 513074 8604 513076
rect 44004 513074 44604 513076
rect 80004 513074 80604 513076
rect 116004 513074 116604 513076
rect 152004 513074 152604 513076
rect 188004 513074 188604 513076
rect 224004 513074 224604 513076
rect 260004 513074 260604 513076
rect 296004 513074 296604 513076
rect 332004 513074 332604 513076
rect 368004 513074 368604 513076
rect 404004 513074 404604 513076
rect 440004 513074 440604 513076
rect 476004 513074 476604 513076
rect 512004 513074 512604 513076
rect 548004 513074 548604 513076
rect 589080 513074 589680 513076
rect -3876 510076 -3276 510078
rect 4404 510076 5004 510078
rect 40404 510076 41004 510078
rect 76404 510076 77004 510078
rect 112404 510076 113004 510078
rect 148404 510076 149004 510078
rect 184404 510076 185004 510078
rect 220404 510076 221004 510078
rect 256404 510076 257004 510078
rect 292404 510076 293004 510078
rect 328404 510076 329004 510078
rect 364404 510076 365004 510078
rect 400404 510076 401004 510078
rect 436404 510076 437004 510078
rect 472404 510076 473004 510078
rect 508404 510076 509004 510078
rect 544404 510076 545004 510078
rect 580404 510076 581004 510078
rect 587200 510076 587800 510078
rect -4816 510054 588740 510076
rect -4816 509818 -3694 510054
rect -3458 509818 4586 510054
rect 4822 509818 40586 510054
rect 40822 509818 76586 510054
rect 76822 509818 112586 510054
rect 112822 509818 148586 510054
rect 148822 509818 184586 510054
rect 184822 509818 220586 510054
rect 220822 509818 256586 510054
rect 256822 509818 292586 510054
rect 292822 509818 328586 510054
rect 328822 509818 364586 510054
rect 364822 509818 400586 510054
rect 400822 509818 436586 510054
rect 436822 509818 472586 510054
rect 472822 509818 508586 510054
rect 508822 509818 544586 510054
rect 544822 509818 580586 510054
rect 580822 509818 587382 510054
rect 587618 509818 588740 510054
rect -4816 509734 588740 509818
rect -4816 509498 -3694 509734
rect -3458 509498 4586 509734
rect 4822 509498 40586 509734
rect 40822 509498 76586 509734
rect 76822 509498 112586 509734
rect 112822 509498 148586 509734
rect 148822 509498 184586 509734
rect 184822 509498 220586 509734
rect 220822 509498 256586 509734
rect 256822 509498 292586 509734
rect 292822 509498 328586 509734
rect 328822 509498 364586 509734
rect 364822 509498 400586 509734
rect 400822 509498 436586 509734
rect 436822 509498 472586 509734
rect 472822 509498 508586 509734
rect 508822 509498 544586 509734
rect 544822 509498 580586 509734
rect 580822 509498 587382 509734
rect 587618 509498 588740 509734
rect -4816 509476 588740 509498
rect -3876 509474 -3276 509476
rect 4404 509474 5004 509476
rect 40404 509474 41004 509476
rect 76404 509474 77004 509476
rect 112404 509474 113004 509476
rect 148404 509474 149004 509476
rect 184404 509474 185004 509476
rect 220404 509474 221004 509476
rect 256404 509474 257004 509476
rect 292404 509474 293004 509476
rect 328404 509474 329004 509476
rect 364404 509474 365004 509476
rect 400404 509474 401004 509476
rect 436404 509474 437004 509476
rect 472404 509474 473004 509476
rect 508404 509474 509004 509476
rect 544404 509474 545004 509476
rect 580404 509474 581004 509476
rect 587200 509474 587800 509476
rect -1996 506476 -1396 506478
rect 804 506476 1404 506478
rect 36804 506476 37404 506478
rect 72804 506476 73404 506478
rect 108804 506476 109404 506478
rect 144804 506476 145404 506478
rect 180804 506476 181404 506478
rect 216804 506476 217404 506478
rect 252804 506476 253404 506478
rect 288804 506476 289404 506478
rect 324804 506476 325404 506478
rect 360804 506476 361404 506478
rect 396804 506476 397404 506478
rect 432804 506476 433404 506478
rect 468804 506476 469404 506478
rect 504804 506476 505404 506478
rect 540804 506476 541404 506478
rect 576804 506476 577404 506478
rect 585320 506476 585920 506478
rect -2936 506454 586860 506476
rect -2936 506218 -1814 506454
rect -1578 506218 986 506454
rect 1222 506218 36986 506454
rect 37222 506218 72986 506454
rect 73222 506218 108986 506454
rect 109222 506218 144986 506454
rect 145222 506218 180986 506454
rect 181222 506218 216986 506454
rect 217222 506218 252986 506454
rect 253222 506218 288986 506454
rect 289222 506218 324986 506454
rect 325222 506218 360986 506454
rect 361222 506218 396986 506454
rect 397222 506218 432986 506454
rect 433222 506218 468986 506454
rect 469222 506218 504986 506454
rect 505222 506218 540986 506454
rect 541222 506218 576986 506454
rect 577222 506218 585502 506454
rect 585738 506218 586860 506454
rect -2936 506134 586860 506218
rect -2936 505898 -1814 506134
rect -1578 505898 986 506134
rect 1222 505898 36986 506134
rect 37222 505898 72986 506134
rect 73222 505898 108986 506134
rect 109222 505898 144986 506134
rect 145222 505898 180986 506134
rect 181222 505898 216986 506134
rect 217222 505898 252986 506134
rect 253222 505898 288986 506134
rect 289222 505898 324986 506134
rect 325222 505898 360986 506134
rect 361222 505898 396986 506134
rect 397222 505898 432986 506134
rect 433222 505898 468986 506134
rect 469222 505898 504986 506134
rect 505222 505898 540986 506134
rect 541222 505898 576986 506134
rect 577222 505898 585502 506134
rect 585738 505898 586860 506134
rect -2936 505876 586860 505898
rect -1996 505874 -1396 505876
rect 804 505874 1404 505876
rect 36804 505874 37404 505876
rect 72804 505874 73404 505876
rect 108804 505874 109404 505876
rect 144804 505874 145404 505876
rect 180804 505874 181404 505876
rect 216804 505874 217404 505876
rect 252804 505874 253404 505876
rect 288804 505874 289404 505876
rect 324804 505874 325404 505876
rect 360804 505874 361404 505876
rect 396804 505874 397404 505876
rect 432804 505874 433404 505876
rect 468804 505874 469404 505876
rect 504804 505874 505404 505876
rect 540804 505874 541404 505876
rect 576804 505874 577404 505876
rect 585320 505874 585920 505876
rect -8576 499276 -7976 499278
rect 29604 499276 30204 499278
rect 65604 499276 66204 499278
rect 101604 499276 102204 499278
rect 137604 499276 138204 499278
rect 173604 499276 174204 499278
rect 209604 499276 210204 499278
rect 245604 499276 246204 499278
rect 281604 499276 282204 499278
rect 317604 499276 318204 499278
rect 353604 499276 354204 499278
rect 389604 499276 390204 499278
rect 425604 499276 426204 499278
rect 461604 499276 462204 499278
rect 497604 499276 498204 499278
rect 533604 499276 534204 499278
rect 569604 499276 570204 499278
rect 591900 499276 592500 499278
rect -8576 499254 592500 499276
rect -8576 499018 -8394 499254
rect -8158 499018 29786 499254
rect 30022 499018 65786 499254
rect 66022 499018 101786 499254
rect 102022 499018 137786 499254
rect 138022 499018 173786 499254
rect 174022 499018 209786 499254
rect 210022 499018 245786 499254
rect 246022 499018 281786 499254
rect 282022 499018 317786 499254
rect 318022 499018 353786 499254
rect 354022 499018 389786 499254
rect 390022 499018 425786 499254
rect 426022 499018 461786 499254
rect 462022 499018 497786 499254
rect 498022 499018 533786 499254
rect 534022 499018 569786 499254
rect 570022 499018 592082 499254
rect 592318 499018 592500 499254
rect -8576 498934 592500 499018
rect -8576 498698 -8394 498934
rect -8158 498698 29786 498934
rect 30022 498698 65786 498934
rect 66022 498698 101786 498934
rect 102022 498698 137786 498934
rect 138022 498698 173786 498934
rect 174022 498698 209786 498934
rect 210022 498698 245786 498934
rect 246022 498698 281786 498934
rect 282022 498698 317786 498934
rect 318022 498698 353786 498934
rect 354022 498698 389786 498934
rect 390022 498698 425786 498934
rect 426022 498698 461786 498934
rect 462022 498698 497786 498934
rect 498022 498698 533786 498934
rect 534022 498698 569786 498934
rect 570022 498698 592082 498934
rect 592318 498698 592500 498934
rect -8576 498676 592500 498698
rect -8576 498674 -7976 498676
rect 29604 498674 30204 498676
rect 65604 498674 66204 498676
rect 101604 498674 102204 498676
rect 137604 498674 138204 498676
rect 173604 498674 174204 498676
rect 209604 498674 210204 498676
rect 245604 498674 246204 498676
rect 281604 498674 282204 498676
rect 317604 498674 318204 498676
rect 353604 498674 354204 498676
rect 389604 498674 390204 498676
rect 425604 498674 426204 498676
rect 461604 498674 462204 498676
rect 497604 498674 498204 498676
rect 533604 498674 534204 498676
rect 569604 498674 570204 498676
rect 591900 498674 592500 498676
rect -6696 495676 -6096 495678
rect 26004 495676 26604 495678
rect 62004 495676 62604 495678
rect 98004 495676 98604 495678
rect 134004 495676 134604 495678
rect 170004 495676 170604 495678
rect 206004 495676 206604 495678
rect 242004 495676 242604 495678
rect 278004 495676 278604 495678
rect 314004 495676 314604 495678
rect 350004 495676 350604 495678
rect 386004 495676 386604 495678
rect 422004 495676 422604 495678
rect 458004 495676 458604 495678
rect 494004 495676 494604 495678
rect 530004 495676 530604 495678
rect 566004 495676 566604 495678
rect 590020 495676 590620 495678
rect -6696 495654 590620 495676
rect -6696 495418 -6514 495654
rect -6278 495418 26186 495654
rect 26422 495418 62186 495654
rect 62422 495418 98186 495654
rect 98422 495418 134186 495654
rect 134422 495418 170186 495654
rect 170422 495418 206186 495654
rect 206422 495418 242186 495654
rect 242422 495418 278186 495654
rect 278422 495418 314186 495654
rect 314422 495418 350186 495654
rect 350422 495418 386186 495654
rect 386422 495418 422186 495654
rect 422422 495418 458186 495654
rect 458422 495418 494186 495654
rect 494422 495418 530186 495654
rect 530422 495418 566186 495654
rect 566422 495418 590202 495654
rect 590438 495418 590620 495654
rect -6696 495334 590620 495418
rect -6696 495098 -6514 495334
rect -6278 495098 26186 495334
rect 26422 495098 62186 495334
rect 62422 495098 98186 495334
rect 98422 495098 134186 495334
rect 134422 495098 170186 495334
rect 170422 495098 206186 495334
rect 206422 495098 242186 495334
rect 242422 495098 278186 495334
rect 278422 495098 314186 495334
rect 314422 495098 350186 495334
rect 350422 495098 386186 495334
rect 386422 495098 422186 495334
rect 422422 495098 458186 495334
rect 458422 495098 494186 495334
rect 494422 495098 530186 495334
rect 530422 495098 566186 495334
rect 566422 495098 590202 495334
rect 590438 495098 590620 495334
rect -6696 495076 590620 495098
rect -6696 495074 -6096 495076
rect 26004 495074 26604 495076
rect 62004 495074 62604 495076
rect 98004 495074 98604 495076
rect 134004 495074 134604 495076
rect 170004 495074 170604 495076
rect 206004 495074 206604 495076
rect 242004 495074 242604 495076
rect 278004 495074 278604 495076
rect 314004 495074 314604 495076
rect 350004 495074 350604 495076
rect 386004 495074 386604 495076
rect 422004 495074 422604 495076
rect 458004 495074 458604 495076
rect 494004 495074 494604 495076
rect 530004 495074 530604 495076
rect 566004 495074 566604 495076
rect 590020 495074 590620 495076
rect -4816 492076 -4216 492078
rect 22404 492076 23004 492078
rect 58404 492076 59004 492078
rect 94404 492076 95004 492078
rect 130404 492076 131004 492078
rect 166404 492076 167004 492078
rect 202404 492076 203004 492078
rect 238404 492076 239004 492078
rect 274404 492076 275004 492078
rect 310404 492076 311004 492078
rect 346404 492076 347004 492078
rect 382404 492076 383004 492078
rect 418404 492076 419004 492078
rect 454404 492076 455004 492078
rect 490404 492076 491004 492078
rect 526404 492076 527004 492078
rect 562404 492076 563004 492078
rect 588140 492076 588740 492078
rect -4816 492054 588740 492076
rect -4816 491818 -4634 492054
rect -4398 491818 22586 492054
rect 22822 491818 58586 492054
rect 58822 491818 94586 492054
rect 94822 491818 130586 492054
rect 130822 491818 166586 492054
rect 166822 491818 202586 492054
rect 202822 491818 238586 492054
rect 238822 491818 274586 492054
rect 274822 491818 310586 492054
rect 310822 491818 346586 492054
rect 346822 491818 382586 492054
rect 382822 491818 418586 492054
rect 418822 491818 454586 492054
rect 454822 491818 490586 492054
rect 490822 491818 526586 492054
rect 526822 491818 562586 492054
rect 562822 491818 588322 492054
rect 588558 491818 588740 492054
rect -4816 491734 588740 491818
rect -4816 491498 -4634 491734
rect -4398 491498 22586 491734
rect 22822 491498 58586 491734
rect 58822 491498 94586 491734
rect 94822 491498 130586 491734
rect 130822 491498 166586 491734
rect 166822 491498 202586 491734
rect 202822 491498 238586 491734
rect 238822 491498 274586 491734
rect 274822 491498 310586 491734
rect 310822 491498 346586 491734
rect 346822 491498 382586 491734
rect 382822 491498 418586 491734
rect 418822 491498 454586 491734
rect 454822 491498 490586 491734
rect 490822 491498 526586 491734
rect 526822 491498 562586 491734
rect 562822 491498 588322 491734
rect 588558 491498 588740 491734
rect -4816 491476 588740 491498
rect -4816 491474 -4216 491476
rect 22404 491474 23004 491476
rect 58404 491474 59004 491476
rect 94404 491474 95004 491476
rect 130404 491474 131004 491476
rect 166404 491474 167004 491476
rect 202404 491474 203004 491476
rect 238404 491474 239004 491476
rect 274404 491474 275004 491476
rect 310404 491474 311004 491476
rect 346404 491474 347004 491476
rect 382404 491474 383004 491476
rect 418404 491474 419004 491476
rect 454404 491474 455004 491476
rect 490404 491474 491004 491476
rect 526404 491474 527004 491476
rect 562404 491474 563004 491476
rect 588140 491474 588740 491476
rect -2936 488476 -2336 488478
rect 18804 488476 19404 488478
rect 54804 488476 55404 488478
rect 90804 488476 91404 488478
rect 126804 488476 127404 488478
rect 162804 488476 163404 488478
rect 198804 488476 199404 488478
rect 234804 488476 235404 488478
rect 270804 488476 271404 488478
rect 306804 488476 307404 488478
rect 342804 488476 343404 488478
rect 378804 488476 379404 488478
rect 414804 488476 415404 488478
rect 450804 488476 451404 488478
rect 486804 488476 487404 488478
rect 522804 488476 523404 488478
rect 558804 488476 559404 488478
rect 586260 488476 586860 488478
rect -2936 488454 586860 488476
rect -2936 488218 -2754 488454
rect -2518 488218 18986 488454
rect 19222 488218 54986 488454
rect 55222 488218 90986 488454
rect 91222 488218 126986 488454
rect 127222 488218 162986 488454
rect 163222 488218 198986 488454
rect 199222 488218 234986 488454
rect 235222 488218 270986 488454
rect 271222 488218 306986 488454
rect 307222 488218 342986 488454
rect 343222 488218 378986 488454
rect 379222 488218 414986 488454
rect 415222 488218 450986 488454
rect 451222 488218 486986 488454
rect 487222 488218 522986 488454
rect 523222 488218 558986 488454
rect 559222 488218 586442 488454
rect 586678 488218 586860 488454
rect -2936 488134 586860 488218
rect -2936 487898 -2754 488134
rect -2518 487898 18986 488134
rect 19222 487898 54986 488134
rect 55222 487898 90986 488134
rect 91222 487898 126986 488134
rect 127222 487898 162986 488134
rect 163222 487898 198986 488134
rect 199222 487898 234986 488134
rect 235222 487898 270986 488134
rect 271222 487898 306986 488134
rect 307222 487898 342986 488134
rect 343222 487898 378986 488134
rect 379222 487898 414986 488134
rect 415222 487898 450986 488134
rect 451222 487898 486986 488134
rect 487222 487898 522986 488134
rect 523222 487898 558986 488134
rect 559222 487898 586442 488134
rect 586678 487898 586860 488134
rect -2936 487876 586860 487898
rect -2936 487874 -2336 487876
rect 18804 487874 19404 487876
rect 54804 487874 55404 487876
rect 90804 487874 91404 487876
rect 126804 487874 127404 487876
rect 162804 487874 163404 487876
rect 198804 487874 199404 487876
rect 234804 487874 235404 487876
rect 270804 487874 271404 487876
rect 306804 487874 307404 487876
rect 342804 487874 343404 487876
rect 378804 487874 379404 487876
rect 414804 487874 415404 487876
rect 450804 487874 451404 487876
rect 486804 487874 487404 487876
rect 522804 487874 523404 487876
rect 558804 487874 559404 487876
rect 586260 487874 586860 487876
rect -7636 481276 -7036 481278
rect 11604 481276 12204 481278
rect 47604 481276 48204 481278
rect 83604 481276 84204 481278
rect 119604 481276 120204 481278
rect 155604 481276 156204 481278
rect 191604 481276 192204 481278
rect 227604 481276 228204 481278
rect 551604 481276 552204 481278
rect 590960 481276 591560 481278
rect -8576 481254 592500 481276
rect -8576 481018 -7454 481254
rect -7218 481018 11786 481254
rect 12022 481018 47786 481254
rect 48022 481018 83786 481254
rect 84022 481018 119786 481254
rect 120022 481018 155786 481254
rect 156022 481018 191786 481254
rect 192022 481018 227786 481254
rect 228022 481018 551786 481254
rect 552022 481018 591142 481254
rect 591378 481018 592500 481254
rect -8576 480934 592500 481018
rect -8576 480698 -7454 480934
rect -7218 480698 11786 480934
rect 12022 480698 47786 480934
rect 48022 480698 83786 480934
rect 84022 480698 119786 480934
rect 120022 480698 155786 480934
rect 156022 480698 191786 480934
rect 192022 480698 227786 480934
rect 228022 480698 551786 480934
rect 552022 480698 591142 480934
rect 591378 480698 592500 480934
rect -8576 480676 592500 480698
rect -7636 480674 -7036 480676
rect 11604 480674 12204 480676
rect 47604 480674 48204 480676
rect 83604 480674 84204 480676
rect 119604 480674 120204 480676
rect 155604 480674 156204 480676
rect 191604 480674 192204 480676
rect 227604 480674 228204 480676
rect 551604 480674 552204 480676
rect 590960 480674 591560 480676
rect -5756 477676 -5156 477678
rect 8004 477676 8604 477678
rect 44004 477676 44604 477678
rect 80004 477676 80604 477678
rect 116004 477676 116604 477678
rect 152004 477676 152604 477678
rect 188004 477676 188604 477678
rect 224004 477676 224604 477678
rect 548004 477676 548604 477678
rect 589080 477676 589680 477678
rect -6696 477654 590620 477676
rect -6696 477418 -5574 477654
rect -5338 477418 8186 477654
rect 8422 477418 44186 477654
rect 44422 477418 80186 477654
rect 80422 477418 116186 477654
rect 116422 477418 152186 477654
rect 152422 477418 188186 477654
rect 188422 477418 224186 477654
rect 224422 477418 548186 477654
rect 548422 477418 589262 477654
rect 589498 477418 590620 477654
rect -6696 477334 590620 477418
rect -6696 477098 -5574 477334
rect -5338 477098 8186 477334
rect 8422 477098 44186 477334
rect 44422 477098 80186 477334
rect 80422 477098 116186 477334
rect 116422 477098 152186 477334
rect 152422 477098 188186 477334
rect 188422 477098 224186 477334
rect 224422 477098 548186 477334
rect 548422 477098 589262 477334
rect 589498 477098 590620 477334
rect -6696 477076 590620 477098
rect -5756 477074 -5156 477076
rect 8004 477074 8604 477076
rect 44004 477074 44604 477076
rect 80004 477074 80604 477076
rect 116004 477074 116604 477076
rect 152004 477074 152604 477076
rect 188004 477074 188604 477076
rect 224004 477074 224604 477076
rect 548004 477074 548604 477076
rect 589080 477074 589680 477076
rect -3876 474076 -3276 474078
rect 4404 474076 5004 474078
rect 40404 474076 41004 474078
rect 76404 474076 77004 474078
rect 112404 474076 113004 474078
rect 148404 474076 149004 474078
rect 184404 474076 185004 474078
rect 220404 474076 221004 474078
rect 544404 474076 545004 474078
rect 580404 474076 581004 474078
rect 587200 474076 587800 474078
rect -4816 474054 588740 474076
rect -4816 473818 -3694 474054
rect -3458 473818 4586 474054
rect 4822 473818 40586 474054
rect 40822 473818 76586 474054
rect 76822 473818 112586 474054
rect 112822 473818 148586 474054
rect 148822 473818 184586 474054
rect 184822 473818 220586 474054
rect 220822 473818 544586 474054
rect 544822 473818 580586 474054
rect 580822 473818 587382 474054
rect 587618 473818 588740 474054
rect -4816 473734 588740 473818
rect -4816 473498 -3694 473734
rect -3458 473498 4586 473734
rect 4822 473498 40586 473734
rect 40822 473498 76586 473734
rect 76822 473498 112586 473734
rect 112822 473498 148586 473734
rect 148822 473498 184586 473734
rect 184822 473498 220586 473734
rect 220822 473498 544586 473734
rect 544822 473498 580586 473734
rect 580822 473498 587382 473734
rect 587618 473498 588740 473734
rect -4816 473476 588740 473498
rect -3876 473474 -3276 473476
rect 4404 473474 5004 473476
rect 40404 473474 41004 473476
rect 76404 473474 77004 473476
rect 112404 473474 113004 473476
rect 148404 473474 149004 473476
rect 184404 473474 185004 473476
rect 220404 473474 221004 473476
rect 544404 473474 545004 473476
rect 580404 473474 581004 473476
rect 587200 473474 587800 473476
rect -1996 470476 -1396 470478
rect 804 470476 1404 470478
rect 36804 470476 37404 470478
rect 72804 470476 73404 470478
rect 108804 470476 109404 470478
rect 144804 470476 145404 470478
rect 180804 470476 181404 470478
rect 216804 470476 217404 470478
rect 252804 470476 253404 470478
rect 264208 470476 264528 470478
rect 576804 470476 577404 470478
rect 585320 470476 585920 470478
rect -2936 470454 586860 470476
rect -2936 470218 -1814 470454
rect -1578 470218 986 470454
rect 1222 470218 36986 470454
rect 37222 470218 72986 470454
rect 73222 470218 108986 470454
rect 109222 470218 144986 470454
rect 145222 470218 180986 470454
rect 181222 470218 216986 470454
rect 217222 470218 252986 470454
rect 253222 470218 264250 470454
rect 264486 470218 576986 470454
rect 577222 470218 585502 470454
rect 585738 470218 586860 470454
rect -2936 470134 586860 470218
rect -2936 469898 -1814 470134
rect -1578 469898 986 470134
rect 1222 469898 36986 470134
rect 37222 469898 72986 470134
rect 73222 469898 108986 470134
rect 109222 469898 144986 470134
rect 145222 469898 180986 470134
rect 181222 469898 216986 470134
rect 217222 469898 252986 470134
rect 253222 469898 264250 470134
rect 264486 469898 576986 470134
rect 577222 469898 585502 470134
rect 585738 469898 586860 470134
rect -2936 469876 586860 469898
rect -1996 469874 -1396 469876
rect 804 469874 1404 469876
rect 36804 469874 37404 469876
rect 72804 469874 73404 469876
rect 108804 469874 109404 469876
rect 144804 469874 145404 469876
rect 180804 469874 181404 469876
rect 216804 469874 217404 469876
rect 252804 469874 253404 469876
rect 264208 469874 264528 469876
rect 576804 469874 577404 469876
rect 585320 469874 585920 469876
rect -8576 463276 -7976 463278
rect 29604 463276 30204 463278
rect 65604 463276 66204 463278
rect 101604 463276 102204 463278
rect 137604 463276 138204 463278
rect 173604 463276 174204 463278
rect 209604 463276 210204 463278
rect 245604 463276 246204 463278
rect 569604 463276 570204 463278
rect 591900 463276 592500 463278
rect -8576 463254 592500 463276
rect -8576 463018 -8394 463254
rect -8158 463018 29786 463254
rect 30022 463018 65786 463254
rect 66022 463018 101786 463254
rect 102022 463018 137786 463254
rect 138022 463018 173786 463254
rect 174022 463018 209786 463254
rect 210022 463018 245786 463254
rect 246022 463018 569786 463254
rect 570022 463018 592082 463254
rect 592318 463018 592500 463254
rect -8576 462934 592500 463018
rect -8576 462698 -8394 462934
rect -8158 462698 29786 462934
rect 30022 462698 65786 462934
rect 66022 462698 101786 462934
rect 102022 462698 137786 462934
rect 138022 462698 173786 462934
rect 174022 462698 209786 462934
rect 210022 462698 245786 462934
rect 246022 462698 569786 462934
rect 570022 462698 592082 462934
rect 592318 462698 592500 462934
rect -8576 462676 592500 462698
rect -8576 462674 -7976 462676
rect 29604 462674 30204 462676
rect 65604 462674 66204 462676
rect 101604 462674 102204 462676
rect 137604 462674 138204 462676
rect 173604 462674 174204 462676
rect 209604 462674 210204 462676
rect 245604 462674 246204 462676
rect 569604 462674 570204 462676
rect 591900 462674 592500 462676
rect -6696 459676 -6096 459678
rect 26004 459676 26604 459678
rect 62004 459676 62604 459678
rect 98004 459676 98604 459678
rect 134004 459676 134604 459678
rect 170004 459676 170604 459678
rect 206004 459676 206604 459678
rect 242004 459676 242604 459678
rect 566004 459676 566604 459678
rect 590020 459676 590620 459678
rect -6696 459654 590620 459676
rect -6696 459418 -6514 459654
rect -6278 459418 26186 459654
rect 26422 459418 62186 459654
rect 62422 459418 98186 459654
rect 98422 459418 134186 459654
rect 134422 459418 170186 459654
rect 170422 459418 206186 459654
rect 206422 459418 242186 459654
rect 242422 459418 566186 459654
rect 566422 459418 590202 459654
rect 590438 459418 590620 459654
rect -6696 459334 590620 459418
rect -6696 459098 -6514 459334
rect -6278 459098 26186 459334
rect 26422 459098 62186 459334
rect 62422 459098 98186 459334
rect 98422 459098 134186 459334
rect 134422 459098 170186 459334
rect 170422 459098 206186 459334
rect 206422 459098 242186 459334
rect 242422 459098 566186 459334
rect 566422 459098 590202 459334
rect 590438 459098 590620 459334
rect -6696 459076 590620 459098
rect -6696 459074 -6096 459076
rect 26004 459074 26604 459076
rect 62004 459074 62604 459076
rect 98004 459074 98604 459076
rect 134004 459074 134604 459076
rect 170004 459074 170604 459076
rect 206004 459074 206604 459076
rect 242004 459074 242604 459076
rect 566004 459074 566604 459076
rect 590020 459074 590620 459076
rect -4816 456076 -4216 456078
rect 22404 456076 23004 456078
rect 58404 456076 59004 456078
rect 94404 456076 95004 456078
rect 130404 456076 131004 456078
rect 166404 456076 167004 456078
rect 202404 456076 203004 456078
rect 238404 456076 239004 456078
rect 562404 456076 563004 456078
rect 588140 456076 588740 456078
rect -4816 456054 588740 456076
rect -4816 455818 -4634 456054
rect -4398 455818 22586 456054
rect 22822 455818 58586 456054
rect 58822 455818 94586 456054
rect 94822 455818 130586 456054
rect 130822 455818 166586 456054
rect 166822 455818 202586 456054
rect 202822 455818 238586 456054
rect 238822 455818 562586 456054
rect 562822 455818 588322 456054
rect 588558 455818 588740 456054
rect -4816 455734 588740 455818
rect -4816 455498 -4634 455734
rect -4398 455498 22586 455734
rect 22822 455498 58586 455734
rect 58822 455498 94586 455734
rect 94822 455498 130586 455734
rect 130822 455498 166586 455734
rect 166822 455498 202586 455734
rect 202822 455498 238586 455734
rect 238822 455498 562586 455734
rect 562822 455498 588322 455734
rect 588558 455498 588740 455734
rect -4816 455476 588740 455498
rect -4816 455474 -4216 455476
rect 22404 455474 23004 455476
rect 58404 455474 59004 455476
rect 94404 455474 95004 455476
rect 130404 455474 131004 455476
rect 166404 455474 167004 455476
rect 202404 455474 203004 455476
rect 238404 455474 239004 455476
rect 562404 455474 563004 455476
rect 588140 455474 588740 455476
rect -2936 452476 -2336 452478
rect 18804 452476 19404 452478
rect 54804 452476 55404 452478
rect 90804 452476 91404 452478
rect 126804 452476 127404 452478
rect 162804 452476 163404 452478
rect 198804 452476 199404 452478
rect 234804 452476 235404 452478
rect 279568 452476 279888 452478
rect 558804 452476 559404 452478
rect 586260 452476 586860 452478
rect -2936 452454 586860 452476
rect -2936 452218 -2754 452454
rect -2518 452218 18986 452454
rect 19222 452218 54986 452454
rect 55222 452218 90986 452454
rect 91222 452218 126986 452454
rect 127222 452218 162986 452454
rect 163222 452218 198986 452454
rect 199222 452218 234986 452454
rect 235222 452218 279610 452454
rect 279846 452218 558986 452454
rect 559222 452218 586442 452454
rect 586678 452218 586860 452454
rect -2936 452134 586860 452218
rect -2936 451898 -2754 452134
rect -2518 451898 18986 452134
rect 19222 451898 54986 452134
rect 55222 451898 90986 452134
rect 91222 451898 126986 452134
rect 127222 451898 162986 452134
rect 163222 451898 198986 452134
rect 199222 451898 234986 452134
rect 235222 451898 279610 452134
rect 279846 451898 558986 452134
rect 559222 451898 586442 452134
rect 586678 451898 586860 452134
rect -2936 451876 586860 451898
rect -2936 451874 -2336 451876
rect 18804 451874 19404 451876
rect 54804 451874 55404 451876
rect 90804 451874 91404 451876
rect 126804 451874 127404 451876
rect 162804 451874 163404 451876
rect 198804 451874 199404 451876
rect 234804 451874 235404 451876
rect 279568 451874 279888 451876
rect 558804 451874 559404 451876
rect 586260 451874 586860 451876
rect -7636 445276 -7036 445278
rect 11604 445276 12204 445278
rect 47604 445276 48204 445278
rect 83604 445276 84204 445278
rect 119604 445276 120204 445278
rect 155604 445276 156204 445278
rect 191604 445276 192204 445278
rect 227604 445276 228204 445278
rect 551604 445276 552204 445278
rect 590960 445276 591560 445278
rect -8576 445254 592500 445276
rect -8576 445018 -7454 445254
rect -7218 445018 11786 445254
rect 12022 445018 47786 445254
rect 48022 445018 83786 445254
rect 84022 445018 119786 445254
rect 120022 445018 155786 445254
rect 156022 445018 191786 445254
rect 192022 445018 227786 445254
rect 228022 445018 551786 445254
rect 552022 445018 591142 445254
rect 591378 445018 592500 445254
rect -8576 444934 592500 445018
rect -8576 444698 -7454 444934
rect -7218 444698 11786 444934
rect 12022 444698 47786 444934
rect 48022 444698 83786 444934
rect 84022 444698 119786 444934
rect 120022 444698 155786 444934
rect 156022 444698 191786 444934
rect 192022 444698 227786 444934
rect 228022 444698 551786 444934
rect 552022 444698 591142 444934
rect 591378 444698 592500 444934
rect -8576 444676 592500 444698
rect -7636 444674 -7036 444676
rect 11604 444674 12204 444676
rect 47604 444674 48204 444676
rect 83604 444674 84204 444676
rect 119604 444674 120204 444676
rect 155604 444674 156204 444676
rect 191604 444674 192204 444676
rect 227604 444674 228204 444676
rect 551604 444674 552204 444676
rect 590960 444674 591560 444676
rect -5756 441676 -5156 441678
rect 8004 441676 8604 441678
rect 44004 441676 44604 441678
rect 80004 441676 80604 441678
rect 116004 441676 116604 441678
rect 152004 441676 152604 441678
rect 188004 441676 188604 441678
rect 224004 441676 224604 441678
rect 548004 441676 548604 441678
rect 589080 441676 589680 441678
rect -6696 441654 590620 441676
rect -6696 441418 -5574 441654
rect -5338 441418 8186 441654
rect 8422 441418 44186 441654
rect 44422 441418 80186 441654
rect 80422 441418 116186 441654
rect 116422 441418 152186 441654
rect 152422 441418 188186 441654
rect 188422 441418 224186 441654
rect 224422 441418 548186 441654
rect 548422 441418 589262 441654
rect 589498 441418 590620 441654
rect -6696 441334 590620 441418
rect -6696 441098 -5574 441334
rect -5338 441098 8186 441334
rect 8422 441098 44186 441334
rect 44422 441098 80186 441334
rect 80422 441098 116186 441334
rect 116422 441098 152186 441334
rect 152422 441098 188186 441334
rect 188422 441098 224186 441334
rect 224422 441098 548186 441334
rect 548422 441098 589262 441334
rect 589498 441098 590620 441334
rect -6696 441076 590620 441098
rect -5756 441074 -5156 441076
rect 8004 441074 8604 441076
rect 44004 441074 44604 441076
rect 80004 441074 80604 441076
rect 116004 441074 116604 441076
rect 152004 441074 152604 441076
rect 188004 441074 188604 441076
rect 224004 441074 224604 441076
rect 548004 441074 548604 441076
rect 589080 441074 589680 441076
rect -3876 438076 -3276 438078
rect 4404 438076 5004 438078
rect 40404 438076 41004 438078
rect 76404 438076 77004 438078
rect 112404 438076 113004 438078
rect 148404 438076 149004 438078
rect 184404 438076 185004 438078
rect 220404 438076 221004 438078
rect 544404 438076 545004 438078
rect 580404 438076 581004 438078
rect 587200 438076 587800 438078
rect -4816 438054 588740 438076
rect -4816 437818 -3694 438054
rect -3458 437818 4586 438054
rect 4822 437818 40586 438054
rect 40822 437818 76586 438054
rect 76822 437818 112586 438054
rect 112822 437818 148586 438054
rect 148822 437818 184586 438054
rect 184822 437818 220586 438054
rect 220822 437818 544586 438054
rect 544822 437818 580586 438054
rect 580822 437818 587382 438054
rect 587618 437818 588740 438054
rect -4816 437734 588740 437818
rect -4816 437498 -3694 437734
rect -3458 437498 4586 437734
rect 4822 437498 40586 437734
rect 40822 437498 76586 437734
rect 76822 437498 112586 437734
rect 112822 437498 148586 437734
rect 148822 437498 184586 437734
rect 184822 437498 220586 437734
rect 220822 437498 544586 437734
rect 544822 437498 580586 437734
rect 580822 437498 587382 437734
rect 587618 437498 588740 437734
rect -4816 437476 588740 437498
rect -3876 437474 -3276 437476
rect 4404 437474 5004 437476
rect 40404 437474 41004 437476
rect 76404 437474 77004 437476
rect 112404 437474 113004 437476
rect 148404 437474 149004 437476
rect 184404 437474 185004 437476
rect 220404 437474 221004 437476
rect 544404 437474 545004 437476
rect 580404 437474 581004 437476
rect 587200 437474 587800 437476
rect -1996 434476 -1396 434478
rect 804 434476 1404 434478
rect 36804 434476 37404 434478
rect 72804 434476 73404 434478
rect 108804 434476 109404 434478
rect 144804 434476 145404 434478
rect 180804 434476 181404 434478
rect 216804 434476 217404 434478
rect 252804 434476 253404 434478
rect 264208 434476 264528 434478
rect 576804 434476 577404 434478
rect 585320 434476 585920 434478
rect -2936 434454 586860 434476
rect -2936 434218 -1814 434454
rect -1578 434218 986 434454
rect 1222 434218 36986 434454
rect 37222 434218 72986 434454
rect 73222 434218 108986 434454
rect 109222 434218 144986 434454
rect 145222 434218 180986 434454
rect 181222 434218 216986 434454
rect 217222 434218 252986 434454
rect 253222 434218 264250 434454
rect 264486 434218 576986 434454
rect 577222 434218 585502 434454
rect 585738 434218 586860 434454
rect -2936 434134 586860 434218
rect -2936 433898 -1814 434134
rect -1578 433898 986 434134
rect 1222 433898 36986 434134
rect 37222 433898 72986 434134
rect 73222 433898 108986 434134
rect 109222 433898 144986 434134
rect 145222 433898 180986 434134
rect 181222 433898 216986 434134
rect 217222 433898 252986 434134
rect 253222 433898 264250 434134
rect 264486 433898 576986 434134
rect 577222 433898 585502 434134
rect 585738 433898 586860 434134
rect -2936 433876 586860 433898
rect -1996 433874 -1396 433876
rect 804 433874 1404 433876
rect 36804 433874 37404 433876
rect 72804 433874 73404 433876
rect 108804 433874 109404 433876
rect 144804 433874 145404 433876
rect 180804 433874 181404 433876
rect 216804 433874 217404 433876
rect 252804 433874 253404 433876
rect 264208 433874 264528 433876
rect 576804 433874 577404 433876
rect 585320 433874 585920 433876
rect -8576 427276 -7976 427278
rect 29604 427276 30204 427278
rect 65604 427276 66204 427278
rect 101604 427276 102204 427278
rect 137604 427276 138204 427278
rect 173604 427276 174204 427278
rect 209604 427276 210204 427278
rect 245604 427276 246204 427278
rect 569604 427276 570204 427278
rect 591900 427276 592500 427278
rect -8576 427254 592500 427276
rect -8576 427018 -8394 427254
rect -8158 427018 29786 427254
rect 30022 427018 65786 427254
rect 66022 427018 101786 427254
rect 102022 427018 137786 427254
rect 138022 427018 173786 427254
rect 174022 427018 209786 427254
rect 210022 427018 245786 427254
rect 246022 427018 569786 427254
rect 570022 427018 592082 427254
rect 592318 427018 592500 427254
rect -8576 426934 592500 427018
rect -8576 426698 -8394 426934
rect -8158 426698 29786 426934
rect 30022 426698 65786 426934
rect 66022 426698 101786 426934
rect 102022 426698 137786 426934
rect 138022 426698 173786 426934
rect 174022 426698 209786 426934
rect 210022 426698 245786 426934
rect 246022 426698 569786 426934
rect 570022 426698 592082 426934
rect 592318 426698 592500 426934
rect -8576 426676 592500 426698
rect -8576 426674 -7976 426676
rect 29604 426674 30204 426676
rect 65604 426674 66204 426676
rect 101604 426674 102204 426676
rect 137604 426674 138204 426676
rect 173604 426674 174204 426676
rect 209604 426674 210204 426676
rect 245604 426674 246204 426676
rect 569604 426674 570204 426676
rect 591900 426674 592500 426676
rect -6696 423676 -6096 423678
rect 26004 423676 26604 423678
rect 62004 423676 62604 423678
rect 98004 423676 98604 423678
rect 134004 423676 134604 423678
rect 170004 423676 170604 423678
rect 206004 423676 206604 423678
rect 242004 423676 242604 423678
rect 566004 423676 566604 423678
rect 590020 423676 590620 423678
rect -6696 423654 590620 423676
rect -6696 423418 -6514 423654
rect -6278 423418 26186 423654
rect 26422 423418 62186 423654
rect 62422 423418 98186 423654
rect 98422 423418 134186 423654
rect 134422 423418 170186 423654
rect 170422 423418 206186 423654
rect 206422 423418 242186 423654
rect 242422 423418 566186 423654
rect 566422 423418 590202 423654
rect 590438 423418 590620 423654
rect -6696 423334 590620 423418
rect -6696 423098 -6514 423334
rect -6278 423098 26186 423334
rect 26422 423098 62186 423334
rect 62422 423098 98186 423334
rect 98422 423098 134186 423334
rect 134422 423098 170186 423334
rect 170422 423098 206186 423334
rect 206422 423098 242186 423334
rect 242422 423098 566186 423334
rect 566422 423098 590202 423334
rect 590438 423098 590620 423334
rect -6696 423076 590620 423098
rect -6696 423074 -6096 423076
rect 26004 423074 26604 423076
rect 62004 423074 62604 423076
rect 98004 423074 98604 423076
rect 134004 423074 134604 423076
rect 170004 423074 170604 423076
rect 206004 423074 206604 423076
rect 242004 423074 242604 423076
rect 566004 423074 566604 423076
rect 590020 423074 590620 423076
rect -4816 420076 -4216 420078
rect 22404 420076 23004 420078
rect 58404 420076 59004 420078
rect 94404 420076 95004 420078
rect 130404 420076 131004 420078
rect 166404 420076 167004 420078
rect 202404 420076 203004 420078
rect 238404 420076 239004 420078
rect 562404 420076 563004 420078
rect 588140 420076 588740 420078
rect -4816 420054 588740 420076
rect -4816 419818 -4634 420054
rect -4398 419818 22586 420054
rect 22822 419818 58586 420054
rect 58822 419818 94586 420054
rect 94822 419818 130586 420054
rect 130822 419818 166586 420054
rect 166822 419818 202586 420054
rect 202822 419818 238586 420054
rect 238822 419818 562586 420054
rect 562822 419818 588322 420054
rect 588558 419818 588740 420054
rect -4816 419734 588740 419818
rect -4816 419498 -4634 419734
rect -4398 419498 22586 419734
rect 22822 419498 58586 419734
rect 58822 419498 94586 419734
rect 94822 419498 130586 419734
rect 130822 419498 166586 419734
rect 166822 419498 202586 419734
rect 202822 419498 238586 419734
rect 238822 419498 562586 419734
rect 562822 419498 588322 419734
rect 588558 419498 588740 419734
rect -4816 419476 588740 419498
rect -4816 419474 -4216 419476
rect 22404 419474 23004 419476
rect 58404 419474 59004 419476
rect 94404 419474 95004 419476
rect 130404 419474 131004 419476
rect 166404 419474 167004 419476
rect 202404 419474 203004 419476
rect 238404 419474 239004 419476
rect 562404 419474 563004 419476
rect 588140 419474 588740 419476
rect -2936 416476 -2336 416478
rect 18804 416476 19404 416478
rect 54804 416476 55404 416478
rect 90804 416476 91404 416478
rect 126804 416476 127404 416478
rect 162804 416476 163404 416478
rect 198804 416476 199404 416478
rect 234804 416476 235404 416478
rect 279568 416476 279888 416478
rect 558804 416476 559404 416478
rect 586260 416476 586860 416478
rect -2936 416454 586860 416476
rect -2936 416218 -2754 416454
rect -2518 416218 18986 416454
rect 19222 416218 54986 416454
rect 55222 416218 90986 416454
rect 91222 416218 126986 416454
rect 127222 416218 162986 416454
rect 163222 416218 198986 416454
rect 199222 416218 234986 416454
rect 235222 416218 279610 416454
rect 279846 416218 558986 416454
rect 559222 416218 586442 416454
rect 586678 416218 586860 416454
rect -2936 416134 586860 416218
rect -2936 415898 -2754 416134
rect -2518 415898 18986 416134
rect 19222 415898 54986 416134
rect 55222 415898 90986 416134
rect 91222 415898 126986 416134
rect 127222 415898 162986 416134
rect 163222 415898 198986 416134
rect 199222 415898 234986 416134
rect 235222 415898 279610 416134
rect 279846 415898 558986 416134
rect 559222 415898 586442 416134
rect 586678 415898 586860 416134
rect -2936 415876 586860 415898
rect -2936 415874 -2336 415876
rect 18804 415874 19404 415876
rect 54804 415874 55404 415876
rect 90804 415874 91404 415876
rect 126804 415874 127404 415876
rect 162804 415874 163404 415876
rect 198804 415874 199404 415876
rect 234804 415874 235404 415876
rect 279568 415874 279888 415876
rect 558804 415874 559404 415876
rect 586260 415874 586860 415876
rect -7636 409276 -7036 409278
rect 11604 409276 12204 409278
rect 47604 409276 48204 409278
rect 83604 409276 84204 409278
rect 119604 409276 120204 409278
rect 155604 409276 156204 409278
rect 191604 409276 192204 409278
rect 227604 409276 228204 409278
rect 551604 409276 552204 409278
rect 590960 409276 591560 409278
rect -8576 409254 592500 409276
rect -8576 409018 -7454 409254
rect -7218 409018 11786 409254
rect 12022 409018 47786 409254
rect 48022 409018 83786 409254
rect 84022 409018 119786 409254
rect 120022 409018 155786 409254
rect 156022 409018 191786 409254
rect 192022 409018 227786 409254
rect 228022 409018 551786 409254
rect 552022 409018 591142 409254
rect 591378 409018 592500 409254
rect -8576 408934 592500 409018
rect -8576 408698 -7454 408934
rect -7218 408698 11786 408934
rect 12022 408698 47786 408934
rect 48022 408698 83786 408934
rect 84022 408698 119786 408934
rect 120022 408698 155786 408934
rect 156022 408698 191786 408934
rect 192022 408698 227786 408934
rect 228022 408698 551786 408934
rect 552022 408698 591142 408934
rect 591378 408698 592500 408934
rect -8576 408676 592500 408698
rect -7636 408674 -7036 408676
rect 11604 408674 12204 408676
rect 47604 408674 48204 408676
rect 83604 408674 84204 408676
rect 119604 408674 120204 408676
rect 155604 408674 156204 408676
rect 191604 408674 192204 408676
rect 227604 408674 228204 408676
rect 551604 408674 552204 408676
rect 590960 408674 591560 408676
rect -5756 405676 -5156 405678
rect 8004 405676 8604 405678
rect 44004 405676 44604 405678
rect 80004 405676 80604 405678
rect 116004 405676 116604 405678
rect 152004 405676 152604 405678
rect 188004 405676 188604 405678
rect 224004 405676 224604 405678
rect 548004 405676 548604 405678
rect 589080 405676 589680 405678
rect -6696 405654 590620 405676
rect -6696 405418 -5574 405654
rect -5338 405418 8186 405654
rect 8422 405418 44186 405654
rect 44422 405418 80186 405654
rect 80422 405418 116186 405654
rect 116422 405418 152186 405654
rect 152422 405418 188186 405654
rect 188422 405418 224186 405654
rect 224422 405418 548186 405654
rect 548422 405418 589262 405654
rect 589498 405418 590620 405654
rect -6696 405334 590620 405418
rect -6696 405098 -5574 405334
rect -5338 405098 8186 405334
rect 8422 405098 44186 405334
rect 44422 405098 80186 405334
rect 80422 405098 116186 405334
rect 116422 405098 152186 405334
rect 152422 405098 188186 405334
rect 188422 405098 224186 405334
rect 224422 405098 548186 405334
rect 548422 405098 589262 405334
rect 589498 405098 590620 405334
rect -6696 405076 590620 405098
rect -5756 405074 -5156 405076
rect 8004 405074 8604 405076
rect 44004 405074 44604 405076
rect 80004 405074 80604 405076
rect 116004 405074 116604 405076
rect 152004 405074 152604 405076
rect 188004 405074 188604 405076
rect 224004 405074 224604 405076
rect 548004 405074 548604 405076
rect 589080 405074 589680 405076
rect -3876 402076 -3276 402078
rect 4404 402076 5004 402078
rect 40404 402076 41004 402078
rect 76404 402076 77004 402078
rect 112404 402076 113004 402078
rect 148404 402076 149004 402078
rect 184404 402076 185004 402078
rect 220404 402076 221004 402078
rect 544404 402076 545004 402078
rect 580404 402076 581004 402078
rect 587200 402076 587800 402078
rect -4816 402054 588740 402076
rect -4816 401818 -3694 402054
rect -3458 401818 4586 402054
rect 4822 401818 40586 402054
rect 40822 401818 76586 402054
rect 76822 401818 112586 402054
rect 112822 401818 148586 402054
rect 148822 401818 184586 402054
rect 184822 401818 220586 402054
rect 220822 401818 544586 402054
rect 544822 401818 580586 402054
rect 580822 401818 587382 402054
rect 587618 401818 588740 402054
rect -4816 401734 588740 401818
rect -4816 401498 -3694 401734
rect -3458 401498 4586 401734
rect 4822 401498 40586 401734
rect 40822 401498 76586 401734
rect 76822 401498 112586 401734
rect 112822 401498 148586 401734
rect 148822 401498 184586 401734
rect 184822 401498 220586 401734
rect 220822 401498 544586 401734
rect 544822 401498 580586 401734
rect 580822 401498 587382 401734
rect 587618 401498 588740 401734
rect -4816 401476 588740 401498
rect -3876 401474 -3276 401476
rect 4404 401474 5004 401476
rect 40404 401474 41004 401476
rect 76404 401474 77004 401476
rect 112404 401474 113004 401476
rect 148404 401474 149004 401476
rect 184404 401474 185004 401476
rect 220404 401474 221004 401476
rect 544404 401474 545004 401476
rect 580404 401474 581004 401476
rect 587200 401474 587800 401476
rect -1996 398476 -1396 398478
rect 804 398476 1404 398478
rect 36804 398476 37404 398478
rect 72804 398476 73404 398478
rect 108804 398476 109404 398478
rect 144804 398476 145404 398478
rect 180804 398476 181404 398478
rect 216804 398476 217404 398478
rect 252804 398476 253404 398478
rect 264208 398476 264528 398478
rect 576804 398476 577404 398478
rect 585320 398476 585920 398478
rect -2936 398454 586860 398476
rect -2936 398218 -1814 398454
rect -1578 398218 986 398454
rect 1222 398218 36986 398454
rect 37222 398218 72986 398454
rect 73222 398218 108986 398454
rect 109222 398218 144986 398454
rect 145222 398218 180986 398454
rect 181222 398218 216986 398454
rect 217222 398218 252986 398454
rect 253222 398218 264250 398454
rect 264486 398218 576986 398454
rect 577222 398218 585502 398454
rect 585738 398218 586860 398454
rect -2936 398134 586860 398218
rect -2936 397898 -1814 398134
rect -1578 397898 986 398134
rect 1222 397898 36986 398134
rect 37222 397898 72986 398134
rect 73222 397898 108986 398134
rect 109222 397898 144986 398134
rect 145222 397898 180986 398134
rect 181222 397898 216986 398134
rect 217222 397898 252986 398134
rect 253222 397898 264250 398134
rect 264486 397898 576986 398134
rect 577222 397898 585502 398134
rect 585738 397898 586860 398134
rect -2936 397876 586860 397898
rect -1996 397874 -1396 397876
rect 804 397874 1404 397876
rect 36804 397874 37404 397876
rect 72804 397874 73404 397876
rect 108804 397874 109404 397876
rect 144804 397874 145404 397876
rect 180804 397874 181404 397876
rect 216804 397874 217404 397876
rect 252804 397874 253404 397876
rect 264208 397874 264528 397876
rect 576804 397874 577404 397876
rect 585320 397874 585920 397876
rect -8576 391276 -7976 391278
rect 29604 391276 30204 391278
rect 65604 391276 66204 391278
rect 101604 391276 102204 391278
rect 137604 391276 138204 391278
rect 173604 391276 174204 391278
rect 209604 391276 210204 391278
rect 245604 391276 246204 391278
rect 569604 391276 570204 391278
rect 591900 391276 592500 391278
rect -8576 391254 592500 391276
rect -8576 391018 -8394 391254
rect -8158 391018 29786 391254
rect 30022 391018 65786 391254
rect 66022 391018 101786 391254
rect 102022 391018 137786 391254
rect 138022 391018 173786 391254
rect 174022 391018 209786 391254
rect 210022 391018 245786 391254
rect 246022 391018 569786 391254
rect 570022 391018 592082 391254
rect 592318 391018 592500 391254
rect -8576 390934 592500 391018
rect -8576 390698 -8394 390934
rect -8158 390698 29786 390934
rect 30022 390698 65786 390934
rect 66022 390698 101786 390934
rect 102022 390698 137786 390934
rect 138022 390698 173786 390934
rect 174022 390698 209786 390934
rect 210022 390698 245786 390934
rect 246022 390698 569786 390934
rect 570022 390698 592082 390934
rect 592318 390698 592500 390934
rect -8576 390676 592500 390698
rect -8576 390674 -7976 390676
rect 29604 390674 30204 390676
rect 65604 390674 66204 390676
rect 101604 390674 102204 390676
rect 137604 390674 138204 390676
rect 173604 390674 174204 390676
rect 209604 390674 210204 390676
rect 245604 390674 246204 390676
rect 569604 390674 570204 390676
rect 591900 390674 592500 390676
rect -6696 387676 -6096 387678
rect 26004 387676 26604 387678
rect 62004 387676 62604 387678
rect 98004 387676 98604 387678
rect 134004 387676 134604 387678
rect 170004 387676 170604 387678
rect 206004 387676 206604 387678
rect 242004 387676 242604 387678
rect 566004 387676 566604 387678
rect 590020 387676 590620 387678
rect -6696 387654 590620 387676
rect -6696 387418 -6514 387654
rect -6278 387418 26186 387654
rect 26422 387418 62186 387654
rect 62422 387418 98186 387654
rect 98422 387418 134186 387654
rect 134422 387418 170186 387654
rect 170422 387418 206186 387654
rect 206422 387418 242186 387654
rect 242422 387418 566186 387654
rect 566422 387418 590202 387654
rect 590438 387418 590620 387654
rect -6696 387334 590620 387418
rect -6696 387098 -6514 387334
rect -6278 387098 26186 387334
rect 26422 387098 62186 387334
rect 62422 387098 98186 387334
rect 98422 387098 134186 387334
rect 134422 387098 170186 387334
rect 170422 387098 206186 387334
rect 206422 387098 242186 387334
rect 242422 387098 566186 387334
rect 566422 387098 590202 387334
rect 590438 387098 590620 387334
rect -6696 387076 590620 387098
rect -6696 387074 -6096 387076
rect 26004 387074 26604 387076
rect 62004 387074 62604 387076
rect 98004 387074 98604 387076
rect 134004 387074 134604 387076
rect 170004 387074 170604 387076
rect 206004 387074 206604 387076
rect 242004 387074 242604 387076
rect 566004 387074 566604 387076
rect 590020 387074 590620 387076
rect -4816 384076 -4216 384078
rect 22404 384076 23004 384078
rect 58404 384076 59004 384078
rect 94404 384076 95004 384078
rect 130404 384076 131004 384078
rect 166404 384076 167004 384078
rect 202404 384076 203004 384078
rect 238404 384076 239004 384078
rect 562404 384076 563004 384078
rect 588140 384076 588740 384078
rect -4816 384054 588740 384076
rect -4816 383818 -4634 384054
rect -4398 383818 22586 384054
rect 22822 383818 58586 384054
rect 58822 383818 94586 384054
rect 94822 383818 130586 384054
rect 130822 383818 166586 384054
rect 166822 383818 202586 384054
rect 202822 383818 238586 384054
rect 238822 383818 562586 384054
rect 562822 383818 588322 384054
rect 588558 383818 588740 384054
rect -4816 383734 588740 383818
rect -4816 383498 -4634 383734
rect -4398 383498 22586 383734
rect 22822 383498 58586 383734
rect 58822 383498 94586 383734
rect 94822 383498 130586 383734
rect 130822 383498 166586 383734
rect 166822 383498 202586 383734
rect 202822 383498 238586 383734
rect 238822 383498 562586 383734
rect 562822 383498 588322 383734
rect 588558 383498 588740 383734
rect -4816 383476 588740 383498
rect -4816 383474 -4216 383476
rect 22404 383474 23004 383476
rect 58404 383474 59004 383476
rect 94404 383474 95004 383476
rect 130404 383474 131004 383476
rect 166404 383474 167004 383476
rect 202404 383474 203004 383476
rect 238404 383474 239004 383476
rect 562404 383474 563004 383476
rect 588140 383474 588740 383476
rect -2936 380476 -2336 380478
rect 18804 380476 19404 380478
rect 54804 380476 55404 380478
rect 90804 380476 91404 380478
rect 126804 380476 127404 380478
rect 162804 380476 163404 380478
rect 198804 380476 199404 380478
rect 234804 380476 235404 380478
rect 279568 380476 279888 380478
rect 558804 380476 559404 380478
rect 586260 380476 586860 380478
rect -2936 380454 586860 380476
rect -2936 380218 -2754 380454
rect -2518 380218 18986 380454
rect 19222 380218 54986 380454
rect 55222 380218 90986 380454
rect 91222 380218 126986 380454
rect 127222 380218 162986 380454
rect 163222 380218 198986 380454
rect 199222 380218 234986 380454
rect 235222 380218 279610 380454
rect 279846 380218 558986 380454
rect 559222 380218 586442 380454
rect 586678 380218 586860 380454
rect -2936 380134 586860 380218
rect -2936 379898 -2754 380134
rect -2518 379898 18986 380134
rect 19222 379898 54986 380134
rect 55222 379898 90986 380134
rect 91222 379898 126986 380134
rect 127222 379898 162986 380134
rect 163222 379898 198986 380134
rect 199222 379898 234986 380134
rect 235222 379898 279610 380134
rect 279846 379898 558986 380134
rect 559222 379898 586442 380134
rect 586678 379898 586860 380134
rect -2936 379876 586860 379898
rect -2936 379874 -2336 379876
rect 18804 379874 19404 379876
rect 54804 379874 55404 379876
rect 90804 379874 91404 379876
rect 126804 379874 127404 379876
rect 162804 379874 163404 379876
rect 198804 379874 199404 379876
rect 234804 379874 235404 379876
rect 279568 379874 279888 379876
rect 558804 379874 559404 379876
rect 586260 379874 586860 379876
rect -7636 373276 -7036 373278
rect 11604 373276 12204 373278
rect 47604 373276 48204 373278
rect 83604 373276 84204 373278
rect 119604 373276 120204 373278
rect 155604 373276 156204 373278
rect 191604 373276 192204 373278
rect 227604 373276 228204 373278
rect 551604 373276 552204 373278
rect 590960 373276 591560 373278
rect -8576 373254 592500 373276
rect -8576 373018 -7454 373254
rect -7218 373018 11786 373254
rect 12022 373018 47786 373254
rect 48022 373018 83786 373254
rect 84022 373018 119786 373254
rect 120022 373018 155786 373254
rect 156022 373018 191786 373254
rect 192022 373018 227786 373254
rect 228022 373018 551786 373254
rect 552022 373018 591142 373254
rect 591378 373018 592500 373254
rect -8576 372934 592500 373018
rect -8576 372698 -7454 372934
rect -7218 372698 11786 372934
rect 12022 372698 47786 372934
rect 48022 372698 83786 372934
rect 84022 372698 119786 372934
rect 120022 372698 155786 372934
rect 156022 372698 191786 372934
rect 192022 372698 227786 372934
rect 228022 372698 551786 372934
rect 552022 372698 591142 372934
rect 591378 372698 592500 372934
rect -8576 372676 592500 372698
rect -7636 372674 -7036 372676
rect 11604 372674 12204 372676
rect 47604 372674 48204 372676
rect 83604 372674 84204 372676
rect 119604 372674 120204 372676
rect 155604 372674 156204 372676
rect 191604 372674 192204 372676
rect 227604 372674 228204 372676
rect 551604 372674 552204 372676
rect 590960 372674 591560 372676
rect -5756 369676 -5156 369678
rect 8004 369676 8604 369678
rect 44004 369676 44604 369678
rect 80004 369676 80604 369678
rect 116004 369676 116604 369678
rect 152004 369676 152604 369678
rect 188004 369676 188604 369678
rect 224004 369676 224604 369678
rect 548004 369676 548604 369678
rect 589080 369676 589680 369678
rect -6696 369654 590620 369676
rect -6696 369418 -5574 369654
rect -5338 369418 8186 369654
rect 8422 369418 44186 369654
rect 44422 369418 80186 369654
rect 80422 369418 116186 369654
rect 116422 369418 152186 369654
rect 152422 369418 188186 369654
rect 188422 369418 224186 369654
rect 224422 369418 548186 369654
rect 548422 369418 589262 369654
rect 589498 369418 590620 369654
rect -6696 369334 590620 369418
rect -6696 369098 -5574 369334
rect -5338 369098 8186 369334
rect 8422 369098 44186 369334
rect 44422 369098 80186 369334
rect 80422 369098 116186 369334
rect 116422 369098 152186 369334
rect 152422 369098 188186 369334
rect 188422 369098 224186 369334
rect 224422 369098 548186 369334
rect 548422 369098 589262 369334
rect 589498 369098 590620 369334
rect -6696 369076 590620 369098
rect -5756 369074 -5156 369076
rect 8004 369074 8604 369076
rect 44004 369074 44604 369076
rect 80004 369074 80604 369076
rect 116004 369074 116604 369076
rect 152004 369074 152604 369076
rect 188004 369074 188604 369076
rect 224004 369074 224604 369076
rect 548004 369074 548604 369076
rect 589080 369074 589680 369076
rect -3876 366076 -3276 366078
rect 4404 366076 5004 366078
rect 40404 366076 41004 366078
rect 76404 366076 77004 366078
rect 112404 366076 113004 366078
rect 148404 366076 149004 366078
rect 184404 366076 185004 366078
rect 220404 366076 221004 366078
rect 544404 366076 545004 366078
rect 580404 366076 581004 366078
rect 587200 366076 587800 366078
rect -4816 366054 588740 366076
rect -4816 365818 -3694 366054
rect -3458 365818 4586 366054
rect 4822 365818 40586 366054
rect 40822 365818 76586 366054
rect 76822 365818 112586 366054
rect 112822 365818 148586 366054
rect 148822 365818 184586 366054
rect 184822 365818 220586 366054
rect 220822 365818 544586 366054
rect 544822 365818 580586 366054
rect 580822 365818 587382 366054
rect 587618 365818 588740 366054
rect -4816 365734 588740 365818
rect -4816 365498 -3694 365734
rect -3458 365498 4586 365734
rect 4822 365498 40586 365734
rect 40822 365498 76586 365734
rect 76822 365498 112586 365734
rect 112822 365498 148586 365734
rect 148822 365498 184586 365734
rect 184822 365498 220586 365734
rect 220822 365498 544586 365734
rect 544822 365498 580586 365734
rect 580822 365498 587382 365734
rect 587618 365498 588740 365734
rect -4816 365476 588740 365498
rect -3876 365474 -3276 365476
rect 4404 365474 5004 365476
rect 40404 365474 41004 365476
rect 76404 365474 77004 365476
rect 112404 365474 113004 365476
rect 148404 365474 149004 365476
rect 184404 365474 185004 365476
rect 220404 365474 221004 365476
rect 544404 365474 545004 365476
rect 580404 365474 581004 365476
rect 587200 365474 587800 365476
rect -1996 362476 -1396 362478
rect 804 362476 1404 362478
rect 36804 362476 37404 362478
rect 72804 362476 73404 362478
rect 108804 362476 109404 362478
rect 144804 362476 145404 362478
rect 180804 362476 181404 362478
rect 216804 362476 217404 362478
rect 252804 362476 253404 362478
rect 264208 362476 264528 362478
rect 576804 362476 577404 362478
rect 585320 362476 585920 362478
rect -2936 362454 586860 362476
rect -2936 362218 -1814 362454
rect -1578 362218 986 362454
rect 1222 362218 36986 362454
rect 37222 362218 72986 362454
rect 73222 362218 108986 362454
rect 109222 362218 144986 362454
rect 145222 362218 180986 362454
rect 181222 362218 216986 362454
rect 217222 362218 252986 362454
rect 253222 362218 264250 362454
rect 264486 362218 576986 362454
rect 577222 362218 585502 362454
rect 585738 362218 586860 362454
rect -2936 362134 586860 362218
rect -2936 361898 -1814 362134
rect -1578 361898 986 362134
rect 1222 361898 36986 362134
rect 37222 361898 72986 362134
rect 73222 361898 108986 362134
rect 109222 361898 144986 362134
rect 145222 361898 180986 362134
rect 181222 361898 216986 362134
rect 217222 361898 252986 362134
rect 253222 361898 264250 362134
rect 264486 361898 576986 362134
rect 577222 361898 585502 362134
rect 585738 361898 586860 362134
rect -2936 361876 586860 361898
rect -1996 361874 -1396 361876
rect 804 361874 1404 361876
rect 36804 361874 37404 361876
rect 72804 361874 73404 361876
rect 108804 361874 109404 361876
rect 144804 361874 145404 361876
rect 180804 361874 181404 361876
rect 216804 361874 217404 361876
rect 252804 361874 253404 361876
rect 264208 361874 264528 361876
rect 576804 361874 577404 361876
rect 585320 361874 585920 361876
rect -8576 355276 -7976 355278
rect 29604 355276 30204 355278
rect 65604 355276 66204 355278
rect 101604 355276 102204 355278
rect 137604 355276 138204 355278
rect 173604 355276 174204 355278
rect 209604 355276 210204 355278
rect 245604 355276 246204 355278
rect 569604 355276 570204 355278
rect 591900 355276 592500 355278
rect -8576 355254 592500 355276
rect -8576 355018 -8394 355254
rect -8158 355018 29786 355254
rect 30022 355018 65786 355254
rect 66022 355018 101786 355254
rect 102022 355018 137786 355254
rect 138022 355018 173786 355254
rect 174022 355018 209786 355254
rect 210022 355018 245786 355254
rect 246022 355018 569786 355254
rect 570022 355018 592082 355254
rect 592318 355018 592500 355254
rect -8576 354934 592500 355018
rect -8576 354698 -8394 354934
rect -8158 354698 29786 354934
rect 30022 354698 65786 354934
rect 66022 354698 101786 354934
rect 102022 354698 137786 354934
rect 138022 354698 173786 354934
rect 174022 354698 209786 354934
rect 210022 354698 245786 354934
rect 246022 354698 569786 354934
rect 570022 354698 592082 354934
rect 592318 354698 592500 354934
rect -8576 354676 592500 354698
rect -8576 354674 -7976 354676
rect 29604 354674 30204 354676
rect 65604 354674 66204 354676
rect 101604 354674 102204 354676
rect 137604 354674 138204 354676
rect 173604 354674 174204 354676
rect 209604 354674 210204 354676
rect 245604 354674 246204 354676
rect 569604 354674 570204 354676
rect 591900 354674 592500 354676
rect -6696 351676 -6096 351678
rect 26004 351676 26604 351678
rect 62004 351676 62604 351678
rect 98004 351676 98604 351678
rect 134004 351676 134604 351678
rect 170004 351676 170604 351678
rect 206004 351676 206604 351678
rect 242004 351676 242604 351678
rect 566004 351676 566604 351678
rect 590020 351676 590620 351678
rect -6696 351654 590620 351676
rect -6696 351418 -6514 351654
rect -6278 351418 26186 351654
rect 26422 351418 62186 351654
rect 62422 351418 98186 351654
rect 98422 351418 134186 351654
rect 134422 351418 170186 351654
rect 170422 351418 206186 351654
rect 206422 351418 242186 351654
rect 242422 351418 566186 351654
rect 566422 351418 590202 351654
rect 590438 351418 590620 351654
rect -6696 351334 590620 351418
rect -6696 351098 -6514 351334
rect -6278 351098 26186 351334
rect 26422 351098 62186 351334
rect 62422 351098 98186 351334
rect 98422 351098 134186 351334
rect 134422 351098 170186 351334
rect 170422 351098 206186 351334
rect 206422 351098 242186 351334
rect 242422 351098 566186 351334
rect 566422 351098 590202 351334
rect 590438 351098 590620 351334
rect -6696 351076 590620 351098
rect -6696 351074 -6096 351076
rect 26004 351074 26604 351076
rect 62004 351074 62604 351076
rect 98004 351074 98604 351076
rect 134004 351074 134604 351076
rect 170004 351074 170604 351076
rect 206004 351074 206604 351076
rect 242004 351074 242604 351076
rect 566004 351074 566604 351076
rect 590020 351074 590620 351076
rect -4816 348076 -4216 348078
rect 22404 348076 23004 348078
rect 58404 348076 59004 348078
rect 94404 348076 95004 348078
rect 130404 348076 131004 348078
rect 166404 348076 167004 348078
rect 202404 348076 203004 348078
rect 238404 348076 239004 348078
rect 562404 348076 563004 348078
rect 588140 348076 588740 348078
rect -4816 348054 588740 348076
rect -4816 347818 -4634 348054
rect -4398 347818 22586 348054
rect 22822 347818 58586 348054
rect 58822 347818 94586 348054
rect 94822 347818 130586 348054
rect 130822 347818 166586 348054
rect 166822 347818 202586 348054
rect 202822 347818 238586 348054
rect 238822 347818 562586 348054
rect 562822 347818 588322 348054
rect 588558 347818 588740 348054
rect -4816 347734 588740 347818
rect -4816 347498 -4634 347734
rect -4398 347498 22586 347734
rect 22822 347498 58586 347734
rect 58822 347498 94586 347734
rect 94822 347498 130586 347734
rect 130822 347498 166586 347734
rect 166822 347498 202586 347734
rect 202822 347498 238586 347734
rect 238822 347498 562586 347734
rect 562822 347498 588322 347734
rect 588558 347498 588740 347734
rect -4816 347476 588740 347498
rect -4816 347474 -4216 347476
rect 22404 347474 23004 347476
rect 58404 347474 59004 347476
rect 94404 347474 95004 347476
rect 130404 347474 131004 347476
rect 166404 347474 167004 347476
rect 202404 347474 203004 347476
rect 238404 347474 239004 347476
rect 562404 347474 563004 347476
rect 588140 347474 588740 347476
rect -2936 344476 -2336 344478
rect 18804 344476 19404 344478
rect 54804 344476 55404 344478
rect 90804 344476 91404 344478
rect 126804 344476 127404 344478
rect 162804 344476 163404 344478
rect 198804 344476 199404 344478
rect 234804 344476 235404 344478
rect 279568 344476 279888 344478
rect 558804 344476 559404 344478
rect 586260 344476 586860 344478
rect -2936 344454 586860 344476
rect -2936 344218 -2754 344454
rect -2518 344218 18986 344454
rect 19222 344218 54986 344454
rect 55222 344218 90986 344454
rect 91222 344218 126986 344454
rect 127222 344218 162986 344454
rect 163222 344218 198986 344454
rect 199222 344218 234986 344454
rect 235222 344218 279610 344454
rect 279846 344218 558986 344454
rect 559222 344218 586442 344454
rect 586678 344218 586860 344454
rect -2936 344134 586860 344218
rect -2936 343898 -2754 344134
rect -2518 343898 18986 344134
rect 19222 343898 54986 344134
rect 55222 343898 90986 344134
rect 91222 343898 126986 344134
rect 127222 343898 162986 344134
rect 163222 343898 198986 344134
rect 199222 343898 234986 344134
rect 235222 343898 279610 344134
rect 279846 343898 558986 344134
rect 559222 343898 586442 344134
rect 586678 343898 586860 344134
rect -2936 343876 586860 343898
rect -2936 343874 -2336 343876
rect 18804 343874 19404 343876
rect 54804 343874 55404 343876
rect 90804 343874 91404 343876
rect 126804 343874 127404 343876
rect 162804 343874 163404 343876
rect 198804 343874 199404 343876
rect 234804 343874 235404 343876
rect 279568 343874 279888 343876
rect 558804 343874 559404 343876
rect 586260 343874 586860 343876
rect -7636 337276 -7036 337278
rect 11604 337276 12204 337278
rect 47604 337276 48204 337278
rect 83604 337276 84204 337278
rect 119604 337276 120204 337278
rect 155604 337276 156204 337278
rect 191604 337276 192204 337278
rect 227604 337276 228204 337278
rect 551604 337276 552204 337278
rect 590960 337276 591560 337278
rect -8576 337254 592500 337276
rect -8576 337018 -7454 337254
rect -7218 337018 11786 337254
rect 12022 337018 47786 337254
rect 48022 337018 83786 337254
rect 84022 337018 119786 337254
rect 120022 337018 155786 337254
rect 156022 337018 191786 337254
rect 192022 337018 227786 337254
rect 228022 337018 551786 337254
rect 552022 337018 591142 337254
rect 591378 337018 592500 337254
rect -8576 336934 592500 337018
rect -8576 336698 -7454 336934
rect -7218 336698 11786 336934
rect 12022 336698 47786 336934
rect 48022 336698 83786 336934
rect 84022 336698 119786 336934
rect 120022 336698 155786 336934
rect 156022 336698 191786 336934
rect 192022 336698 227786 336934
rect 228022 336698 551786 336934
rect 552022 336698 591142 336934
rect 591378 336698 592500 336934
rect -8576 336676 592500 336698
rect -7636 336674 -7036 336676
rect 11604 336674 12204 336676
rect 47604 336674 48204 336676
rect 83604 336674 84204 336676
rect 119604 336674 120204 336676
rect 155604 336674 156204 336676
rect 191604 336674 192204 336676
rect 227604 336674 228204 336676
rect 551604 336674 552204 336676
rect 590960 336674 591560 336676
rect -5756 333676 -5156 333678
rect 8004 333676 8604 333678
rect 44004 333676 44604 333678
rect 80004 333676 80604 333678
rect 116004 333676 116604 333678
rect 152004 333676 152604 333678
rect 188004 333676 188604 333678
rect 224004 333676 224604 333678
rect 548004 333676 548604 333678
rect 589080 333676 589680 333678
rect -6696 333654 590620 333676
rect -6696 333418 -5574 333654
rect -5338 333418 8186 333654
rect 8422 333418 44186 333654
rect 44422 333418 80186 333654
rect 80422 333418 116186 333654
rect 116422 333418 152186 333654
rect 152422 333418 188186 333654
rect 188422 333418 224186 333654
rect 224422 333418 548186 333654
rect 548422 333418 589262 333654
rect 589498 333418 590620 333654
rect -6696 333334 590620 333418
rect -6696 333098 -5574 333334
rect -5338 333098 8186 333334
rect 8422 333098 44186 333334
rect 44422 333098 80186 333334
rect 80422 333098 116186 333334
rect 116422 333098 152186 333334
rect 152422 333098 188186 333334
rect 188422 333098 224186 333334
rect 224422 333098 548186 333334
rect 548422 333098 589262 333334
rect 589498 333098 590620 333334
rect -6696 333076 590620 333098
rect -5756 333074 -5156 333076
rect 8004 333074 8604 333076
rect 44004 333074 44604 333076
rect 80004 333074 80604 333076
rect 116004 333074 116604 333076
rect 152004 333074 152604 333076
rect 188004 333074 188604 333076
rect 224004 333074 224604 333076
rect 548004 333074 548604 333076
rect 589080 333074 589680 333076
rect -3876 330076 -3276 330078
rect 4404 330076 5004 330078
rect 40404 330076 41004 330078
rect 76404 330076 77004 330078
rect 112404 330076 113004 330078
rect 148404 330076 149004 330078
rect 184404 330076 185004 330078
rect 220404 330076 221004 330078
rect 544404 330076 545004 330078
rect 580404 330076 581004 330078
rect 587200 330076 587800 330078
rect -4816 330054 588740 330076
rect -4816 329818 -3694 330054
rect -3458 329818 4586 330054
rect 4822 329818 40586 330054
rect 40822 329818 76586 330054
rect 76822 329818 112586 330054
rect 112822 329818 148586 330054
rect 148822 329818 184586 330054
rect 184822 329818 220586 330054
rect 220822 329818 544586 330054
rect 544822 329818 580586 330054
rect 580822 329818 587382 330054
rect 587618 329818 588740 330054
rect -4816 329734 588740 329818
rect -4816 329498 -3694 329734
rect -3458 329498 4586 329734
rect 4822 329498 40586 329734
rect 40822 329498 76586 329734
rect 76822 329498 112586 329734
rect 112822 329498 148586 329734
rect 148822 329498 184586 329734
rect 184822 329498 220586 329734
rect 220822 329498 544586 329734
rect 544822 329498 580586 329734
rect 580822 329498 587382 329734
rect 587618 329498 588740 329734
rect -4816 329476 588740 329498
rect -3876 329474 -3276 329476
rect 4404 329474 5004 329476
rect 40404 329474 41004 329476
rect 76404 329474 77004 329476
rect 112404 329474 113004 329476
rect 148404 329474 149004 329476
rect 184404 329474 185004 329476
rect 220404 329474 221004 329476
rect 544404 329474 545004 329476
rect 580404 329474 581004 329476
rect 587200 329474 587800 329476
rect -1996 326476 -1396 326478
rect 804 326476 1404 326478
rect 36804 326476 37404 326478
rect 72804 326476 73404 326478
rect 108804 326476 109404 326478
rect 144804 326476 145404 326478
rect 180804 326476 181404 326478
rect 216804 326476 217404 326478
rect 252804 326476 253404 326478
rect 264208 326476 264528 326478
rect 576804 326476 577404 326478
rect 585320 326476 585920 326478
rect -2936 326454 586860 326476
rect -2936 326218 -1814 326454
rect -1578 326218 986 326454
rect 1222 326218 36986 326454
rect 37222 326218 72986 326454
rect 73222 326218 108986 326454
rect 109222 326218 144986 326454
rect 145222 326218 180986 326454
rect 181222 326218 216986 326454
rect 217222 326218 252986 326454
rect 253222 326218 264250 326454
rect 264486 326218 576986 326454
rect 577222 326218 585502 326454
rect 585738 326218 586860 326454
rect -2936 326134 586860 326218
rect -2936 325898 -1814 326134
rect -1578 325898 986 326134
rect 1222 325898 36986 326134
rect 37222 325898 72986 326134
rect 73222 325898 108986 326134
rect 109222 325898 144986 326134
rect 145222 325898 180986 326134
rect 181222 325898 216986 326134
rect 217222 325898 252986 326134
rect 253222 325898 264250 326134
rect 264486 325898 576986 326134
rect 577222 325898 585502 326134
rect 585738 325898 586860 326134
rect -2936 325876 586860 325898
rect -1996 325874 -1396 325876
rect 804 325874 1404 325876
rect 36804 325874 37404 325876
rect 72804 325874 73404 325876
rect 108804 325874 109404 325876
rect 144804 325874 145404 325876
rect 180804 325874 181404 325876
rect 216804 325874 217404 325876
rect 252804 325874 253404 325876
rect 264208 325874 264528 325876
rect 576804 325874 577404 325876
rect 585320 325874 585920 325876
rect -8576 319276 -7976 319278
rect 29604 319276 30204 319278
rect 65604 319276 66204 319278
rect 101604 319276 102204 319278
rect 137604 319276 138204 319278
rect 173604 319276 174204 319278
rect 209604 319276 210204 319278
rect 245604 319276 246204 319278
rect 569604 319276 570204 319278
rect 591900 319276 592500 319278
rect -8576 319254 592500 319276
rect -8576 319018 -8394 319254
rect -8158 319018 29786 319254
rect 30022 319018 65786 319254
rect 66022 319018 101786 319254
rect 102022 319018 137786 319254
rect 138022 319018 173786 319254
rect 174022 319018 209786 319254
rect 210022 319018 245786 319254
rect 246022 319018 569786 319254
rect 570022 319018 592082 319254
rect 592318 319018 592500 319254
rect -8576 318934 592500 319018
rect -8576 318698 -8394 318934
rect -8158 318698 29786 318934
rect 30022 318698 65786 318934
rect 66022 318698 101786 318934
rect 102022 318698 137786 318934
rect 138022 318698 173786 318934
rect 174022 318698 209786 318934
rect 210022 318698 245786 318934
rect 246022 318698 569786 318934
rect 570022 318698 592082 318934
rect 592318 318698 592500 318934
rect -8576 318676 592500 318698
rect -8576 318674 -7976 318676
rect 29604 318674 30204 318676
rect 65604 318674 66204 318676
rect 101604 318674 102204 318676
rect 137604 318674 138204 318676
rect 173604 318674 174204 318676
rect 209604 318674 210204 318676
rect 245604 318674 246204 318676
rect 569604 318674 570204 318676
rect 591900 318674 592500 318676
rect -6696 315676 -6096 315678
rect 26004 315676 26604 315678
rect 62004 315676 62604 315678
rect 98004 315676 98604 315678
rect 134004 315676 134604 315678
rect 170004 315676 170604 315678
rect 206004 315676 206604 315678
rect 242004 315676 242604 315678
rect 566004 315676 566604 315678
rect 590020 315676 590620 315678
rect -6696 315654 590620 315676
rect -6696 315418 -6514 315654
rect -6278 315418 26186 315654
rect 26422 315418 62186 315654
rect 62422 315418 98186 315654
rect 98422 315418 134186 315654
rect 134422 315418 170186 315654
rect 170422 315418 206186 315654
rect 206422 315418 242186 315654
rect 242422 315418 566186 315654
rect 566422 315418 590202 315654
rect 590438 315418 590620 315654
rect -6696 315334 590620 315418
rect -6696 315098 -6514 315334
rect -6278 315098 26186 315334
rect 26422 315098 62186 315334
rect 62422 315098 98186 315334
rect 98422 315098 134186 315334
rect 134422 315098 170186 315334
rect 170422 315098 206186 315334
rect 206422 315098 242186 315334
rect 242422 315098 566186 315334
rect 566422 315098 590202 315334
rect 590438 315098 590620 315334
rect -6696 315076 590620 315098
rect -6696 315074 -6096 315076
rect 26004 315074 26604 315076
rect 62004 315074 62604 315076
rect 98004 315074 98604 315076
rect 134004 315074 134604 315076
rect 170004 315074 170604 315076
rect 206004 315074 206604 315076
rect 242004 315074 242604 315076
rect 566004 315074 566604 315076
rect 590020 315074 590620 315076
rect -4816 312076 -4216 312078
rect 22404 312076 23004 312078
rect 58404 312076 59004 312078
rect 94404 312076 95004 312078
rect 130404 312076 131004 312078
rect 166404 312076 167004 312078
rect 202404 312076 203004 312078
rect 238404 312076 239004 312078
rect 562404 312076 563004 312078
rect 588140 312076 588740 312078
rect -4816 312054 588740 312076
rect -4816 311818 -4634 312054
rect -4398 311818 22586 312054
rect 22822 311818 58586 312054
rect 58822 311818 94586 312054
rect 94822 311818 130586 312054
rect 130822 311818 166586 312054
rect 166822 311818 202586 312054
rect 202822 311818 238586 312054
rect 238822 311818 562586 312054
rect 562822 311818 588322 312054
rect 588558 311818 588740 312054
rect -4816 311734 588740 311818
rect -4816 311498 -4634 311734
rect -4398 311498 22586 311734
rect 22822 311498 58586 311734
rect 58822 311498 94586 311734
rect 94822 311498 130586 311734
rect 130822 311498 166586 311734
rect 166822 311498 202586 311734
rect 202822 311498 238586 311734
rect 238822 311498 562586 311734
rect 562822 311498 588322 311734
rect 588558 311498 588740 311734
rect -4816 311476 588740 311498
rect -4816 311474 -4216 311476
rect 22404 311474 23004 311476
rect 58404 311474 59004 311476
rect 94404 311474 95004 311476
rect 130404 311474 131004 311476
rect 166404 311474 167004 311476
rect 202404 311474 203004 311476
rect 238404 311474 239004 311476
rect 562404 311474 563004 311476
rect 588140 311474 588740 311476
rect -2936 308476 -2336 308478
rect 18804 308476 19404 308478
rect 54804 308476 55404 308478
rect 90804 308476 91404 308478
rect 126804 308476 127404 308478
rect 162804 308476 163404 308478
rect 198804 308476 199404 308478
rect 234804 308476 235404 308478
rect 279568 308476 279888 308478
rect 558804 308476 559404 308478
rect 586260 308476 586860 308478
rect -2936 308454 586860 308476
rect -2936 308218 -2754 308454
rect -2518 308218 18986 308454
rect 19222 308218 54986 308454
rect 55222 308218 90986 308454
rect 91222 308218 126986 308454
rect 127222 308218 162986 308454
rect 163222 308218 198986 308454
rect 199222 308218 234986 308454
rect 235222 308218 279610 308454
rect 279846 308218 558986 308454
rect 559222 308218 586442 308454
rect 586678 308218 586860 308454
rect -2936 308134 586860 308218
rect -2936 307898 -2754 308134
rect -2518 307898 18986 308134
rect 19222 307898 54986 308134
rect 55222 307898 90986 308134
rect 91222 307898 126986 308134
rect 127222 307898 162986 308134
rect 163222 307898 198986 308134
rect 199222 307898 234986 308134
rect 235222 307898 279610 308134
rect 279846 307898 558986 308134
rect 559222 307898 586442 308134
rect 586678 307898 586860 308134
rect -2936 307876 586860 307898
rect -2936 307874 -2336 307876
rect 18804 307874 19404 307876
rect 54804 307874 55404 307876
rect 90804 307874 91404 307876
rect 126804 307874 127404 307876
rect 162804 307874 163404 307876
rect 198804 307874 199404 307876
rect 234804 307874 235404 307876
rect 279568 307874 279888 307876
rect 558804 307874 559404 307876
rect 586260 307874 586860 307876
rect -7636 301276 -7036 301278
rect 11604 301276 12204 301278
rect 47604 301276 48204 301278
rect 83604 301276 84204 301278
rect 119604 301276 120204 301278
rect 155604 301276 156204 301278
rect 191604 301276 192204 301278
rect 227604 301276 228204 301278
rect 551604 301276 552204 301278
rect 590960 301276 591560 301278
rect -8576 301254 592500 301276
rect -8576 301018 -7454 301254
rect -7218 301018 11786 301254
rect 12022 301018 47786 301254
rect 48022 301018 83786 301254
rect 84022 301018 119786 301254
rect 120022 301018 155786 301254
rect 156022 301018 191786 301254
rect 192022 301018 227786 301254
rect 228022 301018 551786 301254
rect 552022 301018 591142 301254
rect 591378 301018 592500 301254
rect -8576 300934 592500 301018
rect -8576 300698 -7454 300934
rect -7218 300698 11786 300934
rect 12022 300698 47786 300934
rect 48022 300698 83786 300934
rect 84022 300698 119786 300934
rect 120022 300698 155786 300934
rect 156022 300698 191786 300934
rect 192022 300698 227786 300934
rect 228022 300698 551786 300934
rect 552022 300698 591142 300934
rect 591378 300698 592500 300934
rect -8576 300676 592500 300698
rect -7636 300674 -7036 300676
rect 11604 300674 12204 300676
rect 47604 300674 48204 300676
rect 83604 300674 84204 300676
rect 119604 300674 120204 300676
rect 155604 300674 156204 300676
rect 191604 300674 192204 300676
rect 227604 300674 228204 300676
rect 551604 300674 552204 300676
rect 590960 300674 591560 300676
rect -5756 297676 -5156 297678
rect 8004 297676 8604 297678
rect 44004 297676 44604 297678
rect 80004 297676 80604 297678
rect 116004 297676 116604 297678
rect 152004 297676 152604 297678
rect 188004 297676 188604 297678
rect 224004 297676 224604 297678
rect 548004 297676 548604 297678
rect 589080 297676 589680 297678
rect -6696 297654 590620 297676
rect -6696 297418 -5574 297654
rect -5338 297418 8186 297654
rect 8422 297418 44186 297654
rect 44422 297418 80186 297654
rect 80422 297418 116186 297654
rect 116422 297418 152186 297654
rect 152422 297418 188186 297654
rect 188422 297418 224186 297654
rect 224422 297418 548186 297654
rect 548422 297418 589262 297654
rect 589498 297418 590620 297654
rect -6696 297334 590620 297418
rect -6696 297098 -5574 297334
rect -5338 297098 8186 297334
rect 8422 297098 44186 297334
rect 44422 297098 80186 297334
rect 80422 297098 116186 297334
rect 116422 297098 152186 297334
rect 152422 297098 188186 297334
rect 188422 297098 224186 297334
rect 224422 297098 548186 297334
rect 548422 297098 589262 297334
rect 589498 297098 590620 297334
rect -6696 297076 590620 297098
rect -5756 297074 -5156 297076
rect 8004 297074 8604 297076
rect 44004 297074 44604 297076
rect 80004 297074 80604 297076
rect 116004 297074 116604 297076
rect 152004 297074 152604 297076
rect 188004 297074 188604 297076
rect 224004 297074 224604 297076
rect 548004 297074 548604 297076
rect 589080 297074 589680 297076
rect -3876 294076 -3276 294078
rect 4404 294076 5004 294078
rect 40404 294076 41004 294078
rect 76404 294076 77004 294078
rect 112404 294076 113004 294078
rect 148404 294076 149004 294078
rect 184404 294076 185004 294078
rect 220404 294076 221004 294078
rect 544404 294076 545004 294078
rect 580404 294076 581004 294078
rect 587200 294076 587800 294078
rect -4816 294054 588740 294076
rect -4816 293818 -3694 294054
rect -3458 293818 4586 294054
rect 4822 293818 40586 294054
rect 40822 293818 76586 294054
rect 76822 293818 112586 294054
rect 112822 293818 148586 294054
rect 148822 293818 184586 294054
rect 184822 293818 220586 294054
rect 220822 293818 544586 294054
rect 544822 293818 580586 294054
rect 580822 293818 587382 294054
rect 587618 293818 588740 294054
rect -4816 293734 588740 293818
rect -4816 293498 -3694 293734
rect -3458 293498 4586 293734
rect 4822 293498 40586 293734
rect 40822 293498 76586 293734
rect 76822 293498 112586 293734
rect 112822 293498 148586 293734
rect 148822 293498 184586 293734
rect 184822 293498 220586 293734
rect 220822 293498 544586 293734
rect 544822 293498 580586 293734
rect 580822 293498 587382 293734
rect 587618 293498 588740 293734
rect -4816 293476 588740 293498
rect -3876 293474 -3276 293476
rect 4404 293474 5004 293476
rect 40404 293474 41004 293476
rect 76404 293474 77004 293476
rect 112404 293474 113004 293476
rect 148404 293474 149004 293476
rect 184404 293474 185004 293476
rect 220404 293474 221004 293476
rect 544404 293474 545004 293476
rect 580404 293474 581004 293476
rect 587200 293474 587800 293476
rect -1996 290476 -1396 290478
rect 804 290476 1404 290478
rect 36804 290476 37404 290478
rect 72804 290476 73404 290478
rect 108804 290476 109404 290478
rect 144804 290476 145404 290478
rect 180804 290476 181404 290478
rect 216804 290476 217404 290478
rect 252804 290476 253404 290478
rect 264208 290476 264528 290478
rect 576804 290476 577404 290478
rect 585320 290476 585920 290478
rect -2936 290454 586860 290476
rect -2936 290218 -1814 290454
rect -1578 290218 986 290454
rect 1222 290218 36986 290454
rect 37222 290218 72986 290454
rect 73222 290218 108986 290454
rect 109222 290218 144986 290454
rect 145222 290218 180986 290454
rect 181222 290218 216986 290454
rect 217222 290218 252986 290454
rect 253222 290218 264250 290454
rect 264486 290218 576986 290454
rect 577222 290218 585502 290454
rect 585738 290218 586860 290454
rect -2936 290134 586860 290218
rect -2936 289898 -1814 290134
rect -1578 289898 986 290134
rect 1222 289898 36986 290134
rect 37222 289898 72986 290134
rect 73222 289898 108986 290134
rect 109222 289898 144986 290134
rect 145222 289898 180986 290134
rect 181222 289898 216986 290134
rect 217222 289898 252986 290134
rect 253222 289898 264250 290134
rect 264486 289898 576986 290134
rect 577222 289898 585502 290134
rect 585738 289898 586860 290134
rect -2936 289876 586860 289898
rect -1996 289874 -1396 289876
rect 804 289874 1404 289876
rect 36804 289874 37404 289876
rect 72804 289874 73404 289876
rect 108804 289874 109404 289876
rect 144804 289874 145404 289876
rect 180804 289874 181404 289876
rect 216804 289874 217404 289876
rect 252804 289874 253404 289876
rect 264208 289874 264528 289876
rect 576804 289874 577404 289876
rect 585320 289874 585920 289876
rect -8576 283276 -7976 283278
rect 29604 283276 30204 283278
rect 65604 283276 66204 283278
rect 101604 283276 102204 283278
rect 137604 283276 138204 283278
rect 173604 283276 174204 283278
rect 209604 283276 210204 283278
rect 245604 283276 246204 283278
rect 569604 283276 570204 283278
rect 591900 283276 592500 283278
rect -8576 283254 592500 283276
rect -8576 283018 -8394 283254
rect -8158 283018 29786 283254
rect 30022 283018 65786 283254
rect 66022 283018 101786 283254
rect 102022 283018 137786 283254
rect 138022 283018 173786 283254
rect 174022 283018 209786 283254
rect 210022 283018 245786 283254
rect 246022 283018 569786 283254
rect 570022 283018 592082 283254
rect 592318 283018 592500 283254
rect -8576 282934 592500 283018
rect -8576 282698 -8394 282934
rect -8158 282698 29786 282934
rect 30022 282698 65786 282934
rect 66022 282698 101786 282934
rect 102022 282698 137786 282934
rect 138022 282698 173786 282934
rect 174022 282698 209786 282934
rect 210022 282698 245786 282934
rect 246022 282698 569786 282934
rect 570022 282698 592082 282934
rect 592318 282698 592500 282934
rect -8576 282676 592500 282698
rect -8576 282674 -7976 282676
rect 29604 282674 30204 282676
rect 65604 282674 66204 282676
rect 101604 282674 102204 282676
rect 137604 282674 138204 282676
rect 173604 282674 174204 282676
rect 209604 282674 210204 282676
rect 245604 282674 246204 282676
rect 569604 282674 570204 282676
rect 591900 282674 592500 282676
rect -6696 279676 -6096 279678
rect 26004 279676 26604 279678
rect 62004 279676 62604 279678
rect 98004 279676 98604 279678
rect 134004 279676 134604 279678
rect 170004 279676 170604 279678
rect 206004 279676 206604 279678
rect 242004 279676 242604 279678
rect 566004 279676 566604 279678
rect 590020 279676 590620 279678
rect -6696 279654 590620 279676
rect -6696 279418 -6514 279654
rect -6278 279418 26186 279654
rect 26422 279418 62186 279654
rect 62422 279418 98186 279654
rect 98422 279418 134186 279654
rect 134422 279418 170186 279654
rect 170422 279418 206186 279654
rect 206422 279418 242186 279654
rect 242422 279418 566186 279654
rect 566422 279418 590202 279654
rect 590438 279418 590620 279654
rect -6696 279334 590620 279418
rect -6696 279098 -6514 279334
rect -6278 279098 26186 279334
rect 26422 279098 62186 279334
rect 62422 279098 98186 279334
rect 98422 279098 134186 279334
rect 134422 279098 170186 279334
rect 170422 279098 206186 279334
rect 206422 279098 242186 279334
rect 242422 279098 566186 279334
rect 566422 279098 590202 279334
rect 590438 279098 590620 279334
rect -6696 279076 590620 279098
rect -6696 279074 -6096 279076
rect 26004 279074 26604 279076
rect 62004 279074 62604 279076
rect 98004 279074 98604 279076
rect 134004 279074 134604 279076
rect 170004 279074 170604 279076
rect 206004 279074 206604 279076
rect 242004 279074 242604 279076
rect 566004 279074 566604 279076
rect 590020 279074 590620 279076
rect -4816 276076 -4216 276078
rect 22404 276076 23004 276078
rect 58404 276076 59004 276078
rect 94404 276076 95004 276078
rect 130404 276076 131004 276078
rect 166404 276076 167004 276078
rect 202404 276076 203004 276078
rect 238404 276076 239004 276078
rect 562404 276076 563004 276078
rect 588140 276076 588740 276078
rect -4816 276054 588740 276076
rect -4816 275818 -4634 276054
rect -4398 275818 22586 276054
rect 22822 275818 58586 276054
rect 58822 275818 94586 276054
rect 94822 275818 130586 276054
rect 130822 275818 166586 276054
rect 166822 275818 202586 276054
rect 202822 275818 238586 276054
rect 238822 275818 562586 276054
rect 562822 275818 588322 276054
rect 588558 275818 588740 276054
rect -4816 275734 588740 275818
rect -4816 275498 -4634 275734
rect -4398 275498 22586 275734
rect 22822 275498 58586 275734
rect 58822 275498 94586 275734
rect 94822 275498 130586 275734
rect 130822 275498 166586 275734
rect 166822 275498 202586 275734
rect 202822 275498 238586 275734
rect 238822 275498 562586 275734
rect 562822 275498 588322 275734
rect 588558 275498 588740 275734
rect -4816 275476 588740 275498
rect -4816 275474 -4216 275476
rect 22404 275474 23004 275476
rect 58404 275474 59004 275476
rect 94404 275474 95004 275476
rect 130404 275474 131004 275476
rect 166404 275474 167004 275476
rect 202404 275474 203004 275476
rect 238404 275474 239004 275476
rect 562404 275474 563004 275476
rect 588140 275474 588740 275476
rect -2936 272476 -2336 272478
rect 18804 272476 19404 272478
rect 54804 272476 55404 272478
rect 90804 272476 91404 272478
rect 126804 272476 127404 272478
rect 162804 272476 163404 272478
rect 198804 272476 199404 272478
rect 234804 272476 235404 272478
rect 279568 272476 279888 272478
rect 558804 272476 559404 272478
rect 586260 272476 586860 272478
rect -2936 272454 586860 272476
rect -2936 272218 -2754 272454
rect -2518 272218 18986 272454
rect 19222 272218 54986 272454
rect 55222 272218 90986 272454
rect 91222 272218 126986 272454
rect 127222 272218 162986 272454
rect 163222 272218 198986 272454
rect 199222 272218 234986 272454
rect 235222 272218 279610 272454
rect 279846 272218 558986 272454
rect 559222 272218 586442 272454
rect 586678 272218 586860 272454
rect -2936 272134 586860 272218
rect -2936 271898 -2754 272134
rect -2518 271898 18986 272134
rect 19222 271898 54986 272134
rect 55222 271898 90986 272134
rect 91222 271898 126986 272134
rect 127222 271898 162986 272134
rect 163222 271898 198986 272134
rect 199222 271898 234986 272134
rect 235222 271898 279610 272134
rect 279846 271898 558986 272134
rect 559222 271898 586442 272134
rect 586678 271898 586860 272134
rect -2936 271876 586860 271898
rect -2936 271874 -2336 271876
rect 18804 271874 19404 271876
rect 54804 271874 55404 271876
rect 90804 271874 91404 271876
rect 126804 271874 127404 271876
rect 162804 271874 163404 271876
rect 198804 271874 199404 271876
rect 234804 271874 235404 271876
rect 279568 271874 279888 271876
rect 558804 271874 559404 271876
rect 586260 271874 586860 271876
rect -7636 265276 -7036 265278
rect 11604 265276 12204 265278
rect 47604 265276 48204 265278
rect 83604 265276 84204 265278
rect 119604 265276 120204 265278
rect 155604 265276 156204 265278
rect 191604 265276 192204 265278
rect 227604 265276 228204 265278
rect 551604 265276 552204 265278
rect 590960 265276 591560 265278
rect -8576 265254 592500 265276
rect -8576 265018 -7454 265254
rect -7218 265018 11786 265254
rect 12022 265018 47786 265254
rect 48022 265018 83786 265254
rect 84022 265018 119786 265254
rect 120022 265018 155786 265254
rect 156022 265018 191786 265254
rect 192022 265018 227786 265254
rect 228022 265018 551786 265254
rect 552022 265018 591142 265254
rect 591378 265018 592500 265254
rect -8576 264934 592500 265018
rect -8576 264698 -7454 264934
rect -7218 264698 11786 264934
rect 12022 264698 47786 264934
rect 48022 264698 83786 264934
rect 84022 264698 119786 264934
rect 120022 264698 155786 264934
rect 156022 264698 191786 264934
rect 192022 264698 227786 264934
rect 228022 264698 551786 264934
rect 552022 264698 591142 264934
rect 591378 264698 592500 264934
rect -8576 264676 592500 264698
rect -7636 264674 -7036 264676
rect 11604 264674 12204 264676
rect 47604 264674 48204 264676
rect 83604 264674 84204 264676
rect 119604 264674 120204 264676
rect 155604 264674 156204 264676
rect 191604 264674 192204 264676
rect 227604 264674 228204 264676
rect 551604 264674 552204 264676
rect 590960 264674 591560 264676
rect -5756 261676 -5156 261678
rect 8004 261676 8604 261678
rect 44004 261676 44604 261678
rect 80004 261676 80604 261678
rect 116004 261676 116604 261678
rect 152004 261676 152604 261678
rect 188004 261676 188604 261678
rect 224004 261676 224604 261678
rect 548004 261676 548604 261678
rect 589080 261676 589680 261678
rect -6696 261654 590620 261676
rect -6696 261418 -5574 261654
rect -5338 261418 8186 261654
rect 8422 261418 44186 261654
rect 44422 261418 80186 261654
rect 80422 261418 116186 261654
rect 116422 261418 152186 261654
rect 152422 261418 188186 261654
rect 188422 261418 224186 261654
rect 224422 261418 548186 261654
rect 548422 261418 589262 261654
rect 589498 261418 590620 261654
rect -6696 261334 590620 261418
rect -6696 261098 -5574 261334
rect -5338 261098 8186 261334
rect 8422 261098 44186 261334
rect 44422 261098 80186 261334
rect 80422 261098 116186 261334
rect 116422 261098 152186 261334
rect 152422 261098 188186 261334
rect 188422 261098 224186 261334
rect 224422 261098 548186 261334
rect 548422 261098 589262 261334
rect 589498 261098 590620 261334
rect -6696 261076 590620 261098
rect -5756 261074 -5156 261076
rect 8004 261074 8604 261076
rect 44004 261074 44604 261076
rect 80004 261074 80604 261076
rect 116004 261074 116604 261076
rect 152004 261074 152604 261076
rect 188004 261074 188604 261076
rect 224004 261074 224604 261076
rect 548004 261074 548604 261076
rect 589080 261074 589680 261076
rect -3876 258076 -3276 258078
rect 4404 258076 5004 258078
rect 40404 258076 41004 258078
rect 76404 258076 77004 258078
rect 112404 258076 113004 258078
rect 148404 258076 149004 258078
rect 184404 258076 185004 258078
rect 220404 258076 221004 258078
rect 544404 258076 545004 258078
rect 580404 258076 581004 258078
rect 587200 258076 587800 258078
rect -4816 258054 588740 258076
rect -4816 257818 -3694 258054
rect -3458 257818 4586 258054
rect 4822 257818 40586 258054
rect 40822 257818 76586 258054
rect 76822 257818 112586 258054
rect 112822 257818 148586 258054
rect 148822 257818 184586 258054
rect 184822 257818 220586 258054
rect 220822 257818 544586 258054
rect 544822 257818 580586 258054
rect 580822 257818 587382 258054
rect 587618 257818 588740 258054
rect -4816 257734 588740 257818
rect -4816 257498 -3694 257734
rect -3458 257498 4586 257734
rect 4822 257498 40586 257734
rect 40822 257498 76586 257734
rect 76822 257498 112586 257734
rect 112822 257498 148586 257734
rect 148822 257498 184586 257734
rect 184822 257498 220586 257734
rect 220822 257498 544586 257734
rect 544822 257498 580586 257734
rect 580822 257498 587382 257734
rect 587618 257498 588740 257734
rect -4816 257476 588740 257498
rect -3876 257474 -3276 257476
rect 4404 257474 5004 257476
rect 40404 257474 41004 257476
rect 76404 257474 77004 257476
rect 112404 257474 113004 257476
rect 148404 257474 149004 257476
rect 184404 257474 185004 257476
rect 220404 257474 221004 257476
rect 544404 257474 545004 257476
rect 580404 257474 581004 257476
rect 587200 257474 587800 257476
rect -1996 254476 -1396 254478
rect 804 254476 1404 254478
rect 36804 254476 37404 254478
rect 72804 254476 73404 254478
rect 108804 254476 109404 254478
rect 144804 254476 145404 254478
rect 180804 254476 181404 254478
rect 216804 254476 217404 254478
rect 252804 254476 253404 254478
rect 264208 254476 264528 254478
rect 576804 254476 577404 254478
rect 585320 254476 585920 254478
rect -2936 254454 586860 254476
rect -2936 254218 -1814 254454
rect -1578 254218 986 254454
rect 1222 254218 36986 254454
rect 37222 254218 72986 254454
rect 73222 254218 108986 254454
rect 109222 254218 144986 254454
rect 145222 254218 180986 254454
rect 181222 254218 216986 254454
rect 217222 254218 252986 254454
rect 253222 254218 264250 254454
rect 264486 254218 576986 254454
rect 577222 254218 585502 254454
rect 585738 254218 586860 254454
rect -2936 254134 586860 254218
rect -2936 253898 -1814 254134
rect -1578 253898 986 254134
rect 1222 253898 36986 254134
rect 37222 253898 72986 254134
rect 73222 253898 108986 254134
rect 109222 253898 144986 254134
rect 145222 253898 180986 254134
rect 181222 253898 216986 254134
rect 217222 253898 252986 254134
rect 253222 253898 264250 254134
rect 264486 253898 576986 254134
rect 577222 253898 585502 254134
rect 585738 253898 586860 254134
rect -2936 253876 586860 253898
rect -1996 253874 -1396 253876
rect 804 253874 1404 253876
rect 36804 253874 37404 253876
rect 72804 253874 73404 253876
rect 108804 253874 109404 253876
rect 144804 253874 145404 253876
rect 180804 253874 181404 253876
rect 216804 253874 217404 253876
rect 252804 253874 253404 253876
rect 264208 253874 264528 253876
rect 576804 253874 577404 253876
rect 585320 253874 585920 253876
rect -8576 247276 -7976 247278
rect 29604 247276 30204 247278
rect 65604 247276 66204 247278
rect 101604 247276 102204 247278
rect 137604 247276 138204 247278
rect 173604 247276 174204 247278
rect 209604 247276 210204 247278
rect 245604 247276 246204 247278
rect 569604 247276 570204 247278
rect 591900 247276 592500 247278
rect -8576 247254 592500 247276
rect -8576 247018 -8394 247254
rect -8158 247018 29786 247254
rect 30022 247018 65786 247254
rect 66022 247018 101786 247254
rect 102022 247018 137786 247254
rect 138022 247018 173786 247254
rect 174022 247018 209786 247254
rect 210022 247018 245786 247254
rect 246022 247018 569786 247254
rect 570022 247018 592082 247254
rect 592318 247018 592500 247254
rect -8576 246934 592500 247018
rect -8576 246698 -8394 246934
rect -8158 246698 29786 246934
rect 30022 246698 65786 246934
rect 66022 246698 101786 246934
rect 102022 246698 137786 246934
rect 138022 246698 173786 246934
rect 174022 246698 209786 246934
rect 210022 246698 245786 246934
rect 246022 246698 569786 246934
rect 570022 246698 592082 246934
rect 592318 246698 592500 246934
rect -8576 246676 592500 246698
rect -8576 246674 -7976 246676
rect 29604 246674 30204 246676
rect 65604 246674 66204 246676
rect 101604 246674 102204 246676
rect 137604 246674 138204 246676
rect 173604 246674 174204 246676
rect 209604 246674 210204 246676
rect 245604 246674 246204 246676
rect 569604 246674 570204 246676
rect 591900 246674 592500 246676
rect -6696 243676 -6096 243678
rect 26004 243676 26604 243678
rect 62004 243676 62604 243678
rect 98004 243676 98604 243678
rect 134004 243676 134604 243678
rect 170004 243676 170604 243678
rect 206004 243676 206604 243678
rect 242004 243676 242604 243678
rect 566004 243676 566604 243678
rect 590020 243676 590620 243678
rect -6696 243654 590620 243676
rect -6696 243418 -6514 243654
rect -6278 243418 26186 243654
rect 26422 243418 62186 243654
rect 62422 243418 98186 243654
rect 98422 243418 134186 243654
rect 134422 243418 170186 243654
rect 170422 243418 206186 243654
rect 206422 243418 242186 243654
rect 242422 243418 566186 243654
rect 566422 243418 590202 243654
rect 590438 243418 590620 243654
rect -6696 243334 590620 243418
rect -6696 243098 -6514 243334
rect -6278 243098 26186 243334
rect 26422 243098 62186 243334
rect 62422 243098 98186 243334
rect 98422 243098 134186 243334
rect 134422 243098 170186 243334
rect 170422 243098 206186 243334
rect 206422 243098 242186 243334
rect 242422 243098 566186 243334
rect 566422 243098 590202 243334
rect 590438 243098 590620 243334
rect -6696 243076 590620 243098
rect -6696 243074 -6096 243076
rect 26004 243074 26604 243076
rect 62004 243074 62604 243076
rect 98004 243074 98604 243076
rect 134004 243074 134604 243076
rect 170004 243074 170604 243076
rect 206004 243074 206604 243076
rect 242004 243074 242604 243076
rect 566004 243074 566604 243076
rect 590020 243074 590620 243076
rect -4816 240076 -4216 240078
rect 22404 240076 23004 240078
rect 58404 240076 59004 240078
rect 94404 240076 95004 240078
rect 130404 240076 131004 240078
rect 166404 240076 167004 240078
rect 202404 240076 203004 240078
rect 238404 240076 239004 240078
rect 562404 240076 563004 240078
rect 588140 240076 588740 240078
rect -4816 240054 588740 240076
rect -4816 239818 -4634 240054
rect -4398 239818 22586 240054
rect 22822 239818 58586 240054
rect 58822 239818 94586 240054
rect 94822 239818 130586 240054
rect 130822 239818 166586 240054
rect 166822 239818 202586 240054
rect 202822 239818 238586 240054
rect 238822 239818 562586 240054
rect 562822 239818 588322 240054
rect 588558 239818 588740 240054
rect -4816 239734 588740 239818
rect -4816 239498 -4634 239734
rect -4398 239498 22586 239734
rect 22822 239498 58586 239734
rect 58822 239498 94586 239734
rect 94822 239498 130586 239734
rect 130822 239498 166586 239734
rect 166822 239498 202586 239734
rect 202822 239498 238586 239734
rect 238822 239498 562586 239734
rect 562822 239498 588322 239734
rect 588558 239498 588740 239734
rect -4816 239476 588740 239498
rect -4816 239474 -4216 239476
rect 22404 239474 23004 239476
rect 58404 239474 59004 239476
rect 94404 239474 95004 239476
rect 130404 239474 131004 239476
rect 166404 239474 167004 239476
rect 202404 239474 203004 239476
rect 238404 239474 239004 239476
rect 562404 239474 563004 239476
rect 588140 239474 588740 239476
rect -2936 236476 -2336 236478
rect 18804 236476 19404 236478
rect 54804 236476 55404 236478
rect 90804 236476 91404 236478
rect 126804 236476 127404 236478
rect 162804 236476 163404 236478
rect 198804 236476 199404 236478
rect 234804 236476 235404 236478
rect 270804 236476 271404 236478
rect 306804 236476 307404 236478
rect 342804 236476 343404 236478
rect 378804 236476 379404 236478
rect 414804 236476 415404 236478
rect 450804 236476 451404 236478
rect 486804 236476 487404 236478
rect 522804 236476 523404 236478
rect 558804 236476 559404 236478
rect 586260 236476 586860 236478
rect -2936 236454 586860 236476
rect -2936 236218 -2754 236454
rect -2518 236218 18986 236454
rect 19222 236218 54986 236454
rect 55222 236218 90986 236454
rect 91222 236218 126986 236454
rect 127222 236218 162986 236454
rect 163222 236218 198986 236454
rect 199222 236218 234986 236454
rect 235222 236218 270986 236454
rect 271222 236218 306986 236454
rect 307222 236218 342986 236454
rect 343222 236218 378986 236454
rect 379222 236218 414986 236454
rect 415222 236218 450986 236454
rect 451222 236218 486986 236454
rect 487222 236218 522986 236454
rect 523222 236218 558986 236454
rect 559222 236218 586442 236454
rect 586678 236218 586860 236454
rect -2936 236134 586860 236218
rect -2936 235898 -2754 236134
rect -2518 235898 18986 236134
rect 19222 235898 54986 236134
rect 55222 235898 90986 236134
rect 91222 235898 126986 236134
rect 127222 235898 162986 236134
rect 163222 235898 198986 236134
rect 199222 235898 234986 236134
rect 235222 235898 270986 236134
rect 271222 235898 306986 236134
rect 307222 235898 342986 236134
rect 343222 235898 378986 236134
rect 379222 235898 414986 236134
rect 415222 235898 450986 236134
rect 451222 235898 486986 236134
rect 487222 235898 522986 236134
rect 523222 235898 558986 236134
rect 559222 235898 586442 236134
rect 586678 235898 586860 236134
rect -2936 235876 586860 235898
rect -2936 235874 -2336 235876
rect 18804 235874 19404 235876
rect 54804 235874 55404 235876
rect 90804 235874 91404 235876
rect 126804 235874 127404 235876
rect 162804 235874 163404 235876
rect 198804 235874 199404 235876
rect 234804 235874 235404 235876
rect 270804 235874 271404 235876
rect 306804 235874 307404 235876
rect 342804 235874 343404 235876
rect 378804 235874 379404 235876
rect 414804 235874 415404 235876
rect 450804 235874 451404 235876
rect 486804 235874 487404 235876
rect 522804 235874 523404 235876
rect 558804 235874 559404 235876
rect 586260 235874 586860 235876
rect -7636 229276 -7036 229278
rect 11604 229276 12204 229278
rect 47604 229276 48204 229278
rect 83604 229276 84204 229278
rect 119604 229276 120204 229278
rect 155604 229276 156204 229278
rect 191604 229276 192204 229278
rect 227604 229276 228204 229278
rect 263604 229276 264204 229278
rect 299604 229276 300204 229278
rect 335604 229276 336204 229278
rect 371604 229276 372204 229278
rect 407604 229276 408204 229278
rect 443604 229276 444204 229278
rect 479604 229276 480204 229278
rect 515604 229276 516204 229278
rect 551604 229276 552204 229278
rect 590960 229276 591560 229278
rect -8576 229254 592500 229276
rect -8576 229018 -7454 229254
rect -7218 229018 11786 229254
rect 12022 229018 47786 229254
rect 48022 229018 83786 229254
rect 84022 229018 119786 229254
rect 120022 229018 155786 229254
rect 156022 229018 191786 229254
rect 192022 229018 227786 229254
rect 228022 229018 263786 229254
rect 264022 229018 299786 229254
rect 300022 229018 335786 229254
rect 336022 229018 371786 229254
rect 372022 229018 407786 229254
rect 408022 229018 443786 229254
rect 444022 229018 479786 229254
rect 480022 229018 515786 229254
rect 516022 229018 551786 229254
rect 552022 229018 591142 229254
rect 591378 229018 592500 229254
rect -8576 228934 592500 229018
rect -8576 228698 -7454 228934
rect -7218 228698 11786 228934
rect 12022 228698 47786 228934
rect 48022 228698 83786 228934
rect 84022 228698 119786 228934
rect 120022 228698 155786 228934
rect 156022 228698 191786 228934
rect 192022 228698 227786 228934
rect 228022 228698 263786 228934
rect 264022 228698 299786 228934
rect 300022 228698 335786 228934
rect 336022 228698 371786 228934
rect 372022 228698 407786 228934
rect 408022 228698 443786 228934
rect 444022 228698 479786 228934
rect 480022 228698 515786 228934
rect 516022 228698 551786 228934
rect 552022 228698 591142 228934
rect 591378 228698 592500 228934
rect -8576 228676 592500 228698
rect -7636 228674 -7036 228676
rect 11604 228674 12204 228676
rect 47604 228674 48204 228676
rect 83604 228674 84204 228676
rect 119604 228674 120204 228676
rect 155604 228674 156204 228676
rect 191604 228674 192204 228676
rect 227604 228674 228204 228676
rect 263604 228674 264204 228676
rect 299604 228674 300204 228676
rect 335604 228674 336204 228676
rect 371604 228674 372204 228676
rect 407604 228674 408204 228676
rect 443604 228674 444204 228676
rect 479604 228674 480204 228676
rect 515604 228674 516204 228676
rect 551604 228674 552204 228676
rect 590960 228674 591560 228676
rect -5756 225676 -5156 225678
rect 8004 225676 8604 225678
rect 44004 225676 44604 225678
rect 80004 225676 80604 225678
rect 116004 225676 116604 225678
rect 152004 225676 152604 225678
rect 188004 225676 188604 225678
rect 224004 225676 224604 225678
rect 260004 225676 260604 225678
rect 296004 225676 296604 225678
rect 332004 225676 332604 225678
rect 368004 225676 368604 225678
rect 404004 225676 404604 225678
rect 440004 225676 440604 225678
rect 476004 225676 476604 225678
rect 512004 225676 512604 225678
rect 548004 225676 548604 225678
rect 589080 225676 589680 225678
rect -6696 225654 590620 225676
rect -6696 225418 -5574 225654
rect -5338 225418 8186 225654
rect 8422 225418 44186 225654
rect 44422 225418 80186 225654
rect 80422 225418 116186 225654
rect 116422 225418 152186 225654
rect 152422 225418 188186 225654
rect 188422 225418 224186 225654
rect 224422 225418 260186 225654
rect 260422 225418 296186 225654
rect 296422 225418 332186 225654
rect 332422 225418 368186 225654
rect 368422 225418 404186 225654
rect 404422 225418 440186 225654
rect 440422 225418 476186 225654
rect 476422 225418 512186 225654
rect 512422 225418 548186 225654
rect 548422 225418 589262 225654
rect 589498 225418 590620 225654
rect -6696 225334 590620 225418
rect -6696 225098 -5574 225334
rect -5338 225098 8186 225334
rect 8422 225098 44186 225334
rect 44422 225098 80186 225334
rect 80422 225098 116186 225334
rect 116422 225098 152186 225334
rect 152422 225098 188186 225334
rect 188422 225098 224186 225334
rect 224422 225098 260186 225334
rect 260422 225098 296186 225334
rect 296422 225098 332186 225334
rect 332422 225098 368186 225334
rect 368422 225098 404186 225334
rect 404422 225098 440186 225334
rect 440422 225098 476186 225334
rect 476422 225098 512186 225334
rect 512422 225098 548186 225334
rect 548422 225098 589262 225334
rect 589498 225098 590620 225334
rect -6696 225076 590620 225098
rect -5756 225074 -5156 225076
rect 8004 225074 8604 225076
rect 44004 225074 44604 225076
rect 80004 225074 80604 225076
rect 116004 225074 116604 225076
rect 152004 225074 152604 225076
rect 188004 225074 188604 225076
rect 224004 225074 224604 225076
rect 260004 225074 260604 225076
rect 296004 225074 296604 225076
rect 332004 225074 332604 225076
rect 368004 225074 368604 225076
rect 404004 225074 404604 225076
rect 440004 225074 440604 225076
rect 476004 225074 476604 225076
rect 512004 225074 512604 225076
rect 548004 225074 548604 225076
rect 589080 225074 589680 225076
rect -3876 222076 -3276 222078
rect 4404 222076 5004 222078
rect 40404 222076 41004 222078
rect 76404 222076 77004 222078
rect 112404 222076 113004 222078
rect 148404 222076 149004 222078
rect 184404 222076 185004 222078
rect 220404 222076 221004 222078
rect 256404 222076 257004 222078
rect 292404 222076 293004 222078
rect 328404 222076 329004 222078
rect 364404 222076 365004 222078
rect 400404 222076 401004 222078
rect 436404 222076 437004 222078
rect 472404 222076 473004 222078
rect 508404 222076 509004 222078
rect 544404 222076 545004 222078
rect 580404 222076 581004 222078
rect 587200 222076 587800 222078
rect -4816 222054 588740 222076
rect -4816 221818 -3694 222054
rect -3458 221818 4586 222054
rect 4822 221818 40586 222054
rect 40822 221818 76586 222054
rect 76822 221818 112586 222054
rect 112822 221818 148586 222054
rect 148822 221818 184586 222054
rect 184822 221818 220586 222054
rect 220822 221818 256586 222054
rect 256822 221818 292586 222054
rect 292822 221818 328586 222054
rect 328822 221818 364586 222054
rect 364822 221818 400586 222054
rect 400822 221818 436586 222054
rect 436822 221818 472586 222054
rect 472822 221818 508586 222054
rect 508822 221818 544586 222054
rect 544822 221818 580586 222054
rect 580822 221818 587382 222054
rect 587618 221818 588740 222054
rect -4816 221734 588740 221818
rect -4816 221498 -3694 221734
rect -3458 221498 4586 221734
rect 4822 221498 40586 221734
rect 40822 221498 76586 221734
rect 76822 221498 112586 221734
rect 112822 221498 148586 221734
rect 148822 221498 184586 221734
rect 184822 221498 220586 221734
rect 220822 221498 256586 221734
rect 256822 221498 292586 221734
rect 292822 221498 328586 221734
rect 328822 221498 364586 221734
rect 364822 221498 400586 221734
rect 400822 221498 436586 221734
rect 436822 221498 472586 221734
rect 472822 221498 508586 221734
rect 508822 221498 544586 221734
rect 544822 221498 580586 221734
rect 580822 221498 587382 221734
rect 587618 221498 588740 221734
rect -4816 221476 588740 221498
rect -3876 221474 -3276 221476
rect 4404 221474 5004 221476
rect 40404 221474 41004 221476
rect 76404 221474 77004 221476
rect 112404 221474 113004 221476
rect 148404 221474 149004 221476
rect 184404 221474 185004 221476
rect 220404 221474 221004 221476
rect 256404 221474 257004 221476
rect 292404 221474 293004 221476
rect 328404 221474 329004 221476
rect 364404 221474 365004 221476
rect 400404 221474 401004 221476
rect 436404 221474 437004 221476
rect 472404 221474 473004 221476
rect 508404 221474 509004 221476
rect 544404 221474 545004 221476
rect 580404 221474 581004 221476
rect 587200 221474 587800 221476
rect -1996 218476 -1396 218478
rect 804 218476 1404 218478
rect 36804 218476 37404 218478
rect 72804 218476 73404 218478
rect 108804 218476 109404 218478
rect 144804 218476 145404 218478
rect 180804 218476 181404 218478
rect 216804 218476 217404 218478
rect 252804 218476 253404 218478
rect 288804 218476 289404 218478
rect 324804 218476 325404 218478
rect 360804 218476 361404 218478
rect 396804 218476 397404 218478
rect 432804 218476 433404 218478
rect 468804 218476 469404 218478
rect 504804 218476 505404 218478
rect 540804 218476 541404 218478
rect 576804 218476 577404 218478
rect 585320 218476 585920 218478
rect -2936 218454 586860 218476
rect -2936 218218 -1814 218454
rect -1578 218218 986 218454
rect 1222 218218 36986 218454
rect 37222 218218 72986 218454
rect 73222 218218 108986 218454
rect 109222 218218 144986 218454
rect 145222 218218 180986 218454
rect 181222 218218 216986 218454
rect 217222 218218 252986 218454
rect 253222 218218 288986 218454
rect 289222 218218 324986 218454
rect 325222 218218 360986 218454
rect 361222 218218 396986 218454
rect 397222 218218 432986 218454
rect 433222 218218 468986 218454
rect 469222 218218 504986 218454
rect 505222 218218 540986 218454
rect 541222 218218 576986 218454
rect 577222 218218 585502 218454
rect 585738 218218 586860 218454
rect -2936 218134 586860 218218
rect -2936 217898 -1814 218134
rect -1578 217898 986 218134
rect 1222 217898 36986 218134
rect 37222 217898 72986 218134
rect 73222 217898 108986 218134
rect 109222 217898 144986 218134
rect 145222 217898 180986 218134
rect 181222 217898 216986 218134
rect 217222 217898 252986 218134
rect 253222 217898 288986 218134
rect 289222 217898 324986 218134
rect 325222 217898 360986 218134
rect 361222 217898 396986 218134
rect 397222 217898 432986 218134
rect 433222 217898 468986 218134
rect 469222 217898 504986 218134
rect 505222 217898 540986 218134
rect 541222 217898 576986 218134
rect 577222 217898 585502 218134
rect 585738 217898 586860 218134
rect -2936 217876 586860 217898
rect -1996 217874 -1396 217876
rect 804 217874 1404 217876
rect 36804 217874 37404 217876
rect 72804 217874 73404 217876
rect 108804 217874 109404 217876
rect 144804 217874 145404 217876
rect 180804 217874 181404 217876
rect 216804 217874 217404 217876
rect 252804 217874 253404 217876
rect 288804 217874 289404 217876
rect 324804 217874 325404 217876
rect 360804 217874 361404 217876
rect 396804 217874 397404 217876
rect 432804 217874 433404 217876
rect 468804 217874 469404 217876
rect 504804 217874 505404 217876
rect 540804 217874 541404 217876
rect 576804 217874 577404 217876
rect 585320 217874 585920 217876
rect -8576 211276 -7976 211278
rect 29604 211276 30204 211278
rect 65604 211276 66204 211278
rect 101604 211276 102204 211278
rect 137604 211276 138204 211278
rect 173604 211276 174204 211278
rect 209604 211276 210204 211278
rect 245604 211276 246204 211278
rect 281604 211276 282204 211278
rect 317604 211276 318204 211278
rect 353604 211276 354204 211278
rect 389604 211276 390204 211278
rect 425604 211276 426204 211278
rect 461604 211276 462204 211278
rect 497604 211276 498204 211278
rect 533604 211276 534204 211278
rect 569604 211276 570204 211278
rect 591900 211276 592500 211278
rect -8576 211254 592500 211276
rect -8576 211018 -8394 211254
rect -8158 211018 29786 211254
rect 30022 211018 65786 211254
rect 66022 211018 101786 211254
rect 102022 211018 137786 211254
rect 138022 211018 173786 211254
rect 174022 211018 209786 211254
rect 210022 211018 245786 211254
rect 246022 211018 281786 211254
rect 282022 211018 317786 211254
rect 318022 211018 353786 211254
rect 354022 211018 389786 211254
rect 390022 211018 425786 211254
rect 426022 211018 461786 211254
rect 462022 211018 497786 211254
rect 498022 211018 533786 211254
rect 534022 211018 569786 211254
rect 570022 211018 592082 211254
rect 592318 211018 592500 211254
rect -8576 210934 592500 211018
rect -8576 210698 -8394 210934
rect -8158 210698 29786 210934
rect 30022 210698 65786 210934
rect 66022 210698 101786 210934
rect 102022 210698 137786 210934
rect 138022 210698 173786 210934
rect 174022 210698 209786 210934
rect 210022 210698 245786 210934
rect 246022 210698 281786 210934
rect 282022 210698 317786 210934
rect 318022 210698 353786 210934
rect 354022 210698 389786 210934
rect 390022 210698 425786 210934
rect 426022 210698 461786 210934
rect 462022 210698 497786 210934
rect 498022 210698 533786 210934
rect 534022 210698 569786 210934
rect 570022 210698 592082 210934
rect 592318 210698 592500 210934
rect -8576 210676 592500 210698
rect -8576 210674 -7976 210676
rect 29604 210674 30204 210676
rect 65604 210674 66204 210676
rect 101604 210674 102204 210676
rect 137604 210674 138204 210676
rect 173604 210674 174204 210676
rect 209604 210674 210204 210676
rect 245604 210674 246204 210676
rect 281604 210674 282204 210676
rect 317604 210674 318204 210676
rect 353604 210674 354204 210676
rect 389604 210674 390204 210676
rect 425604 210674 426204 210676
rect 461604 210674 462204 210676
rect 497604 210674 498204 210676
rect 533604 210674 534204 210676
rect 569604 210674 570204 210676
rect 591900 210674 592500 210676
rect -6696 207676 -6096 207678
rect 26004 207676 26604 207678
rect 62004 207676 62604 207678
rect 98004 207676 98604 207678
rect 134004 207676 134604 207678
rect 170004 207676 170604 207678
rect 206004 207676 206604 207678
rect 242004 207676 242604 207678
rect 278004 207676 278604 207678
rect 314004 207676 314604 207678
rect 350004 207676 350604 207678
rect 386004 207676 386604 207678
rect 422004 207676 422604 207678
rect 458004 207676 458604 207678
rect 494004 207676 494604 207678
rect 530004 207676 530604 207678
rect 566004 207676 566604 207678
rect 590020 207676 590620 207678
rect -6696 207654 590620 207676
rect -6696 207418 -6514 207654
rect -6278 207418 26186 207654
rect 26422 207418 62186 207654
rect 62422 207418 98186 207654
rect 98422 207418 134186 207654
rect 134422 207418 170186 207654
rect 170422 207418 206186 207654
rect 206422 207418 242186 207654
rect 242422 207418 278186 207654
rect 278422 207418 314186 207654
rect 314422 207418 350186 207654
rect 350422 207418 386186 207654
rect 386422 207418 422186 207654
rect 422422 207418 458186 207654
rect 458422 207418 494186 207654
rect 494422 207418 530186 207654
rect 530422 207418 566186 207654
rect 566422 207418 590202 207654
rect 590438 207418 590620 207654
rect -6696 207334 590620 207418
rect -6696 207098 -6514 207334
rect -6278 207098 26186 207334
rect 26422 207098 62186 207334
rect 62422 207098 98186 207334
rect 98422 207098 134186 207334
rect 134422 207098 170186 207334
rect 170422 207098 206186 207334
rect 206422 207098 242186 207334
rect 242422 207098 278186 207334
rect 278422 207098 314186 207334
rect 314422 207098 350186 207334
rect 350422 207098 386186 207334
rect 386422 207098 422186 207334
rect 422422 207098 458186 207334
rect 458422 207098 494186 207334
rect 494422 207098 530186 207334
rect 530422 207098 566186 207334
rect 566422 207098 590202 207334
rect 590438 207098 590620 207334
rect -6696 207076 590620 207098
rect -6696 207074 -6096 207076
rect 26004 207074 26604 207076
rect 62004 207074 62604 207076
rect 98004 207074 98604 207076
rect 134004 207074 134604 207076
rect 170004 207074 170604 207076
rect 206004 207074 206604 207076
rect 242004 207074 242604 207076
rect 278004 207074 278604 207076
rect 314004 207074 314604 207076
rect 350004 207074 350604 207076
rect 386004 207074 386604 207076
rect 422004 207074 422604 207076
rect 458004 207074 458604 207076
rect 494004 207074 494604 207076
rect 530004 207074 530604 207076
rect 566004 207074 566604 207076
rect 590020 207074 590620 207076
rect -4816 204076 -4216 204078
rect 22404 204076 23004 204078
rect 58404 204076 59004 204078
rect 94404 204076 95004 204078
rect 130404 204076 131004 204078
rect 166404 204076 167004 204078
rect 202404 204076 203004 204078
rect 238404 204076 239004 204078
rect 274404 204076 275004 204078
rect 382404 204076 383004 204078
rect 526404 204076 527004 204078
rect 562404 204076 563004 204078
rect 588140 204076 588740 204078
rect -4816 204054 588740 204076
rect -4816 203818 -4634 204054
rect -4398 203818 22586 204054
rect 22822 203818 58586 204054
rect 58822 203818 94586 204054
rect 94822 203818 130586 204054
rect 130822 203818 166586 204054
rect 166822 203818 202586 204054
rect 202822 203818 238586 204054
rect 238822 203818 274586 204054
rect 274822 203818 382586 204054
rect 382822 203818 526586 204054
rect 526822 203818 562586 204054
rect 562822 203818 588322 204054
rect 588558 203818 588740 204054
rect -4816 203734 588740 203818
rect -4816 203498 -4634 203734
rect -4398 203498 22586 203734
rect 22822 203498 58586 203734
rect 58822 203498 94586 203734
rect 94822 203498 130586 203734
rect 130822 203498 166586 203734
rect 166822 203498 202586 203734
rect 202822 203498 238586 203734
rect 238822 203498 274586 203734
rect 274822 203498 382586 203734
rect 382822 203498 526586 203734
rect 526822 203498 562586 203734
rect 562822 203498 588322 203734
rect 588558 203498 588740 203734
rect -4816 203476 588740 203498
rect -4816 203474 -4216 203476
rect 22404 203474 23004 203476
rect 58404 203474 59004 203476
rect 94404 203474 95004 203476
rect 130404 203474 131004 203476
rect 166404 203474 167004 203476
rect 202404 203474 203004 203476
rect 238404 203474 239004 203476
rect 274404 203474 275004 203476
rect 382404 203474 383004 203476
rect 526404 203474 527004 203476
rect 562404 203474 563004 203476
rect 588140 203474 588740 203476
rect -2936 200476 -2336 200478
rect 18804 200476 19404 200478
rect 54804 200476 55404 200478
rect 90804 200476 91404 200478
rect 126804 200476 127404 200478
rect 162804 200476 163404 200478
rect 198804 200476 199404 200478
rect 234804 200476 235404 200478
rect 270804 200476 271404 200478
rect 414804 200476 415404 200478
rect 522804 200476 523404 200478
rect 558804 200476 559404 200478
rect 586260 200476 586860 200478
rect -2936 200454 586860 200476
rect -2936 200218 -2754 200454
rect -2518 200218 18986 200454
rect 19222 200218 54986 200454
rect 55222 200218 90986 200454
rect 91222 200218 126986 200454
rect 127222 200218 162986 200454
rect 163222 200218 198986 200454
rect 199222 200218 234986 200454
rect 235222 200218 270986 200454
rect 271222 200218 414986 200454
rect 415222 200218 522986 200454
rect 523222 200218 558986 200454
rect 559222 200218 586442 200454
rect 586678 200218 586860 200454
rect -2936 200134 586860 200218
rect -2936 199898 -2754 200134
rect -2518 199898 18986 200134
rect 19222 199898 54986 200134
rect 55222 199898 90986 200134
rect 91222 199898 126986 200134
rect 127222 199898 162986 200134
rect 163222 199898 198986 200134
rect 199222 199898 234986 200134
rect 235222 199898 270986 200134
rect 271222 199898 414986 200134
rect 415222 199898 522986 200134
rect 523222 199898 558986 200134
rect 559222 199898 586442 200134
rect 586678 199898 586860 200134
rect -2936 199876 586860 199898
rect -2936 199874 -2336 199876
rect 18804 199874 19404 199876
rect 54804 199874 55404 199876
rect 90804 199874 91404 199876
rect 126804 199874 127404 199876
rect 162804 199874 163404 199876
rect 198804 199874 199404 199876
rect 234804 199874 235404 199876
rect 270804 199874 271404 199876
rect 414804 199874 415404 199876
rect 522804 199874 523404 199876
rect 558804 199874 559404 199876
rect 586260 199874 586860 199876
rect -7636 193276 -7036 193278
rect 11604 193276 12204 193278
rect 47604 193276 48204 193278
rect 83604 193276 84204 193278
rect 119604 193276 120204 193278
rect 155604 193276 156204 193278
rect 191604 193276 192204 193278
rect 227604 193276 228204 193278
rect 263604 193276 264204 193278
rect 407604 193276 408204 193278
rect 515604 193276 516204 193278
rect 551604 193276 552204 193278
rect 590960 193276 591560 193278
rect -8576 193254 592500 193276
rect -8576 193018 -7454 193254
rect -7218 193018 11786 193254
rect 12022 193018 47786 193254
rect 48022 193018 83786 193254
rect 84022 193018 119786 193254
rect 120022 193018 155786 193254
rect 156022 193018 191786 193254
rect 192022 193018 227786 193254
rect 228022 193018 263786 193254
rect 264022 193018 407786 193254
rect 408022 193018 515786 193254
rect 516022 193018 551786 193254
rect 552022 193018 591142 193254
rect 591378 193018 592500 193254
rect -8576 192934 592500 193018
rect -8576 192698 -7454 192934
rect -7218 192698 11786 192934
rect 12022 192698 47786 192934
rect 48022 192698 83786 192934
rect 84022 192698 119786 192934
rect 120022 192698 155786 192934
rect 156022 192698 191786 192934
rect 192022 192698 227786 192934
rect 228022 192698 263786 192934
rect 264022 192698 407786 192934
rect 408022 192698 515786 192934
rect 516022 192698 551786 192934
rect 552022 192698 591142 192934
rect 591378 192698 592500 192934
rect -8576 192676 592500 192698
rect -7636 192674 -7036 192676
rect 11604 192674 12204 192676
rect 47604 192674 48204 192676
rect 83604 192674 84204 192676
rect 119604 192674 120204 192676
rect 155604 192674 156204 192676
rect 191604 192674 192204 192676
rect 227604 192674 228204 192676
rect 263604 192674 264204 192676
rect 407604 192674 408204 192676
rect 515604 192674 516204 192676
rect 551604 192674 552204 192676
rect 590960 192674 591560 192676
rect -5756 189676 -5156 189678
rect 8004 189676 8604 189678
rect 44004 189676 44604 189678
rect 80004 189676 80604 189678
rect 116004 189676 116604 189678
rect 152004 189676 152604 189678
rect 188004 189676 188604 189678
rect 224004 189676 224604 189678
rect 260004 189676 260604 189678
rect 296004 189676 296604 189678
rect 404004 189676 404604 189678
rect 512004 189676 512604 189678
rect 548004 189676 548604 189678
rect 589080 189676 589680 189678
rect -6696 189654 590620 189676
rect -6696 189418 -5574 189654
rect -5338 189418 8186 189654
rect 8422 189418 44186 189654
rect 44422 189418 80186 189654
rect 80422 189418 116186 189654
rect 116422 189418 152186 189654
rect 152422 189418 188186 189654
rect 188422 189418 224186 189654
rect 224422 189418 260186 189654
rect 260422 189418 296186 189654
rect 296422 189418 404186 189654
rect 404422 189418 512186 189654
rect 512422 189418 548186 189654
rect 548422 189418 589262 189654
rect 589498 189418 590620 189654
rect -6696 189334 590620 189418
rect -6696 189098 -5574 189334
rect -5338 189098 8186 189334
rect 8422 189098 44186 189334
rect 44422 189098 80186 189334
rect 80422 189098 116186 189334
rect 116422 189098 152186 189334
rect 152422 189098 188186 189334
rect 188422 189098 224186 189334
rect 224422 189098 260186 189334
rect 260422 189098 296186 189334
rect 296422 189098 404186 189334
rect 404422 189098 512186 189334
rect 512422 189098 548186 189334
rect 548422 189098 589262 189334
rect 589498 189098 590620 189334
rect -6696 189076 590620 189098
rect -5756 189074 -5156 189076
rect 8004 189074 8604 189076
rect 44004 189074 44604 189076
rect 80004 189074 80604 189076
rect 116004 189074 116604 189076
rect 152004 189074 152604 189076
rect 188004 189074 188604 189076
rect 224004 189074 224604 189076
rect 260004 189074 260604 189076
rect 296004 189074 296604 189076
rect 404004 189074 404604 189076
rect 512004 189074 512604 189076
rect 548004 189074 548604 189076
rect 589080 189074 589680 189076
rect -3876 186076 -3276 186078
rect 4404 186076 5004 186078
rect 40404 186076 41004 186078
rect 76404 186076 77004 186078
rect 112404 186076 113004 186078
rect 148404 186076 149004 186078
rect 184404 186076 185004 186078
rect 220404 186076 221004 186078
rect 256404 186076 257004 186078
rect 292404 186076 293004 186078
rect 400404 186076 401004 186078
rect 508404 186076 509004 186078
rect 544404 186076 545004 186078
rect 580404 186076 581004 186078
rect 587200 186076 587800 186078
rect -4816 186054 588740 186076
rect -4816 185818 -3694 186054
rect -3458 185818 4586 186054
rect 4822 185818 40586 186054
rect 40822 185818 76586 186054
rect 76822 185818 112586 186054
rect 112822 185818 148586 186054
rect 148822 185818 184586 186054
rect 184822 185818 220586 186054
rect 220822 185818 256586 186054
rect 256822 185818 292586 186054
rect 292822 185818 400586 186054
rect 400822 185818 508586 186054
rect 508822 185818 544586 186054
rect 544822 185818 580586 186054
rect 580822 185818 587382 186054
rect 587618 185818 588740 186054
rect -4816 185734 588740 185818
rect -4816 185498 -3694 185734
rect -3458 185498 4586 185734
rect 4822 185498 40586 185734
rect 40822 185498 76586 185734
rect 76822 185498 112586 185734
rect 112822 185498 148586 185734
rect 148822 185498 184586 185734
rect 184822 185498 220586 185734
rect 220822 185498 256586 185734
rect 256822 185498 292586 185734
rect 292822 185498 400586 185734
rect 400822 185498 508586 185734
rect 508822 185498 544586 185734
rect 544822 185498 580586 185734
rect 580822 185498 587382 185734
rect 587618 185498 588740 185734
rect -4816 185476 588740 185498
rect -3876 185474 -3276 185476
rect 4404 185474 5004 185476
rect 40404 185474 41004 185476
rect 76404 185474 77004 185476
rect 112404 185474 113004 185476
rect 148404 185474 149004 185476
rect 184404 185474 185004 185476
rect 220404 185474 221004 185476
rect 256404 185474 257004 185476
rect 292404 185474 293004 185476
rect 400404 185474 401004 185476
rect 508404 185474 509004 185476
rect 544404 185474 545004 185476
rect 580404 185474 581004 185476
rect 587200 185474 587800 185476
rect -1996 182476 -1396 182478
rect 804 182476 1404 182478
rect 36804 182476 37404 182478
rect 72804 182476 73404 182478
rect 108804 182476 109404 182478
rect 144804 182476 145404 182478
rect 180804 182476 181404 182478
rect 216804 182476 217404 182478
rect 252804 182476 253404 182478
rect 288804 182476 289404 182478
rect 300482 182476 300802 182478
rect 396804 182476 397404 182478
rect 420482 182476 420802 182478
rect 504804 182476 505404 182478
rect 540804 182476 541404 182478
rect 576804 182476 577404 182478
rect 585320 182476 585920 182478
rect -2936 182454 586860 182476
rect -2936 182218 -1814 182454
rect -1578 182218 986 182454
rect 1222 182218 36986 182454
rect 37222 182218 72986 182454
rect 73222 182218 108986 182454
rect 109222 182218 144986 182454
rect 145222 182218 180986 182454
rect 181222 182218 216986 182454
rect 217222 182218 252986 182454
rect 253222 182218 288986 182454
rect 289222 182218 300524 182454
rect 300760 182218 396986 182454
rect 397222 182218 420524 182454
rect 420760 182218 504986 182454
rect 505222 182218 540986 182454
rect 541222 182218 576986 182454
rect 577222 182218 585502 182454
rect 585738 182218 586860 182454
rect -2936 182134 586860 182218
rect -2936 181898 -1814 182134
rect -1578 181898 986 182134
rect 1222 181898 36986 182134
rect 37222 181898 72986 182134
rect 73222 181898 108986 182134
rect 109222 181898 144986 182134
rect 145222 181898 180986 182134
rect 181222 181898 216986 182134
rect 217222 181898 252986 182134
rect 253222 181898 288986 182134
rect 289222 181898 300524 182134
rect 300760 181898 396986 182134
rect 397222 181898 420524 182134
rect 420760 181898 504986 182134
rect 505222 181898 540986 182134
rect 541222 181898 576986 182134
rect 577222 181898 585502 182134
rect 585738 181898 586860 182134
rect -2936 181876 586860 181898
rect -1996 181874 -1396 181876
rect 804 181874 1404 181876
rect 36804 181874 37404 181876
rect 72804 181874 73404 181876
rect 108804 181874 109404 181876
rect 144804 181874 145404 181876
rect 180804 181874 181404 181876
rect 216804 181874 217404 181876
rect 252804 181874 253404 181876
rect 288804 181874 289404 181876
rect 300482 181874 300802 181876
rect 396804 181874 397404 181876
rect 420482 181874 420802 181876
rect 504804 181874 505404 181876
rect 540804 181874 541404 181876
rect 576804 181874 577404 181876
rect 585320 181874 585920 181876
rect -8576 175276 -7976 175278
rect 29604 175276 30204 175278
rect 65604 175276 66204 175278
rect 101604 175276 102204 175278
rect 137604 175276 138204 175278
rect 173604 175276 174204 175278
rect 209604 175276 210204 175278
rect 245604 175276 246204 175278
rect 281604 175276 282204 175278
rect 389604 175276 390204 175278
rect 533604 175276 534204 175278
rect 569604 175276 570204 175278
rect 591900 175276 592500 175278
rect -8576 175254 592500 175276
rect -8576 175018 -8394 175254
rect -8158 175018 29786 175254
rect 30022 175018 65786 175254
rect 66022 175018 101786 175254
rect 102022 175018 137786 175254
rect 138022 175018 173786 175254
rect 174022 175018 209786 175254
rect 210022 175018 245786 175254
rect 246022 175018 281786 175254
rect 282022 175018 389786 175254
rect 390022 175018 533786 175254
rect 534022 175018 569786 175254
rect 570022 175018 592082 175254
rect 592318 175018 592500 175254
rect -8576 174934 592500 175018
rect -8576 174698 -8394 174934
rect -8158 174698 29786 174934
rect 30022 174698 65786 174934
rect 66022 174698 101786 174934
rect 102022 174698 137786 174934
rect 138022 174698 173786 174934
rect 174022 174698 209786 174934
rect 210022 174698 245786 174934
rect 246022 174698 281786 174934
rect 282022 174698 389786 174934
rect 390022 174698 533786 174934
rect 534022 174698 569786 174934
rect 570022 174698 592082 174934
rect 592318 174698 592500 174934
rect -8576 174676 592500 174698
rect -8576 174674 -7976 174676
rect 29604 174674 30204 174676
rect 65604 174674 66204 174676
rect 101604 174674 102204 174676
rect 137604 174674 138204 174676
rect 173604 174674 174204 174676
rect 209604 174674 210204 174676
rect 245604 174674 246204 174676
rect 281604 174674 282204 174676
rect 389604 174674 390204 174676
rect 533604 174674 534204 174676
rect 569604 174674 570204 174676
rect 591900 174674 592500 174676
rect -6696 171676 -6096 171678
rect 26004 171676 26604 171678
rect 62004 171676 62604 171678
rect 98004 171676 98604 171678
rect 134004 171676 134604 171678
rect 170004 171676 170604 171678
rect 206004 171676 206604 171678
rect 242004 171676 242604 171678
rect 278004 171676 278604 171678
rect 386004 171676 386604 171678
rect 530004 171676 530604 171678
rect 566004 171676 566604 171678
rect 590020 171676 590620 171678
rect -6696 171654 590620 171676
rect -6696 171418 -6514 171654
rect -6278 171418 26186 171654
rect 26422 171418 62186 171654
rect 62422 171418 98186 171654
rect 98422 171418 134186 171654
rect 134422 171418 170186 171654
rect 170422 171418 206186 171654
rect 206422 171418 242186 171654
rect 242422 171418 278186 171654
rect 278422 171418 386186 171654
rect 386422 171418 530186 171654
rect 530422 171418 566186 171654
rect 566422 171418 590202 171654
rect 590438 171418 590620 171654
rect -6696 171334 590620 171418
rect -6696 171098 -6514 171334
rect -6278 171098 26186 171334
rect 26422 171098 62186 171334
rect 62422 171098 98186 171334
rect 98422 171098 134186 171334
rect 134422 171098 170186 171334
rect 170422 171098 206186 171334
rect 206422 171098 242186 171334
rect 242422 171098 278186 171334
rect 278422 171098 386186 171334
rect 386422 171098 530186 171334
rect 530422 171098 566186 171334
rect 566422 171098 590202 171334
rect 590438 171098 590620 171334
rect -6696 171076 590620 171098
rect -6696 171074 -6096 171076
rect 26004 171074 26604 171076
rect 62004 171074 62604 171076
rect 98004 171074 98604 171076
rect 134004 171074 134604 171076
rect 170004 171074 170604 171076
rect 206004 171074 206604 171076
rect 242004 171074 242604 171076
rect 278004 171074 278604 171076
rect 386004 171074 386604 171076
rect 530004 171074 530604 171076
rect 566004 171074 566604 171076
rect 590020 171074 590620 171076
rect -4816 168076 -4216 168078
rect 22404 168076 23004 168078
rect 58404 168076 59004 168078
rect 94404 168076 95004 168078
rect 130404 168076 131004 168078
rect 166404 168076 167004 168078
rect 202404 168076 203004 168078
rect 238404 168076 239004 168078
rect 274404 168076 275004 168078
rect 382404 168076 383004 168078
rect 526404 168076 527004 168078
rect 562404 168076 563004 168078
rect 588140 168076 588740 168078
rect -4816 168054 588740 168076
rect -4816 167818 -4634 168054
rect -4398 167818 22586 168054
rect 22822 167818 58586 168054
rect 58822 167818 94586 168054
rect 94822 167818 130586 168054
rect 130822 167818 166586 168054
rect 166822 167818 202586 168054
rect 202822 167818 238586 168054
rect 238822 167818 274586 168054
rect 274822 167818 382586 168054
rect 382822 167818 526586 168054
rect 526822 167818 562586 168054
rect 562822 167818 588322 168054
rect 588558 167818 588740 168054
rect -4816 167734 588740 167818
rect -4816 167498 -4634 167734
rect -4398 167498 22586 167734
rect 22822 167498 58586 167734
rect 58822 167498 94586 167734
rect 94822 167498 130586 167734
rect 130822 167498 166586 167734
rect 166822 167498 202586 167734
rect 202822 167498 238586 167734
rect 238822 167498 274586 167734
rect 274822 167498 382586 167734
rect 382822 167498 526586 167734
rect 526822 167498 562586 167734
rect 562822 167498 588322 167734
rect 588558 167498 588740 167734
rect -4816 167476 588740 167498
rect -4816 167474 -4216 167476
rect 22404 167474 23004 167476
rect 58404 167474 59004 167476
rect 94404 167474 95004 167476
rect 130404 167474 131004 167476
rect 166404 167474 167004 167476
rect 202404 167474 203004 167476
rect 238404 167474 239004 167476
rect 274404 167474 275004 167476
rect 382404 167474 383004 167476
rect 526404 167474 527004 167476
rect 562404 167474 563004 167476
rect 588140 167474 588740 167476
rect -2936 164476 -2336 164478
rect 18804 164476 19404 164478
rect 54804 164476 55404 164478
rect 90804 164476 91404 164478
rect 126804 164476 127404 164478
rect 162804 164476 163404 164478
rect 198804 164476 199404 164478
rect 234804 164476 235404 164478
rect 270804 164476 271404 164478
rect 300034 164476 300358 164478
rect 414804 164476 415404 164478
rect 420034 164476 420358 164478
rect 522804 164476 523404 164478
rect 558804 164476 559404 164478
rect 586260 164476 586860 164478
rect -2936 164454 586860 164476
rect -2936 164218 -2754 164454
rect -2518 164218 18986 164454
rect 19222 164218 54986 164454
rect 55222 164218 90986 164454
rect 91222 164218 126986 164454
rect 127222 164218 162986 164454
rect 163222 164218 198986 164454
rect 199222 164218 234986 164454
rect 235222 164218 270986 164454
rect 271222 164218 300078 164454
rect 300314 164218 414986 164454
rect 415222 164218 420078 164454
rect 420314 164218 522986 164454
rect 523222 164218 558986 164454
rect 559222 164218 586442 164454
rect 586678 164218 586860 164454
rect -2936 164134 586860 164218
rect -2936 163898 -2754 164134
rect -2518 163898 18986 164134
rect 19222 163898 54986 164134
rect 55222 163898 90986 164134
rect 91222 163898 126986 164134
rect 127222 163898 162986 164134
rect 163222 163898 198986 164134
rect 199222 163898 234986 164134
rect 235222 163898 270986 164134
rect 271222 163898 300078 164134
rect 300314 163898 414986 164134
rect 415222 163898 420078 164134
rect 420314 163898 522986 164134
rect 523222 163898 558986 164134
rect 559222 163898 586442 164134
rect 586678 163898 586860 164134
rect -2936 163876 586860 163898
rect -2936 163874 -2336 163876
rect 18804 163874 19404 163876
rect 54804 163874 55404 163876
rect 90804 163874 91404 163876
rect 126804 163874 127404 163876
rect 162804 163874 163404 163876
rect 198804 163874 199404 163876
rect 234804 163874 235404 163876
rect 270804 163874 271404 163876
rect 300034 163874 300358 163876
rect 414804 163874 415404 163876
rect 420034 163874 420358 163876
rect 522804 163874 523404 163876
rect 558804 163874 559404 163876
rect 586260 163874 586860 163876
rect -7636 157276 -7036 157278
rect 11604 157276 12204 157278
rect 47604 157276 48204 157278
rect 83604 157276 84204 157278
rect 119604 157276 120204 157278
rect 155604 157276 156204 157278
rect 191604 157276 192204 157278
rect 227604 157276 228204 157278
rect 263604 157276 264204 157278
rect 407604 157276 408204 157278
rect 515604 157276 516204 157278
rect 551604 157276 552204 157278
rect 590960 157276 591560 157278
rect -8576 157254 592500 157276
rect -8576 157018 -7454 157254
rect -7218 157018 11786 157254
rect 12022 157018 47786 157254
rect 48022 157018 83786 157254
rect 84022 157018 119786 157254
rect 120022 157018 155786 157254
rect 156022 157018 191786 157254
rect 192022 157018 227786 157254
rect 228022 157018 263786 157254
rect 264022 157018 407786 157254
rect 408022 157018 515786 157254
rect 516022 157018 551786 157254
rect 552022 157018 591142 157254
rect 591378 157018 592500 157254
rect -8576 156934 592500 157018
rect -8576 156698 -7454 156934
rect -7218 156698 11786 156934
rect 12022 156698 47786 156934
rect 48022 156698 83786 156934
rect 84022 156698 119786 156934
rect 120022 156698 155786 156934
rect 156022 156698 191786 156934
rect 192022 156698 227786 156934
rect 228022 156698 263786 156934
rect 264022 156698 407786 156934
rect 408022 156698 515786 156934
rect 516022 156698 551786 156934
rect 552022 156698 591142 156934
rect 591378 156698 592500 156934
rect -8576 156676 592500 156698
rect -7636 156674 -7036 156676
rect 11604 156674 12204 156676
rect 47604 156674 48204 156676
rect 83604 156674 84204 156676
rect 119604 156674 120204 156676
rect 155604 156674 156204 156676
rect 191604 156674 192204 156676
rect 227604 156674 228204 156676
rect 263604 156674 264204 156676
rect 407604 156674 408204 156676
rect 515604 156674 516204 156676
rect 551604 156674 552204 156676
rect 590960 156674 591560 156676
rect -5756 153676 -5156 153678
rect 8004 153676 8604 153678
rect 44004 153676 44604 153678
rect 80004 153676 80604 153678
rect 116004 153676 116604 153678
rect 152004 153676 152604 153678
rect 188004 153676 188604 153678
rect 224004 153676 224604 153678
rect 260004 153676 260604 153678
rect 296004 153676 296604 153678
rect 404004 153676 404604 153678
rect 512004 153676 512604 153678
rect 548004 153676 548604 153678
rect 589080 153676 589680 153678
rect -6696 153654 590620 153676
rect -6696 153418 -5574 153654
rect -5338 153418 8186 153654
rect 8422 153418 44186 153654
rect 44422 153418 80186 153654
rect 80422 153418 116186 153654
rect 116422 153418 152186 153654
rect 152422 153418 188186 153654
rect 188422 153418 224186 153654
rect 224422 153418 260186 153654
rect 260422 153418 296186 153654
rect 296422 153418 404186 153654
rect 404422 153418 512186 153654
rect 512422 153418 548186 153654
rect 548422 153418 589262 153654
rect 589498 153418 590620 153654
rect -6696 153334 590620 153418
rect -6696 153098 -5574 153334
rect -5338 153098 8186 153334
rect 8422 153098 44186 153334
rect 44422 153098 80186 153334
rect 80422 153098 116186 153334
rect 116422 153098 152186 153334
rect 152422 153098 188186 153334
rect 188422 153098 224186 153334
rect 224422 153098 260186 153334
rect 260422 153098 296186 153334
rect 296422 153098 404186 153334
rect 404422 153098 512186 153334
rect 512422 153098 548186 153334
rect 548422 153098 589262 153334
rect 589498 153098 590620 153334
rect -6696 153076 590620 153098
rect -5756 153074 -5156 153076
rect 8004 153074 8604 153076
rect 44004 153074 44604 153076
rect 80004 153074 80604 153076
rect 116004 153074 116604 153076
rect 152004 153074 152604 153076
rect 188004 153074 188604 153076
rect 224004 153074 224604 153076
rect 260004 153074 260604 153076
rect 296004 153074 296604 153076
rect 404004 153074 404604 153076
rect 512004 153074 512604 153076
rect 548004 153074 548604 153076
rect 589080 153074 589680 153076
rect -3876 150076 -3276 150078
rect 4404 150076 5004 150078
rect 40404 150076 41004 150078
rect 76404 150076 77004 150078
rect 112404 150076 113004 150078
rect 148404 150076 149004 150078
rect 184404 150076 185004 150078
rect 220404 150076 221004 150078
rect 256404 150076 257004 150078
rect 292404 150076 293004 150078
rect 400404 150076 401004 150078
rect 508404 150076 509004 150078
rect 544404 150076 545004 150078
rect 580404 150076 581004 150078
rect 587200 150076 587800 150078
rect -4816 150054 588740 150076
rect -4816 149818 -3694 150054
rect -3458 149818 4586 150054
rect 4822 149818 40586 150054
rect 40822 149818 76586 150054
rect 76822 149818 112586 150054
rect 112822 149818 148586 150054
rect 148822 149818 184586 150054
rect 184822 149818 220586 150054
rect 220822 149818 256586 150054
rect 256822 149818 292586 150054
rect 292822 149818 400586 150054
rect 400822 149818 508586 150054
rect 508822 149818 544586 150054
rect 544822 149818 580586 150054
rect 580822 149818 587382 150054
rect 587618 149818 588740 150054
rect -4816 149734 588740 149818
rect -4816 149498 -3694 149734
rect -3458 149498 4586 149734
rect 4822 149498 40586 149734
rect 40822 149498 76586 149734
rect 76822 149498 112586 149734
rect 112822 149498 148586 149734
rect 148822 149498 184586 149734
rect 184822 149498 220586 149734
rect 220822 149498 256586 149734
rect 256822 149498 292586 149734
rect 292822 149498 400586 149734
rect 400822 149498 508586 149734
rect 508822 149498 544586 149734
rect 544822 149498 580586 149734
rect 580822 149498 587382 149734
rect 587618 149498 588740 149734
rect -4816 149476 588740 149498
rect -3876 149474 -3276 149476
rect 4404 149474 5004 149476
rect 40404 149474 41004 149476
rect 76404 149474 77004 149476
rect 112404 149474 113004 149476
rect 148404 149474 149004 149476
rect 184404 149474 185004 149476
rect 220404 149474 221004 149476
rect 256404 149474 257004 149476
rect 292404 149474 293004 149476
rect 400404 149474 401004 149476
rect 508404 149474 509004 149476
rect 544404 149474 545004 149476
rect 580404 149474 581004 149476
rect 587200 149474 587800 149476
rect -1996 146476 -1396 146478
rect 804 146476 1404 146478
rect 36804 146476 37404 146478
rect 72804 146476 73404 146478
rect 108804 146476 109404 146478
rect 144804 146476 145404 146478
rect 180804 146476 181404 146478
rect 216804 146476 217404 146478
rect 252804 146476 253404 146478
rect 288804 146476 289404 146478
rect 300482 146476 300802 146478
rect 396804 146476 397404 146478
rect 420482 146476 420802 146478
rect 504804 146476 505404 146478
rect 540804 146476 541404 146478
rect 576804 146476 577404 146478
rect 585320 146476 585920 146478
rect -2936 146454 586860 146476
rect -2936 146218 -1814 146454
rect -1578 146218 986 146454
rect 1222 146218 36986 146454
rect 37222 146218 72986 146454
rect 73222 146218 108986 146454
rect 109222 146218 144986 146454
rect 145222 146218 180986 146454
rect 181222 146218 216986 146454
rect 217222 146218 252986 146454
rect 253222 146218 288986 146454
rect 289222 146218 300524 146454
rect 300760 146218 396986 146454
rect 397222 146218 420524 146454
rect 420760 146218 504986 146454
rect 505222 146218 540986 146454
rect 541222 146218 576986 146454
rect 577222 146218 585502 146454
rect 585738 146218 586860 146454
rect -2936 146134 586860 146218
rect -2936 145898 -1814 146134
rect -1578 145898 986 146134
rect 1222 145898 36986 146134
rect 37222 145898 72986 146134
rect 73222 145898 108986 146134
rect 109222 145898 144986 146134
rect 145222 145898 180986 146134
rect 181222 145898 216986 146134
rect 217222 145898 252986 146134
rect 253222 145898 288986 146134
rect 289222 145898 300524 146134
rect 300760 145898 396986 146134
rect 397222 145898 420524 146134
rect 420760 145898 504986 146134
rect 505222 145898 540986 146134
rect 541222 145898 576986 146134
rect 577222 145898 585502 146134
rect 585738 145898 586860 146134
rect -2936 145876 586860 145898
rect -1996 145874 -1396 145876
rect 804 145874 1404 145876
rect 36804 145874 37404 145876
rect 72804 145874 73404 145876
rect 108804 145874 109404 145876
rect 144804 145874 145404 145876
rect 180804 145874 181404 145876
rect 216804 145874 217404 145876
rect 252804 145874 253404 145876
rect 288804 145874 289404 145876
rect 300482 145874 300802 145876
rect 396804 145874 397404 145876
rect 420482 145874 420802 145876
rect 504804 145874 505404 145876
rect 540804 145874 541404 145876
rect 576804 145874 577404 145876
rect 585320 145874 585920 145876
rect -8576 139276 -7976 139278
rect 29604 139276 30204 139278
rect 65604 139276 66204 139278
rect 101604 139276 102204 139278
rect 137604 139276 138204 139278
rect 173604 139276 174204 139278
rect 209604 139276 210204 139278
rect 245604 139276 246204 139278
rect 281604 139276 282204 139278
rect 389604 139276 390204 139278
rect 533604 139276 534204 139278
rect 569604 139276 570204 139278
rect 591900 139276 592500 139278
rect -8576 139254 592500 139276
rect -8576 139018 -8394 139254
rect -8158 139018 29786 139254
rect 30022 139018 65786 139254
rect 66022 139018 101786 139254
rect 102022 139018 137786 139254
rect 138022 139018 173786 139254
rect 174022 139018 209786 139254
rect 210022 139018 245786 139254
rect 246022 139018 281786 139254
rect 282022 139018 389786 139254
rect 390022 139018 533786 139254
rect 534022 139018 569786 139254
rect 570022 139018 592082 139254
rect 592318 139018 592500 139254
rect -8576 138934 592500 139018
rect -8576 138698 -8394 138934
rect -8158 138698 29786 138934
rect 30022 138698 65786 138934
rect 66022 138698 101786 138934
rect 102022 138698 137786 138934
rect 138022 138698 173786 138934
rect 174022 138698 209786 138934
rect 210022 138698 245786 138934
rect 246022 138698 281786 138934
rect 282022 138698 389786 138934
rect 390022 138698 533786 138934
rect 534022 138698 569786 138934
rect 570022 138698 592082 138934
rect 592318 138698 592500 138934
rect -8576 138676 592500 138698
rect -8576 138674 -7976 138676
rect 29604 138674 30204 138676
rect 65604 138674 66204 138676
rect 101604 138674 102204 138676
rect 137604 138674 138204 138676
rect 173604 138674 174204 138676
rect 209604 138674 210204 138676
rect 245604 138674 246204 138676
rect 281604 138674 282204 138676
rect 389604 138674 390204 138676
rect 533604 138674 534204 138676
rect 569604 138674 570204 138676
rect 591900 138674 592500 138676
rect -6696 135676 -6096 135678
rect 26004 135676 26604 135678
rect 62004 135676 62604 135678
rect 98004 135676 98604 135678
rect 134004 135676 134604 135678
rect 170004 135676 170604 135678
rect 206004 135676 206604 135678
rect 242004 135676 242604 135678
rect 278004 135676 278604 135678
rect 386004 135676 386604 135678
rect 530004 135676 530604 135678
rect 566004 135676 566604 135678
rect 590020 135676 590620 135678
rect -6696 135654 590620 135676
rect -6696 135418 -6514 135654
rect -6278 135418 26186 135654
rect 26422 135418 62186 135654
rect 62422 135418 98186 135654
rect 98422 135418 134186 135654
rect 134422 135418 170186 135654
rect 170422 135418 206186 135654
rect 206422 135418 242186 135654
rect 242422 135418 278186 135654
rect 278422 135418 386186 135654
rect 386422 135418 530186 135654
rect 530422 135418 566186 135654
rect 566422 135418 590202 135654
rect 590438 135418 590620 135654
rect -6696 135334 590620 135418
rect -6696 135098 -6514 135334
rect -6278 135098 26186 135334
rect 26422 135098 62186 135334
rect 62422 135098 98186 135334
rect 98422 135098 134186 135334
rect 134422 135098 170186 135334
rect 170422 135098 206186 135334
rect 206422 135098 242186 135334
rect 242422 135098 278186 135334
rect 278422 135098 386186 135334
rect 386422 135098 530186 135334
rect 530422 135098 566186 135334
rect 566422 135098 590202 135334
rect 590438 135098 590620 135334
rect -6696 135076 590620 135098
rect -6696 135074 -6096 135076
rect 26004 135074 26604 135076
rect 62004 135074 62604 135076
rect 98004 135074 98604 135076
rect 134004 135074 134604 135076
rect 170004 135074 170604 135076
rect 206004 135074 206604 135076
rect 242004 135074 242604 135076
rect 278004 135074 278604 135076
rect 386004 135074 386604 135076
rect 530004 135074 530604 135076
rect 566004 135074 566604 135076
rect 590020 135074 590620 135076
rect -4816 132076 -4216 132078
rect 22404 132076 23004 132078
rect 58404 132076 59004 132078
rect 94404 132076 95004 132078
rect 130404 132076 131004 132078
rect 166404 132076 167004 132078
rect 202404 132076 203004 132078
rect 238404 132076 239004 132078
rect 274404 132076 275004 132078
rect 382404 132076 383004 132078
rect 526404 132076 527004 132078
rect 562404 132076 563004 132078
rect 588140 132076 588740 132078
rect -4816 132054 588740 132076
rect -4816 131818 -4634 132054
rect -4398 131818 22586 132054
rect 22822 131818 58586 132054
rect 58822 131818 94586 132054
rect 94822 131818 130586 132054
rect 130822 131818 166586 132054
rect 166822 131818 202586 132054
rect 202822 131818 238586 132054
rect 238822 131818 274586 132054
rect 274822 131818 382586 132054
rect 382822 131818 526586 132054
rect 526822 131818 562586 132054
rect 562822 131818 588322 132054
rect 588558 131818 588740 132054
rect -4816 131734 588740 131818
rect -4816 131498 -4634 131734
rect -4398 131498 22586 131734
rect 22822 131498 58586 131734
rect 58822 131498 94586 131734
rect 94822 131498 130586 131734
rect 130822 131498 166586 131734
rect 166822 131498 202586 131734
rect 202822 131498 238586 131734
rect 238822 131498 274586 131734
rect 274822 131498 382586 131734
rect 382822 131498 526586 131734
rect 526822 131498 562586 131734
rect 562822 131498 588322 131734
rect 588558 131498 588740 131734
rect -4816 131476 588740 131498
rect -4816 131474 -4216 131476
rect 22404 131474 23004 131476
rect 58404 131474 59004 131476
rect 94404 131474 95004 131476
rect 130404 131474 131004 131476
rect 166404 131474 167004 131476
rect 202404 131474 203004 131476
rect 238404 131474 239004 131476
rect 274404 131474 275004 131476
rect 382404 131474 383004 131476
rect 526404 131474 527004 131476
rect 562404 131474 563004 131476
rect 588140 131474 588740 131476
rect -2936 128476 -2336 128478
rect 18804 128476 19404 128478
rect 54804 128476 55404 128478
rect 90804 128476 91404 128478
rect 126804 128476 127404 128478
rect 162804 128476 163404 128478
rect 198804 128476 199404 128478
rect 234804 128476 235404 128478
rect 270804 128476 271404 128478
rect 300034 128476 300358 128478
rect 414804 128476 415404 128478
rect 420034 128476 420358 128478
rect 522804 128476 523404 128478
rect 558804 128476 559404 128478
rect 586260 128476 586860 128478
rect -2936 128454 586860 128476
rect -2936 128218 -2754 128454
rect -2518 128218 18986 128454
rect 19222 128218 54986 128454
rect 55222 128218 90986 128454
rect 91222 128218 126986 128454
rect 127222 128218 162986 128454
rect 163222 128218 198986 128454
rect 199222 128218 234986 128454
rect 235222 128218 270986 128454
rect 271222 128218 300078 128454
rect 300314 128218 414986 128454
rect 415222 128218 420078 128454
rect 420314 128218 522986 128454
rect 523222 128218 558986 128454
rect 559222 128218 586442 128454
rect 586678 128218 586860 128454
rect -2936 128134 586860 128218
rect -2936 127898 -2754 128134
rect -2518 127898 18986 128134
rect 19222 127898 54986 128134
rect 55222 127898 90986 128134
rect 91222 127898 126986 128134
rect 127222 127898 162986 128134
rect 163222 127898 198986 128134
rect 199222 127898 234986 128134
rect 235222 127898 270986 128134
rect 271222 127898 300078 128134
rect 300314 127898 414986 128134
rect 415222 127898 420078 128134
rect 420314 127898 522986 128134
rect 523222 127898 558986 128134
rect 559222 127898 586442 128134
rect 586678 127898 586860 128134
rect -2936 127876 586860 127898
rect -2936 127874 -2336 127876
rect 18804 127874 19404 127876
rect 54804 127874 55404 127876
rect 90804 127874 91404 127876
rect 126804 127874 127404 127876
rect 162804 127874 163404 127876
rect 198804 127874 199404 127876
rect 234804 127874 235404 127876
rect 270804 127874 271404 127876
rect 300034 127874 300358 127876
rect 414804 127874 415404 127876
rect 420034 127874 420358 127876
rect 522804 127874 523404 127876
rect 558804 127874 559404 127876
rect 586260 127874 586860 127876
rect -7636 121276 -7036 121278
rect 11604 121276 12204 121278
rect 47604 121276 48204 121278
rect 83604 121276 84204 121278
rect 119604 121276 120204 121278
rect 155604 121276 156204 121278
rect 191604 121276 192204 121278
rect 227604 121276 228204 121278
rect 263604 121276 264204 121278
rect 407604 121276 408204 121278
rect 515604 121276 516204 121278
rect 551604 121276 552204 121278
rect 590960 121276 591560 121278
rect -8576 121254 592500 121276
rect -8576 121018 -7454 121254
rect -7218 121018 11786 121254
rect 12022 121018 47786 121254
rect 48022 121018 83786 121254
rect 84022 121018 119786 121254
rect 120022 121018 155786 121254
rect 156022 121018 191786 121254
rect 192022 121018 227786 121254
rect 228022 121018 263786 121254
rect 264022 121018 407786 121254
rect 408022 121018 515786 121254
rect 516022 121018 551786 121254
rect 552022 121018 591142 121254
rect 591378 121018 592500 121254
rect -8576 120934 592500 121018
rect -8576 120698 -7454 120934
rect -7218 120698 11786 120934
rect 12022 120698 47786 120934
rect 48022 120698 83786 120934
rect 84022 120698 119786 120934
rect 120022 120698 155786 120934
rect 156022 120698 191786 120934
rect 192022 120698 227786 120934
rect 228022 120698 263786 120934
rect 264022 120698 407786 120934
rect 408022 120698 515786 120934
rect 516022 120698 551786 120934
rect 552022 120698 591142 120934
rect 591378 120698 592500 120934
rect -8576 120676 592500 120698
rect -7636 120674 -7036 120676
rect 11604 120674 12204 120676
rect 47604 120674 48204 120676
rect 83604 120674 84204 120676
rect 119604 120674 120204 120676
rect 155604 120674 156204 120676
rect 191604 120674 192204 120676
rect 227604 120674 228204 120676
rect 263604 120674 264204 120676
rect 407604 120674 408204 120676
rect 515604 120674 516204 120676
rect 551604 120674 552204 120676
rect 590960 120674 591560 120676
rect -5756 117676 -5156 117678
rect 8004 117676 8604 117678
rect 44004 117676 44604 117678
rect 80004 117676 80604 117678
rect 116004 117676 116604 117678
rect 152004 117676 152604 117678
rect 188004 117676 188604 117678
rect 224004 117676 224604 117678
rect 260004 117676 260604 117678
rect 296004 117676 296604 117678
rect 404004 117676 404604 117678
rect 512004 117676 512604 117678
rect 548004 117676 548604 117678
rect 589080 117676 589680 117678
rect -6696 117654 590620 117676
rect -6696 117418 -5574 117654
rect -5338 117418 8186 117654
rect 8422 117418 44186 117654
rect 44422 117418 80186 117654
rect 80422 117418 116186 117654
rect 116422 117418 152186 117654
rect 152422 117418 188186 117654
rect 188422 117418 224186 117654
rect 224422 117418 260186 117654
rect 260422 117418 296186 117654
rect 296422 117418 404186 117654
rect 404422 117418 512186 117654
rect 512422 117418 548186 117654
rect 548422 117418 589262 117654
rect 589498 117418 590620 117654
rect -6696 117334 590620 117418
rect -6696 117098 -5574 117334
rect -5338 117098 8186 117334
rect 8422 117098 44186 117334
rect 44422 117098 80186 117334
rect 80422 117098 116186 117334
rect 116422 117098 152186 117334
rect 152422 117098 188186 117334
rect 188422 117098 224186 117334
rect 224422 117098 260186 117334
rect 260422 117098 296186 117334
rect 296422 117098 404186 117334
rect 404422 117098 512186 117334
rect 512422 117098 548186 117334
rect 548422 117098 589262 117334
rect 589498 117098 590620 117334
rect -6696 117076 590620 117098
rect -5756 117074 -5156 117076
rect 8004 117074 8604 117076
rect 44004 117074 44604 117076
rect 80004 117074 80604 117076
rect 116004 117074 116604 117076
rect 152004 117074 152604 117076
rect 188004 117074 188604 117076
rect 224004 117074 224604 117076
rect 260004 117074 260604 117076
rect 296004 117074 296604 117076
rect 404004 117074 404604 117076
rect 512004 117074 512604 117076
rect 548004 117074 548604 117076
rect 589080 117074 589680 117076
rect -3876 114076 -3276 114078
rect 4404 114076 5004 114078
rect 40404 114076 41004 114078
rect 76404 114076 77004 114078
rect 112404 114076 113004 114078
rect 148404 114076 149004 114078
rect 184404 114076 185004 114078
rect 220404 114076 221004 114078
rect 256404 114076 257004 114078
rect 292404 114076 293004 114078
rect 400404 114076 401004 114078
rect 508404 114076 509004 114078
rect 544404 114076 545004 114078
rect 580404 114076 581004 114078
rect 587200 114076 587800 114078
rect -4816 114054 588740 114076
rect -4816 113818 -3694 114054
rect -3458 113818 4586 114054
rect 4822 113818 40586 114054
rect 40822 113818 76586 114054
rect 76822 113818 112586 114054
rect 112822 113818 148586 114054
rect 148822 113818 184586 114054
rect 184822 113818 220586 114054
rect 220822 113818 256586 114054
rect 256822 113818 292586 114054
rect 292822 113818 400586 114054
rect 400822 113818 508586 114054
rect 508822 113818 544586 114054
rect 544822 113818 580586 114054
rect 580822 113818 587382 114054
rect 587618 113818 588740 114054
rect -4816 113734 588740 113818
rect -4816 113498 -3694 113734
rect -3458 113498 4586 113734
rect 4822 113498 40586 113734
rect 40822 113498 76586 113734
rect 76822 113498 112586 113734
rect 112822 113498 148586 113734
rect 148822 113498 184586 113734
rect 184822 113498 220586 113734
rect 220822 113498 256586 113734
rect 256822 113498 292586 113734
rect 292822 113498 400586 113734
rect 400822 113498 508586 113734
rect 508822 113498 544586 113734
rect 544822 113498 580586 113734
rect 580822 113498 587382 113734
rect 587618 113498 588740 113734
rect -4816 113476 588740 113498
rect -3876 113474 -3276 113476
rect 4404 113474 5004 113476
rect 40404 113474 41004 113476
rect 76404 113474 77004 113476
rect 112404 113474 113004 113476
rect 148404 113474 149004 113476
rect 184404 113474 185004 113476
rect 220404 113474 221004 113476
rect 256404 113474 257004 113476
rect 292404 113474 293004 113476
rect 400404 113474 401004 113476
rect 508404 113474 509004 113476
rect 544404 113474 545004 113476
rect 580404 113474 581004 113476
rect 587200 113474 587800 113476
rect -1996 110476 -1396 110478
rect 804 110476 1404 110478
rect 36804 110476 37404 110478
rect 72804 110476 73404 110478
rect 108804 110476 109404 110478
rect 144804 110476 145404 110478
rect 180804 110476 181404 110478
rect 216804 110476 217404 110478
rect 252804 110476 253404 110478
rect 288804 110476 289404 110478
rect 396804 110476 397404 110478
rect 504804 110476 505404 110478
rect 540804 110476 541404 110478
rect 576804 110476 577404 110478
rect 585320 110476 585920 110478
rect -2936 110454 586860 110476
rect -2936 110218 -1814 110454
rect -1578 110218 986 110454
rect 1222 110218 36986 110454
rect 37222 110218 72986 110454
rect 73222 110218 108986 110454
rect 109222 110218 144986 110454
rect 145222 110218 180986 110454
rect 181222 110218 216986 110454
rect 217222 110218 252986 110454
rect 253222 110218 288986 110454
rect 289222 110218 396986 110454
rect 397222 110218 504986 110454
rect 505222 110218 540986 110454
rect 541222 110218 576986 110454
rect 577222 110218 585502 110454
rect 585738 110218 586860 110454
rect -2936 110134 586860 110218
rect -2936 109898 -1814 110134
rect -1578 109898 986 110134
rect 1222 109898 36986 110134
rect 37222 109898 72986 110134
rect 73222 109898 108986 110134
rect 109222 109898 144986 110134
rect 145222 109898 180986 110134
rect 181222 109898 216986 110134
rect 217222 109898 252986 110134
rect 253222 109898 288986 110134
rect 289222 109898 396986 110134
rect 397222 109898 504986 110134
rect 505222 109898 540986 110134
rect 541222 109898 576986 110134
rect 577222 109898 585502 110134
rect 585738 109898 586860 110134
rect -2936 109876 586860 109898
rect -1996 109874 -1396 109876
rect 804 109874 1404 109876
rect 36804 109874 37404 109876
rect 72804 109874 73404 109876
rect 108804 109874 109404 109876
rect 144804 109874 145404 109876
rect 180804 109874 181404 109876
rect 216804 109874 217404 109876
rect 252804 109874 253404 109876
rect 288804 109874 289404 109876
rect 396804 109874 397404 109876
rect 504804 109874 505404 109876
rect 540804 109874 541404 109876
rect 576804 109874 577404 109876
rect 585320 109874 585920 109876
rect -8576 103276 -7976 103278
rect 29604 103276 30204 103278
rect 65604 103276 66204 103278
rect 101604 103276 102204 103278
rect 137604 103276 138204 103278
rect 173604 103276 174204 103278
rect 209604 103276 210204 103278
rect 245604 103276 246204 103278
rect 281604 103276 282204 103278
rect 317604 103276 318204 103278
rect 353604 103276 354204 103278
rect 389604 103276 390204 103278
rect 425604 103276 426204 103278
rect 461604 103276 462204 103278
rect 497604 103276 498204 103278
rect 533604 103276 534204 103278
rect 569604 103276 570204 103278
rect 591900 103276 592500 103278
rect -8576 103254 592500 103276
rect -8576 103018 -8394 103254
rect -8158 103018 29786 103254
rect 30022 103018 65786 103254
rect 66022 103018 101786 103254
rect 102022 103018 137786 103254
rect 138022 103018 173786 103254
rect 174022 103018 209786 103254
rect 210022 103018 245786 103254
rect 246022 103018 281786 103254
rect 282022 103018 317786 103254
rect 318022 103018 353786 103254
rect 354022 103018 389786 103254
rect 390022 103018 425786 103254
rect 426022 103018 461786 103254
rect 462022 103018 497786 103254
rect 498022 103018 533786 103254
rect 534022 103018 569786 103254
rect 570022 103018 592082 103254
rect 592318 103018 592500 103254
rect -8576 102934 592500 103018
rect -8576 102698 -8394 102934
rect -8158 102698 29786 102934
rect 30022 102698 65786 102934
rect 66022 102698 101786 102934
rect 102022 102698 137786 102934
rect 138022 102698 173786 102934
rect 174022 102698 209786 102934
rect 210022 102698 245786 102934
rect 246022 102698 281786 102934
rect 282022 102698 317786 102934
rect 318022 102698 353786 102934
rect 354022 102698 389786 102934
rect 390022 102698 425786 102934
rect 426022 102698 461786 102934
rect 462022 102698 497786 102934
rect 498022 102698 533786 102934
rect 534022 102698 569786 102934
rect 570022 102698 592082 102934
rect 592318 102698 592500 102934
rect -8576 102676 592500 102698
rect -8576 102674 -7976 102676
rect 29604 102674 30204 102676
rect 65604 102674 66204 102676
rect 101604 102674 102204 102676
rect 137604 102674 138204 102676
rect 173604 102674 174204 102676
rect 209604 102674 210204 102676
rect 245604 102674 246204 102676
rect 281604 102674 282204 102676
rect 317604 102674 318204 102676
rect 353604 102674 354204 102676
rect 389604 102674 390204 102676
rect 425604 102674 426204 102676
rect 461604 102674 462204 102676
rect 497604 102674 498204 102676
rect 533604 102674 534204 102676
rect 569604 102674 570204 102676
rect 591900 102674 592500 102676
rect -6696 99676 -6096 99678
rect 26004 99676 26604 99678
rect 62004 99676 62604 99678
rect 98004 99676 98604 99678
rect 134004 99676 134604 99678
rect 170004 99676 170604 99678
rect 206004 99676 206604 99678
rect 242004 99676 242604 99678
rect 278004 99676 278604 99678
rect 314004 99676 314604 99678
rect 350004 99676 350604 99678
rect 386004 99676 386604 99678
rect 422004 99676 422604 99678
rect 458004 99676 458604 99678
rect 494004 99676 494604 99678
rect 530004 99676 530604 99678
rect 566004 99676 566604 99678
rect 590020 99676 590620 99678
rect -6696 99654 590620 99676
rect -6696 99418 -6514 99654
rect -6278 99418 26186 99654
rect 26422 99418 62186 99654
rect 62422 99418 98186 99654
rect 98422 99418 134186 99654
rect 134422 99418 170186 99654
rect 170422 99418 206186 99654
rect 206422 99418 242186 99654
rect 242422 99418 278186 99654
rect 278422 99418 314186 99654
rect 314422 99418 350186 99654
rect 350422 99418 386186 99654
rect 386422 99418 422186 99654
rect 422422 99418 458186 99654
rect 458422 99418 494186 99654
rect 494422 99418 530186 99654
rect 530422 99418 566186 99654
rect 566422 99418 590202 99654
rect 590438 99418 590620 99654
rect -6696 99334 590620 99418
rect -6696 99098 -6514 99334
rect -6278 99098 26186 99334
rect 26422 99098 62186 99334
rect 62422 99098 98186 99334
rect 98422 99098 134186 99334
rect 134422 99098 170186 99334
rect 170422 99098 206186 99334
rect 206422 99098 242186 99334
rect 242422 99098 278186 99334
rect 278422 99098 314186 99334
rect 314422 99098 350186 99334
rect 350422 99098 386186 99334
rect 386422 99098 422186 99334
rect 422422 99098 458186 99334
rect 458422 99098 494186 99334
rect 494422 99098 530186 99334
rect 530422 99098 566186 99334
rect 566422 99098 590202 99334
rect 590438 99098 590620 99334
rect -6696 99076 590620 99098
rect -6696 99074 -6096 99076
rect 26004 99074 26604 99076
rect 62004 99074 62604 99076
rect 98004 99074 98604 99076
rect 134004 99074 134604 99076
rect 170004 99074 170604 99076
rect 206004 99074 206604 99076
rect 242004 99074 242604 99076
rect 278004 99074 278604 99076
rect 314004 99074 314604 99076
rect 350004 99074 350604 99076
rect 386004 99074 386604 99076
rect 422004 99074 422604 99076
rect 458004 99074 458604 99076
rect 494004 99074 494604 99076
rect 530004 99074 530604 99076
rect 566004 99074 566604 99076
rect 590020 99074 590620 99076
rect -4816 96076 -4216 96078
rect 22404 96076 23004 96078
rect 58404 96076 59004 96078
rect 94404 96076 95004 96078
rect 130404 96076 131004 96078
rect 166404 96076 167004 96078
rect 202404 96076 203004 96078
rect 238404 96076 239004 96078
rect 274404 96076 275004 96078
rect 310404 96076 311004 96078
rect 346404 96076 347004 96078
rect 382404 96076 383004 96078
rect 418404 96076 419004 96078
rect 454404 96076 455004 96078
rect 490404 96076 491004 96078
rect 526404 96076 527004 96078
rect 562404 96076 563004 96078
rect 588140 96076 588740 96078
rect -4816 96054 588740 96076
rect -4816 95818 -4634 96054
rect -4398 95818 22586 96054
rect 22822 95818 58586 96054
rect 58822 95818 94586 96054
rect 94822 95818 130586 96054
rect 130822 95818 166586 96054
rect 166822 95818 202586 96054
rect 202822 95818 238586 96054
rect 238822 95818 274586 96054
rect 274822 95818 310586 96054
rect 310822 95818 346586 96054
rect 346822 95818 382586 96054
rect 382822 95818 418586 96054
rect 418822 95818 454586 96054
rect 454822 95818 490586 96054
rect 490822 95818 526586 96054
rect 526822 95818 562586 96054
rect 562822 95818 588322 96054
rect 588558 95818 588740 96054
rect -4816 95734 588740 95818
rect -4816 95498 -4634 95734
rect -4398 95498 22586 95734
rect 22822 95498 58586 95734
rect 58822 95498 94586 95734
rect 94822 95498 130586 95734
rect 130822 95498 166586 95734
rect 166822 95498 202586 95734
rect 202822 95498 238586 95734
rect 238822 95498 274586 95734
rect 274822 95498 310586 95734
rect 310822 95498 346586 95734
rect 346822 95498 382586 95734
rect 382822 95498 418586 95734
rect 418822 95498 454586 95734
rect 454822 95498 490586 95734
rect 490822 95498 526586 95734
rect 526822 95498 562586 95734
rect 562822 95498 588322 95734
rect 588558 95498 588740 95734
rect -4816 95476 588740 95498
rect -4816 95474 -4216 95476
rect 22404 95474 23004 95476
rect 58404 95474 59004 95476
rect 94404 95474 95004 95476
rect 130404 95474 131004 95476
rect 166404 95474 167004 95476
rect 202404 95474 203004 95476
rect 238404 95474 239004 95476
rect 274404 95474 275004 95476
rect 310404 95474 311004 95476
rect 346404 95474 347004 95476
rect 382404 95474 383004 95476
rect 418404 95474 419004 95476
rect 454404 95474 455004 95476
rect 490404 95474 491004 95476
rect 526404 95474 527004 95476
rect 562404 95474 563004 95476
rect 588140 95474 588740 95476
rect -2936 92476 -2336 92478
rect 18804 92476 19404 92478
rect 54804 92476 55404 92478
rect 90804 92476 91404 92478
rect 126804 92476 127404 92478
rect 162804 92476 163404 92478
rect 198804 92476 199404 92478
rect 234804 92476 235404 92478
rect 270804 92476 271404 92478
rect 306804 92476 307404 92478
rect 342804 92476 343404 92478
rect 378804 92476 379404 92478
rect 414804 92476 415404 92478
rect 450804 92476 451404 92478
rect 486804 92476 487404 92478
rect 522804 92476 523404 92478
rect 558804 92476 559404 92478
rect 586260 92476 586860 92478
rect -2936 92454 586860 92476
rect -2936 92218 -2754 92454
rect -2518 92218 18986 92454
rect 19222 92218 54986 92454
rect 55222 92218 90986 92454
rect 91222 92218 126986 92454
rect 127222 92218 162986 92454
rect 163222 92218 198986 92454
rect 199222 92218 234986 92454
rect 235222 92218 270986 92454
rect 271222 92218 306986 92454
rect 307222 92218 342986 92454
rect 343222 92218 378986 92454
rect 379222 92218 414986 92454
rect 415222 92218 450986 92454
rect 451222 92218 486986 92454
rect 487222 92218 522986 92454
rect 523222 92218 558986 92454
rect 559222 92218 586442 92454
rect 586678 92218 586860 92454
rect -2936 92134 586860 92218
rect -2936 91898 -2754 92134
rect -2518 91898 18986 92134
rect 19222 91898 54986 92134
rect 55222 91898 90986 92134
rect 91222 91898 126986 92134
rect 127222 91898 162986 92134
rect 163222 91898 198986 92134
rect 199222 91898 234986 92134
rect 235222 91898 270986 92134
rect 271222 91898 306986 92134
rect 307222 91898 342986 92134
rect 343222 91898 378986 92134
rect 379222 91898 414986 92134
rect 415222 91898 450986 92134
rect 451222 91898 486986 92134
rect 487222 91898 522986 92134
rect 523222 91898 558986 92134
rect 559222 91898 586442 92134
rect 586678 91898 586860 92134
rect -2936 91876 586860 91898
rect -2936 91874 -2336 91876
rect 18804 91874 19404 91876
rect 54804 91874 55404 91876
rect 90804 91874 91404 91876
rect 126804 91874 127404 91876
rect 162804 91874 163404 91876
rect 198804 91874 199404 91876
rect 234804 91874 235404 91876
rect 270804 91874 271404 91876
rect 306804 91874 307404 91876
rect 342804 91874 343404 91876
rect 378804 91874 379404 91876
rect 414804 91874 415404 91876
rect 450804 91874 451404 91876
rect 486804 91874 487404 91876
rect 522804 91874 523404 91876
rect 558804 91874 559404 91876
rect 586260 91874 586860 91876
rect -7636 85276 -7036 85278
rect 11604 85276 12204 85278
rect 47604 85276 48204 85278
rect 83604 85276 84204 85278
rect 119604 85276 120204 85278
rect 155604 85276 156204 85278
rect 191604 85276 192204 85278
rect 227604 85276 228204 85278
rect 263604 85276 264204 85278
rect 299604 85276 300204 85278
rect 335604 85276 336204 85278
rect 371604 85276 372204 85278
rect 407604 85276 408204 85278
rect 443604 85276 444204 85278
rect 479604 85276 480204 85278
rect 515604 85276 516204 85278
rect 551604 85276 552204 85278
rect 590960 85276 591560 85278
rect -8576 85254 592500 85276
rect -8576 85018 -7454 85254
rect -7218 85018 11786 85254
rect 12022 85018 47786 85254
rect 48022 85018 83786 85254
rect 84022 85018 119786 85254
rect 120022 85018 155786 85254
rect 156022 85018 191786 85254
rect 192022 85018 227786 85254
rect 228022 85018 263786 85254
rect 264022 85018 299786 85254
rect 300022 85018 335786 85254
rect 336022 85018 371786 85254
rect 372022 85018 407786 85254
rect 408022 85018 443786 85254
rect 444022 85018 479786 85254
rect 480022 85018 515786 85254
rect 516022 85018 551786 85254
rect 552022 85018 591142 85254
rect 591378 85018 592500 85254
rect -8576 84934 592500 85018
rect -8576 84698 -7454 84934
rect -7218 84698 11786 84934
rect 12022 84698 47786 84934
rect 48022 84698 83786 84934
rect 84022 84698 119786 84934
rect 120022 84698 155786 84934
rect 156022 84698 191786 84934
rect 192022 84698 227786 84934
rect 228022 84698 263786 84934
rect 264022 84698 299786 84934
rect 300022 84698 335786 84934
rect 336022 84698 371786 84934
rect 372022 84698 407786 84934
rect 408022 84698 443786 84934
rect 444022 84698 479786 84934
rect 480022 84698 515786 84934
rect 516022 84698 551786 84934
rect 552022 84698 591142 84934
rect 591378 84698 592500 84934
rect -8576 84676 592500 84698
rect -7636 84674 -7036 84676
rect 11604 84674 12204 84676
rect 47604 84674 48204 84676
rect 83604 84674 84204 84676
rect 119604 84674 120204 84676
rect 155604 84674 156204 84676
rect 191604 84674 192204 84676
rect 227604 84674 228204 84676
rect 263604 84674 264204 84676
rect 299604 84674 300204 84676
rect 335604 84674 336204 84676
rect 371604 84674 372204 84676
rect 407604 84674 408204 84676
rect 443604 84674 444204 84676
rect 479604 84674 480204 84676
rect 515604 84674 516204 84676
rect 551604 84674 552204 84676
rect 590960 84674 591560 84676
rect -5756 81676 -5156 81678
rect 8004 81676 8604 81678
rect 44004 81676 44604 81678
rect 80004 81676 80604 81678
rect 116004 81676 116604 81678
rect 152004 81676 152604 81678
rect 188004 81676 188604 81678
rect 224004 81676 224604 81678
rect 260004 81676 260604 81678
rect 296004 81676 296604 81678
rect 332004 81676 332604 81678
rect 368004 81676 368604 81678
rect 404004 81676 404604 81678
rect 440004 81676 440604 81678
rect 476004 81676 476604 81678
rect 512004 81676 512604 81678
rect 548004 81676 548604 81678
rect 589080 81676 589680 81678
rect -6696 81654 590620 81676
rect -6696 81418 -5574 81654
rect -5338 81418 8186 81654
rect 8422 81418 44186 81654
rect 44422 81418 80186 81654
rect 80422 81418 116186 81654
rect 116422 81418 152186 81654
rect 152422 81418 188186 81654
rect 188422 81418 224186 81654
rect 224422 81418 260186 81654
rect 260422 81418 296186 81654
rect 296422 81418 332186 81654
rect 332422 81418 368186 81654
rect 368422 81418 404186 81654
rect 404422 81418 440186 81654
rect 440422 81418 476186 81654
rect 476422 81418 512186 81654
rect 512422 81418 548186 81654
rect 548422 81418 589262 81654
rect 589498 81418 590620 81654
rect -6696 81334 590620 81418
rect -6696 81098 -5574 81334
rect -5338 81098 8186 81334
rect 8422 81098 44186 81334
rect 44422 81098 80186 81334
rect 80422 81098 116186 81334
rect 116422 81098 152186 81334
rect 152422 81098 188186 81334
rect 188422 81098 224186 81334
rect 224422 81098 260186 81334
rect 260422 81098 296186 81334
rect 296422 81098 332186 81334
rect 332422 81098 368186 81334
rect 368422 81098 404186 81334
rect 404422 81098 440186 81334
rect 440422 81098 476186 81334
rect 476422 81098 512186 81334
rect 512422 81098 548186 81334
rect 548422 81098 589262 81334
rect 589498 81098 590620 81334
rect -6696 81076 590620 81098
rect -5756 81074 -5156 81076
rect 8004 81074 8604 81076
rect 44004 81074 44604 81076
rect 80004 81074 80604 81076
rect 116004 81074 116604 81076
rect 152004 81074 152604 81076
rect 188004 81074 188604 81076
rect 224004 81074 224604 81076
rect 260004 81074 260604 81076
rect 296004 81074 296604 81076
rect 332004 81074 332604 81076
rect 368004 81074 368604 81076
rect 404004 81074 404604 81076
rect 440004 81074 440604 81076
rect 476004 81074 476604 81076
rect 512004 81074 512604 81076
rect 548004 81074 548604 81076
rect 589080 81074 589680 81076
rect -3876 78076 -3276 78078
rect 4404 78076 5004 78078
rect 40404 78076 41004 78078
rect 76404 78076 77004 78078
rect 112404 78076 113004 78078
rect 148404 78076 149004 78078
rect 184404 78076 185004 78078
rect 220404 78076 221004 78078
rect 256404 78076 257004 78078
rect 292404 78076 293004 78078
rect 328404 78076 329004 78078
rect 364404 78076 365004 78078
rect 400404 78076 401004 78078
rect 436404 78076 437004 78078
rect 472404 78076 473004 78078
rect 508404 78076 509004 78078
rect 544404 78076 545004 78078
rect 580404 78076 581004 78078
rect 587200 78076 587800 78078
rect -4816 78054 588740 78076
rect -4816 77818 -3694 78054
rect -3458 77818 4586 78054
rect 4822 77818 40586 78054
rect 40822 77818 76586 78054
rect 76822 77818 112586 78054
rect 112822 77818 148586 78054
rect 148822 77818 184586 78054
rect 184822 77818 220586 78054
rect 220822 77818 256586 78054
rect 256822 77818 292586 78054
rect 292822 77818 328586 78054
rect 328822 77818 364586 78054
rect 364822 77818 400586 78054
rect 400822 77818 436586 78054
rect 436822 77818 472586 78054
rect 472822 77818 508586 78054
rect 508822 77818 544586 78054
rect 544822 77818 580586 78054
rect 580822 77818 587382 78054
rect 587618 77818 588740 78054
rect -4816 77734 588740 77818
rect -4816 77498 -3694 77734
rect -3458 77498 4586 77734
rect 4822 77498 40586 77734
rect 40822 77498 76586 77734
rect 76822 77498 112586 77734
rect 112822 77498 148586 77734
rect 148822 77498 184586 77734
rect 184822 77498 220586 77734
rect 220822 77498 256586 77734
rect 256822 77498 292586 77734
rect 292822 77498 328586 77734
rect 328822 77498 364586 77734
rect 364822 77498 400586 77734
rect 400822 77498 436586 77734
rect 436822 77498 472586 77734
rect 472822 77498 508586 77734
rect 508822 77498 544586 77734
rect 544822 77498 580586 77734
rect 580822 77498 587382 77734
rect 587618 77498 588740 77734
rect -4816 77476 588740 77498
rect -3876 77474 -3276 77476
rect 4404 77474 5004 77476
rect 40404 77474 41004 77476
rect 76404 77474 77004 77476
rect 112404 77474 113004 77476
rect 148404 77474 149004 77476
rect 184404 77474 185004 77476
rect 220404 77474 221004 77476
rect 256404 77474 257004 77476
rect 292404 77474 293004 77476
rect 328404 77474 329004 77476
rect 364404 77474 365004 77476
rect 400404 77474 401004 77476
rect 436404 77474 437004 77476
rect 472404 77474 473004 77476
rect 508404 77474 509004 77476
rect 544404 77474 545004 77476
rect 580404 77474 581004 77476
rect 587200 77474 587800 77476
rect -1996 74476 -1396 74478
rect 804 74476 1404 74478
rect 36804 74476 37404 74478
rect 72804 74476 73404 74478
rect 108804 74476 109404 74478
rect 144804 74476 145404 74478
rect 180804 74476 181404 74478
rect 216804 74476 217404 74478
rect 252804 74476 253404 74478
rect 288804 74476 289404 74478
rect 324804 74476 325404 74478
rect 360804 74476 361404 74478
rect 396804 74476 397404 74478
rect 432804 74476 433404 74478
rect 468804 74476 469404 74478
rect 504804 74476 505404 74478
rect 540804 74476 541404 74478
rect 576804 74476 577404 74478
rect 585320 74476 585920 74478
rect -2936 74454 586860 74476
rect -2936 74218 -1814 74454
rect -1578 74218 986 74454
rect 1222 74218 36986 74454
rect 37222 74218 72986 74454
rect 73222 74218 108986 74454
rect 109222 74218 144986 74454
rect 145222 74218 180986 74454
rect 181222 74218 216986 74454
rect 217222 74218 252986 74454
rect 253222 74218 288986 74454
rect 289222 74218 324986 74454
rect 325222 74218 360986 74454
rect 361222 74218 396986 74454
rect 397222 74218 432986 74454
rect 433222 74218 468986 74454
rect 469222 74218 504986 74454
rect 505222 74218 540986 74454
rect 541222 74218 576986 74454
rect 577222 74218 585502 74454
rect 585738 74218 586860 74454
rect -2936 74134 586860 74218
rect -2936 73898 -1814 74134
rect -1578 73898 986 74134
rect 1222 73898 36986 74134
rect 37222 73898 72986 74134
rect 73222 73898 108986 74134
rect 109222 73898 144986 74134
rect 145222 73898 180986 74134
rect 181222 73898 216986 74134
rect 217222 73898 252986 74134
rect 253222 73898 288986 74134
rect 289222 73898 324986 74134
rect 325222 73898 360986 74134
rect 361222 73898 396986 74134
rect 397222 73898 432986 74134
rect 433222 73898 468986 74134
rect 469222 73898 504986 74134
rect 505222 73898 540986 74134
rect 541222 73898 576986 74134
rect 577222 73898 585502 74134
rect 585738 73898 586860 74134
rect -2936 73876 586860 73898
rect -1996 73874 -1396 73876
rect 804 73874 1404 73876
rect 36804 73874 37404 73876
rect 72804 73874 73404 73876
rect 108804 73874 109404 73876
rect 144804 73874 145404 73876
rect 180804 73874 181404 73876
rect 216804 73874 217404 73876
rect 252804 73874 253404 73876
rect 288804 73874 289404 73876
rect 324804 73874 325404 73876
rect 360804 73874 361404 73876
rect 396804 73874 397404 73876
rect 432804 73874 433404 73876
rect 468804 73874 469404 73876
rect 504804 73874 505404 73876
rect 540804 73874 541404 73876
rect 576804 73874 577404 73876
rect 585320 73874 585920 73876
rect -8576 67276 -7976 67278
rect 29604 67276 30204 67278
rect 65604 67276 66204 67278
rect 101604 67276 102204 67278
rect 137604 67276 138204 67278
rect 173604 67276 174204 67278
rect 209604 67276 210204 67278
rect 245604 67276 246204 67278
rect 281604 67276 282204 67278
rect 317604 67276 318204 67278
rect 353604 67276 354204 67278
rect 389604 67276 390204 67278
rect 425604 67276 426204 67278
rect 461604 67276 462204 67278
rect 497604 67276 498204 67278
rect 533604 67276 534204 67278
rect 569604 67276 570204 67278
rect 591900 67276 592500 67278
rect -8576 67254 592500 67276
rect -8576 67018 -8394 67254
rect -8158 67018 29786 67254
rect 30022 67018 65786 67254
rect 66022 67018 101786 67254
rect 102022 67018 137786 67254
rect 138022 67018 173786 67254
rect 174022 67018 209786 67254
rect 210022 67018 245786 67254
rect 246022 67018 281786 67254
rect 282022 67018 317786 67254
rect 318022 67018 353786 67254
rect 354022 67018 389786 67254
rect 390022 67018 425786 67254
rect 426022 67018 461786 67254
rect 462022 67018 497786 67254
rect 498022 67018 533786 67254
rect 534022 67018 569786 67254
rect 570022 67018 592082 67254
rect 592318 67018 592500 67254
rect -8576 66934 592500 67018
rect -8576 66698 -8394 66934
rect -8158 66698 29786 66934
rect 30022 66698 65786 66934
rect 66022 66698 101786 66934
rect 102022 66698 137786 66934
rect 138022 66698 173786 66934
rect 174022 66698 209786 66934
rect 210022 66698 245786 66934
rect 246022 66698 281786 66934
rect 282022 66698 317786 66934
rect 318022 66698 353786 66934
rect 354022 66698 389786 66934
rect 390022 66698 425786 66934
rect 426022 66698 461786 66934
rect 462022 66698 497786 66934
rect 498022 66698 533786 66934
rect 534022 66698 569786 66934
rect 570022 66698 592082 66934
rect 592318 66698 592500 66934
rect -8576 66676 592500 66698
rect -8576 66674 -7976 66676
rect 29604 66674 30204 66676
rect 65604 66674 66204 66676
rect 101604 66674 102204 66676
rect 137604 66674 138204 66676
rect 173604 66674 174204 66676
rect 209604 66674 210204 66676
rect 245604 66674 246204 66676
rect 281604 66674 282204 66676
rect 317604 66674 318204 66676
rect 353604 66674 354204 66676
rect 389604 66674 390204 66676
rect 425604 66674 426204 66676
rect 461604 66674 462204 66676
rect 497604 66674 498204 66676
rect 533604 66674 534204 66676
rect 569604 66674 570204 66676
rect 591900 66674 592500 66676
rect -6696 63676 -6096 63678
rect 26004 63676 26604 63678
rect 62004 63676 62604 63678
rect 98004 63676 98604 63678
rect 134004 63676 134604 63678
rect 170004 63676 170604 63678
rect 206004 63676 206604 63678
rect 242004 63676 242604 63678
rect 278004 63676 278604 63678
rect 314004 63676 314604 63678
rect 350004 63676 350604 63678
rect 386004 63676 386604 63678
rect 422004 63676 422604 63678
rect 458004 63676 458604 63678
rect 494004 63676 494604 63678
rect 530004 63676 530604 63678
rect 566004 63676 566604 63678
rect 590020 63676 590620 63678
rect -6696 63654 590620 63676
rect -6696 63418 -6514 63654
rect -6278 63418 26186 63654
rect 26422 63418 62186 63654
rect 62422 63418 98186 63654
rect 98422 63418 134186 63654
rect 134422 63418 170186 63654
rect 170422 63418 206186 63654
rect 206422 63418 242186 63654
rect 242422 63418 278186 63654
rect 278422 63418 314186 63654
rect 314422 63418 350186 63654
rect 350422 63418 386186 63654
rect 386422 63418 422186 63654
rect 422422 63418 458186 63654
rect 458422 63418 494186 63654
rect 494422 63418 530186 63654
rect 530422 63418 566186 63654
rect 566422 63418 590202 63654
rect 590438 63418 590620 63654
rect -6696 63334 590620 63418
rect -6696 63098 -6514 63334
rect -6278 63098 26186 63334
rect 26422 63098 62186 63334
rect 62422 63098 98186 63334
rect 98422 63098 134186 63334
rect 134422 63098 170186 63334
rect 170422 63098 206186 63334
rect 206422 63098 242186 63334
rect 242422 63098 278186 63334
rect 278422 63098 314186 63334
rect 314422 63098 350186 63334
rect 350422 63098 386186 63334
rect 386422 63098 422186 63334
rect 422422 63098 458186 63334
rect 458422 63098 494186 63334
rect 494422 63098 530186 63334
rect 530422 63098 566186 63334
rect 566422 63098 590202 63334
rect 590438 63098 590620 63334
rect -6696 63076 590620 63098
rect -6696 63074 -6096 63076
rect 26004 63074 26604 63076
rect 62004 63074 62604 63076
rect 98004 63074 98604 63076
rect 134004 63074 134604 63076
rect 170004 63074 170604 63076
rect 206004 63074 206604 63076
rect 242004 63074 242604 63076
rect 278004 63074 278604 63076
rect 314004 63074 314604 63076
rect 350004 63074 350604 63076
rect 386004 63074 386604 63076
rect 422004 63074 422604 63076
rect 458004 63074 458604 63076
rect 494004 63074 494604 63076
rect 530004 63074 530604 63076
rect 566004 63074 566604 63076
rect 590020 63074 590620 63076
rect -4816 60076 -4216 60078
rect 22404 60076 23004 60078
rect 58404 60076 59004 60078
rect 94404 60076 95004 60078
rect 130404 60076 131004 60078
rect 166404 60076 167004 60078
rect 202404 60076 203004 60078
rect 238404 60076 239004 60078
rect 274404 60076 275004 60078
rect 310404 60076 311004 60078
rect 346404 60076 347004 60078
rect 382404 60076 383004 60078
rect 418404 60076 419004 60078
rect 454404 60076 455004 60078
rect 490404 60076 491004 60078
rect 526404 60076 527004 60078
rect 562404 60076 563004 60078
rect 588140 60076 588740 60078
rect -4816 60054 588740 60076
rect -4816 59818 -4634 60054
rect -4398 59818 22586 60054
rect 22822 59818 58586 60054
rect 58822 59818 94586 60054
rect 94822 59818 130586 60054
rect 130822 59818 166586 60054
rect 166822 59818 202586 60054
rect 202822 59818 238586 60054
rect 238822 59818 274586 60054
rect 274822 59818 310586 60054
rect 310822 59818 346586 60054
rect 346822 59818 382586 60054
rect 382822 59818 418586 60054
rect 418822 59818 454586 60054
rect 454822 59818 490586 60054
rect 490822 59818 526586 60054
rect 526822 59818 562586 60054
rect 562822 59818 588322 60054
rect 588558 59818 588740 60054
rect -4816 59734 588740 59818
rect -4816 59498 -4634 59734
rect -4398 59498 22586 59734
rect 22822 59498 58586 59734
rect 58822 59498 94586 59734
rect 94822 59498 130586 59734
rect 130822 59498 166586 59734
rect 166822 59498 202586 59734
rect 202822 59498 238586 59734
rect 238822 59498 274586 59734
rect 274822 59498 310586 59734
rect 310822 59498 346586 59734
rect 346822 59498 382586 59734
rect 382822 59498 418586 59734
rect 418822 59498 454586 59734
rect 454822 59498 490586 59734
rect 490822 59498 526586 59734
rect 526822 59498 562586 59734
rect 562822 59498 588322 59734
rect 588558 59498 588740 59734
rect -4816 59476 588740 59498
rect -4816 59474 -4216 59476
rect 22404 59474 23004 59476
rect 58404 59474 59004 59476
rect 94404 59474 95004 59476
rect 130404 59474 131004 59476
rect 166404 59474 167004 59476
rect 202404 59474 203004 59476
rect 238404 59474 239004 59476
rect 274404 59474 275004 59476
rect 310404 59474 311004 59476
rect 346404 59474 347004 59476
rect 382404 59474 383004 59476
rect 418404 59474 419004 59476
rect 454404 59474 455004 59476
rect 490404 59474 491004 59476
rect 526404 59474 527004 59476
rect 562404 59474 563004 59476
rect 588140 59474 588740 59476
rect -2936 56476 -2336 56478
rect 18804 56476 19404 56478
rect 54804 56476 55404 56478
rect 90804 56476 91404 56478
rect 126804 56476 127404 56478
rect 162804 56476 163404 56478
rect 198804 56476 199404 56478
rect 234804 56476 235404 56478
rect 270804 56476 271404 56478
rect 306804 56476 307404 56478
rect 342804 56476 343404 56478
rect 378804 56476 379404 56478
rect 414804 56476 415404 56478
rect 450804 56476 451404 56478
rect 486804 56476 487404 56478
rect 522804 56476 523404 56478
rect 558804 56476 559404 56478
rect 586260 56476 586860 56478
rect -2936 56454 586860 56476
rect -2936 56218 -2754 56454
rect -2518 56218 18986 56454
rect 19222 56218 54986 56454
rect 55222 56218 90986 56454
rect 91222 56218 126986 56454
rect 127222 56218 162986 56454
rect 163222 56218 198986 56454
rect 199222 56218 234986 56454
rect 235222 56218 270986 56454
rect 271222 56218 306986 56454
rect 307222 56218 342986 56454
rect 343222 56218 378986 56454
rect 379222 56218 414986 56454
rect 415222 56218 450986 56454
rect 451222 56218 486986 56454
rect 487222 56218 522986 56454
rect 523222 56218 558986 56454
rect 559222 56218 586442 56454
rect 586678 56218 586860 56454
rect -2936 56134 586860 56218
rect -2936 55898 -2754 56134
rect -2518 55898 18986 56134
rect 19222 55898 54986 56134
rect 55222 55898 90986 56134
rect 91222 55898 126986 56134
rect 127222 55898 162986 56134
rect 163222 55898 198986 56134
rect 199222 55898 234986 56134
rect 235222 55898 270986 56134
rect 271222 55898 306986 56134
rect 307222 55898 342986 56134
rect 343222 55898 378986 56134
rect 379222 55898 414986 56134
rect 415222 55898 450986 56134
rect 451222 55898 486986 56134
rect 487222 55898 522986 56134
rect 523222 55898 558986 56134
rect 559222 55898 586442 56134
rect 586678 55898 586860 56134
rect -2936 55876 586860 55898
rect -2936 55874 -2336 55876
rect 18804 55874 19404 55876
rect 54804 55874 55404 55876
rect 90804 55874 91404 55876
rect 126804 55874 127404 55876
rect 162804 55874 163404 55876
rect 198804 55874 199404 55876
rect 234804 55874 235404 55876
rect 270804 55874 271404 55876
rect 306804 55874 307404 55876
rect 342804 55874 343404 55876
rect 378804 55874 379404 55876
rect 414804 55874 415404 55876
rect 450804 55874 451404 55876
rect 486804 55874 487404 55876
rect 522804 55874 523404 55876
rect 558804 55874 559404 55876
rect 586260 55874 586860 55876
rect -7636 49276 -7036 49278
rect 11604 49276 12204 49278
rect 47604 49276 48204 49278
rect 83604 49276 84204 49278
rect 119604 49276 120204 49278
rect 155604 49276 156204 49278
rect 191604 49276 192204 49278
rect 227604 49276 228204 49278
rect 263604 49276 264204 49278
rect 299604 49276 300204 49278
rect 335604 49276 336204 49278
rect 371604 49276 372204 49278
rect 407604 49276 408204 49278
rect 443604 49276 444204 49278
rect 479604 49276 480204 49278
rect 515604 49276 516204 49278
rect 551604 49276 552204 49278
rect 590960 49276 591560 49278
rect -8576 49254 592500 49276
rect -8576 49018 -7454 49254
rect -7218 49018 11786 49254
rect 12022 49018 47786 49254
rect 48022 49018 83786 49254
rect 84022 49018 119786 49254
rect 120022 49018 155786 49254
rect 156022 49018 191786 49254
rect 192022 49018 227786 49254
rect 228022 49018 263786 49254
rect 264022 49018 299786 49254
rect 300022 49018 335786 49254
rect 336022 49018 371786 49254
rect 372022 49018 407786 49254
rect 408022 49018 443786 49254
rect 444022 49018 479786 49254
rect 480022 49018 515786 49254
rect 516022 49018 551786 49254
rect 552022 49018 591142 49254
rect 591378 49018 592500 49254
rect -8576 48934 592500 49018
rect -8576 48698 -7454 48934
rect -7218 48698 11786 48934
rect 12022 48698 47786 48934
rect 48022 48698 83786 48934
rect 84022 48698 119786 48934
rect 120022 48698 155786 48934
rect 156022 48698 191786 48934
rect 192022 48698 227786 48934
rect 228022 48698 263786 48934
rect 264022 48698 299786 48934
rect 300022 48698 335786 48934
rect 336022 48698 371786 48934
rect 372022 48698 407786 48934
rect 408022 48698 443786 48934
rect 444022 48698 479786 48934
rect 480022 48698 515786 48934
rect 516022 48698 551786 48934
rect 552022 48698 591142 48934
rect 591378 48698 592500 48934
rect -8576 48676 592500 48698
rect -7636 48674 -7036 48676
rect 11604 48674 12204 48676
rect 47604 48674 48204 48676
rect 83604 48674 84204 48676
rect 119604 48674 120204 48676
rect 155604 48674 156204 48676
rect 191604 48674 192204 48676
rect 227604 48674 228204 48676
rect 263604 48674 264204 48676
rect 299604 48674 300204 48676
rect 335604 48674 336204 48676
rect 371604 48674 372204 48676
rect 407604 48674 408204 48676
rect 443604 48674 444204 48676
rect 479604 48674 480204 48676
rect 515604 48674 516204 48676
rect 551604 48674 552204 48676
rect 590960 48674 591560 48676
rect -5756 45676 -5156 45678
rect 8004 45676 8604 45678
rect 44004 45676 44604 45678
rect 80004 45676 80604 45678
rect 116004 45676 116604 45678
rect 152004 45676 152604 45678
rect 188004 45676 188604 45678
rect 224004 45676 224604 45678
rect 260004 45676 260604 45678
rect 296004 45676 296604 45678
rect 332004 45676 332604 45678
rect 368004 45676 368604 45678
rect 404004 45676 404604 45678
rect 440004 45676 440604 45678
rect 476004 45676 476604 45678
rect 512004 45676 512604 45678
rect 548004 45676 548604 45678
rect 589080 45676 589680 45678
rect -6696 45654 590620 45676
rect -6696 45418 -5574 45654
rect -5338 45418 8186 45654
rect 8422 45418 44186 45654
rect 44422 45418 80186 45654
rect 80422 45418 116186 45654
rect 116422 45418 152186 45654
rect 152422 45418 188186 45654
rect 188422 45418 224186 45654
rect 224422 45418 260186 45654
rect 260422 45418 296186 45654
rect 296422 45418 332186 45654
rect 332422 45418 368186 45654
rect 368422 45418 404186 45654
rect 404422 45418 440186 45654
rect 440422 45418 476186 45654
rect 476422 45418 512186 45654
rect 512422 45418 548186 45654
rect 548422 45418 589262 45654
rect 589498 45418 590620 45654
rect -6696 45334 590620 45418
rect -6696 45098 -5574 45334
rect -5338 45098 8186 45334
rect 8422 45098 44186 45334
rect 44422 45098 80186 45334
rect 80422 45098 116186 45334
rect 116422 45098 152186 45334
rect 152422 45098 188186 45334
rect 188422 45098 224186 45334
rect 224422 45098 260186 45334
rect 260422 45098 296186 45334
rect 296422 45098 332186 45334
rect 332422 45098 368186 45334
rect 368422 45098 404186 45334
rect 404422 45098 440186 45334
rect 440422 45098 476186 45334
rect 476422 45098 512186 45334
rect 512422 45098 548186 45334
rect 548422 45098 589262 45334
rect 589498 45098 590620 45334
rect -6696 45076 590620 45098
rect -5756 45074 -5156 45076
rect 8004 45074 8604 45076
rect 44004 45074 44604 45076
rect 80004 45074 80604 45076
rect 116004 45074 116604 45076
rect 152004 45074 152604 45076
rect 188004 45074 188604 45076
rect 224004 45074 224604 45076
rect 260004 45074 260604 45076
rect 296004 45074 296604 45076
rect 332004 45074 332604 45076
rect 368004 45074 368604 45076
rect 404004 45074 404604 45076
rect 440004 45074 440604 45076
rect 476004 45074 476604 45076
rect 512004 45074 512604 45076
rect 548004 45074 548604 45076
rect 589080 45074 589680 45076
rect -3876 42076 -3276 42078
rect 4404 42076 5004 42078
rect 40404 42076 41004 42078
rect 76404 42076 77004 42078
rect 112404 42076 113004 42078
rect 148404 42076 149004 42078
rect 184404 42076 185004 42078
rect 220404 42076 221004 42078
rect 256404 42076 257004 42078
rect 292404 42076 293004 42078
rect 328404 42076 329004 42078
rect 364404 42076 365004 42078
rect 400404 42076 401004 42078
rect 436404 42076 437004 42078
rect 472404 42076 473004 42078
rect 508404 42076 509004 42078
rect 544404 42076 545004 42078
rect 580404 42076 581004 42078
rect 587200 42076 587800 42078
rect -4816 42054 588740 42076
rect -4816 41818 -3694 42054
rect -3458 41818 4586 42054
rect 4822 41818 40586 42054
rect 40822 41818 76586 42054
rect 76822 41818 112586 42054
rect 112822 41818 148586 42054
rect 148822 41818 184586 42054
rect 184822 41818 220586 42054
rect 220822 41818 256586 42054
rect 256822 41818 292586 42054
rect 292822 41818 328586 42054
rect 328822 41818 364586 42054
rect 364822 41818 400586 42054
rect 400822 41818 436586 42054
rect 436822 41818 472586 42054
rect 472822 41818 508586 42054
rect 508822 41818 544586 42054
rect 544822 41818 580586 42054
rect 580822 41818 587382 42054
rect 587618 41818 588740 42054
rect -4816 41734 588740 41818
rect -4816 41498 -3694 41734
rect -3458 41498 4586 41734
rect 4822 41498 40586 41734
rect 40822 41498 76586 41734
rect 76822 41498 112586 41734
rect 112822 41498 148586 41734
rect 148822 41498 184586 41734
rect 184822 41498 220586 41734
rect 220822 41498 256586 41734
rect 256822 41498 292586 41734
rect 292822 41498 328586 41734
rect 328822 41498 364586 41734
rect 364822 41498 400586 41734
rect 400822 41498 436586 41734
rect 436822 41498 472586 41734
rect 472822 41498 508586 41734
rect 508822 41498 544586 41734
rect 544822 41498 580586 41734
rect 580822 41498 587382 41734
rect 587618 41498 588740 41734
rect -4816 41476 588740 41498
rect -3876 41474 -3276 41476
rect 4404 41474 5004 41476
rect 40404 41474 41004 41476
rect 76404 41474 77004 41476
rect 112404 41474 113004 41476
rect 148404 41474 149004 41476
rect 184404 41474 185004 41476
rect 220404 41474 221004 41476
rect 256404 41474 257004 41476
rect 292404 41474 293004 41476
rect 328404 41474 329004 41476
rect 364404 41474 365004 41476
rect 400404 41474 401004 41476
rect 436404 41474 437004 41476
rect 472404 41474 473004 41476
rect 508404 41474 509004 41476
rect 544404 41474 545004 41476
rect 580404 41474 581004 41476
rect 587200 41474 587800 41476
rect -1996 38476 -1396 38478
rect 804 38476 1404 38478
rect 36804 38476 37404 38478
rect 72804 38476 73404 38478
rect 108804 38476 109404 38478
rect 144804 38476 145404 38478
rect 180804 38476 181404 38478
rect 216804 38476 217404 38478
rect 252804 38476 253404 38478
rect 288804 38476 289404 38478
rect 324804 38476 325404 38478
rect 360804 38476 361404 38478
rect 396804 38476 397404 38478
rect 432804 38476 433404 38478
rect 468804 38476 469404 38478
rect 504804 38476 505404 38478
rect 540804 38476 541404 38478
rect 576804 38476 577404 38478
rect 585320 38476 585920 38478
rect -2936 38454 586860 38476
rect -2936 38218 -1814 38454
rect -1578 38218 986 38454
rect 1222 38218 36986 38454
rect 37222 38218 72986 38454
rect 73222 38218 108986 38454
rect 109222 38218 144986 38454
rect 145222 38218 180986 38454
rect 181222 38218 216986 38454
rect 217222 38218 252986 38454
rect 253222 38218 288986 38454
rect 289222 38218 324986 38454
rect 325222 38218 360986 38454
rect 361222 38218 396986 38454
rect 397222 38218 432986 38454
rect 433222 38218 468986 38454
rect 469222 38218 504986 38454
rect 505222 38218 540986 38454
rect 541222 38218 576986 38454
rect 577222 38218 585502 38454
rect 585738 38218 586860 38454
rect -2936 38134 586860 38218
rect -2936 37898 -1814 38134
rect -1578 37898 986 38134
rect 1222 37898 36986 38134
rect 37222 37898 72986 38134
rect 73222 37898 108986 38134
rect 109222 37898 144986 38134
rect 145222 37898 180986 38134
rect 181222 37898 216986 38134
rect 217222 37898 252986 38134
rect 253222 37898 288986 38134
rect 289222 37898 324986 38134
rect 325222 37898 360986 38134
rect 361222 37898 396986 38134
rect 397222 37898 432986 38134
rect 433222 37898 468986 38134
rect 469222 37898 504986 38134
rect 505222 37898 540986 38134
rect 541222 37898 576986 38134
rect 577222 37898 585502 38134
rect 585738 37898 586860 38134
rect -2936 37876 586860 37898
rect -1996 37874 -1396 37876
rect 804 37874 1404 37876
rect 36804 37874 37404 37876
rect 72804 37874 73404 37876
rect 108804 37874 109404 37876
rect 144804 37874 145404 37876
rect 180804 37874 181404 37876
rect 216804 37874 217404 37876
rect 252804 37874 253404 37876
rect 288804 37874 289404 37876
rect 324804 37874 325404 37876
rect 360804 37874 361404 37876
rect 396804 37874 397404 37876
rect 432804 37874 433404 37876
rect 468804 37874 469404 37876
rect 504804 37874 505404 37876
rect 540804 37874 541404 37876
rect 576804 37874 577404 37876
rect 585320 37874 585920 37876
rect -8576 31276 -7976 31278
rect 29604 31276 30204 31278
rect 65604 31276 66204 31278
rect 101604 31276 102204 31278
rect 137604 31276 138204 31278
rect 173604 31276 174204 31278
rect 209604 31276 210204 31278
rect 245604 31276 246204 31278
rect 281604 31276 282204 31278
rect 317604 31276 318204 31278
rect 353604 31276 354204 31278
rect 389604 31276 390204 31278
rect 425604 31276 426204 31278
rect 461604 31276 462204 31278
rect 497604 31276 498204 31278
rect 533604 31276 534204 31278
rect 569604 31276 570204 31278
rect 591900 31276 592500 31278
rect -8576 31254 592500 31276
rect -8576 31018 -8394 31254
rect -8158 31018 29786 31254
rect 30022 31018 65786 31254
rect 66022 31018 101786 31254
rect 102022 31018 137786 31254
rect 138022 31018 173786 31254
rect 174022 31018 209786 31254
rect 210022 31018 245786 31254
rect 246022 31018 281786 31254
rect 282022 31018 317786 31254
rect 318022 31018 353786 31254
rect 354022 31018 389786 31254
rect 390022 31018 425786 31254
rect 426022 31018 461786 31254
rect 462022 31018 497786 31254
rect 498022 31018 533786 31254
rect 534022 31018 569786 31254
rect 570022 31018 592082 31254
rect 592318 31018 592500 31254
rect -8576 30934 592500 31018
rect -8576 30698 -8394 30934
rect -8158 30698 29786 30934
rect 30022 30698 65786 30934
rect 66022 30698 101786 30934
rect 102022 30698 137786 30934
rect 138022 30698 173786 30934
rect 174022 30698 209786 30934
rect 210022 30698 245786 30934
rect 246022 30698 281786 30934
rect 282022 30698 317786 30934
rect 318022 30698 353786 30934
rect 354022 30698 389786 30934
rect 390022 30698 425786 30934
rect 426022 30698 461786 30934
rect 462022 30698 497786 30934
rect 498022 30698 533786 30934
rect 534022 30698 569786 30934
rect 570022 30698 592082 30934
rect 592318 30698 592500 30934
rect -8576 30676 592500 30698
rect -8576 30674 -7976 30676
rect 29604 30674 30204 30676
rect 65604 30674 66204 30676
rect 101604 30674 102204 30676
rect 137604 30674 138204 30676
rect 173604 30674 174204 30676
rect 209604 30674 210204 30676
rect 245604 30674 246204 30676
rect 281604 30674 282204 30676
rect 317604 30674 318204 30676
rect 353604 30674 354204 30676
rect 389604 30674 390204 30676
rect 425604 30674 426204 30676
rect 461604 30674 462204 30676
rect 497604 30674 498204 30676
rect 533604 30674 534204 30676
rect 569604 30674 570204 30676
rect 591900 30674 592500 30676
rect -6696 27676 -6096 27678
rect 26004 27676 26604 27678
rect 62004 27676 62604 27678
rect 98004 27676 98604 27678
rect 134004 27676 134604 27678
rect 170004 27676 170604 27678
rect 206004 27676 206604 27678
rect 242004 27676 242604 27678
rect 278004 27676 278604 27678
rect 314004 27676 314604 27678
rect 350004 27676 350604 27678
rect 386004 27676 386604 27678
rect 422004 27676 422604 27678
rect 458004 27676 458604 27678
rect 494004 27676 494604 27678
rect 530004 27676 530604 27678
rect 566004 27676 566604 27678
rect 590020 27676 590620 27678
rect -6696 27654 590620 27676
rect -6696 27418 -6514 27654
rect -6278 27418 26186 27654
rect 26422 27418 62186 27654
rect 62422 27418 98186 27654
rect 98422 27418 134186 27654
rect 134422 27418 170186 27654
rect 170422 27418 206186 27654
rect 206422 27418 242186 27654
rect 242422 27418 278186 27654
rect 278422 27418 314186 27654
rect 314422 27418 350186 27654
rect 350422 27418 386186 27654
rect 386422 27418 422186 27654
rect 422422 27418 458186 27654
rect 458422 27418 494186 27654
rect 494422 27418 530186 27654
rect 530422 27418 566186 27654
rect 566422 27418 590202 27654
rect 590438 27418 590620 27654
rect -6696 27334 590620 27418
rect -6696 27098 -6514 27334
rect -6278 27098 26186 27334
rect 26422 27098 62186 27334
rect 62422 27098 98186 27334
rect 98422 27098 134186 27334
rect 134422 27098 170186 27334
rect 170422 27098 206186 27334
rect 206422 27098 242186 27334
rect 242422 27098 278186 27334
rect 278422 27098 314186 27334
rect 314422 27098 350186 27334
rect 350422 27098 386186 27334
rect 386422 27098 422186 27334
rect 422422 27098 458186 27334
rect 458422 27098 494186 27334
rect 494422 27098 530186 27334
rect 530422 27098 566186 27334
rect 566422 27098 590202 27334
rect 590438 27098 590620 27334
rect -6696 27076 590620 27098
rect -6696 27074 -6096 27076
rect 26004 27074 26604 27076
rect 62004 27074 62604 27076
rect 98004 27074 98604 27076
rect 134004 27074 134604 27076
rect 170004 27074 170604 27076
rect 206004 27074 206604 27076
rect 242004 27074 242604 27076
rect 278004 27074 278604 27076
rect 314004 27074 314604 27076
rect 350004 27074 350604 27076
rect 386004 27074 386604 27076
rect 422004 27074 422604 27076
rect 458004 27074 458604 27076
rect 494004 27074 494604 27076
rect 530004 27074 530604 27076
rect 566004 27074 566604 27076
rect 590020 27074 590620 27076
rect -4816 24076 -4216 24078
rect 22404 24076 23004 24078
rect 58404 24076 59004 24078
rect 94404 24076 95004 24078
rect 130404 24076 131004 24078
rect 166404 24076 167004 24078
rect 202404 24076 203004 24078
rect 238404 24076 239004 24078
rect 274404 24076 275004 24078
rect 310404 24076 311004 24078
rect 346404 24076 347004 24078
rect 382404 24076 383004 24078
rect 418404 24076 419004 24078
rect 454404 24076 455004 24078
rect 490404 24076 491004 24078
rect 526404 24076 527004 24078
rect 562404 24076 563004 24078
rect 588140 24076 588740 24078
rect -4816 24054 588740 24076
rect -4816 23818 -4634 24054
rect -4398 23818 22586 24054
rect 22822 23818 58586 24054
rect 58822 23818 94586 24054
rect 94822 23818 130586 24054
rect 130822 23818 166586 24054
rect 166822 23818 202586 24054
rect 202822 23818 238586 24054
rect 238822 23818 274586 24054
rect 274822 23818 310586 24054
rect 310822 23818 346586 24054
rect 346822 23818 382586 24054
rect 382822 23818 418586 24054
rect 418822 23818 454586 24054
rect 454822 23818 490586 24054
rect 490822 23818 526586 24054
rect 526822 23818 562586 24054
rect 562822 23818 588322 24054
rect 588558 23818 588740 24054
rect -4816 23734 588740 23818
rect -4816 23498 -4634 23734
rect -4398 23498 22586 23734
rect 22822 23498 58586 23734
rect 58822 23498 94586 23734
rect 94822 23498 130586 23734
rect 130822 23498 166586 23734
rect 166822 23498 202586 23734
rect 202822 23498 238586 23734
rect 238822 23498 274586 23734
rect 274822 23498 310586 23734
rect 310822 23498 346586 23734
rect 346822 23498 382586 23734
rect 382822 23498 418586 23734
rect 418822 23498 454586 23734
rect 454822 23498 490586 23734
rect 490822 23498 526586 23734
rect 526822 23498 562586 23734
rect 562822 23498 588322 23734
rect 588558 23498 588740 23734
rect -4816 23476 588740 23498
rect -4816 23474 -4216 23476
rect 22404 23474 23004 23476
rect 58404 23474 59004 23476
rect 94404 23474 95004 23476
rect 130404 23474 131004 23476
rect 166404 23474 167004 23476
rect 202404 23474 203004 23476
rect 238404 23474 239004 23476
rect 274404 23474 275004 23476
rect 310404 23474 311004 23476
rect 346404 23474 347004 23476
rect 382404 23474 383004 23476
rect 418404 23474 419004 23476
rect 454404 23474 455004 23476
rect 490404 23474 491004 23476
rect 526404 23474 527004 23476
rect 562404 23474 563004 23476
rect 588140 23474 588740 23476
rect -2936 20476 -2336 20478
rect 18804 20476 19404 20478
rect 54804 20476 55404 20478
rect 90804 20476 91404 20478
rect 126804 20476 127404 20478
rect 162804 20476 163404 20478
rect 198804 20476 199404 20478
rect 234804 20476 235404 20478
rect 270804 20476 271404 20478
rect 306804 20476 307404 20478
rect 342804 20476 343404 20478
rect 378804 20476 379404 20478
rect 414804 20476 415404 20478
rect 450804 20476 451404 20478
rect 486804 20476 487404 20478
rect 522804 20476 523404 20478
rect 558804 20476 559404 20478
rect 586260 20476 586860 20478
rect -2936 20454 586860 20476
rect -2936 20218 -2754 20454
rect -2518 20218 18986 20454
rect 19222 20218 54986 20454
rect 55222 20218 90986 20454
rect 91222 20218 126986 20454
rect 127222 20218 162986 20454
rect 163222 20218 198986 20454
rect 199222 20218 234986 20454
rect 235222 20218 270986 20454
rect 271222 20218 306986 20454
rect 307222 20218 342986 20454
rect 343222 20218 378986 20454
rect 379222 20218 414986 20454
rect 415222 20218 450986 20454
rect 451222 20218 486986 20454
rect 487222 20218 522986 20454
rect 523222 20218 558986 20454
rect 559222 20218 586442 20454
rect 586678 20218 586860 20454
rect -2936 20134 586860 20218
rect -2936 19898 -2754 20134
rect -2518 19898 18986 20134
rect 19222 19898 54986 20134
rect 55222 19898 90986 20134
rect 91222 19898 126986 20134
rect 127222 19898 162986 20134
rect 163222 19898 198986 20134
rect 199222 19898 234986 20134
rect 235222 19898 270986 20134
rect 271222 19898 306986 20134
rect 307222 19898 342986 20134
rect 343222 19898 378986 20134
rect 379222 19898 414986 20134
rect 415222 19898 450986 20134
rect 451222 19898 486986 20134
rect 487222 19898 522986 20134
rect 523222 19898 558986 20134
rect 559222 19898 586442 20134
rect 586678 19898 586860 20134
rect -2936 19876 586860 19898
rect -2936 19874 -2336 19876
rect 18804 19874 19404 19876
rect 54804 19874 55404 19876
rect 90804 19874 91404 19876
rect 126804 19874 127404 19876
rect 162804 19874 163404 19876
rect 198804 19874 199404 19876
rect 234804 19874 235404 19876
rect 270804 19874 271404 19876
rect 306804 19874 307404 19876
rect 342804 19874 343404 19876
rect 378804 19874 379404 19876
rect 414804 19874 415404 19876
rect 450804 19874 451404 19876
rect 486804 19874 487404 19876
rect 522804 19874 523404 19876
rect 558804 19874 559404 19876
rect 586260 19874 586860 19876
rect -7636 13276 -7036 13278
rect 11604 13276 12204 13278
rect 47604 13276 48204 13278
rect 83604 13276 84204 13278
rect 119604 13276 120204 13278
rect 155604 13276 156204 13278
rect 191604 13276 192204 13278
rect 227604 13276 228204 13278
rect 263604 13276 264204 13278
rect 299604 13276 300204 13278
rect 335604 13276 336204 13278
rect 371604 13276 372204 13278
rect 407604 13276 408204 13278
rect 443604 13276 444204 13278
rect 479604 13276 480204 13278
rect 515604 13276 516204 13278
rect 551604 13276 552204 13278
rect 590960 13276 591560 13278
rect -8576 13254 592500 13276
rect -8576 13018 -7454 13254
rect -7218 13018 11786 13254
rect 12022 13018 47786 13254
rect 48022 13018 83786 13254
rect 84022 13018 119786 13254
rect 120022 13018 155786 13254
rect 156022 13018 191786 13254
rect 192022 13018 227786 13254
rect 228022 13018 263786 13254
rect 264022 13018 299786 13254
rect 300022 13018 335786 13254
rect 336022 13018 371786 13254
rect 372022 13018 407786 13254
rect 408022 13018 443786 13254
rect 444022 13018 479786 13254
rect 480022 13018 515786 13254
rect 516022 13018 551786 13254
rect 552022 13018 591142 13254
rect 591378 13018 592500 13254
rect -8576 12934 592500 13018
rect -8576 12698 -7454 12934
rect -7218 12698 11786 12934
rect 12022 12698 47786 12934
rect 48022 12698 83786 12934
rect 84022 12698 119786 12934
rect 120022 12698 155786 12934
rect 156022 12698 191786 12934
rect 192022 12698 227786 12934
rect 228022 12698 263786 12934
rect 264022 12698 299786 12934
rect 300022 12698 335786 12934
rect 336022 12698 371786 12934
rect 372022 12698 407786 12934
rect 408022 12698 443786 12934
rect 444022 12698 479786 12934
rect 480022 12698 515786 12934
rect 516022 12698 551786 12934
rect 552022 12698 591142 12934
rect 591378 12698 592500 12934
rect -8576 12676 592500 12698
rect -7636 12674 -7036 12676
rect 11604 12674 12204 12676
rect 47604 12674 48204 12676
rect 83604 12674 84204 12676
rect 119604 12674 120204 12676
rect 155604 12674 156204 12676
rect 191604 12674 192204 12676
rect 227604 12674 228204 12676
rect 263604 12674 264204 12676
rect 299604 12674 300204 12676
rect 335604 12674 336204 12676
rect 371604 12674 372204 12676
rect 407604 12674 408204 12676
rect 443604 12674 444204 12676
rect 479604 12674 480204 12676
rect 515604 12674 516204 12676
rect 551604 12674 552204 12676
rect 590960 12674 591560 12676
rect -5756 9676 -5156 9678
rect 8004 9676 8604 9678
rect 44004 9676 44604 9678
rect 80004 9676 80604 9678
rect 116004 9676 116604 9678
rect 152004 9676 152604 9678
rect 188004 9676 188604 9678
rect 224004 9676 224604 9678
rect 260004 9676 260604 9678
rect 296004 9676 296604 9678
rect 332004 9676 332604 9678
rect 368004 9676 368604 9678
rect 404004 9676 404604 9678
rect 440004 9676 440604 9678
rect 476004 9676 476604 9678
rect 512004 9676 512604 9678
rect 548004 9676 548604 9678
rect 589080 9676 589680 9678
rect -6696 9654 590620 9676
rect -6696 9418 -5574 9654
rect -5338 9418 8186 9654
rect 8422 9418 44186 9654
rect 44422 9418 80186 9654
rect 80422 9418 116186 9654
rect 116422 9418 152186 9654
rect 152422 9418 188186 9654
rect 188422 9418 224186 9654
rect 224422 9418 260186 9654
rect 260422 9418 296186 9654
rect 296422 9418 332186 9654
rect 332422 9418 368186 9654
rect 368422 9418 404186 9654
rect 404422 9418 440186 9654
rect 440422 9418 476186 9654
rect 476422 9418 512186 9654
rect 512422 9418 548186 9654
rect 548422 9418 589262 9654
rect 589498 9418 590620 9654
rect -6696 9334 590620 9418
rect -6696 9098 -5574 9334
rect -5338 9098 8186 9334
rect 8422 9098 44186 9334
rect 44422 9098 80186 9334
rect 80422 9098 116186 9334
rect 116422 9098 152186 9334
rect 152422 9098 188186 9334
rect 188422 9098 224186 9334
rect 224422 9098 260186 9334
rect 260422 9098 296186 9334
rect 296422 9098 332186 9334
rect 332422 9098 368186 9334
rect 368422 9098 404186 9334
rect 404422 9098 440186 9334
rect 440422 9098 476186 9334
rect 476422 9098 512186 9334
rect 512422 9098 548186 9334
rect 548422 9098 589262 9334
rect 589498 9098 590620 9334
rect -6696 9076 590620 9098
rect -5756 9074 -5156 9076
rect 8004 9074 8604 9076
rect 44004 9074 44604 9076
rect 80004 9074 80604 9076
rect 116004 9074 116604 9076
rect 152004 9074 152604 9076
rect 188004 9074 188604 9076
rect 224004 9074 224604 9076
rect 260004 9074 260604 9076
rect 296004 9074 296604 9076
rect 332004 9074 332604 9076
rect 368004 9074 368604 9076
rect 404004 9074 404604 9076
rect 440004 9074 440604 9076
rect 476004 9074 476604 9076
rect 512004 9074 512604 9076
rect 548004 9074 548604 9076
rect 589080 9074 589680 9076
rect -3876 6076 -3276 6078
rect 4404 6076 5004 6078
rect 40404 6076 41004 6078
rect 76404 6076 77004 6078
rect 112404 6076 113004 6078
rect 148404 6076 149004 6078
rect 184404 6076 185004 6078
rect 220404 6076 221004 6078
rect 256404 6076 257004 6078
rect 292404 6076 293004 6078
rect 328404 6076 329004 6078
rect 364404 6076 365004 6078
rect 400404 6076 401004 6078
rect 436404 6076 437004 6078
rect 472404 6076 473004 6078
rect 508404 6076 509004 6078
rect 544404 6076 545004 6078
rect 580404 6076 581004 6078
rect 587200 6076 587800 6078
rect -4816 6054 588740 6076
rect -4816 5818 -3694 6054
rect -3458 5818 4586 6054
rect 4822 5818 40586 6054
rect 40822 5818 76586 6054
rect 76822 5818 112586 6054
rect 112822 5818 148586 6054
rect 148822 5818 184586 6054
rect 184822 5818 220586 6054
rect 220822 5818 256586 6054
rect 256822 5818 292586 6054
rect 292822 5818 328586 6054
rect 328822 5818 364586 6054
rect 364822 5818 400586 6054
rect 400822 5818 436586 6054
rect 436822 5818 472586 6054
rect 472822 5818 508586 6054
rect 508822 5818 544586 6054
rect 544822 5818 580586 6054
rect 580822 5818 587382 6054
rect 587618 5818 588740 6054
rect -4816 5734 588740 5818
rect -4816 5498 -3694 5734
rect -3458 5498 4586 5734
rect 4822 5498 40586 5734
rect 40822 5498 76586 5734
rect 76822 5498 112586 5734
rect 112822 5498 148586 5734
rect 148822 5498 184586 5734
rect 184822 5498 220586 5734
rect 220822 5498 256586 5734
rect 256822 5498 292586 5734
rect 292822 5498 328586 5734
rect 328822 5498 364586 5734
rect 364822 5498 400586 5734
rect 400822 5498 436586 5734
rect 436822 5498 472586 5734
rect 472822 5498 508586 5734
rect 508822 5498 544586 5734
rect 544822 5498 580586 5734
rect 580822 5498 587382 5734
rect 587618 5498 588740 5734
rect -4816 5476 588740 5498
rect -3876 5474 -3276 5476
rect 4404 5474 5004 5476
rect 40404 5474 41004 5476
rect 76404 5474 77004 5476
rect 112404 5474 113004 5476
rect 148404 5474 149004 5476
rect 184404 5474 185004 5476
rect 220404 5474 221004 5476
rect 256404 5474 257004 5476
rect 292404 5474 293004 5476
rect 328404 5474 329004 5476
rect 364404 5474 365004 5476
rect 400404 5474 401004 5476
rect 436404 5474 437004 5476
rect 472404 5474 473004 5476
rect 508404 5474 509004 5476
rect 544404 5474 545004 5476
rect 580404 5474 581004 5476
rect 587200 5474 587800 5476
rect -1996 2476 -1396 2478
rect 804 2476 1404 2478
rect 36804 2476 37404 2478
rect 72804 2476 73404 2478
rect 108804 2476 109404 2478
rect 144804 2476 145404 2478
rect 180804 2476 181404 2478
rect 216804 2476 217404 2478
rect 252804 2476 253404 2478
rect 288804 2476 289404 2478
rect 324804 2476 325404 2478
rect 360804 2476 361404 2478
rect 396804 2476 397404 2478
rect 432804 2476 433404 2478
rect 468804 2476 469404 2478
rect 504804 2476 505404 2478
rect 540804 2476 541404 2478
rect 576804 2476 577404 2478
rect 585320 2476 585920 2478
rect -2936 2454 586860 2476
rect -2936 2218 -1814 2454
rect -1578 2218 986 2454
rect 1222 2218 36986 2454
rect 37222 2218 72986 2454
rect 73222 2218 108986 2454
rect 109222 2218 144986 2454
rect 145222 2218 180986 2454
rect 181222 2218 216986 2454
rect 217222 2218 252986 2454
rect 253222 2218 288986 2454
rect 289222 2218 324986 2454
rect 325222 2218 360986 2454
rect 361222 2218 396986 2454
rect 397222 2218 432986 2454
rect 433222 2218 468986 2454
rect 469222 2218 504986 2454
rect 505222 2218 540986 2454
rect 541222 2218 576986 2454
rect 577222 2218 585502 2454
rect 585738 2218 586860 2454
rect -2936 2134 586860 2218
rect -2936 1898 -1814 2134
rect -1578 1898 986 2134
rect 1222 1898 36986 2134
rect 37222 1898 72986 2134
rect 73222 1898 108986 2134
rect 109222 1898 144986 2134
rect 145222 1898 180986 2134
rect 181222 1898 216986 2134
rect 217222 1898 252986 2134
rect 253222 1898 288986 2134
rect 289222 1898 324986 2134
rect 325222 1898 360986 2134
rect 361222 1898 396986 2134
rect 397222 1898 432986 2134
rect 433222 1898 468986 2134
rect 469222 1898 504986 2134
rect 505222 1898 540986 2134
rect 541222 1898 576986 2134
rect 577222 1898 585502 2134
rect 585738 1898 586860 2134
rect -2936 1876 586860 1898
rect -1996 1874 -1396 1876
rect 804 1874 1404 1876
rect 36804 1874 37404 1876
rect 72804 1874 73404 1876
rect 108804 1874 109404 1876
rect 144804 1874 145404 1876
rect 180804 1874 181404 1876
rect 216804 1874 217404 1876
rect 252804 1874 253404 1876
rect 288804 1874 289404 1876
rect 324804 1874 325404 1876
rect 360804 1874 361404 1876
rect 396804 1874 397404 1876
rect 432804 1874 433404 1876
rect 468804 1874 469404 1876
rect 504804 1874 505404 1876
rect 540804 1874 541404 1876
rect 576804 1874 577404 1876
rect 585320 1874 585920 1876
rect -1996 -324 -1396 -322
rect 804 -324 1404 -322
rect 36804 -324 37404 -322
rect 72804 -324 73404 -322
rect 108804 -324 109404 -322
rect 144804 -324 145404 -322
rect 180804 -324 181404 -322
rect 216804 -324 217404 -322
rect 252804 -324 253404 -322
rect 288804 -324 289404 -322
rect 324804 -324 325404 -322
rect 360804 -324 361404 -322
rect 396804 -324 397404 -322
rect 432804 -324 433404 -322
rect 468804 -324 469404 -322
rect 504804 -324 505404 -322
rect 540804 -324 541404 -322
rect 576804 -324 577404 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 986 -346
rect 1222 -582 36986 -346
rect 37222 -582 72986 -346
rect 73222 -582 108986 -346
rect 109222 -582 144986 -346
rect 145222 -582 180986 -346
rect 181222 -582 216986 -346
rect 217222 -582 252986 -346
rect 253222 -582 288986 -346
rect 289222 -582 324986 -346
rect 325222 -582 360986 -346
rect 361222 -582 396986 -346
rect 397222 -582 432986 -346
rect 433222 -582 468986 -346
rect 469222 -582 504986 -346
rect 505222 -582 540986 -346
rect 541222 -582 576986 -346
rect 577222 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 986 -666
rect 1222 -902 36986 -666
rect 37222 -902 72986 -666
rect 73222 -902 108986 -666
rect 109222 -902 144986 -666
rect 145222 -902 180986 -666
rect 181222 -902 216986 -666
rect 217222 -902 252986 -666
rect 253222 -902 288986 -666
rect 289222 -902 324986 -666
rect 325222 -902 360986 -666
rect 361222 -902 396986 -666
rect 397222 -902 432986 -666
rect 433222 -902 468986 -666
rect 469222 -902 504986 -666
rect 505222 -902 540986 -666
rect 541222 -902 576986 -666
rect 577222 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 108804 -926 109404 -924
rect 144804 -926 145404 -924
rect 180804 -926 181404 -924
rect 216804 -926 217404 -924
rect 252804 -926 253404 -924
rect 288804 -926 289404 -924
rect 324804 -926 325404 -924
rect 360804 -926 361404 -924
rect 396804 -926 397404 -924
rect 432804 -926 433404 -924
rect 468804 -926 469404 -924
rect 504804 -926 505404 -924
rect 540804 -926 541404 -924
rect 576804 -926 577404 -924
rect 585320 -926 585920 -924
rect -2936 -1264 -2336 -1262
rect 18804 -1264 19404 -1262
rect 54804 -1264 55404 -1262
rect 90804 -1264 91404 -1262
rect 126804 -1264 127404 -1262
rect 162804 -1264 163404 -1262
rect 198804 -1264 199404 -1262
rect 234804 -1264 235404 -1262
rect 270804 -1264 271404 -1262
rect 306804 -1264 307404 -1262
rect 342804 -1264 343404 -1262
rect 378804 -1264 379404 -1262
rect 414804 -1264 415404 -1262
rect 450804 -1264 451404 -1262
rect 486804 -1264 487404 -1262
rect 522804 -1264 523404 -1262
rect 558804 -1264 559404 -1262
rect 586260 -1264 586860 -1262
rect -2936 -1286 586860 -1264
rect -2936 -1522 -2754 -1286
rect -2518 -1522 18986 -1286
rect 19222 -1522 54986 -1286
rect 55222 -1522 90986 -1286
rect 91222 -1522 126986 -1286
rect 127222 -1522 162986 -1286
rect 163222 -1522 198986 -1286
rect 199222 -1522 234986 -1286
rect 235222 -1522 270986 -1286
rect 271222 -1522 306986 -1286
rect 307222 -1522 342986 -1286
rect 343222 -1522 378986 -1286
rect 379222 -1522 414986 -1286
rect 415222 -1522 450986 -1286
rect 451222 -1522 486986 -1286
rect 487222 -1522 522986 -1286
rect 523222 -1522 558986 -1286
rect 559222 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect -2936 -1606 586860 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 18986 -1606
rect 19222 -1842 54986 -1606
rect 55222 -1842 90986 -1606
rect 91222 -1842 126986 -1606
rect 127222 -1842 162986 -1606
rect 163222 -1842 198986 -1606
rect 199222 -1842 234986 -1606
rect 235222 -1842 270986 -1606
rect 271222 -1842 306986 -1606
rect 307222 -1842 342986 -1606
rect 343222 -1842 378986 -1606
rect 379222 -1842 414986 -1606
rect 415222 -1842 450986 -1606
rect 451222 -1842 486986 -1606
rect 487222 -1842 522986 -1606
rect 523222 -1842 558986 -1606
rect 559222 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect -2936 -1864 586860 -1842
rect -2936 -1866 -2336 -1864
rect 18804 -1866 19404 -1864
rect 54804 -1866 55404 -1864
rect 90804 -1866 91404 -1864
rect 126804 -1866 127404 -1864
rect 162804 -1866 163404 -1864
rect 198804 -1866 199404 -1864
rect 234804 -1866 235404 -1864
rect 270804 -1866 271404 -1864
rect 306804 -1866 307404 -1864
rect 342804 -1866 343404 -1864
rect 378804 -1866 379404 -1864
rect 414804 -1866 415404 -1864
rect 450804 -1866 451404 -1864
rect 486804 -1866 487404 -1864
rect 522804 -1866 523404 -1864
rect 558804 -1866 559404 -1864
rect 586260 -1866 586860 -1864
rect -3876 -2204 -3276 -2202
rect 4404 -2204 5004 -2202
rect 40404 -2204 41004 -2202
rect 76404 -2204 77004 -2202
rect 112404 -2204 113004 -2202
rect 148404 -2204 149004 -2202
rect 184404 -2204 185004 -2202
rect 220404 -2204 221004 -2202
rect 256404 -2204 257004 -2202
rect 292404 -2204 293004 -2202
rect 328404 -2204 329004 -2202
rect 364404 -2204 365004 -2202
rect 400404 -2204 401004 -2202
rect 436404 -2204 437004 -2202
rect 472404 -2204 473004 -2202
rect 508404 -2204 509004 -2202
rect 544404 -2204 545004 -2202
rect 580404 -2204 581004 -2202
rect 587200 -2204 587800 -2202
rect -3876 -2226 587800 -2204
rect -3876 -2462 -3694 -2226
rect -3458 -2462 4586 -2226
rect 4822 -2462 40586 -2226
rect 40822 -2462 76586 -2226
rect 76822 -2462 112586 -2226
rect 112822 -2462 148586 -2226
rect 148822 -2462 184586 -2226
rect 184822 -2462 220586 -2226
rect 220822 -2462 256586 -2226
rect 256822 -2462 292586 -2226
rect 292822 -2462 328586 -2226
rect 328822 -2462 364586 -2226
rect 364822 -2462 400586 -2226
rect 400822 -2462 436586 -2226
rect 436822 -2462 472586 -2226
rect 472822 -2462 508586 -2226
rect 508822 -2462 544586 -2226
rect 544822 -2462 580586 -2226
rect 580822 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect -3876 -2546 587800 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 4586 -2546
rect 4822 -2782 40586 -2546
rect 40822 -2782 76586 -2546
rect 76822 -2782 112586 -2546
rect 112822 -2782 148586 -2546
rect 148822 -2782 184586 -2546
rect 184822 -2782 220586 -2546
rect 220822 -2782 256586 -2546
rect 256822 -2782 292586 -2546
rect 292822 -2782 328586 -2546
rect 328822 -2782 364586 -2546
rect 364822 -2782 400586 -2546
rect 400822 -2782 436586 -2546
rect 436822 -2782 472586 -2546
rect 472822 -2782 508586 -2546
rect 508822 -2782 544586 -2546
rect 544822 -2782 580586 -2546
rect 580822 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect -3876 -2804 587800 -2782
rect -3876 -2806 -3276 -2804
rect 4404 -2806 5004 -2804
rect 40404 -2806 41004 -2804
rect 76404 -2806 77004 -2804
rect 112404 -2806 113004 -2804
rect 148404 -2806 149004 -2804
rect 184404 -2806 185004 -2804
rect 220404 -2806 221004 -2804
rect 256404 -2806 257004 -2804
rect 292404 -2806 293004 -2804
rect 328404 -2806 329004 -2804
rect 364404 -2806 365004 -2804
rect 400404 -2806 401004 -2804
rect 436404 -2806 437004 -2804
rect 472404 -2806 473004 -2804
rect 508404 -2806 509004 -2804
rect 544404 -2806 545004 -2804
rect 580404 -2806 581004 -2804
rect 587200 -2806 587800 -2804
rect -4816 -3144 -4216 -3142
rect 22404 -3144 23004 -3142
rect 58404 -3144 59004 -3142
rect 94404 -3144 95004 -3142
rect 130404 -3144 131004 -3142
rect 166404 -3144 167004 -3142
rect 202404 -3144 203004 -3142
rect 238404 -3144 239004 -3142
rect 274404 -3144 275004 -3142
rect 310404 -3144 311004 -3142
rect 346404 -3144 347004 -3142
rect 382404 -3144 383004 -3142
rect 418404 -3144 419004 -3142
rect 454404 -3144 455004 -3142
rect 490404 -3144 491004 -3142
rect 526404 -3144 527004 -3142
rect 562404 -3144 563004 -3142
rect 588140 -3144 588740 -3142
rect -4816 -3166 588740 -3144
rect -4816 -3402 -4634 -3166
rect -4398 -3402 22586 -3166
rect 22822 -3402 58586 -3166
rect 58822 -3402 94586 -3166
rect 94822 -3402 130586 -3166
rect 130822 -3402 166586 -3166
rect 166822 -3402 202586 -3166
rect 202822 -3402 238586 -3166
rect 238822 -3402 274586 -3166
rect 274822 -3402 310586 -3166
rect 310822 -3402 346586 -3166
rect 346822 -3402 382586 -3166
rect 382822 -3402 418586 -3166
rect 418822 -3402 454586 -3166
rect 454822 -3402 490586 -3166
rect 490822 -3402 526586 -3166
rect 526822 -3402 562586 -3166
rect 562822 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect -4816 -3486 588740 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 22586 -3486
rect 22822 -3722 58586 -3486
rect 58822 -3722 94586 -3486
rect 94822 -3722 130586 -3486
rect 130822 -3722 166586 -3486
rect 166822 -3722 202586 -3486
rect 202822 -3722 238586 -3486
rect 238822 -3722 274586 -3486
rect 274822 -3722 310586 -3486
rect 310822 -3722 346586 -3486
rect 346822 -3722 382586 -3486
rect 382822 -3722 418586 -3486
rect 418822 -3722 454586 -3486
rect 454822 -3722 490586 -3486
rect 490822 -3722 526586 -3486
rect 526822 -3722 562586 -3486
rect 562822 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect -4816 -3744 588740 -3722
rect -4816 -3746 -4216 -3744
rect 22404 -3746 23004 -3744
rect 58404 -3746 59004 -3744
rect 94404 -3746 95004 -3744
rect 130404 -3746 131004 -3744
rect 166404 -3746 167004 -3744
rect 202404 -3746 203004 -3744
rect 238404 -3746 239004 -3744
rect 274404 -3746 275004 -3744
rect 310404 -3746 311004 -3744
rect 346404 -3746 347004 -3744
rect 382404 -3746 383004 -3744
rect 418404 -3746 419004 -3744
rect 454404 -3746 455004 -3744
rect 490404 -3746 491004 -3744
rect 526404 -3746 527004 -3744
rect 562404 -3746 563004 -3744
rect 588140 -3746 588740 -3744
rect -5756 -4084 -5156 -4082
rect 8004 -4084 8604 -4082
rect 44004 -4084 44604 -4082
rect 80004 -4084 80604 -4082
rect 116004 -4084 116604 -4082
rect 152004 -4084 152604 -4082
rect 188004 -4084 188604 -4082
rect 224004 -4084 224604 -4082
rect 260004 -4084 260604 -4082
rect 296004 -4084 296604 -4082
rect 332004 -4084 332604 -4082
rect 368004 -4084 368604 -4082
rect 404004 -4084 404604 -4082
rect 440004 -4084 440604 -4082
rect 476004 -4084 476604 -4082
rect 512004 -4084 512604 -4082
rect 548004 -4084 548604 -4082
rect 589080 -4084 589680 -4082
rect -5756 -4106 589680 -4084
rect -5756 -4342 -5574 -4106
rect -5338 -4342 8186 -4106
rect 8422 -4342 44186 -4106
rect 44422 -4342 80186 -4106
rect 80422 -4342 116186 -4106
rect 116422 -4342 152186 -4106
rect 152422 -4342 188186 -4106
rect 188422 -4342 224186 -4106
rect 224422 -4342 260186 -4106
rect 260422 -4342 296186 -4106
rect 296422 -4342 332186 -4106
rect 332422 -4342 368186 -4106
rect 368422 -4342 404186 -4106
rect 404422 -4342 440186 -4106
rect 440422 -4342 476186 -4106
rect 476422 -4342 512186 -4106
rect 512422 -4342 548186 -4106
rect 548422 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect -5756 -4426 589680 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 8186 -4426
rect 8422 -4662 44186 -4426
rect 44422 -4662 80186 -4426
rect 80422 -4662 116186 -4426
rect 116422 -4662 152186 -4426
rect 152422 -4662 188186 -4426
rect 188422 -4662 224186 -4426
rect 224422 -4662 260186 -4426
rect 260422 -4662 296186 -4426
rect 296422 -4662 332186 -4426
rect 332422 -4662 368186 -4426
rect 368422 -4662 404186 -4426
rect 404422 -4662 440186 -4426
rect 440422 -4662 476186 -4426
rect 476422 -4662 512186 -4426
rect 512422 -4662 548186 -4426
rect 548422 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect -5756 -4684 589680 -4662
rect -5756 -4686 -5156 -4684
rect 8004 -4686 8604 -4684
rect 44004 -4686 44604 -4684
rect 80004 -4686 80604 -4684
rect 116004 -4686 116604 -4684
rect 152004 -4686 152604 -4684
rect 188004 -4686 188604 -4684
rect 224004 -4686 224604 -4684
rect 260004 -4686 260604 -4684
rect 296004 -4686 296604 -4684
rect 332004 -4686 332604 -4684
rect 368004 -4686 368604 -4684
rect 404004 -4686 404604 -4684
rect 440004 -4686 440604 -4684
rect 476004 -4686 476604 -4684
rect 512004 -4686 512604 -4684
rect 548004 -4686 548604 -4684
rect 589080 -4686 589680 -4684
rect -6696 -5024 -6096 -5022
rect 26004 -5024 26604 -5022
rect 62004 -5024 62604 -5022
rect 98004 -5024 98604 -5022
rect 134004 -5024 134604 -5022
rect 170004 -5024 170604 -5022
rect 206004 -5024 206604 -5022
rect 242004 -5024 242604 -5022
rect 278004 -5024 278604 -5022
rect 314004 -5024 314604 -5022
rect 350004 -5024 350604 -5022
rect 386004 -5024 386604 -5022
rect 422004 -5024 422604 -5022
rect 458004 -5024 458604 -5022
rect 494004 -5024 494604 -5022
rect 530004 -5024 530604 -5022
rect 566004 -5024 566604 -5022
rect 590020 -5024 590620 -5022
rect -6696 -5046 590620 -5024
rect -6696 -5282 -6514 -5046
rect -6278 -5282 26186 -5046
rect 26422 -5282 62186 -5046
rect 62422 -5282 98186 -5046
rect 98422 -5282 134186 -5046
rect 134422 -5282 170186 -5046
rect 170422 -5282 206186 -5046
rect 206422 -5282 242186 -5046
rect 242422 -5282 278186 -5046
rect 278422 -5282 314186 -5046
rect 314422 -5282 350186 -5046
rect 350422 -5282 386186 -5046
rect 386422 -5282 422186 -5046
rect 422422 -5282 458186 -5046
rect 458422 -5282 494186 -5046
rect 494422 -5282 530186 -5046
rect 530422 -5282 566186 -5046
rect 566422 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect -6696 -5366 590620 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 26186 -5366
rect 26422 -5602 62186 -5366
rect 62422 -5602 98186 -5366
rect 98422 -5602 134186 -5366
rect 134422 -5602 170186 -5366
rect 170422 -5602 206186 -5366
rect 206422 -5602 242186 -5366
rect 242422 -5602 278186 -5366
rect 278422 -5602 314186 -5366
rect 314422 -5602 350186 -5366
rect 350422 -5602 386186 -5366
rect 386422 -5602 422186 -5366
rect 422422 -5602 458186 -5366
rect 458422 -5602 494186 -5366
rect 494422 -5602 530186 -5366
rect 530422 -5602 566186 -5366
rect 566422 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect -6696 -5624 590620 -5602
rect -6696 -5626 -6096 -5624
rect 26004 -5626 26604 -5624
rect 62004 -5626 62604 -5624
rect 98004 -5626 98604 -5624
rect 134004 -5626 134604 -5624
rect 170004 -5626 170604 -5624
rect 206004 -5626 206604 -5624
rect 242004 -5626 242604 -5624
rect 278004 -5626 278604 -5624
rect 314004 -5626 314604 -5624
rect 350004 -5626 350604 -5624
rect 386004 -5626 386604 -5624
rect 422004 -5626 422604 -5624
rect 458004 -5626 458604 -5624
rect 494004 -5626 494604 -5624
rect 530004 -5626 530604 -5624
rect 566004 -5626 566604 -5624
rect 590020 -5626 590620 -5624
rect -7636 -5964 -7036 -5962
rect 11604 -5964 12204 -5962
rect 47604 -5964 48204 -5962
rect 83604 -5964 84204 -5962
rect 119604 -5964 120204 -5962
rect 155604 -5964 156204 -5962
rect 191604 -5964 192204 -5962
rect 227604 -5964 228204 -5962
rect 263604 -5964 264204 -5962
rect 299604 -5964 300204 -5962
rect 335604 -5964 336204 -5962
rect 371604 -5964 372204 -5962
rect 407604 -5964 408204 -5962
rect 443604 -5964 444204 -5962
rect 479604 -5964 480204 -5962
rect 515604 -5964 516204 -5962
rect 551604 -5964 552204 -5962
rect 590960 -5964 591560 -5962
rect -7636 -5986 591560 -5964
rect -7636 -6222 -7454 -5986
rect -7218 -6222 11786 -5986
rect 12022 -6222 47786 -5986
rect 48022 -6222 83786 -5986
rect 84022 -6222 119786 -5986
rect 120022 -6222 155786 -5986
rect 156022 -6222 191786 -5986
rect 192022 -6222 227786 -5986
rect 228022 -6222 263786 -5986
rect 264022 -6222 299786 -5986
rect 300022 -6222 335786 -5986
rect 336022 -6222 371786 -5986
rect 372022 -6222 407786 -5986
rect 408022 -6222 443786 -5986
rect 444022 -6222 479786 -5986
rect 480022 -6222 515786 -5986
rect 516022 -6222 551786 -5986
rect 552022 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect -7636 -6306 591560 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 11786 -6306
rect 12022 -6542 47786 -6306
rect 48022 -6542 83786 -6306
rect 84022 -6542 119786 -6306
rect 120022 -6542 155786 -6306
rect 156022 -6542 191786 -6306
rect 192022 -6542 227786 -6306
rect 228022 -6542 263786 -6306
rect 264022 -6542 299786 -6306
rect 300022 -6542 335786 -6306
rect 336022 -6542 371786 -6306
rect 372022 -6542 407786 -6306
rect 408022 -6542 443786 -6306
rect 444022 -6542 479786 -6306
rect 480022 -6542 515786 -6306
rect 516022 -6542 551786 -6306
rect 552022 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect -7636 -6564 591560 -6542
rect -7636 -6566 -7036 -6564
rect 11604 -6566 12204 -6564
rect 47604 -6566 48204 -6564
rect 83604 -6566 84204 -6564
rect 119604 -6566 120204 -6564
rect 155604 -6566 156204 -6564
rect 191604 -6566 192204 -6564
rect 227604 -6566 228204 -6564
rect 263604 -6566 264204 -6564
rect 299604 -6566 300204 -6564
rect 335604 -6566 336204 -6564
rect 371604 -6566 372204 -6564
rect 407604 -6566 408204 -6564
rect 443604 -6566 444204 -6564
rect 479604 -6566 480204 -6564
rect 515604 -6566 516204 -6564
rect 551604 -6566 552204 -6564
rect 590960 -6566 591560 -6564
rect -8576 -6904 -7976 -6902
rect 29604 -6904 30204 -6902
rect 65604 -6904 66204 -6902
rect 101604 -6904 102204 -6902
rect 137604 -6904 138204 -6902
rect 173604 -6904 174204 -6902
rect 209604 -6904 210204 -6902
rect 245604 -6904 246204 -6902
rect 281604 -6904 282204 -6902
rect 317604 -6904 318204 -6902
rect 353604 -6904 354204 -6902
rect 389604 -6904 390204 -6902
rect 425604 -6904 426204 -6902
rect 461604 -6904 462204 -6902
rect 497604 -6904 498204 -6902
rect 533604 -6904 534204 -6902
rect 569604 -6904 570204 -6902
rect 591900 -6904 592500 -6902
rect -8576 -6926 592500 -6904
rect -8576 -7162 -8394 -6926
rect -8158 -7162 29786 -6926
rect 30022 -7162 65786 -6926
rect 66022 -7162 101786 -6926
rect 102022 -7162 137786 -6926
rect 138022 -7162 173786 -6926
rect 174022 -7162 209786 -6926
rect 210022 -7162 245786 -6926
rect 246022 -7162 281786 -6926
rect 282022 -7162 317786 -6926
rect 318022 -7162 353786 -6926
rect 354022 -7162 389786 -6926
rect 390022 -7162 425786 -6926
rect 426022 -7162 461786 -6926
rect 462022 -7162 497786 -6926
rect 498022 -7162 533786 -6926
rect 534022 -7162 569786 -6926
rect 570022 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect -8576 -7246 592500 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 29786 -7246
rect 30022 -7482 65786 -7246
rect 66022 -7482 101786 -7246
rect 102022 -7482 137786 -7246
rect 138022 -7482 173786 -7246
rect 174022 -7482 209786 -7246
rect 210022 -7482 245786 -7246
rect 246022 -7482 281786 -7246
rect 282022 -7482 317786 -7246
rect 318022 -7482 353786 -7246
rect 354022 -7482 389786 -7246
rect 390022 -7482 425786 -7246
rect 426022 -7482 461786 -7246
rect 462022 -7482 497786 -7246
rect 498022 -7482 533786 -7246
rect 534022 -7482 569786 -7246
rect 570022 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect -8576 -7504 592500 -7482
rect -8576 -7506 -7976 -7504
rect 29604 -7506 30204 -7504
rect 65604 -7506 66204 -7504
rect 101604 -7506 102204 -7504
rect 137604 -7506 138204 -7504
rect 173604 -7506 174204 -7504
rect 209604 -7506 210204 -7504
rect 245604 -7506 246204 -7504
rect 281604 -7506 282204 -7504
rect 317604 -7506 318204 -7504
rect 353604 -7506 354204 -7504
rect 389604 -7506 390204 -7504
rect 425604 -7506 426204 -7504
rect 461604 -7506 462204 -7504
rect 497604 -7506 498204 -7504
rect 533604 -7506 534204 -7504
rect 569604 -7506 570204 -7504
rect 591900 -7506 592500 -7504
use sram_1rw1r_32_256_8_sky130  sram3
timestamp 1612306080
transform -1 0 497296 0 -1 201247
box 0 0 77296 91247
use sram_1rw1r_32_256_8_sky130  sram2
timestamp 1612306080
transform -1 0 377296 0 -1 201247
box 0 0 77296 91247
use sram_1rw1r_32_256_8_sky130  sram1
timestamp 1612306080
transform 1 0 420000 0 1 520000
box 0 0 77296 91247
use sram_1rw1r_32_256_8_sky130  sram0
timestamp 1612306080
transform 1 0 300000 0 1 520000
box 0 0 77296 91247
use hs32_core1  core1
timestamp 1612306080
transform 1 0 260000 0 1 240000
box 0 0 280000 240000
<< labels >>
rlabel metal3 s 583520 5796 584960 6036 6 analog_io[0]
port 0 nsew default bidirectional
rlabel metal3 s 583520 474996 584960 475236 6 analog_io[10]
port 1 nsew default bidirectional
rlabel metal3 s 583520 521916 584960 522156 6 analog_io[11]
port 2 nsew default bidirectional
rlabel metal3 s 583520 568836 584960 569076 6 analog_io[12]
port 3 nsew default bidirectional
rlabel metal3 s 583520 615756 584960 615996 6 analog_io[13]
port 4 nsew default bidirectional
rlabel metal3 s 583520 662676 584960 662916 6 analog_io[14]
port 5 nsew default bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[15]
port 6 nsew default bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[16]
port 7 nsew default bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[17]
port 8 nsew default bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[18]
port 9 nsew default bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[19]
port 10 nsew default bidirectional
rlabel metal3 s 583520 52716 584960 52956 6 analog_io[1]
port 11 nsew default bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[20]
port 12 nsew default bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[21]
port 13 nsew default bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[22]
port 14 nsew default bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[23]
port 15 nsew default bidirectional
rlabel metal3 s -960 696540 480 696780 4 analog_io[24]
port 16 nsew default bidirectional
rlabel metal3 s -960 639012 480 639252 4 analog_io[25]
port 17 nsew default bidirectional
rlabel metal3 s -960 581620 480 581860 4 analog_io[26]
port 18 nsew default bidirectional
rlabel metal3 s -960 524092 480 524332 4 analog_io[27]
port 19 nsew default bidirectional
rlabel metal3 s -960 466700 480 466940 4 analog_io[28]
port 20 nsew default bidirectional
rlabel metal3 s -960 409172 480 409412 4 analog_io[29]
port 21 nsew default bidirectional
rlabel metal3 s 583520 99636 584960 99876 6 analog_io[2]
port 22 nsew default bidirectional
rlabel metal3 s -960 351780 480 352020 4 analog_io[30]
port 23 nsew default bidirectional
rlabel metal3 s 583520 146556 584960 146796 6 analog_io[3]
port 24 nsew default bidirectional
rlabel metal3 s 583520 193476 584960 193716 6 analog_io[4]
port 25 nsew default bidirectional
rlabel metal3 s 583520 240396 584960 240636 6 analog_io[5]
port 26 nsew default bidirectional
rlabel metal3 s 583520 287316 584960 287556 6 analog_io[6]
port 27 nsew default bidirectional
rlabel metal3 s 583520 334236 584960 334476 6 analog_io[7]
port 28 nsew default bidirectional
rlabel metal3 s 583520 381156 584960 381396 6 analog_io[8]
port 29 nsew default bidirectional
rlabel metal3 s 583520 428076 584960 428316 6 analog_io[9]
port 30 nsew default bidirectional
rlabel metal3 s 583520 17492 584960 17732 6 io_in[0]
port 31 nsew default input
rlabel metal3 s 583520 486692 584960 486932 6 io_in[10]
port 32 nsew default input
rlabel metal3 s 583520 533748 584960 533988 6 io_in[11]
port 33 nsew default input
rlabel metal3 s 583520 580668 584960 580908 6 io_in[12]
port 34 nsew default input
rlabel metal3 s 583520 627588 584960 627828 6 io_in[13]
port 35 nsew default input
rlabel metal3 s 583520 674508 584960 674748 6 io_in[14]
port 36 nsew default input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 37 nsew default input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 38 nsew default input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 39 nsew default input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 40 nsew default input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 41 nsew default input
rlabel metal3 s 583520 64412 584960 64652 6 io_in[1]
port 42 nsew default input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 43 nsew default input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 44 nsew default input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 45 nsew default input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 46 nsew default input
rlabel metal3 s -960 682124 480 682364 4 io_in[24]
port 47 nsew default input
rlabel metal3 s -960 624732 480 624972 4 io_in[25]
port 48 nsew default input
rlabel metal3 s -960 567204 480 567444 4 io_in[26]
port 49 nsew default input
rlabel metal3 s -960 509812 480 510052 4 io_in[27]
port 50 nsew default input
rlabel metal3 s -960 452284 480 452524 4 io_in[28]
port 51 nsew default input
rlabel metal3 s -960 394892 480 395132 4 io_in[29]
port 52 nsew default input
rlabel metal3 s 583520 111332 584960 111572 6 io_in[2]
port 53 nsew default input
rlabel metal3 s -960 337364 480 337604 4 io_in[30]
port 54 nsew default input
rlabel metal3 s -960 294252 480 294492 4 io_in[31]
port 55 nsew default input
rlabel metal3 s -960 251140 480 251380 4 io_in[32]
port 56 nsew default input
rlabel metal3 s -960 208028 480 208268 4 io_in[33]
port 57 nsew default input
rlabel metal3 s -960 164916 480 165156 4 io_in[34]
port 58 nsew default input
rlabel metal3 s -960 121940 480 122180 4 io_in[35]
port 59 nsew default input
rlabel metal3 s -960 78828 480 79068 4 io_in[36]
port 60 nsew default input
rlabel metal3 s -960 35716 480 35956 4 io_in[37]
port 61 nsew default input
rlabel metal3 s 583520 158252 584960 158492 6 io_in[3]
port 62 nsew default input
rlabel metal3 s 583520 205172 584960 205412 6 io_in[4]
port 63 nsew default input
rlabel metal3 s 583520 252092 584960 252332 6 io_in[5]
port 64 nsew default input
rlabel metal3 s 583520 299012 584960 299252 6 io_in[6]
port 65 nsew default input
rlabel metal3 s 583520 345932 584960 346172 6 io_in[7]
port 66 nsew default input
rlabel metal3 s 583520 392852 584960 393092 6 io_in[8]
port 67 nsew default input
rlabel metal3 s 583520 439772 584960 440012 6 io_in[9]
port 68 nsew default input
rlabel metal3 s 583520 40884 584960 41124 6 io_oeb[0]
port 69 nsew default tristate
rlabel metal3 s 583520 510220 584960 510460 6 io_oeb[10]
port 70 nsew default tristate
rlabel metal3 s 583520 557140 584960 557380 6 io_oeb[11]
port 71 nsew default tristate
rlabel metal3 s 583520 604060 584960 604300 6 io_oeb[12]
port 72 nsew default tristate
rlabel metal3 s 583520 650980 584960 651220 6 io_oeb[13]
port 73 nsew default tristate
rlabel metal3 s 583520 697900 584960 698140 6 io_oeb[14]
port 74 nsew default tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 75 nsew default tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 76 nsew default tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 77 nsew default tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 78 nsew default tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 79 nsew default tristate
rlabel metal3 s 583520 87804 584960 88044 6 io_oeb[1]
port 80 nsew default tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 81 nsew default tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 82 nsew default tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 83 nsew default tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 84 nsew default tristate
rlabel metal3 s -960 653428 480 653668 4 io_oeb[24]
port 85 nsew default tristate
rlabel metal3 s -960 595900 480 596140 4 io_oeb[25]
port 86 nsew default tristate
rlabel metal3 s -960 538508 480 538748 4 io_oeb[26]
port 87 nsew default tristate
rlabel metal3 s -960 480980 480 481220 4 io_oeb[27]
port 88 nsew default tristate
rlabel metal3 s -960 423588 480 423828 4 io_oeb[28]
port 89 nsew default tristate
rlabel metal3 s -960 366060 480 366300 4 io_oeb[29]
port 90 nsew default tristate
rlabel metal3 s 583520 134724 584960 134964 6 io_oeb[2]
port 91 nsew default tristate
rlabel metal3 s -960 308668 480 308908 4 io_oeb[30]
port 92 nsew default tristate
rlabel metal3 s -960 265556 480 265796 4 io_oeb[31]
port 93 nsew default tristate
rlabel metal3 s -960 222444 480 222684 4 io_oeb[32]
port 94 nsew default tristate
rlabel metal3 s -960 179332 480 179572 4 io_oeb[33]
port 95 nsew default tristate
rlabel metal3 s -960 136220 480 136460 4 io_oeb[34]
port 96 nsew default tristate
rlabel metal3 s -960 93108 480 93348 4 io_oeb[35]
port 97 nsew default tristate
rlabel metal3 s -960 49996 480 50236 4 io_oeb[36]
port 98 nsew default tristate
rlabel metal3 s -960 7020 480 7260 4 io_oeb[37]
port 99 nsew default tristate
rlabel metal3 s 583520 181780 584960 182020 6 io_oeb[3]
port 100 nsew default tristate
rlabel metal3 s 583520 228700 584960 228940 6 io_oeb[4]
port 101 nsew default tristate
rlabel metal3 s 583520 275620 584960 275860 6 io_oeb[5]
port 102 nsew default tristate
rlabel metal3 s 583520 322540 584960 322780 6 io_oeb[6]
port 103 nsew default tristate
rlabel metal3 s 583520 369460 584960 369700 6 io_oeb[7]
port 104 nsew default tristate
rlabel metal3 s 583520 416380 584960 416620 6 io_oeb[8]
port 105 nsew default tristate
rlabel metal3 s 583520 463300 584960 463540 6 io_oeb[9]
port 106 nsew default tristate
rlabel metal3 s 583520 29188 584960 29428 6 io_out[0]
port 107 nsew default tristate
rlabel metal3 s 583520 498524 584960 498764 6 io_out[10]
port 108 nsew default tristate
rlabel metal3 s 583520 545444 584960 545684 6 io_out[11]
port 109 nsew default tristate
rlabel metal3 s 583520 592364 584960 592604 6 io_out[12]
port 110 nsew default tristate
rlabel metal3 s 583520 639284 584960 639524 6 io_out[13]
port 111 nsew default tristate
rlabel metal3 s 583520 686204 584960 686444 6 io_out[14]
port 112 nsew default tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 113 nsew default tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 114 nsew default tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 115 nsew default tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 116 nsew default tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 117 nsew default tristate
rlabel metal3 s 583520 76108 584960 76348 6 io_out[1]
port 118 nsew default tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 119 nsew default tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 120 nsew default tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 121 nsew default tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 122 nsew default tristate
rlabel metal3 s -960 667844 480 668084 4 io_out[24]
port 123 nsew default tristate
rlabel metal3 s -960 610316 480 610556 4 io_out[25]
port 124 nsew default tristate
rlabel metal3 s -960 552924 480 553164 4 io_out[26]
port 125 nsew default tristate
rlabel metal3 s -960 495396 480 495636 4 io_out[27]
port 126 nsew default tristate
rlabel metal3 s -960 437868 480 438108 4 io_out[28]
port 127 nsew default tristate
rlabel metal3 s -960 380476 480 380716 4 io_out[29]
port 128 nsew default tristate
rlabel metal3 s 583520 123028 584960 123268 6 io_out[2]
port 129 nsew default tristate
rlabel metal3 s -960 322948 480 323188 4 io_out[30]
port 130 nsew default tristate
rlabel metal3 s -960 279972 480 280212 4 io_out[31]
port 131 nsew default tristate
rlabel metal3 s -960 236860 480 237100 4 io_out[32]
port 132 nsew default tristate
rlabel metal3 s -960 193748 480 193988 4 io_out[33]
port 133 nsew default tristate
rlabel metal3 s -960 150636 480 150876 4 io_out[34]
port 134 nsew default tristate
rlabel metal3 s -960 107524 480 107764 4 io_out[35]
port 135 nsew default tristate
rlabel metal3 s -960 64412 480 64652 4 io_out[36]
port 136 nsew default tristate
rlabel metal3 s -960 21300 480 21540 4 io_out[37]
port 137 nsew default tristate
rlabel metal3 s 583520 169948 584960 170188 6 io_out[3]
port 138 nsew default tristate
rlabel metal3 s 583520 216868 584960 217108 6 io_out[4]
port 139 nsew default tristate
rlabel metal3 s 583520 263788 584960 264028 6 io_out[5]
port 140 nsew default tristate
rlabel metal3 s 583520 310708 584960 310948 6 io_out[6]
port 141 nsew default tristate
rlabel metal3 s 583520 357764 584960 358004 6 io_out[7]
port 142 nsew default tristate
rlabel metal3 s 583520 404684 584960 404924 6 io_out[8]
port 143 nsew default tristate
rlabel metal3 s 583520 451604 584960 451844 6 io_out[9]
port 144 nsew default tristate
rlabel metal2 s 126582 -960 126694 480 8 la_data_in[0]
port 145 nsew default input
rlabel metal2 s 483450 -960 483562 480 8 la_data_in[100]
port 146 nsew default input
rlabel metal2 s 486946 -960 487058 480 8 la_data_in[101]
port 147 nsew default input
rlabel metal2 s 490534 -960 490646 480 8 la_data_in[102]
port 148 nsew default input
rlabel metal2 s 494122 -960 494234 480 8 la_data_in[103]
port 149 nsew default input
rlabel metal2 s 497710 -960 497822 480 8 la_data_in[104]
port 150 nsew default input
rlabel metal2 s 501206 -960 501318 480 8 la_data_in[105]
port 151 nsew default input
rlabel metal2 s 504794 -960 504906 480 8 la_data_in[106]
port 152 nsew default input
rlabel metal2 s 508382 -960 508494 480 8 la_data_in[107]
port 153 nsew default input
rlabel metal2 s 511970 -960 512082 480 8 la_data_in[108]
port 154 nsew default input
rlabel metal2 s 515558 -960 515670 480 8 la_data_in[109]
port 155 nsew default input
rlabel metal2 s 162278 -960 162390 480 8 la_data_in[10]
port 156 nsew default input
rlabel metal2 s 519054 -960 519166 480 8 la_data_in[110]
port 157 nsew default input
rlabel metal2 s 522642 -960 522754 480 8 la_data_in[111]
port 158 nsew default input
rlabel metal2 s 526230 -960 526342 480 8 la_data_in[112]
port 159 nsew default input
rlabel metal2 s 529818 -960 529930 480 8 la_data_in[113]
port 160 nsew default input
rlabel metal2 s 533406 -960 533518 480 8 la_data_in[114]
port 161 nsew default input
rlabel metal2 s 536902 -960 537014 480 8 la_data_in[115]
port 162 nsew default input
rlabel metal2 s 540490 -960 540602 480 8 la_data_in[116]
port 163 nsew default input
rlabel metal2 s 544078 -960 544190 480 8 la_data_in[117]
port 164 nsew default input
rlabel metal2 s 547666 -960 547778 480 8 la_data_in[118]
port 165 nsew default input
rlabel metal2 s 551162 -960 551274 480 8 la_data_in[119]
port 166 nsew default input
rlabel metal2 s 165866 -960 165978 480 8 la_data_in[11]
port 167 nsew default input
rlabel metal2 s 554750 -960 554862 480 8 la_data_in[120]
port 168 nsew default input
rlabel metal2 s 558338 -960 558450 480 8 la_data_in[121]
port 169 nsew default input
rlabel metal2 s 561926 -960 562038 480 8 la_data_in[122]
port 170 nsew default input
rlabel metal2 s 565514 -960 565626 480 8 la_data_in[123]
port 171 nsew default input
rlabel metal2 s 569010 -960 569122 480 8 la_data_in[124]
port 172 nsew default input
rlabel metal2 s 572598 -960 572710 480 8 la_data_in[125]
port 173 nsew default input
rlabel metal2 s 576186 -960 576298 480 8 la_data_in[126]
port 174 nsew default input
rlabel metal2 s 579774 -960 579886 480 8 la_data_in[127]
port 175 nsew default input
rlabel metal2 s 169362 -960 169474 480 8 la_data_in[12]
port 176 nsew default input
rlabel metal2 s 172950 -960 173062 480 8 la_data_in[13]
port 177 nsew default input
rlabel metal2 s 176538 -960 176650 480 8 la_data_in[14]
port 178 nsew default input
rlabel metal2 s 180126 -960 180238 480 8 la_data_in[15]
port 179 nsew default input
rlabel metal2 s 183714 -960 183826 480 8 la_data_in[16]
port 180 nsew default input
rlabel metal2 s 187210 -960 187322 480 8 la_data_in[17]
port 181 nsew default input
rlabel metal2 s 190798 -960 190910 480 8 la_data_in[18]
port 182 nsew default input
rlabel metal2 s 194386 -960 194498 480 8 la_data_in[19]
port 183 nsew default input
rlabel metal2 s 130170 -960 130282 480 8 la_data_in[1]
port 184 nsew default input
rlabel metal2 s 197974 -960 198086 480 8 la_data_in[20]
port 185 nsew default input
rlabel metal2 s 201470 -960 201582 480 8 la_data_in[21]
port 186 nsew default input
rlabel metal2 s 205058 -960 205170 480 8 la_data_in[22]
port 187 nsew default input
rlabel metal2 s 208646 -960 208758 480 8 la_data_in[23]
port 188 nsew default input
rlabel metal2 s 212234 -960 212346 480 8 la_data_in[24]
port 189 nsew default input
rlabel metal2 s 215822 -960 215934 480 8 la_data_in[25]
port 190 nsew default input
rlabel metal2 s 219318 -960 219430 480 8 la_data_in[26]
port 191 nsew default input
rlabel metal2 s 222906 -960 223018 480 8 la_data_in[27]
port 192 nsew default input
rlabel metal2 s 226494 -960 226606 480 8 la_data_in[28]
port 193 nsew default input
rlabel metal2 s 230082 -960 230194 480 8 la_data_in[29]
port 194 nsew default input
rlabel metal2 s 133758 -960 133870 480 8 la_data_in[2]
port 195 nsew default input
rlabel metal2 s 233670 -960 233782 480 8 la_data_in[30]
port 196 nsew default input
rlabel metal2 s 237166 -960 237278 480 8 la_data_in[31]
port 197 nsew default input
rlabel metal2 s 240754 -960 240866 480 8 la_data_in[32]
port 198 nsew default input
rlabel metal2 s 244342 -960 244454 480 8 la_data_in[33]
port 199 nsew default input
rlabel metal2 s 247930 -960 248042 480 8 la_data_in[34]
port 200 nsew default input
rlabel metal2 s 251426 -960 251538 480 8 la_data_in[35]
port 201 nsew default input
rlabel metal2 s 255014 -960 255126 480 8 la_data_in[36]
port 202 nsew default input
rlabel metal2 s 258602 -960 258714 480 8 la_data_in[37]
port 203 nsew default input
rlabel metal2 s 262190 -960 262302 480 8 la_data_in[38]
port 204 nsew default input
rlabel metal2 s 265778 -960 265890 480 8 la_data_in[39]
port 205 nsew default input
rlabel metal2 s 137254 -960 137366 480 8 la_data_in[3]
port 206 nsew default input
rlabel metal2 s 269274 -960 269386 480 8 la_data_in[40]
port 207 nsew default input
rlabel metal2 s 272862 -960 272974 480 8 la_data_in[41]
port 208 nsew default input
rlabel metal2 s 276450 -960 276562 480 8 la_data_in[42]
port 209 nsew default input
rlabel metal2 s 280038 -960 280150 480 8 la_data_in[43]
port 210 nsew default input
rlabel metal2 s 283626 -960 283738 480 8 la_data_in[44]
port 211 nsew default input
rlabel metal2 s 287122 -960 287234 480 8 la_data_in[45]
port 212 nsew default input
rlabel metal2 s 290710 -960 290822 480 8 la_data_in[46]
port 213 nsew default input
rlabel metal2 s 294298 -960 294410 480 8 la_data_in[47]
port 214 nsew default input
rlabel metal2 s 297886 -960 297998 480 8 la_data_in[48]
port 215 nsew default input
rlabel metal2 s 301382 -960 301494 480 8 la_data_in[49]
port 216 nsew default input
rlabel metal2 s 140842 -960 140954 480 8 la_data_in[4]
port 217 nsew default input
rlabel metal2 s 304970 -960 305082 480 8 la_data_in[50]
port 218 nsew default input
rlabel metal2 s 308558 -960 308670 480 8 la_data_in[51]
port 219 nsew default input
rlabel metal2 s 312146 -960 312258 480 8 la_data_in[52]
port 220 nsew default input
rlabel metal2 s 315734 -960 315846 480 8 la_data_in[53]
port 221 nsew default input
rlabel metal2 s 319230 -960 319342 480 8 la_data_in[54]
port 222 nsew default input
rlabel metal2 s 322818 -960 322930 480 8 la_data_in[55]
port 223 nsew default input
rlabel metal2 s 326406 -960 326518 480 8 la_data_in[56]
port 224 nsew default input
rlabel metal2 s 329994 -960 330106 480 8 la_data_in[57]
port 225 nsew default input
rlabel metal2 s 333582 -960 333694 480 8 la_data_in[58]
port 226 nsew default input
rlabel metal2 s 337078 -960 337190 480 8 la_data_in[59]
port 227 nsew default input
rlabel metal2 s 144430 -960 144542 480 8 la_data_in[5]
port 228 nsew default input
rlabel metal2 s 340666 -960 340778 480 8 la_data_in[60]
port 229 nsew default input
rlabel metal2 s 344254 -960 344366 480 8 la_data_in[61]
port 230 nsew default input
rlabel metal2 s 347842 -960 347954 480 8 la_data_in[62]
port 231 nsew default input
rlabel metal2 s 351338 -960 351450 480 8 la_data_in[63]
port 232 nsew default input
rlabel metal2 s 354926 -960 355038 480 8 la_data_in[64]
port 233 nsew default input
rlabel metal2 s 358514 -960 358626 480 8 la_data_in[65]
port 234 nsew default input
rlabel metal2 s 362102 -960 362214 480 8 la_data_in[66]
port 235 nsew default input
rlabel metal2 s 365690 -960 365802 480 8 la_data_in[67]
port 236 nsew default input
rlabel metal2 s 369186 -960 369298 480 8 la_data_in[68]
port 237 nsew default input
rlabel metal2 s 372774 -960 372886 480 8 la_data_in[69]
port 238 nsew default input
rlabel metal2 s 148018 -960 148130 480 8 la_data_in[6]
port 239 nsew default input
rlabel metal2 s 376362 -960 376474 480 8 la_data_in[70]
port 240 nsew default input
rlabel metal2 s 379950 -960 380062 480 8 la_data_in[71]
port 241 nsew default input
rlabel metal2 s 383538 -960 383650 480 8 la_data_in[72]
port 242 nsew default input
rlabel metal2 s 387034 -960 387146 480 8 la_data_in[73]
port 243 nsew default input
rlabel metal2 s 390622 -960 390734 480 8 la_data_in[74]
port 244 nsew default input
rlabel metal2 s 394210 -960 394322 480 8 la_data_in[75]
port 245 nsew default input
rlabel metal2 s 397798 -960 397910 480 8 la_data_in[76]
port 246 nsew default input
rlabel metal2 s 401294 -960 401406 480 8 la_data_in[77]
port 247 nsew default input
rlabel metal2 s 404882 -960 404994 480 8 la_data_in[78]
port 248 nsew default input
rlabel metal2 s 408470 -960 408582 480 8 la_data_in[79]
port 249 nsew default input
rlabel metal2 s 151514 -960 151626 480 8 la_data_in[7]
port 250 nsew default input
rlabel metal2 s 412058 -960 412170 480 8 la_data_in[80]
port 251 nsew default input
rlabel metal2 s 415646 -960 415758 480 8 la_data_in[81]
port 252 nsew default input
rlabel metal2 s 419142 -960 419254 480 8 la_data_in[82]
port 253 nsew default input
rlabel metal2 s 422730 -960 422842 480 8 la_data_in[83]
port 254 nsew default input
rlabel metal2 s 426318 -960 426430 480 8 la_data_in[84]
port 255 nsew default input
rlabel metal2 s 429906 -960 430018 480 8 la_data_in[85]
port 256 nsew default input
rlabel metal2 s 433494 -960 433606 480 8 la_data_in[86]
port 257 nsew default input
rlabel metal2 s 436990 -960 437102 480 8 la_data_in[87]
port 258 nsew default input
rlabel metal2 s 440578 -960 440690 480 8 la_data_in[88]
port 259 nsew default input
rlabel metal2 s 444166 -960 444278 480 8 la_data_in[89]
port 260 nsew default input
rlabel metal2 s 155102 -960 155214 480 8 la_data_in[8]
port 261 nsew default input
rlabel metal2 s 447754 -960 447866 480 8 la_data_in[90]
port 262 nsew default input
rlabel metal2 s 451250 -960 451362 480 8 la_data_in[91]
port 263 nsew default input
rlabel metal2 s 454838 -960 454950 480 8 la_data_in[92]
port 264 nsew default input
rlabel metal2 s 458426 -960 458538 480 8 la_data_in[93]
port 265 nsew default input
rlabel metal2 s 462014 -960 462126 480 8 la_data_in[94]
port 266 nsew default input
rlabel metal2 s 465602 -960 465714 480 8 la_data_in[95]
port 267 nsew default input
rlabel metal2 s 469098 -960 469210 480 8 la_data_in[96]
port 268 nsew default input
rlabel metal2 s 472686 -960 472798 480 8 la_data_in[97]
port 269 nsew default input
rlabel metal2 s 476274 -960 476386 480 8 la_data_in[98]
port 270 nsew default input
rlabel metal2 s 479862 -960 479974 480 8 la_data_in[99]
port 271 nsew default input
rlabel metal2 s 158690 -960 158802 480 8 la_data_in[9]
port 272 nsew default input
rlabel metal2 s 127778 -960 127890 480 8 la_data_out[0]
port 273 nsew default tristate
rlabel metal2 s 131366 -960 131478 480 8 la_data_out[1]
port 274 nsew default tristate
rlabel metal2 s 134862 -960 134974 480 8 la_data_out[2]
port 275 nsew default tristate
rlabel metal2 s 128974 -960 129086 480 8 la_oen[0]
port 276 nsew default input
rlabel metal2 s 485750 -960 485862 480 8 la_oen[100]
port 277 nsew default input
rlabel metal2 s 489338 -960 489450 480 8 la_oen[101]
port 278 nsew default input
rlabel metal2 s 492926 -960 493038 480 8 la_oen[102]
port 279 nsew default input
rlabel metal2 s 496514 -960 496626 480 8 la_oen[103]
port 280 nsew default input
rlabel metal2 s 500102 -960 500214 480 8 la_oen[104]
port 281 nsew default input
rlabel metal2 s 503598 -960 503710 480 8 la_oen[105]
port 282 nsew default input
rlabel metal2 s 507186 -960 507298 480 8 la_oen[106]
port 283 nsew default input
rlabel metal2 s 510774 -960 510886 480 8 la_oen[107]
port 284 nsew default input
rlabel metal2 s 514362 -960 514474 480 8 la_oen[108]
port 285 nsew default input
rlabel metal2 s 517858 -960 517970 480 8 la_oen[109]
port 286 nsew default input
rlabel metal2 s 164670 -960 164782 480 8 la_oen[10]
port 287 nsew default input
rlabel metal2 s 521446 -960 521558 480 8 la_oen[110]
port 288 nsew default input
rlabel metal2 s 525034 -960 525146 480 8 la_oen[111]
port 289 nsew default input
rlabel metal2 s 528622 -960 528734 480 8 la_oen[112]
port 290 nsew default input
rlabel metal2 s 532210 -960 532322 480 8 la_oen[113]
port 291 nsew default input
rlabel metal2 s 535706 -960 535818 480 8 la_oen[114]
port 292 nsew default input
rlabel metal2 s 539294 -960 539406 480 8 la_oen[115]
port 293 nsew default input
rlabel metal2 s 542882 -960 542994 480 8 la_oen[116]
port 294 nsew default input
rlabel metal2 s 546470 -960 546582 480 8 la_oen[117]
port 295 nsew default input
rlabel metal2 s 550058 -960 550170 480 8 la_oen[118]
port 296 nsew default input
rlabel metal2 s 553554 -960 553666 480 8 la_oen[119]
port 297 nsew default input
rlabel metal2 s 168166 -960 168278 480 8 la_oen[11]
port 298 nsew default input
rlabel metal2 s 557142 -960 557254 480 8 la_oen[120]
port 299 nsew default input
rlabel metal2 s 560730 -960 560842 480 8 la_oen[121]
port 300 nsew default input
rlabel metal2 s 564318 -960 564430 480 8 la_oen[122]
port 301 nsew default input
rlabel metal2 s 567814 -960 567926 480 8 la_oen[123]
port 302 nsew default input
rlabel metal2 s 571402 -960 571514 480 8 la_oen[124]
port 303 nsew default input
rlabel metal2 s 574990 -960 575102 480 8 la_oen[125]
port 304 nsew default input
rlabel metal2 s 578578 -960 578690 480 8 la_oen[126]
port 305 nsew default input
rlabel metal2 s 582166 -960 582278 480 8 la_oen[127]
port 306 nsew default input
rlabel metal2 s 171754 -960 171866 480 8 la_oen[12]
port 307 nsew default input
rlabel metal2 s 175342 -960 175454 480 8 la_oen[13]
port 308 nsew default input
rlabel metal2 s 178930 -960 179042 480 8 la_oen[14]
port 309 nsew default input
rlabel metal2 s 182518 -960 182630 480 8 la_oen[15]
port 310 nsew default input
rlabel metal2 s 186014 -960 186126 480 8 la_oen[16]
port 311 nsew default input
rlabel metal2 s 189602 -960 189714 480 8 la_oen[17]
port 312 nsew default input
rlabel metal2 s 193190 -960 193302 480 8 la_oen[18]
port 313 nsew default input
rlabel metal2 s 196778 -960 196890 480 8 la_oen[19]
port 314 nsew default input
rlabel metal2 s 132562 -960 132674 480 8 la_oen[1]
port 315 nsew default input
rlabel metal2 s 200366 -960 200478 480 8 la_oen[20]
port 316 nsew default input
rlabel metal2 s 203862 -960 203974 480 8 la_oen[21]
port 317 nsew default input
rlabel metal2 s 207450 -960 207562 480 8 la_oen[22]
port 318 nsew default input
rlabel metal2 s 211038 -960 211150 480 8 la_oen[23]
port 319 nsew default input
rlabel metal2 s 214626 -960 214738 480 8 la_oen[24]
port 320 nsew default input
rlabel metal2 s 218122 -960 218234 480 8 la_oen[25]
port 321 nsew default input
rlabel metal2 s 221710 -960 221822 480 8 la_oen[26]
port 322 nsew default input
rlabel metal2 s 225298 -960 225410 480 8 la_oen[27]
port 323 nsew default input
rlabel metal2 s 228886 -960 228998 480 8 la_oen[28]
port 324 nsew default input
rlabel metal2 s 232474 -960 232586 480 8 la_oen[29]
port 325 nsew default input
rlabel metal2 s 136058 -960 136170 480 8 la_oen[2]
port 326 nsew default input
rlabel metal2 s 235970 -960 236082 480 8 la_oen[30]
port 327 nsew default input
rlabel metal2 s 239558 -960 239670 480 8 la_oen[31]
port 328 nsew default input
rlabel metal2 s 243146 -960 243258 480 8 la_oen[32]
port 329 nsew default input
rlabel metal2 s 246734 -960 246846 480 8 la_oen[33]
port 330 nsew default input
rlabel metal2 s 250322 -960 250434 480 8 la_oen[34]
port 331 nsew default input
rlabel metal2 s 253818 -960 253930 480 8 la_oen[35]
port 332 nsew default input
rlabel metal2 s 257406 -960 257518 480 8 la_oen[36]
port 333 nsew default input
rlabel metal2 s 260994 -960 261106 480 8 la_oen[37]
port 334 nsew default input
rlabel metal2 s 264582 -960 264694 480 8 la_oen[38]
port 335 nsew default input
rlabel metal2 s 268078 -960 268190 480 8 la_oen[39]
port 336 nsew default input
rlabel metal2 s 139646 -960 139758 480 8 la_oen[3]
port 337 nsew default input
rlabel metal2 s 271666 -960 271778 480 8 la_oen[40]
port 338 nsew default input
rlabel metal2 s 275254 -960 275366 480 8 la_oen[41]
port 339 nsew default input
rlabel metal2 s 278842 -960 278954 480 8 la_oen[42]
port 340 nsew default input
rlabel metal2 s 282430 -960 282542 480 8 la_oen[43]
port 341 nsew default input
rlabel metal2 s 285926 -960 286038 480 8 la_oen[44]
port 342 nsew default input
rlabel metal2 s 289514 -960 289626 480 8 la_oen[45]
port 343 nsew default input
rlabel metal2 s 293102 -960 293214 480 8 la_oen[46]
port 344 nsew default input
rlabel metal2 s 296690 -960 296802 480 8 la_oen[47]
port 345 nsew default input
rlabel metal2 s 300278 -960 300390 480 8 la_oen[48]
port 346 nsew default input
rlabel metal2 s 303774 -960 303886 480 8 la_oen[49]
port 347 nsew default input
rlabel metal2 s 143234 -960 143346 480 8 la_oen[4]
port 348 nsew default input
rlabel metal2 s 307362 -960 307474 480 8 la_oen[50]
port 349 nsew default input
rlabel metal2 s 310950 -960 311062 480 8 la_oen[51]
port 350 nsew default input
rlabel metal2 s 314538 -960 314650 480 8 la_oen[52]
port 351 nsew default input
rlabel metal2 s 318034 -960 318146 480 8 la_oen[53]
port 352 nsew default input
rlabel metal2 s 321622 -960 321734 480 8 la_oen[54]
port 353 nsew default input
rlabel metal2 s 325210 -960 325322 480 8 la_oen[55]
port 354 nsew default input
rlabel metal2 s 328798 -960 328910 480 8 la_oen[56]
port 355 nsew default input
rlabel metal2 s 332386 -960 332498 480 8 la_oen[57]
port 356 nsew default input
rlabel metal2 s 335882 -960 335994 480 8 la_oen[58]
port 357 nsew default input
rlabel metal2 s 339470 -960 339582 480 8 la_oen[59]
port 358 nsew default input
rlabel metal2 s 146822 -960 146934 480 8 la_oen[5]
port 359 nsew default input
rlabel metal2 s 343058 -960 343170 480 8 la_oen[60]
port 360 nsew default input
rlabel metal2 s 346646 -960 346758 480 8 la_oen[61]
port 361 nsew default input
rlabel metal2 s 350234 -960 350346 480 8 la_oen[62]
port 362 nsew default input
rlabel metal2 s 353730 -960 353842 480 8 la_oen[63]
port 363 nsew default input
rlabel metal2 s 357318 -960 357430 480 8 la_oen[64]
port 364 nsew default input
rlabel metal2 s 360906 -960 361018 480 8 la_oen[65]
port 365 nsew default input
rlabel metal2 s 364494 -960 364606 480 8 la_oen[66]
port 366 nsew default input
rlabel metal2 s 367990 -960 368102 480 8 la_oen[67]
port 367 nsew default input
rlabel metal2 s 371578 -960 371690 480 8 la_oen[68]
port 368 nsew default input
rlabel metal2 s 375166 -960 375278 480 8 la_oen[69]
port 369 nsew default input
rlabel metal2 s 150410 -960 150522 480 8 la_oen[6]
port 370 nsew default input
rlabel metal2 s 378754 -960 378866 480 8 la_oen[70]
port 371 nsew default input
rlabel metal2 s 382342 -960 382454 480 8 la_oen[71]
port 372 nsew default input
rlabel metal2 s 385838 -960 385950 480 8 la_oen[72]
port 373 nsew default input
rlabel metal2 s 389426 -960 389538 480 8 la_oen[73]
port 374 nsew default input
rlabel metal2 s 393014 -960 393126 480 8 la_oen[74]
port 375 nsew default input
rlabel metal2 s 396602 -960 396714 480 8 la_oen[75]
port 376 nsew default input
rlabel metal2 s 400190 -960 400302 480 8 la_oen[76]
port 377 nsew default input
rlabel metal2 s 403686 -960 403798 480 8 la_oen[77]
port 378 nsew default input
rlabel metal2 s 407274 -960 407386 480 8 la_oen[78]
port 379 nsew default input
rlabel metal2 s 410862 -960 410974 480 8 la_oen[79]
port 380 nsew default input
rlabel metal2 s 153906 -960 154018 480 8 la_oen[7]
port 381 nsew default input
rlabel metal2 s 414450 -960 414562 480 8 la_oen[80]
port 382 nsew default input
rlabel metal2 s 417946 -960 418058 480 8 la_oen[81]
port 383 nsew default input
rlabel metal2 s 421534 -960 421646 480 8 la_oen[82]
port 384 nsew default input
rlabel metal2 s 425122 -960 425234 480 8 la_oen[83]
port 385 nsew default input
rlabel metal2 s 428710 -960 428822 480 8 la_oen[84]
port 386 nsew default input
rlabel metal2 s 432298 -960 432410 480 8 la_oen[85]
port 387 nsew default input
rlabel metal2 s 435794 -960 435906 480 8 la_oen[86]
port 388 nsew default input
rlabel metal2 s 439382 -960 439494 480 8 la_oen[87]
port 389 nsew default input
rlabel metal2 s 442970 -960 443082 480 8 la_oen[88]
port 390 nsew default input
rlabel metal2 s 446558 -960 446670 480 8 la_oen[89]
port 391 nsew default input
rlabel metal2 s 157494 -960 157606 480 8 la_oen[8]
port 392 nsew default input
rlabel metal2 s 450146 -960 450258 480 8 la_oen[90]
port 393 nsew default input
rlabel metal2 s 453642 -960 453754 480 8 la_oen[91]
port 394 nsew default input
rlabel metal2 s 457230 -960 457342 480 8 la_oen[92]
port 395 nsew default input
rlabel metal2 s 460818 -960 460930 480 8 la_oen[93]
port 396 nsew default input
rlabel metal2 s 464406 -960 464518 480 8 la_oen[94]
port 397 nsew default input
rlabel metal2 s 467902 -960 468014 480 8 la_oen[95]
port 398 nsew default input
rlabel metal2 s 471490 -960 471602 480 8 la_oen[96]
port 399 nsew default input
rlabel metal2 s 475078 -960 475190 480 8 la_oen[97]
port 400 nsew default input
rlabel metal2 s 478666 -960 478778 480 8 la_oen[98]
port 401 nsew default input
rlabel metal2 s 482254 -960 482366 480 8 la_oen[99]
port 402 nsew default input
rlabel metal2 s 161082 -960 161194 480 8 la_oen[9]
port 403 nsew default input
rlabel metal2 s 583362 -960 583474 480 8 user_clock2
port 404 nsew default input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 405 nsew default input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 406 nsew default input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 407 nsew default tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 408 nsew default input
rlabel metal2 s 48106 -960 48218 480 8 wbs_adr_i[10]
port 409 nsew default input
rlabel metal2 s 51602 -960 51714 480 8 wbs_adr_i[11]
port 410 nsew default input
rlabel metal2 s 55190 -960 55302 480 8 wbs_adr_i[12]
port 411 nsew default input
rlabel metal2 s 58778 -960 58890 480 8 wbs_adr_i[13]
port 412 nsew default input
rlabel metal2 s 62366 -960 62478 480 8 wbs_adr_i[14]
port 413 nsew default input
rlabel metal2 s 65954 -960 66066 480 8 wbs_adr_i[15]
port 414 nsew default input
rlabel metal2 s 69450 -960 69562 480 8 wbs_adr_i[16]
port 415 nsew default input
rlabel metal2 s 73038 -960 73150 480 8 wbs_adr_i[17]
port 416 nsew default input
rlabel metal2 s 76626 -960 76738 480 8 wbs_adr_i[18]
port 417 nsew default input
rlabel metal2 s 80214 -960 80326 480 8 wbs_adr_i[19]
port 418 nsew default input
rlabel metal2 s 12410 -960 12522 480 8 wbs_adr_i[1]
port 419 nsew default input
rlabel metal2 s 83802 -960 83914 480 8 wbs_adr_i[20]
port 420 nsew default input
rlabel metal2 s 87298 -960 87410 480 8 wbs_adr_i[21]
port 421 nsew default input
rlabel metal2 s 90886 -960 90998 480 8 wbs_adr_i[22]
port 422 nsew default input
rlabel metal2 s 94474 -960 94586 480 8 wbs_adr_i[23]
port 423 nsew default input
rlabel metal2 s 98062 -960 98174 480 8 wbs_adr_i[24]
port 424 nsew default input
rlabel metal2 s 101558 -960 101670 480 8 wbs_adr_i[25]
port 425 nsew default input
rlabel metal2 s 105146 -960 105258 480 8 wbs_adr_i[26]
port 426 nsew default input
rlabel metal2 s 108734 -960 108846 480 8 wbs_adr_i[27]
port 427 nsew default input
rlabel metal2 s 112322 -960 112434 480 8 wbs_adr_i[28]
port 428 nsew default input
rlabel metal2 s 115910 -960 116022 480 8 wbs_adr_i[29]
port 429 nsew default input
rlabel metal2 s 17194 -960 17306 480 8 wbs_adr_i[2]
port 430 nsew default input
rlabel metal2 s 119406 -960 119518 480 8 wbs_adr_i[30]
port 431 nsew default input
rlabel metal2 s 122994 -960 123106 480 8 wbs_adr_i[31]
port 432 nsew default input
rlabel metal2 s 21886 -960 21998 480 8 wbs_adr_i[3]
port 433 nsew default input
rlabel metal2 s 26670 -960 26782 480 8 wbs_adr_i[4]
port 434 nsew default input
rlabel metal2 s 30258 -960 30370 480 8 wbs_adr_i[5]
port 435 nsew default input
rlabel metal2 s 33846 -960 33958 480 8 wbs_adr_i[6]
port 436 nsew default input
rlabel metal2 s 37342 -960 37454 480 8 wbs_adr_i[7]
port 437 nsew default input
rlabel metal2 s 40930 -960 41042 480 8 wbs_adr_i[8]
port 438 nsew default input
rlabel metal2 s 44518 -960 44630 480 8 wbs_adr_i[9]
port 439 nsew default input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 440 nsew default input
rlabel metal2 s 8822 -960 8934 480 8 wbs_dat_i[0]
port 441 nsew default input
rlabel metal2 s 49302 -960 49414 480 8 wbs_dat_i[10]
port 442 nsew default input
rlabel metal2 s 52798 -960 52910 480 8 wbs_dat_i[11]
port 443 nsew default input
rlabel metal2 s 56386 -960 56498 480 8 wbs_dat_i[12]
port 444 nsew default input
rlabel metal2 s 59974 -960 60086 480 8 wbs_dat_i[13]
port 445 nsew default input
rlabel metal2 s 63562 -960 63674 480 8 wbs_dat_i[14]
port 446 nsew default input
rlabel metal2 s 67150 -960 67262 480 8 wbs_dat_i[15]
port 447 nsew default input
rlabel metal2 s 70646 -960 70758 480 8 wbs_dat_i[16]
port 448 nsew default input
rlabel metal2 s 74234 -960 74346 480 8 wbs_dat_i[17]
port 449 nsew default input
rlabel metal2 s 77822 -960 77934 480 8 wbs_dat_i[18]
port 450 nsew default input
rlabel metal2 s 81410 -960 81522 480 8 wbs_dat_i[19]
port 451 nsew default input
rlabel metal2 s 13606 -960 13718 480 8 wbs_dat_i[1]
port 452 nsew default input
rlabel metal2 s 84906 -960 85018 480 8 wbs_dat_i[20]
port 453 nsew default input
rlabel metal2 s 88494 -960 88606 480 8 wbs_dat_i[21]
port 454 nsew default input
rlabel metal2 s 92082 -960 92194 480 8 wbs_dat_i[22]
port 455 nsew default input
rlabel metal2 s 95670 -960 95782 480 8 wbs_dat_i[23]
port 456 nsew default input
rlabel metal2 s 99258 -960 99370 480 8 wbs_dat_i[24]
port 457 nsew default input
rlabel metal2 s 102754 -960 102866 480 8 wbs_dat_i[25]
port 458 nsew default input
rlabel metal2 s 106342 -960 106454 480 8 wbs_dat_i[26]
port 459 nsew default input
rlabel metal2 s 109930 -960 110042 480 8 wbs_dat_i[27]
port 460 nsew default input
rlabel metal2 s 113518 -960 113630 480 8 wbs_dat_i[28]
port 461 nsew default input
rlabel metal2 s 117106 -960 117218 480 8 wbs_dat_i[29]
port 462 nsew default input
rlabel metal2 s 18298 -960 18410 480 8 wbs_dat_i[2]
port 463 nsew default input
rlabel metal2 s 120602 -960 120714 480 8 wbs_dat_i[30]
port 464 nsew default input
rlabel metal2 s 124190 -960 124302 480 8 wbs_dat_i[31]
port 465 nsew default input
rlabel metal2 s 23082 -960 23194 480 8 wbs_dat_i[3]
port 466 nsew default input
rlabel metal2 s 27866 -960 27978 480 8 wbs_dat_i[4]
port 467 nsew default input
rlabel metal2 s 31454 -960 31566 480 8 wbs_dat_i[5]
port 468 nsew default input
rlabel metal2 s 34950 -960 35062 480 8 wbs_dat_i[6]
port 469 nsew default input
rlabel metal2 s 38538 -960 38650 480 8 wbs_dat_i[7]
port 470 nsew default input
rlabel metal2 s 42126 -960 42238 480 8 wbs_dat_i[8]
port 471 nsew default input
rlabel metal2 s 45714 -960 45826 480 8 wbs_dat_i[9]
port 472 nsew default input
rlabel metal2 s 10018 -960 10130 480 8 wbs_dat_o[0]
port 473 nsew default tristate
rlabel metal2 s 50498 -960 50610 480 8 wbs_dat_o[10]
port 474 nsew default tristate
rlabel metal2 s 53994 -960 54106 480 8 wbs_dat_o[11]
port 475 nsew default tristate
rlabel metal2 s 57582 -960 57694 480 8 wbs_dat_o[12]
port 476 nsew default tristate
rlabel metal2 s 61170 -960 61282 480 8 wbs_dat_o[13]
port 477 nsew default tristate
rlabel metal2 s 64758 -960 64870 480 8 wbs_dat_o[14]
port 478 nsew default tristate
rlabel metal2 s 68254 -960 68366 480 8 wbs_dat_o[15]
port 479 nsew default tristate
rlabel metal2 s 71842 -960 71954 480 8 wbs_dat_o[16]
port 480 nsew default tristate
rlabel metal2 s 75430 -960 75542 480 8 wbs_dat_o[17]
port 481 nsew default tristate
rlabel metal2 s 79018 -960 79130 480 8 wbs_dat_o[18]
port 482 nsew default tristate
rlabel metal2 s 82606 -960 82718 480 8 wbs_dat_o[19]
port 483 nsew default tristate
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[1]
port 484 nsew default tristate
rlabel metal2 s 86102 -960 86214 480 8 wbs_dat_o[20]
port 485 nsew default tristate
rlabel metal2 s 89690 -960 89802 480 8 wbs_dat_o[21]
port 486 nsew default tristate
rlabel metal2 s 93278 -960 93390 480 8 wbs_dat_o[22]
port 487 nsew default tristate
rlabel metal2 s 96866 -960 96978 480 8 wbs_dat_o[23]
port 488 nsew default tristate
rlabel metal2 s 100454 -960 100566 480 8 wbs_dat_o[24]
port 489 nsew default tristate
rlabel metal2 s 103950 -960 104062 480 8 wbs_dat_o[25]
port 490 nsew default tristate
rlabel metal2 s 107538 -960 107650 480 8 wbs_dat_o[26]
port 491 nsew default tristate
rlabel metal2 s 111126 -960 111238 480 8 wbs_dat_o[27]
port 492 nsew default tristate
rlabel metal2 s 114714 -960 114826 480 8 wbs_dat_o[28]
port 493 nsew default tristate
rlabel metal2 s 118210 -960 118322 480 8 wbs_dat_o[29]
port 494 nsew default tristate
rlabel metal2 s 19494 -960 19606 480 8 wbs_dat_o[2]
port 495 nsew default tristate
rlabel metal2 s 121798 -960 121910 480 8 wbs_dat_o[30]
port 496 nsew default tristate
rlabel metal2 s 125386 -960 125498 480 8 wbs_dat_o[31]
port 497 nsew default tristate
rlabel metal2 s 24278 -960 24390 480 8 wbs_dat_o[3]
port 498 nsew default tristate
rlabel metal2 s 29062 -960 29174 480 8 wbs_dat_o[4]
port 499 nsew default tristate
rlabel metal2 s 32650 -960 32762 480 8 wbs_dat_o[5]
port 500 nsew default tristate
rlabel metal2 s 36146 -960 36258 480 8 wbs_dat_o[6]
port 501 nsew default tristate
rlabel metal2 s 39734 -960 39846 480 8 wbs_dat_o[7]
port 502 nsew default tristate
rlabel metal2 s 43322 -960 43434 480 8 wbs_dat_o[8]
port 503 nsew default tristate
rlabel metal2 s 46910 -960 47022 480 8 wbs_dat_o[9]
port 504 nsew default tristate
rlabel metal2 s 11214 -960 11326 480 8 wbs_sel_i[0]
port 505 nsew default input
rlabel metal2 s 15998 -960 16110 480 8 wbs_sel_i[1]
port 506 nsew default input
rlabel metal2 s 20690 -960 20802 480 8 wbs_sel_i[2]
port 507 nsew default input
rlabel metal2 s 25474 -960 25586 480 8 wbs_sel_i[3]
port 508 nsew default input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 509 nsew default input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 510 nsew default input
rlabel metal2 s 484554 -960 484666 480 8 la_data_out[100]
port 511 nsew default tristate
rlabel metal2 s 488142 -960 488254 480 8 la_data_out[101]
port 512 nsew default tristate
rlabel metal2 s 491730 -960 491842 480 8 la_data_out[102]
port 513 nsew default tristate
rlabel metal2 s 495318 -960 495430 480 8 la_data_out[103]
port 514 nsew default tristate
rlabel metal2 s 498906 -960 499018 480 8 la_data_out[104]
port 515 nsew default tristate
rlabel metal2 s 502402 -960 502514 480 8 la_data_out[105]
port 516 nsew default tristate
rlabel metal2 s 505990 -960 506102 480 8 la_data_out[106]
port 517 nsew default tristate
rlabel metal2 s 509578 -960 509690 480 8 la_data_out[107]
port 518 nsew default tristate
rlabel metal2 s 513166 -960 513278 480 8 la_data_out[108]
port 519 nsew default tristate
rlabel metal2 s 516754 -960 516866 480 8 la_data_out[109]
port 520 nsew default tristate
rlabel metal2 s 163474 -960 163586 480 8 la_data_out[10]
port 521 nsew default tristate
rlabel metal2 s 520250 -960 520362 480 8 la_data_out[110]
port 522 nsew default tristate
rlabel metal2 s 523838 -960 523950 480 8 la_data_out[111]
port 523 nsew default tristate
rlabel metal2 s 527426 -960 527538 480 8 la_data_out[112]
port 524 nsew default tristate
rlabel metal2 s 531014 -960 531126 480 8 la_data_out[113]
port 525 nsew default tristate
rlabel metal2 s 534510 -960 534622 480 8 la_data_out[114]
port 526 nsew default tristate
rlabel metal2 s 538098 -960 538210 480 8 la_data_out[115]
port 527 nsew default tristate
rlabel metal2 s 541686 -960 541798 480 8 la_data_out[116]
port 528 nsew default tristate
rlabel metal2 s 545274 -960 545386 480 8 la_data_out[117]
port 529 nsew default tristate
rlabel metal2 s 548862 -960 548974 480 8 la_data_out[118]
port 530 nsew default tristate
rlabel metal2 s 552358 -960 552470 480 8 la_data_out[119]
port 531 nsew default tristate
rlabel metal2 s 167062 -960 167174 480 8 la_data_out[11]
port 532 nsew default tristate
rlabel metal2 s 555946 -960 556058 480 8 la_data_out[120]
port 533 nsew default tristate
rlabel metal2 s 559534 -960 559646 480 8 la_data_out[121]
port 534 nsew default tristate
rlabel metal2 s 563122 -960 563234 480 8 la_data_out[122]
port 535 nsew default tristate
rlabel metal2 s 566710 -960 566822 480 8 la_data_out[123]
port 536 nsew default tristate
rlabel metal2 s 570206 -960 570318 480 8 la_data_out[124]
port 537 nsew default tristate
rlabel metal2 s 573794 -960 573906 480 8 la_data_out[125]
port 538 nsew default tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[126]
port 539 nsew default tristate
rlabel metal2 s 580970 -960 581082 480 8 la_data_out[127]
port 540 nsew default tristate
rlabel metal2 s 170558 -960 170670 480 8 la_data_out[12]
port 541 nsew default tristate
rlabel metal2 s 174146 -960 174258 480 8 la_data_out[13]
port 542 nsew default tristate
rlabel metal2 s 177734 -960 177846 480 8 la_data_out[14]
port 543 nsew default tristate
rlabel metal2 s 181322 -960 181434 480 8 la_data_out[15]
port 544 nsew default tristate
rlabel metal2 s 184818 -960 184930 480 8 la_data_out[16]
port 545 nsew default tristate
rlabel metal2 s 188406 -960 188518 480 8 la_data_out[17]
port 546 nsew default tristate
rlabel metal2 s 191994 -960 192106 480 8 la_data_out[18]
port 547 nsew default tristate
rlabel metal2 s 195582 -960 195694 480 8 la_data_out[19]
port 548 nsew default tristate
rlabel metal2 s 199170 -960 199282 480 8 la_data_out[20]
port 549 nsew default tristate
rlabel metal2 s 202666 -960 202778 480 8 la_data_out[21]
port 550 nsew default tristate
rlabel metal2 s 206254 -960 206366 480 8 la_data_out[22]
port 551 nsew default tristate
rlabel metal2 s 209842 -960 209954 480 8 la_data_out[23]
port 552 nsew default tristate
rlabel metal2 s 213430 -960 213542 480 8 la_data_out[24]
port 553 nsew default tristate
rlabel metal2 s 217018 -960 217130 480 8 la_data_out[25]
port 554 nsew default tristate
rlabel metal2 s 220514 -960 220626 480 8 la_data_out[26]
port 555 nsew default tristate
rlabel metal2 s 224102 -960 224214 480 8 la_data_out[27]
port 556 nsew default tristate
rlabel metal2 s 227690 -960 227802 480 8 la_data_out[28]
port 557 nsew default tristate
rlabel metal2 s 231278 -960 231390 480 8 la_data_out[29]
port 558 nsew default tristate
rlabel metal2 s 234774 -960 234886 480 8 la_data_out[30]
port 559 nsew default tristate
rlabel metal2 s 238362 -960 238474 480 8 la_data_out[31]
port 560 nsew default tristate
rlabel metal2 s 241950 -960 242062 480 8 la_data_out[32]
port 561 nsew default tristate
rlabel metal2 s 245538 -960 245650 480 8 la_data_out[33]
port 562 nsew default tristate
rlabel metal2 s 249126 -960 249238 480 8 la_data_out[34]
port 563 nsew default tristate
rlabel metal2 s 252622 -960 252734 480 8 la_data_out[35]
port 564 nsew default tristate
rlabel metal2 s 256210 -960 256322 480 8 la_data_out[36]
port 565 nsew default tristate
rlabel metal2 s 259798 -960 259910 480 8 la_data_out[37]
port 566 nsew default tristate
rlabel metal2 s 263386 -960 263498 480 8 la_data_out[38]
port 567 nsew default tristate
rlabel metal2 s 266974 -960 267086 480 8 la_data_out[39]
port 568 nsew default tristate
rlabel metal2 s 138450 -960 138562 480 8 la_data_out[3]
port 569 nsew default tristate
rlabel metal2 s 270470 -960 270582 480 8 la_data_out[40]
port 570 nsew default tristate
rlabel metal2 s 274058 -960 274170 480 8 la_data_out[41]
port 571 nsew default tristate
rlabel metal2 s 277646 -960 277758 480 8 la_data_out[42]
port 572 nsew default tristate
rlabel metal2 s 281234 -960 281346 480 8 la_data_out[43]
port 573 nsew default tristate
rlabel metal2 s 284730 -960 284842 480 8 la_data_out[44]
port 574 nsew default tristate
rlabel metal2 s 288318 -960 288430 480 8 la_data_out[45]
port 575 nsew default tristate
rlabel metal2 s 291906 -960 292018 480 8 la_data_out[46]
port 576 nsew default tristate
rlabel metal2 s 295494 -960 295606 480 8 la_data_out[47]
port 577 nsew default tristate
rlabel metal2 s 299082 -960 299194 480 8 la_data_out[48]
port 578 nsew default tristate
rlabel metal2 s 302578 -960 302690 480 8 la_data_out[49]
port 579 nsew default tristate
rlabel metal2 s 142038 -960 142150 480 8 la_data_out[4]
port 580 nsew default tristate
rlabel metal2 s 306166 -960 306278 480 8 la_data_out[50]
port 581 nsew default tristate
rlabel metal2 s 309754 -960 309866 480 8 la_data_out[51]
port 582 nsew default tristate
rlabel metal2 s 313342 -960 313454 480 8 la_data_out[52]
port 583 nsew default tristate
rlabel metal2 s 316930 -960 317042 480 8 la_data_out[53]
port 584 nsew default tristate
rlabel metal2 s 320426 -960 320538 480 8 la_data_out[54]
port 585 nsew default tristate
rlabel metal2 s 324014 -960 324126 480 8 la_data_out[55]
port 586 nsew default tristate
rlabel metal2 s 327602 -960 327714 480 8 la_data_out[56]
port 587 nsew default tristate
rlabel metal2 s 331190 -960 331302 480 8 la_data_out[57]
port 588 nsew default tristate
rlabel metal2 s 334686 -960 334798 480 8 la_data_out[58]
port 589 nsew default tristate
rlabel metal2 s 338274 -960 338386 480 8 la_data_out[59]
port 590 nsew default tristate
rlabel metal2 s 145626 -960 145738 480 8 la_data_out[5]
port 591 nsew default tristate
rlabel metal2 s 341862 -960 341974 480 8 la_data_out[60]
port 592 nsew default tristate
rlabel metal2 s 345450 -960 345562 480 8 la_data_out[61]
port 593 nsew default tristate
rlabel metal2 s 349038 -960 349150 480 8 la_data_out[62]
port 594 nsew default tristate
rlabel metal2 s 352534 -960 352646 480 8 la_data_out[63]
port 595 nsew default tristate
rlabel metal2 s 356122 -960 356234 480 8 la_data_out[64]
port 596 nsew default tristate
rlabel metal2 s 359710 -960 359822 480 8 la_data_out[65]
port 597 nsew default tristate
rlabel metal2 s 363298 -960 363410 480 8 la_data_out[66]
port 598 nsew default tristate
rlabel metal2 s 366886 -960 366998 480 8 la_data_out[67]
port 599 nsew default tristate
rlabel metal2 s 370382 -960 370494 480 8 la_data_out[68]
port 600 nsew default tristate
rlabel metal2 s 373970 -960 374082 480 8 la_data_out[69]
port 601 nsew default tristate
rlabel metal2 s 149214 -960 149326 480 8 la_data_out[6]
port 602 nsew default tristate
rlabel metal2 s 377558 -960 377670 480 8 la_data_out[70]
port 603 nsew default tristate
rlabel metal2 s 381146 -960 381258 480 8 la_data_out[71]
port 604 nsew default tristate
rlabel metal2 s 384642 -960 384754 480 8 la_data_out[72]
port 605 nsew default tristate
rlabel metal2 s 388230 -960 388342 480 8 la_data_out[73]
port 606 nsew default tristate
rlabel metal2 s 391818 -960 391930 480 8 la_data_out[74]
port 607 nsew default tristate
rlabel metal2 s 395406 -960 395518 480 8 la_data_out[75]
port 608 nsew default tristate
rlabel metal2 s 398994 -960 399106 480 8 la_data_out[76]
port 609 nsew default tristate
rlabel metal2 s 402490 -960 402602 480 8 la_data_out[77]
port 610 nsew default tristate
rlabel metal2 s 406078 -960 406190 480 8 la_data_out[78]
port 611 nsew default tristate
rlabel metal2 s 409666 -960 409778 480 8 la_data_out[79]
port 612 nsew default tristate
rlabel metal2 s 152710 -960 152822 480 8 la_data_out[7]
port 613 nsew default tristate
rlabel metal2 s 413254 -960 413366 480 8 la_data_out[80]
port 614 nsew default tristate
rlabel metal2 s 416842 -960 416954 480 8 la_data_out[81]
port 615 nsew default tristate
rlabel metal2 s 420338 -960 420450 480 8 la_data_out[82]
port 616 nsew default tristate
rlabel metal2 s 423926 -960 424038 480 8 la_data_out[83]
port 617 nsew default tristate
rlabel metal2 s 427514 -960 427626 480 8 la_data_out[84]
port 618 nsew default tristate
rlabel metal2 s 431102 -960 431214 480 8 la_data_out[85]
port 619 nsew default tristate
rlabel metal2 s 434598 -960 434710 480 8 la_data_out[86]
port 620 nsew default tristate
rlabel metal2 s 438186 -960 438298 480 8 la_data_out[87]
port 621 nsew default tristate
rlabel metal2 s 441774 -960 441886 480 8 la_data_out[88]
port 622 nsew default tristate
rlabel metal2 s 445362 -960 445474 480 8 la_data_out[89]
port 623 nsew default tristate
rlabel metal2 s 156298 -960 156410 480 8 la_data_out[8]
port 624 nsew default tristate
rlabel metal2 s 448950 -960 449062 480 8 la_data_out[90]
port 625 nsew default tristate
rlabel metal2 s 452446 -960 452558 480 8 la_data_out[91]
port 626 nsew default tristate
rlabel metal2 s 456034 -960 456146 480 8 la_data_out[92]
port 627 nsew default tristate
rlabel metal2 s 459622 -960 459734 480 8 la_data_out[93]
port 628 nsew default tristate
rlabel metal2 s 463210 -960 463322 480 8 la_data_out[94]
port 629 nsew default tristate
rlabel metal2 s 466798 -960 466910 480 8 la_data_out[95]
port 630 nsew default tristate
rlabel metal2 s 470294 -960 470406 480 8 la_data_out[96]
port 631 nsew default tristate
rlabel metal2 s 473882 -960 473994 480 8 la_data_out[97]
port 632 nsew default tristate
rlabel metal2 s 477470 -960 477582 480 8 la_data_out[98]
port 633 nsew default tristate
rlabel metal2 s 481058 -960 481170 480 8 la_data_out[99]
port 634 nsew default tristate
rlabel metal2 s 159886 -960 159998 480 8 la_data_out[9]
port 635 nsew default tristate
rlabel metal5 s -1996 -924 585920 -324 8 vccd1
port 636 nsew default input
rlabel metal5 s -2936 -1864 586860 -1264 8 vssd1
port 637 nsew default input
rlabel metal5 s -3876 -2804 587800 -2204 8 vccd2
port 638 nsew default input
rlabel metal5 s -4816 -3744 588740 -3144 8 vssd2
port 639 nsew default input
rlabel metal5 s -5756 -4684 589680 -4084 8 vdda1
port 640 nsew default input
rlabel metal5 s -6696 -5624 590620 -5024 8 vssa1
port 641 nsew default input
rlabel metal5 s -7636 -6564 591560 -5964 8 vdda2
port 642 nsew default input
rlabel metal5 s -8576 -7504 592500 -6904 8 vssa2
port 643 nsew default input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
