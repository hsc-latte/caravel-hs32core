magic
tech sky130A
magscale 1 2
timestamp 1608410898
<< obsli1 >>
rect 1104 2159 219023 217617
<< obsm1 >>
rect 14 892 219038 219156
<< metal2 >>
rect 1030 219200 1086 220000
rect 3054 219200 3110 220000
rect 5170 219200 5226 220000
rect 7194 219200 7250 220000
rect 9310 219200 9366 220000
rect 11334 219200 11390 220000
rect 13450 219200 13506 220000
rect 15474 219200 15530 220000
rect 17590 219200 17646 220000
rect 19706 219200 19762 220000
rect 21730 219200 21786 220000
rect 23846 219200 23902 220000
rect 25870 219200 25926 220000
rect 27986 219200 28042 220000
rect 30010 219200 30066 220000
rect 32126 219200 32182 220000
rect 34150 219200 34206 220000
rect 36266 219200 36322 220000
rect 38382 219200 38438 220000
rect 40406 219200 40462 220000
rect 42522 219200 42578 220000
rect 44546 219200 44602 220000
rect 46662 219200 46718 220000
rect 48686 219200 48742 220000
rect 50802 219200 50858 220000
rect 52826 219200 52882 220000
rect 54942 219200 54998 220000
rect 57058 219200 57114 220000
rect 59082 219200 59138 220000
rect 61198 219200 61254 220000
rect 63222 219200 63278 220000
rect 65338 219200 65394 220000
rect 67362 219200 67418 220000
rect 69478 219200 69534 220000
rect 71502 219200 71558 220000
rect 73618 219200 73674 220000
rect 75734 219200 75790 220000
rect 77758 219200 77814 220000
rect 79874 219200 79930 220000
rect 81898 219200 81954 220000
rect 84014 219200 84070 220000
rect 86038 219200 86094 220000
rect 88154 219200 88210 220000
rect 90178 219200 90234 220000
rect 92294 219200 92350 220000
rect 94410 219200 94466 220000
rect 96434 219200 96490 220000
rect 98550 219200 98606 220000
rect 100574 219200 100630 220000
rect 102690 219200 102746 220000
rect 104714 219200 104770 220000
rect 106830 219200 106886 220000
rect 108854 219200 108910 220000
rect 110970 219200 111026 220000
rect 113086 219200 113142 220000
rect 115110 219200 115166 220000
rect 117226 219200 117282 220000
rect 119250 219200 119306 220000
rect 121366 219200 121422 220000
rect 123390 219200 123446 220000
rect 125506 219200 125562 220000
rect 127530 219200 127586 220000
rect 129646 219200 129702 220000
rect 131762 219200 131818 220000
rect 133786 219200 133842 220000
rect 135902 219200 135958 220000
rect 137926 219200 137982 220000
rect 140042 219200 140098 220000
rect 142066 219200 142122 220000
rect 144182 219200 144238 220000
rect 146206 219200 146262 220000
rect 148322 219200 148378 220000
rect 150438 219200 150494 220000
rect 152462 219200 152518 220000
rect 154578 219200 154634 220000
rect 156602 219200 156658 220000
rect 158718 219200 158774 220000
rect 160742 219200 160798 220000
rect 162858 219200 162914 220000
rect 164882 219200 164938 220000
rect 166998 219200 167054 220000
rect 169114 219200 169170 220000
rect 171138 219200 171194 220000
rect 173254 219200 173310 220000
rect 175278 219200 175334 220000
rect 177394 219200 177450 220000
rect 179418 219200 179474 220000
rect 181534 219200 181590 220000
rect 183558 219200 183614 220000
rect 185674 219200 185730 220000
rect 187790 219200 187846 220000
rect 189814 219200 189870 220000
rect 191930 219200 191986 220000
rect 193954 219200 194010 220000
rect 196070 219200 196126 220000
rect 198094 219200 198150 220000
rect 200210 219200 200266 220000
rect 202234 219200 202290 220000
rect 204350 219200 204406 220000
rect 206466 219200 206522 220000
rect 208490 219200 208546 220000
rect 210606 219200 210662 220000
rect 212630 219200 212686 220000
rect 214746 219200 214802 220000
rect 216770 219200 216826 220000
rect 218886 219200 218942 220000
rect 938 0 994 800
rect 2870 0 2926 800
rect 4802 0 4858 800
rect 6734 0 6790 800
rect 8666 0 8722 800
rect 10598 0 10654 800
rect 12530 0 12586 800
rect 14554 0 14610 800
rect 16486 0 16542 800
rect 18418 0 18474 800
rect 20350 0 20406 800
rect 22282 0 22338 800
rect 24214 0 24270 800
rect 26238 0 26294 800
rect 28170 0 28226 800
rect 30102 0 30158 800
rect 32034 0 32090 800
rect 33966 0 34022 800
rect 35898 0 35954 800
rect 37922 0 37978 800
rect 39854 0 39910 800
rect 41786 0 41842 800
rect 43718 0 43774 800
rect 45650 0 45706 800
rect 47582 0 47638 800
rect 49514 0 49570 800
rect 51538 0 51594 800
rect 53470 0 53526 800
rect 55402 0 55458 800
rect 57334 0 57390 800
rect 59266 0 59322 800
rect 61198 0 61254 800
rect 63222 0 63278 800
rect 65154 0 65210 800
rect 67086 0 67142 800
rect 69018 0 69074 800
rect 70950 0 71006 800
rect 72882 0 72938 800
rect 74906 0 74962 800
rect 76838 0 76894 800
rect 78770 0 78826 800
rect 80702 0 80758 800
rect 82634 0 82690 800
rect 84566 0 84622 800
rect 86590 0 86646 800
rect 88522 0 88578 800
rect 90454 0 90510 800
rect 92386 0 92442 800
rect 94318 0 94374 800
rect 96250 0 96306 800
rect 98182 0 98238 800
rect 100206 0 100262 800
rect 102138 0 102194 800
rect 104070 0 104126 800
rect 106002 0 106058 800
rect 107934 0 107990 800
rect 109866 0 109922 800
rect 111890 0 111946 800
rect 113822 0 113878 800
rect 115754 0 115810 800
rect 117686 0 117742 800
rect 119618 0 119674 800
rect 121550 0 121606 800
rect 123574 0 123630 800
rect 125506 0 125562 800
rect 127438 0 127494 800
rect 129370 0 129426 800
rect 131302 0 131358 800
rect 133234 0 133290 800
rect 135166 0 135222 800
rect 137190 0 137246 800
rect 139122 0 139178 800
rect 141054 0 141110 800
rect 142986 0 143042 800
rect 144918 0 144974 800
rect 146850 0 146906 800
rect 148874 0 148930 800
rect 150806 0 150862 800
rect 152738 0 152794 800
rect 154670 0 154726 800
rect 156602 0 156658 800
rect 158534 0 158590 800
rect 160558 0 160614 800
rect 162490 0 162546 800
rect 164422 0 164478 800
rect 166354 0 166410 800
rect 168286 0 168342 800
rect 170218 0 170274 800
rect 172242 0 172298 800
rect 174174 0 174230 800
rect 176106 0 176162 800
rect 178038 0 178094 800
rect 179970 0 180026 800
rect 181902 0 181958 800
rect 183834 0 183890 800
rect 185858 0 185914 800
rect 187790 0 187846 800
rect 189722 0 189778 800
rect 191654 0 191710 800
rect 193586 0 193642 800
rect 195518 0 195574 800
rect 197542 0 197598 800
rect 199474 0 199530 800
rect 201406 0 201462 800
rect 203338 0 203394 800
rect 205270 0 205326 800
rect 207202 0 207258 800
rect 209226 0 209282 800
rect 211158 0 211214 800
rect 213090 0 213146 800
rect 215022 0 215078 800
rect 216954 0 217010 800
rect 218886 0 218942 800
<< obsm2 >>
rect 18 219144 974 219200
rect 1142 219144 2998 219200
rect 3166 219144 5114 219200
rect 5282 219144 7138 219200
rect 7306 219144 9254 219200
rect 9422 219144 11278 219200
rect 11446 219144 13394 219200
rect 13562 219144 15418 219200
rect 15586 219144 17534 219200
rect 17702 219144 19650 219200
rect 19818 219144 21674 219200
rect 21842 219144 23790 219200
rect 23958 219144 25814 219200
rect 25982 219144 27930 219200
rect 28098 219144 29954 219200
rect 30122 219144 32070 219200
rect 32238 219144 34094 219200
rect 34262 219144 36210 219200
rect 36378 219144 38326 219200
rect 38494 219144 40350 219200
rect 40518 219144 42466 219200
rect 42634 219144 44490 219200
rect 44658 219144 46606 219200
rect 46774 219144 48630 219200
rect 48798 219144 50746 219200
rect 50914 219144 52770 219200
rect 52938 219144 54886 219200
rect 55054 219144 57002 219200
rect 57170 219144 59026 219200
rect 59194 219144 61142 219200
rect 61310 219144 63166 219200
rect 63334 219144 65282 219200
rect 65450 219144 67306 219200
rect 67474 219144 69422 219200
rect 69590 219144 71446 219200
rect 71614 219144 73562 219200
rect 73730 219144 75678 219200
rect 75846 219144 77702 219200
rect 77870 219144 79818 219200
rect 79986 219144 81842 219200
rect 82010 219144 83958 219200
rect 84126 219144 85982 219200
rect 86150 219144 88098 219200
rect 88266 219144 90122 219200
rect 90290 219144 92238 219200
rect 92406 219144 94354 219200
rect 94522 219144 96378 219200
rect 96546 219144 98494 219200
rect 98662 219144 100518 219200
rect 100686 219144 102634 219200
rect 102802 219144 104658 219200
rect 104826 219144 106774 219200
rect 106942 219144 108798 219200
rect 108966 219144 110914 219200
rect 111082 219144 113030 219200
rect 113198 219144 115054 219200
rect 115222 219144 117170 219200
rect 117338 219144 119194 219200
rect 119362 219144 121310 219200
rect 121478 219144 123334 219200
rect 123502 219144 125450 219200
rect 125618 219144 127474 219200
rect 127642 219144 129590 219200
rect 129758 219144 131706 219200
rect 131874 219144 133730 219200
rect 133898 219144 135846 219200
rect 136014 219144 137870 219200
rect 138038 219144 139986 219200
rect 140154 219144 142010 219200
rect 142178 219144 144126 219200
rect 144294 219144 146150 219200
rect 146318 219144 148266 219200
rect 148434 219144 150382 219200
rect 150550 219144 152406 219200
rect 152574 219144 154522 219200
rect 154690 219144 156546 219200
rect 156714 219144 158662 219200
rect 158830 219144 160686 219200
rect 160854 219144 162802 219200
rect 162970 219144 164826 219200
rect 164994 219144 166942 219200
rect 167110 219144 169058 219200
rect 169226 219144 171082 219200
rect 171250 219144 173198 219200
rect 173366 219144 175222 219200
rect 175390 219144 177338 219200
rect 177506 219144 179362 219200
rect 179530 219144 181478 219200
rect 181646 219144 183502 219200
rect 183670 219144 185618 219200
rect 185786 219144 187734 219200
rect 187902 219144 189758 219200
rect 189926 219144 191874 219200
rect 192042 219144 193898 219200
rect 194066 219144 196014 219200
rect 196182 219144 198038 219200
rect 198206 219144 200154 219200
rect 200322 219144 202178 219200
rect 202346 219144 204294 219200
rect 204462 219144 206410 219200
rect 206578 219144 208434 219200
rect 208602 219144 210550 219200
rect 210718 219144 212574 219200
rect 212742 219144 214690 219200
rect 214858 219144 216714 219200
rect 216882 219144 218830 219200
rect 218998 219144 219126 219200
rect 18 856 219126 219144
rect 18 439 882 856
rect 1050 439 2814 856
rect 2982 439 4746 856
rect 4914 439 6678 856
rect 6846 439 8610 856
rect 8778 439 10542 856
rect 10710 439 12474 856
rect 12642 439 14498 856
rect 14666 439 16430 856
rect 16598 439 18362 856
rect 18530 439 20294 856
rect 20462 439 22226 856
rect 22394 439 24158 856
rect 24326 439 26182 856
rect 26350 439 28114 856
rect 28282 439 30046 856
rect 30214 439 31978 856
rect 32146 439 33910 856
rect 34078 439 35842 856
rect 36010 439 37866 856
rect 38034 439 39798 856
rect 39966 439 41730 856
rect 41898 439 43662 856
rect 43830 439 45594 856
rect 45762 439 47526 856
rect 47694 439 49458 856
rect 49626 439 51482 856
rect 51650 439 53414 856
rect 53582 439 55346 856
rect 55514 439 57278 856
rect 57446 439 59210 856
rect 59378 439 61142 856
rect 61310 439 63166 856
rect 63334 439 65098 856
rect 65266 439 67030 856
rect 67198 439 68962 856
rect 69130 439 70894 856
rect 71062 439 72826 856
rect 72994 439 74850 856
rect 75018 439 76782 856
rect 76950 439 78714 856
rect 78882 439 80646 856
rect 80814 439 82578 856
rect 82746 439 84510 856
rect 84678 439 86534 856
rect 86702 439 88466 856
rect 88634 439 90398 856
rect 90566 439 92330 856
rect 92498 439 94262 856
rect 94430 439 96194 856
rect 96362 439 98126 856
rect 98294 439 100150 856
rect 100318 439 102082 856
rect 102250 439 104014 856
rect 104182 439 105946 856
rect 106114 439 107878 856
rect 108046 439 109810 856
rect 109978 439 111834 856
rect 112002 439 113766 856
rect 113934 439 115698 856
rect 115866 439 117630 856
rect 117798 439 119562 856
rect 119730 439 121494 856
rect 121662 439 123518 856
rect 123686 439 125450 856
rect 125618 439 127382 856
rect 127550 439 129314 856
rect 129482 439 131246 856
rect 131414 439 133178 856
rect 133346 439 135110 856
rect 135278 439 137134 856
rect 137302 439 139066 856
rect 139234 439 140998 856
rect 141166 439 142930 856
rect 143098 439 144862 856
rect 145030 439 146794 856
rect 146962 439 148818 856
rect 148986 439 150750 856
rect 150918 439 152682 856
rect 152850 439 154614 856
rect 154782 439 156546 856
rect 156714 439 158478 856
rect 158646 439 160502 856
rect 160670 439 162434 856
rect 162602 439 164366 856
rect 164534 439 166298 856
rect 166466 439 168230 856
rect 168398 439 170162 856
rect 170330 439 172186 856
rect 172354 439 174118 856
rect 174286 439 176050 856
rect 176218 439 177982 856
rect 178150 439 179914 856
rect 180082 439 181846 856
rect 182014 439 183778 856
rect 183946 439 185802 856
rect 185970 439 187734 856
rect 187902 439 189666 856
rect 189834 439 191598 856
rect 191766 439 193530 856
rect 193698 439 195462 856
rect 195630 439 197486 856
rect 197654 439 199418 856
rect 199586 439 201350 856
rect 201518 439 203282 856
rect 203450 439 205214 856
rect 205382 439 207146 856
rect 207314 439 209170 856
rect 209338 439 211102 856
rect 211270 439 213034 856
rect 213202 439 214966 856
rect 215134 439 216898 856
rect 217066 439 218830 856
rect 218998 439 219126 856
<< metal3 >>
rect 219200 219376 220000 219496
rect 0 218968 800 219088
rect 219200 218424 220000 218544
rect 219200 217336 220000 217456
rect 0 217064 800 217184
rect 219200 216384 220000 216504
rect 0 215160 800 215280
rect 219200 215296 220000 215416
rect 219200 214344 220000 214464
rect 0 213256 800 213376
rect 219200 213392 220000 213512
rect 219200 212304 220000 212424
rect 0 211352 800 211472
rect 219200 211352 220000 211472
rect 219200 210264 220000 210384
rect 0 209312 800 209432
rect 219200 209312 220000 209432
rect 219200 208224 220000 208344
rect 0 207408 800 207528
rect 219200 207272 220000 207392
rect 219200 206320 220000 206440
rect 0 205504 800 205624
rect 219200 205232 220000 205352
rect 219200 204280 220000 204400
rect 0 203600 800 203720
rect 219200 203192 220000 203312
rect 219200 202240 220000 202360
rect 0 201696 800 201816
rect 219200 201152 220000 201272
rect 219200 200200 220000 200320
rect 0 199656 800 199776
rect 219200 199248 220000 199368
rect 219200 198160 220000 198280
rect 0 197752 800 197872
rect 219200 197208 220000 197328
rect 219200 196120 220000 196240
rect 0 195848 800 195968
rect 219200 195168 220000 195288
rect 219200 194216 220000 194336
rect 0 193944 800 194064
rect 219200 193128 220000 193248
rect 0 192040 800 192160
rect 219200 192176 220000 192296
rect 219200 191088 220000 191208
rect 0 190000 800 190120
rect 219200 190136 220000 190256
rect 219200 189048 220000 189168
rect 0 188096 800 188216
rect 219200 188096 220000 188216
rect 219200 187144 220000 187264
rect 0 186192 800 186312
rect 219200 186056 220000 186176
rect 219200 185104 220000 185224
rect 0 184288 800 184408
rect 219200 184016 220000 184136
rect 219200 183064 220000 183184
rect 0 182384 800 182504
rect 219200 181976 220000 182096
rect 219200 181024 220000 181144
rect 0 180344 800 180464
rect 219200 180072 220000 180192
rect 219200 178984 220000 179104
rect 0 178440 800 178560
rect 219200 178032 220000 178152
rect 219200 176944 220000 177064
rect 0 176536 800 176656
rect 219200 175992 220000 176112
rect 219200 175040 220000 175160
rect 0 174632 800 174752
rect 219200 173952 220000 174072
rect 219200 173000 220000 173120
rect 0 172728 800 172848
rect 219200 171912 220000 172032
rect 219200 170960 220000 171080
rect 0 170688 800 170808
rect 219200 169872 220000 169992
rect 0 168784 800 168904
rect 219200 168920 220000 169040
rect 219200 167968 220000 168088
rect 0 166880 800 167000
rect 219200 166880 220000 167000
rect 219200 165928 220000 166048
rect 0 164976 800 165096
rect 219200 164840 220000 164960
rect 219200 163888 220000 164008
rect 0 163072 800 163192
rect 219200 162800 220000 162920
rect 219200 161848 220000 161968
rect 0 161168 800 161288
rect 219200 160896 220000 161016
rect 219200 159808 220000 159928
rect 0 159128 800 159248
rect 219200 158856 220000 158976
rect 219200 157768 220000 157888
rect 0 157224 800 157344
rect 219200 156816 220000 156936
rect 219200 155728 220000 155848
rect 0 155320 800 155440
rect 219200 154776 220000 154896
rect 219200 153824 220000 153944
rect 0 153416 800 153536
rect 219200 152736 220000 152856
rect 219200 151784 220000 151904
rect 0 151512 800 151632
rect 219200 150696 220000 150816
rect 219200 149744 220000 149864
rect 0 149472 800 149592
rect 219200 148792 220000 148912
rect 0 147568 800 147688
rect 219200 147704 220000 147824
rect 219200 146752 220000 146872
rect 0 145664 800 145784
rect 219200 145664 220000 145784
rect 219200 144712 220000 144832
rect 0 143760 800 143880
rect 219200 143624 220000 143744
rect 219200 142672 220000 142792
rect 0 141856 800 141976
rect 219200 141720 220000 141840
rect 219200 140632 220000 140752
rect 0 139816 800 139936
rect 219200 139680 220000 139800
rect 219200 138592 220000 138712
rect 0 137912 800 138032
rect 219200 137640 220000 137760
rect 219200 136552 220000 136672
rect 0 136008 800 136128
rect 219200 135600 220000 135720
rect 219200 134648 220000 134768
rect 0 134104 800 134224
rect 219200 133560 220000 133680
rect 219200 132608 220000 132728
rect 0 132200 800 132320
rect 219200 131520 220000 131640
rect 219200 130568 220000 130688
rect 0 130160 800 130280
rect 219200 129616 220000 129736
rect 219200 128528 220000 128648
rect 0 128256 800 128376
rect 219200 127576 220000 127696
rect 0 126352 800 126472
rect 219200 126488 220000 126608
rect 219200 125536 220000 125656
rect 0 124448 800 124568
rect 219200 124448 220000 124568
rect 219200 123496 220000 123616
rect 0 122544 800 122664
rect 219200 122544 220000 122664
rect 219200 121456 220000 121576
rect 0 120504 800 120624
rect 219200 120504 220000 120624
rect 219200 119416 220000 119536
rect 0 118600 800 118720
rect 219200 118464 220000 118584
rect 219200 117376 220000 117496
rect 0 116696 800 116816
rect 219200 116424 220000 116544
rect 219200 115472 220000 115592
rect 0 114792 800 114912
rect 219200 114384 220000 114504
rect 219200 113432 220000 113552
rect 0 112888 800 113008
rect 219200 112344 220000 112464
rect 219200 111392 220000 111512
rect 0 110984 800 111104
rect 219200 110440 220000 110560
rect 219200 109352 220000 109472
rect 0 108944 800 109064
rect 219200 108400 220000 108520
rect 219200 107312 220000 107432
rect 0 107040 800 107160
rect 219200 106360 220000 106480
rect 0 105136 800 105256
rect 219200 105272 220000 105392
rect 219200 104320 220000 104440
rect 0 103232 800 103352
rect 219200 103368 220000 103488
rect 219200 102280 220000 102400
rect 0 101328 800 101448
rect 219200 101328 220000 101448
rect 219200 100240 220000 100360
rect 0 99288 800 99408
rect 219200 99288 220000 99408
rect 219200 98200 220000 98320
rect 0 97384 800 97504
rect 219200 97248 220000 97368
rect 219200 96296 220000 96416
rect 0 95480 800 95600
rect 219200 95208 220000 95328
rect 219200 94256 220000 94376
rect 0 93576 800 93696
rect 219200 93168 220000 93288
rect 219200 92216 220000 92336
rect 0 91672 800 91792
rect 219200 91128 220000 91248
rect 219200 90176 220000 90296
rect 0 89632 800 89752
rect 219200 89224 220000 89344
rect 219200 88136 220000 88256
rect 0 87728 800 87848
rect 219200 87184 220000 87304
rect 219200 86096 220000 86216
rect 0 85824 800 85944
rect 219200 85144 220000 85264
rect 219200 84192 220000 84312
rect 0 83920 800 84040
rect 219200 83104 220000 83224
rect 0 82016 800 82136
rect 219200 82152 220000 82272
rect 219200 81064 220000 81184
rect 0 79976 800 80096
rect 219200 80112 220000 80232
rect 219200 79024 220000 79144
rect 0 78072 800 78192
rect 219200 78072 220000 78192
rect 219200 77120 220000 77240
rect 0 76168 800 76288
rect 219200 76032 220000 76152
rect 219200 75080 220000 75200
rect 0 74264 800 74384
rect 219200 73992 220000 74112
rect 219200 73040 220000 73160
rect 0 72360 800 72480
rect 219200 71952 220000 72072
rect 219200 71000 220000 71120
rect 0 70320 800 70440
rect 219200 70048 220000 70168
rect 219200 68960 220000 69080
rect 0 68416 800 68536
rect 219200 68008 220000 68128
rect 219200 66920 220000 67040
rect 0 66512 800 66632
rect 219200 65968 220000 66088
rect 219200 65016 220000 65136
rect 0 64608 800 64728
rect 219200 63928 220000 64048
rect 219200 62976 220000 63096
rect 0 62704 800 62824
rect 219200 61888 220000 62008
rect 219200 60936 220000 61056
rect 0 60664 800 60784
rect 219200 59848 220000 59968
rect 0 58760 800 58880
rect 219200 58896 220000 59016
rect 219200 57944 220000 58064
rect 0 56856 800 56976
rect 219200 56856 220000 56976
rect 219200 55904 220000 56024
rect 0 54952 800 55072
rect 219200 54816 220000 54936
rect 219200 53864 220000 53984
rect 0 53048 800 53168
rect 219200 52776 220000 52896
rect 219200 51824 220000 51944
rect 0 51144 800 51264
rect 219200 50872 220000 50992
rect 219200 49784 220000 49904
rect 0 49104 800 49224
rect 219200 48832 220000 48952
rect 219200 47744 220000 47864
rect 0 47200 800 47320
rect 219200 46792 220000 46912
rect 219200 45704 220000 45824
rect 0 45296 800 45416
rect 219200 44752 220000 44872
rect 219200 43800 220000 43920
rect 0 43392 800 43512
rect 219200 42712 220000 42832
rect 219200 41760 220000 41880
rect 0 41488 800 41608
rect 219200 40672 220000 40792
rect 219200 39720 220000 39840
rect 0 39448 800 39568
rect 219200 38768 220000 38888
rect 0 37544 800 37664
rect 219200 37680 220000 37800
rect 219200 36728 220000 36848
rect 0 35640 800 35760
rect 219200 35640 220000 35760
rect 219200 34688 220000 34808
rect 0 33736 800 33856
rect 219200 33600 220000 33720
rect 219200 32648 220000 32768
rect 0 31832 800 31952
rect 219200 31696 220000 31816
rect 219200 30608 220000 30728
rect 0 29792 800 29912
rect 219200 29656 220000 29776
rect 219200 28568 220000 28688
rect 0 27888 800 28008
rect 219200 27616 220000 27736
rect 219200 26528 220000 26648
rect 0 25984 800 26104
rect 219200 25576 220000 25696
rect 219200 24624 220000 24744
rect 0 24080 800 24200
rect 219200 23536 220000 23656
rect 219200 22584 220000 22704
rect 0 22176 800 22296
rect 219200 21496 220000 21616
rect 219200 20544 220000 20664
rect 0 20136 800 20256
rect 219200 19592 220000 19712
rect 219200 18504 220000 18624
rect 0 18232 800 18352
rect 219200 17552 220000 17672
rect 0 16328 800 16448
rect 219200 16464 220000 16584
rect 219200 15512 220000 15632
rect 0 14424 800 14544
rect 219200 14424 220000 14544
rect 219200 13472 220000 13592
rect 0 12520 800 12640
rect 219200 12520 220000 12640
rect 219200 11432 220000 11552
rect 0 10480 800 10600
rect 219200 10480 220000 10600
rect 219200 9392 220000 9512
rect 0 8576 800 8696
rect 219200 8440 220000 8560
rect 219200 7352 220000 7472
rect 0 6672 800 6792
rect 219200 6400 220000 6520
rect 219200 5448 220000 5568
rect 0 4768 800 4888
rect 219200 4360 220000 4480
rect 219200 3408 220000 3528
rect 0 2864 800 2984
rect 219200 2320 220000 2440
rect 219200 1368 220000 1488
rect 0 960 800 1080
rect 219200 416 220000 536
<< obsm3 >>
rect 13 219296 219120 219468
rect 13 219168 219200 219296
rect 880 218888 219200 219168
rect 13 218624 219200 218888
rect 13 218344 219120 218624
rect 13 217536 219200 218344
rect 13 217264 219120 217536
rect 880 217256 219120 217264
rect 880 216984 219200 217256
rect 13 216584 219200 216984
rect 13 216304 219120 216584
rect 13 215496 219200 216304
rect 13 215360 219120 215496
rect 880 215216 219120 215360
rect 880 215080 219200 215216
rect 13 214544 219200 215080
rect 13 214264 219120 214544
rect 13 213592 219200 214264
rect 13 213456 219120 213592
rect 880 213312 219120 213456
rect 880 213176 219200 213312
rect 13 212504 219200 213176
rect 13 212224 219120 212504
rect 13 211552 219200 212224
rect 880 211272 219120 211552
rect 13 210464 219200 211272
rect 13 210184 219120 210464
rect 13 209512 219200 210184
rect 880 209232 219120 209512
rect 13 208424 219200 209232
rect 13 208144 219120 208424
rect 13 207608 219200 208144
rect 880 207472 219200 207608
rect 880 207328 219120 207472
rect 13 207192 219120 207328
rect 13 206520 219200 207192
rect 13 206240 219120 206520
rect 13 205704 219200 206240
rect 880 205432 219200 205704
rect 880 205424 219120 205432
rect 13 205152 219120 205424
rect 13 204480 219200 205152
rect 13 204200 219120 204480
rect 13 203800 219200 204200
rect 880 203520 219200 203800
rect 13 203392 219200 203520
rect 13 203112 219120 203392
rect 13 202440 219200 203112
rect 13 202160 219120 202440
rect 13 201896 219200 202160
rect 880 201616 219200 201896
rect 13 201352 219200 201616
rect 13 201072 219120 201352
rect 13 200400 219200 201072
rect 13 200120 219120 200400
rect 13 199856 219200 200120
rect 880 199576 219200 199856
rect 13 199448 219200 199576
rect 13 199168 219120 199448
rect 13 198360 219200 199168
rect 13 198080 219120 198360
rect 13 197952 219200 198080
rect 880 197672 219200 197952
rect 13 197408 219200 197672
rect 13 197128 219120 197408
rect 13 196320 219200 197128
rect 13 196048 219120 196320
rect 880 196040 219120 196048
rect 880 195768 219200 196040
rect 13 195368 219200 195768
rect 13 195088 219120 195368
rect 13 194416 219200 195088
rect 13 194144 219120 194416
rect 880 194136 219120 194144
rect 880 193864 219200 194136
rect 13 193328 219200 193864
rect 13 193048 219120 193328
rect 13 192376 219200 193048
rect 13 192240 219120 192376
rect 880 192096 219120 192240
rect 880 191960 219200 192096
rect 13 191288 219200 191960
rect 13 191008 219120 191288
rect 13 190336 219200 191008
rect 13 190200 219120 190336
rect 880 190056 219120 190200
rect 880 189920 219200 190056
rect 13 189248 219200 189920
rect 13 188968 219120 189248
rect 13 188296 219200 188968
rect 880 188016 219120 188296
rect 13 187344 219200 188016
rect 13 187064 219120 187344
rect 13 186392 219200 187064
rect 880 186256 219200 186392
rect 880 186112 219120 186256
rect 13 185976 219120 186112
rect 13 185304 219200 185976
rect 13 185024 219120 185304
rect 13 184488 219200 185024
rect 880 184216 219200 184488
rect 880 184208 219120 184216
rect 13 183936 219120 184208
rect 13 183264 219200 183936
rect 13 182984 219120 183264
rect 13 182584 219200 182984
rect 880 182304 219200 182584
rect 13 182176 219200 182304
rect 13 181896 219120 182176
rect 13 181224 219200 181896
rect 13 180944 219120 181224
rect 13 180544 219200 180944
rect 880 180272 219200 180544
rect 880 180264 219120 180272
rect 13 179992 219120 180264
rect 13 179184 219200 179992
rect 13 178904 219120 179184
rect 13 178640 219200 178904
rect 880 178360 219200 178640
rect 13 178232 219200 178360
rect 13 177952 219120 178232
rect 13 177144 219200 177952
rect 13 176864 219120 177144
rect 13 176736 219200 176864
rect 880 176456 219200 176736
rect 13 176192 219200 176456
rect 13 175912 219120 176192
rect 13 175240 219200 175912
rect 13 174960 219120 175240
rect 13 174832 219200 174960
rect 880 174552 219200 174832
rect 13 174152 219200 174552
rect 13 173872 219120 174152
rect 13 173200 219200 173872
rect 13 172928 219120 173200
rect 880 172920 219120 172928
rect 880 172648 219200 172920
rect 13 172112 219200 172648
rect 13 171832 219120 172112
rect 13 171160 219200 171832
rect 13 170888 219120 171160
rect 880 170880 219120 170888
rect 880 170608 219200 170880
rect 13 170072 219200 170608
rect 13 169792 219120 170072
rect 13 169120 219200 169792
rect 13 168984 219120 169120
rect 880 168840 219120 168984
rect 880 168704 219200 168840
rect 13 168168 219200 168704
rect 13 167888 219120 168168
rect 13 167080 219200 167888
rect 880 166800 219120 167080
rect 13 166128 219200 166800
rect 13 165848 219120 166128
rect 13 165176 219200 165848
rect 880 165040 219200 165176
rect 880 164896 219120 165040
rect 13 164760 219120 164896
rect 13 164088 219200 164760
rect 13 163808 219120 164088
rect 13 163272 219200 163808
rect 880 163000 219200 163272
rect 880 162992 219120 163000
rect 13 162720 219120 162992
rect 13 162048 219200 162720
rect 13 161768 219120 162048
rect 13 161368 219200 161768
rect 880 161096 219200 161368
rect 880 161088 219120 161096
rect 13 160816 219120 161088
rect 13 160008 219200 160816
rect 13 159728 219120 160008
rect 13 159328 219200 159728
rect 880 159056 219200 159328
rect 880 159048 219120 159056
rect 13 158776 219120 159048
rect 13 157968 219200 158776
rect 13 157688 219120 157968
rect 13 157424 219200 157688
rect 880 157144 219200 157424
rect 13 157016 219200 157144
rect 13 156736 219120 157016
rect 13 155928 219200 156736
rect 13 155648 219120 155928
rect 13 155520 219200 155648
rect 880 155240 219200 155520
rect 13 154976 219200 155240
rect 13 154696 219120 154976
rect 13 154024 219200 154696
rect 13 153744 219120 154024
rect 13 153616 219200 153744
rect 880 153336 219200 153616
rect 13 152936 219200 153336
rect 13 152656 219120 152936
rect 13 151984 219200 152656
rect 13 151712 219120 151984
rect 880 151704 219120 151712
rect 880 151432 219200 151704
rect 13 150896 219200 151432
rect 13 150616 219120 150896
rect 13 149944 219200 150616
rect 13 149672 219120 149944
rect 880 149664 219120 149672
rect 880 149392 219200 149664
rect 13 148992 219200 149392
rect 13 148712 219120 148992
rect 13 147904 219200 148712
rect 13 147768 219120 147904
rect 880 147624 219120 147768
rect 880 147488 219200 147624
rect 13 146952 219200 147488
rect 13 146672 219120 146952
rect 13 145864 219200 146672
rect 880 145584 219120 145864
rect 13 144912 219200 145584
rect 13 144632 219120 144912
rect 13 143960 219200 144632
rect 880 143824 219200 143960
rect 880 143680 219120 143824
rect 13 143544 219120 143680
rect 13 142872 219200 143544
rect 13 142592 219120 142872
rect 13 142056 219200 142592
rect 880 141920 219200 142056
rect 880 141776 219120 141920
rect 13 141640 219120 141776
rect 13 140832 219200 141640
rect 13 140552 219120 140832
rect 13 140016 219200 140552
rect 880 139880 219200 140016
rect 880 139736 219120 139880
rect 13 139600 219120 139736
rect 13 138792 219200 139600
rect 13 138512 219120 138792
rect 13 138112 219200 138512
rect 880 137840 219200 138112
rect 880 137832 219120 137840
rect 13 137560 219120 137832
rect 13 136752 219200 137560
rect 13 136472 219120 136752
rect 13 136208 219200 136472
rect 880 135928 219200 136208
rect 13 135800 219200 135928
rect 13 135520 219120 135800
rect 13 134848 219200 135520
rect 13 134568 219120 134848
rect 13 134304 219200 134568
rect 880 134024 219200 134304
rect 13 133760 219200 134024
rect 13 133480 219120 133760
rect 13 132808 219200 133480
rect 13 132528 219120 132808
rect 13 132400 219200 132528
rect 880 132120 219200 132400
rect 13 131720 219200 132120
rect 13 131440 219120 131720
rect 13 130768 219200 131440
rect 13 130488 219120 130768
rect 13 130360 219200 130488
rect 880 130080 219200 130360
rect 13 129816 219200 130080
rect 13 129536 219120 129816
rect 13 128728 219200 129536
rect 13 128456 219120 128728
rect 880 128448 219120 128456
rect 880 128176 219200 128448
rect 13 127776 219200 128176
rect 13 127496 219120 127776
rect 13 126688 219200 127496
rect 13 126552 219120 126688
rect 880 126408 219120 126552
rect 880 126272 219200 126408
rect 13 125736 219200 126272
rect 13 125456 219120 125736
rect 13 124648 219200 125456
rect 880 124368 219120 124648
rect 13 123696 219200 124368
rect 13 123416 219120 123696
rect 13 122744 219200 123416
rect 880 122464 219120 122744
rect 13 121656 219200 122464
rect 13 121376 219120 121656
rect 13 120704 219200 121376
rect 880 120424 219120 120704
rect 13 119616 219200 120424
rect 13 119336 219120 119616
rect 13 118800 219200 119336
rect 880 118664 219200 118800
rect 880 118520 219120 118664
rect 13 118384 219120 118520
rect 13 117576 219200 118384
rect 13 117296 219120 117576
rect 13 116896 219200 117296
rect 880 116624 219200 116896
rect 880 116616 219120 116624
rect 13 116344 219120 116616
rect 13 115672 219200 116344
rect 13 115392 219120 115672
rect 13 114992 219200 115392
rect 880 114712 219200 114992
rect 13 114584 219200 114712
rect 13 114304 219120 114584
rect 13 113632 219200 114304
rect 13 113352 219120 113632
rect 13 113088 219200 113352
rect 880 112808 219200 113088
rect 13 112544 219200 112808
rect 13 112264 219120 112544
rect 13 111592 219200 112264
rect 13 111312 219120 111592
rect 13 111184 219200 111312
rect 880 110904 219200 111184
rect 13 110640 219200 110904
rect 13 110360 219120 110640
rect 13 109552 219200 110360
rect 13 109272 219120 109552
rect 13 109144 219200 109272
rect 880 108864 219200 109144
rect 13 108600 219200 108864
rect 13 108320 219120 108600
rect 13 107512 219200 108320
rect 13 107240 219120 107512
rect 880 107232 219120 107240
rect 880 106960 219200 107232
rect 13 106560 219200 106960
rect 13 106280 219120 106560
rect 13 105472 219200 106280
rect 13 105336 219120 105472
rect 880 105192 219120 105336
rect 880 105056 219200 105192
rect 13 104520 219200 105056
rect 13 104240 219120 104520
rect 13 103568 219200 104240
rect 13 103432 219120 103568
rect 880 103288 219120 103432
rect 880 103152 219200 103288
rect 13 102480 219200 103152
rect 13 102200 219120 102480
rect 13 101528 219200 102200
rect 880 101248 219120 101528
rect 13 100440 219200 101248
rect 13 100160 219120 100440
rect 13 99488 219200 100160
rect 880 99208 219120 99488
rect 13 98400 219200 99208
rect 13 98120 219120 98400
rect 13 97584 219200 98120
rect 880 97448 219200 97584
rect 880 97304 219120 97448
rect 13 97168 219120 97304
rect 13 96496 219200 97168
rect 13 96216 219120 96496
rect 13 95680 219200 96216
rect 880 95408 219200 95680
rect 880 95400 219120 95408
rect 13 95128 219120 95400
rect 13 94456 219200 95128
rect 13 94176 219120 94456
rect 13 93776 219200 94176
rect 880 93496 219200 93776
rect 13 93368 219200 93496
rect 13 93088 219120 93368
rect 13 92416 219200 93088
rect 13 92136 219120 92416
rect 13 91872 219200 92136
rect 880 91592 219200 91872
rect 13 91328 219200 91592
rect 13 91048 219120 91328
rect 13 90376 219200 91048
rect 13 90096 219120 90376
rect 13 89832 219200 90096
rect 880 89552 219200 89832
rect 13 89424 219200 89552
rect 13 89144 219120 89424
rect 13 88336 219200 89144
rect 13 88056 219120 88336
rect 13 87928 219200 88056
rect 880 87648 219200 87928
rect 13 87384 219200 87648
rect 13 87104 219120 87384
rect 13 86296 219200 87104
rect 13 86024 219120 86296
rect 880 86016 219120 86024
rect 880 85744 219200 86016
rect 13 85344 219200 85744
rect 13 85064 219120 85344
rect 13 84392 219200 85064
rect 13 84120 219120 84392
rect 880 84112 219120 84120
rect 880 83840 219200 84112
rect 13 83304 219200 83840
rect 13 83024 219120 83304
rect 13 82352 219200 83024
rect 13 82216 219120 82352
rect 880 82072 219120 82216
rect 880 81936 219200 82072
rect 13 81264 219200 81936
rect 13 80984 219120 81264
rect 13 80312 219200 80984
rect 13 80176 219120 80312
rect 880 80032 219120 80176
rect 880 79896 219200 80032
rect 13 79224 219200 79896
rect 13 78944 219120 79224
rect 13 78272 219200 78944
rect 880 77992 219120 78272
rect 13 77320 219200 77992
rect 13 77040 219120 77320
rect 13 76368 219200 77040
rect 880 76232 219200 76368
rect 880 76088 219120 76232
rect 13 75952 219120 76088
rect 13 75280 219200 75952
rect 13 75000 219120 75280
rect 13 74464 219200 75000
rect 880 74192 219200 74464
rect 880 74184 219120 74192
rect 13 73912 219120 74184
rect 13 73240 219200 73912
rect 13 72960 219120 73240
rect 13 72560 219200 72960
rect 880 72280 219200 72560
rect 13 72152 219200 72280
rect 13 71872 219120 72152
rect 13 71200 219200 71872
rect 13 70920 219120 71200
rect 13 70520 219200 70920
rect 880 70248 219200 70520
rect 880 70240 219120 70248
rect 13 69968 219120 70240
rect 13 69160 219200 69968
rect 13 68880 219120 69160
rect 13 68616 219200 68880
rect 880 68336 219200 68616
rect 13 68208 219200 68336
rect 13 67928 219120 68208
rect 13 67120 219200 67928
rect 13 66840 219120 67120
rect 13 66712 219200 66840
rect 880 66432 219200 66712
rect 13 66168 219200 66432
rect 13 65888 219120 66168
rect 13 65216 219200 65888
rect 13 64936 219120 65216
rect 13 64808 219200 64936
rect 880 64528 219200 64808
rect 13 64128 219200 64528
rect 13 63848 219120 64128
rect 13 63176 219200 63848
rect 13 62904 219120 63176
rect 880 62896 219120 62904
rect 880 62624 219200 62896
rect 13 62088 219200 62624
rect 13 61808 219120 62088
rect 13 61136 219200 61808
rect 13 60864 219120 61136
rect 880 60856 219120 60864
rect 880 60584 219200 60856
rect 13 60048 219200 60584
rect 13 59768 219120 60048
rect 13 59096 219200 59768
rect 13 58960 219120 59096
rect 880 58816 219120 58960
rect 880 58680 219200 58816
rect 13 58144 219200 58680
rect 13 57864 219120 58144
rect 13 57056 219200 57864
rect 880 56776 219120 57056
rect 13 56104 219200 56776
rect 13 55824 219120 56104
rect 13 55152 219200 55824
rect 880 55016 219200 55152
rect 880 54872 219120 55016
rect 13 54736 219120 54872
rect 13 54064 219200 54736
rect 13 53784 219120 54064
rect 13 53248 219200 53784
rect 880 52976 219200 53248
rect 880 52968 219120 52976
rect 13 52696 219120 52968
rect 13 52024 219200 52696
rect 13 51744 219120 52024
rect 13 51344 219200 51744
rect 880 51072 219200 51344
rect 880 51064 219120 51072
rect 13 50792 219120 51064
rect 13 49984 219200 50792
rect 13 49704 219120 49984
rect 13 49304 219200 49704
rect 880 49032 219200 49304
rect 880 49024 219120 49032
rect 13 48752 219120 49024
rect 13 47944 219200 48752
rect 13 47664 219120 47944
rect 13 47400 219200 47664
rect 880 47120 219200 47400
rect 13 46992 219200 47120
rect 13 46712 219120 46992
rect 13 45904 219200 46712
rect 13 45624 219120 45904
rect 13 45496 219200 45624
rect 880 45216 219200 45496
rect 13 44952 219200 45216
rect 13 44672 219120 44952
rect 13 44000 219200 44672
rect 13 43720 219120 44000
rect 13 43592 219200 43720
rect 880 43312 219200 43592
rect 13 42912 219200 43312
rect 13 42632 219120 42912
rect 13 41960 219200 42632
rect 13 41688 219120 41960
rect 880 41680 219120 41688
rect 880 41408 219200 41680
rect 13 40872 219200 41408
rect 13 40592 219120 40872
rect 13 39920 219200 40592
rect 13 39648 219120 39920
rect 880 39640 219120 39648
rect 880 39368 219200 39640
rect 13 38968 219200 39368
rect 13 38688 219120 38968
rect 13 37880 219200 38688
rect 13 37744 219120 37880
rect 880 37600 219120 37744
rect 880 37464 219200 37600
rect 13 36928 219200 37464
rect 13 36648 219120 36928
rect 13 35840 219200 36648
rect 880 35560 219120 35840
rect 13 34888 219200 35560
rect 13 34608 219120 34888
rect 13 33936 219200 34608
rect 880 33800 219200 33936
rect 880 33656 219120 33800
rect 13 33520 219120 33656
rect 13 32848 219200 33520
rect 13 32568 219120 32848
rect 13 32032 219200 32568
rect 880 31896 219200 32032
rect 880 31752 219120 31896
rect 13 31616 219120 31752
rect 13 30808 219200 31616
rect 13 30528 219120 30808
rect 13 29992 219200 30528
rect 880 29856 219200 29992
rect 880 29712 219120 29856
rect 13 29576 219120 29712
rect 13 28768 219200 29576
rect 13 28488 219120 28768
rect 13 28088 219200 28488
rect 880 27816 219200 28088
rect 880 27808 219120 27816
rect 13 27536 219120 27808
rect 13 26728 219200 27536
rect 13 26448 219120 26728
rect 13 26184 219200 26448
rect 880 25904 219200 26184
rect 13 25776 219200 25904
rect 13 25496 219120 25776
rect 13 24824 219200 25496
rect 13 24544 219120 24824
rect 13 24280 219200 24544
rect 880 24000 219200 24280
rect 13 23736 219200 24000
rect 13 23456 219120 23736
rect 13 22784 219200 23456
rect 13 22504 219120 22784
rect 13 22376 219200 22504
rect 880 22096 219200 22376
rect 13 21696 219200 22096
rect 13 21416 219120 21696
rect 13 20744 219200 21416
rect 13 20464 219120 20744
rect 13 20336 219200 20464
rect 880 20056 219200 20336
rect 13 19792 219200 20056
rect 13 19512 219120 19792
rect 13 18704 219200 19512
rect 13 18432 219120 18704
rect 880 18424 219120 18432
rect 880 18152 219200 18424
rect 13 17752 219200 18152
rect 13 17472 219120 17752
rect 13 16664 219200 17472
rect 13 16528 219120 16664
rect 880 16384 219120 16528
rect 880 16248 219200 16384
rect 13 15712 219200 16248
rect 13 15432 219120 15712
rect 13 14624 219200 15432
rect 880 14344 219120 14624
rect 13 13672 219200 14344
rect 13 13392 219120 13672
rect 13 12720 219200 13392
rect 880 12440 219120 12720
rect 13 11632 219200 12440
rect 13 11352 219120 11632
rect 13 10680 219200 11352
rect 880 10400 219120 10680
rect 13 9592 219200 10400
rect 13 9312 219120 9592
rect 13 8776 219200 9312
rect 880 8640 219200 8776
rect 880 8496 219120 8640
rect 13 8360 219120 8496
rect 13 7552 219200 8360
rect 13 7272 219120 7552
rect 13 6872 219200 7272
rect 880 6600 219200 6872
rect 880 6592 219120 6600
rect 13 6320 219120 6592
rect 13 5648 219200 6320
rect 13 5368 219120 5648
rect 13 4968 219200 5368
rect 880 4688 219200 4968
rect 13 4560 219200 4688
rect 13 4280 219120 4560
rect 13 3608 219200 4280
rect 13 3328 219120 3608
rect 13 3064 219200 3328
rect 880 2784 219200 3064
rect 13 2520 219200 2784
rect 13 2240 219120 2520
rect 13 1568 219200 2240
rect 13 1288 219120 1568
rect 13 1160 219200 1288
rect 880 880 219200 1160
rect 13 616 219200 880
rect 13 443 219120 616
<< metal4 >>
rect 4208 2128 4528 217648
rect 19568 2128 19888 217648
<< obsm4 >>
rect 4659 217728 217981 219469
rect 4659 2048 19488 217728
rect 19968 2048 217981 217728
rect 4659 1395 217981 2048
<< labels >>
rlabel metal3 s 219200 13472 220000 13592 6 cpu_addr_e[0]
port 1 nsew default output
rlabel metal3 s 219200 23536 220000 23656 6 cpu_addr_e[10]
port 2 nsew default output
rlabel metal3 s 219200 24624 220000 24744 6 cpu_addr_e[11]
port 3 nsew default output
rlabel metal3 s 219200 25576 220000 25696 6 cpu_addr_e[12]
port 4 nsew default output
rlabel metal3 s 219200 26528 220000 26648 6 cpu_addr_e[13]
port 5 nsew default output
rlabel metal3 s 219200 27616 220000 27736 6 cpu_addr_e[14]
port 6 nsew default output
rlabel metal3 s 219200 28568 220000 28688 6 cpu_addr_e[15]
port 7 nsew default output
rlabel metal3 s 219200 14424 220000 14544 6 cpu_addr_e[1]
port 8 nsew default output
rlabel metal3 s 219200 15512 220000 15632 6 cpu_addr_e[2]
port 9 nsew default output
rlabel metal3 s 219200 16464 220000 16584 6 cpu_addr_e[3]
port 10 nsew default output
rlabel metal3 s 219200 17552 220000 17672 6 cpu_addr_e[4]
port 11 nsew default output
rlabel metal3 s 219200 18504 220000 18624 6 cpu_addr_e[5]
port 12 nsew default output
rlabel metal3 s 219200 19592 220000 19712 6 cpu_addr_e[6]
port 13 nsew default output
rlabel metal3 s 219200 20544 220000 20664 6 cpu_addr_e[7]
port 14 nsew default output
rlabel metal3 s 219200 21496 220000 21616 6 cpu_addr_e[8]
port 15 nsew default output
rlabel metal3 s 219200 22584 220000 22704 6 cpu_addr_e[9]
port 16 nsew default output
rlabel metal2 s 21730 219200 21786 220000 6 cpu_addr_n[0]
port 17 nsew default output
rlabel metal2 s 42522 219200 42578 220000 6 cpu_addr_n[10]
port 18 nsew default output
rlabel metal2 s 44546 219200 44602 220000 6 cpu_addr_n[11]
port 19 nsew default output
rlabel metal2 s 46662 219200 46718 220000 6 cpu_addr_n[12]
port 20 nsew default output
rlabel metal2 s 48686 219200 48742 220000 6 cpu_addr_n[13]
port 21 nsew default output
rlabel metal2 s 50802 219200 50858 220000 6 cpu_addr_n[14]
port 22 nsew default output
rlabel metal2 s 52826 219200 52882 220000 6 cpu_addr_n[15]
port 23 nsew default output
rlabel metal2 s 23846 219200 23902 220000 6 cpu_addr_n[1]
port 24 nsew default output
rlabel metal2 s 25870 219200 25926 220000 6 cpu_addr_n[2]
port 25 nsew default output
rlabel metal2 s 27986 219200 28042 220000 6 cpu_addr_n[3]
port 26 nsew default output
rlabel metal2 s 30010 219200 30066 220000 6 cpu_addr_n[4]
port 27 nsew default output
rlabel metal2 s 32126 219200 32182 220000 6 cpu_addr_n[5]
port 28 nsew default output
rlabel metal2 s 34150 219200 34206 220000 6 cpu_addr_n[6]
port 29 nsew default output
rlabel metal2 s 36266 219200 36322 220000 6 cpu_addr_n[7]
port 30 nsew default output
rlabel metal2 s 38382 219200 38438 220000 6 cpu_addr_n[8]
port 31 nsew default output
rlabel metal2 s 40406 219200 40462 220000 6 cpu_addr_n[9]
port 32 nsew default output
rlabel metal3 s 219200 45704 220000 45824 6 cpu_dtr_e0[0]
port 33 nsew default input
rlabel metal3 s 219200 55904 220000 56024 6 cpu_dtr_e0[10]
port 34 nsew default input
rlabel metal3 s 219200 56856 220000 56976 6 cpu_dtr_e0[11]
port 35 nsew default input
rlabel metal3 s 219200 57944 220000 58064 6 cpu_dtr_e0[12]
port 36 nsew default input
rlabel metal3 s 219200 58896 220000 59016 6 cpu_dtr_e0[13]
port 37 nsew default input
rlabel metal3 s 219200 59848 220000 59968 6 cpu_dtr_e0[14]
port 38 nsew default input
rlabel metal3 s 219200 60936 220000 61056 6 cpu_dtr_e0[15]
port 39 nsew default input
rlabel metal3 s 219200 61888 220000 62008 6 cpu_dtr_e0[16]
port 40 nsew default input
rlabel metal3 s 219200 62976 220000 63096 6 cpu_dtr_e0[17]
port 41 nsew default input
rlabel metal3 s 219200 63928 220000 64048 6 cpu_dtr_e0[18]
port 42 nsew default input
rlabel metal3 s 219200 65016 220000 65136 6 cpu_dtr_e0[19]
port 43 nsew default input
rlabel metal3 s 219200 46792 220000 46912 6 cpu_dtr_e0[1]
port 44 nsew default input
rlabel metal3 s 219200 65968 220000 66088 6 cpu_dtr_e0[20]
port 45 nsew default input
rlabel metal3 s 219200 66920 220000 67040 6 cpu_dtr_e0[21]
port 46 nsew default input
rlabel metal3 s 219200 68008 220000 68128 6 cpu_dtr_e0[22]
port 47 nsew default input
rlabel metal3 s 219200 68960 220000 69080 6 cpu_dtr_e0[23]
port 48 nsew default input
rlabel metal3 s 219200 70048 220000 70168 6 cpu_dtr_e0[24]
port 49 nsew default input
rlabel metal3 s 219200 71000 220000 71120 6 cpu_dtr_e0[25]
port 50 nsew default input
rlabel metal3 s 219200 71952 220000 72072 6 cpu_dtr_e0[26]
port 51 nsew default input
rlabel metal3 s 219200 73040 220000 73160 6 cpu_dtr_e0[27]
port 52 nsew default input
rlabel metal3 s 219200 73992 220000 74112 6 cpu_dtr_e0[28]
port 53 nsew default input
rlabel metal3 s 219200 75080 220000 75200 6 cpu_dtr_e0[29]
port 54 nsew default input
rlabel metal3 s 219200 47744 220000 47864 6 cpu_dtr_e0[2]
port 55 nsew default input
rlabel metal3 s 219200 76032 220000 76152 6 cpu_dtr_e0[30]
port 56 nsew default input
rlabel metal3 s 219200 77120 220000 77240 6 cpu_dtr_e0[31]
port 57 nsew default input
rlabel metal3 s 219200 48832 220000 48952 6 cpu_dtr_e0[3]
port 58 nsew default input
rlabel metal3 s 219200 49784 220000 49904 6 cpu_dtr_e0[4]
port 59 nsew default input
rlabel metal3 s 219200 50872 220000 50992 6 cpu_dtr_e0[5]
port 60 nsew default input
rlabel metal3 s 219200 51824 220000 51944 6 cpu_dtr_e0[6]
port 61 nsew default input
rlabel metal3 s 219200 52776 220000 52896 6 cpu_dtr_e0[7]
port 62 nsew default input
rlabel metal3 s 219200 53864 220000 53984 6 cpu_dtr_e0[8]
port 63 nsew default input
rlabel metal3 s 219200 54816 220000 54936 6 cpu_dtr_e0[9]
port 64 nsew default input
rlabel metal3 s 219200 78072 220000 78192 6 cpu_dtr_e1[0]
port 65 nsew default input
rlabel metal3 s 219200 88136 220000 88256 6 cpu_dtr_e1[10]
port 66 nsew default input
rlabel metal3 s 219200 89224 220000 89344 6 cpu_dtr_e1[11]
port 67 nsew default input
rlabel metal3 s 219200 90176 220000 90296 6 cpu_dtr_e1[12]
port 68 nsew default input
rlabel metal3 s 219200 91128 220000 91248 6 cpu_dtr_e1[13]
port 69 nsew default input
rlabel metal3 s 219200 92216 220000 92336 6 cpu_dtr_e1[14]
port 70 nsew default input
rlabel metal3 s 219200 93168 220000 93288 6 cpu_dtr_e1[15]
port 71 nsew default input
rlabel metal3 s 219200 94256 220000 94376 6 cpu_dtr_e1[16]
port 72 nsew default input
rlabel metal3 s 219200 95208 220000 95328 6 cpu_dtr_e1[17]
port 73 nsew default input
rlabel metal3 s 219200 96296 220000 96416 6 cpu_dtr_e1[18]
port 74 nsew default input
rlabel metal3 s 219200 97248 220000 97368 6 cpu_dtr_e1[19]
port 75 nsew default input
rlabel metal3 s 219200 79024 220000 79144 6 cpu_dtr_e1[1]
port 76 nsew default input
rlabel metal3 s 219200 98200 220000 98320 6 cpu_dtr_e1[20]
port 77 nsew default input
rlabel metal3 s 219200 99288 220000 99408 6 cpu_dtr_e1[21]
port 78 nsew default input
rlabel metal3 s 219200 100240 220000 100360 6 cpu_dtr_e1[22]
port 79 nsew default input
rlabel metal3 s 219200 101328 220000 101448 6 cpu_dtr_e1[23]
port 80 nsew default input
rlabel metal3 s 219200 102280 220000 102400 6 cpu_dtr_e1[24]
port 81 nsew default input
rlabel metal3 s 219200 103368 220000 103488 6 cpu_dtr_e1[25]
port 82 nsew default input
rlabel metal3 s 219200 104320 220000 104440 6 cpu_dtr_e1[26]
port 83 nsew default input
rlabel metal3 s 219200 105272 220000 105392 6 cpu_dtr_e1[27]
port 84 nsew default input
rlabel metal3 s 219200 106360 220000 106480 6 cpu_dtr_e1[28]
port 85 nsew default input
rlabel metal3 s 219200 107312 220000 107432 6 cpu_dtr_e1[29]
port 86 nsew default input
rlabel metal3 s 219200 80112 220000 80232 6 cpu_dtr_e1[2]
port 87 nsew default input
rlabel metal3 s 219200 108400 220000 108520 6 cpu_dtr_e1[30]
port 88 nsew default input
rlabel metal3 s 219200 109352 220000 109472 6 cpu_dtr_e1[31]
port 89 nsew default input
rlabel metal3 s 219200 81064 220000 81184 6 cpu_dtr_e1[3]
port 90 nsew default input
rlabel metal3 s 219200 82152 220000 82272 6 cpu_dtr_e1[4]
port 91 nsew default input
rlabel metal3 s 219200 83104 220000 83224 6 cpu_dtr_e1[5]
port 92 nsew default input
rlabel metal3 s 219200 84192 220000 84312 6 cpu_dtr_e1[6]
port 93 nsew default input
rlabel metal3 s 219200 85144 220000 85264 6 cpu_dtr_e1[7]
port 94 nsew default input
rlabel metal3 s 219200 86096 220000 86216 6 cpu_dtr_e1[8]
port 95 nsew default input
rlabel metal3 s 219200 87184 220000 87304 6 cpu_dtr_e1[9]
port 96 nsew default input
rlabel metal2 s 88154 219200 88210 220000 6 cpu_dtr_n0[0]
port 97 nsew default input
rlabel metal2 s 108854 219200 108910 220000 6 cpu_dtr_n0[10]
port 98 nsew default input
rlabel metal2 s 110970 219200 111026 220000 6 cpu_dtr_n0[11]
port 99 nsew default input
rlabel metal2 s 113086 219200 113142 220000 6 cpu_dtr_n0[12]
port 100 nsew default input
rlabel metal2 s 115110 219200 115166 220000 6 cpu_dtr_n0[13]
port 101 nsew default input
rlabel metal2 s 117226 219200 117282 220000 6 cpu_dtr_n0[14]
port 102 nsew default input
rlabel metal2 s 119250 219200 119306 220000 6 cpu_dtr_n0[15]
port 103 nsew default input
rlabel metal2 s 121366 219200 121422 220000 6 cpu_dtr_n0[16]
port 104 nsew default input
rlabel metal2 s 123390 219200 123446 220000 6 cpu_dtr_n0[17]
port 105 nsew default input
rlabel metal2 s 125506 219200 125562 220000 6 cpu_dtr_n0[18]
port 106 nsew default input
rlabel metal2 s 127530 219200 127586 220000 6 cpu_dtr_n0[19]
port 107 nsew default input
rlabel metal2 s 90178 219200 90234 220000 6 cpu_dtr_n0[1]
port 108 nsew default input
rlabel metal2 s 129646 219200 129702 220000 6 cpu_dtr_n0[20]
port 109 nsew default input
rlabel metal2 s 131762 219200 131818 220000 6 cpu_dtr_n0[21]
port 110 nsew default input
rlabel metal2 s 133786 219200 133842 220000 6 cpu_dtr_n0[22]
port 111 nsew default input
rlabel metal2 s 135902 219200 135958 220000 6 cpu_dtr_n0[23]
port 112 nsew default input
rlabel metal2 s 137926 219200 137982 220000 6 cpu_dtr_n0[24]
port 113 nsew default input
rlabel metal2 s 140042 219200 140098 220000 6 cpu_dtr_n0[25]
port 114 nsew default input
rlabel metal2 s 142066 219200 142122 220000 6 cpu_dtr_n0[26]
port 115 nsew default input
rlabel metal2 s 144182 219200 144238 220000 6 cpu_dtr_n0[27]
port 116 nsew default input
rlabel metal2 s 146206 219200 146262 220000 6 cpu_dtr_n0[28]
port 117 nsew default input
rlabel metal2 s 148322 219200 148378 220000 6 cpu_dtr_n0[29]
port 118 nsew default input
rlabel metal2 s 92294 219200 92350 220000 6 cpu_dtr_n0[2]
port 119 nsew default input
rlabel metal2 s 150438 219200 150494 220000 6 cpu_dtr_n0[30]
port 120 nsew default input
rlabel metal2 s 152462 219200 152518 220000 6 cpu_dtr_n0[31]
port 121 nsew default input
rlabel metal2 s 94410 219200 94466 220000 6 cpu_dtr_n0[3]
port 122 nsew default input
rlabel metal2 s 96434 219200 96490 220000 6 cpu_dtr_n0[4]
port 123 nsew default input
rlabel metal2 s 98550 219200 98606 220000 6 cpu_dtr_n0[5]
port 124 nsew default input
rlabel metal2 s 100574 219200 100630 220000 6 cpu_dtr_n0[6]
port 125 nsew default input
rlabel metal2 s 102690 219200 102746 220000 6 cpu_dtr_n0[7]
port 126 nsew default input
rlabel metal2 s 104714 219200 104770 220000 6 cpu_dtr_n0[8]
port 127 nsew default input
rlabel metal2 s 106830 219200 106886 220000 6 cpu_dtr_n0[9]
port 128 nsew default input
rlabel metal2 s 154578 219200 154634 220000 6 cpu_dtr_n1[0]
port 129 nsew default input
rlabel metal2 s 175278 219200 175334 220000 6 cpu_dtr_n1[10]
port 130 nsew default input
rlabel metal2 s 177394 219200 177450 220000 6 cpu_dtr_n1[11]
port 131 nsew default input
rlabel metal2 s 179418 219200 179474 220000 6 cpu_dtr_n1[12]
port 132 nsew default input
rlabel metal2 s 181534 219200 181590 220000 6 cpu_dtr_n1[13]
port 133 nsew default input
rlabel metal2 s 183558 219200 183614 220000 6 cpu_dtr_n1[14]
port 134 nsew default input
rlabel metal2 s 185674 219200 185730 220000 6 cpu_dtr_n1[15]
port 135 nsew default input
rlabel metal2 s 187790 219200 187846 220000 6 cpu_dtr_n1[16]
port 136 nsew default input
rlabel metal2 s 189814 219200 189870 220000 6 cpu_dtr_n1[17]
port 137 nsew default input
rlabel metal2 s 191930 219200 191986 220000 6 cpu_dtr_n1[18]
port 138 nsew default input
rlabel metal2 s 193954 219200 194010 220000 6 cpu_dtr_n1[19]
port 139 nsew default input
rlabel metal2 s 156602 219200 156658 220000 6 cpu_dtr_n1[1]
port 140 nsew default input
rlabel metal2 s 196070 219200 196126 220000 6 cpu_dtr_n1[20]
port 141 nsew default input
rlabel metal2 s 198094 219200 198150 220000 6 cpu_dtr_n1[21]
port 142 nsew default input
rlabel metal2 s 200210 219200 200266 220000 6 cpu_dtr_n1[22]
port 143 nsew default input
rlabel metal2 s 202234 219200 202290 220000 6 cpu_dtr_n1[23]
port 144 nsew default input
rlabel metal2 s 204350 219200 204406 220000 6 cpu_dtr_n1[24]
port 145 nsew default input
rlabel metal2 s 206466 219200 206522 220000 6 cpu_dtr_n1[25]
port 146 nsew default input
rlabel metal2 s 208490 219200 208546 220000 6 cpu_dtr_n1[26]
port 147 nsew default input
rlabel metal2 s 210606 219200 210662 220000 6 cpu_dtr_n1[27]
port 148 nsew default input
rlabel metal2 s 212630 219200 212686 220000 6 cpu_dtr_n1[28]
port 149 nsew default input
rlabel metal2 s 214746 219200 214802 220000 6 cpu_dtr_n1[29]
port 150 nsew default input
rlabel metal2 s 158718 219200 158774 220000 6 cpu_dtr_n1[2]
port 151 nsew default input
rlabel metal2 s 216770 219200 216826 220000 6 cpu_dtr_n1[30]
port 152 nsew default input
rlabel metal2 s 218886 219200 218942 220000 6 cpu_dtr_n1[31]
port 153 nsew default input
rlabel metal2 s 160742 219200 160798 220000 6 cpu_dtr_n1[3]
port 154 nsew default input
rlabel metal2 s 162858 219200 162914 220000 6 cpu_dtr_n1[4]
port 155 nsew default input
rlabel metal2 s 164882 219200 164938 220000 6 cpu_dtr_n1[5]
port 156 nsew default input
rlabel metal2 s 166998 219200 167054 220000 6 cpu_dtr_n1[6]
port 157 nsew default input
rlabel metal2 s 169114 219200 169170 220000 6 cpu_dtr_n1[7]
port 158 nsew default input
rlabel metal2 s 171138 219200 171194 220000 6 cpu_dtr_n1[8]
port 159 nsew default input
rlabel metal2 s 173254 219200 173310 220000 6 cpu_dtr_n1[9]
port 160 nsew default input
rlabel metal3 s 219200 29656 220000 29776 6 cpu_dtw_e[0]
port 161 nsew default output
rlabel metal3 s 219200 39720 220000 39840 6 cpu_dtw_e[10]
port 162 nsew default output
rlabel metal3 s 219200 40672 220000 40792 6 cpu_dtw_e[11]
port 163 nsew default output
rlabel metal3 s 219200 41760 220000 41880 6 cpu_dtw_e[12]
port 164 nsew default output
rlabel metal3 s 219200 42712 220000 42832 6 cpu_dtw_e[13]
port 165 nsew default output
rlabel metal3 s 219200 43800 220000 43920 6 cpu_dtw_e[14]
port 166 nsew default output
rlabel metal3 s 219200 44752 220000 44872 6 cpu_dtw_e[15]
port 167 nsew default output
rlabel metal3 s 219200 30608 220000 30728 6 cpu_dtw_e[1]
port 168 nsew default output
rlabel metal3 s 219200 31696 220000 31816 6 cpu_dtw_e[2]
port 169 nsew default output
rlabel metal3 s 219200 32648 220000 32768 6 cpu_dtw_e[3]
port 170 nsew default output
rlabel metal3 s 219200 33600 220000 33720 6 cpu_dtw_e[4]
port 171 nsew default output
rlabel metal3 s 219200 34688 220000 34808 6 cpu_dtw_e[5]
port 172 nsew default output
rlabel metal3 s 219200 35640 220000 35760 6 cpu_dtw_e[6]
port 173 nsew default output
rlabel metal3 s 219200 36728 220000 36848 6 cpu_dtw_e[7]
port 174 nsew default output
rlabel metal3 s 219200 37680 220000 37800 6 cpu_dtw_e[8]
port 175 nsew default output
rlabel metal3 s 219200 38768 220000 38888 6 cpu_dtw_e[9]
port 176 nsew default output
rlabel metal2 s 54942 219200 54998 220000 6 cpu_dtw_n[0]
port 177 nsew default output
rlabel metal2 s 75734 219200 75790 220000 6 cpu_dtw_n[10]
port 178 nsew default output
rlabel metal2 s 77758 219200 77814 220000 6 cpu_dtw_n[11]
port 179 nsew default output
rlabel metal2 s 79874 219200 79930 220000 6 cpu_dtw_n[12]
port 180 nsew default output
rlabel metal2 s 81898 219200 81954 220000 6 cpu_dtw_n[13]
port 181 nsew default output
rlabel metal2 s 84014 219200 84070 220000 6 cpu_dtw_n[14]
port 182 nsew default output
rlabel metal2 s 86038 219200 86094 220000 6 cpu_dtw_n[15]
port 183 nsew default output
rlabel metal2 s 57058 219200 57114 220000 6 cpu_dtw_n[1]
port 184 nsew default output
rlabel metal2 s 59082 219200 59138 220000 6 cpu_dtw_n[2]
port 185 nsew default output
rlabel metal2 s 61198 219200 61254 220000 6 cpu_dtw_n[3]
port 186 nsew default output
rlabel metal2 s 63222 219200 63278 220000 6 cpu_dtw_n[4]
port 187 nsew default output
rlabel metal2 s 65338 219200 65394 220000 6 cpu_dtw_n[5]
port 188 nsew default output
rlabel metal2 s 67362 219200 67418 220000 6 cpu_dtw_n[6]
port 189 nsew default output
rlabel metal2 s 69478 219200 69534 220000 6 cpu_dtw_n[7]
port 190 nsew default output
rlabel metal2 s 71502 219200 71558 220000 6 cpu_dtw_n[8]
port 191 nsew default output
rlabel metal2 s 73618 219200 73674 220000 6 cpu_dtw_n[9]
port 192 nsew default output
rlabel metal3 s 219200 3408 220000 3528 6 cpu_mask_e[0]
port 193 nsew default output
rlabel metal3 s 219200 4360 220000 4480 6 cpu_mask_e[1]
port 194 nsew default output
rlabel metal3 s 219200 5448 220000 5568 6 cpu_mask_e[2]
port 195 nsew default output
rlabel metal3 s 219200 6400 220000 6520 6 cpu_mask_e[3]
port 196 nsew default output
rlabel metal3 s 219200 7352 220000 7472 6 cpu_mask_e[4]
port 197 nsew default output
rlabel metal3 s 219200 8440 220000 8560 6 cpu_mask_e[5]
port 198 nsew default output
rlabel metal3 s 219200 9392 220000 9512 6 cpu_mask_e[6]
port 199 nsew default output
rlabel metal3 s 219200 10480 220000 10600 6 cpu_mask_e[7]
port 200 nsew default output
rlabel metal2 s 1030 219200 1086 220000 6 cpu_mask_n[0]
port 201 nsew default output
rlabel metal2 s 3054 219200 3110 220000 6 cpu_mask_n[1]
port 202 nsew default output
rlabel metal2 s 5170 219200 5226 220000 6 cpu_mask_n[2]
port 203 nsew default output
rlabel metal2 s 7194 219200 7250 220000 6 cpu_mask_n[3]
port 204 nsew default output
rlabel metal2 s 9310 219200 9366 220000 6 cpu_mask_n[4]
port 205 nsew default output
rlabel metal2 s 11334 219200 11390 220000 6 cpu_mask_n[5]
port 206 nsew default output
rlabel metal2 s 13450 219200 13506 220000 6 cpu_mask_n[6]
port 207 nsew default output
rlabel metal2 s 15474 219200 15530 220000 6 cpu_mask_n[7]
port 208 nsew default output
rlabel metal3 s 219200 11432 220000 11552 6 cpu_wen_e[0]
port 209 nsew default output
rlabel metal3 s 219200 12520 220000 12640 6 cpu_wen_e[1]
port 210 nsew default output
rlabel metal2 s 17590 219200 17646 220000 6 cpu_wen_n[0]
port 211 nsew default output
rlabel metal2 s 19706 219200 19762 220000 6 cpu_wen_n[1]
port 212 nsew default output
rlabel metal3 s 0 960 800 1080 6 io_in[0]
port 213 nsew default input
rlabel metal3 s 0 58760 800 58880 6 io_in[10]
port 214 nsew default input
rlabel metal3 s 0 64608 800 64728 6 io_in[11]
port 215 nsew default input
rlabel metal3 s 0 70320 800 70440 6 io_in[12]
port 216 nsew default input
rlabel metal3 s 0 76168 800 76288 6 io_in[13]
port 217 nsew default input
rlabel metal3 s 0 82016 800 82136 6 io_in[14]
port 218 nsew default input
rlabel metal3 s 0 87728 800 87848 6 io_in[15]
port 219 nsew default input
rlabel metal3 s 0 93576 800 93696 6 io_in[16]
port 220 nsew default input
rlabel metal3 s 0 99288 800 99408 6 io_in[17]
port 221 nsew default input
rlabel metal3 s 0 105136 800 105256 6 io_in[18]
port 222 nsew default input
rlabel metal3 s 0 110984 800 111104 6 io_in[19]
port 223 nsew default input
rlabel metal3 s 0 6672 800 6792 6 io_in[1]
port 224 nsew default input
rlabel metal3 s 0 116696 800 116816 6 io_in[20]
port 225 nsew default input
rlabel metal3 s 0 122544 800 122664 6 io_in[21]
port 226 nsew default input
rlabel metal3 s 0 128256 800 128376 6 io_in[22]
port 227 nsew default input
rlabel metal3 s 0 134104 800 134224 6 io_in[23]
port 228 nsew default input
rlabel metal3 s 0 139816 800 139936 6 io_in[24]
port 229 nsew default input
rlabel metal3 s 0 145664 800 145784 6 io_in[25]
port 230 nsew default input
rlabel metal3 s 0 151512 800 151632 6 io_in[26]
port 231 nsew default input
rlabel metal3 s 0 157224 800 157344 6 io_in[27]
port 232 nsew default input
rlabel metal3 s 0 163072 800 163192 6 io_in[28]
port 233 nsew default input
rlabel metal3 s 0 168784 800 168904 6 io_in[29]
port 234 nsew default input
rlabel metal3 s 0 12520 800 12640 6 io_in[2]
port 235 nsew default input
rlabel metal3 s 0 174632 800 174752 6 io_in[30]
port 236 nsew default input
rlabel metal3 s 0 180344 800 180464 6 io_in[31]
port 237 nsew default input
rlabel metal3 s 0 186192 800 186312 6 io_in[32]
port 238 nsew default input
rlabel metal3 s 0 192040 800 192160 6 io_in[33]
port 239 nsew default input
rlabel metal3 s 0 197752 800 197872 6 io_in[34]
port 240 nsew default input
rlabel metal3 s 0 203600 800 203720 6 io_in[35]
port 241 nsew default input
rlabel metal3 s 0 209312 800 209432 6 io_in[36]
port 242 nsew default input
rlabel metal3 s 0 215160 800 215280 6 io_in[37]
port 243 nsew default input
rlabel metal3 s 0 18232 800 18352 6 io_in[3]
port 244 nsew default input
rlabel metal3 s 0 24080 800 24200 6 io_in[4]
port 245 nsew default input
rlabel metal3 s 0 29792 800 29912 6 io_in[5]
port 246 nsew default input
rlabel metal3 s 0 35640 800 35760 6 io_in[6]
port 247 nsew default input
rlabel metal3 s 0 41488 800 41608 6 io_in[7]
port 248 nsew default input
rlabel metal3 s 0 47200 800 47320 6 io_in[8]
port 249 nsew default input
rlabel metal3 s 0 53048 800 53168 6 io_in[9]
port 250 nsew default input
rlabel metal3 s 0 2864 800 2984 6 io_oeb[0]
port 251 nsew default output
rlabel metal3 s 0 60664 800 60784 6 io_oeb[10]
port 252 nsew default output
rlabel metal3 s 0 66512 800 66632 6 io_oeb[11]
port 253 nsew default output
rlabel metal3 s 0 72360 800 72480 6 io_oeb[12]
port 254 nsew default output
rlabel metal3 s 0 78072 800 78192 6 io_oeb[13]
port 255 nsew default output
rlabel metal3 s 0 83920 800 84040 6 io_oeb[14]
port 256 nsew default output
rlabel metal3 s 0 89632 800 89752 6 io_oeb[15]
port 257 nsew default output
rlabel metal3 s 0 95480 800 95600 6 io_oeb[16]
port 258 nsew default output
rlabel metal3 s 0 101328 800 101448 6 io_oeb[17]
port 259 nsew default output
rlabel metal3 s 0 107040 800 107160 6 io_oeb[18]
port 260 nsew default output
rlabel metal3 s 0 112888 800 113008 6 io_oeb[19]
port 261 nsew default output
rlabel metal3 s 0 8576 800 8696 6 io_oeb[1]
port 262 nsew default output
rlabel metal3 s 0 118600 800 118720 6 io_oeb[20]
port 263 nsew default output
rlabel metal3 s 0 124448 800 124568 6 io_oeb[21]
port 264 nsew default output
rlabel metal3 s 0 130160 800 130280 6 io_oeb[22]
port 265 nsew default output
rlabel metal3 s 0 136008 800 136128 6 io_oeb[23]
port 266 nsew default output
rlabel metal3 s 0 141856 800 141976 6 io_oeb[24]
port 267 nsew default output
rlabel metal3 s 0 147568 800 147688 6 io_oeb[25]
port 268 nsew default output
rlabel metal3 s 0 153416 800 153536 6 io_oeb[26]
port 269 nsew default output
rlabel metal3 s 0 159128 800 159248 6 io_oeb[27]
port 270 nsew default output
rlabel metal3 s 0 164976 800 165096 6 io_oeb[28]
port 271 nsew default output
rlabel metal3 s 0 170688 800 170808 6 io_oeb[29]
port 272 nsew default output
rlabel metal3 s 0 14424 800 14544 6 io_oeb[2]
port 273 nsew default output
rlabel metal3 s 0 176536 800 176656 6 io_oeb[30]
port 274 nsew default output
rlabel metal3 s 0 182384 800 182504 6 io_oeb[31]
port 275 nsew default output
rlabel metal3 s 0 188096 800 188216 6 io_oeb[32]
port 276 nsew default output
rlabel metal3 s 0 193944 800 194064 6 io_oeb[33]
port 277 nsew default output
rlabel metal3 s 0 199656 800 199776 6 io_oeb[34]
port 278 nsew default output
rlabel metal3 s 0 205504 800 205624 6 io_oeb[35]
port 279 nsew default output
rlabel metal3 s 0 211352 800 211472 6 io_oeb[36]
port 280 nsew default output
rlabel metal3 s 0 217064 800 217184 6 io_oeb[37]
port 281 nsew default output
rlabel metal3 s 0 20136 800 20256 6 io_oeb[3]
port 282 nsew default output
rlabel metal3 s 0 25984 800 26104 6 io_oeb[4]
port 283 nsew default output
rlabel metal3 s 0 31832 800 31952 6 io_oeb[5]
port 284 nsew default output
rlabel metal3 s 0 37544 800 37664 6 io_oeb[6]
port 285 nsew default output
rlabel metal3 s 0 43392 800 43512 6 io_oeb[7]
port 286 nsew default output
rlabel metal3 s 0 49104 800 49224 6 io_oeb[8]
port 287 nsew default output
rlabel metal3 s 0 54952 800 55072 6 io_oeb[9]
port 288 nsew default output
rlabel metal3 s 0 4768 800 4888 6 io_out[0]
port 289 nsew default output
rlabel metal3 s 0 62704 800 62824 6 io_out[10]
port 290 nsew default output
rlabel metal3 s 0 68416 800 68536 6 io_out[11]
port 291 nsew default output
rlabel metal3 s 0 74264 800 74384 6 io_out[12]
port 292 nsew default output
rlabel metal3 s 0 79976 800 80096 6 io_out[13]
port 293 nsew default output
rlabel metal3 s 0 85824 800 85944 6 io_out[14]
port 294 nsew default output
rlabel metal3 s 0 91672 800 91792 6 io_out[15]
port 295 nsew default output
rlabel metal3 s 0 97384 800 97504 6 io_out[16]
port 296 nsew default output
rlabel metal3 s 0 103232 800 103352 6 io_out[17]
port 297 nsew default output
rlabel metal3 s 0 108944 800 109064 6 io_out[18]
port 298 nsew default output
rlabel metal3 s 0 114792 800 114912 6 io_out[19]
port 299 nsew default output
rlabel metal3 s 0 10480 800 10600 6 io_out[1]
port 300 nsew default output
rlabel metal3 s 0 120504 800 120624 6 io_out[20]
port 301 nsew default output
rlabel metal3 s 0 126352 800 126472 6 io_out[21]
port 302 nsew default output
rlabel metal3 s 0 132200 800 132320 6 io_out[22]
port 303 nsew default output
rlabel metal3 s 0 137912 800 138032 6 io_out[23]
port 304 nsew default output
rlabel metal3 s 0 143760 800 143880 6 io_out[24]
port 305 nsew default output
rlabel metal3 s 0 149472 800 149592 6 io_out[25]
port 306 nsew default output
rlabel metal3 s 0 155320 800 155440 6 io_out[26]
port 307 nsew default output
rlabel metal3 s 0 161168 800 161288 6 io_out[27]
port 308 nsew default output
rlabel metal3 s 0 166880 800 167000 6 io_out[28]
port 309 nsew default output
rlabel metal3 s 0 172728 800 172848 6 io_out[29]
port 310 nsew default output
rlabel metal3 s 0 16328 800 16448 6 io_out[2]
port 311 nsew default output
rlabel metal3 s 0 178440 800 178560 6 io_out[30]
port 312 nsew default output
rlabel metal3 s 0 184288 800 184408 6 io_out[31]
port 313 nsew default output
rlabel metal3 s 0 190000 800 190120 6 io_out[32]
port 314 nsew default output
rlabel metal3 s 0 195848 800 195968 6 io_out[33]
port 315 nsew default output
rlabel metal3 s 0 201696 800 201816 6 io_out[34]
port 316 nsew default output
rlabel metal3 s 0 207408 800 207528 6 io_out[35]
port 317 nsew default output
rlabel metal3 s 0 213256 800 213376 6 io_out[36]
port 318 nsew default output
rlabel metal3 s 0 218968 800 219088 6 io_out[37]
port 319 nsew default output
rlabel metal3 s 0 22176 800 22296 6 io_out[3]
port 320 nsew default output
rlabel metal3 s 0 27888 800 28008 6 io_out[4]
port 321 nsew default output
rlabel metal3 s 0 33736 800 33856 6 io_out[5]
port 322 nsew default output
rlabel metal3 s 0 39448 800 39568 6 io_out[6]
port 323 nsew default output
rlabel metal3 s 0 45296 800 45416 6 io_out[7]
port 324 nsew default output
rlabel metal3 s 0 51144 800 51264 6 io_out[8]
port 325 nsew default output
rlabel metal3 s 0 56856 800 56976 6 io_out[9]
port 326 nsew default output
rlabel metal2 s 207202 0 207258 800 6 la_data_in[0]
port 327 nsew default input
rlabel metal2 s 213090 0 213146 800 6 la_data_in[1]
port 328 nsew default input
rlabel metal2 s 209226 0 209282 800 6 la_data_out[0]
port 329 nsew default output
rlabel metal2 s 215022 0 215078 800 6 la_data_out[1]
port 330 nsew default output
rlabel metal2 s 218886 0 218942 800 6 la_data_out[2]
port 331 nsew default output
rlabel metal2 s 211158 0 211214 800 6 la_oen[0]
port 332 nsew default input
rlabel metal2 s 216954 0 217010 800 6 la_oen[1]
port 333 nsew default input
rlabel metal3 s 219200 1368 220000 1488 6 one
port 334 nsew default output
rlabel metal3 s 219200 2320 220000 2440 6 ram_ce
port 335 nsew default output
rlabel metal3 s 219200 110440 220000 110560 6 sr0_ce
port 336 nsew default output
rlabel metal3 s 219200 111392 220000 111512 6 sr0_dtr[0]
port 337 nsew default input
rlabel metal3 s 219200 121456 220000 121576 6 sr0_dtr[10]
port 338 nsew default input
rlabel metal3 s 219200 122544 220000 122664 6 sr0_dtr[11]
port 339 nsew default input
rlabel metal3 s 219200 123496 220000 123616 6 sr0_dtr[12]
port 340 nsew default input
rlabel metal3 s 219200 124448 220000 124568 6 sr0_dtr[13]
port 341 nsew default input
rlabel metal3 s 219200 125536 220000 125656 6 sr0_dtr[14]
port 342 nsew default input
rlabel metal3 s 219200 126488 220000 126608 6 sr0_dtr[15]
port 343 nsew default input
rlabel metal3 s 219200 127576 220000 127696 6 sr0_dtr[16]
port 344 nsew default input
rlabel metal3 s 219200 128528 220000 128648 6 sr0_dtr[17]
port 345 nsew default input
rlabel metal3 s 219200 129616 220000 129736 6 sr0_dtr[18]
port 346 nsew default input
rlabel metal3 s 219200 130568 220000 130688 6 sr0_dtr[19]
port 347 nsew default input
rlabel metal3 s 219200 112344 220000 112464 6 sr0_dtr[1]
port 348 nsew default input
rlabel metal3 s 219200 131520 220000 131640 6 sr0_dtr[20]
port 349 nsew default input
rlabel metal3 s 219200 132608 220000 132728 6 sr0_dtr[21]
port 350 nsew default input
rlabel metal3 s 219200 133560 220000 133680 6 sr0_dtr[22]
port 351 nsew default input
rlabel metal3 s 219200 134648 220000 134768 6 sr0_dtr[23]
port 352 nsew default input
rlabel metal3 s 219200 135600 220000 135720 6 sr0_dtr[24]
port 353 nsew default input
rlabel metal3 s 219200 136552 220000 136672 6 sr0_dtr[25]
port 354 nsew default input
rlabel metal3 s 219200 137640 220000 137760 6 sr0_dtr[26]
port 355 nsew default input
rlabel metal3 s 219200 138592 220000 138712 6 sr0_dtr[27]
port 356 nsew default input
rlabel metal3 s 219200 139680 220000 139800 6 sr0_dtr[28]
port 357 nsew default input
rlabel metal3 s 219200 140632 220000 140752 6 sr0_dtr[29]
port 358 nsew default input
rlabel metal3 s 219200 113432 220000 113552 6 sr0_dtr[2]
port 359 nsew default input
rlabel metal3 s 219200 141720 220000 141840 6 sr0_dtr[30]
port 360 nsew default input
rlabel metal3 s 219200 142672 220000 142792 6 sr0_dtr[31]
port 361 nsew default input
rlabel metal3 s 219200 114384 220000 114504 6 sr0_dtr[3]
port 362 nsew default input
rlabel metal3 s 219200 115472 220000 115592 6 sr0_dtr[4]
port 363 nsew default input
rlabel metal3 s 219200 116424 220000 116544 6 sr0_dtr[5]
port 364 nsew default input
rlabel metal3 s 219200 117376 220000 117496 6 sr0_dtr[6]
port 365 nsew default input
rlabel metal3 s 219200 118464 220000 118584 6 sr0_dtr[7]
port 366 nsew default input
rlabel metal3 s 219200 119416 220000 119536 6 sr0_dtr[8]
port 367 nsew default input
rlabel metal3 s 219200 120504 220000 120624 6 sr0_dtr[9]
port 368 nsew default input
rlabel metal3 s 219200 143624 220000 143744 6 sr1_ce
port 369 nsew default output
rlabel metal3 s 219200 144712 220000 144832 6 sr1_dtr[0]
port 370 nsew default input
rlabel metal3 s 219200 154776 220000 154896 6 sr1_dtr[10]
port 371 nsew default input
rlabel metal3 s 219200 155728 220000 155848 6 sr1_dtr[11]
port 372 nsew default input
rlabel metal3 s 219200 156816 220000 156936 6 sr1_dtr[12]
port 373 nsew default input
rlabel metal3 s 219200 157768 220000 157888 6 sr1_dtr[13]
port 374 nsew default input
rlabel metal3 s 219200 158856 220000 158976 6 sr1_dtr[14]
port 375 nsew default input
rlabel metal3 s 219200 159808 220000 159928 6 sr1_dtr[15]
port 376 nsew default input
rlabel metal3 s 219200 160896 220000 161016 6 sr1_dtr[16]
port 377 nsew default input
rlabel metal3 s 219200 161848 220000 161968 6 sr1_dtr[17]
port 378 nsew default input
rlabel metal3 s 219200 162800 220000 162920 6 sr1_dtr[18]
port 379 nsew default input
rlabel metal3 s 219200 163888 220000 164008 6 sr1_dtr[19]
port 380 nsew default input
rlabel metal3 s 219200 145664 220000 145784 6 sr1_dtr[1]
port 381 nsew default input
rlabel metal3 s 219200 164840 220000 164960 6 sr1_dtr[20]
port 382 nsew default input
rlabel metal3 s 219200 165928 220000 166048 6 sr1_dtr[21]
port 383 nsew default input
rlabel metal3 s 219200 166880 220000 167000 6 sr1_dtr[22]
port 384 nsew default input
rlabel metal3 s 219200 167968 220000 168088 6 sr1_dtr[23]
port 385 nsew default input
rlabel metal3 s 219200 168920 220000 169040 6 sr1_dtr[24]
port 386 nsew default input
rlabel metal3 s 219200 169872 220000 169992 6 sr1_dtr[25]
port 387 nsew default input
rlabel metal3 s 219200 170960 220000 171080 6 sr1_dtr[26]
port 388 nsew default input
rlabel metal3 s 219200 171912 220000 172032 6 sr1_dtr[27]
port 389 nsew default input
rlabel metal3 s 219200 173000 220000 173120 6 sr1_dtr[28]
port 390 nsew default input
rlabel metal3 s 219200 173952 220000 174072 6 sr1_dtr[29]
port 391 nsew default input
rlabel metal3 s 219200 146752 220000 146872 6 sr1_dtr[2]
port 392 nsew default input
rlabel metal3 s 219200 175040 220000 175160 6 sr1_dtr[30]
port 393 nsew default input
rlabel metal3 s 219200 175992 220000 176112 6 sr1_dtr[31]
port 394 nsew default input
rlabel metal3 s 219200 147704 220000 147824 6 sr1_dtr[3]
port 395 nsew default input
rlabel metal3 s 219200 148792 220000 148912 6 sr1_dtr[4]
port 396 nsew default input
rlabel metal3 s 219200 149744 220000 149864 6 sr1_dtr[5]
port 397 nsew default input
rlabel metal3 s 219200 150696 220000 150816 6 sr1_dtr[6]
port 398 nsew default input
rlabel metal3 s 219200 151784 220000 151904 6 sr1_dtr[7]
port 399 nsew default input
rlabel metal3 s 219200 152736 220000 152856 6 sr1_dtr[8]
port 400 nsew default input
rlabel metal3 s 219200 153824 220000 153944 6 sr1_dtr[9]
port 401 nsew default input
rlabel metal3 s 219200 178032 220000 178152 6 srx_addr[0]
port 402 nsew default output
rlabel metal3 s 219200 180072 220000 180192 6 srx_addr[1]
port 403 nsew default output
rlabel metal3 s 219200 181976 220000 182096 6 srx_addr[2]
port 404 nsew default output
rlabel metal3 s 219200 184016 220000 184136 6 srx_addr[3]
port 405 nsew default output
rlabel metal3 s 219200 186056 220000 186176 6 srx_addr[4]
port 406 nsew default output
rlabel metal3 s 219200 188096 220000 188216 6 srx_addr[5]
port 407 nsew default output
rlabel metal3 s 219200 190136 220000 190256 6 srx_addr[6]
port 408 nsew default output
rlabel metal3 s 219200 192176 220000 192296 6 srx_addr[7]
port 409 nsew default output
rlabel metal3 s 219200 194216 220000 194336 6 srx_addr[8]
port 410 nsew default output
rlabel metal3 s 219200 196120 220000 196240 6 srx_addr[9]
port 411 nsew default output
rlabel metal3 s 219200 178984 220000 179104 6 srx_dtw[0]
port 412 nsew default output
rlabel metal3 s 219200 198160 220000 198280 6 srx_dtw[10]
port 413 nsew default output
rlabel metal3 s 219200 199248 220000 199368 6 srx_dtw[11]
port 414 nsew default output
rlabel metal3 s 219200 200200 220000 200320 6 srx_dtw[12]
port 415 nsew default output
rlabel metal3 s 219200 201152 220000 201272 6 srx_dtw[13]
port 416 nsew default output
rlabel metal3 s 219200 202240 220000 202360 6 srx_dtw[14]
port 417 nsew default output
rlabel metal3 s 219200 203192 220000 203312 6 srx_dtw[15]
port 418 nsew default output
rlabel metal3 s 219200 204280 220000 204400 6 srx_dtw[16]
port 419 nsew default output
rlabel metal3 s 219200 205232 220000 205352 6 srx_dtw[17]
port 420 nsew default output
rlabel metal3 s 219200 206320 220000 206440 6 srx_dtw[18]
port 421 nsew default output
rlabel metal3 s 219200 207272 220000 207392 6 srx_dtw[19]
port 422 nsew default output
rlabel metal3 s 219200 181024 220000 181144 6 srx_dtw[1]
port 423 nsew default output
rlabel metal3 s 219200 208224 220000 208344 6 srx_dtw[20]
port 424 nsew default output
rlabel metal3 s 219200 209312 220000 209432 6 srx_dtw[21]
port 425 nsew default output
rlabel metal3 s 219200 210264 220000 210384 6 srx_dtw[22]
port 426 nsew default output
rlabel metal3 s 219200 211352 220000 211472 6 srx_dtw[23]
port 427 nsew default output
rlabel metal3 s 219200 212304 220000 212424 6 srx_dtw[24]
port 428 nsew default output
rlabel metal3 s 219200 213392 220000 213512 6 srx_dtw[25]
port 429 nsew default output
rlabel metal3 s 219200 214344 220000 214464 6 srx_dtw[26]
port 430 nsew default output
rlabel metal3 s 219200 215296 220000 215416 6 srx_dtw[27]
port 431 nsew default output
rlabel metal3 s 219200 216384 220000 216504 6 srx_dtw[28]
port 432 nsew default output
rlabel metal3 s 219200 217336 220000 217456 6 srx_dtw[29]
port 433 nsew default output
rlabel metal3 s 219200 183064 220000 183184 6 srx_dtw[2]
port 434 nsew default output
rlabel metal3 s 219200 218424 220000 218544 6 srx_dtw[30]
port 435 nsew default output
rlabel metal3 s 219200 219376 220000 219496 6 srx_dtw[31]
port 436 nsew default output
rlabel metal3 s 219200 185104 220000 185224 6 srx_dtw[3]
port 437 nsew default output
rlabel metal3 s 219200 187144 220000 187264 6 srx_dtw[4]
port 438 nsew default output
rlabel metal3 s 219200 189048 220000 189168 6 srx_dtw[5]
port 439 nsew default output
rlabel metal3 s 219200 191088 220000 191208 6 srx_dtw[6]
port 440 nsew default output
rlabel metal3 s 219200 193128 220000 193248 6 srx_dtw[7]
port 441 nsew default output
rlabel metal3 s 219200 195168 220000 195288 6 srx_dtw[8]
port 442 nsew default output
rlabel metal3 s 219200 197208 220000 197328 6 srx_dtw[9]
port 443 nsew default output
rlabel metal3 s 219200 176944 220000 177064 6 srx_we
port 444 nsew default output
rlabel metal2 s 938 0 994 800 6 wb_clk_i
port 445 nsew default input
rlabel metal2 s 2870 0 2926 800 6 wb_rst_i
port 446 nsew default input
rlabel metal2 s 4802 0 4858 800 6 wbs_ack_o
port 447 nsew default output
rlabel metal2 s 12530 0 12586 800 6 wbs_adr_i[0]
port 448 nsew default input
rlabel metal2 s 78770 0 78826 800 6 wbs_adr_i[10]
port 449 nsew default input
rlabel metal2 s 84566 0 84622 800 6 wbs_adr_i[11]
port 450 nsew default input
rlabel metal2 s 90454 0 90510 800 6 wbs_adr_i[12]
port 451 nsew default input
rlabel metal2 s 96250 0 96306 800 6 wbs_adr_i[13]
port 452 nsew default input
rlabel metal2 s 102138 0 102194 800 6 wbs_adr_i[14]
port 453 nsew default input
rlabel metal2 s 107934 0 107990 800 6 wbs_adr_i[15]
port 454 nsew default input
rlabel metal2 s 113822 0 113878 800 6 wbs_adr_i[16]
port 455 nsew default input
rlabel metal2 s 119618 0 119674 800 6 wbs_adr_i[17]
port 456 nsew default input
rlabel metal2 s 125506 0 125562 800 6 wbs_adr_i[18]
port 457 nsew default input
rlabel metal2 s 131302 0 131358 800 6 wbs_adr_i[19]
port 458 nsew default input
rlabel metal2 s 20350 0 20406 800 6 wbs_adr_i[1]
port 459 nsew default input
rlabel metal2 s 137190 0 137246 800 6 wbs_adr_i[20]
port 460 nsew default input
rlabel metal2 s 142986 0 143042 800 6 wbs_adr_i[21]
port 461 nsew default input
rlabel metal2 s 148874 0 148930 800 6 wbs_adr_i[22]
port 462 nsew default input
rlabel metal2 s 154670 0 154726 800 6 wbs_adr_i[23]
port 463 nsew default input
rlabel metal2 s 160558 0 160614 800 6 wbs_adr_i[24]
port 464 nsew default input
rlabel metal2 s 166354 0 166410 800 6 wbs_adr_i[25]
port 465 nsew default input
rlabel metal2 s 172242 0 172298 800 6 wbs_adr_i[26]
port 466 nsew default input
rlabel metal2 s 178038 0 178094 800 6 wbs_adr_i[27]
port 467 nsew default input
rlabel metal2 s 183834 0 183890 800 6 wbs_adr_i[28]
port 468 nsew default input
rlabel metal2 s 189722 0 189778 800 6 wbs_adr_i[29]
port 469 nsew default input
rlabel metal2 s 28170 0 28226 800 6 wbs_adr_i[2]
port 470 nsew default input
rlabel metal2 s 195518 0 195574 800 6 wbs_adr_i[30]
port 471 nsew default input
rlabel metal2 s 201406 0 201462 800 6 wbs_adr_i[31]
port 472 nsew default input
rlabel metal2 s 35898 0 35954 800 6 wbs_adr_i[3]
port 473 nsew default input
rlabel metal2 s 43718 0 43774 800 6 wbs_adr_i[4]
port 474 nsew default input
rlabel metal2 s 49514 0 49570 800 6 wbs_adr_i[5]
port 475 nsew default input
rlabel metal2 s 55402 0 55458 800 6 wbs_adr_i[6]
port 476 nsew default input
rlabel metal2 s 61198 0 61254 800 6 wbs_adr_i[7]
port 477 nsew default input
rlabel metal2 s 67086 0 67142 800 6 wbs_adr_i[8]
port 478 nsew default input
rlabel metal2 s 72882 0 72938 800 6 wbs_adr_i[9]
port 479 nsew default input
rlabel metal2 s 6734 0 6790 800 6 wbs_cyc_i
port 480 nsew default input
rlabel metal2 s 14554 0 14610 800 6 wbs_dat_i[0]
port 481 nsew default input
rlabel metal2 s 80702 0 80758 800 6 wbs_dat_i[10]
port 482 nsew default input
rlabel metal2 s 86590 0 86646 800 6 wbs_dat_i[11]
port 483 nsew default input
rlabel metal2 s 92386 0 92442 800 6 wbs_dat_i[12]
port 484 nsew default input
rlabel metal2 s 98182 0 98238 800 6 wbs_dat_i[13]
port 485 nsew default input
rlabel metal2 s 104070 0 104126 800 6 wbs_dat_i[14]
port 486 nsew default input
rlabel metal2 s 109866 0 109922 800 6 wbs_dat_i[15]
port 487 nsew default input
rlabel metal2 s 115754 0 115810 800 6 wbs_dat_i[16]
port 488 nsew default input
rlabel metal2 s 121550 0 121606 800 6 wbs_dat_i[17]
port 489 nsew default input
rlabel metal2 s 127438 0 127494 800 6 wbs_dat_i[18]
port 490 nsew default input
rlabel metal2 s 133234 0 133290 800 6 wbs_dat_i[19]
port 491 nsew default input
rlabel metal2 s 22282 0 22338 800 6 wbs_dat_i[1]
port 492 nsew default input
rlabel metal2 s 139122 0 139178 800 6 wbs_dat_i[20]
port 493 nsew default input
rlabel metal2 s 144918 0 144974 800 6 wbs_dat_i[21]
port 494 nsew default input
rlabel metal2 s 150806 0 150862 800 6 wbs_dat_i[22]
port 495 nsew default input
rlabel metal2 s 156602 0 156658 800 6 wbs_dat_i[23]
port 496 nsew default input
rlabel metal2 s 162490 0 162546 800 6 wbs_dat_i[24]
port 497 nsew default input
rlabel metal2 s 168286 0 168342 800 6 wbs_dat_i[25]
port 498 nsew default input
rlabel metal2 s 174174 0 174230 800 6 wbs_dat_i[26]
port 499 nsew default input
rlabel metal2 s 179970 0 180026 800 6 wbs_dat_i[27]
port 500 nsew default input
rlabel metal2 s 185858 0 185914 800 6 wbs_dat_i[28]
port 501 nsew default input
rlabel metal2 s 191654 0 191710 800 6 wbs_dat_i[29]
port 502 nsew default input
rlabel metal2 s 30102 0 30158 800 6 wbs_dat_i[2]
port 503 nsew default input
rlabel metal2 s 197542 0 197598 800 6 wbs_dat_i[30]
port 504 nsew default input
rlabel metal2 s 203338 0 203394 800 6 wbs_dat_i[31]
port 505 nsew default input
rlabel metal2 s 37922 0 37978 800 6 wbs_dat_i[3]
port 506 nsew default input
rlabel metal2 s 45650 0 45706 800 6 wbs_dat_i[4]
port 507 nsew default input
rlabel metal2 s 51538 0 51594 800 6 wbs_dat_i[5]
port 508 nsew default input
rlabel metal2 s 57334 0 57390 800 6 wbs_dat_i[6]
port 509 nsew default input
rlabel metal2 s 63222 0 63278 800 6 wbs_dat_i[7]
port 510 nsew default input
rlabel metal2 s 69018 0 69074 800 6 wbs_dat_i[8]
port 511 nsew default input
rlabel metal2 s 74906 0 74962 800 6 wbs_dat_i[9]
port 512 nsew default input
rlabel metal2 s 16486 0 16542 800 6 wbs_dat_o[0]
port 513 nsew default output
rlabel metal2 s 82634 0 82690 800 6 wbs_dat_o[10]
port 514 nsew default output
rlabel metal2 s 88522 0 88578 800 6 wbs_dat_o[11]
port 515 nsew default output
rlabel metal2 s 94318 0 94374 800 6 wbs_dat_o[12]
port 516 nsew default output
rlabel metal2 s 100206 0 100262 800 6 wbs_dat_o[13]
port 517 nsew default output
rlabel metal2 s 106002 0 106058 800 6 wbs_dat_o[14]
port 518 nsew default output
rlabel metal2 s 111890 0 111946 800 6 wbs_dat_o[15]
port 519 nsew default output
rlabel metal2 s 117686 0 117742 800 6 wbs_dat_o[16]
port 520 nsew default output
rlabel metal2 s 123574 0 123630 800 6 wbs_dat_o[17]
port 521 nsew default output
rlabel metal2 s 129370 0 129426 800 6 wbs_dat_o[18]
port 522 nsew default output
rlabel metal2 s 135166 0 135222 800 6 wbs_dat_o[19]
port 523 nsew default output
rlabel metal2 s 24214 0 24270 800 6 wbs_dat_o[1]
port 524 nsew default output
rlabel metal2 s 141054 0 141110 800 6 wbs_dat_o[20]
port 525 nsew default output
rlabel metal2 s 146850 0 146906 800 6 wbs_dat_o[21]
port 526 nsew default output
rlabel metal2 s 152738 0 152794 800 6 wbs_dat_o[22]
port 527 nsew default output
rlabel metal2 s 158534 0 158590 800 6 wbs_dat_o[23]
port 528 nsew default output
rlabel metal2 s 164422 0 164478 800 6 wbs_dat_o[24]
port 529 nsew default output
rlabel metal2 s 170218 0 170274 800 6 wbs_dat_o[25]
port 530 nsew default output
rlabel metal2 s 176106 0 176162 800 6 wbs_dat_o[26]
port 531 nsew default output
rlabel metal2 s 181902 0 181958 800 6 wbs_dat_o[27]
port 532 nsew default output
rlabel metal2 s 187790 0 187846 800 6 wbs_dat_o[28]
port 533 nsew default output
rlabel metal2 s 193586 0 193642 800 6 wbs_dat_o[29]
port 534 nsew default output
rlabel metal2 s 32034 0 32090 800 6 wbs_dat_o[2]
port 535 nsew default output
rlabel metal2 s 199474 0 199530 800 6 wbs_dat_o[30]
port 536 nsew default output
rlabel metal2 s 205270 0 205326 800 6 wbs_dat_o[31]
port 537 nsew default output
rlabel metal2 s 39854 0 39910 800 6 wbs_dat_o[3]
port 538 nsew default output
rlabel metal2 s 47582 0 47638 800 6 wbs_dat_o[4]
port 539 nsew default output
rlabel metal2 s 53470 0 53526 800 6 wbs_dat_o[5]
port 540 nsew default output
rlabel metal2 s 59266 0 59322 800 6 wbs_dat_o[6]
port 541 nsew default output
rlabel metal2 s 65154 0 65210 800 6 wbs_dat_o[7]
port 542 nsew default output
rlabel metal2 s 70950 0 71006 800 6 wbs_dat_o[8]
port 543 nsew default output
rlabel metal2 s 76838 0 76894 800 6 wbs_dat_o[9]
port 544 nsew default output
rlabel metal2 s 18418 0 18474 800 6 wbs_sel_i[0]
port 545 nsew default input
rlabel metal2 s 26238 0 26294 800 6 wbs_sel_i[1]
port 546 nsew default input
rlabel metal2 s 33966 0 34022 800 6 wbs_sel_i[2]
port 547 nsew default input
rlabel metal2 s 41786 0 41842 800 6 wbs_sel_i[3]
port 548 nsew default input
rlabel metal2 s 8666 0 8722 800 6 wbs_stb_i
port 549 nsew default input
rlabel metal2 s 10598 0 10654 800 6 wbs_we_i
port 550 nsew default input
rlabel metal3 s 219200 416 220000 536 6 zero
port 551 nsew default output
rlabel metal4 s 4208 2128 4528 217648 6 VPWR
port 552 nsew power input
rlabel metal4 s 19568 2128 19888 217648 6 VGND
port 553 nsew ground input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 220000 220000
string LEFview TRUE
<< end >>
