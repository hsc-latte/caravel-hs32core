magic
tech sky130A
magscale 1 2
timestamp 1607833730
<< obsli1 >>
rect 1090 2159 218854 217617
<< obsm1 >>
rect 0 2128 219300 219156
<< metal2 >>
rect 1016 219200 1072 220000
rect 3040 219200 3096 220000
rect 5156 219200 5212 220000
rect 7180 219200 7236 220000
rect 9296 219200 9352 220000
rect 11320 219200 11376 220000
rect 13436 219200 13492 220000
rect 15460 219200 15516 220000
rect 17576 219200 17632 220000
rect 19692 219200 19748 220000
rect 21716 219200 21772 220000
rect 23832 219200 23888 220000
rect 25856 219200 25912 220000
rect 27972 219200 28028 220000
rect 29996 219200 30052 220000
rect 32112 219200 32168 220000
rect 34136 219200 34192 220000
rect 36252 219200 36308 220000
rect 38368 219200 38424 220000
rect 40392 219200 40448 220000
rect 42508 219200 42564 220000
rect 44532 219200 44588 220000
rect 46648 219200 46704 220000
rect 48672 219200 48728 220000
rect 50788 219200 50844 220000
rect 52812 219200 52868 220000
rect 54928 219200 54984 220000
rect 57044 219200 57100 220000
rect 59068 219200 59124 220000
rect 61184 219200 61240 220000
rect 63208 219200 63264 220000
rect 65324 219200 65380 220000
rect 67348 219200 67404 220000
rect 69464 219200 69520 220000
rect 71488 219200 71544 220000
rect 73604 219200 73660 220000
rect 75720 219200 75776 220000
rect 77744 219200 77800 220000
rect 79860 219200 79916 220000
rect 81884 219200 81940 220000
rect 84000 219200 84056 220000
rect 86024 219200 86080 220000
rect 88140 219200 88196 220000
rect 90164 219200 90220 220000
rect 92280 219200 92336 220000
rect 94396 219200 94452 220000
rect 96420 219200 96476 220000
rect 98536 219200 98592 220000
rect 100560 219200 100616 220000
rect 102676 219200 102732 220000
rect 104700 219200 104756 220000
rect 106816 219200 106872 220000
rect 108840 219200 108896 220000
rect 110956 219200 111012 220000
rect 113072 219200 113128 220000
rect 115096 219200 115152 220000
rect 117212 219200 117268 220000
rect 119236 219200 119292 220000
rect 121352 219200 121408 220000
rect 123376 219200 123432 220000
rect 125492 219200 125548 220000
rect 127516 219200 127572 220000
rect 129632 219200 129688 220000
rect 131748 219200 131804 220000
rect 133772 219200 133828 220000
rect 135888 219200 135944 220000
rect 137912 219200 137968 220000
rect 140028 219200 140084 220000
rect 142052 219200 142108 220000
rect 144168 219200 144224 220000
rect 146192 219200 146248 220000
rect 148308 219200 148364 220000
rect 150424 219200 150480 220000
rect 152448 219200 152504 220000
rect 154564 219200 154620 220000
rect 156588 219200 156644 220000
rect 158704 219200 158760 220000
rect 160728 219200 160784 220000
rect 162844 219200 162900 220000
rect 164868 219200 164924 220000
rect 166984 219200 167040 220000
rect 169100 219200 169156 220000
rect 171124 219200 171180 220000
rect 173240 219200 173296 220000
rect 175264 219200 175320 220000
rect 177380 219200 177436 220000
rect 179404 219200 179460 220000
rect 181520 219200 181576 220000
rect 183544 219200 183600 220000
rect 185660 219200 185716 220000
rect 187776 219200 187832 220000
rect 189800 219200 189856 220000
rect 191916 219200 191972 220000
rect 193940 219200 193996 220000
rect 196056 219200 196112 220000
rect 198080 219200 198136 220000
rect 200196 219200 200252 220000
rect 202220 219200 202276 220000
rect 204336 219200 204392 220000
rect 206452 219200 206508 220000
rect 208476 219200 208532 220000
rect 210592 219200 210648 220000
rect 212616 219200 212672 220000
rect 214732 219200 214788 220000
rect 216756 219200 216812 220000
rect 218872 219200 218928 220000
rect 188 0 244 800
rect 556 0 612 800
rect 1016 0 1072 800
rect 1476 0 1532 800
rect 1936 0 1992 800
rect 2396 0 2452 800
rect 2856 0 2912 800
rect 3316 0 3372 800
rect 3776 0 3832 800
rect 4144 0 4200 800
rect 4604 0 4660 800
rect 5064 0 5120 800
rect 5524 0 5580 800
rect 5984 0 6040 800
rect 6444 0 6500 800
rect 6904 0 6960 800
rect 7364 0 7420 800
rect 7732 0 7788 800
rect 8192 0 8248 800
rect 8652 0 8708 800
rect 9112 0 9168 800
rect 9572 0 9628 800
rect 10032 0 10088 800
rect 10492 0 10548 800
rect 10952 0 11008 800
rect 11320 0 11376 800
rect 11780 0 11836 800
rect 12240 0 12296 800
rect 12700 0 12756 800
rect 13160 0 13216 800
rect 13620 0 13676 800
rect 14080 0 14136 800
rect 14540 0 14596 800
rect 15000 0 15056 800
rect 15368 0 15424 800
rect 15828 0 15884 800
rect 16288 0 16344 800
rect 16748 0 16804 800
rect 17208 0 17264 800
rect 17668 0 17724 800
rect 18128 0 18184 800
rect 18588 0 18644 800
rect 18956 0 19012 800
rect 19416 0 19472 800
rect 19876 0 19932 800
rect 20336 0 20392 800
rect 20796 0 20852 800
rect 21256 0 21312 800
rect 21716 0 21772 800
rect 22176 0 22232 800
rect 22544 0 22600 800
rect 23004 0 23060 800
rect 23464 0 23520 800
rect 23924 0 23980 800
rect 24384 0 24440 800
rect 24844 0 24900 800
rect 25304 0 25360 800
rect 25764 0 25820 800
rect 26224 0 26280 800
rect 26592 0 26648 800
rect 27052 0 27108 800
rect 27512 0 27568 800
rect 27972 0 28028 800
rect 28432 0 28488 800
rect 28892 0 28948 800
rect 29352 0 29408 800
rect 29812 0 29868 800
rect 30180 0 30236 800
rect 30640 0 30696 800
rect 31100 0 31156 800
rect 31560 0 31616 800
rect 32020 0 32076 800
rect 32480 0 32536 800
rect 32940 0 32996 800
rect 33400 0 33456 800
rect 33768 0 33824 800
rect 34228 0 34284 800
rect 34688 0 34744 800
rect 35148 0 35204 800
rect 35608 0 35664 800
rect 36068 0 36124 800
rect 36528 0 36584 800
rect 36988 0 37044 800
rect 37448 0 37504 800
rect 37816 0 37872 800
rect 38276 0 38332 800
rect 38736 0 38792 800
rect 39196 0 39252 800
rect 39656 0 39712 800
rect 40116 0 40172 800
rect 40576 0 40632 800
rect 41036 0 41092 800
rect 41404 0 41460 800
rect 41864 0 41920 800
rect 42324 0 42380 800
rect 42784 0 42840 800
rect 43244 0 43300 800
rect 43704 0 43760 800
rect 44164 0 44220 800
rect 44624 0 44680 800
rect 44992 0 45048 800
rect 45452 0 45508 800
rect 45912 0 45968 800
rect 46372 0 46428 800
rect 46832 0 46888 800
rect 47292 0 47348 800
rect 47752 0 47808 800
rect 48212 0 48268 800
rect 48580 0 48636 800
rect 49040 0 49096 800
rect 49500 0 49556 800
rect 49960 0 50016 800
rect 50420 0 50476 800
rect 50880 0 50936 800
rect 51340 0 51396 800
rect 51800 0 51856 800
rect 52260 0 52316 800
rect 52628 0 52684 800
rect 53088 0 53144 800
rect 53548 0 53604 800
rect 54008 0 54064 800
rect 54468 0 54524 800
rect 54928 0 54984 800
rect 55388 0 55444 800
rect 55848 0 55904 800
rect 56216 0 56272 800
rect 56676 0 56732 800
rect 57136 0 57192 800
rect 57596 0 57652 800
rect 58056 0 58112 800
rect 58516 0 58572 800
rect 58976 0 59032 800
rect 59436 0 59492 800
rect 59804 0 59860 800
rect 60264 0 60320 800
rect 60724 0 60780 800
rect 61184 0 61240 800
rect 61644 0 61700 800
rect 62104 0 62160 800
rect 62564 0 62620 800
rect 63024 0 63080 800
rect 63484 0 63540 800
rect 63852 0 63908 800
rect 64312 0 64368 800
rect 64772 0 64828 800
rect 65232 0 65288 800
rect 65692 0 65748 800
rect 66152 0 66208 800
rect 66612 0 66668 800
rect 67072 0 67128 800
rect 67440 0 67496 800
rect 67900 0 67956 800
rect 68360 0 68416 800
rect 68820 0 68876 800
rect 69280 0 69336 800
rect 69740 0 69796 800
rect 70200 0 70256 800
rect 70660 0 70716 800
rect 71028 0 71084 800
rect 71488 0 71544 800
rect 71948 0 72004 800
rect 72408 0 72464 800
rect 72868 0 72924 800
rect 73328 0 73384 800
rect 73788 0 73844 800
rect 74248 0 74304 800
rect 74708 0 74764 800
rect 75076 0 75132 800
rect 75536 0 75592 800
rect 75996 0 76052 800
rect 76456 0 76512 800
rect 76916 0 76972 800
rect 77376 0 77432 800
rect 77836 0 77892 800
rect 78296 0 78352 800
rect 78664 0 78720 800
rect 79124 0 79180 800
rect 79584 0 79640 800
rect 80044 0 80100 800
rect 80504 0 80560 800
rect 80964 0 81020 800
rect 81424 0 81480 800
rect 81884 0 81940 800
rect 82252 0 82308 800
rect 82712 0 82768 800
rect 83172 0 83228 800
rect 83632 0 83688 800
rect 84092 0 84148 800
rect 84552 0 84608 800
rect 85012 0 85068 800
rect 85472 0 85528 800
rect 85932 0 85988 800
rect 86300 0 86356 800
rect 86760 0 86816 800
rect 87220 0 87276 800
rect 87680 0 87736 800
rect 88140 0 88196 800
rect 88600 0 88656 800
rect 89060 0 89116 800
rect 89520 0 89576 800
rect 89888 0 89944 800
rect 90348 0 90404 800
rect 90808 0 90864 800
rect 91268 0 91324 800
rect 91728 0 91784 800
rect 92188 0 92244 800
rect 92648 0 92704 800
rect 93108 0 93164 800
rect 93476 0 93532 800
rect 93936 0 93992 800
rect 94396 0 94452 800
rect 94856 0 94912 800
rect 95316 0 95372 800
rect 95776 0 95832 800
rect 96236 0 96292 800
rect 96696 0 96752 800
rect 97064 0 97120 800
rect 97524 0 97580 800
rect 97984 0 98040 800
rect 98444 0 98500 800
rect 98904 0 98960 800
rect 99364 0 99420 800
rect 99824 0 99880 800
rect 100284 0 100340 800
rect 100744 0 100800 800
rect 101112 0 101168 800
rect 101572 0 101628 800
rect 102032 0 102088 800
rect 102492 0 102548 800
rect 102952 0 103008 800
rect 103412 0 103468 800
rect 103872 0 103928 800
rect 104332 0 104388 800
rect 104700 0 104756 800
rect 105160 0 105216 800
rect 105620 0 105676 800
rect 106080 0 106136 800
rect 106540 0 106596 800
rect 107000 0 107056 800
rect 107460 0 107516 800
rect 107920 0 107976 800
rect 108288 0 108344 800
rect 108748 0 108804 800
rect 109208 0 109264 800
rect 109668 0 109724 800
rect 110128 0 110184 800
rect 110588 0 110644 800
rect 111048 0 111104 800
rect 111508 0 111564 800
rect 111968 0 112024 800
rect 112336 0 112392 800
rect 112796 0 112852 800
rect 113256 0 113312 800
rect 113716 0 113772 800
rect 114176 0 114232 800
rect 114636 0 114692 800
rect 115096 0 115152 800
rect 115556 0 115612 800
rect 115924 0 115980 800
rect 116384 0 116440 800
rect 116844 0 116900 800
rect 117304 0 117360 800
rect 117764 0 117820 800
rect 118224 0 118280 800
rect 118684 0 118740 800
rect 119144 0 119200 800
rect 119512 0 119568 800
rect 119972 0 120028 800
rect 120432 0 120488 800
rect 120892 0 120948 800
rect 121352 0 121408 800
rect 121812 0 121868 800
rect 122272 0 122328 800
rect 122732 0 122788 800
rect 123192 0 123248 800
rect 123560 0 123616 800
rect 124020 0 124076 800
rect 124480 0 124536 800
rect 124940 0 124996 800
rect 125400 0 125456 800
rect 125860 0 125916 800
rect 126320 0 126376 800
rect 126780 0 126836 800
rect 127148 0 127204 800
rect 127608 0 127664 800
rect 128068 0 128124 800
rect 128528 0 128584 800
rect 128988 0 129044 800
rect 129448 0 129504 800
rect 129908 0 129964 800
rect 130368 0 130424 800
rect 130736 0 130792 800
rect 131196 0 131252 800
rect 131656 0 131712 800
rect 132116 0 132172 800
rect 132576 0 132632 800
rect 133036 0 133092 800
rect 133496 0 133552 800
rect 133956 0 134012 800
rect 134324 0 134380 800
rect 134784 0 134840 800
rect 135244 0 135300 800
rect 135704 0 135760 800
rect 136164 0 136220 800
rect 136624 0 136680 800
rect 137084 0 137140 800
rect 137544 0 137600 800
rect 138004 0 138060 800
rect 138372 0 138428 800
rect 138832 0 138888 800
rect 139292 0 139348 800
rect 139752 0 139808 800
rect 140212 0 140268 800
rect 140672 0 140728 800
rect 141132 0 141188 800
rect 141592 0 141648 800
rect 141960 0 142016 800
rect 142420 0 142476 800
rect 142880 0 142936 800
rect 143340 0 143396 800
rect 143800 0 143856 800
rect 144260 0 144316 800
rect 144720 0 144776 800
rect 145180 0 145236 800
rect 145548 0 145604 800
rect 146008 0 146064 800
rect 146468 0 146524 800
rect 146928 0 146984 800
rect 147388 0 147444 800
rect 147848 0 147904 800
rect 148308 0 148364 800
rect 148768 0 148824 800
rect 149228 0 149284 800
rect 149596 0 149652 800
rect 150056 0 150112 800
rect 150516 0 150572 800
rect 150976 0 151032 800
rect 151436 0 151492 800
rect 151896 0 151952 800
rect 152356 0 152412 800
rect 152816 0 152872 800
rect 153184 0 153240 800
rect 153644 0 153700 800
rect 154104 0 154160 800
rect 154564 0 154620 800
rect 155024 0 155080 800
rect 155484 0 155540 800
rect 155944 0 156000 800
rect 156404 0 156460 800
rect 156772 0 156828 800
rect 157232 0 157288 800
rect 157692 0 157748 800
rect 158152 0 158208 800
rect 158612 0 158668 800
rect 159072 0 159128 800
rect 159532 0 159588 800
rect 159992 0 160048 800
rect 160452 0 160508 800
rect 160820 0 160876 800
rect 161280 0 161336 800
rect 161740 0 161796 800
rect 162200 0 162256 800
rect 162660 0 162716 800
rect 163120 0 163176 800
rect 163580 0 163636 800
rect 164040 0 164096 800
rect 164408 0 164464 800
rect 164868 0 164924 800
rect 165328 0 165384 800
rect 165788 0 165844 800
rect 166248 0 166304 800
rect 166708 0 166764 800
rect 167168 0 167224 800
rect 167628 0 167684 800
rect 167996 0 168052 800
rect 168456 0 168512 800
rect 168916 0 168972 800
rect 169376 0 169432 800
rect 169836 0 169892 800
rect 170296 0 170352 800
rect 170756 0 170812 800
rect 171216 0 171272 800
rect 171676 0 171732 800
rect 172044 0 172100 800
rect 172504 0 172560 800
rect 172964 0 173020 800
rect 173424 0 173480 800
rect 173884 0 173940 800
rect 174344 0 174400 800
rect 174804 0 174860 800
rect 175264 0 175320 800
rect 175632 0 175688 800
rect 176092 0 176148 800
rect 176552 0 176608 800
rect 177012 0 177068 800
rect 177472 0 177528 800
rect 177932 0 177988 800
rect 178392 0 178448 800
rect 178852 0 178908 800
rect 179220 0 179276 800
rect 179680 0 179736 800
rect 180140 0 180196 800
rect 180600 0 180656 800
rect 181060 0 181116 800
rect 181520 0 181576 800
rect 181980 0 182036 800
rect 182440 0 182496 800
rect 182808 0 182864 800
rect 183268 0 183324 800
rect 183728 0 183784 800
rect 184188 0 184244 800
rect 184648 0 184704 800
rect 185108 0 185164 800
rect 185568 0 185624 800
rect 186028 0 186084 800
rect 186488 0 186544 800
rect 186856 0 186912 800
rect 187316 0 187372 800
rect 187776 0 187832 800
rect 188236 0 188292 800
rect 188696 0 188752 800
rect 189156 0 189212 800
rect 189616 0 189672 800
rect 190076 0 190132 800
rect 190444 0 190500 800
rect 190904 0 190960 800
rect 191364 0 191420 800
rect 191824 0 191880 800
rect 192284 0 192340 800
rect 192744 0 192800 800
rect 193204 0 193260 800
rect 193664 0 193720 800
rect 194032 0 194088 800
rect 194492 0 194548 800
rect 194952 0 195008 800
rect 195412 0 195468 800
rect 195872 0 195928 800
rect 196332 0 196388 800
rect 196792 0 196848 800
rect 197252 0 197308 800
rect 197712 0 197768 800
rect 198080 0 198136 800
rect 198540 0 198596 800
rect 199000 0 199056 800
rect 199460 0 199516 800
rect 199920 0 199976 800
rect 200380 0 200436 800
rect 200840 0 200896 800
rect 201300 0 201356 800
rect 201668 0 201724 800
rect 202128 0 202184 800
rect 202588 0 202644 800
rect 203048 0 203104 800
rect 203508 0 203564 800
rect 203968 0 204024 800
rect 204428 0 204484 800
rect 204888 0 204944 800
rect 205256 0 205312 800
rect 205716 0 205772 800
rect 206176 0 206232 800
rect 206636 0 206692 800
rect 207096 0 207152 800
rect 207556 0 207612 800
rect 208016 0 208072 800
rect 208476 0 208532 800
rect 208936 0 208992 800
rect 209304 0 209360 800
rect 209764 0 209820 800
rect 210224 0 210280 800
rect 210684 0 210740 800
rect 211144 0 211200 800
rect 211604 0 211660 800
rect 212064 0 212120 800
rect 212524 0 212580 800
rect 212892 0 212948 800
rect 213352 0 213408 800
rect 213812 0 213868 800
rect 214272 0 214328 800
rect 214732 0 214788 800
rect 215192 0 215248 800
rect 215652 0 215708 800
rect 216112 0 216168 800
rect 216480 0 216536 800
rect 216940 0 216996 800
rect 217400 0 217456 800
rect 217860 0 217916 800
rect 218320 0 218376 800
rect 218780 0 218836 800
rect 219240 0 219296 800
rect 219700 0 219756 800
<< obsm2 >>
rect 6 219144 960 219200
rect 1128 219144 2984 219200
rect 3152 219144 5100 219200
rect 5268 219144 7124 219200
rect 7292 219144 9240 219200
rect 9408 219144 11264 219200
rect 11432 219144 13380 219200
rect 13548 219144 15404 219200
rect 15572 219144 17520 219200
rect 17688 219144 19636 219200
rect 19804 219144 21660 219200
rect 21828 219144 23776 219200
rect 23944 219144 25800 219200
rect 25968 219144 27916 219200
rect 28084 219144 29940 219200
rect 30108 219144 32056 219200
rect 32224 219144 34080 219200
rect 34248 219144 36196 219200
rect 36364 219144 38312 219200
rect 38480 219144 40336 219200
rect 40504 219144 42452 219200
rect 42620 219144 44476 219200
rect 44644 219144 46592 219200
rect 46760 219144 48616 219200
rect 48784 219144 50732 219200
rect 50900 219144 52756 219200
rect 52924 219144 54872 219200
rect 55040 219144 56988 219200
rect 57156 219144 59012 219200
rect 59180 219144 61128 219200
rect 61296 219144 63152 219200
rect 63320 219144 65268 219200
rect 65436 219144 67292 219200
rect 67460 219144 69408 219200
rect 69576 219144 71432 219200
rect 71600 219144 73548 219200
rect 73716 219144 75664 219200
rect 75832 219144 77688 219200
rect 77856 219144 79804 219200
rect 79972 219144 81828 219200
rect 81996 219144 83944 219200
rect 84112 219144 85968 219200
rect 86136 219144 88084 219200
rect 88252 219144 90108 219200
rect 90276 219144 92224 219200
rect 92392 219144 94340 219200
rect 94508 219144 96364 219200
rect 96532 219144 98480 219200
rect 98648 219144 100504 219200
rect 100672 219144 102620 219200
rect 102788 219144 104644 219200
rect 104812 219144 106760 219200
rect 106928 219144 108784 219200
rect 108952 219144 110900 219200
rect 111068 219144 113016 219200
rect 113184 219144 115040 219200
rect 115208 219144 117156 219200
rect 117324 219144 119180 219200
rect 119348 219144 121296 219200
rect 121464 219144 123320 219200
rect 123488 219144 125436 219200
rect 125604 219144 127460 219200
rect 127628 219144 129576 219200
rect 129744 219144 131692 219200
rect 131860 219144 133716 219200
rect 133884 219144 135832 219200
rect 136000 219144 137856 219200
rect 138024 219144 139972 219200
rect 140140 219144 141996 219200
rect 142164 219144 144112 219200
rect 144280 219144 146136 219200
rect 146304 219144 148252 219200
rect 148420 219144 150368 219200
rect 150536 219144 152392 219200
rect 152560 219144 154508 219200
rect 154676 219144 156532 219200
rect 156700 219144 158648 219200
rect 158816 219144 160672 219200
rect 160840 219144 162788 219200
rect 162956 219144 164812 219200
rect 164980 219144 166928 219200
rect 167096 219144 169044 219200
rect 169212 219144 171068 219200
rect 171236 219144 173184 219200
rect 173352 219144 175208 219200
rect 175376 219144 177324 219200
rect 177492 219144 179348 219200
rect 179516 219144 181464 219200
rect 181632 219144 183488 219200
rect 183656 219144 185604 219200
rect 185772 219144 187720 219200
rect 187888 219144 189744 219200
rect 189912 219144 191860 219200
rect 192028 219144 193884 219200
rect 194052 219144 196000 219200
rect 196168 219144 198024 219200
rect 198192 219144 200140 219200
rect 200308 219144 202164 219200
rect 202332 219144 204280 219200
rect 204448 219144 206396 219200
rect 206564 219144 208420 219200
rect 208588 219144 210536 219200
rect 210704 219144 212560 219200
rect 212728 219144 214676 219200
rect 214844 219144 216700 219200
rect 216868 219144 218816 219200
rect 218984 219144 219294 219200
rect 6 856 219294 219144
rect 6 800 132 856
rect 300 800 500 856
rect 668 800 960 856
rect 1128 800 1420 856
rect 1588 800 1880 856
rect 2048 800 2340 856
rect 2508 800 2800 856
rect 2968 800 3260 856
rect 3428 800 3720 856
rect 3888 800 4088 856
rect 4256 800 4548 856
rect 4716 800 5008 856
rect 5176 800 5468 856
rect 5636 800 5928 856
rect 6096 800 6388 856
rect 6556 800 6848 856
rect 7016 800 7308 856
rect 7476 800 7676 856
rect 7844 800 8136 856
rect 8304 800 8596 856
rect 8764 800 9056 856
rect 9224 800 9516 856
rect 9684 800 9976 856
rect 10144 800 10436 856
rect 10604 800 10896 856
rect 11064 800 11264 856
rect 11432 800 11724 856
rect 11892 800 12184 856
rect 12352 800 12644 856
rect 12812 800 13104 856
rect 13272 800 13564 856
rect 13732 800 14024 856
rect 14192 800 14484 856
rect 14652 800 14944 856
rect 15112 800 15312 856
rect 15480 800 15772 856
rect 15940 800 16232 856
rect 16400 800 16692 856
rect 16860 800 17152 856
rect 17320 800 17612 856
rect 17780 800 18072 856
rect 18240 800 18532 856
rect 18700 800 18900 856
rect 19068 800 19360 856
rect 19528 800 19820 856
rect 19988 800 20280 856
rect 20448 800 20740 856
rect 20908 800 21200 856
rect 21368 800 21660 856
rect 21828 800 22120 856
rect 22288 800 22488 856
rect 22656 800 22948 856
rect 23116 800 23408 856
rect 23576 800 23868 856
rect 24036 800 24328 856
rect 24496 800 24788 856
rect 24956 800 25248 856
rect 25416 800 25708 856
rect 25876 800 26168 856
rect 26336 800 26536 856
rect 26704 800 26996 856
rect 27164 800 27456 856
rect 27624 800 27916 856
rect 28084 800 28376 856
rect 28544 800 28836 856
rect 29004 800 29296 856
rect 29464 800 29756 856
rect 29924 800 30124 856
rect 30292 800 30584 856
rect 30752 800 31044 856
rect 31212 800 31504 856
rect 31672 800 31964 856
rect 32132 800 32424 856
rect 32592 800 32884 856
rect 33052 800 33344 856
rect 33512 800 33712 856
rect 33880 800 34172 856
rect 34340 800 34632 856
rect 34800 800 35092 856
rect 35260 800 35552 856
rect 35720 800 36012 856
rect 36180 800 36472 856
rect 36640 800 36932 856
rect 37100 800 37392 856
rect 37560 800 37760 856
rect 37928 800 38220 856
rect 38388 800 38680 856
rect 38848 800 39140 856
rect 39308 800 39600 856
rect 39768 800 40060 856
rect 40228 800 40520 856
rect 40688 800 40980 856
rect 41148 800 41348 856
rect 41516 800 41808 856
rect 41976 800 42268 856
rect 42436 800 42728 856
rect 42896 800 43188 856
rect 43356 800 43648 856
rect 43816 800 44108 856
rect 44276 800 44568 856
rect 44736 800 44936 856
rect 45104 800 45396 856
rect 45564 800 45856 856
rect 46024 800 46316 856
rect 46484 800 46776 856
rect 46944 800 47236 856
rect 47404 800 47696 856
rect 47864 800 48156 856
rect 48324 800 48524 856
rect 48692 800 48984 856
rect 49152 800 49444 856
rect 49612 800 49904 856
rect 50072 800 50364 856
rect 50532 800 50824 856
rect 50992 800 51284 856
rect 51452 800 51744 856
rect 51912 800 52204 856
rect 52372 800 52572 856
rect 52740 800 53032 856
rect 53200 800 53492 856
rect 53660 800 53952 856
rect 54120 800 54412 856
rect 54580 800 54872 856
rect 55040 800 55332 856
rect 55500 800 55792 856
rect 55960 800 56160 856
rect 56328 800 56620 856
rect 56788 800 57080 856
rect 57248 800 57540 856
rect 57708 800 58000 856
rect 58168 800 58460 856
rect 58628 800 58920 856
rect 59088 800 59380 856
rect 59548 800 59748 856
rect 59916 800 60208 856
rect 60376 800 60668 856
rect 60836 800 61128 856
rect 61296 800 61588 856
rect 61756 800 62048 856
rect 62216 800 62508 856
rect 62676 800 62968 856
rect 63136 800 63428 856
rect 63596 800 63796 856
rect 63964 800 64256 856
rect 64424 800 64716 856
rect 64884 800 65176 856
rect 65344 800 65636 856
rect 65804 800 66096 856
rect 66264 800 66556 856
rect 66724 800 67016 856
rect 67184 800 67384 856
rect 67552 800 67844 856
rect 68012 800 68304 856
rect 68472 800 68764 856
rect 68932 800 69224 856
rect 69392 800 69684 856
rect 69852 800 70144 856
rect 70312 800 70604 856
rect 70772 800 70972 856
rect 71140 800 71432 856
rect 71600 800 71892 856
rect 72060 800 72352 856
rect 72520 800 72812 856
rect 72980 800 73272 856
rect 73440 800 73732 856
rect 73900 800 74192 856
rect 74360 800 74652 856
rect 74820 800 75020 856
rect 75188 800 75480 856
rect 75648 800 75940 856
rect 76108 800 76400 856
rect 76568 800 76860 856
rect 77028 800 77320 856
rect 77488 800 77780 856
rect 77948 800 78240 856
rect 78408 800 78608 856
rect 78776 800 79068 856
rect 79236 800 79528 856
rect 79696 800 79988 856
rect 80156 800 80448 856
rect 80616 800 80908 856
rect 81076 800 81368 856
rect 81536 800 81828 856
rect 81996 800 82196 856
rect 82364 800 82656 856
rect 82824 800 83116 856
rect 83284 800 83576 856
rect 83744 800 84036 856
rect 84204 800 84496 856
rect 84664 800 84956 856
rect 85124 800 85416 856
rect 85584 800 85876 856
rect 86044 800 86244 856
rect 86412 800 86704 856
rect 86872 800 87164 856
rect 87332 800 87624 856
rect 87792 800 88084 856
rect 88252 800 88544 856
rect 88712 800 89004 856
rect 89172 800 89464 856
rect 89632 800 89832 856
rect 90000 800 90292 856
rect 90460 800 90752 856
rect 90920 800 91212 856
rect 91380 800 91672 856
rect 91840 800 92132 856
rect 92300 800 92592 856
rect 92760 800 93052 856
rect 93220 800 93420 856
rect 93588 800 93880 856
rect 94048 800 94340 856
rect 94508 800 94800 856
rect 94968 800 95260 856
rect 95428 800 95720 856
rect 95888 800 96180 856
rect 96348 800 96640 856
rect 96808 800 97008 856
rect 97176 800 97468 856
rect 97636 800 97928 856
rect 98096 800 98388 856
rect 98556 800 98848 856
rect 99016 800 99308 856
rect 99476 800 99768 856
rect 99936 800 100228 856
rect 100396 800 100688 856
rect 100856 800 101056 856
rect 101224 800 101516 856
rect 101684 800 101976 856
rect 102144 800 102436 856
rect 102604 800 102896 856
rect 103064 800 103356 856
rect 103524 800 103816 856
rect 103984 800 104276 856
rect 104444 800 104644 856
rect 104812 800 105104 856
rect 105272 800 105564 856
rect 105732 800 106024 856
rect 106192 800 106484 856
rect 106652 800 106944 856
rect 107112 800 107404 856
rect 107572 800 107864 856
rect 108032 800 108232 856
rect 108400 800 108692 856
rect 108860 800 109152 856
rect 109320 800 109612 856
rect 109780 800 110072 856
rect 110240 800 110532 856
rect 110700 800 110992 856
rect 111160 800 111452 856
rect 111620 800 111912 856
rect 112080 800 112280 856
rect 112448 800 112740 856
rect 112908 800 113200 856
rect 113368 800 113660 856
rect 113828 800 114120 856
rect 114288 800 114580 856
rect 114748 800 115040 856
rect 115208 800 115500 856
rect 115668 800 115868 856
rect 116036 800 116328 856
rect 116496 800 116788 856
rect 116956 800 117248 856
rect 117416 800 117708 856
rect 117876 800 118168 856
rect 118336 800 118628 856
rect 118796 800 119088 856
rect 119256 800 119456 856
rect 119624 800 119916 856
rect 120084 800 120376 856
rect 120544 800 120836 856
rect 121004 800 121296 856
rect 121464 800 121756 856
rect 121924 800 122216 856
rect 122384 800 122676 856
rect 122844 800 123136 856
rect 123304 800 123504 856
rect 123672 800 123964 856
rect 124132 800 124424 856
rect 124592 800 124884 856
rect 125052 800 125344 856
rect 125512 800 125804 856
rect 125972 800 126264 856
rect 126432 800 126724 856
rect 126892 800 127092 856
rect 127260 800 127552 856
rect 127720 800 128012 856
rect 128180 800 128472 856
rect 128640 800 128932 856
rect 129100 800 129392 856
rect 129560 800 129852 856
rect 130020 800 130312 856
rect 130480 800 130680 856
rect 130848 800 131140 856
rect 131308 800 131600 856
rect 131768 800 132060 856
rect 132228 800 132520 856
rect 132688 800 132980 856
rect 133148 800 133440 856
rect 133608 800 133900 856
rect 134068 800 134268 856
rect 134436 800 134728 856
rect 134896 800 135188 856
rect 135356 800 135648 856
rect 135816 800 136108 856
rect 136276 800 136568 856
rect 136736 800 137028 856
rect 137196 800 137488 856
rect 137656 800 137948 856
rect 138116 800 138316 856
rect 138484 800 138776 856
rect 138944 800 139236 856
rect 139404 800 139696 856
rect 139864 800 140156 856
rect 140324 800 140616 856
rect 140784 800 141076 856
rect 141244 800 141536 856
rect 141704 800 141904 856
rect 142072 800 142364 856
rect 142532 800 142824 856
rect 142992 800 143284 856
rect 143452 800 143744 856
rect 143912 800 144204 856
rect 144372 800 144664 856
rect 144832 800 145124 856
rect 145292 800 145492 856
rect 145660 800 145952 856
rect 146120 800 146412 856
rect 146580 800 146872 856
rect 147040 800 147332 856
rect 147500 800 147792 856
rect 147960 800 148252 856
rect 148420 800 148712 856
rect 148880 800 149172 856
rect 149340 800 149540 856
rect 149708 800 150000 856
rect 150168 800 150460 856
rect 150628 800 150920 856
rect 151088 800 151380 856
rect 151548 800 151840 856
rect 152008 800 152300 856
rect 152468 800 152760 856
rect 152928 800 153128 856
rect 153296 800 153588 856
rect 153756 800 154048 856
rect 154216 800 154508 856
rect 154676 800 154968 856
rect 155136 800 155428 856
rect 155596 800 155888 856
rect 156056 800 156348 856
rect 156516 800 156716 856
rect 156884 800 157176 856
rect 157344 800 157636 856
rect 157804 800 158096 856
rect 158264 800 158556 856
rect 158724 800 159016 856
rect 159184 800 159476 856
rect 159644 800 159936 856
rect 160104 800 160396 856
rect 160564 800 160764 856
rect 160932 800 161224 856
rect 161392 800 161684 856
rect 161852 800 162144 856
rect 162312 800 162604 856
rect 162772 800 163064 856
rect 163232 800 163524 856
rect 163692 800 163984 856
rect 164152 800 164352 856
rect 164520 800 164812 856
rect 164980 800 165272 856
rect 165440 800 165732 856
rect 165900 800 166192 856
rect 166360 800 166652 856
rect 166820 800 167112 856
rect 167280 800 167572 856
rect 167740 800 167940 856
rect 168108 800 168400 856
rect 168568 800 168860 856
rect 169028 800 169320 856
rect 169488 800 169780 856
rect 169948 800 170240 856
rect 170408 800 170700 856
rect 170868 800 171160 856
rect 171328 800 171620 856
rect 171788 800 171988 856
rect 172156 800 172448 856
rect 172616 800 172908 856
rect 173076 800 173368 856
rect 173536 800 173828 856
rect 173996 800 174288 856
rect 174456 800 174748 856
rect 174916 800 175208 856
rect 175376 800 175576 856
rect 175744 800 176036 856
rect 176204 800 176496 856
rect 176664 800 176956 856
rect 177124 800 177416 856
rect 177584 800 177876 856
rect 178044 800 178336 856
rect 178504 800 178796 856
rect 178964 800 179164 856
rect 179332 800 179624 856
rect 179792 800 180084 856
rect 180252 800 180544 856
rect 180712 800 181004 856
rect 181172 800 181464 856
rect 181632 800 181924 856
rect 182092 800 182384 856
rect 182552 800 182752 856
rect 182920 800 183212 856
rect 183380 800 183672 856
rect 183840 800 184132 856
rect 184300 800 184592 856
rect 184760 800 185052 856
rect 185220 800 185512 856
rect 185680 800 185972 856
rect 186140 800 186432 856
rect 186600 800 186800 856
rect 186968 800 187260 856
rect 187428 800 187720 856
rect 187888 800 188180 856
rect 188348 800 188640 856
rect 188808 800 189100 856
rect 189268 800 189560 856
rect 189728 800 190020 856
rect 190188 800 190388 856
rect 190556 800 190848 856
rect 191016 800 191308 856
rect 191476 800 191768 856
rect 191936 800 192228 856
rect 192396 800 192688 856
rect 192856 800 193148 856
rect 193316 800 193608 856
rect 193776 800 193976 856
rect 194144 800 194436 856
rect 194604 800 194896 856
rect 195064 800 195356 856
rect 195524 800 195816 856
rect 195984 800 196276 856
rect 196444 800 196736 856
rect 196904 800 197196 856
rect 197364 800 197656 856
rect 197824 800 198024 856
rect 198192 800 198484 856
rect 198652 800 198944 856
rect 199112 800 199404 856
rect 199572 800 199864 856
rect 200032 800 200324 856
rect 200492 800 200784 856
rect 200952 800 201244 856
rect 201412 800 201612 856
rect 201780 800 202072 856
rect 202240 800 202532 856
rect 202700 800 202992 856
rect 203160 800 203452 856
rect 203620 800 203912 856
rect 204080 800 204372 856
rect 204540 800 204832 856
rect 205000 800 205200 856
rect 205368 800 205660 856
rect 205828 800 206120 856
rect 206288 800 206580 856
rect 206748 800 207040 856
rect 207208 800 207500 856
rect 207668 800 207960 856
rect 208128 800 208420 856
rect 208588 800 208880 856
rect 209048 800 209248 856
rect 209416 800 209708 856
rect 209876 800 210168 856
rect 210336 800 210628 856
rect 210796 800 211088 856
rect 211256 800 211548 856
rect 211716 800 212008 856
rect 212176 800 212468 856
rect 212636 800 212836 856
rect 213004 800 213296 856
rect 213464 800 213756 856
rect 213924 800 214216 856
rect 214384 800 214676 856
rect 214844 800 215136 856
rect 215304 800 215596 856
rect 215764 800 216056 856
rect 216224 800 216424 856
rect 216592 800 216884 856
rect 217052 800 217344 856
rect 217512 800 217804 856
rect 217972 800 218264 856
rect 218432 800 218724 856
rect 218892 800 219184 856
<< metal3 >>
rect 219186 218968 219986 219088
rect 219186 216928 219986 217048
rect 219186 214888 219986 215008
rect 219186 212848 219986 212968
rect 219186 210808 219986 210928
rect 219186 208768 219986 208888
rect 219186 206728 219986 206848
rect 219186 204688 219986 204808
rect 219186 202648 219986 202768
rect 219186 200608 219986 200728
rect 219186 198568 219986 198688
rect 219186 196528 219986 196648
rect 219186 194488 219986 194608
rect 219186 192448 219986 192568
rect 219186 190408 219986 190528
rect 219186 188368 219986 188488
rect 219186 186328 219986 186448
rect 219186 184288 219986 184408
rect 219186 182248 219986 182368
rect 219186 180208 219986 180328
rect 219186 178168 219986 178288
rect 219186 176128 219986 176248
rect 219186 174088 219986 174208
rect 219186 172048 219986 172168
rect 219186 170008 219986 170128
rect 219186 167968 219986 168088
rect 219186 165928 219986 166048
rect 219186 163888 219986 164008
rect 219186 161848 219986 161968
rect 219186 159808 219986 159928
rect 219186 157768 219986 157888
rect 219186 155728 219986 155848
rect 219186 153688 219986 153808
rect 219186 151648 219986 151768
rect 219186 149608 219986 149728
rect 219186 147568 219986 147688
rect 219186 145528 219986 145648
rect 219186 143488 219986 143608
rect 219186 141448 219986 141568
rect 219186 139408 219986 139528
rect 219186 137368 219986 137488
rect 219186 135328 219986 135448
rect 219186 133288 219986 133408
rect 219186 131248 219986 131368
rect 219186 129208 219986 129328
rect 219186 127168 219986 127288
rect 219186 125128 219986 125248
rect 219186 123088 219986 123208
rect 219186 121048 219986 121168
rect 219186 119008 219986 119128
rect 219186 116968 219986 117088
rect 219186 114928 219986 115048
rect 219186 112888 219986 113008
rect 219186 110984 219986 111104
rect 219186 108944 219986 109064
rect 219186 106904 219986 107024
rect 219186 104864 219986 104984
rect 219186 102824 219986 102944
rect 219186 100784 219986 100904
rect 219186 98744 219986 98864
rect 219186 96704 219986 96824
rect 219186 94664 219986 94784
rect 219186 92624 219986 92744
rect 219186 90584 219986 90704
rect 219186 88544 219986 88664
rect 219186 86504 219986 86624
rect 219186 84464 219986 84584
rect 219186 82424 219986 82544
rect 219186 80384 219986 80504
rect 219186 78344 219986 78464
rect 219186 76304 219986 76424
rect 219186 74264 219986 74384
rect 219186 72224 219986 72344
rect 219186 70184 219986 70304
rect 219186 68144 219986 68264
rect 219186 66104 219986 66224
rect 219186 64064 219986 64184
rect 219186 62024 219986 62144
rect 219186 59984 219986 60104
rect 219186 57944 219986 58064
rect 219186 55904 219986 56024
rect 219186 53864 219986 53984
rect 219186 51824 219986 51944
rect 219186 49784 219986 49904
rect 219186 47744 219986 47864
rect 219186 45704 219986 45824
rect 219186 43664 219986 43784
rect 219186 41624 219986 41744
rect 219186 39584 219986 39704
rect 219186 37544 219986 37664
rect 219186 35504 219986 35624
rect 219186 33464 219986 33584
rect 219186 31424 219986 31544
rect 219186 29384 219986 29504
rect 219186 27344 219986 27464
rect 219186 25304 219986 25424
rect 219186 23264 219986 23384
rect 219186 21224 219986 21344
rect 219186 19184 219986 19304
rect 219186 17144 219986 17264
rect 219186 15104 219986 15224
rect 219186 13064 219986 13184
rect 219186 11024 219986 11144
rect 219186 8984 219986 9104
rect 219186 6944 219986 7064
rect 219186 4904 219986 5024
rect 219186 2864 219986 2984
rect 219186 960 219986 1080
<< obsm3 >>
rect 183 218888 219106 219061
rect 183 217128 219186 218888
rect 183 216848 219106 217128
rect 183 215088 219186 216848
rect 183 214808 219106 215088
rect 183 213048 219186 214808
rect 183 212768 219106 213048
rect 183 211008 219186 212768
rect 183 210728 219106 211008
rect 183 208968 219186 210728
rect 183 208688 219106 208968
rect 183 206928 219186 208688
rect 183 206648 219106 206928
rect 183 204888 219186 206648
rect 183 204608 219106 204888
rect 183 202848 219186 204608
rect 183 202568 219106 202848
rect 183 200808 219186 202568
rect 183 200528 219106 200808
rect 183 198768 219186 200528
rect 183 198488 219106 198768
rect 183 196728 219186 198488
rect 183 196448 219106 196728
rect 183 194688 219186 196448
rect 183 194408 219106 194688
rect 183 192648 219186 194408
rect 183 192368 219106 192648
rect 183 190608 219186 192368
rect 183 190328 219106 190608
rect 183 188568 219186 190328
rect 183 188288 219106 188568
rect 183 186528 219186 188288
rect 183 186248 219106 186528
rect 183 184488 219186 186248
rect 183 184208 219106 184488
rect 183 182448 219186 184208
rect 183 182168 219106 182448
rect 183 180408 219186 182168
rect 183 180128 219106 180408
rect 183 178368 219186 180128
rect 183 178088 219106 178368
rect 183 176328 219186 178088
rect 183 176048 219106 176328
rect 183 174288 219186 176048
rect 183 174008 219106 174288
rect 183 172248 219186 174008
rect 183 171968 219106 172248
rect 183 170208 219186 171968
rect 183 169928 219106 170208
rect 183 168168 219186 169928
rect 183 167888 219106 168168
rect 183 166128 219186 167888
rect 183 165848 219106 166128
rect 183 164088 219186 165848
rect 183 163808 219106 164088
rect 183 162048 219186 163808
rect 183 161768 219106 162048
rect 183 160008 219186 161768
rect 183 159728 219106 160008
rect 183 157968 219186 159728
rect 183 157688 219106 157968
rect 183 155928 219186 157688
rect 183 155648 219106 155928
rect 183 153888 219186 155648
rect 183 153608 219106 153888
rect 183 151848 219186 153608
rect 183 151568 219106 151848
rect 183 149808 219186 151568
rect 183 149528 219106 149808
rect 183 147768 219186 149528
rect 183 147488 219106 147768
rect 183 145728 219186 147488
rect 183 145448 219106 145728
rect 183 143688 219186 145448
rect 183 143408 219106 143688
rect 183 141648 219186 143408
rect 183 141368 219106 141648
rect 183 139608 219186 141368
rect 183 139328 219106 139608
rect 183 137568 219186 139328
rect 183 137288 219106 137568
rect 183 135528 219186 137288
rect 183 135248 219106 135528
rect 183 133488 219186 135248
rect 183 133208 219106 133488
rect 183 131448 219186 133208
rect 183 131168 219106 131448
rect 183 129408 219186 131168
rect 183 129128 219106 129408
rect 183 127368 219186 129128
rect 183 127088 219106 127368
rect 183 125328 219186 127088
rect 183 125048 219106 125328
rect 183 123288 219186 125048
rect 183 123008 219106 123288
rect 183 121248 219186 123008
rect 183 120968 219106 121248
rect 183 119208 219186 120968
rect 183 118928 219106 119208
rect 183 117168 219186 118928
rect 183 116888 219106 117168
rect 183 115128 219186 116888
rect 183 114848 219106 115128
rect 183 113088 219186 114848
rect 183 112808 219106 113088
rect 183 111184 219186 112808
rect 183 110904 219106 111184
rect 183 109144 219186 110904
rect 183 108864 219106 109144
rect 183 107104 219186 108864
rect 183 106824 219106 107104
rect 183 105064 219186 106824
rect 183 104784 219106 105064
rect 183 103024 219186 104784
rect 183 102744 219106 103024
rect 183 100984 219186 102744
rect 183 100704 219106 100984
rect 183 98944 219186 100704
rect 183 98664 219106 98944
rect 183 96904 219186 98664
rect 183 96624 219106 96904
rect 183 94864 219186 96624
rect 183 94584 219106 94864
rect 183 92824 219186 94584
rect 183 92544 219106 92824
rect 183 90784 219186 92544
rect 183 90504 219106 90784
rect 183 88744 219186 90504
rect 183 88464 219106 88744
rect 183 86704 219186 88464
rect 183 86424 219106 86704
rect 183 84664 219186 86424
rect 183 84384 219106 84664
rect 183 82624 219186 84384
rect 183 82344 219106 82624
rect 183 80584 219186 82344
rect 183 80304 219106 80584
rect 183 78544 219186 80304
rect 183 78264 219106 78544
rect 183 76504 219186 78264
rect 183 76224 219106 76504
rect 183 74464 219186 76224
rect 183 74184 219106 74464
rect 183 72424 219186 74184
rect 183 72144 219106 72424
rect 183 70384 219186 72144
rect 183 70104 219106 70384
rect 183 68344 219186 70104
rect 183 68064 219106 68344
rect 183 66304 219186 68064
rect 183 66024 219106 66304
rect 183 64264 219186 66024
rect 183 63984 219106 64264
rect 183 62224 219186 63984
rect 183 61944 219106 62224
rect 183 60184 219186 61944
rect 183 59904 219106 60184
rect 183 58144 219186 59904
rect 183 57864 219106 58144
rect 183 56104 219186 57864
rect 183 55824 219106 56104
rect 183 54064 219186 55824
rect 183 53784 219106 54064
rect 183 52024 219186 53784
rect 183 51744 219106 52024
rect 183 49984 219186 51744
rect 183 49704 219106 49984
rect 183 47944 219186 49704
rect 183 47664 219106 47944
rect 183 45904 219186 47664
rect 183 45624 219106 45904
rect 183 43864 219186 45624
rect 183 43584 219106 43864
rect 183 41824 219186 43584
rect 183 41544 219106 41824
rect 183 39784 219186 41544
rect 183 39504 219106 39784
rect 183 37744 219186 39504
rect 183 37464 219106 37744
rect 183 35704 219186 37464
rect 183 35424 219106 35704
rect 183 33664 219186 35424
rect 183 33384 219106 33664
rect 183 31624 219186 33384
rect 183 31344 219106 31624
rect 183 29584 219186 31344
rect 183 29304 219106 29584
rect 183 27544 219186 29304
rect 183 27264 219106 27544
rect 183 25504 219186 27264
rect 183 25224 219106 25504
rect 183 23464 219186 25224
rect 183 23184 219106 23464
rect 183 21424 219186 23184
rect 183 21144 219106 21424
rect 183 19384 219186 21144
rect 183 19104 219106 19384
rect 183 17344 219186 19104
rect 183 17064 219106 17344
rect 183 15304 219186 17064
rect 183 15024 219106 15304
rect 183 13264 219186 15024
rect 183 12984 219106 13264
rect 183 11224 219186 12984
rect 183 10944 219106 11224
rect 183 9184 219186 10944
rect 183 8904 219106 9184
rect 183 7144 219186 8904
rect 183 6864 219106 7144
rect 183 5104 219186 6864
rect 183 4824 219106 5104
rect 183 3064 219186 4824
rect 183 2784 219106 3064
rect 183 1160 219186 2784
rect 183 987 219106 1160
<< metal4 >>
rect 4194 2128 4514 217648
rect 19554 2128 19874 217648
<< obsm4 >>
rect 13293 2128 19474 217648
rect 19954 2128 217599 217648
<< labels >>
rlabel metal3 s 219186 25304 219986 25424 6 cpu_addr_e[0]
port 1 nsew default output
rlabel metal3 s 219186 45704 219986 45824 6 cpu_addr_e[10]
port 2 nsew default output
rlabel metal3 s 219186 47744 219986 47864 6 cpu_addr_e[11]
port 3 nsew default output
rlabel metal3 s 219186 49784 219986 49904 6 cpu_addr_e[12]
port 4 nsew default output
rlabel metal3 s 219186 51824 219986 51944 6 cpu_addr_e[13]
port 5 nsew default output
rlabel metal3 s 219186 53864 219986 53984 6 cpu_addr_e[14]
port 6 nsew default output
rlabel metal3 s 219186 55904 219986 56024 6 cpu_addr_e[15]
port 7 nsew default output
rlabel metal3 s 219186 27344 219986 27464 6 cpu_addr_e[1]
port 8 nsew default output
rlabel metal3 s 219186 29384 219986 29504 6 cpu_addr_e[2]
port 9 nsew default output
rlabel metal3 s 219186 31424 219986 31544 6 cpu_addr_e[3]
port 10 nsew default output
rlabel metal3 s 219186 33464 219986 33584 6 cpu_addr_e[4]
port 11 nsew default output
rlabel metal3 s 219186 35504 219986 35624 6 cpu_addr_e[5]
port 12 nsew default output
rlabel metal3 s 219186 37544 219986 37664 6 cpu_addr_e[6]
port 13 nsew default output
rlabel metal3 s 219186 39584 219986 39704 6 cpu_addr_e[7]
port 14 nsew default output
rlabel metal3 s 219186 41624 219986 41744 6 cpu_addr_e[8]
port 15 nsew default output
rlabel metal3 s 219186 43664 219986 43784 6 cpu_addr_e[9]
port 16 nsew default output
rlabel metal2 s 21716 219200 21772 220000 6 cpu_addr_n[0]
port 17 nsew default output
rlabel metal2 s 42508 219200 42564 220000 6 cpu_addr_n[10]
port 18 nsew default output
rlabel metal2 s 44532 219200 44588 220000 6 cpu_addr_n[11]
port 19 nsew default output
rlabel metal2 s 46648 219200 46704 220000 6 cpu_addr_n[12]
port 20 nsew default output
rlabel metal2 s 48672 219200 48728 220000 6 cpu_addr_n[13]
port 21 nsew default output
rlabel metal2 s 50788 219200 50844 220000 6 cpu_addr_n[14]
port 22 nsew default output
rlabel metal2 s 52812 219200 52868 220000 6 cpu_addr_n[15]
port 23 nsew default output
rlabel metal2 s 23832 219200 23888 220000 6 cpu_addr_n[1]
port 24 nsew default output
rlabel metal2 s 25856 219200 25912 220000 6 cpu_addr_n[2]
port 25 nsew default output
rlabel metal2 s 27972 219200 28028 220000 6 cpu_addr_n[3]
port 26 nsew default output
rlabel metal2 s 29996 219200 30052 220000 6 cpu_addr_n[4]
port 27 nsew default output
rlabel metal2 s 32112 219200 32168 220000 6 cpu_addr_n[5]
port 28 nsew default output
rlabel metal2 s 34136 219200 34192 220000 6 cpu_addr_n[6]
port 29 nsew default output
rlabel metal2 s 36252 219200 36308 220000 6 cpu_addr_n[7]
port 30 nsew default output
rlabel metal2 s 38368 219200 38424 220000 6 cpu_addr_n[8]
port 31 nsew default output
rlabel metal2 s 40392 219200 40448 220000 6 cpu_addr_n[9]
port 32 nsew default output
rlabel metal3 s 219186 90584 219986 90704 6 cpu_dtr_e0[0]
port 33 nsew default input
rlabel metal3 s 219186 110984 219986 111104 6 cpu_dtr_e0[10]
port 34 nsew default input
rlabel metal3 s 219186 112888 219986 113008 6 cpu_dtr_e0[11]
port 35 nsew default input
rlabel metal3 s 219186 114928 219986 115048 6 cpu_dtr_e0[12]
port 36 nsew default input
rlabel metal3 s 219186 116968 219986 117088 6 cpu_dtr_e0[13]
port 37 nsew default input
rlabel metal3 s 219186 119008 219986 119128 6 cpu_dtr_e0[14]
port 38 nsew default input
rlabel metal3 s 219186 121048 219986 121168 6 cpu_dtr_e0[15]
port 39 nsew default input
rlabel metal3 s 219186 123088 219986 123208 6 cpu_dtr_e0[16]
port 40 nsew default input
rlabel metal3 s 219186 125128 219986 125248 6 cpu_dtr_e0[17]
port 41 nsew default input
rlabel metal3 s 219186 127168 219986 127288 6 cpu_dtr_e0[18]
port 42 nsew default input
rlabel metal3 s 219186 129208 219986 129328 6 cpu_dtr_e0[19]
port 43 nsew default input
rlabel metal3 s 219186 92624 219986 92744 6 cpu_dtr_e0[1]
port 44 nsew default input
rlabel metal3 s 219186 131248 219986 131368 6 cpu_dtr_e0[20]
port 45 nsew default input
rlabel metal3 s 219186 133288 219986 133408 6 cpu_dtr_e0[21]
port 46 nsew default input
rlabel metal3 s 219186 135328 219986 135448 6 cpu_dtr_e0[22]
port 47 nsew default input
rlabel metal3 s 219186 137368 219986 137488 6 cpu_dtr_e0[23]
port 48 nsew default input
rlabel metal3 s 219186 139408 219986 139528 6 cpu_dtr_e0[24]
port 49 nsew default input
rlabel metal3 s 219186 141448 219986 141568 6 cpu_dtr_e0[25]
port 50 nsew default input
rlabel metal3 s 219186 143488 219986 143608 6 cpu_dtr_e0[26]
port 51 nsew default input
rlabel metal3 s 219186 145528 219986 145648 6 cpu_dtr_e0[27]
port 52 nsew default input
rlabel metal3 s 219186 147568 219986 147688 6 cpu_dtr_e0[28]
port 53 nsew default input
rlabel metal3 s 219186 149608 219986 149728 6 cpu_dtr_e0[29]
port 54 nsew default input
rlabel metal3 s 219186 94664 219986 94784 6 cpu_dtr_e0[2]
port 55 nsew default input
rlabel metal3 s 219186 151648 219986 151768 6 cpu_dtr_e0[30]
port 56 nsew default input
rlabel metal3 s 219186 153688 219986 153808 6 cpu_dtr_e0[31]
port 57 nsew default input
rlabel metal3 s 219186 96704 219986 96824 6 cpu_dtr_e0[3]
port 58 nsew default input
rlabel metal3 s 219186 98744 219986 98864 6 cpu_dtr_e0[4]
port 59 nsew default input
rlabel metal3 s 219186 100784 219986 100904 6 cpu_dtr_e0[5]
port 60 nsew default input
rlabel metal3 s 219186 102824 219986 102944 6 cpu_dtr_e0[6]
port 61 nsew default input
rlabel metal3 s 219186 104864 219986 104984 6 cpu_dtr_e0[7]
port 62 nsew default input
rlabel metal3 s 219186 106904 219986 107024 6 cpu_dtr_e0[8]
port 63 nsew default input
rlabel metal3 s 219186 108944 219986 109064 6 cpu_dtr_e0[9]
port 64 nsew default input
rlabel metal3 s 219186 155728 219986 155848 6 cpu_dtr_e1[0]
port 65 nsew default input
rlabel metal3 s 219186 176128 219986 176248 6 cpu_dtr_e1[10]
port 66 nsew default input
rlabel metal3 s 219186 178168 219986 178288 6 cpu_dtr_e1[11]
port 67 nsew default input
rlabel metal3 s 219186 180208 219986 180328 6 cpu_dtr_e1[12]
port 68 nsew default input
rlabel metal3 s 219186 182248 219986 182368 6 cpu_dtr_e1[13]
port 69 nsew default input
rlabel metal3 s 219186 184288 219986 184408 6 cpu_dtr_e1[14]
port 70 nsew default input
rlabel metal3 s 219186 186328 219986 186448 6 cpu_dtr_e1[15]
port 71 nsew default input
rlabel metal3 s 219186 188368 219986 188488 6 cpu_dtr_e1[16]
port 72 nsew default input
rlabel metal3 s 219186 190408 219986 190528 6 cpu_dtr_e1[17]
port 73 nsew default input
rlabel metal3 s 219186 192448 219986 192568 6 cpu_dtr_e1[18]
port 74 nsew default input
rlabel metal3 s 219186 194488 219986 194608 6 cpu_dtr_e1[19]
port 75 nsew default input
rlabel metal3 s 219186 157768 219986 157888 6 cpu_dtr_e1[1]
port 76 nsew default input
rlabel metal3 s 219186 196528 219986 196648 6 cpu_dtr_e1[20]
port 77 nsew default input
rlabel metal3 s 219186 198568 219986 198688 6 cpu_dtr_e1[21]
port 78 nsew default input
rlabel metal3 s 219186 200608 219986 200728 6 cpu_dtr_e1[22]
port 79 nsew default input
rlabel metal3 s 219186 202648 219986 202768 6 cpu_dtr_e1[23]
port 80 nsew default input
rlabel metal3 s 219186 204688 219986 204808 6 cpu_dtr_e1[24]
port 81 nsew default input
rlabel metal3 s 219186 206728 219986 206848 6 cpu_dtr_e1[25]
port 82 nsew default input
rlabel metal3 s 219186 208768 219986 208888 6 cpu_dtr_e1[26]
port 83 nsew default input
rlabel metal3 s 219186 210808 219986 210928 6 cpu_dtr_e1[27]
port 84 nsew default input
rlabel metal3 s 219186 212848 219986 212968 6 cpu_dtr_e1[28]
port 85 nsew default input
rlabel metal3 s 219186 214888 219986 215008 6 cpu_dtr_e1[29]
port 86 nsew default input
rlabel metal3 s 219186 159808 219986 159928 6 cpu_dtr_e1[2]
port 87 nsew default input
rlabel metal3 s 219186 216928 219986 217048 6 cpu_dtr_e1[30]
port 88 nsew default input
rlabel metal3 s 219186 218968 219986 219088 6 cpu_dtr_e1[31]
port 89 nsew default input
rlabel metal3 s 219186 161848 219986 161968 6 cpu_dtr_e1[3]
port 90 nsew default input
rlabel metal3 s 219186 163888 219986 164008 6 cpu_dtr_e1[4]
port 91 nsew default input
rlabel metal3 s 219186 165928 219986 166048 6 cpu_dtr_e1[5]
port 92 nsew default input
rlabel metal3 s 219186 167968 219986 168088 6 cpu_dtr_e1[6]
port 93 nsew default input
rlabel metal3 s 219186 170008 219986 170128 6 cpu_dtr_e1[7]
port 94 nsew default input
rlabel metal3 s 219186 172048 219986 172168 6 cpu_dtr_e1[8]
port 95 nsew default input
rlabel metal3 s 219186 174088 219986 174208 6 cpu_dtr_e1[9]
port 96 nsew default input
rlabel metal2 s 88140 219200 88196 220000 6 cpu_dtr_n0[0]
port 97 nsew default input
rlabel metal2 s 108840 219200 108896 220000 6 cpu_dtr_n0[10]
port 98 nsew default input
rlabel metal2 s 110956 219200 111012 220000 6 cpu_dtr_n0[11]
port 99 nsew default input
rlabel metal2 s 113072 219200 113128 220000 6 cpu_dtr_n0[12]
port 100 nsew default input
rlabel metal2 s 115096 219200 115152 220000 6 cpu_dtr_n0[13]
port 101 nsew default input
rlabel metal2 s 117212 219200 117268 220000 6 cpu_dtr_n0[14]
port 102 nsew default input
rlabel metal2 s 119236 219200 119292 220000 6 cpu_dtr_n0[15]
port 103 nsew default input
rlabel metal2 s 121352 219200 121408 220000 6 cpu_dtr_n0[16]
port 104 nsew default input
rlabel metal2 s 123376 219200 123432 220000 6 cpu_dtr_n0[17]
port 105 nsew default input
rlabel metal2 s 125492 219200 125548 220000 6 cpu_dtr_n0[18]
port 106 nsew default input
rlabel metal2 s 127516 219200 127572 220000 6 cpu_dtr_n0[19]
port 107 nsew default input
rlabel metal2 s 90164 219200 90220 220000 6 cpu_dtr_n0[1]
port 108 nsew default input
rlabel metal2 s 129632 219200 129688 220000 6 cpu_dtr_n0[20]
port 109 nsew default input
rlabel metal2 s 131748 219200 131804 220000 6 cpu_dtr_n0[21]
port 110 nsew default input
rlabel metal2 s 133772 219200 133828 220000 6 cpu_dtr_n0[22]
port 111 nsew default input
rlabel metal2 s 135888 219200 135944 220000 6 cpu_dtr_n0[23]
port 112 nsew default input
rlabel metal2 s 137912 219200 137968 220000 6 cpu_dtr_n0[24]
port 113 nsew default input
rlabel metal2 s 140028 219200 140084 220000 6 cpu_dtr_n0[25]
port 114 nsew default input
rlabel metal2 s 142052 219200 142108 220000 6 cpu_dtr_n0[26]
port 115 nsew default input
rlabel metal2 s 144168 219200 144224 220000 6 cpu_dtr_n0[27]
port 116 nsew default input
rlabel metal2 s 146192 219200 146248 220000 6 cpu_dtr_n0[28]
port 117 nsew default input
rlabel metal2 s 148308 219200 148364 220000 6 cpu_dtr_n0[29]
port 118 nsew default input
rlabel metal2 s 92280 219200 92336 220000 6 cpu_dtr_n0[2]
port 119 nsew default input
rlabel metal2 s 150424 219200 150480 220000 6 cpu_dtr_n0[30]
port 120 nsew default input
rlabel metal2 s 152448 219200 152504 220000 6 cpu_dtr_n0[31]
port 121 nsew default input
rlabel metal2 s 94396 219200 94452 220000 6 cpu_dtr_n0[3]
port 122 nsew default input
rlabel metal2 s 96420 219200 96476 220000 6 cpu_dtr_n0[4]
port 123 nsew default input
rlabel metal2 s 98536 219200 98592 220000 6 cpu_dtr_n0[5]
port 124 nsew default input
rlabel metal2 s 100560 219200 100616 220000 6 cpu_dtr_n0[6]
port 125 nsew default input
rlabel metal2 s 102676 219200 102732 220000 6 cpu_dtr_n0[7]
port 126 nsew default input
rlabel metal2 s 104700 219200 104756 220000 6 cpu_dtr_n0[8]
port 127 nsew default input
rlabel metal2 s 106816 219200 106872 220000 6 cpu_dtr_n0[9]
port 128 nsew default input
rlabel metal2 s 154564 219200 154620 220000 6 cpu_dtr_n1[0]
port 129 nsew default input
rlabel metal2 s 175264 219200 175320 220000 6 cpu_dtr_n1[10]
port 130 nsew default input
rlabel metal2 s 177380 219200 177436 220000 6 cpu_dtr_n1[11]
port 131 nsew default input
rlabel metal2 s 179404 219200 179460 220000 6 cpu_dtr_n1[12]
port 132 nsew default input
rlabel metal2 s 181520 219200 181576 220000 6 cpu_dtr_n1[13]
port 133 nsew default input
rlabel metal2 s 183544 219200 183600 220000 6 cpu_dtr_n1[14]
port 134 nsew default input
rlabel metal2 s 185660 219200 185716 220000 6 cpu_dtr_n1[15]
port 135 nsew default input
rlabel metal2 s 187776 219200 187832 220000 6 cpu_dtr_n1[16]
port 136 nsew default input
rlabel metal2 s 189800 219200 189856 220000 6 cpu_dtr_n1[17]
port 137 nsew default input
rlabel metal2 s 191916 219200 191972 220000 6 cpu_dtr_n1[18]
port 138 nsew default input
rlabel metal2 s 193940 219200 193996 220000 6 cpu_dtr_n1[19]
port 139 nsew default input
rlabel metal2 s 156588 219200 156644 220000 6 cpu_dtr_n1[1]
port 140 nsew default input
rlabel metal2 s 196056 219200 196112 220000 6 cpu_dtr_n1[20]
port 141 nsew default input
rlabel metal2 s 198080 219200 198136 220000 6 cpu_dtr_n1[21]
port 142 nsew default input
rlabel metal2 s 200196 219200 200252 220000 6 cpu_dtr_n1[22]
port 143 nsew default input
rlabel metal2 s 202220 219200 202276 220000 6 cpu_dtr_n1[23]
port 144 nsew default input
rlabel metal2 s 204336 219200 204392 220000 6 cpu_dtr_n1[24]
port 145 nsew default input
rlabel metal2 s 206452 219200 206508 220000 6 cpu_dtr_n1[25]
port 146 nsew default input
rlabel metal2 s 208476 219200 208532 220000 6 cpu_dtr_n1[26]
port 147 nsew default input
rlabel metal2 s 210592 219200 210648 220000 6 cpu_dtr_n1[27]
port 148 nsew default input
rlabel metal2 s 212616 219200 212672 220000 6 cpu_dtr_n1[28]
port 149 nsew default input
rlabel metal2 s 214732 219200 214788 220000 6 cpu_dtr_n1[29]
port 150 nsew default input
rlabel metal2 s 158704 219200 158760 220000 6 cpu_dtr_n1[2]
port 151 nsew default input
rlabel metal2 s 216756 219200 216812 220000 6 cpu_dtr_n1[30]
port 152 nsew default input
rlabel metal2 s 218872 219200 218928 220000 6 cpu_dtr_n1[31]
port 153 nsew default input
rlabel metal2 s 160728 219200 160784 220000 6 cpu_dtr_n1[3]
port 154 nsew default input
rlabel metal2 s 162844 219200 162900 220000 6 cpu_dtr_n1[4]
port 155 nsew default input
rlabel metal2 s 164868 219200 164924 220000 6 cpu_dtr_n1[5]
port 156 nsew default input
rlabel metal2 s 166984 219200 167040 220000 6 cpu_dtr_n1[6]
port 157 nsew default input
rlabel metal2 s 169100 219200 169156 220000 6 cpu_dtr_n1[7]
port 158 nsew default input
rlabel metal2 s 171124 219200 171180 220000 6 cpu_dtr_n1[8]
port 159 nsew default input
rlabel metal2 s 173240 219200 173296 220000 6 cpu_dtr_n1[9]
port 160 nsew default input
rlabel metal3 s 219186 57944 219986 58064 6 cpu_dtw_e[0]
port 161 nsew default output
rlabel metal3 s 219186 78344 219986 78464 6 cpu_dtw_e[10]
port 162 nsew default output
rlabel metal3 s 219186 80384 219986 80504 6 cpu_dtw_e[11]
port 163 nsew default output
rlabel metal3 s 219186 82424 219986 82544 6 cpu_dtw_e[12]
port 164 nsew default output
rlabel metal3 s 219186 84464 219986 84584 6 cpu_dtw_e[13]
port 165 nsew default output
rlabel metal3 s 219186 86504 219986 86624 6 cpu_dtw_e[14]
port 166 nsew default output
rlabel metal3 s 219186 88544 219986 88664 6 cpu_dtw_e[15]
port 167 nsew default output
rlabel metal3 s 219186 59984 219986 60104 6 cpu_dtw_e[1]
port 168 nsew default output
rlabel metal3 s 219186 62024 219986 62144 6 cpu_dtw_e[2]
port 169 nsew default output
rlabel metal3 s 219186 64064 219986 64184 6 cpu_dtw_e[3]
port 170 nsew default output
rlabel metal3 s 219186 66104 219986 66224 6 cpu_dtw_e[4]
port 171 nsew default output
rlabel metal3 s 219186 68144 219986 68264 6 cpu_dtw_e[5]
port 172 nsew default output
rlabel metal3 s 219186 70184 219986 70304 6 cpu_dtw_e[6]
port 173 nsew default output
rlabel metal3 s 219186 72224 219986 72344 6 cpu_dtw_e[7]
port 174 nsew default output
rlabel metal3 s 219186 74264 219986 74384 6 cpu_dtw_e[8]
port 175 nsew default output
rlabel metal3 s 219186 76304 219986 76424 6 cpu_dtw_e[9]
port 176 nsew default output
rlabel metal2 s 54928 219200 54984 220000 6 cpu_dtw_n[0]
port 177 nsew default output
rlabel metal2 s 75720 219200 75776 220000 6 cpu_dtw_n[10]
port 178 nsew default output
rlabel metal2 s 77744 219200 77800 220000 6 cpu_dtw_n[11]
port 179 nsew default output
rlabel metal2 s 79860 219200 79916 220000 6 cpu_dtw_n[12]
port 180 nsew default output
rlabel metal2 s 81884 219200 81940 220000 6 cpu_dtw_n[13]
port 181 nsew default output
rlabel metal2 s 84000 219200 84056 220000 6 cpu_dtw_n[14]
port 182 nsew default output
rlabel metal2 s 86024 219200 86080 220000 6 cpu_dtw_n[15]
port 183 nsew default output
rlabel metal2 s 57044 219200 57100 220000 6 cpu_dtw_n[1]
port 184 nsew default output
rlabel metal2 s 59068 219200 59124 220000 6 cpu_dtw_n[2]
port 185 nsew default output
rlabel metal2 s 61184 219200 61240 220000 6 cpu_dtw_n[3]
port 186 nsew default output
rlabel metal2 s 63208 219200 63264 220000 6 cpu_dtw_n[4]
port 187 nsew default output
rlabel metal2 s 65324 219200 65380 220000 6 cpu_dtw_n[5]
port 188 nsew default output
rlabel metal2 s 67348 219200 67404 220000 6 cpu_dtw_n[6]
port 189 nsew default output
rlabel metal2 s 69464 219200 69520 220000 6 cpu_dtw_n[7]
port 190 nsew default output
rlabel metal2 s 71488 219200 71544 220000 6 cpu_dtw_n[8]
port 191 nsew default output
rlabel metal2 s 73604 219200 73660 220000 6 cpu_dtw_n[9]
port 192 nsew default output
rlabel metal3 s 219186 4904 219986 5024 6 cpu_mask_e[0]
port 193 nsew default output
rlabel metal3 s 219186 6944 219986 7064 6 cpu_mask_e[1]
port 194 nsew default output
rlabel metal3 s 219186 8984 219986 9104 6 cpu_mask_e[2]
port 195 nsew default output
rlabel metal3 s 219186 11024 219986 11144 6 cpu_mask_e[3]
port 196 nsew default output
rlabel metal3 s 219186 13064 219986 13184 6 cpu_mask_e[4]
port 197 nsew default output
rlabel metal3 s 219186 15104 219986 15224 6 cpu_mask_e[5]
port 198 nsew default output
rlabel metal3 s 219186 17144 219986 17264 6 cpu_mask_e[6]
port 199 nsew default output
rlabel metal3 s 219186 19184 219986 19304 6 cpu_mask_e[7]
port 200 nsew default output
rlabel metal2 s 1016 219200 1072 220000 6 cpu_mask_n[0]
port 201 nsew default output
rlabel metal2 s 3040 219200 3096 220000 6 cpu_mask_n[1]
port 202 nsew default output
rlabel metal2 s 5156 219200 5212 220000 6 cpu_mask_n[2]
port 203 nsew default output
rlabel metal2 s 7180 219200 7236 220000 6 cpu_mask_n[3]
port 204 nsew default output
rlabel metal2 s 9296 219200 9352 220000 6 cpu_mask_n[4]
port 205 nsew default output
rlabel metal2 s 11320 219200 11376 220000 6 cpu_mask_n[5]
port 206 nsew default output
rlabel metal2 s 13436 219200 13492 220000 6 cpu_mask_n[6]
port 207 nsew default output
rlabel metal2 s 15460 219200 15516 220000 6 cpu_mask_n[7]
port 208 nsew default output
rlabel metal3 s 219186 21224 219986 21344 6 cpu_wen_e[0]
port 209 nsew default output
rlabel metal3 s 219186 23264 219986 23384 6 cpu_wen_e[1]
port 210 nsew default output
rlabel metal2 s 17576 219200 17632 220000 6 cpu_wen_n[0]
port 211 nsew default output
rlabel metal2 s 19692 219200 19748 220000 6 cpu_wen_n[1]
port 212 nsew default output
rlabel metal2 s 47752 0 47808 800 6 la_data_in[0]
port 213 nsew default input
rlabel metal2 s 182440 0 182496 800 6 la_data_in[100]
port 214 nsew default input
rlabel metal2 s 183728 0 183784 800 6 la_data_in[101]
port 215 nsew default input
rlabel metal2 s 185108 0 185164 800 6 la_data_in[102]
port 216 nsew default input
rlabel metal2 s 186488 0 186544 800 6 la_data_in[103]
port 217 nsew default input
rlabel metal2 s 187776 0 187832 800 6 la_data_in[104]
port 218 nsew default input
rlabel metal2 s 189156 0 189212 800 6 la_data_in[105]
port 219 nsew default input
rlabel metal2 s 190444 0 190500 800 6 la_data_in[106]
port 220 nsew default input
rlabel metal2 s 191824 0 191880 800 6 la_data_in[107]
port 221 nsew default input
rlabel metal2 s 193204 0 193260 800 6 la_data_in[108]
port 222 nsew default input
rlabel metal2 s 194492 0 194548 800 6 la_data_in[109]
port 223 nsew default input
rlabel metal2 s 61184 0 61240 800 6 la_data_in[10]
port 224 nsew default input
rlabel metal2 s 195872 0 195928 800 6 la_data_in[110]
port 225 nsew default input
rlabel metal2 s 197252 0 197308 800 6 la_data_in[111]
port 226 nsew default input
rlabel metal2 s 198540 0 198596 800 6 la_data_in[112]
port 227 nsew default input
rlabel metal2 s 199920 0 199976 800 6 la_data_in[113]
port 228 nsew default input
rlabel metal2 s 201300 0 201356 800 6 la_data_in[114]
port 229 nsew default input
rlabel metal2 s 202588 0 202644 800 6 la_data_in[115]
port 230 nsew default input
rlabel metal2 s 203968 0 204024 800 6 la_data_in[116]
port 231 nsew default input
rlabel metal2 s 205256 0 205312 800 6 la_data_in[117]
port 232 nsew default input
rlabel metal2 s 206636 0 206692 800 6 la_data_in[118]
port 233 nsew default input
rlabel metal2 s 208016 0 208072 800 6 la_data_in[119]
port 234 nsew default input
rlabel metal2 s 62564 0 62620 800 6 la_data_in[11]
port 235 nsew default input
rlabel metal2 s 209304 0 209360 800 6 la_data_in[120]
port 236 nsew default input
rlabel metal2 s 210684 0 210740 800 6 la_data_in[121]
port 237 nsew default input
rlabel metal2 s 212064 0 212120 800 6 la_data_in[122]
port 238 nsew default input
rlabel metal2 s 213352 0 213408 800 6 la_data_in[123]
port 239 nsew default input
rlabel metal2 s 214732 0 214788 800 6 la_data_in[124]
port 240 nsew default input
rlabel metal2 s 216112 0 216168 800 6 la_data_in[125]
port 241 nsew default input
rlabel metal2 s 217400 0 217456 800 6 la_data_in[126]
port 242 nsew default input
rlabel metal2 s 218780 0 218836 800 6 la_data_in[127]
port 243 nsew default input
rlabel metal2 s 63852 0 63908 800 6 la_data_in[12]
port 244 nsew default input
rlabel metal2 s 65232 0 65288 800 6 la_data_in[13]
port 245 nsew default input
rlabel metal2 s 66612 0 66668 800 6 la_data_in[14]
port 246 nsew default input
rlabel metal2 s 67900 0 67956 800 6 la_data_in[15]
port 247 nsew default input
rlabel metal2 s 69280 0 69336 800 6 la_data_in[16]
port 248 nsew default input
rlabel metal2 s 70660 0 70716 800 6 la_data_in[17]
port 249 nsew default input
rlabel metal2 s 71948 0 72004 800 6 la_data_in[18]
port 250 nsew default input
rlabel metal2 s 73328 0 73384 800 6 la_data_in[19]
port 251 nsew default input
rlabel metal2 s 49040 0 49096 800 6 la_data_in[1]
port 252 nsew default input
rlabel metal2 s 74708 0 74764 800 6 la_data_in[20]
port 253 nsew default input
rlabel metal2 s 75996 0 76052 800 6 la_data_in[21]
port 254 nsew default input
rlabel metal2 s 77376 0 77432 800 6 la_data_in[22]
port 255 nsew default input
rlabel metal2 s 78664 0 78720 800 6 la_data_in[23]
port 256 nsew default input
rlabel metal2 s 80044 0 80100 800 6 la_data_in[24]
port 257 nsew default input
rlabel metal2 s 81424 0 81480 800 6 la_data_in[25]
port 258 nsew default input
rlabel metal2 s 82712 0 82768 800 6 la_data_in[26]
port 259 nsew default input
rlabel metal2 s 84092 0 84148 800 6 la_data_in[27]
port 260 nsew default input
rlabel metal2 s 85472 0 85528 800 6 la_data_in[28]
port 261 nsew default input
rlabel metal2 s 86760 0 86816 800 6 la_data_in[29]
port 262 nsew default input
rlabel metal2 s 50420 0 50476 800 6 la_data_in[2]
port 263 nsew default input
rlabel metal2 s 88140 0 88196 800 6 la_data_in[30]
port 264 nsew default input
rlabel metal2 s 89520 0 89576 800 6 la_data_in[31]
port 265 nsew default input
rlabel metal2 s 90808 0 90864 800 6 la_data_in[32]
port 266 nsew default input
rlabel metal2 s 92188 0 92244 800 6 la_data_in[33]
port 267 nsew default input
rlabel metal2 s 93476 0 93532 800 6 la_data_in[34]
port 268 nsew default input
rlabel metal2 s 94856 0 94912 800 6 la_data_in[35]
port 269 nsew default input
rlabel metal2 s 96236 0 96292 800 6 la_data_in[36]
port 270 nsew default input
rlabel metal2 s 97524 0 97580 800 6 la_data_in[37]
port 271 nsew default input
rlabel metal2 s 98904 0 98960 800 6 la_data_in[38]
port 272 nsew default input
rlabel metal2 s 100284 0 100340 800 6 la_data_in[39]
port 273 nsew default input
rlabel metal2 s 51800 0 51856 800 6 la_data_in[3]
port 274 nsew default input
rlabel metal2 s 101572 0 101628 800 6 la_data_in[40]
port 275 nsew default input
rlabel metal2 s 102952 0 103008 800 6 la_data_in[41]
port 276 nsew default input
rlabel metal2 s 104332 0 104388 800 6 la_data_in[42]
port 277 nsew default input
rlabel metal2 s 105620 0 105676 800 6 la_data_in[43]
port 278 nsew default input
rlabel metal2 s 107000 0 107056 800 6 la_data_in[44]
port 279 nsew default input
rlabel metal2 s 108288 0 108344 800 6 la_data_in[45]
port 280 nsew default input
rlabel metal2 s 109668 0 109724 800 6 la_data_in[46]
port 281 nsew default input
rlabel metal2 s 111048 0 111104 800 6 la_data_in[47]
port 282 nsew default input
rlabel metal2 s 112336 0 112392 800 6 la_data_in[48]
port 283 nsew default input
rlabel metal2 s 113716 0 113772 800 6 la_data_in[49]
port 284 nsew default input
rlabel metal2 s 53088 0 53144 800 6 la_data_in[4]
port 285 nsew default input
rlabel metal2 s 115096 0 115152 800 6 la_data_in[50]
port 286 nsew default input
rlabel metal2 s 116384 0 116440 800 6 la_data_in[51]
port 287 nsew default input
rlabel metal2 s 117764 0 117820 800 6 la_data_in[52]
port 288 nsew default input
rlabel metal2 s 119144 0 119200 800 6 la_data_in[53]
port 289 nsew default input
rlabel metal2 s 120432 0 120488 800 6 la_data_in[54]
port 290 nsew default input
rlabel metal2 s 121812 0 121868 800 6 la_data_in[55]
port 291 nsew default input
rlabel metal2 s 123192 0 123248 800 6 la_data_in[56]
port 292 nsew default input
rlabel metal2 s 124480 0 124536 800 6 la_data_in[57]
port 293 nsew default input
rlabel metal2 s 125860 0 125916 800 6 la_data_in[58]
port 294 nsew default input
rlabel metal2 s 127148 0 127204 800 6 la_data_in[59]
port 295 nsew default input
rlabel metal2 s 54468 0 54524 800 6 la_data_in[5]
port 296 nsew default input
rlabel metal2 s 128528 0 128584 800 6 la_data_in[60]
port 297 nsew default input
rlabel metal2 s 129908 0 129964 800 6 la_data_in[61]
port 298 nsew default input
rlabel metal2 s 131196 0 131252 800 6 la_data_in[62]
port 299 nsew default input
rlabel metal2 s 132576 0 132632 800 6 la_data_in[63]
port 300 nsew default input
rlabel metal2 s 133956 0 134012 800 6 la_data_in[64]
port 301 nsew default input
rlabel metal2 s 135244 0 135300 800 6 la_data_in[65]
port 302 nsew default input
rlabel metal2 s 136624 0 136680 800 6 la_data_in[66]
port 303 nsew default input
rlabel metal2 s 138004 0 138060 800 6 la_data_in[67]
port 304 nsew default input
rlabel metal2 s 139292 0 139348 800 6 la_data_in[68]
port 305 nsew default input
rlabel metal2 s 140672 0 140728 800 6 la_data_in[69]
port 306 nsew default input
rlabel metal2 s 55848 0 55904 800 6 la_data_in[6]
port 307 nsew default input
rlabel metal2 s 141960 0 142016 800 6 la_data_in[70]
port 308 nsew default input
rlabel metal2 s 143340 0 143396 800 6 la_data_in[71]
port 309 nsew default input
rlabel metal2 s 144720 0 144776 800 6 la_data_in[72]
port 310 nsew default input
rlabel metal2 s 146008 0 146064 800 6 la_data_in[73]
port 311 nsew default input
rlabel metal2 s 147388 0 147444 800 6 la_data_in[74]
port 312 nsew default input
rlabel metal2 s 148768 0 148824 800 6 la_data_in[75]
port 313 nsew default input
rlabel metal2 s 150056 0 150112 800 6 la_data_in[76]
port 314 nsew default input
rlabel metal2 s 151436 0 151492 800 6 la_data_in[77]
port 315 nsew default input
rlabel metal2 s 152816 0 152872 800 6 la_data_in[78]
port 316 nsew default input
rlabel metal2 s 154104 0 154160 800 6 la_data_in[79]
port 317 nsew default input
rlabel metal2 s 57136 0 57192 800 6 la_data_in[7]
port 318 nsew default input
rlabel metal2 s 155484 0 155540 800 6 la_data_in[80]
port 319 nsew default input
rlabel metal2 s 156772 0 156828 800 6 la_data_in[81]
port 320 nsew default input
rlabel metal2 s 158152 0 158208 800 6 la_data_in[82]
port 321 nsew default input
rlabel metal2 s 159532 0 159588 800 6 la_data_in[83]
port 322 nsew default input
rlabel metal2 s 160820 0 160876 800 6 la_data_in[84]
port 323 nsew default input
rlabel metal2 s 162200 0 162256 800 6 la_data_in[85]
port 324 nsew default input
rlabel metal2 s 163580 0 163636 800 6 la_data_in[86]
port 325 nsew default input
rlabel metal2 s 164868 0 164924 800 6 la_data_in[87]
port 326 nsew default input
rlabel metal2 s 166248 0 166304 800 6 la_data_in[88]
port 327 nsew default input
rlabel metal2 s 167628 0 167684 800 6 la_data_in[89]
port 328 nsew default input
rlabel metal2 s 58516 0 58572 800 6 la_data_in[8]
port 329 nsew default input
rlabel metal2 s 168916 0 168972 800 6 la_data_in[90]
port 330 nsew default input
rlabel metal2 s 170296 0 170352 800 6 la_data_in[91]
port 331 nsew default input
rlabel metal2 s 171676 0 171732 800 6 la_data_in[92]
port 332 nsew default input
rlabel metal2 s 172964 0 173020 800 6 la_data_in[93]
port 333 nsew default input
rlabel metal2 s 174344 0 174400 800 6 la_data_in[94]
port 334 nsew default input
rlabel metal2 s 175632 0 175688 800 6 la_data_in[95]
port 335 nsew default input
rlabel metal2 s 177012 0 177068 800 6 la_data_in[96]
port 336 nsew default input
rlabel metal2 s 178392 0 178448 800 6 la_data_in[97]
port 337 nsew default input
rlabel metal2 s 179680 0 179736 800 6 la_data_in[98]
port 338 nsew default input
rlabel metal2 s 181060 0 181116 800 6 la_data_in[99]
port 339 nsew default input
rlabel metal2 s 59804 0 59860 800 6 la_data_in[9]
port 340 nsew default input
rlabel metal2 s 48212 0 48268 800 6 la_data_out[0]
port 341 nsew default output
rlabel metal2 s 182808 0 182864 800 6 la_data_out[100]
port 342 nsew default output
rlabel metal2 s 184188 0 184244 800 6 la_data_out[101]
port 343 nsew default output
rlabel metal2 s 185568 0 185624 800 6 la_data_out[102]
port 344 nsew default output
rlabel metal2 s 186856 0 186912 800 6 la_data_out[103]
port 345 nsew default output
rlabel metal2 s 188236 0 188292 800 6 la_data_out[104]
port 346 nsew default output
rlabel metal2 s 189616 0 189672 800 6 la_data_out[105]
port 347 nsew default output
rlabel metal2 s 190904 0 190960 800 6 la_data_out[106]
port 348 nsew default output
rlabel metal2 s 192284 0 192340 800 6 la_data_out[107]
port 349 nsew default output
rlabel metal2 s 193664 0 193720 800 6 la_data_out[108]
port 350 nsew default output
rlabel metal2 s 194952 0 195008 800 6 la_data_out[109]
port 351 nsew default output
rlabel metal2 s 61644 0 61700 800 6 la_data_out[10]
port 352 nsew default output
rlabel metal2 s 196332 0 196388 800 6 la_data_out[110]
port 353 nsew default output
rlabel metal2 s 197712 0 197768 800 6 la_data_out[111]
port 354 nsew default output
rlabel metal2 s 199000 0 199056 800 6 la_data_out[112]
port 355 nsew default output
rlabel metal2 s 200380 0 200436 800 6 la_data_out[113]
port 356 nsew default output
rlabel metal2 s 201668 0 201724 800 6 la_data_out[114]
port 357 nsew default output
rlabel metal2 s 203048 0 203104 800 6 la_data_out[115]
port 358 nsew default output
rlabel metal2 s 204428 0 204484 800 6 la_data_out[116]
port 359 nsew default output
rlabel metal2 s 205716 0 205772 800 6 la_data_out[117]
port 360 nsew default output
rlabel metal2 s 207096 0 207152 800 6 la_data_out[118]
port 361 nsew default output
rlabel metal2 s 208476 0 208532 800 6 la_data_out[119]
port 362 nsew default output
rlabel metal2 s 63024 0 63080 800 6 la_data_out[11]
port 363 nsew default output
rlabel metal2 s 209764 0 209820 800 6 la_data_out[120]
port 364 nsew default output
rlabel metal2 s 211144 0 211200 800 6 la_data_out[121]
port 365 nsew default output
rlabel metal2 s 212524 0 212580 800 6 la_data_out[122]
port 366 nsew default output
rlabel metal2 s 213812 0 213868 800 6 la_data_out[123]
port 367 nsew default output
rlabel metal2 s 215192 0 215248 800 6 la_data_out[124]
port 368 nsew default output
rlabel metal2 s 216480 0 216536 800 6 la_data_out[125]
port 369 nsew default output
rlabel metal2 s 217860 0 217916 800 6 la_data_out[126]
port 370 nsew default output
rlabel metal2 s 219240 0 219296 800 6 la_data_out[127]
port 371 nsew default output
rlabel metal2 s 64312 0 64368 800 6 la_data_out[12]
port 372 nsew default output
rlabel metal2 s 65692 0 65748 800 6 la_data_out[13]
port 373 nsew default output
rlabel metal2 s 67072 0 67128 800 6 la_data_out[14]
port 374 nsew default output
rlabel metal2 s 68360 0 68416 800 6 la_data_out[15]
port 375 nsew default output
rlabel metal2 s 69740 0 69796 800 6 la_data_out[16]
port 376 nsew default output
rlabel metal2 s 71028 0 71084 800 6 la_data_out[17]
port 377 nsew default output
rlabel metal2 s 72408 0 72464 800 6 la_data_out[18]
port 378 nsew default output
rlabel metal2 s 73788 0 73844 800 6 la_data_out[19]
port 379 nsew default output
rlabel metal2 s 49500 0 49556 800 6 la_data_out[1]
port 380 nsew default output
rlabel metal2 s 75076 0 75132 800 6 la_data_out[20]
port 381 nsew default output
rlabel metal2 s 76456 0 76512 800 6 la_data_out[21]
port 382 nsew default output
rlabel metal2 s 77836 0 77892 800 6 la_data_out[22]
port 383 nsew default output
rlabel metal2 s 79124 0 79180 800 6 la_data_out[23]
port 384 nsew default output
rlabel metal2 s 80504 0 80560 800 6 la_data_out[24]
port 385 nsew default output
rlabel metal2 s 81884 0 81940 800 6 la_data_out[25]
port 386 nsew default output
rlabel metal2 s 83172 0 83228 800 6 la_data_out[26]
port 387 nsew default output
rlabel metal2 s 84552 0 84608 800 6 la_data_out[27]
port 388 nsew default output
rlabel metal2 s 85932 0 85988 800 6 la_data_out[28]
port 389 nsew default output
rlabel metal2 s 87220 0 87276 800 6 la_data_out[29]
port 390 nsew default output
rlabel metal2 s 50880 0 50936 800 6 la_data_out[2]
port 391 nsew default output
rlabel metal2 s 88600 0 88656 800 6 la_data_out[30]
port 392 nsew default output
rlabel metal2 s 89888 0 89944 800 6 la_data_out[31]
port 393 nsew default output
rlabel metal2 s 91268 0 91324 800 6 la_data_out[32]
port 394 nsew default output
rlabel metal2 s 92648 0 92704 800 6 la_data_out[33]
port 395 nsew default output
rlabel metal2 s 93936 0 93992 800 6 la_data_out[34]
port 396 nsew default output
rlabel metal2 s 95316 0 95372 800 6 la_data_out[35]
port 397 nsew default output
rlabel metal2 s 96696 0 96752 800 6 la_data_out[36]
port 398 nsew default output
rlabel metal2 s 97984 0 98040 800 6 la_data_out[37]
port 399 nsew default output
rlabel metal2 s 99364 0 99420 800 6 la_data_out[38]
port 400 nsew default output
rlabel metal2 s 100744 0 100800 800 6 la_data_out[39]
port 401 nsew default output
rlabel metal2 s 52260 0 52316 800 6 la_data_out[3]
port 402 nsew default output
rlabel metal2 s 102032 0 102088 800 6 la_data_out[40]
port 403 nsew default output
rlabel metal2 s 103412 0 103468 800 6 la_data_out[41]
port 404 nsew default output
rlabel metal2 s 104700 0 104756 800 6 la_data_out[42]
port 405 nsew default output
rlabel metal2 s 106080 0 106136 800 6 la_data_out[43]
port 406 nsew default output
rlabel metal2 s 107460 0 107516 800 6 la_data_out[44]
port 407 nsew default output
rlabel metal2 s 108748 0 108804 800 6 la_data_out[45]
port 408 nsew default output
rlabel metal2 s 110128 0 110184 800 6 la_data_out[46]
port 409 nsew default output
rlabel metal2 s 111508 0 111564 800 6 la_data_out[47]
port 410 nsew default output
rlabel metal2 s 112796 0 112852 800 6 la_data_out[48]
port 411 nsew default output
rlabel metal2 s 114176 0 114232 800 6 la_data_out[49]
port 412 nsew default output
rlabel metal2 s 53548 0 53604 800 6 la_data_out[4]
port 413 nsew default output
rlabel metal2 s 115556 0 115612 800 6 la_data_out[50]
port 414 nsew default output
rlabel metal2 s 116844 0 116900 800 6 la_data_out[51]
port 415 nsew default output
rlabel metal2 s 118224 0 118280 800 6 la_data_out[52]
port 416 nsew default output
rlabel metal2 s 119512 0 119568 800 6 la_data_out[53]
port 417 nsew default output
rlabel metal2 s 120892 0 120948 800 6 la_data_out[54]
port 418 nsew default output
rlabel metal2 s 122272 0 122328 800 6 la_data_out[55]
port 419 nsew default output
rlabel metal2 s 123560 0 123616 800 6 la_data_out[56]
port 420 nsew default output
rlabel metal2 s 124940 0 124996 800 6 la_data_out[57]
port 421 nsew default output
rlabel metal2 s 126320 0 126376 800 6 la_data_out[58]
port 422 nsew default output
rlabel metal2 s 127608 0 127664 800 6 la_data_out[59]
port 423 nsew default output
rlabel metal2 s 54928 0 54984 800 6 la_data_out[5]
port 424 nsew default output
rlabel metal2 s 128988 0 129044 800 6 la_data_out[60]
port 425 nsew default output
rlabel metal2 s 130368 0 130424 800 6 la_data_out[61]
port 426 nsew default output
rlabel metal2 s 131656 0 131712 800 6 la_data_out[62]
port 427 nsew default output
rlabel metal2 s 133036 0 133092 800 6 la_data_out[63]
port 428 nsew default output
rlabel metal2 s 134324 0 134380 800 6 la_data_out[64]
port 429 nsew default output
rlabel metal2 s 135704 0 135760 800 6 la_data_out[65]
port 430 nsew default output
rlabel metal2 s 137084 0 137140 800 6 la_data_out[66]
port 431 nsew default output
rlabel metal2 s 138372 0 138428 800 6 la_data_out[67]
port 432 nsew default output
rlabel metal2 s 139752 0 139808 800 6 la_data_out[68]
port 433 nsew default output
rlabel metal2 s 141132 0 141188 800 6 la_data_out[69]
port 434 nsew default output
rlabel metal2 s 56216 0 56272 800 6 la_data_out[6]
port 435 nsew default output
rlabel metal2 s 142420 0 142476 800 6 la_data_out[70]
port 436 nsew default output
rlabel metal2 s 143800 0 143856 800 6 la_data_out[71]
port 437 nsew default output
rlabel metal2 s 145180 0 145236 800 6 la_data_out[72]
port 438 nsew default output
rlabel metal2 s 146468 0 146524 800 6 la_data_out[73]
port 439 nsew default output
rlabel metal2 s 147848 0 147904 800 6 la_data_out[74]
port 440 nsew default output
rlabel metal2 s 149228 0 149284 800 6 la_data_out[75]
port 441 nsew default output
rlabel metal2 s 150516 0 150572 800 6 la_data_out[76]
port 442 nsew default output
rlabel metal2 s 151896 0 151952 800 6 la_data_out[77]
port 443 nsew default output
rlabel metal2 s 153184 0 153240 800 6 la_data_out[78]
port 444 nsew default output
rlabel metal2 s 154564 0 154620 800 6 la_data_out[79]
port 445 nsew default output
rlabel metal2 s 57596 0 57652 800 6 la_data_out[7]
port 446 nsew default output
rlabel metal2 s 155944 0 156000 800 6 la_data_out[80]
port 447 nsew default output
rlabel metal2 s 157232 0 157288 800 6 la_data_out[81]
port 448 nsew default output
rlabel metal2 s 158612 0 158668 800 6 la_data_out[82]
port 449 nsew default output
rlabel metal2 s 159992 0 160048 800 6 la_data_out[83]
port 450 nsew default output
rlabel metal2 s 161280 0 161336 800 6 la_data_out[84]
port 451 nsew default output
rlabel metal2 s 162660 0 162716 800 6 la_data_out[85]
port 452 nsew default output
rlabel metal2 s 164040 0 164096 800 6 la_data_out[86]
port 453 nsew default output
rlabel metal2 s 165328 0 165384 800 6 la_data_out[87]
port 454 nsew default output
rlabel metal2 s 166708 0 166764 800 6 la_data_out[88]
port 455 nsew default output
rlabel metal2 s 167996 0 168052 800 6 la_data_out[89]
port 456 nsew default output
rlabel metal2 s 58976 0 59032 800 6 la_data_out[8]
port 457 nsew default output
rlabel metal2 s 169376 0 169432 800 6 la_data_out[90]
port 458 nsew default output
rlabel metal2 s 170756 0 170812 800 6 la_data_out[91]
port 459 nsew default output
rlabel metal2 s 172044 0 172100 800 6 la_data_out[92]
port 460 nsew default output
rlabel metal2 s 173424 0 173480 800 6 la_data_out[93]
port 461 nsew default output
rlabel metal2 s 174804 0 174860 800 6 la_data_out[94]
port 462 nsew default output
rlabel metal2 s 176092 0 176148 800 6 la_data_out[95]
port 463 nsew default output
rlabel metal2 s 177472 0 177528 800 6 la_data_out[96]
port 464 nsew default output
rlabel metal2 s 178852 0 178908 800 6 la_data_out[97]
port 465 nsew default output
rlabel metal2 s 180140 0 180196 800 6 la_data_out[98]
port 466 nsew default output
rlabel metal2 s 181520 0 181576 800 6 la_data_out[99]
port 467 nsew default output
rlabel metal2 s 60264 0 60320 800 6 la_data_out[9]
port 468 nsew default output
rlabel metal2 s 48580 0 48636 800 6 la_oen[0]
port 469 nsew default input
rlabel metal2 s 183268 0 183324 800 6 la_oen[100]
port 470 nsew default input
rlabel metal2 s 184648 0 184704 800 6 la_oen[101]
port 471 nsew default input
rlabel metal2 s 186028 0 186084 800 6 la_oen[102]
port 472 nsew default input
rlabel metal2 s 187316 0 187372 800 6 la_oen[103]
port 473 nsew default input
rlabel metal2 s 188696 0 188752 800 6 la_oen[104]
port 474 nsew default input
rlabel metal2 s 190076 0 190132 800 6 la_oen[105]
port 475 nsew default input
rlabel metal2 s 191364 0 191420 800 6 la_oen[106]
port 476 nsew default input
rlabel metal2 s 192744 0 192800 800 6 la_oen[107]
port 477 nsew default input
rlabel metal2 s 194032 0 194088 800 6 la_oen[108]
port 478 nsew default input
rlabel metal2 s 195412 0 195468 800 6 la_oen[109]
port 479 nsew default input
rlabel metal2 s 62104 0 62160 800 6 la_oen[10]
port 480 nsew default input
rlabel metal2 s 196792 0 196848 800 6 la_oen[110]
port 481 nsew default input
rlabel metal2 s 198080 0 198136 800 6 la_oen[111]
port 482 nsew default input
rlabel metal2 s 199460 0 199516 800 6 la_oen[112]
port 483 nsew default input
rlabel metal2 s 200840 0 200896 800 6 la_oen[113]
port 484 nsew default input
rlabel metal2 s 202128 0 202184 800 6 la_oen[114]
port 485 nsew default input
rlabel metal2 s 203508 0 203564 800 6 la_oen[115]
port 486 nsew default input
rlabel metal2 s 204888 0 204944 800 6 la_oen[116]
port 487 nsew default input
rlabel metal2 s 206176 0 206232 800 6 la_oen[117]
port 488 nsew default input
rlabel metal2 s 207556 0 207612 800 6 la_oen[118]
port 489 nsew default input
rlabel metal2 s 208936 0 208992 800 6 la_oen[119]
port 490 nsew default input
rlabel metal2 s 63484 0 63540 800 6 la_oen[11]
port 491 nsew default input
rlabel metal2 s 210224 0 210280 800 6 la_oen[120]
port 492 nsew default input
rlabel metal2 s 211604 0 211660 800 6 la_oen[121]
port 493 nsew default input
rlabel metal2 s 212892 0 212948 800 6 la_oen[122]
port 494 nsew default input
rlabel metal2 s 214272 0 214328 800 6 la_oen[123]
port 495 nsew default input
rlabel metal2 s 215652 0 215708 800 6 la_oen[124]
port 496 nsew default input
rlabel metal2 s 216940 0 216996 800 6 la_oen[125]
port 497 nsew default input
rlabel metal2 s 218320 0 218376 800 6 la_oen[126]
port 498 nsew default input
rlabel metal2 s 219700 0 219756 800 6 la_oen[127]
port 499 nsew default input
rlabel metal2 s 64772 0 64828 800 6 la_oen[12]
port 500 nsew default input
rlabel metal2 s 66152 0 66208 800 6 la_oen[13]
port 501 nsew default input
rlabel metal2 s 67440 0 67496 800 6 la_oen[14]
port 502 nsew default input
rlabel metal2 s 68820 0 68876 800 6 la_oen[15]
port 503 nsew default input
rlabel metal2 s 70200 0 70256 800 6 la_oen[16]
port 504 nsew default input
rlabel metal2 s 71488 0 71544 800 6 la_oen[17]
port 505 nsew default input
rlabel metal2 s 72868 0 72924 800 6 la_oen[18]
port 506 nsew default input
rlabel metal2 s 74248 0 74304 800 6 la_oen[19]
port 507 nsew default input
rlabel metal2 s 49960 0 50016 800 6 la_oen[1]
port 508 nsew default input
rlabel metal2 s 75536 0 75592 800 6 la_oen[20]
port 509 nsew default input
rlabel metal2 s 76916 0 76972 800 6 la_oen[21]
port 510 nsew default input
rlabel metal2 s 78296 0 78352 800 6 la_oen[22]
port 511 nsew default input
rlabel metal2 s 79584 0 79640 800 6 la_oen[23]
port 512 nsew default input
rlabel metal2 s 80964 0 81020 800 6 la_oen[24]
port 513 nsew default input
rlabel metal2 s 82252 0 82308 800 6 la_oen[25]
port 514 nsew default input
rlabel metal2 s 83632 0 83688 800 6 la_oen[26]
port 515 nsew default input
rlabel metal2 s 85012 0 85068 800 6 la_oen[27]
port 516 nsew default input
rlabel metal2 s 86300 0 86356 800 6 la_oen[28]
port 517 nsew default input
rlabel metal2 s 87680 0 87736 800 6 la_oen[29]
port 518 nsew default input
rlabel metal2 s 51340 0 51396 800 6 la_oen[2]
port 519 nsew default input
rlabel metal2 s 89060 0 89116 800 6 la_oen[30]
port 520 nsew default input
rlabel metal2 s 90348 0 90404 800 6 la_oen[31]
port 521 nsew default input
rlabel metal2 s 91728 0 91784 800 6 la_oen[32]
port 522 nsew default input
rlabel metal2 s 93108 0 93164 800 6 la_oen[33]
port 523 nsew default input
rlabel metal2 s 94396 0 94452 800 6 la_oen[34]
port 524 nsew default input
rlabel metal2 s 95776 0 95832 800 6 la_oen[35]
port 525 nsew default input
rlabel metal2 s 97064 0 97120 800 6 la_oen[36]
port 526 nsew default input
rlabel metal2 s 98444 0 98500 800 6 la_oen[37]
port 527 nsew default input
rlabel metal2 s 99824 0 99880 800 6 la_oen[38]
port 528 nsew default input
rlabel metal2 s 101112 0 101168 800 6 la_oen[39]
port 529 nsew default input
rlabel metal2 s 52628 0 52684 800 6 la_oen[3]
port 530 nsew default input
rlabel metal2 s 102492 0 102548 800 6 la_oen[40]
port 531 nsew default input
rlabel metal2 s 103872 0 103928 800 6 la_oen[41]
port 532 nsew default input
rlabel metal2 s 105160 0 105216 800 6 la_oen[42]
port 533 nsew default input
rlabel metal2 s 106540 0 106596 800 6 la_oen[43]
port 534 nsew default input
rlabel metal2 s 107920 0 107976 800 6 la_oen[44]
port 535 nsew default input
rlabel metal2 s 109208 0 109264 800 6 la_oen[45]
port 536 nsew default input
rlabel metal2 s 110588 0 110644 800 6 la_oen[46]
port 537 nsew default input
rlabel metal2 s 111968 0 112024 800 6 la_oen[47]
port 538 nsew default input
rlabel metal2 s 113256 0 113312 800 6 la_oen[48]
port 539 nsew default input
rlabel metal2 s 114636 0 114692 800 6 la_oen[49]
port 540 nsew default input
rlabel metal2 s 54008 0 54064 800 6 la_oen[4]
port 541 nsew default input
rlabel metal2 s 115924 0 115980 800 6 la_oen[50]
port 542 nsew default input
rlabel metal2 s 117304 0 117360 800 6 la_oen[51]
port 543 nsew default input
rlabel metal2 s 118684 0 118740 800 6 la_oen[52]
port 544 nsew default input
rlabel metal2 s 119972 0 120028 800 6 la_oen[53]
port 545 nsew default input
rlabel metal2 s 121352 0 121408 800 6 la_oen[54]
port 546 nsew default input
rlabel metal2 s 122732 0 122788 800 6 la_oen[55]
port 547 nsew default input
rlabel metal2 s 124020 0 124076 800 6 la_oen[56]
port 548 nsew default input
rlabel metal2 s 125400 0 125456 800 6 la_oen[57]
port 549 nsew default input
rlabel metal2 s 126780 0 126836 800 6 la_oen[58]
port 550 nsew default input
rlabel metal2 s 128068 0 128124 800 6 la_oen[59]
port 551 nsew default input
rlabel metal2 s 55388 0 55444 800 6 la_oen[5]
port 552 nsew default input
rlabel metal2 s 129448 0 129504 800 6 la_oen[60]
port 553 nsew default input
rlabel metal2 s 130736 0 130792 800 6 la_oen[61]
port 554 nsew default input
rlabel metal2 s 132116 0 132172 800 6 la_oen[62]
port 555 nsew default input
rlabel metal2 s 133496 0 133552 800 6 la_oen[63]
port 556 nsew default input
rlabel metal2 s 134784 0 134840 800 6 la_oen[64]
port 557 nsew default input
rlabel metal2 s 136164 0 136220 800 6 la_oen[65]
port 558 nsew default input
rlabel metal2 s 137544 0 137600 800 6 la_oen[66]
port 559 nsew default input
rlabel metal2 s 138832 0 138888 800 6 la_oen[67]
port 560 nsew default input
rlabel metal2 s 140212 0 140268 800 6 la_oen[68]
port 561 nsew default input
rlabel metal2 s 141592 0 141648 800 6 la_oen[69]
port 562 nsew default input
rlabel metal2 s 56676 0 56732 800 6 la_oen[6]
port 563 nsew default input
rlabel metal2 s 142880 0 142936 800 6 la_oen[70]
port 564 nsew default input
rlabel metal2 s 144260 0 144316 800 6 la_oen[71]
port 565 nsew default input
rlabel metal2 s 145548 0 145604 800 6 la_oen[72]
port 566 nsew default input
rlabel metal2 s 146928 0 146984 800 6 la_oen[73]
port 567 nsew default input
rlabel metal2 s 148308 0 148364 800 6 la_oen[74]
port 568 nsew default input
rlabel metal2 s 149596 0 149652 800 6 la_oen[75]
port 569 nsew default input
rlabel metal2 s 150976 0 151032 800 6 la_oen[76]
port 570 nsew default input
rlabel metal2 s 152356 0 152412 800 6 la_oen[77]
port 571 nsew default input
rlabel metal2 s 153644 0 153700 800 6 la_oen[78]
port 572 nsew default input
rlabel metal2 s 155024 0 155080 800 6 la_oen[79]
port 573 nsew default input
rlabel metal2 s 58056 0 58112 800 6 la_oen[7]
port 574 nsew default input
rlabel metal2 s 156404 0 156460 800 6 la_oen[80]
port 575 nsew default input
rlabel metal2 s 157692 0 157748 800 6 la_oen[81]
port 576 nsew default input
rlabel metal2 s 159072 0 159128 800 6 la_oen[82]
port 577 nsew default input
rlabel metal2 s 160452 0 160508 800 6 la_oen[83]
port 578 nsew default input
rlabel metal2 s 161740 0 161796 800 6 la_oen[84]
port 579 nsew default input
rlabel metal2 s 163120 0 163176 800 6 la_oen[85]
port 580 nsew default input
rlabel metal2 s 164408 0 164464 800 6 la_oen[86]
port 581 nsew default input
rlabel metal2 s 165788 0 165844 800 6 la_oen[87]
port 582 nsew default input
rlabel metal2 s 167168 0 167224 800 6 la_oen[88]
port 583 nsew default input
rlabel metal2 s 168456 0 168512 800 6 la_oen[89]
port 584 nsew default input
rlabel metal2 s 59436 0 59492 800 6 la_oen[8]
port 585 nsew default input
rlabel metal2 s 169836 0 169892 800 6 la_oen[90]
port 586 nsew default input
rlabel metal2 s 171216 0 171272 800 6 la_oen[91]
port 587 nsew default input
rlabel metal2 s 172504 0 172560 800 6 la_oen[92]
port 588 nsew default input
rlabel metal2 s 173884 0 173940 800 6 la_oen[93]
port 589 nsew default input
rlabel metal2 s 175264 0 175320 800 6 la_oen[94]
port 590 nsew default input
rlabel metal2 s 176552 0 176608 800 6 la_oen[95]
port 591 nsew default input
rlabel metal2 s 177932 0 177988 800 6 la_oen[96]
port 592 nsew default input
rlabel metal2 s 179220 0 179276 800 6 la_oen[97]
port 593 nsew default input
rlabel metal2 s 180600 0 180656 800 6 la_oen[98]
port 594 nsew default input
rlabel metal2 s 181980 0 182036 800 6 la_oen[99]
port 595 nsew default input
rlabel metal2 s 60724 0 60780 800 6 la_oen[9]
port 596 nsew default input
rlabel metal3 s 219186 2864 219986 2984 6 one
port 597 nsew default output
rlabel metal2 s 188 0 244 800 6 wb_clk_i
port 598 nsew default input
rlabel metal2 s 556 0 612 800 6 wb_rst_i
port 599 nsew default input
rlabel metal2 s 1016 0 1072 800 6 wbs_ack_o
port 600 nsew default output
rlabel metal2 s 2856 0 2912 800 6 wbs_adr_i[0]
port 601 nsew default input
rlabel metal2 s 18128 0 18184 800 6 wbs_adr_i[10]
port 602 nsew default input
rlabel metal2 s 19416 0 19472 800 6 wbs_adr_i[11]
port 603 nsew default input
rlabel metal2 s 20796 0 20852 800 6 wbs_adr_i[12]
port 604 nsew default input
rlabel metal2 s 22176 0 22232 800 6 wbs_adr_i[13]
port 605 nsew default input
rlabel metal2 s 23464 0 23520 800 6 wbs_adr_i[14]
port 606 nsew default input
rlabel metal2 s 24844 0 24900 800 6 wbs_adr_i[15]
port 607 nsew default input
rlabel metal2 s 26224 0 26280 800 6 wbs_adr_i[16]
port 608 nsew default input
rlabel metal2 s 27512 0 27568 800 6 wbs_adr_i[17]
port 609 nsew default input
rlabel metal2 s 28892 0 28948 800 6 wbs_adr_i[18]
port 610 nsew default input
rlabel metal2 s 30180 0 30236 800 6 wbs_adr_i[19]
port 611 nsew default input
rlabel metal2 s 4604 0 4660 800 6 wbs_adr_i[1]
port 612 nsew default input
rlabel metal2 s 31560 0 31616 800 6 wbs_adr_i[20]
port 613 nsew default input
rlabel metal2 s 32940 0 32996 800 6 wbs_adr_i[21]
port 614 nsew default input
rlabel metal2 s 34228 0 34284 800 6 wbs_adr_i[22]
port 615 nsew default input
rlabel metal2 s 35608 0 35664 800 6 wbs_adr_i[23]
port 616 nsew default input
rlabel metal2 s 36988 0 37044 800 6 wbs_adr_i[24]
port 617 nsew default input
rlabel metal2 s 38276 0 38332 800 6 wbs_adr_i[25]
port 618 nsew default input
rlabel metal2 s 39656 0 39712 800 6 wbs_adr_i[26]
port 619 nsew default input
rlabel metal2 s 41036 0 41092 800 6 wbs_adr_i[27]
port 620 nsew default input
rlabel metal2 s 42324 0 42380 800 6 wbs_adr_i[28]
port 621 nsew default input
rlabel metal2 s 43704 0 43760 800 6 wbs_adr_i[29]
port 622 nsew default input
rlabel metal2 s 6444 0 6500 800 6 wbs_adr_i[2]
port 623 nsew default input
rlabel metal2 s 44992 0 45048 800 6 wbs_adr_i[30]
port 624 nsew default input
rlabel metal2 s 46372 0 46428 800 6 wbs_adr_i[31]
port 625 nsew default input
rlabel metal2 s 8192 0 8248 800 6 wbs_adr_i[3]
port 626 nsew default input
rlabel metal2 s 10032 0 10088 800 6 wbs_adr_i[4]
port 627 nsew default input
rlabel metal2 s 11320 0 11376 800 6 wbs_adr_i[5]
port 628 nsew default input
rlabel metal2 s 12700 0 12756 800 6 wbs_adr_i[6]
port 629 nsew default input
rlabel metal2 s 14080 0 14136 800 6 wbs_adr_i[7]
port 630 nsew default input
rlabel metal2 s 15368 0 15424 800 6 wbs_adr_i[8]
port 631 nsew default input
rlabel metal2 s 16748 0 16804 800 6 wbs_adr_i[9]
port 632 nsew default input
rlabel metal2 s 1476 0 1532 800 6 wbs_cyc_i
port 633 nsew default input
rlabel metal2 s 3316 0 3372 800 6 wbs_dat_i[0]
port 634 nsew default input
rlabel metal2 s 18588 0 18644 800 6 wbs_dat_i[10]
port 635 nsew default input
rlabel metal2 s 19876 0 19932 800 6 wbs_dat_i[11]
port 636 nsew default input
rlabel metal2 s 21256 0 21312 800 6 wbs_dat_i[12]
port 637 nsew default input
rlabel metal2 s 22544 0 22600 800 6 wbs_dat_i[13]
port 638 nsew default input
rlabel metal2 s 23924 0 23980 800 6 wbs_dat_i[14]
port 639 nsew default input
rlabel metal2 s 25304 0 25360 800 6 wbs_dat_i[15]
port 640 nsew default input
rlabel metal2 s 26592 0 26648 800 6 wbs_dat_i[16]
port 641 nsew default input
rlabel metal2 s 27972 0 28028 800 6 wbs_dat_i[17]
port 642 nsew default input
rlabel metal2 s 29352 0 29408 800 6 wbs_dat_i[18]
port 643 nsew default input
rlabel metal2 s 30640 0 30696 800 6 wbs_dat_i[19]
port 644 nsew default input
rlabel metal2 s 5064 0 5120 800 6 wbs_dat_i[1]
port 645 nsew default input
rlabel metal2 s 32020 0 32076 800 6 wbs_dat_i[20]
port 646 nsew default input
rlabel metal2 s 33400 0 33456 800 6 wbs_dat_i[21]
port 647 nsew default input
rlabel metal2 s 34688 0 34744 800 6 wbs_dat_i[22]
port 648 nsew default input
rlabel metal2 s 36068 0 36124 800 6 wbs_dat_i[23]
port 649 nsew default input
rlabel metal2 s 37448 0 37504 800 6 wbs_dat_i[24]
port 650 nsew default input
rlabel metal2 s 38736 0 38792 800 6 wbs_dat_i[25]
port 651 nsew default input
rlabel metal2 s 40116 0 40172 800 6 wbs_dat_i[26]
port 652 nsew default input
rlabel metal2 s 41404 0 41460 800 6 wbs_dat_i[27]
port 653 nsew default input
rlabel metal2 s 42784 0 42840 800 6 wbs_dat_i[28]
port 654 nsew default input
rlabel metal2 s 44164 0 44220 800 6 wbs_dat_i[29]
port 655 nsew default input
rlabel metal2 s 6904 0 6960 800 6 wbs_dat_i[2]
port 656 nsew default input
rlabel metal2 s 45452 0 45508 800 6 wbs_dat_i[30]
port 657 nsew default input
rlabel metal2 s 46832 0 46888 800 6 wbs_dat_i[31]
port 658 nsew default input
rlabel metal2 s 8652 0 8708 800 6 wbs_dat_i[3]
port 659 nsew default input
rlabel metal2 s 10492 0 10548 800 6 wbs_dat_i[4]
port 660 nsew default input
rlabel metal2 s 11780 0 11836 800 6 wbs_dat_i[5]
port 661 nsew default input
rlabel metal2 s 13160 0 13216 800 6 wbs_dat_i[6]
port 662 nsew default input
rlabel metal2 s 14540 0 14596 800 6 wbs_dat_i[7]
port 663 nsew default input
rlabel metal2 s 15828 0 15884 800 6 wbs_dat_i[8]
port 664 nsew default input
rlabel metal2 s 17208 0 17264 800 6 wbs_dat_i[9]
port 665 nsew default input
rlabel metal2 s 3776 0 3832 800 6 wbs_dat_o[0]
port 666 nsew default output
rlabel metal2 s 18956 0 19012 800 6 wbs_dat_o[10]
port 667 nsew default output
rlabel metal2 s 20336 0 20392 800 6 wbs_dat_o[11]
port 668 nsew default output
rlabel metal2 s 21716 0 21772 800 6 wbs_dat_o[12]
port 669 nsew default output
rlabel metal2 s 23004 0 23060 800 6 wbs_dat_o[13]
port 670 nsew default output
rlabel metal2 s 24384 0 24440 800 6 wbs_dat_o[14]
port 671 nsew default output
rlabel metal2 s 25764 0 25820 800 6 wbs_dat_o[15]
port 672 nsew default output
rlabel metal2 s 27052 0 27108 800 6 wbs_dat_o[16]
port 673 nsew default output
rlabel metal2 s 28432 0 28488 800 6 wbs_dat_o[17]
port 674 nsew default output
rlabel metal2 s 29812 0 29868 800 6 wbs_dat_o[18]
port 675 nsew default output
rlabel metal2 s 31100 0 31156 800 6 wbs_dat_o[19]
port 676 nsew default output
rlabel metal2 s 5524 0 5580 800 6 wbs_dat_o[1]
port 677 nsew default output
rlabel metal2 s 32480 0 32536 800 6 wbs_dat_o[20]
port 678 nsew default output
rlabel metal2 s 33768 0 33824 800 6 wbs_dat_o[21]
port 679 nsew default output
rlabel metal2 s 35148 0 35204 800 6 wbs_dat_o[22]
port 680 nsew default output
rlabel metal2 s 36528 0 36584 800 6 wbs_dat_o[23]
port 681 nsew default output
rlabel metal2 s 37816 0 37872 800 6 wbs_dat_o[24]
port 682 nsew default output
rlabel metal2 s 39196 0 39252 800 6 wbs_dat_o[25]
port 683 nsew default output
rlabel metal2 s 40576 0 40632 800 6 wbs_dat_o[26]
port 684 nsew default output
rlabel metal2 s 41864 0 41920 800 6 wbs_dat_o[27]
port 685 nsew default output
rlabel metal2 s 43244 0 43300 800 6 wbs_dat_o[28]
port 686 nsew default output
rlabel metal2 s 44624 0 44680 800 6 wbs_dat_o[29]
port 687 nsew default output
rlabel metal2 s 7364 0 7420 800 6 wbs_dat_o[2]
port 688 nsew default output
rlabel metal2 s 45912 0 45968 800 6 wbs_dat_o[30]
port 689 nsew default output
rlabel metal2 s 47292 0 47348 800 6 wbs_dat_o[31]
port 690 nsew default output
rlabel metal2 s 9112 0 9168 800 6 wbs_dat_o[3]
port 691 nsew default output
rlabel metal2 s 10952 0 11008 800 6 wbs_dat_o[4]
port 692 nsew default output
rlabel metal2 s 12240 0 12296 800 6 wbs_dat_o[5]
port 693 nsew default output
rlabel metal2 s 13620 0 13676 800 6 wbs_dat_o[6]
port 694 nsew default output
rlabel metal2 s 15000 0 15056 800 6 wbs_dat_o[7]
port 695 nsew default output
rlabel metal2 s 16288 0 16344 800 6 wbs_dat_o[8]
port 696 nsew default output
rlabel metal2 s 17668 0 17724 800 6 wbs_dat_o[9]
port 697 nsew default output
rlabel metal2 s 4144 0 4200 800 6 wbs_sel_i[0]
port 698 nsew default input
rlabel metal2 s 5984 0 6040 800 6 wbs_sel_i[1]
port 699 nsew default input
rlabel metal2 s 7732 0 7788 800 6 wbs_sel_i[2]
port 700 nsew default input
rlabel metal2 s 9572 0 9628 800 6 wbs_sel_i[3]
port 701 nsew default input
rlabel metal2 s 1936 0 1992 800 6 wbs_stb_i
port 702 nsew default input
rlabel metal2 s 2396 0 2452 800 6 wbs_we_i
port 703 nsew default input
rlabel metal3 s 219186 960 219986 1080 6 zero
port 704 nsew default output
rlabel metal4 s 4194 2128 4514 217648 6 VPWR
port 705 nsew power input
rlabel metal4 s 19554 2128 19874 217648 6 VGND
port 706 nsew ground input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 219986 220000
string LEFview TRUE
<< end >>
