magic
tech sky130A
magscale 1 2
timestamp 1607539949
<< obsli1 >>
rect 1104 2159 200836 199665
<< obsm1 >>
rect 198 2128 201834 199696
<< metal2 >>
rect 2962 201200 3018 202000
rect 8850 201200 8906 202000
rect 14830 201200 14886 202000
rect 20718 201200 20774 202000
rect 26698 201200 26754 202000
rect 32586 201200 32642 202000
rect 38566 201200 38622 202000
rect 44546 201200 44602 202000
rect 50434 201200 50490 202000
rect 56414 201200 56470 202000
rect 62302 201200 62358 202000
rect 68282 201200 68338 202000
rect 74262 201200 74318 202000
rect 80150 201200 80206 202000
rect 86130 201200 86186 202000
rect 92018 201200 92074 202000
rect 97998 201200 98054 202000
rect 103978 201200 104034 202000
rect 109866 201200 109922 202000
rect 115846 201200 115902 202000
rect 121734 201200 121790 202000
rect 127714 201200 127770 202000
rect 133602 201200 133658 202000
rect 139582 201200 139638 202000
rect 145562 201200 145618 202000
rect 151450 201200 151506 202000
rect 157430 201200 157486 202000
rect 163318 201200 163374 202000
rect 169298 201200 169354 202000
rect 175278 201200 175334 202000
rect 181166 201200 181222 202000
rect 187146 201200 187202 202000
rect 193034 201200 193090 202000
rect 199014 201200 199070 202000
rect 202 0 258 800
rect 570 0 626 800
rect 938 0 994 800
rect 1306 0 1362 800
rect 1674 0 1730 800
rect 2042 0 2098 800
rect 2502 0 2558 800
rect 2870 0 2926 800
rect 3238 0 3294 800
rect 3606 0 3662 800
rect 3974 0 4030 800
rect 4434 0 4490 800
rect 4802 0 4858 800
rect 5170 0 5226 800
rect 5538 0 5594 800
rect 5906 0 5962 800
rect 6366 0 6422 800
rect 6734 0 6790 800
rect 7102 0 7158 800
rect 7470 0 7526 800
rect 7838 0 7894 800
rect 8298 0 8354 800
rect 8666 0 8722 800
rect 9034 0 9090 800
rect 9402 0 9458 800
rect 9770 0 9826 800
rect 10230 0 10286 800
rect 10598 0 10654 800
rect 10966 0 11022 800
rect 11334 0 11390 800
rect 11702 0 11758 800
rect 12162 0 12218 800
rect 12530 0 12586 800
rect 12898 0 12954 800
rect 13266 0 13322 800
rect 13634 0 13690 800
rect 14094 0 14150 800
rect 14462 0 14518 800
rect 14830 0 14886 800
rect 15198 0 15254 800
rect 15566 0 15622 800
rect 16026 0 16082 800
rect 16394 0 16450 800
rect 16762 0 16818 800
rect 17130 0 17186 800
rect 17498 0 17554 800
rect 17958 0 18014 800
rect 18326 0 18382 800
rect 18694 0 18750 800
rect 19062 0 19118 800
rect 19430 0 19486 800
rect 19890 0 19946 800
rect 20258 0 20314 800
rect 20626 0 20682 800
rect 20994 0 21050 800
rect 21362 0 21418 800
rect 21822 0 21878 800
rect 22190 0 22246 800
rect 22558 0 22614 800
rect 22926 0 22982 800
rect 23294 0 23350 800
rect 23754 0 23810 800
rect 24122 0 24178 800
rect 24490 0 24546 800
rect 24858 0 24914 800
rect 25226 0 25282 800
rect 25686 0 25742 800
rect 26054 0 26110 800
rect 26422 0 26478 800
rect 26790 0 26846 800
rect 27158 0 27214 800
rect 27618 0 27674 800
rect 27986 0 28042 800
rect 28354 0 28410 800
rect 28722 0 28778 800
rect 29090 0 29146 800
rect 29550 0 29606 800
rect 29918 0 29974 800
rect 30286 0 30342 800
rect 30654 0 30710 800
rect 31022 0 31078 800
rect 31482 0 31538 800
rect 31850 0 31906 800
rect 32218 0 32274 800
rect 32586 0 32642 800
rect 32954 0 33010 800
rect 33414 0 33470 800
rect 33782 0 33838 800
rect 34150 0 34206 800
rect 34518 0 34574 800
rect 34886 0 34942 800
rect 35346 0 35402 800
rect 35714 0 35770 800
rect 36082 0 36138 800
rect 36450 0 36506 800
rect 36818 0 36874 800
rect 37278 0 37334 800
rect 37646 0 37702 800
rect 38014 0 38070 800
rect 38382 0 38438 800
rect 38750 0 38806 800
rect 39210 0 39266 800
rect 39578 0 39634 800
rect 39946 0 40002 800
rect 40314 0 40370 800
rect 40682 0 40738 800
rect 41142 0 41198 800
rect 41510 0 41566 800
rect 41878 0 41934 800
rect 42246 0 42302 800
rect 42614 0 42670 800
rect 43074 0 43130 800
rect 43442 0 43498 800
rect 43810 0 43866 800
rect 44178 0 44234 800
rect 44546 0 44602 800
rect 45006 0 45062 800
rect 45374 0 45430 800
rect 45742 0 45798 800
rect 46110 0 46166 800
rect 46478 0 46534 800
rect 46938 0 46994 800
rect 47306 0 47362 800
rect 47674 0 47730 800
rect 48042 0 48098 800
rect 48410 0 48466 800
rect 48870 0 48926 800
rect 49238 0 49294 800
rect 49606 0 49662 800
rect 49974 0 50030 800
rect 50342 0 50398 800
rect 50802 0 50858 800
rect 51170 0 51226 800
rect 51538 0 51594 800
rect 51906 0 51962 800
rect 52274 0 52330 800
rect 52734 0 52790 800
rect 53102 0 53158 800
rect 53470 0 53526 800
rect 53838 0 53894 800
rect 54206 0 54262 800
rect 54666 0 54722 800
rect 55034 0 55090 800
rect 55402 0 55458 800
rect 55770 0 55826 800
rect 56138 0 56194 800
rect 56598 0 56654 800
rect 56966 0 57022 800
rect 57334 0 57390 800
rect 57702 0 57758 800
rect 58070 0 58126 800
rect 58530 0 58586 800
rect 58898 0 58954 800
rect 59266 0 59322 800
rect 59634 0 59690 800
rect 60002 0 60058 800
rect 60462 0 60518 800
rect 60830 0 60886 800
rect 61198 0 61254 800
rect 61566 0 61622 800
rect 61934 0 61990 800
rect 62394 0 62450 800
rect 62762 0 62818 800
rect 63130 0 63186 800
rect 63498 0 63554 800
rect 63866 0 63922 800
rect 64326 0 64382 800
rect 64694 0 64750 800
rect 65062 0 65118 800
rect 65430 0 65486 800
rect 65798 0 65854 800
rect 66258 0 66314 800
rect 66626 0 66682 800
rect 66994 0 67050 800
rect 67362 0 67418 800
rect 67730 0 67786 800
rect 68098 0 68154 800
rect 68558 0 68614 800
rect 68926 0 68982 800
rect 69294 0 69350 800
rect 69662 0 69718 800
rect 70030 0 70086 800
rect 70490 0 70546 800
rect 70858 0 70914 800
rect 71226 0 71282 800
rect 71594 0 71650 800
rect 71962 0 72018 800
rect 72422 0 72478 800
rect 72790 0 72846 800
rect 73158 0 73214 800
rect 73526 0 73582 800
rect 73894 0 73950 800
rect 74354 0 74410 800
rect 74722 0 74778 800
rect 75090 0 75146 800
rect 75458 0 75514 800
rect 75826 0 75882 800
rect 76286 0 76342 800
rect 76654 0 76710 800
rect 77022 0 77078 800
rect 77390 0 77446 800
rect 77758 0 77814 800
rect 78218 0 78274 800
rect 78586 0 78642 800
rect 78954 0 79010 800
rect 79322 0 79378 800
rect 79690 0 79746 800
rect 80150 0 80206 800
rect 80518 0 80574 800
rect 80886 0 80942 800
rect 81254 0 81310 800
rect 81622 0 81678 800
rect 82082 0 82138 800
rect 82450 0 82506 800
rect 82818 0 82874 800
rect 83186 0 83242 800
rect 83554 0 83610 800
rect 84014 0 84070 800
rect 84382 0 84438 800
rect 84750 0 84806 800
rect 85118 0 85174 800
rect 85486 0 85542 800
rect 85946 0 86002 800
rect 86314 0 86370 800
rect 86682 0 86738 800
rect 87050 0 87106 800
rect 87418 0 87474 800
rect 87878 0 87934 800
rect 88246 0 88302 800
rect 88614 0 88670 800
rect 88982 0 89038 800
rect 89350 0 89406 800
rect 89810 0 89866 800
rect 90178 0 90234 800
rect 90546 0 90602 800
rect 90914 0 90970 800
rect 91282 0 91338 800
rect 91742 0 91798 800
rect 92110 0 92166 800
rect 92478 0 92534 800
rect 92846 0 92902 800
rect 93214 0 93270 800
rect 93674 0 93730 800
rect 94042 0 94098 800
rect 94410 0 94466 800
rect 94778 0 94834 800
rect 95146 0 95202 800
rect 95606 0 95662 800
rect 95974 0 96030 800
rect 96342 0 96398 800
rect 96710 0 96766 800
rect 97078 0 97134 800
rect 97538 0 97594 800
rect 97906 0 97962 800
rect 98274 0 98330 800
rect 98642 0 98698 800
rect 99010 0 99066 800
rect 99470 0 99526 800
rect 99838 0 99894 800
rect 100206 0 100262 800
rect 100574 0 100630 800
rect 100942 0 100998 800
rect 101402 0 101458 800
rect 101770 0 101826 800
rect 102138 0 102194 800
rect 102506 0 102562 800
rect 102874 0 102930 800
rect 103334 0 103390 800
rect 103702 0 103758 800
rect 104070 0 104126 800
rect 104438 0 104494 800
rect 104806 0 104862 800
rect 105266 0 105322 800
rect 105634 0 105690 800
rect 106002 0 106058 800
rect 106370 0 106426 800
rect 106738 0 106794 800
rect 107198 0 107254 800
rect 107566 0 107622 800
rect 107934 0 107990 800
rect 108302 0 108358 800
rect 108670 0 108726 800
rect 109130 0 109186 800
rect 109498 0 109554 800
rect 109866 0 109922 800
rect 110234 0 110290 800
rect 110602 0 110658 800
rect 111062 0 111118 800
rect 111430 0 111486 800
rect 111798 0 111854 800
rect 112166 0 112222 800
rect 112534 0 112590 800
rect 112994 0 113050 800
rect 113362 0 113418 800
rect 113730 0 113786 800
rect 114098 0 114154 800
rect 114466 0 114522 800
rect 114926 0 114982 800
rect 115294 0 115350 800
rect 115662 0 115718 800
rect 116030 0 116086 800
rect 116398 0 116454 800
rect 116858 0 116914 800
rect 117226 0 117282 800
rect 117594 0 117650 800
rect 117962 0 118018 800
rect 118330 0 118386 800
rect 118790 0 118846 800
rect 119158 0 119214 800
rect 119526 0 119582 800
rect 119894 0 119950 800
rect 120262 0 120318 800
rect 120722 0 120778 800
rect 121090 0 121146 800
rect 121458 0 121514 800
rect 121826 0 121882 800
rect 122194 0 122250 800
rect 122654 0 122710 800
rect 123022 0 123078 800
rect 123390 0 123446 800
rect 123758 0 123814 800
rect 124126 0 124182 800
rect 124586 0 124642 800
rect 124954 0 125010 800
rect 125322 0 125378 800
rect 125690 0 125746 800
rect 126058 0 126114 800
rect 126518 0 126574 800
rect 126886 0 126942 800
rect 127254 0 127310 800
rect 127622 0 127678 800
rect 127990 0 128046 800
rect 128450 0 128506 800
rect 128818 0 128874 800
rect 129186 0 129242 800
rect 129554 0 129610 800
rect 129922 0 129978 800
rect 130382 0 130438 800
rect 130750 0 130806 800
rect 131118 0 131174 800
rect 131486 0 131542 800
rect 131854 0 131910 800
rect 132314 0 132370 800
rect 132682 0 132738 800
rect 133050 0 133106 800
rect 133418 0 133474 800
rect 133786 0 133842 800
rect 134246 0 134302 800
rect 134614 0 134670 800
rect 134982 0 135038 800
rect 135350 0 135406 800
rect 135718 0 135774 800
rect 136086 0 136142 800
rect 136546 0 136602 800
rect 136914 0 136970 800
rect 137282 0 137338 800
rect 137650 0 137706 800
rect 138018 0 138074 800
rect 138478 0 138534 800
rect 138846 0 138902 800
rect 139214 0 139270 800
rect 139582 0 139638 800
rect 139950 0 140006 800
rect 140410 0 140466 800
rect 140778 0 140834 800
rect 141146 0 141202 800
rect 141514 0 141570 800
rect 141882 0 141938 800
rect 142342 0 142398 800
rect 142710 0 142766 800
rect 143078 0 143134 800
rect 143446 0 143502 800
rect 143814 0 143870 800
rect 144274 0 144330 800
rect 144642 0 144698 800
rect 145010 0 145066 800
rect 145378 0 145434 800
rect 145746 0 145802 800
rect 146206 0 146262 800
rect 146574 0 146630 800
rect 146942 0 146998 800
rect 147310 0 147366 800
rect 147678 0 147734 800
rect 148138 0 148194 800
rect 148506 0 148562 800
rect 148874 0 148930 800
rect 149242 0 149298 800
rect 149610 0 149666 800
rect 150070 0 150126 800
rect 150438 0 150494 800
rect 150806 0 150862 800
rect 151174 0 151230 800
rect 151542 0 151598 800
rect 152002 0 152058 800
rect 152370 0 152426 800
rect 152738 0 152794 800
rect 153106 0 153162 800
rect 153474 0 153530 800
rect 153934 0 153990 800
rect 154302 0 154358 800
rect 154670 0 154726 800
rect 155038 0 155094 800
rect 155406 0 155462 800
rect 155866 0 155922 800
rect 156234 0 156290 800
rect 156602 0 156658 800
rect 156970 0 157026 800
rect 157338 0 157394 800
rect 157798 0 157854 800
rect 158166 0 158222 800
rect 158534 0 158590 800
rect 158902 0 158958 800
rect 159270 0 159326 800
rect 159730 0 159786 800
rect 160098 0 160154 800
rect 160466 0 160522 800
rect 160834 0 160890 800
rect 161202 0 161258 800
rect 161662 0 161718 800
rect 162030 0 162086 800
rect 162398 0 162454 800
rect 162766 0 162822 800
rect 163134 0 163190 800
rect 163594 0 163650 800
rect 163962 0 164018 800
rect 164330 0 164386 800
rect 164698 0 164754 800
rect 165066 0 165122 800
rect 165526 0 165582 800
rect 165894 0 165950 800
rect 166262 0 166318 800
rect 166630 0 166686 800
rect 166998 0 167054 800
rect 167458 0 167514 800
rect 167826 0 167882 800
rect 168194 0 168250 800
rect 168562 0 168618 800
rect 168930 0 168986 800
rect 169390 0 169446 800
rect 169758 0 169814 800
rect 170126 0 170182 800
rect 170494 0 170550 800
rect 170862 0 170918 800
rect 171322 0 171378 800
rect 171690 0 171746 800
rect 172058 0 172114 800
rect 172426 0 172482 800
rect 172794 0 172850 800
rect 173254 0 173310 800
rect 173622 0 173678 800
rect 173990 0 174046 800
rect 174358 0 174414 800
rect 174726 0 174782 800
rect 175186 0 175242 800
rect 175554 0 175610 800
rect 175922 0 175978 800
rect 176290 0 176346 800
rect 176658 0 176714 800
rect 177118 0 177174 800
rect 177486 0 177542 800
rect 177854 0 177910 800
rect 178222 0 178278 800
rect 178590 0 178646 800
rect 179050 0 179106 800
rect 179418 0 179474 800
rect 179786 0 179842 800
rect 180154 0 180210 800
rect 180522 0 180578 800
rect 180982 0 181038 800
rect 181350 0 181406 800
rect 181718 0 181774 800
rect 182086 0 182142 800
rect 182454 0 182510 800
rect 182914 0 182970 800
rect 183282 0 183338 800
rect 183650 0 183706 800
rect 184018 0 184074 800
rect 184386 0 184442 800
rect 184846 0 184902 800
rect 185214 0 185270 800
rect 185582 0 185638 800
rect 185950 0 186006 800
rect 186318 0 186374 800
rect 186778 0 186834 800
rect 187146 0 187202 800
rect 187514 0 187570 800
rect 187882 0 187938 800
rect 188250 0 188306 800
rect 188710 0 188766 800
rect 189078 0 189134 800
rect 189446 0 189502 800
rect 189814 0 189870 800
rect 190182 0 190238 800
rect 190642 0 190698 800
rect 191010 0 191066 800
rect 191378 0 191434 800
rect 191746 0 191802 800
rect 192114 0 192170 800
rect 192574 0 192630 800
rect 192942 0 192998 800
rect 193310 0 193366 800
rect 193678 0 193734 800
rect 194046 0 194102 800
rect 194506 0 194562 800
rect 194874 0 194930 800
rect 195242 0 195298 800
rect 195610 0 195666 800
rect 195978 0 196034 800
rect 196438 0 196494 800
rect 196806 0 196862 800
rect 197174 0 197230 800
rect 197542 0 197598 800
rect 197910 0 197966 800
rect 198370 0 198426 800
rect 198738 0 198794 800
rect 199106 0 199162 800
rect 199474 0 199530 800
rect 199842 0 199898 800
rect 200302 0 200358 800
rect 200670 0 200726 800
rect 201038 0 201094 800
rect 201406 0 201462 800
rect 201774 0 201830 800
<< obsm2 >>
rect 204 201144 2906 201200
rect 3074 201144 8794 201200
rect 8962 201144 14774 201200
rect 14942 201144 20662 201200
rect 20830 201144 26642 201200
rect 26810 201144 32530 201200
rect 32698 201144 38510 201200
rect 38678 201144 44490 201200
rect 44658 201144 50378 201200
rect 50546 201144 56358 201200
rect 56526 201144 62246 201200
rect 62414 201144 68226 201200
rect 68394 201144 74206 201200
rect 74374 201144 80094 201200
rect 80262 201144 86074 201200
rect 86242 201144 91962 201200
rect 92130 201144 97942 201200
rect 98110 201144 103922 201200
rect 104090 201144 109810 201200
rect 109978 201144 115790 201200
rect 115958 201144 121678 201200
rect 121846 201144 127658 201200
rect 127826 201144 133546 201200
rect 133714 201144 139526 201200
rect 139694 201144 145506 201200
rect 145674 201144 151394 201200
rect 151562 201144 157374 201200
rect 157542 201144 163262 201200
rect 163430 201144 169242 201200
rect 169410 201144 175222 201200
rect 175390 201144 181110 201200
rect 181278 201144 187090 201200
rect 187258 201144 192978 201200
rect 193146 201144 198958 201200
rect 199126 201144 201828 201200
rect 204 856 201828 201144
rect 314 800 514 856
rect 682 800 882 856
rect 1050 800 1250 856
rect 1418 800 1618 856
rect 1786 800 1986 856
rect 2154 800 2446 856
rect 2614 800 2814 856
rect 2982 800 3182 856
rect 3350 800 3550 856
rect 3718 800 3918 856
rect 4086 800 4378 856
rect 4546 800 4746 856
rect 4914 800 5114 856
rect 5282 800 5482 856
rect 5650 800 5850 856
rect 6018 800 6310 856
rect 6478 800 6678 856
rect 6846 800 7046 856
rect 7214 800 7414 856
rect 7582 800 7782 856
rect 7950 800 8242 856
rect 8410 800 8610 856
rect 8778 800 8978 856
rect 9146 800 9346 856
rect 9514 800 9714 856
rect 9882 800 10174 856
rect 10342 800 10542 856
rect 10710 800 10910 856
rect 11078 800 11278 856
rect 11446 800 11646 856
rect 11814 800 12106 856
rect 12274 800 12474 856
rect 12642 800 12842 856
rect 13010 800 13210 856
rect 13378 800 13578 856
rect 13746 800 14038 856
rect 14206 800 14406 856
rect 14574 800 14774 856
rect 14942 800 15142 856
rect 15310 800 15510 856
rect 15678 800 15970 856
rect 16138 800 16338 856
rect 16506 800 16706 856
rect 16874 800 17074 856
rect 17242 800 17442 856
rect 17610 800 17902 856
rect 18070 800 18270 856
rect 18438 800 18638 856
rect 18806 800 19006 856
rect 19174 800 19374 856
rect 19542 800 19834 856
rect 20002 800 20202 856
rect 20370 800 20570 856
rect 20738 800 20938 856
rect 21106 800 21306 856
rect 21474 800 21766 856
rect 21934 800 22134 856
rect 22302 800 22502 856
rect 22670 800 22870 856
rect 23038 800 23238 856
rect 23406 800 23698 856
rect 23866 800 24066 856
rect 24234 800 24434 856
rect 24602 800 24802 856
rect 24970 800 25170 856
rect 25338 800 25630 856
rect 25798 800 25998 856
rect 26166 800 26366 856
rect 26534 800 26734 856
rect 26902 800 27102 856
rect 27270 800 27562 856
rect 27730 800 27930 856
rect 28098 800 28298 856
rect 28466 800 28666 856
rect 28834 800 29034 856
rect 29202 800 29494 856
rect 29662 800 29862 856
rect 30030 800 30230 856
rect 30398 800 30598 856
rect 30766 800 30966 856
rect 31134 800 31426 856
rect 31594 800 31794 856
rect 31962 800 32162 856
rect 32330 800 32530 856
rect 32698 800 32898 856
rect 33066 800 33358 856
rect 33526 800 33726 856
rect 33894 800 34094 856
rect 34262 800 34462 856
rect 34630 800 34830 856
rect 34998 800 35290 856
rect 35458 800 35658 856
rect 35826 800 36026 856
rect 36194 800 36394 856
rect 36562 800 36762 856
rect 36930 800 37222 856
rect 37390 800 37590 856
rect 37758 800 37958 856
rect 38126 800 38326 856
rect 38494 800 38694 856
rect 38862 800 39154 856
rect 39322 800 39522 856
rect 39690 800 39890 856
rect 40058 800 40258 856
rect 40426 800 40626 856
rect 40794 800 41086 856
rect 41254 800 41454 856
rect 41622 800 41822 856
rect 41990 800 42190 856
rect 42358 800 42558 856
rect 42726 800 43018 856
rect 43186 800 43386 856
rect 43554 800 43754 856
rect 43922 800 44122 856
rect 44290 800 44490 856
rect 44658 800 44950 856
rect 45118 800 45318 856
rect 45486 800 45686 856
rect 45854 800 46054 856
rect 46222 800 46422 856
rect 46590 800 46882 856
rect 47050 800 47250 856
rect 47418 800 47618 856
rect 47786 800 47986 856
rect 48154 800 48354 856
rect 48522 800 48814 856
rect 48982 800 49182 856
rect 49350 800 49550 856
rect 49718 800 49918 856
rect 50086 800 50286 856
rect 50454 800 50746 856
rect 50914 800 51114 856
rect 51282 800 51482 856
rect 51650 800 51850 856
rect 52018 800 52218 856
rect 52386 800 52678 856
rect 52846 800 53046 856
rect 53214 800 53414 856
rect 53582 800 53782 856
rect 53950 800 54150 856
rect 54318 800 54610 856
rect 54778 800 54978 856
rect 55146 800 55346 856
rect 55514 800 55714 856
rect 55882 800 56082 856
rect 56250 800 56542 856
rect 56710 800 56910 856
rect 57078 800 57278 856
rect 57446 800 57646 856
rect 57814 800 58014 856
rect 58182 800 58474 856
rect 58642 800 58842 856
rect 59010 800 59210 856
rect 59378 800 59578 856
rect 59746 800 59946 856
rect 60114 800 60406 856
rect 60574 800 60774 856
rect 60942 800 61142 856
rect 61310 800 61510 856
rect 61678 800 61878 856
rect 62046 800 62338 856
rect 62506 800 62706 856
rect 62874 800 63074 856
rect 63242 800 63442 856
rect 63610 800 63810 856
rect 63978 800 64270 856
rect 64438 800 64638 856
rect 64806 800 65006 856
rect 65174 800 65374 856
rect 65542 800 65742 856
rect 65910 800 66202 856
rect 66370 800 66570 856
rect 66738 800 66938 856
rect 67106 800 67306 856
rect 67474 800 67674 856
rect 67842 800 68042 856
rect 68210 800 68502 856
rect 68670 800 68870 856
rect 69038 800 69238 856
rect 69406 800 69606 856
rect 69774 800 69974 856
rect 70142 800 70434 856
rect 70602 800 70802 856
rect 70970 800 71170 856
rect 71338 800 71538 856
rect 71706 800 71906 856
rect 72074 800 72366 856
rect 72534 800 72734 856
rect 72902 800 73102 856
rect 73270 800 73470 856
rect 73638 800 73838 856
rect 74006 800 74298 856
rect 74466 800 74666 856
rect 74834 800 75034 856
rect 75202 800 75402 856
rect 75570 800 75770 856
rect 75938 800 76230 856
rect 76398 800 76598 856
rect 76766 800 76966 856
rect 77134 800 77334 856
rect 77502 800 77702 856
rect 77870 800 78162 856
rect 78330 800 78530 856
rect 78698 800 78898 856
rect 79066 800 79266 856
rect 79434 800 79634 856
rect 79802 800 80094 856
rect 80262 800 80462 856
rect 80630 800 80830 856
rect 80998 800 81198 856
rect 81366 800 81566 856
rect 81734 800 82026 856
rect 82194 800 82394 856
rect 82562 800 82762 856
rect 82930 800 83130 856
rect 83298 800 83498 856
rect 83666 800 83958 856
rect 84126 800 84326 856
rect 84494 800 84694 856
rect 84862 800 85062 856
rect 85230 800 85430 856
rect 85598 800 85890 856
rect 86058 800 86258 856
rect 86426 800 86626 856
rect 86794 800 86994 856
rect 87162 800 87362 856
rect 87530 800 87822 856
rect 87990 800 88190 856
rect 88358 800 88558 856
rect 88726 800 88926 856
rect 89094 800 89294 856
rect 89462 800 89754 856
rect 89922 800 90122 856
rect 90290 800 90490 856
rect 90658 800 90858 856
rect 91026 800 91226 856
rect 91394 800 91686 856
rect 91854 800 92054 856
rect 92222 800 92422 856
rect 92590 800 92790 856
rect 92958 800 93158 856
rect 93326 800 93618 856
rect 93786 800 93986 856
rect 94154 800 94354 856
rect 94522 800 94722 856
rect 94890 800 95090 856
rect 95258 800 95550 856
rect 95718 800 95918 856
rect 96086 800 96286 856
rect 96454 800 96654 856
rect 96822 800 97022 856
rect 97190 800 97482 856
rect 97650 800 97850 856
rect 98018 800 98218 856
rect 98386 800 98586 856
rect 98754 800 98954 856
rect 99122 800 99414 856
rect 99582 800 99782 856
rect 99950 800 100150 856
rect 100318 800 100518 856
rect 100686 800 100886 856
rect 101054 800 101346 856
rect 101514 800 101714 856
rect 101882 800 102082 856
rect 102250 800 102450 856
rect 102618 800 102818 856
rect 102986 800 103278 856
rect 103446 800 103646 856
rect 103814 800 104014 856
rect 104182 800 104382 856
rect 104550 800 104750 856
rect 104918 800 105210 856
rect 105378 800 105578 856
rect 105746 800 105946 856
rect 106114 800 106314 856
rect 106482 800 106682 856
rect 106850 800 107142 856
rect 107310 800 107510 856
rect 107678 800 107878 856
rect 108046 800 108246 856
rect 108414 800 108614 856
rect 108782 800 109074 856
rect 109242 800 109442 856
rect 109610 800 109810 856
rect 109978 800 110178 856
rect 110346 800 110546 856
rect 110714 800 111006 856
rect 111174 800 111374 856
rect 111542 800 111742 856
rect 111910 800 112110 856
rect 112278 800 112478 856
rect 112646 800 112938 856
rect 113106 800 113306 856
rect 113474 800 113674 856
rect 113842 800 114042 856
rect 114210 800 114410 856
rect 114578 800 114870 856
rect 115038 800 115238 856
rect 115406 800 115606 856
rect 115774 800 115974 856
rect 116142 800 116342 856
rect 116510 800 116802 856
rect 116970 800 117170 856
rect 117338 800 117538 856
rect 117706 800 117906 856
rect 118074 800 118274 856
rect 118442 800 118734 856
rect 118902 800 119102 856
rect 119270 800 119470 856
rect 119638 800 119838 856
rect 120006 800 120206 856
rect 120374 800 120666 856
rect 120834 800 121034 856
rect 121202 800 121402 856
rect 121570 800 121770 856
rect 121938 800 122138 856
rect 122306 800 122598 856
rect 122766 800 122966 856
rect 123134 800 123334 856
rect 123502 800 123702 856
rect 123870 800 124070 856
rect 124238 800 124530 856
rect 124698 800 124898 856
rect 125066 800 125266 856
rect 125434 800 125634 856
rect 125802 800 126002 856
rect 126170 800 126462 856
rect 126630 800 126830 856
rect 126998 800 127198 856
rect 127366 800 127566 856
rect 127734 800 127934 856
rect 128102 800 128394 856
rect 128562 800 128762 856
rect 128930 800 129130 856
rect 129298 800 129498 856
rect 129666 800 129866 856
rect 130034 800 130326 856
rect 130494 800 130694 856
rect 130862 800 131062 856
rect 131230 800 131430 856
rect 131598 800 131798 856
rect 131966 800 132258 856
rect 132426 800 132626 856
rect 132794 800 132994 856
rect 133162 800 133362 856
rect 133530 800 133730 856
rect 133898 800 134190 856
rect 134358 800 134558 856
rect 134726 800 134926 856
rect 135094 800 135294 856
rect 135462 800 135662 856
rect 135830 800 136030 856
rect 136198 800 136490 856
rect 136658 800 136858 856
rect 137026 800 137226 856
rect 137394 800 137594 856
rect 137762 800 137962 856
rect 138130 800 138422 856
rect 138590 800 138790 856
rect 138958 800 139158 856
rect 139326 800 139526 856
rect 139694 800 139894 856
rect 140062 800 140354 856
rect 140522 800 140722 856
rect 140890 800 141090 856
rect 141258 800 141458 856
rect 141626 800 141826 856
rect 141994 800 142286 856
rect 142454 800 142654 856
rect 142822 800 143022 856
rect 143190 800 143390 856
rect 143558 800 143758 856
rect 143926 800 144218 856
rect 144386 800 144586 856
rect 144754 800 144954 856
rect 145122 800 145322 856
rect 145490 800 145690 856
rect 145858 800 146150 856
rect 146318 800 146518 856
rect 146686 800 146886 856
rect 147054 800 147254 856
rect 147422 800 147622 856
rect 147790 800 148082 856
rect 148250 800 148450 856
rect 148618 800 148818 856
rect 148986 800 149186 856
rect 149354 800 149554 856
rect 149722 800 150014 856
rect 150182 800 150382 856
rect 150550 800 150750 856
rect 150918 800 151118 856
rect 151286 800 151486 856
rect 151654 800 151946 856
rect 152114 800 152314 856
rect 152482 800 152682 856
rect 152850 800 153050 856
rect 153218 800 153418 856
rect 153586 800 153878 856
rect 154046 800 154246 856
rect 154414 800 154614 856
rect 154782 800 154982 856
rect 155150 800 155350 856
rect 155518 800 155810 856
rect 155978 800 156178 856
rect 156346 800 156546 856
rect 156714 800 156914 856
rect 157082 800 157282 856
rect 157450 800 157742 856
rect 157910 800 158110 856
rect 158278 800 158478 856
rect 158646 800 158846 856
rect 159014 800 159214 856
rect 159382 800 159674 856
rect 159842 800 160042 856
rect 160210 800 160410 856
rect 160578 800 160778 856
rect 160946 800 161146 856
rect 161314 800 161606 856
rect 161774 800 161974 856
rect 162142 800 162342 856
rect 162510 800 162710 856
rect 162878 800 163078 856
rect 163246 800 163538 856
rect 163706 800 163906 856
rect 164074 800 164274 856
rect 164442 800 164642 856
rect 164810 800 165010 856
rect 165178 800 165470 856
rect 165638 800 165838 856
rect 166006 800 166206 856
rect 166374 800 166574 856
rect 166742 800 166942 856
rect 167110 800 167402 856
rect 167570 800 167770 856
rect 167938 800 168138 856
rect 168306 800 168506 856
rect 168674 800 168874 856
rect 169042 800 169334 856
rect 169502 800 169702 856
rect 169870 800 170070 856
rect 170238 800 170438 856
rect 170606 800 170806 856
rect 170974 800 171266 856
rect 171434 800 171634 856
rect 171802 800 172002 856
rect 172170 800 172370 856
rect 172538 800 172738 856
rect 172906 800 173198 856
rect 173366 800 173566 856
rect 173734 800 173934 856
rect 174102 800 174302 856
rect 174470 800 174670 856
rect 174838 800 175130 856
rect 175298 800 175498 856
rect 175666 800 175866 856
rect 176034 800 176234 856
rect 176402 800 176602 856
rect 176770 800 177062 856
rect 177230 800 177430 856
rect 177598 800 177798 856
rect 177966 800 178166 856
rect 178334 800 178534 856
rect 178702 800 178994 856
rect 179162 800 179362 856
rect 179530 800 179730 856
rect 179898 800 180098 856
rect 180266 800 180466 856
rect 180634 800 180926 856
rect 181094 800 181294 856
rect 181462 800 181662 856
rect 181830 800 182030 856
rect 182198 800 182398 856
rect 182566 800 182858 856
rect 183026 800 183226 856
rect 183394 800 183594 856
rect 183762 800 183962 856
rect 184130 800 184330 856
rect 184498 800 184790 856
rect 184958 800 185158 856
rect 185326 800 185526 856
rect 185694 800 185894 856
rect 186062 800 186262 856
rect 186430 800 186722 856
rect 186890 800 187090 856
rect 187258 800 187458 856
rect 187626 800 187826 856
rect 187994 800 188194 856
rect 188362 800 188654 856
rect 188822 800 189022 856
rect 189190 800 189390 856
rect 189558 800 189758 856
rect 189926 800 190126 856
rect 190294 800 190586 856
rect 190754 800 190954 856
rect 191122 800 191322 856
rect 191490 800 191690 856
rect 191858 800 192058 856
rect 192226 800 192518 856
rect 192686 800 192886 856
rect 193054 800 193254 856
rect 193422 800 193622 856
rect 193790 800 193990 856
rect 194158 800 194450 856
rect 194618 800 194818 856
rect 194986 800 195186 856
rect 195354 800 195554 856
rect 195722 800 195922 856
rect 196090 800 196382 856
rect 196550 800 196750 856
rect 196918 800 197118 856
rect 197286 800 197486 856
rect 197654 800 197854 856
rect 198022 800 198314 856
rect 198482 800 198682 856
rect 198850 800 199050 856
rect 199218 800 199418 856
rect 199586 800 199786 856
rect 199954 800 200246 856
rect 200414 800 200614 856
rect 200782 800 200982 856
rect 201150 800 201350 856
rect 201518 800 201718 856
<< metal3 >>
rect 0 197888 800 198008
rect 201200 197480 202000 197600
rect 0 190136 800 190256
rect 201200 188640 202000 188760
rect 0 182384 800 182504
rect 201200 179936 202000 180056
rect 0 174632 800 174752
rect 201200 171096 202000 171216
rect 0 166880 800 167000
rect 201200 162392 202000 162512
rect 0 159128 800 159248
rect 201200 153552 202000 153672
rect 0 151376 800 151496
rect 201200 144848 202000 144968
rect 0 143624 800 143744
rect 201200 136008 202000 136128
rect 0 135736 800 135856
rect 0 127984 800 128104
rect 201200 127168 202000 127288
rect 0 120232 800 120352
rect 201200 118464 202000 118584
rect 0 112480 800 112600
rect 201200 109624 202000 109744
rect 0 104728 800 104848
rect 201200 100920 202000 101040
rect 0 96976 800 97096
rect 201200 92080 202000 92200
rect 0 89224 800 89344
rect 201200 83376 202000 83496
rect 0 81472 800 81592
rect 201200 74536 202000 74656
rect 0 73720 800 73840
rect 0 65832 800 65952
rect 201200 65696 202000 65816
rect 0 58080 800 58200
rect 201200 56992 202000 57112
rect 0 50328 800 50448
rect 201200 48152 202000 48272
rect 0 42576 800 42696
rect 201200 39448 202000 39568
rect 0 34824 800 34944
rect 201200 30608 202000 30728
rect 0 27072 800 27192
rect 201200 21904 202000 22024
rect 0 19320 800 19440
rect 201200 13064 202000 13184
rect 0 11568 800 11688
rect 201200 4360 202000 4480
rect 0 3816 800 3936
<< obsm3 >>
rect 798 198088 201200 199681
rect 880 197808 201200 198088
rect 798 197680 201200 197808
rect 798 197400 201120 197680
rect 798 190336 201200 197400
rect 880 190056 201200 190336
rect 798 188840 201200 190056
rect 798 188560 201120 188840
rect 798 182584 201200 188560
rect 880 182304 201200 182584
rect 798 180136 201200 182304
rect 798 179856 201120 180136
rect 798 174832 201200 179856
rect 880 174552 201200 174832
rect 798 171296 201200 174552
rect 798 171016 201120 171296
rect 798 167080 201200 171016
rect 880 166800 201200 167080
rect 798 162592 201200 166800
rect 798 162312 201120 162592
rect 798 159328 201200 162312
rect 880 159048 201200 159328
rect 798 153752 201200 159048
rect 798 153472 201120 153752
rect 798 151576 201200 153472
rect 880 151296 201200 151576
rect 798 145048 201200 151296
rect 798 144768 201120 145048
rect 798 143824 201200 144768
rect 880 143544 201200 143824
rect 798 136208 201200 143544
rect 798 135936 201120 136208
rect 880 135928 201120 135936
rect 880 135656 201200 135928
rect 798 128184 201200 135656
rect 880 127904 201200 128184
rect 798 127368 201200 127904
rect 798 127088 201120 127368
rect 798 120432 201200 127088
rect 880 120152 201200 120432
rect 798 118664 201200 120152
rect 798 118384 201120 118664
rect 798 112680 201200 118384
rect 880 112400 201200 112680
rect 798 109824 201200 112400
rect 798 109544 201120 109824
rect 798 104928 201200 109544
rect 880 104648 201200 104928
rect 798 101120 201200 104648
rect 798 100840 201120 101120
rect 798 97176 201200 100840
rect 880 96896 201200 97176
rect 798 92280 201200 96896
rect 798 92000 201120 92280
rect 798 89424 201200 92000
rect 880 89144 201200 89424
rect 798 83576 201200 89144
rect 798 83296 201120 83576
rect 798 81672 201200 83296
rect 880 81392 201200 81672
rect 798 74736 201200 81392
rect 798 74456 201120 74736
rect 798 73920 201200 74456
rect 880 73640 201200 73920
rect 798 66032 201200 73640
rect 880 65896 201200 66032
rect 880 65752 201120 65896
rect 798 65616 201120 65752
rect 798 58280 201200 65616
rect 880 58000 201200 58280
rect 798 57192 201200 58000
rect 798 56912 201120 57192
rect 798 50528 201200 56912
rect 880 50248 201200 50528
rect 798 48352 201200 50248
rect 798 48072 201120 48352
rect 798 42776 201200 48072
rect 880 42496 201200 42776
rect 798 39648 201200 42496
rect 798 39368 201120 39648
rect 798 35024 201200 39368
rect 880 34744 201200 35024
rect 798 30808 201200 34744
rect 798 30528 201120 30808
rect 798 27272 201200 30528
rect 880 26992 201200 27272
rect 798 22104 201200 26992
rect 798 21824 201120 22104
rect 798 19520 201200 21824
rect 880 19240 201200 19520
rect 798 13264 201200 19240
rect 798 12984 201120 13264
rect 798 11768 201200 12984
rect 880 11488 201200 11768
rect 798 4560 201200 11488
rect 798 4280 201120 4560
rect 798 4016 201200 4280
rect 880 3736 201200 4016
rect 798 851 201200 3736
<< metal4 >>
rect 4208 2128 4528 199696
rect 19568 2128 19888 199696
<< obsm4 >>
rect 3739 2128 4128 199696
rect 4608 2128 19488 199696
rect 19968 2128 198661 199696
<< labels >>
rlabel metal2 s 2962 201200 3018 202000 6 cpu_addr_e[0]
port 1 nsew default output
rlabel metal3 s 0 104728 800 104848 6 cpu_addr_e[10]
port 2 nsew default output
rlabel metal2 s 197542 0 197598 800 6 cpu_addr_e[11]
port 3 nsew default output
rlabel metal2 s 198370 0 198426 800 6 cpu_addr_e[12]
port 4 nsew default output
rlabel metal2 s 187146 201200 187202 202000 6 cpu_addr_e[13]
port 5 nsew default output
rlabel metal3 s 0 166880 800 167000 6 cpu_addr_e[14]
port 6 nsew default output
rlabel metal2 s 200670 0 200726 800 6 cpu_addr_e[15]
port 7 nsew default output
rlabel metal3 s 201200 21904 202000 22024 6 cpu_addr_e[1]
port 8 nsew default output
rlabel metal3 s 0 42576 800 42696 6 cpu_addr_e[2]
port 9 nsew default output
rlabel metal2 s 44546 201200 44602 202000 6 cpu_addr_e[3]
port 10 nsew default output
rlabel metal2 s 62302 201200 62358 202000 6 cpu_addr_e[4]
port 11 nsew default output
rlabel metal2 s 193310 0 193366 800 6 cpu_addr_e[5]
port 12 nsew default output
rlabel metal3 s 0 73720 800 73840 6 cpu_addr_e[6]
port 13 nsew default output
rlabel metal3 s 201200 109624 202000 109744 6 cpu_addr_e[7]
port 14 nsew default output
rlabel metal2 s 145562 201200 145618 202000 6 cpu_addr_e[8]
port 15 nsew default output
rlabel metal3 s 201200 162392 202000 162512 6 cpu_addr_e[9]
port 16 nsew default output
rlabel metal2 s 8850 201200 8906 202000 6 cpu_addr_n[0]
port 17 nsew default output
rlabel metal2 s 157430 201200 157486 202000 6 cpu_addr_n[10]
port 18 nsew default output
rlabel metal2 s 169298 201200 169354 202000 6 cpu_addr_n[11]
port 19 nsew default output
rlabel metal3 s 0 143624 800 143744 6 cpu_addr_n[12]
port 20 nsew default output
rlabel metal2 s 199474 0 199530 800 6 cpu_addr_n[13]
port 21 nsew default output
rlabel metal3 s 201200 188640 202000 188760 6 cpu_addr_n[14]
port 22 nsew default output
rlabel metal2 s 201038 0 201094 800 6 cpu_addr_n[15]
port 23 nsew default output
rlabel metal2 s 26698 201200 26754 202000 6 cpu_addr_n[1]
port 24 nsew default output
rlabel metal3 s 201200 56992 202000 57112 6 cpu_addr_n[2]
port 25 nsew default output
rlabel metal2 s 191378 0 191434 800 6 cpu_addr_n[3]
port 26 nsew default output
rlabel metal2 s 68282 201200 68338 202000 6 cpu_addr_n[4]
port 27 nsew default output
rlabel metal2 s 86130 201200 86186 202000 6 cpu_addr_n[5]
port 28 nsew default output
rlabel metal2 s 115846 201200 115902 202000 6 cpu_addr_n[6]
port 29 nsew default output
rlabel metal2 s 194874 0 194930 800 6 cpu_addr_n[7]
port 30 nsew default output
rlabel metal3 s 201200 127168 202000 127288 6 cpu_addr_n[8]
port 31 nsew default output
rlabel metal3 s 201200 171096 202000 171216 6 cpu_addr_n[9]
port 32 nsew default output
rlabel metal3 s 0 3816 800 3936 6 cpu_dtr_e[0]
port 33 nsew default input
rlabel metal2 s 163318 201200 163374 202000 6 cpu_dtr_e[10]
port 34 nsew default input
rlabel metal2 s 175278 201200 175334 202000 6 cpu_dtr_e[11]
port 35 nsew default input
rlabel metal3 s 0 151376 800 151496 6 cpu_dtr_e[12]
port 36 nsew default input
rlabel metal2 s 199842 0 199898 800 6 cpu_dtr_e[13]
port 37 nsew default input
rlabel metal2 s 199014 201200 199070 202000 6 cpu_dtr_e[14]
port 38 nsew default input
rlabel metal2 s 201406 0 201462 800 6 cpu_dtr_e[15]
port 39 nsew default input
rlabel metal2 s 189814 0 189870 800 6 cpu_dtr_e[1]
port 40 nsew default input
rlabel metal2 s 190182 0 190238 800 6 cpu_dtr_e[2]
port 41 nsew default input
rlabel metal2 s 191746 0 191802 800 6 cpu_dtr_e[3]
port 42 nsew default input
rlabel metal2 s 192574 0 192630 800 6 cpu_dtr_e[4]
port 43 nsew default input
rlabel metal2 s 92018 201200 92074 202000 6 cpu_dtr_e[5]
port 44 nsew default input
rlabel metal3 s 201200 100920 202000 101040 6 cpu_dtr_e[6]
port 45 nsew default input
rlabel metal2 s 195242 0 195298 800 6 cpu_dtr_e[7]
port 46 nsew default input
rlabel metal3 s 201200 136008 202000 136128 6 cpu_dtr_e[8]
port 47 nsew default input
rlabel metal2 s 196438 0 196494 800 6 cpu_dtr_e[9]
port 48 nsew default input
rlabel metal2 s 189446 0 189502 800 6 cpu_dtr_n[0]
port 49 nsew default input
rlabel metal3 s 0 112480 800 112600 6 cpu_dtr_n[10]
port 50 nsew default input
rlabel metal3 s 0 135736 800 135856 6 cpu_dtr_n[11]
port 51 nsew default input
rlabel metal3 s 201200 179936 202000 180056 6 cpu_dtr_n[12]
port 52 nsew default input
rlabel metal3 s 0 159128 800 159248 6 cpu_dtr_n[13]
port 53 nsew default input
rlabel metal3 s 0 174632 800 174752 6 cpu_dtr_n[14]
port 54 nsew default input
rlabel metal2 s 201774 0 201830 800 6 cpu_dtr_n[15]
port 55 nsew default input
rlabel metal3 s 201200 30608 202000 30728 6 cpu_dtr_n[1]
port 56 nsew default input
rlabel metal3 s 201200 65696 202000 65816 6 cpu_dtr_n[2]
port 57 nsew default input
rlabel metal2 s 192114 0 192170 800 6 cpu_dtr_n[3]
port 58 nsew default input
rlabel metal3 s 201200 92080 202000 92200 6 cpu_dtr_n[4]
port 59 nsew default input
rlabel metal2 s 97998 201200 98054 202000 6 cpu_dtr_n[5]
port 60 nsew default input
rlabel metal3 s 0 81472 800 81592 6 cpu_dtr_n[6]
port 61 nsew default input
rlabel metal3 s 201200 118464 202000 118584 6 cpu_dtr_n[7]
port 62 nsew default input
rlabel metal2 s 151450 201200 151506 202000 6 cpu_dtr_n[8]
port 63 nsew default input
rlabel metal2 s 196806 0 196862 800 6 cpu_dtr_n[9]
port 64 nsew default input
rlabel metal2 s 14830 201200 14886 202000 6 cpu_dtw_e[0]
port 65 nsew default output
rlabel metal3 s 0 120232 800 120352 6 cpu_dtw_e[10]
port 66 nsew default output
rlabel metal2 s 197910 0 197966 800 6 cpu_dtw_e[11]
port 67 nsew default output
rlabel metal2 s 198738 0 198794 800 6 cpu_dtw_e[12]
port 68 nsew default output
rlabel metal2 s 200302 0 200358 800 6 cpu_dtw_e[13]
port 69 nsew default output
rlabel metal3 s 0 182384 800 182504 6 cpu_dtw_e[14]
port 70 nsew default output
rlabel metal3 s 0 197888 800 198008 6 cpu_dtw_e[15]
port 71 nsew default output
rlabel metal3 s 201200 39448 202000 39568 6 cpu_dtw_e[1]
port 72 nsew default output
rlabel metal2 s 190642 0 190698 800 6 cpu_dtw_e[2]
port 73 nsew default output
rlabel metal3 s 0 50328 800 50448 6 cpu_dtw_e[3]
port 74 nsew default output
rlabel metal2 s 74262 201200 74318 202000 6 cpu_dtw_e[4]
port 75 nsew default output
rlabel metal2 s 193678 0 193734 800 6 cpu_dtw_e[5]
port 76 nsew default output
rlabel metal2 s 194506 0 194562 800 6 cpu_dtw_e[6]
port 77 nsew default output
rlabel metal2 s 195610 0 195666 800 6 cpu_dtw_e[7]
port 78 nsew default output
rlabel metal3 s 201200 144848 202000 144968 6 cpu_dtw_e[8]
port 79 nsew default output
rlabel metal2 s 197174 0 197230 800 6 cpu_dtw_e[9]
port 80 nsew default output
rlabel metal3 s 201200 4360 202000 4480 6 cpu_dtw_n[0]
port 81 nsew default output
rlabel metal3 s 0 127984 800 128104 6 cpu_dtw_n[10]
port 82 nsew default output
rlabel metal2 s 181166 201200 181222 202000 6 cpu_dtw_n[11]
port 83 nsew default output
rlabel metal2 s 199106 0 199162 800 6 cpu_dtw_n[12]
port 84 nsew default output
rlabel metal2 s 193034 201200 193090 202000 6 cpu_dtw_n[13]
port 85 nsew default output
rlabel metal3 s 0 190136 800 190256 6 cpu_dtw_n[14]
port 86 nsew default output
rlabel metal3 s 201200 197480 202000 197600 6 cpu_dtw_n[15]
port 87 nsew default output
rlabel metal2 s 32586 201200 32642 202000 6 cpu_dtw_n[1]
port 88 nsew default output
rlabel metal2 s 191010 0 191066 800 6 cpu_dtw_n[2]
port 89 nsew default output
rlabel metal3 s 0 58080 800 58200 6 cpu_dtw_n[3]
port 90 nsew default output
rlabel metal2 s 80150 201200 80206 202000 6 cpu_dtw_n[4]
port 91 nsew default output
rlabel metal2 s 194046 0 194102 800 6 cpu_dtw_n[5]
port 92 nsew default output
rlabel metal2 s 121734 201200 121790 202000 6 cpu_dtw_n[6]
port 93 nsew default output
rlabel metal2 s 133602 201200 133658 202000 6 cpu_dtw_n[7]
port 94 nsew default output
rlabel metal3 s 201200 153552 202000 153672 6 cpu_dtw_n[8]
port 95 nsew default output
rlabel metal3 s 0 96976 800 97096 6 cpu_dtw_n[9]
port 96 nsew default output
rlabel metal3 s 0 11568 800 11688 6 cpu_mask_e[0]
port 97 nsew default output
rlabel metal2 s 38566 201200 38622 202000 6 cpu_mask_e[1]
port 98 nsew default output
rlabel metal3 s 201200 74536 202000 74656 6 cpu_mask_e[2]
port 99 nsew default output
rlabel metal2 s 50434 201200 50490 202000 6 cpu_mask_e[3]
port 100 nsew default output
rlabel metal3 s 0 65832 800 65952 6 cpu_mask_e[4]
port 101 nsew default output
rlabel metal2 s 103978 201200 104034 202000 6 cpu_mask_e[5]
port 102 nsew default output
rlabel metal3 s 0 89224 800 89344 6 cpu_mask_e[6]
port 103 nsew default output
rlabel metal2 s 139582 201200 139638 202000 6 cpu_mask_e[7]
port 104 nsew default output
rlabel metal3 s 201200 13064 202000 13184 6 cpu_mask_n[0]
port 105 nsew default output
rlabel metal3 s 201200 48152 202000 48272 6 cpu_mask_n[1]
port 106 nsew default output
rlabel metal3 s 201200 83376 202000 83496 6 cpu_mask_n[2]
port 107 nsew default output
rlabel metal2 s 56414 201200 56470 202000 6 cpu_mask_n[3]
port 108 nsew default output
rlabel metal2 s 192942 0 192998 800 6 cpu_mask_n[4]
port 109 nsew default output
rlabel metal2 s 109866 201200 109922 202000 6 cpu_mask_n[5]
port 110 nsew default output
rlabel metal2 s 127714 201200 127770 202000 6 cpu_mask_n[6]
port 111 nsew default output
rlabel metal2 s 195978 0 196034 800 6 cpu_mask_n[7]
port 112 nsew default output
rlabel metal2 s 20718 201200 20774 202000 6 cpu_wen_e[0]
port 113 nsew default output
rlabel metal3 s 0 27072 800 27192 6 cpu_wen_e[1]
port 114 nsew default output
rlabel metal3 s 0 19320 800 19440 6 cpu_wen_n[0]
port 115 nsew default output
rlabel metal3 s 0 34824 800 34944 6 cpu_wen_n[1]
port 116 nsew default output
rlabel metal2 s 41142 0 41198 800 6 la_data_in[0]
port 117 nsew default input
rlabel metal2 s 156970 0 157026 800 6 la_data_in[100]
port 118 nsew default input
rlabel metal2 s 158166 0 158222 800 6 la_data_in[101]
port 119 nsew default input
rlabel metal2 s 159270 0 159326 800 6 la_data_in[102]
port 120 nsew default input
rlabel metal2 s 160466 0 160522 800 6 la_data_in[103]
port 121 nsew default input
rlabel metal2 s 161662 0 161718 800 6 la_data_in[104]
port 122 nsew default input
rlabel metal2 s 162766 0 162822 800 6 la_data_in[105]
port 123 nsew default input
rlabel metal2 s 163962 0 164018 800 6 la_data_in[106]
port 124 nsew default input
rlabel metal2 s 165066 0 165122 800 6 la_data_in[107]
port 125 nsew default input
rlabel metal2 s 166262 0 166318 800 6 la_data_in[108]
port 126 nsew default input
rlabel metal2 s 167458 0 167514 800 6 la_data_in[109]
port 127 nsew default input
rlabel metal2 s 52734 0 52790 800 6 la_data_in[10]
port 128 nsew default input
rlabel metal2 s 168562 0 168618 800 6 la_data_in[110]
port 129 nsew default input
rlabel metal2 s 169758 0 169814 800 6 la_data_in[111]
port 130 nsew default input
rlabel metal2 s 170862 0 170918 800 6 la_data_in[112]
port 131 nsew default input
rlabel metal2 s 172058 0 172114 800 6 la_data_in[113]
port 132 nsew default input
rlabel metal2 s 173254 0 173310 800 6 la_data_in[114]
port 133 nsew default input
rlabel metal2 s 174358 0 174414 800 6 la_data_in[115]
port 134 nsew default input
rlabel metal2 s 175554 0 175610 800 6 la_data_in[116]
port 135 nsew default input
rlabel metal2 s 176658 0 176714 800 6 la_data_in[117]
port 136 nsew default input
rlabel metal2 s 177854 0 177910 800 6 la_data_in[118]
port 137 nsew default input
rlabel metal2 s 179050 0 179106 800 6 la_data_in[119]
port 138 nsew default input
rlabel metal2 s 53838 0 53894 800 6 la_data_in[11]
port 139 nsew default input
rlabel metal2 s 180154 0 180210 800 6 la_data_in[120]
port 140 nsew default input
rlabel metal2 s 181350 0 181406 800 6 la_data_in[121]
port 141 nsew default input
rlabel metal2 s 182454 0 182510 800 6 la_data_in[122]
port 142 nsew default input
rlabel metal2 s 183650 0 183706 800 6 la_data_in[123]
port 143 nsew default input
rlabel metal2 s 184846 0 184902 800 6 la_data_in[124]
port 144 nsew default input
rlabel metal2 s 185950 0 186006 800 6 la_data_in[125]
port 145 nsew default input
rlabel metal2 s 187146 0 187202 800 6 la_data_in[126]
port 146 nsew default input
rlabel metal2 s 188250 0 188306 800 6 la_data_in[127]
port 147 nsew default input
rlabel metal2 s 55034 0 55090 800 6 la_data_in[12]
port 148 nsew default input
rlabel metal2 s 56138 0 56194 800 6 la_data_in[13]
port 149 nsew default input
rlabel metal2 s 57334 0 57390 800 6 la_data_in[14]
port 150 nsew default input
rlabel metal2 s 58530 0 58586 800 6 la_data_in[15]
port 151 nsew default input
rlabel metal2 s 59634 0 59690 800 6 la_data_in[16]
port 152 nsew default input
rlabel metal2 s 60830 0 60886 800 6 la_data_in[17]
port 153 nsew default input
rlabel metal2 s 61934 0 61990 800 6 la_data_in[18]
port 154 nsew default input
rlabel metal2 s 63130 0 63186 800 6 la_data_in[19]
port 155 nsew default input
rlabel metal2 s 42246 0 42302 800 6 la_data_in[1]
port 156 nsew default input
rlabel metal2 s 64326 0 64382 800 6 la_data_in[20]
port 157 nsew default input
rlabel metal2 s 65430 0 65486 800 6 la_data_in[21]
port 158 nsew default input
rlabel metal2 s 66626 0 66682 800 6 la_data_in[22]
port 159 nsew default input
rlabel metal2 s 67730 0 67786 800 6 la_data_in[23]
port 160 nsew default input
rlabel metal2 s 68926 0 68982 800 6 la_data_in[24]
port 161 nsew default input
rlabel metal2 s 70030 0 70086 800 6 la_data_in[25]
port 162 nsew default input
rlabel metal2 s 71226 0 71282 800 6 la_data_in[26]
port 163 nsew default input
rlabel metal2 s 72422 0 72478 800 6 la_data_in[27]
port 164 nsew default input
rlabel metal2 s 73526 0 73582 800 6 la_data_in[28]
port 165 nsew default input
rlabel metal2 s 74722 0 74778 800 6 la_data_in[29]
port 166 nsew default input
rlabel metal2 s 43442 0 43498 800 6 la_data_in[2]
port 167 nsew default input
rlabel metal2 s 75826 0 75882 800 6 la_data_in[30]
port 168 nsew default input
rlabel metal2 s 77022 0 77078 800 6 la_data_in[31]
port 169 nsew default input
rlabel metal2 s 78218 0 78274 800 6 la_data_in[32]
port 170 nsew default input
rlabel metal2 s 79322 0 79378 800 6 la_data_in[33]
port 171 nsew default input
rlabel metal2 s 80518 0 80574 800 6 la_data_in[34]
port 172 nsew default input
rlabel metal2 s 81622 0 81678 800 6 la_data_in[35]
port 173 nsew default input
rlabel metal2 s 82818 0 82874 800 6 la_data_in[36]
port 174 nsew default input
rlabel metal2 s 84014 0 84070 800 6 la_data_in[37]
port 175 nsew default input
rlabel metal2 s 85118 0 85174 800 6 la_data_in[38]
port 176 nsew default input
rlabel metal2 s 86314 0 86370 800 6 la_data_in[39]
port 177 nsew default input
rlabel metal2 s 44546 0 44602 800 6 la_data_in[3]
port 178 nsew default input
rlabel metal2 s 87418 0 87474 800 6 la_data_in[40]
port 179 nsew default input
rlabel metal2 s 88614 0 88670 800 6 la_data_in[41]
port 180 nsew default input
rlabel metal2 s 89810 0 89866 800 6 la_data_in[42]
port 181 nsew default input
rlabel metal2 s 90914 0 90970 800 6 la_data_in[43]
port 182 nsew default input
rlabel metal2 s 92110 0 92166 800 6 la_data_in[44]
port 183 nsew default input
rlabel metal2 s 93214 0 93270 800 6 la_data_in[45]
port 184 nsew default input
rlabel metal2 s 94410 0 94466 800 6 la_data_in[46]
port 185 nsew default input
rlabel metal2 s 95606 0 95662 800 6 la_data_in[47]
port 186 nsew default input
rlabel metal2 s 96710 0 96766 800 6 la_data_in[48]
port 187 nsew default input
rlabel metal2 s 97906 0 97962 800 6 la_data_in[49]
port 188 nsew default input
rlabel metal2 s 45742 0 45798 800 6 la_data_in[4]
port 189 nsew default input
rlabel metal2 s 99010 0 99066 800 6 la_data_in[50]
port 190 nsew default input
rlabel metal2 s 100206 0 100262 800 6 la_data_in[51]
port 191 nsew default input
rlabel metal2 s 101402 0 101458 800 6 la_data_in[52]
port 192 nsew default input
rlabel metal2 s 102506 0 102562 800 6 la_data_in[53]
port 193 nsew default input
rlabel metal2 s 103702 0 103758 800 6 la_data_in[54]
port 194 nsew default input
rlabel metal2 s 104806 0 104862 800 6 la_data_in[55]
port 195 nsew default input
rlabel metal2 s 106002 0 106058 800 6 la_data_in[56]
port 196 nsew default input
rlabel metal2 s 107198 0 107254 800 6 la_data_in[57]
port 197 nsew default input
rlabel metal2 s 108302 0 108358 800 6 la_data_in[58]
port 198 nsew default input
rlabel metal2 s 109498 0 109554 800 6 la_data_in[59]
port 199 nsew default input
rlabel metal2 s 46938 0 46994 800 6 la_data_in[5]
port 200 nsew default input
rlabel metal2 s 110602 0 110658 800 6 la_data_in[60]
port 201 nsew default input
rlabel metal2 s 111798 0 111854 800 6 la_data_in[61]
port 202 nsew default input
rlabel metal2 s 112994 0 113050 800 6 la_data_in[62]
port 203 nsew default input
rlabel metal2 s 114098 0 114154 800 6 la_data_in[63]
port 204 nsew default input
rlabel metal2 s 115294 0 115350 800 6 la_data_in[64]
port 205 nsew default input
rlabel metal2 s 116398 0 116454 800 6 la_data_in[65]
port 206 nsew default input
rlabel metal2 s 117594 0 117650 800 6 la_data_in[66]
port 207 nsew default input
rlabel metal2 s 118790 0 118846 800 6 la_data_in[67]
port 208 nsew default input
rlabel metal2 s 119894 0 119950 800 6 la_data_in[68]
port 209 nsew default input
rlabel metal2 s 121090 0 121146 800 6 la_data_in[69]
port 210 nsew default input
rlabel metal2 s 48042 0 48098 800 6 la_data_in[6]
port 211 nsew default input
rlabel metal2 s 122194 0 122250 800 6 la_data_in[70]
port 212 nsew default input
rlabel metal2 s 123390 0 123446 800 6 la_data_in[71]
port 213 nsew default input
rlabel metal2 s 124586 0 124642 800 6 la_data_in[72]
port 214 nsew default input
rlabel metal2 s 125690 0 125746 800 6 la_data_in[73]
port 215 nsew default input
rlabel metal2 s 126886 0 126942 800 6 la_data_in[74]
port 216 nsew default input
rlabel metal2 s 127990 0 128046 800 6 la_data_in[75]
port 217 nsew default input
rlabel metal2 s 129186 0 129242 800 6 la_data_in[76]
port 218 nsew default input
rlabel metal2 s 130382 0 130438 800 6 la_data_in[77]
port 219 nsew default input
rlabel metal2 s 131486 0 131542 800 6 la_data_in[78]
port 220 nsew default input
rlabel metal2 s 132682 0 132738 800 6 la_data_in[79]
port 221 nsew default input
rlabel metal2 s 49238 0 49294 800 6 la_data_in[7]
port 222 nsew default input
rlabel metal2 s 133786 0 133842 800 6 la_data_in[80]
port 223 nsew default input
rlabel metal2 s 134982 0 135038 800 6 la_data_in[81]
port 224 nsew default input
rlabel metal2 s 136086 0 136142 800 6 la_data_in[82]
port 225 nsew default input
rlabel metal2 s 137282 0 137338 800 6 la_data_in[83]
port 226 nsew default input
rlabel metal2 s 138478 0 138534 800 6 la_data_in[84]
port 227 nsew default input
rlabel metal2 s 139582 0 139638 800 6 la_data_in[85]
port 228 nsew default input
rlabel metal2 s 140778 0 140834 800 6 la_data_in[86]
port 229 nsew default input
rlabel metal2 s 141882 0 141938 800 6 la_data_in[87]
port 230 nsew default input
rlabel metal2 s 143078 0 143134 800 6 la_data_in[88]
port 231 nsew default input
rlabel metal2 s 144274 0 144330 800 6 la_data_in[89]
port 232 nsew default input
rlabel metal2 s 50342 0 50398 800 6 la_data_in[8]
port 233 nsew default input
rlabel metal2 s 145378 0 145434 800 6 la_data_in[90]
port 234 nsew default input
rlabel metal2 s 146574 0 146630 800 6 la_data_in[91]
port 235 nsew default input
rlabel metal2 s 147678 0 147734 800 6 la_data_in[92]
port 236 nsew default input
rlabel metal2 s 148874 0 148930 800 6 la_data_in[93]
port 237 nsew default input
rlabel metal2 s 150070 0 150126 800 6 la_data_in[94]
port 238 nsew default input
rlabel metal2 s 151174 0 151230 800 6 la_data_in[95]
port 239 nsew default input
rlabel metal2 s 152370 0 152426 800 6 la_data_in[96]
port 240 nsew default input
rlabel metal2 s 153474 0 153530 800 6 la_data_in[97]
port 241 nsew default input
rlabel metal2 s 154670 0 154726 800 6 la_data_in[98]
port 242 nsew default input
rlabel metal2 s 155866 0 155922 800 6 la_data_in[99]
port 243 nsew default input
rlabel metal2 s 51538 0 51594 800 6 la_data_in[9]
port 244 nsew default input
rlabel metal2 s 41510 0 41566 800 6 la_data_out[0]
port 245 nsew default output
rlabel metal2 s 157338 0 157394 800 6 la_data_out[100]
port 246 nsew default output
rlabel metal2 s 158534 0 158590 800 6 la_data_out[101]
port 247 nsew default output
rlabel metal2 s 159730 0 159786 800 6 la_data_out[102]
port 248 nsew default output
rlabel metal2 s 160834 0 160890 800 6 la_data_out[103]
port 249 nsew default output
rlabel metal2 s 162030 0 162086 800 6 la_data_out[104]
port 250 nsew default output
rlabel metal2 s 163134 0 163190 800 6 la_data_out[105]
port 251 nsew default output
rlabel metal2 s 164330 0 164386 800 6 la_data_out[106]
port 252 nsew default output
rlabel metal2 s 165526 0 165582 800 6 la_data_out[107]
port 253 nsew default output
rlabel metal2 s 166630 0 166686 800 6 la_data_out[108]
port 254 nsew default output
rlabel metal2 s 167826 0 167882 800 6 la_data_out[109]
port 255 nsew default output
rlabel metal2 s 53102 0 53158 800 6 la_data_out[10]
port 256 nsew default output
rlabel metal2 s 168930 0 168986 800 6 la_data_out[110]
port 257 nsew default output
rlabel metal2 s 170126 0 170182 800 6 la_data_out[111]
port 258 nsew default output
rlabel metal2 s 171322 0 171378 800 6 la_data_out[112]
port 259 nsew default output
rlabel metal2 s 172426 0 172482 800 6 la_data_out[113]
port 260 nsew default output
rlabel metal2 s 173622 0 173678 800 6 la_data_out[114]
port 261 nsew default output
rlabel metal2 s 174726 0 174782 800 6 la_data_out[115]
port 262 nsew default output
rlabel metal2 s 175922 0 175978 800 6 la_data_out[116]
port 263 nsew default output
rlabel metal2 s 177118 0 177174 800 6 la_data_out[117]
port 264 nsew default output
rlabel metal2 s 178222 0 178278 800 6 la_data_out[118]
port 265 nsew default output
rlabel metal2 s 179418 0 179474 800 6 la_data_out[119]
port 266 nsew default output
rlabel metal2 s 54206 0 54262 800 6 la_data_out[11]
port 267 nsew default output
rlabel metal2 s 180522 0 180578 800 6 la_data_out[120]
port 268 nsew default output
rlabel metal2 s 181718 0 181774 800 6 la_data_out[121]
port 269 nsew default output
rlabel metal2 s 182914 0 182970 800 6 la_data_out[122]
port 270 nsew default output
rlabel metal2 s 184018 0 184074 800 6 la_data_out[123]
port 271 nsew default output
rlabel metal2 s 185214 0 185270 800 6 la_data_out[124]
port 272 nsew default output
rlabel metal2 s 186318 0 186374 800 6 la_data_out[125]
port 273 nsew default output
rlabel metal2 s 187514 0 187570 800 6 la_data_out[126]
port 274 nsew default output
rlabel metal2 s 188710 0 188766 800 6 la_data_out[127]
port 275 nsew default output
rlabel metal2 s 55402 0 55458 800 6 la_data_out[12]
port 276 nsew default output
rlabel metal2 s 56598 0 56654 800 6 la_data_out[13]
port 277 nsew default output
rlabel metal2 s 57702 0 57758 800 6 la_data_out[14]
port 278 nsew default output
rlabel metal2 s 58898 0 58954 800 6 la_data_out[15]
port 279 nsew default output
rlabel metal2 s 60002 0 60058 800 6 la_data_out[16]
port 280 nsew default output
rlabel metal2 s 61198 0 61254 800 6 la_data_out[17]
port 281 nsew default output
rlabel metal2 s 62394 0 62450 800 6 la_data_out[18]
port 282 nsew default output
rlabel metal2 s 63498 0 63554 800 6 la_data_out[19]
port 283 nsew default output
rlabel metal2 s 42614 0 42670 800 6 la_data_out[1]
port 284 nsew default output
rlabel metal2 s 64694 0 64750 800 6 la_data_out[20]
port 285 nsew default output
rlabel metal2 s 65798 0 65854 800 6 la_data_out[21]
port 286 nsew default output
rlabel metal2 s 66994 0 67050 800 6 la_data_out[22]
port 287 nsew default output
rlabel metal2 s 68098 0 68154 800 6 la_data_out[23]
port 288 nsew default output
rlabel metal2 s 69294 0 69350 800 6 la_data_out[24]
port 289 nsew default output
rlabel metal2 s 70490 0 70546 800 6 la_data_out[25]
port 290 nsew default output
rlabel metal2 s 71594 0 71650 800 6 la_data_out[26]
port 291 nsew default output
rlabel metal2 s 72790 0 72846 800 6 la_data_out[27]
port 292 nsew default output
rlabel metal2 s 73894 0 73950 800 6 la_data_out[28]
port 293 nsew default output
rlabel metal2 s 75090 0 75146 800 6 la_data_out[29]
port 294 nsew default output
rlabel metal2 s 43810 0 43866 800 6 la_data_out[2]
port 295 nsew default output
rlabel metal2 s 76286 0 76342 800 6 la_data_out[30]
port 296 nsew default output
rlabel metal2 s 77390 0 77446 800 6 la_data_out[31]
port 297 nsew default output
rlabel metal2 s 78586 0 78642 800 6 la_data_out[32]
port 298 nsew default output
rlabel metal2 s 79690 0 79746 800 6 la_data_out[33]
port 299 nsew default output
rlabel metal2 s 80886 0 80942 800 6 la_data_out[34]
port 300 nsew default output
rlabel metal2 s 82082 0 82138 800 6 la_data_out[35]
port 301 nsew default output
rlabel metal2 s 83186 0 83242 800 6 la_data_out[36]
port 302 nsew default output
rlabel metal2 s 84382 0 84438 800 6 la_data_out[37]
port 303 nsew default output
rlabel metal2 s 85486 0 85542 800 6 la_data_out[38]
port 304 nsew default output
rlabel metal2 s 86682 0 86738 800 6 la_data_out[39]
port 305 nsew default output
rlabel metal2 s 45006 0 45062 800 6 la_data_out[3]
port 306 nsew default output
rlabel metal2 s 87878 0 87934 800 6 la_data_out[40]
port 307 nsew default output
rlabel metal2 s 88982 0 89038 800 6 la_data_out[41]
port 308 nsew default output
rlabel metal2 s 90178 0 90234 800 6 la_data_out[42]
port 309 nsew default output
rlabel metal2 s 91282 0 91338 800 6 la_data_out[43]
port 310 nsew default output
rlabel metal2 s 92478 0 92534 800 6 la_data_out[44]
port 311 nsew default output
rlabel metal2 s 93674 0 93730 800 6 la_data_out[45]
port 312 nsew default output
rlabel metal2 s 94778 0 94834 800 6 la_data_out[46]
port 313 nsew default output
rlabel metal2 s 95974 0 96030 800 6 la_data_out[47]
port 314 nsew default output
rlabel metal2 s 97078 0 97134 800 6 la_data_out[48]
port 315 nsew default output
rlabel metal2 s 98274 0 98330 800 6 la_data_out[49]
port 316 nsew default output
rlabel metal2 s 46110 0 46166 800 6 la_data_out[4]
port 317 nsew default output
rlabel metal2 s 99470 0 99526 800 6 la_data_out[50]
port 318 nsew default output
rlabel metal2 s 100574 0 100630 800 6 la_data_out[51]
port 319 nsew default output
rlabel metal2 s 101770 0 101826 800 6 la_data_out[52]
port 320 nsew default output
rlabel metal2 s 102874 0 102930 800 6 la_data_out[53]
port 321 nsew default output
rlabel metal2 s 104070 0 104126 800 6 la_data_out[54]
port 322 nsew default output
rlabel metal2 s 105266 0 105322 800 6 la_data_out[55]
port 323 nsew default output
rlabel metal2 s 106370 0 106426 800 6 la_data_out[56]
port 324 nsew default output
rlabel metal2 s 107566 0 107622 800 6 la_data_out[57]
port 325 nsew default output
rlabel metal2 s 108670 0 108726 800 6 la_data_out[58]
port 326 nsew default output
rlabel metal2 s 109866 0 109922 800 6 la_data_out[59]
port 327 nsew default output
rlabel metal2 s 47306 0 47362 800 6 la_data_out[5]
port 328 nsew default output
rlabel metal2 s 111062 0 111118 800 6 la_data_out[60]
port 329 nsew default output
rlabel metal2 s 112166 0 112222 800 6 la_data_out[61]
port 330 nsew default output
rlabel metal2 s 113362 0 113418 800 6 la_data_out[62]
port 331 nsew default output
rlabel metal2 s 114466 0 114522 800 6 la_data_out[63]
port 332 nsew default output
rlabel metal2 s 115662 0 115718 800 6 la_data_out[64]
port 333 nsew default output
rlabel metal2 s 116858 0 116914 800 6 la_data_out[65]
port 334 nsew default output
rlabel metal2 s 117962 0 118018 800 6 la_data_out[66]
port 335 nsew default output
rlabel metal2 s 119158 0 119214 800 6 la_data_out[67]
port 336 nsew default output
rlabel metal2 s 120262 0 120318 800 6 la_data_out[68]
port 337 nsew default output
rlabel metal2 s 121458 0 121514 800 6 la_data_out[69]
port 338 nsew default output
rlabel metal2 s 48410 0 48466 800 6 la_data_out[6]
port 339 nsew default output
rlabel metal2 s 122654 0 122710 800 6 la_data_out[70]
port 340 nsew default output
rlabel metal2 s 123758 0 123814 800 6 la_data_out[71]
port 341 nsew default output
rlabel metal2 s 124954 0 125010 800 6 la_data_out[72]
port 342 nsew default output
rlabel metal2 s 126058 0 126114 800 6 la_data_out[73]
port 343 nsew default output
rlabel metal2 s 127254 0 127310 800 6 la_data_out[74]
port 344 nsew default output
rlabel metal2 s 128450 0 128506 800 6 la_data_out[75]
port 345 nsew default output
rlabel metal2 s 129554 0 129610 800 6 la_data_out[76]
port 346 nsew default output
rlabel metal2 s 130750 0 130806 800 6 la_data_out[77]
port 347 nsew default output
rlabel metal2 s 131854 0 131910 800 6 la_data_out[78]
port 348 nsew default output
rlabel metal2 s 133050 0 133106 800 6 la_data_out[79]
port 349 nsew default output
rlabel metal2 s 49606 0 49662 800 6 la_data_out[7]
port 350 nsew default output
rlabel metal2 s 134246 0 134302 800 6 la_data_out[80]
port 351 nsew default output
rlabel metal2 s 135350 0 135406 800 6 la_data_out[81]
port 352 nsew default output
rlabel metal2 s 136546 0 136602 800 6 la_data_out[82]
port 353 nsew default output
rlabel metal2 s 137650 0 137706 800 6 la_data_out[83]
port 354 nsew default output
rlabel metal2 s 138846 0 138902 800 6 la_data_out[84]
port 355 nsew default output
rlabel metal2 s 139950 0 140006 800 6 la_data_out[85]
port 356 nsew default output
rlabel metal2 s 141146 0 141202 800 6 la_data_out[86]
port 357 nsew default output
rlabel metal2 s 142342 0 142398 800 6 la_data_out[87]
port 358 nsew default output
rlabel metal2 s 143446 0 143502 800 6 la_data_out[88]
port 359 nsew default output
rlabel metal2 s 144642 0 144698 800 6 la_data_out[89]
port 360 nsew default output
rlabel metal2 s 50802 0 50858 800 6 la_data_out[8]
port 361 nsew default output
rlabel metal2 s 145746 0 145802 800 6 la_data_out[90]
port 362 nsew default output
rlabel metal2 s 146942 0 146998 800 6 la_data_out[91]
port 363 nsew default output
rlabel metal2 s 148138 0 148194 800 6 la_data_out[92]
port 364 nsew default output
rlabel metal2 s 149242 0 149298 800 6 la_data_out[93]
port 365 nsew default output
rlabel metal2 s 150438 0 150494 800 6 la_data_out[94]
port 366 nsew default output
rlabel metal2 s 151542 0 151598 800 6 la_data_out[95]
port 367 nsew default output
rlabel metal2 s 152738 0 152794 800 6 la_data_out[96]
port 368 nsew default output
rlabel metal2 s 153934 0 153990 800 6 la_data_out[97]
port 369 nsew default output
rlabel metal2 s 155038 0 155094 800 6 la_data_out[98]
port 370 nsew default output
rlabel metal2 s 156234 0 156290 800 6 la_data_out[99]
port 371 nsew default output
rlabel metal2 s 51906 0 51962 800 6 la_data_out[9]
port 372 nsew default output
rlabel metal2 s 41878 0 41934 800 6 la_oen[0]
port 373 nsew default input
rlabel metal2 s 157798 0 157854 800 6 la_oen[100]
port 374 nsew default input
rlabel metal2 s 158902 0 158958 800 6 la_oen[101]
port 375 nsew default input
rlabel metal2 s 160098 0 160154 800 6 la_oen[102]
port 376 nsew default input
rlabel metal2 s 161202 0 161258 800 6 la_oen[103]
port 377 nsew default input
rlabel metal2 s 162398 0 162454 800 6 la_oen[104]
port 378 nsew default input
rlabel metal2 s 163594 0 163650 800 6 la_oen[105]
port 379 nsew default input
rlabel metal2 s 164698 0 164754 800 6 la_oen[106]
port 380 nsew default input
rlabel metal2 s 165894 0 165950 800 6 la_oen[107]
port 381 nsew default input
rlabel metal2 s 166998 0 167054 800 6 la_oen[108]
port 382 nsew default input
rlabel metal2 s 168194 0 168250 800 6 la_oen[109]
port 383 nsew default input
rlabel metal2 s 53470 0 53526 800 6 la_oen[10]
port 384 nsew default input
rlabel metal2 s 169390 0 169446 800 6 la_oen[110]
port 385 nsew default input
rlabel metal2 s 170494 0 170550 800 6 la_oen[111]
port 386 nsew default input
rlabel metal2 s 171690 0 171746 800 6 la_oen[112]
port 387 nsew default input
rlabel metal2 s 172794 0 172850 800 6 la_oen[113]
port 388 nsew default input
rlabel metal2 s 173990 0 174046 800 6 la_oen[114]
port 389 nsew default input
rlabel metal2 s 175186 0 175242 800 6 la_oen[115]
port 390 nsew default input
rlabel metal2 s 176290 0 176346 800 6 la_oen[116]
port 391 nsew default input
rlabel metal2 s 177486 0 177542 800 6 la_oen[117]
port 392 nsew default input
rlabel metal2 s 178590 0 178646 800 6 la_oen[118]
port 393 nsew default input
rlabel metal2 s 179786 0 179842 800 6 la_oen[119]
port 394 nsew default input
rlabel metal2 s 54666 0 54722 800 6 la_oen[11]
port 395 nsew default input
rlabel metal2 s 180982 0 181038 800 6 la_oen[120]
port 396 nsew default input
rlabel metal2 s 182086 0 182142 800 6 la_oen[121]
port 397 nsew default input
rlabel metal2 s 183282 0 183338 800 6 la_oen[122]
port 398 nsew default input
rlabel metal2 s 184386 0 184442 800 6 la_oen[123]
port 399 nsew default input
rlabel metal2 s 185582 0 185638 800 6 la_oen[124]
port 400 nsew default input
rlabel metal2 s 186778 0 186834 800 6 la_oen[125]
port 401 nsew default input
rlabel metal2 s 187882 0 187938 800 6 la_oen[126]
port 402 nsew default input
rlabel metal2 s 189078 0 189134 800 6 la_oen[127]
port 403 nsew default input
rlabel metal2 s 55770 0 55826 800 6 la_oen[12]
port 404 nsew default input
rlabel metal2 s 56966 0 57022 800 6 la_oen[13]
port 405 nsew default input
rlabel metal2 s 58070 0 58126 800 6 la_oen[14]
port 406 nsew default input
rlabel metal2 s 59266 0 59322 800 6 la_oen[15]
port 407 nsew default input
rlabel metal2 s 60462 0 60518 800 6 la_oen[16]
port 408 nsew default input
rlabel metal2 s 61566 0 61622 800 6 la_oen[17]
port 409 nsew default input
rlabel metal2 s 62762 0 62818 800 6 la_oen[18]
port 410 nsew default input
rlabel metal2 s 63866 0 63922 800 6 la_oen[19]
port 411 nsew default input
rlabel metal2 s 43074 0 43130 800 6 la_oen[1]
port 412 nsew default input
rlabel metal2 s 65062 0 65118 800 6 la_oen[20]
port 413 nsew default input
rlabel metal2 s 66258 0 66314 800 6 la_oen[21]
port 414 nsew default input
rlabel metal2 s 67362 0 67418 800 6 la_oen[22]
port 415 nsew default input
rlabel metal2 s 68558 0 68614 800 6 la_oen[23]
port 416 nsew default input
rlabel metal2 s 69662 0 69718 800 6 la_oen[24]
port 417 nsew default input
rlabel metal2 s 70858 0 70914 800 6 la_oen[25]
port 418 nsew default input
rlabel metal2 s 71962 0 72018 800 6 la_oen[26]
port 419 nsew default input
rlabel metal2 s 73158 0 73214 800 6 la_oen[27]
port 420 nsew default input
rlabel metal2 s 74354 0 74410 800 6 la_oen[28]
port 421 nsew default input
rlabel metal2 s 75458 0 75514 800 6 la_oen[29]
port 422 nsew default input
rlabel metal2 s 44178 0 44234 800 6 la_oen[2]
port 423 nsew default input
rlabel metal2 s 76654 0 76710 800 6 la_oen[30]
port 424 nsew default input
rlabel metal2 s 77758 0 77814 800 6 la_oen[31]
port 425 nsew default input
rlabel metal2 s 78954 0 79010 800 6 la_oen[32]
port 426 nsew default input
rlabel metal2 s 80150 0 80206 800 6 la_oen[33]
port 427 nsew default input
rlabel metal2 s 81254 0 81310 800 6 la_oen[34]
port 428 nsew default input
rlabel metal2 s 82450 0 82506 800 6 la_oen[35]
port 429 nsew default input
rlabel metal2 s 83554 0 83610 800 6 la_oen[36]
port 430 nsew default input
rlabel metal2 s 84750 0 84806 800 6 la_oen[37]
port 431 nsew default input
rlabel metal2 s 85946 0 86002 800 6 la_oen[38]
port 432 nsew default input
rlabel metal2 s 87050 0 87106 800 6 la_oen[39]
port 433 nsew default input
rlabel metal2 s 45374 0 45430 800 6 la_oen[3]
port 434 nsew default input
rlabel metal2 s 88246 0 88302 800 6 la_oen[40]
port 435 nsew default input
rlabel metal2 s 89350 0 89406 800 6 la_oen[41]
port 436 nsew default input
rlabel metal2 s 90546 0 90602 800 6 la_oen[42]
port 437 nsew default input
rlabel metal2 s 91742 0 91798 800 6 la_oen[43]
port 438 nsew default input
rlabel metal2 s 92846 0 92902 800 6 la_oen[44]
port 439 nsew default input
rlabel metal2 s 94042 0 94098 800 6 la_oen[45]
port 440 nsew default input
rlabel metal2 s 95146 0 95202 800 6 la_oen[46]
port 441 nsew default input
rlabel metal2 s 96342 0 96398 800 6 la_oen[47]
port 442 nsew default input
rlabel metal2 s 97538 0 97594 800 6 la_oen[48]
port 443 nsew default input
rlabel metal2 s 98642 0 98698 800 6 la_oen[49]
port 444 nsew default input
rlabel metal2 s 46478 0 46534 800 6 la_oen[4]
port 445 nsew default input
rlabel metal2 s 99838 0 99894 800 6 la_oen[50]
port 446 nsew default input
rlabel metal2 s 100942 0 100998 800 6 la_oen[51]
port 447 nsew default input
rlabel metal2 s 102138 0 102194 800 6 la_oen[52]
port 448 nsew default input
rlabel metal2 s 103334 0 103390 800 6 la_oen[53]
port 449 nsew default input
rlabel metal2 s 104438 0 104494 800 6 la_oen[54]
port 450 nsew default input
rlabel metal2 s 105634 0 105690 800 6 la_oen[55]
port 451 nsew default input
rlabel metal2 s 106738 0 106794 800 6 la_oen[56]
port 452 nsew default input
rlabel metal2 s 107934 0 107990 800 6 la_oen[57]
port 453 nsew default input
rlabel metal2 s 109130 0 109186 800 6 la_oen[58]
port 454 nsew default input
rlabel metal2 s 110234 0 110290 800 6 la_oen[59]
port 455 nsew default input
rlabel metal2 s 47674 0 47730 800 6 la_oen[5]
port 456 nsew default input
rlabel metal2 s 111430 0 111486 800 6 la_oen[60]
port 457 nsew default input
rlabel metal2 s 112534 0 112590 800 6 la_oen[61]
port 458 nsew default input
rlabel metal2 s 113730 0 113786 800 6 la_oen[62]
port 459 nsew default input
rlabel metal2 s 114926 0 114982 800 6 la_oen[63]
port 460 nsew default input
rlabel metal2 s 116030 0 116086 800 6 la_oen[64]
port 461 nsew default input
rlabel metal2 s 117226 0 117282 800 6 la_oen[65]
port 462 nsew default input
rlabel metal2 s 118330 0 118386 800 6 la_oen[66]
port 463 nsew default input
rlabel metal2 s 119526 0 119582 800 6 la_oen[67]
port 464 nsew default input
rlabel metal2 s 120722 0 120778 800 6 la_oen[68]
port 465 nsew default input
rlabel metal2 s 121826 0 121882 800 6 la_oen[69]
port 466 nsew default input
rlabel metal2 s 48870 0 48926 800 6 la_oen[6]
port 467 nsew default input
rlabel metal2 s 123022 0 123078 800 6 la_oen[70]
port 468 nsew default input
rlabel metal2 s 124126 0 124182 800 6 la_oen[71]
port 469 nsew default input
rlabel metal2 s 125322 0 125378 800 6 la_oen[72]
port 470 nsew default input
rlabel metal2 s 126518 0 126574 800 6 la_oen[73]
port 471 nsew default input
rlabel metal2 s 127622 0 127678 800 6 la_oen[74]
port 472 nsew default input
rlabel metal2 s 128818 0 128874 800 6 la_oen[75]
port 473 nsew default input
rlabel metal2 s 129922 0 129978 800 6 la_oen[76]
port 474 nsew default input
rlabel metal2 s 131118 0 131174 800 6 la_oen[77]
port 475 nsew default input
rlabel metal2 s 132314 0 132370 800 6 la_oen[78]
port 476 nsew default input
rlabel metal2 s 133418 0 133474 800 6 la_oen[79]
port 477 nsew default input
rlabel metal2 s 49974 0 50030 800 6 la_oen[7]
port 478 nsew default input
rlabel metal2 s 134614 0 134670 800 6 la_oen[80]
port 479 nsew default input
rlabel metal2 s 135718 0 135774 800 6 la_oen[81]
port 480 nsew default input
rlabel metal2 s 136914 0 136970 800 6 la_oen[82]
port 481 nsew default input
rlabel metal2 s 138018 0 138074 800 6 la_oen[83]
port 482 nsew default input
rlabel metal2 s 139214 0 139270 800 6 la_oen[84]
port 483 nsew default input
rlabel metal2 s 140410 0 140466 800 6 la_oen[85]
port 484 nsew default input
rlabel metal2 s 141514 0 141570 800 6 la_oen[86]
port 485 nsew default input
rlabel metal2 s 142710 0 142766 800 6 la_oen[87]
port 486 nsew default input
rlabel metal2 s 143814 0 143870 800 6 la_oen[88]
port 487 nsew default input
rlabel metal2 s 145010 0 145066 800 6 la_oen[89]
port 488 nsew default input
rlabel metal2 s 51170 0 51226 800 6 la_oen[8]
port 489 nsew default input
rlabel metal2 s 146206 0 146262 800 6 la_oen[90]
port 490 nsew default input
rlabel metal2 s 147310 0 147366 800 6 la_oen[91]
port 491 nsew default input
rlabel metal2 s 148506 0 148562 800 6 la_oen[92]
port 492 nsew default input
rlabel metal2 s 149610 0 149666 800 6 la_oen[93]
port 493 nsew default input
rlabel metal2 s 150806 0 150862 800 6 la_oen[94]
port 494 nsew default input
rlabel metal2 s 152002 0 152058 800 6 la_oen[95]
port 495 nsew default input
rlabel metal2 s 153106 0 153162 800 6 la_oen[96]
port 496 nsew default input
rlabel metal2 s 154302 0 154358 800 6 la_oen[97]
port 497 nsew default input
rlabel metal2 s 155406 0 155462 800 6 la_oen[98]
port 498 nsew default input
rlabel metal2 s 156602 0 156658 800 6 la_oen[99]
port 499 nsew default input
rlabel metal2 s 52274 0 52330 800 6 la_oen[9]
port 500 nsew default input
rlabel metal2 s 202 0 258 800 6 wb_clk_i
port 501 nsew default input
rlabel metal2 s 570 0 626 800 6 wb_rst_i
port 502 nsew default input
rlabel metal2 s 938 0 994 800 6 wbs_ack_o
port 503 nsew default output
rlabel metal2 s 2502 0 2558 800 6 wbs_adr_i[0]
port 504 nsew default input
rlabel metal2 s 15566 0 15622 800 6 wbs_adr_i[10]
port 505 nsew default input
rlabel metal2 s 16762 0 16818 800 6 wbs_adr_i[11]
port 506 nsew default input
rlabel metal2 s 17958 0 18014 800 6 wbs_adr_i[12]
port 507 nsew default input
rlabel metal2 s 19062 0 19118 800 6 wbs_adr_i[13]
port 508 nsew default input
rlabel metal2 s 20258 0 20314 800 6 wbs_adr_i[14]
port 509 nsew default input
rlabel metal2 s 21362 0 21418 800 6 wbs_adr_i[15]
port 510 nsew default input
rlabel metal2 s 22558 0 22614 800 6 wbs_adr_i[16]
port 511 nsew default input
rlabel metal2 s 23754 0 23810 800 6 wbs_adr_i[17]
port 512 nsew default input
rlabel metal2 s 24858 0 24914 800 6 wbs_adr_i[18]
port 513 nsew default input
rlabel metal2 s 26054 0 26110 800 6 wbs_adr_i[19]
port 514 nsew default input
rlabel metal2 s 3974 0 4030 800 6 wbs_adr_i[1]
port 515 nsew default input
rlabel metal2 s 27158 0 27214 800 6 wbs_adr_i[20]
port 516 nsew default input
rlabel metal2 s 28354 0 28410 800 6 wbs_adr_i[21]
port 517 nsew default input
rlabel metal2 s 29550 0 29606 800 6 wbs_adr_i[22]
port 518 nsew default input
rlabel metal2 s 30654 0 30710 800 6 wbs_adr_i[23]
port 519 nsew default input
rlabel metal2 s 31850 0 31906 800 6 wbs_adr_i[24]
port 520 nsew default input
rlabel metal2 s 32954 0 33010 800 6 wbs_adr_i[25]
port 521 nsew default input
rlabel metal2 s 34150 0 34206 800 6 wbs_adr_i[26]
port 522 nsew default input
rlabel metal2 s 35346 0 35402 800 6 wbs_adr_i[27]
port 523 nsew default input
rlabel metal2 s 36450 0 36506 800 6 wbs_adr_i[28]
port 524 nsew default input
rlabel metal2 s 37646 0 37702 800 6 wbs_adr_i[29]
port 525 nsew default input
rlabel metal2 s 5538 0 5594 800 6 wbs_adr_i[2]
port 526 nsew default input
rlabel metal2 s 38750 0 38806 800 6 wbs_adr_i[30]
port 527 nsew default input
rlabel metal2 s 39946 0 40002 800 6 wbs_adr_i[31]
port 528 nsew default input
rlabel metal2 s 7102 0 7158 800 6 wbs_adr_i[3]
port 529 nsew default input
rlabel metal2 s 8666 0 8722 800 6 wbs_adr_i[4]
port 530 nsew default input
rlabel metal2 s 9770 0 9826 800 6 wbs_adr_i[5]
port 531 nsew default input
rlabel metal2 s 10966 0 11022 800 6 wbs_adr_i[6]
port 532 nsew default input
rlabel metal2 s 12162 0 12218 800 6 wbs_adr_i[7]
port 533 nsew default input
rlabel metal2 s 13266 0 13322 800 6 wbs_adr_i[8]
port 534 nsew default input
rlabel metal2 s 14462 0 14518 800 6 wbs_adr_i[9]
port 535 nsew default input
rlabel metal2 s 1306 0 1362 800 6 wbs_cyc_i
port 536 nsew default input
rlabel metal2 s 2870 0 2926 800 6 wbs_dat_i[0]
port 537 nsew default input
rlabel metal2 s 16026 0 16082 800 6 wbs_dat_i[10]
port 538 nsew default input
rlabel metal2 s 17130 0 17186 800 6 wbs_dat_i[11]
port 539 nsew default input
rlabel metal2 s 18326 0 18382 800 6 wbs_dat_i[12]
port 540 nsew default input
rlabel metal2 s 19430 0 19486 800 6 wbs_dat_i[13]
port 541 nsew default input
rlabel metal2 s 20626 0 20682 800 6 wbs_dat_i[14]
port 542 nsew default input
rlabel metal2 s 21822 0 21878 800 6 wbs_dat_i[15]
port 543 nsew default input
rlabel metal2 s 22926 0 22982 800 6 wbs_dat_i[16]
port 544 nsew default input
rlabel metal2 s 24122 0 24178 800 6 wbs_dat_i[17]
port 545 nsew default input
rlabel metal2 s 25226 0 25282 800 6 wbs_dat_i[18]
port 546 nsew default input
rlabel metal2 s 26422 0 26478 800 6 wbs_dat_i[19]
port 547 nsew default input
rlabel metal2 s 4434 0 4490 800 6 wbs_dat_i[1]
port 548 nsew default input
rlabel metal2 s 27618 0 27674 800 6 wbs_dat_i[20]
port 549 nsew default input
rlabel metal2 s 28722 0 28778 800 6 wbs_dat_i[21]
port 550 nsew default input
rlabel metal2 s 29918 0 29974 800 6 wbs_dat_i[22]
port 551 nsew default input
rlabel metal2 s 31022 0 31078 800 6 wbs_dat_i[23]
port 552 nsew default input
rlabel metal2 s 32218 0 32274 800 6 wbs_dat_i[24]
port 553 nsew default input
rlabel metal2 s 33414 0 33470 800 6 wbs_dat_i[25]
port 554 nsew default input
rlabel metal2 s 34518 0 34574 800 6 wbs_dat_i[26]
port 555 nsew default input
rlabel metal2 s 35714 0 35770 800 6 wbs_dat_i[27]
port 556 nsew default input
rlabel metal2 s 36818 0 36874 800 6 wbs_dat_i[28]
port 557 nsew default input
rlabel metal2 s 38014 0 38070 800 6 wbs_dat_i[29]
port 558 nsew default input
rlabel metal2 s 5906 0 5962 800 6 wbs_dat_i[2]
port 559 nsew default input
rlabel metal2 s 39210 0 39266 800 6 wbs_dat_i[30]
port 560 nsew default input
rlabel metal2 s 40314 0 40370 800 6 wbs_dat_i[31]
port 561 nsew default input
rlabel metal2 s 7470 0 7526 800 6 wbs_dat_i[3]
port 562 nsew default input
rlabel metal2 s 9034 0 9090 800 6 wbs_dat_i[4]
port 563 nsew default input
rlabel metal2 s 10230 0 10286 800 6 wbs_dat_i[5]
port 564 nsew default input
rlabel metal2 s 11334 0 11390 800 6 wbs_dat_i[6]
port 565 nsew default input
rlabel metal2 s 12530 0 12586 800 6 wbs_dat_i[7]
port 566 nsew default input
rlabel metal2 s 13634 0 13690 800 6 wbs_dat_i[8]
port 567 nsew default input
rlabel metal2 s 14830 0 14886 800 6 wbs_dat_i[9]
port 568 nsew default input
rlabel metal2 s 3238 0 3294 800 6 wbs_dat_o[0]
port 569 nsew default output
rlabel metal2 s 16394 0 16450 800 6 wbs_dat_o[10]
port 570 nsew default output
rlabel metal2 s 17498 0 17554 800 6 wbs_dat_o[11]
port 571 nsew default output
rlabel metal2 s 18694 0 18750 800 6 wbs_dat_o[12]
port 572 nsew default output
rlabel metal2 s 19890 0 19946 800 6 wbs_dat_o[13]
port 573 nsew default output
rlabel metal2 s 20994 0 21050 800 6 wbs_dat_o[14]
port 574 nsew default output
rlabel metal2 s 22190 0 22246 800 6 wbs_dat_o[15]
port 575 nsew default output
rlabel metal2 s 23294 0 23350 800 6 wbs_dat_o[16]
port 576 nsew default output
rlabel metal2 s 24490 0 24546 800 6 wbs_dat_o[17]
port 577 nsew default output
rlabel metal2 s 25686 0 25742 800 6 wbs_dat_o[18]
port 578 nsew default output
rlabel metal2 s 26790 0 26846 800 6 wbs_dat_o[19]
port 579 nsew default output
rlabel metal2 s 4802 0 4858 800 6 wbs_dat_o[1]
port 580 nsew default output
rlabel metal2 s 27986 0 28042 800 6 wbs_dat_o[20]
port 581 nsew default output
rlabel metal2 s 29090 0 29146 800 6 wbs_dat_o[21]
port 582 nsew default output
rlabel metal2 s 30286 0 30342 800 6 wbs_dat_o[22]
port 583 nsew default output
rlabel metal2 s 31482 0 31538 800 6 wbs_dat_o[23]
port 584 nsew default output
rlabel metal2 s 32586 0 32642 800 6 wbs_dat_o[24]
port 585 nsew default output
rlabel metal2 s 33782 0 33838 800 6 wbs_dat_o[25]
port 586 nsew default output
rlabel metal2 s 34886 0 34942 800 6 wbs_dat_o[26]
port 587 nsew default output
rlabel metal2 s 36082 0 36138 800 6 wbs_dat_o[27]
port 588 nsew default output
rlabel metal2 s 37278 0 37334 800 6 wbs_dat_o[28]
port 589 nsew default output
rlabel metal2 s 38382 0 38438 800 6 wbs_dat_o[29]
port 590 nsew default output
rlabel metal2 s 6366 0 6422 800 6 wbs_dat_o[2]
port 591 nsew default output
rlabel metal2 s 39578 0 39634 800 6 wbs_dat_o[30]
port 592 nsew default output
rlabel metal2 s 40682 0 40738 800 6 wbs_dat_o[31]
port 593 nsew default output
rlabel metal2 s 7838 0 7894 800 6 wbs_dat_o[3]
port 594 nsew default output
rlabel metal2 s 9402 0 9458 800 6 wbs_dat_o[4]
port 595 nsew default output
rlabel metal2 s 10598 0 10654 800 6 wbs_dat_o[5]
port 596 nsew default output
rlabel metal2 s 11702 0 11758 800 6 wbs_dat_o[6]
port 597 nsew default output
rlabel metal2 s 12898 0 12954 800 6 wbs_dat_o[7]
port 598 nsew default output
rlabel metal2 s 14094 0 14150 800 6 wbs_dat_o[8]
port 599 nsew default output
rlabel metal2 s 15198 0 15254 800 6 wbs_dat_o[9]
port 600 nsew default output
rlabel metal2 s 3606 0 3662 800 6 wbs_sel_i[0]
port 601 nsew default input
rlabel metal2 s 5170 0 5226 800 6 wbs_sel_i[1]
port 602 nsew default input
rlabel metal2 s 6734 0 6790 800 6 wbs_sel_i[2]
port 603 nsew default input
rlabel metal2 s 8298 0 8354 800 6 wbs_sel_i[3]
port 604 nsew default input
rlabel metal2 s 1674 0 1730 800 6 wbs_stb_i
port 605 nsew default input
rlabel metal2 s 2042 0 2098 800 6 wbs_we_i
port 606 nsew default input
rlabel metal4 s 4208 2128 4528 199696 6 VPWR
port 607 nsew power input
rlabel metal4 s 19568 2128 19888 199696 6 VGND
port 608 nsew ground input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 202000 202000
string LEFview TRUE
<< end >>
