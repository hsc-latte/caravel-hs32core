VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO hs32_core1
  CLASS BLOCK ;
  FOREIGN hs32_core1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1099.930 BY 1100.000 ;
  PIN cpu_addr_e[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 67.360 1099.930 67.960 ;
    END
  END cpu_addr_e[0]
  PIN cpu_addr_e[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 117.680 1099.930 118.280 ;
    END
  END cpu_addr_e[10]
  PIN cpu_addr_e[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 123.120 1099.930 123.720 ;
    END
  END cpu_addr_e[11]
  PIN cpu_addr_e[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 127.880 1099.930 128.480 ;
    END
  END cpu_addr_e[12]
  PIN cpu_addr_e[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 132.640 1099.930 133.240 ;
    END
  END cpu_addr_e[13]
  PIN cpu_addr_e[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 138.080 1099.930 138.680 ;
    END
  END cpu_addr_e[14]
  PIN cpu_addr_e[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 142.840 1099.930 143.440 ;
    END
  END cpu_addr_e[15]
  PIN cpu_addr_e[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 72.120 1099.930 72.720 ;
    END
  END cpu_addr_e[1]
  PIN cpu_addr_e[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 77.560 1099.930 78.160 ;
    END
  END cpu_addr_e[2]
  PIN cpu_addr_e[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 82.320 1099.930 82.920 ;
    END
  END cpu_addr_e[3]
  PIN cpu_addr_e[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 87.760 1099.930 88.360 ;
    END
  END cpu_addr_e[4]
  PIN cpu_addr_e[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 92.520 1099.930 93.120 ;
    END
  END cpu_addr_e[5]
  PIN cpu_addr_e[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 97.960 1099.930 98.560 ;
    END
  END cpu_addr_e[6]
  PIN cpu_addr_e[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 102.720 1099.930 103.320 ;
    END
  END cpu_addr_e[7]
  PIN cpu_addr_e[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 107.480 1099.930 108.080 ;
    END
  END cpu_addr_e[8]
  PIN cpu_addr_e[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 112.920 1099.930 113.520 ;
    END
  END cpu_addr_e[9]
  PIN cpu_addr_n[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 108.580 1096.000 108.860 1100.000 ;
    END
  END cpu_addr_n[0]
  PIN cpu_addr_n[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 212.540 1096.000 212.820 1100.000 ;
    END
  END cpu_addr_n[10]
  PIN cpu_addr_n[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 222.660 1096.000 222.940 1100.000 ;
    END
  END cpu_addr_n[11]
  PIN cpu_addr_n[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 233.240 1096.000 233.520 1100.000 ;
    END
  END cpu_addr_n[12]
  PIN cpu_addr_n[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 243.360 1096.000 243.640 1100.000 ;
    END
  END cpu_addr_n[13]
  PIN cpu_addr_n[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 253.940 1096.000 254.220 1100.000 ;
    END
  END cpu_addr_n[14]
  PIN cpu_addr_n[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 264.060 1096.000 264.340 1100.000 ;
    END
  END cpu_addr_n[15]
  PIN cpu_addr_n[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 119.160 1096.000 119.440 1100.000 ;
    END
  END cpu_addr_n[1]
  PIN cpu_addr_n[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 129.280 1096.000 129.560 1100.000 ;
    END
  END cpu_addr_n[2]
  PIN cpu_addr_n[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 139.860 1096.000 140.140 1100.000 ;
    END
  END cpu_addr_n[3]
  PIN cpu_addr_n[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 149.980 1096.000 150.260 1100.000 ;
    END
  END cpu_addr_n[4]
  PIN cpu_addr_n[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 160.560 1096.000 160.840 1100.000 ;
    END
  END cpu_addr_n[5]
  PIN cpu_addr_n[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 170.680 1096.000 170.960 1100.000 ;
    END
  END cpu_addr_n[6]
  PIN cpu_addr_n[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 181.260 1096.000 181.540 1100.000 ;
    END
  END cpu_addr_n[7]
  PIN cpu_addr_n[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 191.840 1096.000 192.120 1100.000 ;
    END
  END cpu_addr_n[8]
  PIN cpu_addr_n[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 201.960 1096.000 202.240 1100.000 ;
    END
  END cpu_addr_n[9]
  PIN cpu_dtr_e0[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 228.520 1099.930 229.120 ;
    END
  END cpu_dtr_e0[0]
  PIN cpu_dtr_e0[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 279.520 1099.930 280.120 ;
    END
  END cpu_dtr_e0[10]
  PIN cpu_dtr_e0[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 284.280 1099.930 284.880 ;
    END
  END cpu_dtr_e0[11]
  PIN cpu_dtr_e0[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 289.720 1099.930 290.320 ;
    END
  END cpu_dtr_e0[12]
  PIN cpu_dtr_e0[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 294.480 1099.930 295.080 ;
    END
  END cpu_dtr_e0[13]
  PIN cpu_dtr_e0[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 299.240 1099.930 299.840 ;
    END
  END cpu_dtr_e0[14]
  PIN cpu_dtr_e0[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 304.680 1099.930 305.280 ;
    END
  END cpu_dtr_e0[15]
  PIN cpu_dtr_e0[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 309.440 1099.930 310.040 ;
    END
  END cpu_dtr_e0[16]
  PIN cpu_dtr_e0[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 314.880 1099.930 315.480 ;
    END
  END cpu_dtr_e0[17]
  PIN cpu_dtr_e0[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 319.640 1099.930 320.240 ;
    END
  END cpu_dtr_e0[18]
  PIN cpu_dtr_e0[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 325.080 1099.930 325.680 ;
    END
  END cpu_dtr_e0[19]
  PIN cpu_dtr_e0[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 233.960 1099.930 234.560 ;
    END
  END cpu_dtr_e0[1]
  PIN cpu_dtr_e0[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 329.840 1099.930 330.440 ;
    END
  END cpu_dtr_e0[20]
  PIN cpu_dtr_e0[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 334.600 1099.930 335.200 ;
    END
  END cpu_dtr_e0[21]
  PIN cpu_dtr_e0[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 340.040 1099.930 340.640 ;
    END
  END cpu_dtr_e0[22]
  PIN cpu_dtr_e0[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 344.800 1099.930 345.400 ;
    END
  END cpu_dtr_e0[23]
  PIN cpu_dtr_e0[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 350.240 1099.930 350.840 ;
    END
  END cpu_dtr_e0[24]
  PIN cpu_dtr_e0[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 355.000 1099.930 355.600 ;
    END
  END cpu_dtr_e0[25]
  PIN cpu_dtr_e0[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 359.760 1099.930 360.360 ;
    END
  END cpu_dtr_e0[26]
  PIN cpu_dtr_e0[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 365.200 1099.930 365.800 ;
    END
  END cpu_dtr_e0[27]
  PIN cpu_dtr_e0[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 369.960 1099.930 370.560 ;
    END
  END cpu_dtr_e0[28]
  PIN cpu_dtr_e0[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 375.400 1099.930 376.000 ;
    END
  END cpu_dtr_e0[29]
  PIN cpu_dtr_e0[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 238.720 1099.930 239.320 ;
    END
  END cpu_dtr_e0[2]
  PIN cpu_dtr_e0[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 380.160 1099.930 380.760 ;
    END
  END cpu_dtr_e0[30]
  PIN cpu_dtr_e0[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 385.600 1099.930 386.200 ;
    END
  END cpu_dtr_e0[31]
  PIN cpu_dtr_e0[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 244.160 1099.930 244.760 ;
    END
  END cpu_dtr_e0[3]
  PIN cpu_dtr_e0[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 248.920 1099.930 249.520 ;
    END
  END cpu_dtr_e0[4]
  PIN cpu_dtr_e0[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 254.360 1099.930 254.960 ;
    END
  END cpu_dtr_e0[5]
  PIN cpu_dtr_e0[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 259.120 1099.930 259.720 ;
    END
  END cpu_dtr_e0[6]
  PIN cpu_dtr_e0[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 263.880 1099.930 264.480 ;
    END
  END cpu_dtr_e0[7]
  PIN cpu_dtr_e0[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 269.320 1099.930 269.920 ;
    END
  END cpu_dtr_e0[8]
  PIN cpu_dtr_e0[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 274.080 1099.930 274.680 ;
    END
  END cpu_dtr_e0[9]
  PIN cpu_dtr_e1[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 390.360 1099.930 390.960 ;
    END
  END cpu_dtr_e1[0]
  PIN cpu_dtr_e1[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 440.680 1099.930 441.280 ;
    END
  END cpu_dtr_e1[10]
  PIN cpu_dtr_e1[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 446.120 1099.930 446.720 ;
    END
  END cpu_dtr_e1[11]
  PIN cpu_dtr_e1[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 450.880 1099.930 451.480 ;
    END
  END cpu_dtr_e1[12]
  PIN cpu_dtr_e1[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 455.640 1099.930 456.240 ;
    END
  END cpu_dtr_e1[13]
  PIN cpu_dtr_e1[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 461.080 1099.930 461.680 ;
    END
  END cpu_dtr_e1[14]
  PIN cpu_dtr_e1[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 465.840 1099.930 466.440 ;
    END
  END cpu_dtr_e1[15]
  PIN cpu_dtr_e1[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 471.280 1099.930 471.880 ;
    END
  END cpu_dtr_e1[16]
  PIN cpu_dtr_e1[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 476.040 1099.930 476.640 ;
    END
  END cpu_dtr_e1[17]
  PIN cpu_dtr_e1[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 481.480 1099.930 482.080 ;
    END
  END cpu_dtr_e1[18]
  PIN cpu_dtr_e1[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 486.240 1099.930 486.840 ;
    END
  END cpu_dtr_e1[19]
  PIN cpu_dtr_e1[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 395.120 1099.930 395.720 ;
    END
  END cpu_dtr_e1[1]
  PIN cpu_dtr_e1[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 491.000 1099.930 491.600 ;
    END
  END cpu_dtr_e1[20]
  PIN cpu_dtr_e1[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 496.440 1099.930 497.040 ;
    END
  END cpu_dtr_e1[21]
  PIN cpu_dtr_e1[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 501.200 1099.930 501.800 ;
    END
  END cpu_dtr_e1[22]
  PIN cpu_dtr_e1[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 506.640 1099.930 507.240 ;
    END
  END cpu_dtr_e1[23]
  PIN cpu_dtr_e1[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 511.400 1099.930 512.000 ;
    END
  END cpu_dtr_e1[24]
  PIN cpu_dtr_e1[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 516.840 1099.930 517.440 ;
    END
  END cpu_dtr_e1[25]
  PIN cpu_dtr_e1[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 521.600 1099.930 522.200 ;
    END
  END cpu_dtr_e1[26]
  PIN cpu_dtr_e1[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 526.360 1099.930 526.960 ;
    END
  END cpu_dtr_e1[27]
  PIN cpu_dtr_e1[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 531.800 1099.930 532.400 ;
    END
  END cpu_dtr_e1[28]
  PIN cpu_dtr_e1[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 536.560 1099.930 537.160 ;
    END
  END cpu_dtr_e1[29]
  PIN cpu_dtr_e1[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 400.560 1099.930 401.160 ;
    END
  END cpu_dtr_e1[2]
  PIN cpu_dtr_e1[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 542.000 1099.930 542.600 ;
    END
  END cpu_dtr_e1[30]
  PIN cpu_dtr_e1[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 546.760 1099.930 547.360 ;
    END
  END cpu_dtr_e1[31]
  PIN cpu_dtr_e1[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 405.320 1099.930 405.920 ;
    END
  END cpu_dtr_e1[3]
  PIN cpu_dtr_e1[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 410.760 1099.930 411.360 ;
    END
  END cpu_dtr_e1[4]
  PIN cpu_dtr_e1[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 415.520 1099.930 416.120 ;
    END
  END cpu_dtr_e1[5]
  PIN cpu_dtr_e1[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 420.960 1099.930 421.560 ;
    END
  END cpu_dtr_e1[6]
  PIN cpu_dtr_e1[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 425.720 1099.930 426.320 ;
    END
  END cpu_dtr_e1[7]
  PIN cpu_dtr_e1[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 430.480 1099.930 431.080 ;
    END
  END cpu_dtr_e1[8]
  PIN cpu_dtr_e1[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 435.920 1099.930 436.520 ;
    END
  END cpu_dtr_e1[9]
  PIN cpu_dtr_n0[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 440.700 1096.000 440.980 1100.000 ;
    END
  END cpu_dtr_n0[0]
  PIN cpu_dtr_n0[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 544.200 1096.000 544.480 1100.000 ;
    END
  END cpu_dtr_n0[10]
  PIN cpu_dtr_n0[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 554.780 1096.000 555.060 1100.000 ;
    END
  END cpu_dtr_n0[11]
  PIN cpu_dtr_n0[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 565.360 1096.000 565.640 1100.000 ;
    END
  END cpu_dtr_n0[12]
  PIN cpu_dtr_n0[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 575.480 1096.000 575.760 1100.000 ;
    END
  END cpu_dtr_n0[13]
  PIN cpu_dtr_n0[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 586.060 1096.000 586.340 1100.000 ;
    END
  END cpu_dtr_n0[14]
  PIN cpu_dtr_n0[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 596.180 1096.000 596.460 1100.000 ;
    END
  END cpu_dtr_n0[15]
  PIN cpu_dtr_n0[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 606.760 1096.000 607.040 1100.000 ;
    END
  END cpu_dtr_n0[16]
  PIN cpu_dtr_n0[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 616.880 1096.000 617.160 1100.000 ;
    END
  END cpu_dtr_n0[17]
  PIN cpu_dtr_n0[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 627.460 1096.000 627.740 1100.000 ;
    END
  END cpu_dtr_n0[18]
  PIN cpu_dtr_n0[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 637.580 1096.000 637.860 1100.000 ;
    END
  END cpu_dtr_n0[19]
  PIN cpu_dtr_n0[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 450.820 1096.000 451.100 1100.000 ;
    END
  END cpu_dtr_n0[1]
  PIN cpu_dtr_n0[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 648.160 1096.000 648.440 1100.000 ;
    END
  END cpu_dtr_n0[20]
  PIN cpu_dtr_n0[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 658.740 1096.000 659.020 1100.000 ;
    END
  END cpu_dtr_n0[21]
  PIN cpu_dtr_n0[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 668.860 1096.000 669.140 1100.000 ;
    END
  END cpu_dtr_n0[22]
  PIN cpu_dtr_n0[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 679.440 1096.000 679.720 1100.000 ;
    END
  END cpu_dtr_n0[23]
  PIN cpu_dtr_n0[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 689.560 1096.000 689.840 1100.000 ;
    END
  END cpu_dtr_n0[24]
  PIN cpu_dtr_n0[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 700.140 1096.000 700.420 1100.000 ;
    END
  END cpu_dtr_n0[25]
  PIN cpu_dtr_n0[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 710.260 1096.000 710.540 1100.000 ;
    END
  END cpu_dtr_n0[26]
  PIN cpu_dtr_n0[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 720.840 1096.000 721.120 1100.000 ;
    END
  END cpu_dtr_n0[27]
  PIN cpu_dtr_n0[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 730.960 1096.000 731.240 1100.000 ;
    END
  END cpu_dtr_n0[28]
  PIN cpu_dtr_n0[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 741.540 1096.000 741.820 1100.000 ;
    END
  END cpu_dtr_n0[29]
  PIN cpu_dtr_n0[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 461.400 1096.000 461.680 1100.000 ;
    END
  END cpu_dtr_n0[2]
  PIN cpu_dtr_n0[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 752.120 1096.000 752.400 1100.000 ;
    END
  END cpu_dtr_n0[30]
  PIN cpu_dtr_n0[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 762.240 1096.000 762.520 1100.000 ;
    END
  END cpu_dtr_n0[31]
  PIN cpu_dtr_n0[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 471.980 1096.000 472.260 1100.000 ;
    END
  END cpu_dtr_n0[3]
  PIN cpu_dtr_n0[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 482.100 1096.000 482.380 1100.000 ;
    END
  END cpu_dtr_n0[4]
  PIN cpu_dtr_n0[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 492.680 1096.000 492.960 1100.000 ;
    END
  END cpu_dtr_n0[5]
  PIN cpu_dtr_n0[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 502.800 1096.000 503.080 1100.000 ;
    END
  END cpu_dtr_n0[6]
  PIN cpu_dtr_n0[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 513.380 1096.000 513.660 1100.000 ;
    END
  END cpu_dtr_n0[7]
  PIN cpu_dtr_n0[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 523.500 1096.000 523.780 1100.000 ;
    END
  END cpu_dtr_n0[8]
  PIN cpu_dtr_n0[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 534.080 1096.000 534.360 1100.000 ;
    END
  END cpu_dtr_n0[9]
  PIN cpu_dtr_n1[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 772.820 1096.000 773.100 1100.000 ;
    END
  END cpu_dtr_n1[0]
  PIN cpu_dtr_n1[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 876.320 1096.000 876.600 1100.000 ;
    END
  END cpu_dtr_n1[10]
  PIN cpu_dtr_n1[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 886.900 1096.000 887.180 1100.000 ;
    END
  END cpu_dtr_n1[11]
  PIN cpu_dtr_n1[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 897.020 1096.000 897.300 1100.000 ;
    END
  END cpu_dtr_n1[12]
  PIN cpu_dtr_n1[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 907.600 1096.000 907.880 1100.000 ;
    END
  END cpu_dtr_n1[13]
  PIN cpu_dtr_n1[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 917.720 1096.000 918.000 1100.000 ;
    END
  END cpu_dtr_n1[14]
  PIN cpu_dtr_n1[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 928.300 1096.000 928.580 1100.000 ;
    END
  END cpu_dtr_n1[15]
  PIN cpu_dtr_n1[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 938.880 1096.000 939.160 1100.000 ;
    END
  END cpu_dtr_n1[16]
  PIN cpu_dtr_n1[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 949.000 1096.000 949.280 1100.000 ;
    END
  END cpu_dtr_n1[17]
  PIN cpu_dtr_n1[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 959.580 1096.000 959.860 1100.000 ;
    END
  END cpu_dtr_n1[18]
  PIN cpu_dtr_n1[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 969.700 1096.000 969.980 1100.000 ;
    END
  END cpu_dtr_n1[19]
  PIN cpu_dtr_n1[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 782.940 1096.000 783.220 1100.000 ;
    END
  END cpu_dtr_n1[1]
  PIN cpu_dtr_n1[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 980.280 1096.000 980.560 1100.000 ;
    END
  END cpu_dtr_n1[20]
  PIN cpu_dtr_n1[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 990.400 1096.000 990.680 1100.000 ;
    END
  END cpu_dtr_n1[21]
  PIN cpu_dtr_n1[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1000.980 1096.000 1001.260 1100.000 ;
    END
  END cpu_dtr_n1[22]
  PIN cpu_dtr_n1[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1011.100 1096.000 1011.380 1100.000 ;
    END
  END cpu_dtr_n1[23]
  PIN cpu_dtr_n1[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1021.680 1096.000 1021.960 1100.000 ;
    END
  END cpu_dtr_n1[24]
  PIN cpu_dtr_n1[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1032.260 1096.000 1032.540 1100.000 ;
    END
  END cpu_dtr_n1[25]
  PIN cpu_dtr_n1[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1042.380 1096.000 1042.660 1100.000 ;
    END
  END cpu_dtr_n1[26]
  PIN cpu_dtr_n1[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1052.960 1096.000 1053.240 1100.000 ;
    END
  END cpu_dtr_n1[27]
  PIN cpu_dtr_n1[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1063.080 1096.000 1063.360 1100.000 ;
    END
  END cpu_dtr_n1[28]
  PIN cpu_dtr_n1[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1073.660 1096.000 1073.940 1100.000 ;
    END
  END cpu_dtr_n1[29]
  PIN cpu_dtr_n1[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 793.520 1096.000 793.800 1100.000 ;
    END
  END cpu_dtr_n1[2]
  PIN cpu_dtr_n1[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1083.780 1096.000 1084.060 1100.000 ;
    END
  END cpu_dtr_n1[30]
  PIN cpu_dtr_n1[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1094.360 1096.000 1094.640 1100.000 ;
    END
  END cpu_dtr_n1[31]
  PIN cpu_dtr_n1[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 803.640 1096.000 803.920 1100.000 ;
    END
  END cpu_dtr_n1[3]
  PIN cpu_dtr_n1[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 814.220 1096.000 814.500 1100.000 ;
    END
  END cpu_dtr_n1[4]
  PIN cpu_dtr_n1[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 824.340 1096.000 824.620 1100.000 ;
    END
  END cpu_dtr_n1[5]
  PIN cpu_dtr_n1[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 834.920 1096.000 835.200 1100.000 ;
    END
  END cpu_dtr_n1[6]
  PIN cpu_dtr_n1[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 845.500 1096.000 845.780 1100.000 ;
    END
  END cpu_dtr_n1[7]
  PIN cpu_dtr_n1[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 855.620 1096.000 855.900 1100.000 ;
    END
  END cpu_dtr_n1[8]
  PIN cpu_dtr_n1[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 866.200 1096.000 866.480 1100.000 ;
    END
  END cpu_dtr_n1[9]
  PIN cpu_dtw_e[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 148.280 1099.930 148.880 ;
    END
  END cpu_dtw_e[0]
  PIN cpu_dtw_e[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 198.600 1099.930 199.200 ;
    END
  END cpu_dtw_e[10]
  PIN cpu_dtw_e[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 203.360 1099.930 203.960 ;
    END
  END cpu_dtw_e[11]
  PIN cpu_dtw_e[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 208.800 1099.930 209.400 ;
    END
  END cpu_dtw_e[12]
  PIN cpu_dtw_e[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 213.560 1099.930 214.160 ;
    END
  END cpu_dtw_e[13]
  PIN cpu_dtw_e[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 219.000 1099.930 219.600 ;
    END
  END cpu_dtw_e[14]
  PIN cpu_dtw_e[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 223.760 1099.930 224.360 ;
    END
  END cpu_dtw_e[15]
  PIN cpu_dtw_e[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 153.040 1099.930 153.640 ;
    END
  END cpu_dtw_e[1]
  PIN cpu_dtw_e[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 158.480 1099.930 159.080 ;
    END
  END cpu_dtw_e[2]
  PIN cpu_dtw_e[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 163.240 1099.930 163.840 ;
    END
  END cpu_dtw_e[3]
  PIN cpu_dtw_e[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 168.000 1099.930 168.600 ;
    END
  END cpu_dtw_e[4]
  PIN cpu_dtw_e[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 173.440 1099.930 174.040 ;
    END
  END cpu_dtw_e[5]
  PIN cpu_dtw_e[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 178.200 1099.930 178.800 ;
    END
  END cpu_dtw_e[6]
  PIN cpu_dtw_e[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 183.640 1099.930 184.240 ;
    END
  END cpu_dtw_e[7]
  PIN cpu_dtw_e[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 188.400 1099.930 189.000 ;
    END
  END cpu_dtw_e[8]
  PIN cpu_dtw_e[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 193.840 1099.930 194.440 ;
    END
  END cpu_dtw_e[9]
  PIN cpu_dtw_n[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 274.640 1096.000 274.920 1100.000 ;
    END
  END cpu_dtw_n[0]
  PIN cpu_dtw_n[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 378.600 1096.000 378.880 1100.000 ;
    END
  END cpu_dtw_n[10]
  PIN cpu_dtw_n[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 388.720 1096.000 389.000 1100.000 ;
    END
  END cpu_dtw_n[11]
  PIN cpu_dtw_n[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 399.300 1096.000 399.580 1100.000 ;
    END
  END cpu_dtw_n[12]
  PIN cpu_dtw_n[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 409.420 1096.000 409.700 1100.000 ;
    END
  END cpu_dtw_n[13]
  PIN cpu_dtw_n[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 420.000 1096.000 420.280 1100.000 ;
    END
  END cpu_dtw_n[14]
  PIN cpu_dtw_n[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 430.120 1096.000 430.400 1100.000 ;
    END
  END cpu_dtw_n[15]
  PIN cpu_dtw_n[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 285.220 1096.000 285.500 1100.000 ;
    END
  END cpu_dtw_n[1]
  PIN cpu_dtw_n[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 295.340 1096.000 295.620 1100.000 ;
    END
  END cpu_dtw_n[2]
  PIN cpu_dtw_n[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 305.920 1096.000 306.200 1100.000 ;
    END
  END cpu_dtw_n[3]
  PIN cpu_dtw_n[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 316.040 1096.000 316.320 1100.000 ;
    END
  END cpu_dtw_n[4]
  PIN cpu_dtw_n[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 326.620 1096.000 326.900 1100.000 ;
    END
  END cpu_dtw_n[5]
  PIN cpu_dtw_n[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 336.740 1096.000 337.020 1100.000 ;
    END
  END cpu_dtw_n[6]
  PIN cpu_dtw_n[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 347.320 1096.000 347.600 1100.000 ;
    END
  END cpu_dtw_n[7]
  PIN cpu_dtw_n[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 357.440 1096.000 357.720 1100.000 ;
    END
  END cpu_dtw_n[8]
  PIN cpu_dtw_n[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 368.020 1096.000 368.300 1100.000 ;
    END
  END cpu_dtw_n[9]
  PIN cpu_mask_e[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 17.040 1099.930 17.640 ;
    END
  END cpu_mask_e[0]
  PIN cpu_mask_e[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 21.800 1099.930 22.400 ;
    END
  END cpu_mask_e[1]
  PIN cpu_mask_e[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 27.240 1099.930 27.840 ;
    END
  END cpu_mask_e[2]
  PIN cpu_mask_e[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 32.000 1099.930 32.600 ;
    END
  END cpu_mask_e[3]
  PIN cpu_mask_e[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 36.760 1099.930 37.360 ;
    END
  END cpu_mask_e[4]
  PIN cpu_mask_e[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 42.200 1099.930 42.800 ;
    END
  END cpu_mask_e[5]
  PIN cpu_mask_e[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 46.960 1099.930 47.560 ;
    END
  END cpu_mask_e[6]
  PIN cpu_mask_e[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 52.400 1099.930 53.000 ;
    END
  END cpu_mask_e[7]
  PIN cpu_mask_n[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 5.080 1096.000 5.360 1100.000 ;
    END
  END cpu_mask_n[0]
  PIN cpu_mask_n[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 15.200 1096.000 15.480 1100.000 ;
    END
  END cpu_mask_n[1]
  PIN cpu_mask_n[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 25.780 1096.000 26.060 1100.000 ;
    END
  END cpu_mask_n[2]
  PIN cpu_mask_n[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 35.900 1096.000 36.180 1100.000 ;
    END
  END cpu_mask_n[3]
  PIN cpu_mask_n[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 46.480 1096.000 46.760 1100.000 ;
    END
  END cpu_mask_n[4]
  PIN cpu_mask_n[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 56.600 1096.000 56.880 1100.000 ;
    END
  END cpu_mask_n[5]
  PIN cpu_mask_n[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 67.180 1096.000 67.460 1100.000 ;
    END
  END cpu_mask_n[6]
  PIN cpu_mask_n[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 77.300 1096.000 77.580 1100.000 ;
    END
  END cpu_mask_n[7]
  PIN cpu_wen_e[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 57.160 1099.930 57.760 ;
    END
  END cpu_wen_e[0]
  PIN cpu_wen_e[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 62.600 1099.930 63.200 ;
    END
  END cpu_wen_e[1]
  PIN cpu_wen_n[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 87.880 1096.000 88.160 1100.000 ;
    END
  END cpu_wen_n[0]
  PIN cpu_wen_n[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 98.460 1096.000 98.740 1100.000 ;
    END
  END cpu_wen_n[1]
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 549.720 0.000 550.000 4.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 695.080 0.000 695.360 4.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 709.340 0.000 709.620 4.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 724.060 0.000 724.340 4.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 738.780 0.000 739.060 4.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 753.040 0.000 753.320 4.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 767.760 0.000 768.040 4.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 782.020 0.000 782.300 4.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 796.740 0.000 797.020 4.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 811.460 0.000 811.740 4.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 825.720 0.000 826.000 4.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 563.980 0.000 564.260 4.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 840.440 0.000 840.720 4.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 854.700 0.000 854.980 4.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 869.420 0.000 869.700 4.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 884.140 0.000 884.420 4.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 898.400 0.000 898.680 4.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 913.120 0.000 913.400 4.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 927.380 0.000 927.660 4.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 942.100 0.000 942.380 4.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 956.820 0.000 957.100 4.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 971.080 0.000 971.360 4.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 578.700 0.000 578.980 4.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 985.800 0.000 986.080 4.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1000.060 0.000 1000.340 4.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1014.780 0.000 1015.060 4.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1029.500 0.000 1029.780 4.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1043.760 0.000 1044.040 4.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1058.480 0.000 1058.760 4.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1072.740 0.000 1073.020 4.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1087.460 0.000 1087.740 4.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 593.420 0.000 593.700 4.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 607.680 0.000 607.960 4.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 622.400 0.000 622.680 4.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 636.660 0.000 636.940 4.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 651.380 0.000 651.660 4.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 666.100 0.000 666.380 4.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 680.360 0.000 680.640 4.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 554.320 0.000 554.600 4.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 699.680 0.000 699.960 4.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 714.400 0.000 714.680 4.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 728.660 0.000 728.940 4.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 743.380 0.000 743.660 4.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 758.100 0.000 758.380 4.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 772.360 0.000 772.640 4.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 787.080 0.000 787.360 4.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 801.340 0.000 801.620 4.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 816.060 0.000 816.340 4.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 830.780 0.000 831.060 4.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 569.040 0.000 569.320 4.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 845.040 0.000 845.320 4.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 859.760 0.000 860.040 4.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 874.020 0.000 874.300 4.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 888.740 0.000 889.020 4.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 903.460 0.000 903.740 4.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 917.720 0.000 918.000 4.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 932.440 0.000 932.720 4.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 946.700 0.000 946.980 4.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 961.420 0.000 961.700 4.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 976.140 0.000 976.420 4.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 583.300 0.000 583.580 4.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 990.400 0.000 990.680 4.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1005.120 0.000 1005.400 4.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1019.380 0.000 1019.660 4.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1034.100 0.000 1034.380 4.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1048.820 0.000 1049.100 4.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1063.080 0.000 1063.360 4.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1077.800 0.000 1078.080 4.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1092.060 0.000 1092.340 4.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 598.020 0.000 598.300 4.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 612.740 0.000 613.020 4.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 627.000 0.000 627.280 4.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 641.720 0.000 642.000 4.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 655.980 0.000 656.260 4.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 670.700 0.000 670.980 4.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 685.420 0.000 685.700 4.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 559.380 0.000 559.660 4.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 704.740 0.000 705.020 4.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 719.000 0.000 719.280 4.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 733.720 0.000 734.000 4.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 748.440 0.000 748.720 4.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 762.700 0.000 762.980 4.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 777.420 0.000 777.700 4.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 791.680 0.000 791.960 4.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 806.400 0.000 806.680 4.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 821.120 0.000 821.400 4.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 835.380 0.000 835.660 4.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 573.640 0.000 573.920 4.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 850.100 0.000 850.380 4.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 864.360 0.000 864.640 4.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 879.080 0.000 879.360 4.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 893.800 0.000 894.080 4.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 908.060 0.000 908.340 4.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 922.780 0.000 923.060 4.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 937.040 0.000 937.320 4.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 951.760 0.000 952.040 4.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 966.480 0.000 966.760 4.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 980.740 0.000 981.020 4.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 588.360 0.000 588.640 4.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 995.460 0.000 995.740 4.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1009.720 0.000 1010.000 4.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1024.440 0.000 1024.720 4.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1039.160 0.000 1039.440 4.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1053.420 0.000 1053.700 4.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1068.140 0.000 1068.420 4.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1082.400 0.000 1082.680 4.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1097.120 0.000 1097.400 4.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 603.080 0.000 603.360 4.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 617.340 0.000 617.620 4.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 632.060 0.000 632.340 4.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 646.320 0.000 646.600 4.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 661.040 0.000 661.320 4.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 675.760 0.000 676.040 4.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 690.020 0.000 690.300 4.000 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 515.680 0.000 515.960 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 530.400 0.000 530.680 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 520.740 0.000 521.020 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 535.000 0.000 535.280 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 544.660 0.000 544.940 4.000 ;
    END
  END la_data_out[2]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 525.340 0.000 525.620 4.000 ;
    END
  END la_oen[0]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 540.060 0.000 540.340 4.000 ;
    END
  END la_oen[1]
  PIN one
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 6.840 1099.930 7.440 ;
    END
  END one
  PIN ram_ce
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 11.600 1099.930 12.200 ;
    END
  END ram_ce
  PIN sr0_ce
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 552.200 1099.930 552.800 ;
    END
  END sr0_ce
  PIN sr0_dtr[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 556.960 1099.930 557.560 ;
    END
  END sr0_dtr[0]
  PIN sr0_dtr[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 607.280 1099.930 607.880 ;
    END
  END sr0_dtr[10]
  PIN sr0_dtr[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 612.720 1099.930 613.320 ;
    END
  END sr0_dtr[11]
  PIN sr0_dtr[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 617.480 1099.930 618.080 ;
    END
  END sr0_dtr[12]
  PIN sr0_dtr[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 622.240 1099.930 622.840 ;
    END
  END sr0_dtr[13]
  PIN sr0_dtr[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 627.680 1099.930 628.280 ;
    END
  END sr0_dtr[14]
  PIN sr0_dtr[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 632.440 1099.930 633.040 ;
    END
  END sr0_dtr[15]
  PIN sr0_dtr[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 637.880 1099.930 638.480 ;
    END
  END sr0_dtr[16]
  PIN sr0_dtr[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 642.640 1099.930 643.240 ;
    END
  END sr0_dtr[17]
  PIN sr0_dtr[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 648.080 1099.930 648.680 ;
    END
  END sr0_dtr[18]
  PIN sr0_dtr[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 652.840 1099.930 653.440 ;
    END
  END sr0_dtr[19]
  PIN sr0_dtr[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 561.720 1099.930 562.320 ;
    END
  END sr0_dtr[1]
  PIN sr0_dtr[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 657.600 1099.930 658.200 ;
    END
  END sr0_dtr[20]
  PIN sr0_dtr[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 663.040 1099.930 663.640 ;
    END
  END sr0_dtr[21]
  PIN sr0_dtr[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 667.800 1099.930 668.400 ;
    END
  END sr0_dtr[22]
  PIN sr0_dtr[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 673.240 1099.930 673.840 ;
    END
  END sr0_dtr[23]
  PIN sr0_dtr[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 678.000 1099.930 678.600 ;
    END
  END sr0_dtr[24]
  PIN sr0_dtr[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 682.760 1099.930 683.360 ;
    END
  END sr0_dtr[25]
  PIN sr0_dtr[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 688.200 1099.930 688.800 ;
    END
  END sr0_dtr[26]
  PIN sr0_dtr[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 692.960 1099.930 693.560 ;
    END
  END sr0_dtr[27]
  PIN sr0_dtr[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 698.400 1099.930 699.000 ;
    END
  END sr0_dtr[28]
  PIN sr0_dtr[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 703.160 1099.930 703.760 ;
    END
  END sr0_dtr[29]
  PIN sr0_dtr[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 567.160 1099.930 567.760 ;
    END
  END sr0_dtr[2]
  PIN sr0_dtr[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 708.600 1099.930 709.200 ;
    END
  END sr0_dtr[30]
  PIN sr0_dtr[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 713.360 1099.930 713.960 ;
    END
  END sr0_dtr[31]
  PIN sr0_dtr[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 571.920 1099.930 572.520 ;
    END
  END sr0_dtr[3]
  PIN sr0_dtr[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 577.360 1099.930 577.960 ;
    END
  END sr0_dtr[4]
  PIN sr0_dtr[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 582.120 1099.930 582.720 ;
    END
  END sr0_dtr[5]
  PIN sr0_dtr[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 586.880 1099.930 587.480 ;
    END
  END sr0_dtr[6]
  PIN sr0_dtr[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 592.320 1099.930 592.920 ;
    END
  END sr0_dtr[7]
  PIN sr0_dtr[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 597.080 1099.930 597.680 ;
    END
  END sr0_dtr[8]
  PIN sr0_dtr[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 602.520 1099.930 603.120 ;
    END
  END sr0_dtr[9]
  PIN sr1_ce
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 718.120 1099.930 718.720 ;
    END
  END sr1_ce
  PIN sr1_dtr[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 723.560 1099.930 724.160 ;
    END
  END sr1_dtr[0]
  PIN sr1_dtr[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 773.880 1099.930 774.480 ;
    END
  END sr1_dtr[10]
  PIN sr1_dtr[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 778.640 1099.930 779.240 ;
    END
  END sr1_dtr[11]
  PIN sr1_dtr[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 784.080 1099.930 784.680 ;
    END
  END sr1_dtr[12]
  PIN sr1_dtr[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 788.840 1099.930 789.440 ;
    END
  END sr1_dtr[13]
  PIN sr1_dtr[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 794.280 1099.930 794.880 ;
    END
  END sr1_dtr[14]
  PIN sr1_dtr[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 799.040 1099.930 799.640 ;
    END
  END sr1_dtr[15]
  PIN sr1_dtr[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 804.480 1099.930 805.080 ;
    END
  END sr1_dtr[16]
  PIN sr1_dtr[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 809.240 1099.930 809.840 ;
    END
  END sr1_dtr[17]
  PIN sr1_dtr[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 814.000 1099.930 814.600 ;
    END
  END sr1_dtr[18]
  PIN sr1_dtr[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 819.440 1099.930 820.040 ;
    END
  END sr1_dtr[19]
  PIN sr1_dtr[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 728.320 1099.930 728.920 ;
    END
  END sr1_dtr[1]
  PIN sr1_dtr[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 824.200 1099.930 824.800 ;
    END
  END sr1_dtr[20]
  PIN sr1_dtr[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 829.640 1099.930 830.240 ;
    END
  END sr1_dtr[21]
  PIN sr1_dtr[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 834.400 1099.930 835.000 ;
    END
  END sr1_dtr[22]
  PIN sr1_dtr[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 839.840 1099.930 840.440 ;
    END
  END sr1_dtr[23]
  PIN sr1_dtr[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 844.600 1099.930 845.200 ;
    END
  END sr1_dtr[24]
  PIN sr1_dtr[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 849.360 1099.930 849.960 ;
    END
  END sr1_dtr[25]
  PIN sr1_dtr[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 854.800 1099.930 855.400 ;
    END
  END sr1_dtr[26]
  PIN sr1_dtr[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 859.560 1099.930 860.160 ;
    END
  END sr1_dtr[27]
  PIN sr1_dtr[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 865.000 1099.930 865.600 ;
    END
  END sr1_dtr[28]
  PIN sr1_dtr[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 869.760 1099.930 870.360 ;
    END
  END sr1_dtr[29]
  PIN sr1_dtr[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 733.760 1099.930 734.360 ;
    END
  END sr1_dtr[2]
  PIN sr1_dtr[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 875.200 1099.930 875.800 ;
    END
  END sr1_dtr[30]
  PIN sr1_dtr[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 879.960 1099.930 880.560 ;
    END
  END sr1_dtr[31]
  PIN sr1_dtr[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 738.520 1099.930 739.120 ;
    END
  END sr1_dtr[3]
  PIN sr1_dtr[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 743.960 1099.930 744.560 ;
    END
  END sr1_dtr[4]
  PIN sr1_dtr[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 748.720 1099.930 749.320 ;
    END
  END sr1_dtr[5]
  PIN sr1_dtr[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 753.480 1099.930 754.080 ;
    END
  END sr1_dtr[6]
  PIN sr1_dtr[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 758.920 1099.930 759.520 ;
    END
  END sr1_dtr[7]
  PIN sr1_dtr[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 763.680 1099.930 764.280 ;
    END
  END sr1_dtr[8]
  PIN sr1_dtr[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 769.120 1099.930 769.720 ;
    END
  END sr1_dtr[9]
  PIN srx_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 890.160 1099.930 890.760 ;
    END
  END srx_addr[0]
  PIN srx_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 900.360 1099.930 900.960 ;
    END
  END srx_addr[1]
  PIN srx_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 909.880 1099.930 910.480 ;
    END
  END srx_addr[2]
  PIN srx_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 920.080 1099.930 920.680 ;
    END
  END srx_addr[3]
  PIN srx_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 930.280 1099.930 930.880 ;
    END
  END srx_addr[4]
  PIN srx_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 940.480 1099.930 941.080 ;
    END
  END srx_addr[5]
  PIN srx_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 950.680 1099.930 951.280 ;
    END
  END srx_addr[6]
  PIN srx_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 960.880 1099.930 961.480 ;
    END
  END srx_addr[7]
  PIN srx_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 971.080 1099.930 971.680 ;
    END
  END srx_addr[8]
  PIN srx_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 980.600 1099.930 981.200 ;
    END
  END srx_addr[9]
  PIN srx_dtw[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 894.920 1099.930 895.520 ;
    END
  END srx_dtw[0]
  PIN srx_dtw[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 990.800 1099.930 991.400 ;
    END
  END srx_dtw[10]
  PIN srx_dtw[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 996.240 1099.930 996.840 ;
    END
  END srx_dtw[11]
  PIN srx_dtw[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 1001.000 1099.930 1001.600 ;
    END
  END srx_dtw[12]
  PIN srx_dtw[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 1005.760 1099.930 1006.360 ;
    END
  END srx_dtw[13]
  PIN srx_dtw[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 1011.200 1099.930 1011.800 ;
    END
  END srx_dtw[14]
  PIN srx_dtw[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 1015.960 1099.930 1016.560 ;
    END
  END srx_dtw[15]
  PIN srx_dtw[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 1021.400 1099.930 1022.000 ;
    END
  END srx_dtw[16]
  PIN srx_dtw[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 1026.160 1099.930 1026.760 ;
    END
  END srx_dtw[17]
  PIN srx_dtw[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 1031.600 1099.930 1032.200 ;
    END
  END srx_dtw[18]
  PIN srx_dtw[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 1036.360 1099.930 1036.960 ;
    END
  END srx_dtw[19]
  PIN srx_dtw[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 905.120 1099.930 905.720 ;
    END
  END srx_dtw[1]
  PIN srx_dtw[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 1041.120 1099.930 1041.720 ;
    END
  END srx_dtw[20]
  PIN srx_dtw[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 1046.560 1099.930 1047.160 ;
    END
  END srx_dtw[21]
  PIN srx_dtw[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 1051.320 1099.930 1051.920 ;
    END
  END srx_dtw[22]
  PIN srx_dtw[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 1056.760 1099.930 1057.360 ;
    END
  END srx_dtw[23]
  PIN srx_dtw[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 1061.520 1099.930 1062.120 ;
    END
  END srx_dtw[24]
  PIN srx_dtw[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 1066.960 1099.930 1067.560 ;
    END
  END srx_dtw[25]
  PIN srx_dtw[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 1071.720 1099.930 1072.320 ;
    END
  END srx_dtw[26]
  PIN srx_dtw[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 1076.480 1099.930 1077.080 ;
    END
  END srx_dtw[27]
  PIN srx_dtw[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 1081.920 1099.930 1082.520 ;
    END
  END srx_dtw[28]
  PIN srx_dtw[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 1086.680 1099.930 1087.280 ;
    END
  END srx_dtw[29]
  PIN srx_dtw[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 915.320 1099.930 915.920 ;
    END
  END srx_dtw[2]
  PIN srx_dtw[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 1092.120 1099.930 1092.720 ;
    END
  END srx_dtw[30]
  PIN srx_dtw[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 1096.880 1099.930 1097.480 ;
    END
  END srx_dtw[31]
  PIN srx_dtw[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 925.520 1099.930 926.120 ;
    END
  END srx_dtw[3]
  PIN srx_dtw[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 935.720 1099.930 936.320 ;
    END
  END srx_dtw[4]
  PIN srx_dtw[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 945.240 1099.930 945.840 ;
    END
  END srx_dtw[5]
  PIN srx_dtw[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 955.440 1099.930 956.040 ;
    END
  END srx_dtw[6]
  PIN srx_dtw[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 965.640 1099.930 966.240 ;
    END
  END srx_dtw[7]
  PIN srx_dtw[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 975.840 1099.930 976.440 ;
    END
  END srx_dtw[8]
  PIN srx_dtw[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 986.040 1099.930 986.640 ;
    END
  END srx_dtw[9]
  PIN srx_we
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 884.720 1099.930 885.320 ;
    END
  END srx_we
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.320 0.000 2.600 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.920 0.000 7.200 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 11.980 0.000 12.260 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 31.300 0.000 31.580 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 195.980 0.000 196.260 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 210.240 0.000 210.520 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 224.960 0.000 225.240 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 239.680 0.000 239.960 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 253.940 0.000 254.220 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 268.660 0.000 268.940 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 282.920 0.000 283.200 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 297.640 0.000 297.920 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 312.360 0.000 312.640 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 326.620 0.000 326.900 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 50.620 0.000 50.900 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 341.340 0.000 341.620 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 355.600 0.000 355.880 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 370.320 0.000 370.600 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 385.040 0.000 385.320 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 399.300 0.000 399.580 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 414.020 0.000 414.300 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 428.280 0.000 428.560 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 443.000 0.000 443.280 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 457.720 0.000 458.000 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 471.980 0.000 472.260 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 69.940 0.000 70.220 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 486.700 0.000 486.980 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 500.960 0.000 501.240 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 89.260 0.000 89.540 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 108.580 0.000 108.860 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 123.300 0.000 123.580 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 137.560 0.000 137.840 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 152.280 0.000 152.560 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 167.000 0.000 167.280 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 181.260 0.000 181.540 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 16.580 0.000 16.860 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.900 0.000 36.180 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 200.580 0.000 200.860 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 215.300 0.000 215.580 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 230.020 0.000 230.300 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 244.280 0.000 244.560 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 259.000 0.000 259.280 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 273.260 0.000 273.540 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 287.980 0.000 288.260 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 302.700 0.000 302.980 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 316.960 0.000 317.240 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 331.680 0.000 331.960 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 55.220 0.000 55.500 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 345.940 0.000 346.220 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 360.660 0.000 360.940 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 375.380 0.000 375.660 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 389.640 0.000 389.920 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 404.360 0.000 404.640 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 418.620 0.000 418.900 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 433.340 0.000 433.620 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 448.060 0.000 448.340 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 462.320 0.000 462.600 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 477.040 0.000 477.320 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 74.540 0.000 74.820 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 491.300 0.000 491.580 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 506.020 0.000 506.300 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 94.320 0.000 94.600 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 113.640 0.000 113.920 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 127.900 0.000 128.180 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 142.620 0.000 142.900 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 157.340 0.000 157.620 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 171.600 0.000 171.880 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 186.320 0.000 186.600 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 40.960 0.000 41.240 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 205.640 0.000 205.920 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 219.900 0.000 220.180 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 234.620 0.000 234.900 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 249.340 0.000 249.620 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 263.600 0.000 263.880 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 278.320 0.000 278.600 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 292.580 0.000 292.860 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 307.300 0.000 307.580 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 322.020 0.000 322.300 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 336.280 0.000 336.560 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 60.280 0.000 60.560 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 351.000 0.000 351.280 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 365.260 0.000 365.540 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 379.980 0.000 380.260 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 394.700 0.000 394.980 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 408.960 0.000 409.240 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 423.680 0.000 423.960 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 437.940 0.000 438.220 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 452.660 0.000 452.940 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 467.380 0.000 467.660 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 481.640 0.000 481.920 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 79.600 0.000 79.880 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 496.360 0.000 496.640 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 510.620 0.000 510.900 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 98.920 0.000 99.200 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 118.240 0.000 118.520 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 132.960 0.000 133.240 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 147.220 0.000 147.500 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 161.940 0.000 162.220 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 176.660 0.000 176.940 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 190.920 0.000 191.200 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 45.560 0.000 45.840 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 64.880 0.000 65.160 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 84.660 0.000 84.940 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 103.980 0.000 104.260 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 21.640 0.000 21.920 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.240 0.000 26.520 4.000 ;
    END
  END wbs_we_i
  PIN zero
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 2.080 1099.930 2.680 ;
    END
  END zero
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 20.970 10.640 22.570 1088.240 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.770 10.640 99.370 1088.240 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.450 10.795 1095.045 1088.085 ;
      LAYER met1 ;
        RECT 0.000 7.860 1097.420 1089.320 ;
      LAYER met2 ;
        RECT 0.030 1095.720 4.800 1097.365 ;
        RECT 5.640 1095.720 14.920 1097.365 ;
        RECT 15.760 1095.720 25.500 1097.365 ;
        RECT 26.340 1095.720 35.620 1097.365 ;
        RECT 36.460 1095.720 46.200 1097.365 ;
        RECT 47.040 1095.720 56.320 1097.365 ;
        RECT 57.160 1095.720 66.900 1097.365 ;
        RECT 67.740 1095.720 77.020 1097.365 ;
        RECT 77.860 1095.720 87.600 1097.365 ;
        RECT 88.440 1095.720 98.180 1097.365 ;
        RECT 99.020 1095.720 108.300 1097.365 ;
        RECT 109.140 1095.720 118.880 1097.365 ;
        RECT 119.720 1095.720 129.000 1097.365 ;
        RECT 129.840 1095.720 139.580 1097.365 ;
        RECT 140.420 1095.720 149.700 1097.365 ;
        RECT 150.540 1095.720 160.280 1097.365 ;
        RECT 161.120 1095.720 170.400 1097.365 ;
        RECT 171.240 1095.720 180.980 1097.365 ;
        RECT 181.820 1095.720 191.560 1097.365 ;
        RECT 192.400 1095.720 201.680 1097.365 ;
        RECT 202.520 1095.720 212.260 1097.365 ;
        RECT 213.100 1095.720 222.380 1097.365 ;
        RECT 223.220 1095.720 232.960 1097.365 ;
        RECT 233.800 1095.720 243.080 1097.365 ;
        RECT 243.920 1095.720 253.660 1097.365 ;
        RECT 254.500 1095.720 263.780 1097.365 ;
        RECT 264.620 1095.720 274.360 1097.365 ;
        RECT 275.200 1095.720 284.940 1097.365 ;
        RECT 285.780 1095.720 295.060 1097.365 ;
        RECT 295.900 1095.720 305.640 1097.365 ;
        RECT 306.480 1095.720 315.760 1097.365 ;
        RECT 316.600 1095.720 326.340 1097.365 ;
        RECT 327.180 1095.720 336.460 1097.365 ;
        RECT 337.300 1095.720 347.040 1097.365 ;
        RECT 347.880 1095.720 357.160 1097.365 ;
        RECT 358.000 1095.720 367.740 1097.365 ;
        RECT 368.580 1095.720 378.320 1097.365 ;
        RECT 379.160 1095.720 388.440 1097.365 ;
        RECT 389.280 1095.720 399.020 1097.365 ;
        RECT 399.860 1095.720 409.140 1097.365 ;
        RECT 409.980 1095.720 419.720 1097.365 ;
        RECT 420.560 1095.720 429.840 1097.365 ;
        RECT 430.680 1095.720 440.420 1097.365 ;
        RECT 441.260 1095.720 450.540 1097.365 ;
        RECT 451.380 1095.720 461.120 1097.365 ;
        RECT 461.960 1095.720 471.700 1097.365 ;
        RECT 472.540 1095.720 481.820 1097.365 ;
        RECT 482.660 1095.720 492.400 1097.365 ;
        RECT 493.240 1095.720 502.520 1097.365 ;
        RECT 503.360 1095.720 513.100 1097.365 ;
        RECT 513.940 1095.720 523.220 1097.365 ;
        RECT 524.060 1095.720 533.800 1097.365 ;
        RECT 534.640 1095.720 543.920 1097.365 ;
        RECT 544.760 1095.720 554.500 1097.365 ;
        RECT 555.340 1095.720 565.080 1097.365 ;
        RECT 565.920 1095.720 575.200 1097.365 ;
        RECT 576.040 1095.720 585.780 1097.365 ;
        RECT 586.620 1095.720 595.900 1097.365 ;
        RECT 596.740 1095.720 606.480 1097.365 ;
        RECT 607.320 1095.720 616.600 1097.365 ;
        RECT 617.440 1095.720 627.180 1097.365 ;
        RECT 628.020 1095.720 637.300 1097.365 ;
        RECT 638.140 1095.720 647.880 1097.365 ;
        RECT 648.720 1095.720 658.460 1097.365 ;
        RECT 659.300 1095.720 668.580 1097.365 ;
        RECT 669.420 1095.720 679.160 1097.365 ;
        RECT 680.000 1095.720 689.280 1097.365 ;
        RECT 690.120 1095.720 699.860 1097.365 ;
        RECT 700.700 1095.720 709.980 1097.365 ;
        RECT 710.820 1095.720 720.560 1097.365 ;
        RECT 721.400 1095.720 730.680 1097.365 ;
        RECT 731.520 1095.720 741.260 1097.365 ;
        RECT 742.100 1095.720 751.840 1097.365 ;
        RECT 752.680 1095.720 761.960 1097.365 ;
        RECT 762.800 1095.720 772.540 1097.365 ;
        RECT 773.380 1095.720 782.660 1097.365 ;
        RECT 783.500 1095.720 793.240 1097.365 ;
        RECT 794.080 1095.720 803.360 1097.365 ;
        RECT 804.200 1095.720 813.940 1097.365 ;
        RECT 814.780 1095.720 824.060 1097.365 ;
        RECT 824.900 1095.720 834.640 1097.365 ;
        RECT 835.480 1095.720 845.220 1097.365 ;
        RECT 846.060 1095.720 855.340 1097.365 ;
        RECT 856.180 1095.720 865.920 1097.365 ;
        RECT 866.760 1095.720 876.040 1097.365 ;
        RECT 876.880 1095.720 886.620 1097.365 ;
        RECT 887.460 1095.720 896.740 1097.365 ;
        RECT 897.580 1095.720 907.320 1097.365 ;
        RECT 908.160 1095.720 917.440 1097.365 ;
        RECT 918.280 1095.720 928.020 1097.365 ;
        RECT 928.860 1095.720 938.600 1097.365 ;
        RECT 939.440 1095.720 948.720 1097.365 ;
        RECT 949.560 1095.720 959.300 1097.365 ;
        RECT 960.140 1095.720 969.420 1097.365 ;
        RECT 970.260 1095.720 980.000 1097.365 ;
        RECT 980.840 1095.720 990.120 1097.365 ;
        RECT 990.960 1095.720 1000.700 1097.365 ;
        RECT 1001.540 1095.720 1010.820 1097.365 ;
        RECT 1011.660 1095.720 1021.400 1097.365 ;
        RECT 1022.240 1095.720 1031.980 1097.365 ;
        RECT 1032.820 1095.720 1042.100 1097.365 ;
        RECT 1042.940 1095.720 1052.680 1097.365 ;
        RECT 1053.520 1095.720 1062.800 1097.365 ;
        RECT 1063.640 1095.720 1073.380 1097.365 ;
        RECT 1074.220 1095.720 1083.500 1097.365 ;
        RECT 1084.340 1095.720 1094.080 1097.365 ;
        RECT 1094.920 1095.720 1097.390 1097.365 ;
        RECT 0.030 4.280 1097.390 1095.720 ;
        RECT 0.030 2.195 2.040 4.280 ;
        RECT 2.880 2.195 6.640 4.280 ;
        RECT 7.480 2.195 11.700 4.280 ;
        RECT 12.540 2.195 16.300 4.280 ;
        RECT 17.140 2.195 21.360 4.280 ;
        RECT 22.200 2.195 25.960 4.280 ;
        RECT 26.800 2.195 31.020 4.280 ;
        RECT 31.860 2.195 35.620 4.280 ;
        RECT 36.460 2.195 40.680 4.280 ;
        RECT 41.520 2.195 45.280 4.280 ;
        RECT 46.120 2.195 50.340 4.280 ;
        RECT 51.180 2.195 54.940 4.280 ;
        RECT 55.780 2.195 60.000 4.280 ;
        RECT 60.840 2.195 64.600 4.280 ;
        RECT 65.440 2.195 69.660 4.280 ;
        RECT 70.500 2.195 74.260 4.280 ;
        RECT 75.100 2.195 79.320 4.280 ;
        RECT 80.160 2.195 84.380 4.280 ;
        RECT 85.220 2.195 88.980 4.280 ;
        RECT 89.820 2.195 94.040 4.280 ;
        RECT 94.880 2.195 98.640 4.280 ;
        RECT 99.480 2.195 103.700 4.280 ;
        RECT 104.540 2.195 108.300 4.280 ;
        RECT 109.140 2.195 113.360 4.280 ;
        RECT 114.200 2.195 117.960 4.280 ;
        RECT 118.800 2.195 123.020 4.280 ;
        RECT 123.860 2.195 127.620 4.280 ;
        RECT 128.460 2.195 132.680 4.280 ;
        RECT 133.520 2.195 137.280 4.280 ;
        RECT 138.120 2.195 142.340 4.280 ;
        RECT 143.180 2.195 146.940 4.280 ;
        RECT 147.780 2.195 152.000 4.280 ;
        RECT 152.840 2.195 157.060 4.280 ;
        RECT 157.900 2.195 161.660 4.280 ;
        RECT 162.500 2.195 166.720 4.280 ;
        RECT 167.560 2.195 171.320 4.280 ;
        RECT 172.160 2.195 176.380 4.280 ;
        RECT 177.220 2.195 180.980 4.280 ;
        RECT 181.820 2.195 186.040 4.280 ;
        RECT 186.880 2.195 190.640 4.280 ;
        RECT 191.480 2.195 195.700 4.280 ;
        RECT 196.540 2.195 200.300 4.280 ;
        RECT 201.140 2.195 205.360 4.280 ;
        RECT 206.200 2.195 209.960 4.280 ;
        RECT 210.800 2.195 215.020 4.280 ;
        RECT 215.860 2.195 219.620 4.280 ;
        RECT 220.460 2.195 224.680 4.280 ;
        RECT 225.520 2.195 229.740 4.280 ;
        RECT 230.580 2.195 234.340 4.280 ;
        RECT 235.180 2.195 239.400 4.280 ;
        RECT 240.240 2.195 244.000 4.280 ;
        RECT 244.840 2.195 249.060 4.280 ;
        RECT 249.900 2.195 253.660 4.280 ;
        RECT 254.500 2.195 258.720 4.280 ;
        RECT 259.560 2.195 263.320 4.280 ;
        RECT 264.160 2.195 268.380 4.280 ;
        RECT 269.220 2.195 272.980 4.280 ;
        RECT 273.820 2.195 278.040 4.280 ;
        RECT 278.880 2.195 282.640 4.280 ;
        RECT 283.480 2.195 287.700 4.280 ;
        RECT 288.540 2.195 292.300 4.280 ;
        RECT 293.140 2.195 297.360 4.280 ;
        RECT 298.200 2.195 302.420 4.280 ;
        RECT 303.260 2.195 307.020 4.280 ;
        RECT 307.860 2.195 312.080 4.280 ;
        RECT 312.920 2.195 316.680 4.280 ;
        RECT 317.520 2.195 321.740 4.280 ;
        RECT 322.580 2.195 326.340 4.280 ;
        RECT 327.180 2.195 331.400 4.280 ;
        RECT 332.240 2.195 336.000 4.280 ;
        RECT 336.840 2.195 341.060 4.280 ;
        RECT 341.900 2.195 345.660 4.280 ;
        RECT 346.500 2.195 350.720 4.280 ;
        RECT 351.560 2.195 355.320 4.280 ;
        RECT 356.160 2.195 360.380 4.280 ;
        RECT 361.220 2.195 364.980 4.280 ;
        RECT 365.820 2.195 370.040 4.280 ;
        RECT 370.880 2.195 375.100 4.280 ;
        RECT 375.940 2.195 379.700 4.280 ;
        RECT 380.540 2.195 384.760 4.280 ;
        RECT 385.600 2.195 389.360 4.280 ;
        RECT 390.200 2.195 394.420 4.280 ;
        RECT 395.260 2.195 399.020 4.280 ;
        RECT 399.860 2.195 404.080 4.280 ;
        RECT 404.920 2.195 408.680 4.280 ;
        RECT 409.520 2.195 413.740 4.280 ;
        RECT 414.580 2.195 418.340 4.280 ;
        RECT 419.180 2.195 423.400 4.280 ;
        RECT 424.240 2.195 428.000 4.280 ;
        RECT 428.840 2.195 433.060 4.280 ;
        RECT 433.900 2.195 437.660 4.280 ;
        RECT 438.500 2.195 442.720 4.280 ;
        RECT 443.560 2.195 447.780 4.280 ;
        RECT 448.620 2.195 452.380 4.280 ;
        RECT 453.220 2.195 457.440 4.280 ;
        RECT 458.280 2.195 462.040 4.280 ;
        RECT 462.880 2.195 467.100 4.280 ;
        RECT 467.940 2.195 471.700 4.280 ;
        RECT 472.540 2.195 476.760 4.280 ;
        RECT 477.600 2.195 481.360 4.280 ;
        RECT 482.200 2.195 486.420 4.280 ;
        RECT 487.260 2.195 491.020 4.280 ;
        RECT 491.860 2.195 496.080 4.280 ;
        RECT 496.920 2.195 500.680 4.280 ;
        RECT 501.520 2.195 505.740 4.280 ;
        RECT 506.580 2.195 510.340 4.280 ;
        RECT 511.180 2.195 515.400 4.280 ;
        RECT 516.240 2.195 520.460 4.280 ;
        RECT 521.300 2.195 525.060 4.280 ;
        RECT 525.900 2.195 530.120 4.280 ;
        RECT 530.960 2.195 534.720 4.280 ;
        RECT 535.560 2.195 539.780 4.280 ;
        RECT 540.620 2.195 544.380 4.280 ;
        RECT 545.220 2.195 549.440 4.280 ;
        RECT 550.280 2.195 554.040 4.280 ;
        RECT 554.880 2.195 559.100 4.280 ;
        RECT 559.940 2.195 563.700 4.280 ;
        RECT 564.540 2.195 568.760 4.280 ;
        RECT 569.600 2.195 573.360 4.280 ;
        RECT 574.200 2.195 578.420 4.280 ;
        RECT 579.260 2.195 583.020 4.280 ;
        RECT 583.860 2.195 588.080 4.280 ;
        RECT 588.920 2.195 593.140 4.280 ;
        RECT 593.980 2.195 597.740 4.280 ;
        RECT 598.580 2.195 602.800 4.280 ;
        RECT 603.640 2.195 607.400 4.280 ;
        RECT 608.240 2.195 612.460 4.280 ;
        RECT 613.300 2.195 617.060 4.280 ;
        RECT 617.900 2.195 622.120 4.280 ;
        RECT 622.960 2.195 626.720 4.280 ;
        RECT 627.560 2.195 631.780 4.280 ;
        RECT 632.620 2.195 636.380 4.280 ;
        RECT 637.220 2.195 641.440 4.280 ;
        RECT 642.280 2.195 646.040 4.280 ;
        RECT 646.880 2.195 651.100 4.280 ;
        RECT 651.940 2.195 655.700 4.280 ;
        RECT 656.540 2.195 660.760 4.280 ;
        RECT 661.600 2.195 665.820 4.280 ;
        RECT 666.660 2.195 670.420 4.280 ;
        RECT 671.260 2.195 675.480 4.280 ;
        RECT 676.320 2.195 680.080 4.280 ;
        RECT 680.920 2.195 685.140 4.280 ;
        RECT 685.980 2.195 689.740 4.280 ;
        RECT 690.580 2.195 694.800 4.280 ;
        RECT 695.640 2.195 699.400 4.280 ;
        RECT 700.240 2.195 704.460 4.280 ;
        RECT 705.300 2.195 709.060 4.280 ;
        RECT 709.900 2.195 714.120 4.280 ;
        RECT 714.960 2.195 718.720 4.280 ;
        RECT 719.560 2.195 723.780 4.280 ;
        RECT 724.620 2.195 728.380 4.280 ;
        RECT 729.220 2.195 733.440 4.280 ;
        RECT 734.280 2.195 738.500 4.280 ;
        RECT 739.340 2.195 743.100 4.280 ;
        RECT 743.940 2.195 748.160 4.280 ;
        RECT 749.000 2.195 752.760 4.280 ;
        RECT 753.600 2.195 757.820 4.280 ;
        RECT 758.660 2.195 762.420 4.280 ;
        RECT 763.260 2.195 767.480 4.280 ;
        RECT 768.320 2.195 772.080 4.280 ;
        RECT 772.920 2.195 777.140 4.280 ;
        RECT 777.980 2.195 781.740 4.280 ;
        RECT 782.580 2.195 786.800 4.280 ;
        RECT 787.640 2.195 791.400 4.280 ;
        RECT 792.240 2.195 796.460 4.280 ;
        RECT 797.300 2.195 801.060 4.280 ;
        RECT 801.900 2.195 806.120 4.280 ;
        RECT 806.960 2.195 811.180 4.280 ;
        RECT 812.020 2.195 815.780 4.280 ;
        RECT 816.620 2.195 820.840 4.280 ;
        RECT 821.680 2.195 825.440 4.280 ;
        RECT 826.280 2.195 830.500 4.280 ;
        RECT 831.340 2.195 835.100 4.280 ;
        RECT 835.940 2.195 840.160 4.280 ;
        RECT 841.000 2.195 844.760 4.280 ;
        RECT 845.600 2.195 849.820 4.280 ;
        RECT 850.660 2.195 854.420 4.280 ;
        RECT 855.260 2.195 859.480 4.280 ;
        RECT 860.320 2.195 864.080 4.280 ;
        RECT 864.920 2.195 869.140 4.280 ;
        RECT 869.980 2.195 873.740 4.280 ;
        RECT 874.580 2.195 878.800 4.280 ;
        RECT 879.640 2.195 883.860 4.280 ;
        RECT 884.700 2.195 888.460 4.280 ;
        RECT 889.300 2.195 893.520 4.280 ;
        RECT 894.360 2.195 898.120 4.280 ;
        RECT 898.960 2.195 903.180 4.280 ;
        RECT 904.020 2.195 907.780 4.280 ;
        RECT 908.620 2.195 912.840 4.280 ;
        RECT 913.680 2.195 917.440 4.280 ;
        RECT 918.280 2.195 922.500 4.280 ;
        RECT 923.340 2.195 927.100 4.280 ;
        RECT 927.940 2.195 932.160 4.280 ;
        RECT 933.000 2.195 936.760 4.280 ;
        RECT 937.600 2.195 941.820 4.280 ;
        RECT 942.660 2.195 946.420 4.280 ;
        RECT 947.260 2.195 951.480 4.280 ;
        RECT 952.320 2.195 956.540 4.280 ;
        RECT 957.380 2.195 961.140 4.280 ;
        RECT 961.980 2.195 966.200 4.280 ;
        RECT 967.040 2.195 970.800 4.280 ;
        RECT 971.640 2.195 975.860 4.280 ;
        RECT 976.700 2.195 980.460 4.280 ;
        RECT 981.300 2.195 985.520 4.280 ;
        RECT 986.360 2.195 990.120 4.280 ;
        RECT 990.960 2.195 995.180 4.280 ;
        RECT 996.020 2.195 999.780 4.280 ;
        RECT 1000.620 2.195 1004.840 4.280 ;
        RECT 1005.680 2.195 1009.440 4.280 ;
        RECT 1010.280 2.195 1014.500 4.280 ;
        RECT 1015.340 2.195 1019.100 4.280 ;
        RECT 1019.940 2.195 1024.160 4.280 ;
        RECT 1025.000 2.195 1029.220 4.280 ;
        RECT 1030.060 2.195 1033.820 4.280 ;
        RECT 1034.660 2.195 1038.880 4.280 ;
        RECT 1039.720 2.195 1043.480 4.280 ;
        RECT 1044.320 2.195 1048.540 4.280 ;
        RECT 1049.380 2.195 1053.140 4.280 ;
        RECT 1053.980 2.195 1058.200 4.280 ;
        RECT 1059.040 2.195 1062.800 4.280 ;
        RECT 1063.640 2.195 1067.860 4.280 ;
        RECT 1068.700 2.195 1072.460 4.280 ;
        RECT 1073.300 2.195 1077.520 4.280 ;
        RECT 1078.360 2.195 1082.120 4.280 ;
        RECT 1082.960 2.195 1087.180 4.280 ;
        RECT 1088.020 2.195 1091.780 4.280 ;
        RECT 1092.620 2.195 1096.840 4.280 ;
      LAYER met3 ;
        RECT 5.055 1096.480 1095.530 1097.345 ;
        RECT 5.055 1093.120 1095.930 1096.480 ;
        RECT 5.055 1091.720 1095.530 1093.120 ;
        RECT 5.055 1087.680 1095.930 1091.720 ;
        RECT 5.055 1086.280 1095.530 1087.680 ;
        RECT 5.055 1082.920 1095.930 1086.280 ;
        RECT 5.055 1081.520 1095.530 1082.920 ;
        RECT 5.055 1077.480 1095.930 1081.520 ;
        RECT 5.055 1076.080 1095.530 1077.480 ;
        RECT 5.055 1072.720 1095.930 1076.080 ;
        RECT 5.055 1071.320 1095.530 1072.720 ;
        RECT 5.055 1067.960 1095.930 1071.320 ;
        RECT 5.055 1066.560 1095.530 1067.960 ;
        RECT 5.055 1062.520 1095.930 1066.560 ;
        RECT 5.055 1061.120 1095.530 1062.520 ;
        RECT 5.055 1057.760 1095.930 1061.120 ;
        RECT 5.055 1056.360 1095.530 1057.760 ;
        RECT 5.055 1052.320 1095.930 1056.360 ;
        RECT 5.055 1050.920 1095.530 1052.320 ;
        RECT 5.055 1047.560 1095.930 1050.920 ;
        RECT 5.055 1046.160 1095.530 1047.560 ;
        RECT 5.055 1042.120 1095.930 1046.160 ;
        RECT 5.055 1040.720 1095.530 1042.120 ;
        RECT 5.055 1037.360 1095.930 1040.720 ;
        RECT 5.055 1035.960 1095.530 1037.360 ;
        RECT 5.055 1032.600 1095.930 1035.960 ;
        RECT 5.055 1031.200 1095.530 1032.600 ;
        RECT 5.055 1027.160 1095.930 1031.200 ;
        RECT 5.055 1025.760 1095.530 1027.160 ;
        RECT 5.055 1022.400 1095.930 1025.760 ;
        RECT 5.055 1021.000 1095.530 1022.400 ;
        RECT 5.055 1016.960 1095.930 1021.000 ;
        RECT 5.055 1015.560 1095.530 1016.960 ;
        RECT 5.055 1012.200 1095.930 1015.560 ;
        RECT 5.055 1010.800 1095.530 1012.200 ;
        RECT 5.055 1006.760 1095.930 1010.800 ;
        RECT 5.055 1005.360 1095.530 1006.760 ;
        RECT 5.055 1002.000 1095.930 1005.360 ;
        RECT 5.055 1000.600 1095.530 1002.000 ;
        RECT 5.055 997.240 1095.930 1000.600 ;
        RECT 5.055 995.840 1095.530 997.240 ;
        RECT 5.055 991.800 1095.930 995.840 ;
        RECT 5.055 990.400 1095.530 991.800 ;
        RECT 5.055 987.040 1095.930 990.400 ;
        RECT 5.055 985.640 1095.530 987.040 ;
        RECT 5.055 981.600 1095.930 985.640 ;
        RECT 5.055 980.200 1095.530 981.600 ;
        RECT 5.055 976.840 1095.930 980.200 ;
        RECT 5.055 975.440 1095.530 976.840 ;
        RECT 5.055 972.080 1095.930 975.440 ;
        RECT 5.055 970.680 1095.530 972.080 ;
        RECT 5.055 966.640 1095.930 970.680 ;
        RECT 5.055 965.240 1095.530 966.640 ;
        RECT 5.055 961.880 1095.930 965.240 ;
        RECT 5.055 960.480 1095.530 961.880 ;
        RECT 5.055 956.440 1095.930 960.480 ;
        RECT 5.055 955.040 1095.530 956.440 ;
        RECT 5.055 951.680 1095.930 955.040 ;
        RECT 5.055 950.280 1095.530 951.680 ;
        RECT 5.055 946.240 1095.930 950.280 ;
        RECT 5.055 944.840 1095.530 946.240 ;
        RECT 5.055 941.480 1095.930 944.840 ;
        RECT 5.055 940.080 1095.530 941.480 ;
        RECT 5.055 936.720 1095.930 940.080 ;
        RECT 5.055 935.320 1095.530 936.720 ;
        RECT 5.055 931.280 1095.930 935.320 ;
        RECT 5.055 929.880 1095.530 931.280 ;
        RECT 5.055 926.520 1095.930 929.880 ;
        RECT 5.055 925.120 1095.530 926.520 ;
        RECT 5.055 921.080 1095.930 925.120 ;
        RECT 5.055 919.680 1095.530 921.080 ;
        RECT 5.055 916.320 1095.930 919.680 ;
        RECT 5.055 914.920 1095.530 916.320 ;
        RECT 5.055 910.880 1095.930 914.920 ;
        RECT 5.055 909.480 1095.530 910.880 ;
        RECT 5.055 906.120 1095.930 909.480 ;
        RECT 5.055 904.720 1095.530 906.120 ;
        RECT 5.055 901.360 1095.930 904.720 ;
        RECT 5.055 899.960 1095.530 901.360 ;
        RECT 5.055 895.920 1095.930 899.960 ;
        RECT 5.055 894.520 1095.530 895.920 ;
        RECT 5.055 891.160 1095.930 894.520 ;
        RECT 5.055 889.760 1095.530 891.160 ;
        RECT 5.055 885.720 1095.930 889.760 ;
        RECT 5.055 884.320 1095.530 885.720 ;
        RECT 5.055 880.960 1095.930 884.320 ;
        RECT 5.055 879.560 1095.530 880.960 ;
        RECT 5.055 876.200 1095.930 879.560 ;
        RECT 5.055 874.800 1095.530 876.200 ;
        RECT 5.055 870.760 1095.930 874.800 ;
        RECT 5.055 869.360 1095.530 870.760 ;
        RECT 5.055 866.000 1095.930 869.360 ;
        RECT 5.055 864.600 1095.530 866.000 ;
        RECT 5.055 860.560 1095.930 864.600 ;
        RECT 5.055 859.160 1095.530 860.560 ;
        RECT 5.055 855.800 1095.930 859.160 ;
        RECT 5.055 854.400 1095.530 855.800 ;
        RECT 5.055 850.360 1095.930 854.400 ;
        RECT 5.055 848.960 1095.530 850.360 ;
        RECT 5.055 845.600 1095.930 848.960 ;
        RECT 5.055 844.200 1095.530 845.600 ;
        RECT 5.055 840.840 1095.930 844.200 ;
        RECT 5.055 839.440 1095.530 840.840 ;
        RECT 5.055 835.400 1095.930 839.440 ;
        RECT 5.055 834.000 1095.530 835.400 ;
        RECT 5.055 830.640 1095.930 834.000 ;
        RECT 5.055 829.240 1095.530 830.640 ;
        RECT 5.055 825.200 1095.930 829.240 ;
        RECT 5.055 823.800 1095.530 825.200 ;
        RECT 5.055 820.440 1095.930 823.800 ;
        RECT 5.055 819.040 1095.530 820.440 ;
        RECT 5.055 815.000 1095.930 819.040 ;
        RECT 5.055 813.600 1095.530 815.000 ;
        RECT 5.055 810.240 1095.930 813.600 ;
        RECT 5.055 808.840 1095.530 810.240 ;
        RECT 5.055 805.480 1095.930 808.840 ;
        RECT 5.055 804.080 1095.530 805.480 ;
        RECT 5.055 800.040 1095.930 804.080 ;
        RECT 5.055 798.640 1095.530 800.040 ;
        RECT 5.055 795.280 1095.930 798.640 ;
        RECT 5.055 793.880 1095.530 795.280 ;
        RECT 5.055 789.840 1095.930 793.880 ;
        RECT 5.055 788.440 1095.530 789.840 ;
        RECT 5.055 785.080 1095.930 788.440 ;
        RECT 5.055 783.680 1095.530 785.080 ;
        RECT 5.055 779.640 1095.930 783.680 ;
        RECT 5.055 778.240 1095.530 779.640 ;
        RECT 5.055 774.880 1095.930 778.240 ;
        RECT 5.055 773.480 1095.530 774.880 ;
        RECT 5.055 770.120 1095.930 773.480 ;
        RECT 5.055 768.720 1095.530 770.120 ;
        RECT 5.055 764.680 1095.930 768.720 ;
        RECT 5.055 763.280 1095.530 764.680 ;
        RECT 5.055 759.920 1095.930 763.280 ;
        RECT 5.055 758.520 1095.530 759.920 ;
        RECT 5.055 754.480 1095.930 758.520 ;
        RECT 5.055 753.080 1095.530 754.480 ;
        RECT 5.055 749.720 1095.930 753.080 ;
        RECT 5.055 748.320 1095.530 749.720 ;
        RECT 5.055 744.960 1095.930 748.320 ;
        RECT 5.055 743.560 1095.530 744.960 ;
        RECT 5.055 739.520 1095.930 743.560 ;
        RECT 5.055 738.120 1095.530 739.520 ;
        RECT 5.055 734.760 1095.930 738.120 ;
        RECT 5.055 733.360 1095.530 734.760 ;
        RECT 5.055 729.320 1095.930 733.360 ;
        RECT 5.055 727.920 1095.530 729.320 ;
        RECT 5.055 724.560 1095.930 727.920 ;
        RECT 5.055 723.160 1095.530 724.560 ;
        RECT 5.055 719.120 1095.930 723.160 ;
        RECT 5.055 717.720 1095.530 719.120 ;
        RECT 5.055 714.360 1095.930 717.720 ;
        RECT 5.055 712.960 1095.530 714.360 ;
        RECT 5.055 709.600 1095.930 712.960 ;
        RECT 5.055 708.200 1095.530 709.600 ;
        RECT 5.055 704.160 1095.930 708.200 ;
        RECT 5.055 702.760 1095.530 704.160 ;
        RECT 5.055 699.400 1095.930 702.760 ;
        RECT 5.055 698.000 1095.530 699.400 ;
        RECT 5.055 693.960 1095.930 698.000 ;
        RECT 5.055 692.560 1095.530 693.960 ;
        RECT 5.055 689.200 1095.930 692.560 ;
        RECT 5.055 687.800 1095.530 689.200 ;
        RECT 5.055 683.760 1095.930 687.800 ;
        RECT 5.055 682.360 1095.530 683.760 ;
        RECT 5.055 679.000 1095.930 682.360 ;
        RECT 5.055 677.600 1095.530 679.000 ;
        RECT 5.055 674.240 1095.930 677.600 ;
        RECT 5.055 672.840 1095.530 674.240 ;
        RECT 5.055 668.800 1095.930 672.840 ;
        RECT 5.055 667.400 1095.530 668.800 ;
        RECT 5.055 664.040 1095.930 667.400 ;
        RECT 5.055 662.640 1095.530 664.040 ;
        RECT 5.055 658.600 1095.930 662.640 ;
        RECT 5.055 657.200 1095.530 658.600 ;
        RECT 5.055 653.840 1095.930 657.200 ;
        RECT 5.055 652.440 1095.530 653.840 ;
        RECT 5.055 649.080 1095.930 652.440 ;
        RECT 5.055 647.680 1095.530 649.080 ;
        RECT 5.055 643.640 1095.930 647.680 ;
        RECT 5.055 642.240 1095.530 643.640 ;
        RECT 5.055 638.880 1095.930 642.240 ;
        RECT 5.055 637.480 1095.530 638.880 ;
        RECT 5.055 633.440 1095.930 637.480 ;
        RECT 5.055 632.040 1095.530 633.440 ;
        RECT 5.055 628.680 1095.930 632.040 ;
        RECT 5.055 627.280 1095.530 628.680 ;
        RECT 5.055 623.240 1095.930 627.280 ;
        RECT 5.055 621.840 1095.530 623.240 ;
        RECT 5.055 618.480 1095.930 621.840 ;
        RECT 5.055 617.080 1095.530 618.480 ;
        RECT 5.055 613.720 1095.930 617.080 ;
        RECT 5.055 612.320 1095.530 613.720 ;
        RECT 5.055 608.280 1095.930 612.320 ;
        RECT 5.055 606.880 1095.530 608.280 ;
        RECT 5.055 603.520 1095.930 606.880 ;
        RECT 5.055 602.120 1095.530 603.520 ;
        RECT 5.055 598.080 1095.930 602.120 ;
        RECT 5.055 596.680 1095.530 598.080 ;
        RECT 5.055 593.320 1095.930 596.680 ;
        RECT 5.055 591.920 1095.530 593.320 ;
        RECT 5.055 587.880 1095.930 591.920 ;
        RECT 5.055 586.480 1095.530 587.880 ;
        RECT 5.055 583.120 1095.930 586.480 ;
        RECT 5.055 581.720 1095.530 583.120 ;
        RECT 5.055 578.360 1095.930 581.720 ;
        RECT 5.055 576.960 1095.530 578.360 ;
        RECT 5.055 572.920 1095.930 576.960 ;
        RECT 5.055 571.520 1095.530 572.920 ;
        RECT 5.055 568.160 1095.930 571.520 ;
        RECT 5.055 566.760 1095.530 568.160 ;
        RECT 5.055 562.720 1095.930 566.760 ;
        RECT 5.055 561.320 1095.530 562.720 ;
        RECT 5.055 557.960 1095.930 561.320 ;
        RECT 5.055 556.560 1095.530 557.960 ;
        RECT 5.055 553.200 1095.930 556.560 ;
        RECT 5.055 551.800 1095.530 553.200 ;
        RECT 5.055 547.760 1095.930 551.800 ;
        RECT 5.055 546.360 1095.530 547.760 ;
        RECT 5.055 543.000 1095.930 546.360 ;
        RECT 5.055 541.600 1095.530 543.000 ;
        RECT 5.055 537.560 1095.930 541.600 ;
        RECT 5.055 536.160 1095.530 537.560 ;
        RECT 5.055 532.800 1095.930 536.160 ;
        RECT 5.055 531.400 1095.530 532.800 ;
        RECT 5.055 527.360 1095.930 531.400 ;
        RECT 5.055 525.960 1095.530 527.360 ;
        RECT 5.055 522.600 1095.930 525.960 ;
        RECT 5.055 521.200 1095.530 522.600 ;
        RECT 5.055 517.840 1095.930 521.200 ;
        RECT 5.055 516.440 1095.530 517.840 ;
        RECT 5.055 512.400 1095.930 516.440 ;
        RECT 5.055 511.000 1095.530 512.400 ;
        RECT 5.055 507.640 1095.930 511.000 ;
        RECT 5.055 506.240 1095.530 507.640 ;
        RECT 5.055 502.200 1095.930 506.240 ;
        RECT 5.055 500.800 1095.530 502.200 ;
        RECT 5.055 497.440 1095.930 500.800 ;
        RECT 5.055 496.040 1095.530 497.440 ;
        RECT 5.055 492.000 1095.930 496.040 ;
        RECT 5.055 490.600 1095.530 492.000 ;
        RECT 5.055 487.240 1095.930 490.600 ;
        RECT 5.055 485.840 1095.530 487.240 ;
        RECT 5.055 482.480 1095.930 485.840 ;
        RECT 5.055 481.080 1095.530 482.480 ;
        RECT 5.055 477.040 1095.930 481.080 ;
        RECT 5.055 475.640 1095.530 477.040 ;
        RECT 5.055 472.280 1095.930 475.640 ;
        RECT 5.055 470.880 1095.530 472.280 ;
        RECT 5.055 466.840 1095.930 470.880 ;
        RECT 5.055 465.440 1095.530 466.840 ;
        RECT 5.055 462.080 1095.930 465.440 ;
        RECT 5.055 460.680 1095.530 462.080 ;
        RECT 5.055 456.640 1095.930 460.680 ;
        RECT 5.055 455.240 1095.530 456.640 ;
        RECT 5.055 451.880 1095.930 455.240 ;
        RECT 5.055 450.480 1095.530 451.880 ;
        RECT 5.055 447.120 1095.930 450.480 ;
        RECT 5.055 445.720 1095.530 447.120 ;
        RECT 5.055 441.680 1095.930 445.720 ;
        RECT 5.055 440.280 1095.530 441.680 ;
        RECT 5.055 436.920 1095.930 440.280 ;
        RECT 5.055 435.520 1095.530 436.920 ;
        RECT 5.055 431.480 1095.930 435.520 ;
        RECT 5.055 430.080 1095.530 431.480 ;
        RECT 5.055 426.720 1095.930 430.080 ;
        RECT 5.055 425.320 1095.530 426.720 ;
        RECT 5.055 421.960 1095.930 425.320 ;
        RECT 5.055 420.560 1095.530 421.960 ;
        RECT 5.055 416.520 1095.930 420.560 ;
        RECT 5.055 415.120 1095.530 416.520 ;
        RECT 5.055 411.760 1095.930 415.120 ;
        RECT 5.055 410.360 1095.530 411.760 ;
        RECT 5.055 406.320 1095.930 410.360 ;
        RECT 5.055 404.920 1095.530 406.320 ;
        RECT 5.055 401.560 1095.930 404.920 ;
        RECT 5.055 400.160 1095.530 401.560 ;
        RECT 5.055 396.120 1095.930 400.160 ;
        RECT 5.055 394.720 1095.530 396.120 ;
        RECT 5.055 391.360 1095.930 394.720 ;
        RECT 5.055 389.960 1095.530 391.360 ;
        RECT 5.055 386.600 1095.930 389.960 ;
        RECT 5.055 385.200 1095.530 386.600 ;
        RECT 5.055 381.160 1095.930 385.200 ;
        RECT 5.055 379.760 1095.530 381.160 ;
        RECT 5.055 376.400 1095.930 379.760 ;
        RECT 5.055 375.000 1095.530 376.400 ;
        RECT 5.055 370.960 1095.930 375.000 ;
        RECT 5.055 369.560 1095.530 370.960 ;
        RECT 5.055 366.200 1095.930 369.560 ;
        RECT 5.055 364.800 1095.530 366.200 ;
        RECT 5.055 360.760 1095.930 364.800 ;
        RECT 5.055 359.360 1095.530 360.760 ;
        RECT 5.055 356.000 1095.930 359.360 ;
        RECT 5.055 354.600 1095.530 356.000 ;
        RECT 5.055 351.240 1095.930 354.600 ;
        RECT 5.055 349.840 1095.530 351.240 ;
        RECT 5.055 345.800 1095.930 349.840 ;
        RECT 5.055 344.400 1095.530 345.800 ;
        RECT 5.055 341.040 1095.930 344.400 ;
        RECT 5.055 339.640 1095.530 341.040 ;
        RECT 5.055 335.600 1095.930 339.640 ;
        RECT 5.055 334.200 1095.530 335.600 ;
        RECT 5.055 330.840 1095.930 334.200 ;
        RECT 5.055 329.440 1095.530 330.840 ;
        RECT 5.055 326.080 1095.930 329.440 ;
        RECT 5.055 324.680 1095.530 326.080 ;
        RECT 5.055 320.640 1095.930 324.680 ;
        RECT 5.055 319.240 1095.530 320.640 ;
        RECT 5.055 315.880 1095.930 319.240 ;
        RECT 5.055 314.480 1095.530 315.880 ;
        RECT 5.055 310.440 1095.930 314.480 ;
        RECT 5.055 309.040 1095.530 310.440 ;
        RECT 5.055 305.680 1095.930 309.040 ;
        RECT 5.055 304.280 1095.530 305.680 ;
        RECT 5.055 300.240 1095.930 304.280 ;
        RECT 5.055 298.840 1095.530 300.240 ;
        RECT 5.055 295.480 1095.930 298.840 ;
        RECT 5.055 294.080 1095.530 295.480 ;
        RECT 5.055 290.720 1095.930 294.080 ;
        RECT 5.055 289.320 1095.530 290.720 ;
        RECT 5.055 285.280 1095.930 289.320 ;
        RECT 5.055 283.880 1095.530 285.280 ;
        RECT 5.055 280.520 1095.930 283.880 ;
        RECT 5.055 279.120 1095.530 280.520 ;
        RECT 5.055 275.080 1095.930 279.120 ;
        RECT 5.055 273.680 1095.530 275.080 ;
        RECT 5.055 270.320 1095.930 273.680 ;
        RECT 5.055 268.920 1095.530 270.320 ;
        RECT 5.055 264.880 1095.930 268.920 ;
        RECT 5.055 263.480 1095.530 264.880 ;
        RECT 5.055 260.120 1095.930 263.480 ;
        RECT 5.055 258.720 1095.530 260.120 ;
        RECT 5.055 255.360 1095.930 258.720 ;
        RECT 5.055 253.960 1095.530 255.360 ;
        RECT 5.055 249.920 1095.930 253.960 ;
        RECT 5.055 248.520 1095.530 249.920 ;
        RECT 5.055 245.160 1095.930 248.520 ;
        RECT 5.055 243.760 1095.530 245.160 ;
        RECT 5.055 239.720 1095.930 243.760 ;
        RECT 5.055 238.320 1095.530 239.720 ;
        RECT 5.055 234.960 1095.930 238.320 ;
        RECT 5.055 233.560 1095.530 234.960 ;
        RECT 5.055 229.520 1095.930 233.560 ;
        RECT 5.055 228.120 1095.530 229.520 ;
        RECT 5.055 224.760 1095.930 228.120 ;
        RECT 5.055 223.360 1095.530 224.760 ;
        RECT 5.055 220.000 1095.930 223.360 ;
        RECT 5.055 218.600 1095.530 220.000 ;
        RECT 5.055 214.560 1095.930 218.600 ;
        RECT 5.055 213.160 1095.530 214.560 ;
        RECT 5.055 209.800 1095.930 213.160 ;
        RECT 5.055 208.400 1095.530 209.800 ;
        RECT 5.055 204.360 1095.930 208.400 ;
        RECT 5.055 202.960 1095.530 204.360 ;
        RECT 5.055 199.600 1095.930 202.960 ;
        RECT 5.055 198.200 1095.530 199.600 ;
        RECT 5.055 194.840 1095.930 198.200 ;
        RECT 5.055 193.440 1095.530 194.840 ;
        RECT 5.055 189.400 1095.930 193.440 ;
        RECT 5.055 188.000 1095.530 189.400 ;
        RECT 5.055 184.640 1095.930 188.000 ;
        RECT 5.055 183.240 1095.530 184.640 ;
        RECT 5.055 179.200 1095.930 183.240 ;
        RECT 5.055 177.800 1095.530 179.200 ;
        RECT 5.055 174.440 1095.930 177.800 ;
        RECT 5.055 173.040 1095.530 174.440 ;
        RECT 5.055 169.000 1095.930 173.040 ;
        RECT 5.055 167.600 1095.530 169.000 ;
        RECT 5.055 164.240 1095.930 167.600 ;
        RECT 5.055 162.840 1095.530 164.240 ;
        RECT 5.055 159.480 1095.930 162.840 ;
        RECT 5.055 158.080 1095.530 159.480 ;
        RECT 5.055 154.040 1095.930 158.080 ;
        RECT 5.055 152.640 1095.530 154.040 ;
        RECT 5.055 149.280 1095.930 152.640 ;
        RECT 5.055 147.880 1095.530 149.280 ;
        RECT 5.055 143.840 1095.930 147.880 ;
        RECT 5.055 142.440 1095.530 143.840 ;
        RECT 5.055 139.080 1095.930 142.440 ;
        RECT 5.055 137.680 1095.530 139.080 ;
        RECT 5.055 133.640 1095.930 137.680 ;
        RECT 5.055 132.240 1095.530 133.640 ;
        RECT 5.055 128.880 1095.930 132.240 ;
        RECT 5.055 127.480 1095.530 128.880 ;
        RECT 5.055 124.120 1095.930 127.480 ;
        RECT 5.055 122.720 1095.530 124.120 ;
        RECT 5.055 118.680 1095.930 122.720 ;
        RECT 5.055 117.280 1095.530 118.680 ;
        RECT 5.055 113.920 1095.930 117.280 ;
        RECT 5.055 112.520 1095.530 113.920 ;
        RECT 5.055 108.480 1095.930 112.520 ;
        RECT 5.055 107.080 1095.530 108.480 ;
        RECT 5.055 103.720 1095.930 107.080 ;
        RECT 5.055 102.320 1095.530 103.720 ;
        RECT 5.055 98.960 1095.930 102.320 ;
        RECT 5.055 97.560 1095.530 98.960 ;
        RECT 5.055 93.520 1095.930 97.560 ;
        RECT 5.055 92.120 1095.530 93.520 ;
        RECT 5.055 88.760 1095.930 92.120 ;
        RECT 5.055 87.360 1095.530 88.760 ;
        RECT 5.055 83.320 1095.930 87.360 ;
        RECT 5.055 81.920 1095.530 83.320 ;
        RECT 5.055 78.560 1095.930 81.920 ;
        RECT 5.055 77.160 1095.530 78.560 ;
        RECT 5.055 73.120 1095.930 77.160 ;
        RECT 5.055 71.720 1095.530 73.120 ;
        RECT 5.055 68.360 1095.930 71.720 ;
        RECT 5.055 66.960 1095.530 68.360 ;
        RECT 5.055 63.600 1095.930 66.960 ;
        RECT 5.055 62.200 1095.530 63.600 ;
        RECT 5.055 58.160 1095.930 62.200 ;
        RECT 5.055 56.760 1095.530 58.160 ;
        RECT 5.055 53.400 1095.930 56.760 ;
        RECT 5.055 52.000 1095.530 53.400 ;
        RECT 5.055 47.960 1095.930 52.000 ;
        RECT 5.055 46.560 1095.530 47.960 ;
        RECT 5.055 43.200 1095.930 46.560 ;
        RECT 5.055 41.800 1095.530 43.200 ;
        RECT 5.055 37.760 1095.930 41.800 ;
        RECT 5.055 36.360 1095.530 37.760 ;
        RECT 5.055 33.000 1095.930 36.360 ;
        RECT 5.055 31.600 1095.530 33.000 ;
        RECT 5.055 28.240 1095.930 31.600 ;
        RECT 5.055 26.840 1095.530 28.240 ;
        RECT 5.055 22.800 1095.930 26.840 ;
        RECT 5.055 21.400 1095.530 22.800 ;
        RECT 5.055 18.040 1095.930 21.400 ;
        RECT 5.055 16.640 1095.530 18.040 ;
        RECT 5.055 12.600 1095.930 16.640 ;
        RECT 5.055 11.200 1095.530 12.600 ;
        RECT 5.055 7.840 1095.930 11.200 ;
        RECT 5.055 6.440 1095.530 7.840 ;
        RECT 5.055 3.080 1095.930 6.440 ;
        RECT 5.055 2.215 1095.530 3.080 ;
      LAYER met4 ;
        RECT 25.065 10.640 97.370 1088.240 ;
        RECT 99.770 10.640 1088.915 1088.240 ;
  END
END hs32_core1
END LIBRARY

