magic
tech sky130A
magscale 1 2
timestamp 1608368632
<< obsli1 >>
rect 1090 2159 219009 217617
<< obsm1 >>
rect 0 1572 219484 217864
<< metal2 >>
rect 1016 219200 1072 220000
rect 3040 219200 3096 220000
rect 5156 219200 5212 220000
rect 7180 219200 7236 220000
rect 9296 219200 9352 220000
rect 11320 219200 11376 220000
rect 13436 219200 13492 220000
rect 15460 219200 15516 220000
rect 17576 219200 17632 220000
rect 19692 219200 19748 220000
rect 21716 219200 21772 220000
rect 23832 219200 23888 220000
rect 25856 219200 25912 220000
rect 27972 219200 28028 220000
rect 29996 219200 30052 220000
rect 32112 219200 32168 220000
rect 34136 219200 34192 220000
rect 36252 219200 36308 220000
rect 38368 219200 38424 220000
rect 40392 219200 40448 220000
rect 42508 219200 42564 220000
rect 44532 219200 44588 220000
rect 46648 219200 46704 220000
rect 48672 219200 48728 220000
rect 50788 219200 50844 220000
rect 52812 219200 52868 220000
rect 54928 219200 54984 220000
rect 57044 219200 57100 220000
rect 59068 219200 59124 220000
rect 61184 219200 61240 220000
rect 63208 219200 63264 220000
rect 65324 219200 65380 220000
rect 67348 219200 67404 220000
rect 69464 219200 69520 220000
rect 71488 219200 71544 220000
rect 73604 219200 73660 220000
rect 75720 219200 75776 220000
rect 77744 219200 77800 220000
rect 79860 219200 79916 220000
rect 81884 219200 81940 220000
rect 84000 219200 84056 220000
rect 86024 219200 86080 220000
rect 88140 219200 88196 220000
rect 90164 219200 90220 220000
rect 92280 219200 92336 220000
rect 94396 219200 94452 220000
rect 96420 219200 96476 220000
rect 98536 219200 98592 220000
rect 100560 219200 100616 220000
rect 102676 219200 102732 220000
rect 104700 219200 104756 220000
rect 106816 219200 106872 220000
rect 108840 219200 108896 220000
rect 110956 219200 111012 220000
rect 113072 219200 113128 220000
rect 115096 219200 115152 220000
rect 117212 219200 117268 220000
rect 119236 219200 119292 220000
rect 121352 219200 121408 220000
rect 123376 219200 123432 220000
rect 125492 219200 125548 220000
rect 127516 219200 127572 220000
rect 129632 219200 129688 220000
rect 131748 219200 131804 220000
rect 133772 219200 133828 220000
rect 135888 219200 135944 220000
rect 137912 219200 137968 220000
rect 140028 219200 140084 220000
rect 142052 219200 142108 220000
rect 144168 219200 144224 220000
rect 146192 219200 146248 220000
rect 148308 219200 148364 220000
rect 150424 219200 150480 220000
rect 152448 219200 152504 220000
rect 154564 219200 154620 220000
rect 156588 219200 156644 220000
rect 158704 219200 158760 220000
rect 160728 219200 160784 220000
rect 162844 219200 162900 220000
rect 164868 219200 164924 220000
rect 166984 219200 167040 220000
rect 169100 219200 169156 220000
rect 171124 219200 171180 220000
rect 173240 219200 173296 220000
rect 175264 219200 175320 220000
rect 177380 219200 177436 220000
rect 179404 219200 179460 220000
rect 181520 219200 181576 220000
rect 183544 219200 183600 220000
rect 185660 219200 185716 220000
rect 187776 219200 187832 220000
rect 189800 219200 189856 220000
rect 191916 219200 191972 220000
rect 193940 219200 193996 220000
rect 196056 219200 196112 220000
rect 198080 219200 198136 220000
rect 200196 219200 200252 220000
rect 202220 219200 202276 220000
rect 204336 219200 204392 220000
rect 206452 219200 206508 220000
rect 208476 219200 208532 220000
rect 210592 219200 210648 220000
rect 212616 219200 212672 220000
rect 214732 219200 214788 220000
rect 216756 219200 216812 220000
rect 218872 219200 218928 220000
rect 464 0 520 800
rect 1384 0 1440 800
rect 2396 0 2452 800
rect 3316 0 3372 800
rect 4328 0 4384 800
rect 5248 0 5304 800
rect 6260 0 6316 800
rect 7180 0 7236 800
rect 8192 0 8248 800
rect 9112 0 9168 800
rect 10124 0 10180 800
rect 11044 0 11100 800
rect 12056 0 12112 800
rect 12976 0 13032 800
rect 13988 0 14044 800
rect 14908 0 14964 800
rect 15920 0 15976 800
rect 16932 0 16988 800
rect 17852 0 17908 800
rect 18864 0 18920 800
rect 19784 0 19840 800
rect 20796 0 20852 800
rect 21716 0 21772 800
rect 22728 0 22784 800
rect 23648 0 23704 800
rect 24660 0 24716 800
rect 25580 0 25636 800
rect 26592 0 26648 800
rect 27512 0 27568 800
rect 28524 0 28580 800
rect 29444 0 29500 800
rect 30456 0 30512 800
rect 31468 0 31524 800
rect 32388 0 32444 800
rect 33400 0 33456 800
rect 34320 0 34376 800
rect 35332 0 35388 800
rect 36252 0 36308 800
rect 37264 0 37320 800
rect 38184 0 38240 800
rect 39196 0 39252 800
rect 40116 0 40172 800
rect 41128 0 41184 800
rect 42048 0 42104 800
rect 43060 0 43116 800
rect 43980 0 44036 800
rect 44992 0 45048 800
rect 46004 0 46060 800
rect 46924 0 46980 800
rect 47936 0 47992 800
rect 48856 0 48912 800
rect 49868 0 49924 800
rect 50788 0 50844 800
rect 51800 0 51856 800
rect 52720 0 52776 800
rect 53732 0 53788 800
rect 54652 0 54708 800
rect 55664 0 55720 800
rect 56584 0 56640 800
rect 57596 0 57652 800
rect 58516 0 58572 800
rect 59528 0 59584 800
rect 60540 0 60596 800
rect 61460 0 61516 800
rect 62472 0 62528 800
rect 63392 0 63448 800
rect 64404 0 64460 800
rect 65324 0 65380 800
rect 66336 0 66392 800
rect 67256 0 67312 800
rect 68268 0 68324 800
rect 69188 0 69244 800
rect 70200 0 70256 800
rect 71120 0 71176 800
rect 72132 0 72188 800
rect 73052 0 73108 800
rect 74064 0 74120 800
rect 75076 0 75132 800
rect 75996 0 76052 800
rect 77008 0 77064 800
rect 77928 0 77984 800
rect 78940 0 78996 800
rect 79860 0 79916 800
rect 80872 0 80928 800
rect 81792 0 81848 800
rect 82804 0 82860 800
rect 83724 0 83780 800
rect 84736 0 84792 800
rect 85656 0 85712 800
rect 86668 0 86724 800
rect 87588 0 87644 800
rect 88600 0 88656 800
rect 89612 0 89668 800
rect 90532 0 90588 800
rect 91544 0 91600 800
rect 92464 0 92520 800
rect 93476 0 93532 800
rect 94396 0 94452 800
rect 95408 0 95464 800
rect 96328 0 96384 800
rect 97340 0 97396 800
rect 98260 0 98316 800
rect 99272 0 99328 800
rect 100192 0 100248 800
rect 101204 0 101260 800
rect 102124 0 102180 800
rect 103136 0 103192 800
rect 104148 0 104204 800
rect 105068 0 105124 800
rect 106080 0 106136 800
rect 107000 0 107056 800
rect 108012 0 108068 800
rect 108932 0 108988 800
rect 109944 0 110000 800
rect 110864 0 110920 800
rect 111876 0 111932 800
rect 112796 0 112852 800
rect 113808 0 113864 800
rect 114728 0 114784 800
rect 115740 0 115796 800
rect 116660 0 116716 800
rect 117672 0 117728 800
rect 118684 0 118740 800
rect 119604 0 119660 800
rect 120616 0 120672 800
rect 121536 0 121592 800
rect 122548 0 122604 800
rect 123468 0 123524 800
rect 124480 0 124536 800
rect 125400 0 125456 800
rect 126412 0 126468 800
rect 127332 0 127388 800
rect 128344 0 128400 800
rect 129264 0 129320 800
rect 130276 0 130332 800
rect 131196 0 131252 800
rect 132208 0 132264 800
rect 133220 0 133276 800
rect 134140 0 134196 800
rect 135152 0 135208 800
rect 136072 0 136128 800
rect 137084 0 137140 800
rect 138004 0 138060 800
rect 139016 0 139072 800
rect 139936 0 139992 800
rect 140948 0 141004 800
rect 141868 0 141924 800
rect 142880 0 142936 800
rect 143800 0 143856 800
rect 144812 0 144868 800
rect 145732 0 145788 800
rect 146744 0 146800 800
rect 147756 0 147812 800
rect 148676 0 148732 800
rect 149688 0 149744 800
rect 150608 0 150664 800
rect 151620 0 151676 800
rect 152540 0 152596 800
rect 153552 0 153608 800
rect 154472 0 154528 800
rect 155484 0 155540 800
rect 156404 0 156460 800
rect 157416 0 157472 800
rect 158336 0 158392 800
rect 159348 0 159404 800
rect 160268 0 160324 800
rect 161280 0 161336 800
rect 162292 0 162348 800
rect 163212 0 163268 800
rect 164224 0 164280 800
rect 165144 0 165200 800
rect 166156 0 166212 800
rect 167076 0 167132 800
rect 168088 0 168144 800
rect 169008 0 169064 800
rect 170020 0 170076 800
rect 170940 0 170996 800
rect 171952 0 172008 800
rect 172872 0 172928 800
rect 173884 0 173940 800
rect 174804 0 174860 800
rect 175816 0 175872 800
rect 176828 0 176884 800
rect 177748 0 177804 800
rect 178760 0 178816 800
rect 179680 0 179736 800
rect 180692 0 180748 800
rect 181612 0 181668 800
rect 182624 0 182680 800
rect 183544 0 183600 800
rect 184556 0 184612 800
rect 185476 0 185532 800
rect 186488 0 186544 800
rect 187408 0 187464 800
rect 188420 0 188476 800
rect 189340 0 189396 800
rect 190352 0 190408 800
rect 191364 0 191420 800
rect 192284 0 192340 800
rect 193296 0 193352 800
rect 194216 0 194272 800
rect 195228 0 195284 800
rect 196148 0 196204 800
rect 197160 0 197216 800
rect 198080 0 198136 800
rect 199092 0 199148 800
rect 200012 0 200068 800
rect 201024 0 201080 800
rect 201944 0 202000 800
rect 202956 0 203012 800
rect 203876 0 203932 800
rect 204888 0 204944 800
rect 205900 0 205956 800
rect 206820 0 206876 800
rect 207832 0 207888 800
rect 208752 0 208808 800
rect 209764 0 209820 800
rect 210684 0 210740 800
rect 211696 0 211752 800
rect 212616 0 212672 800
rect 213628 0 213684 800
rect 214548 0 214604 800
rect 215560 0 215616 800
rect 216480 0 216536 800
rect 217492 0 217548 800
rect 218412 0 218468 800
rect 219424 0 219480 800
<< obsm2 >>
rect 6 219144 960 219473
rect 1128 219144 2984 219473
rect 3152 219144 5100 219473
rect 5268 219144 7124 219473
rect 7292 219144 9240 219473
rect 9408 219144 11264 219473
rect 11432 219144 13380 219473
rect 13548 219144 15404 219473
rect 15572 219144 17520 219473
rect 17688 219144 19636 219473
rect 19804 219144 21660 219473
rect 21828 219144 23776 219473
rect 23944 219144 25800 219473
rect 25968 219144 27916 219473
rect 28084 219144 29940 219473
rect 30108 219144 32056 219473
rect 32224 219144 34080 219473
rect 34248 219144 36196 219473
rect 36364 219144 38312 219473
rect 38480 219144 40336 219473
rect 40504 219144 42452 219473
rect 42620 219144 44476 219473
rect 44644 219144 46592 219473
rect 46760 219144 48616 219473
rect 48784 219144 50732 219473
rect 50900 219144 52756 219473
rect 52924 219144 54872 219473
rect 55040 219144 56988 219473
rect 57156 219144 59012 219473
rect 59180 219144 61128 219473
rect 61296 219144 63152 219473
rect 63320 219144 65268 219473
rect 65436 219144 67292 219473
rect 67460 219144 69408 219473
rect 69576 219144 71432 219473
rect 71600 219144 73548 219473
rect 73716 219144 75664 219473
rect 75832 219144 77688 219473
rect 77856 219144 79804 219473
rect 79972 219144 81828 219473
rect 81996 219144 83944 219473
rect 84112 219144 85968 219473
rect 86136 219144 88084 219473
rect 88252 219144 90108 219473
rect 90276 219144 92224 219473
rect 92392 219144 94340 219473
rect 94508 219144 96364 219473
rect 96532 219144 98480 219473
rect 98648 219144 100504 219473
rect 100672 219144 102620 219473
rect 102788 219144 104644 219473
rect 104812 219144 106760 219473
rect 106928 219144 108784 219473
rect 108952 219144 110900 219473
rect 111068 219144 113016 219473
rect 113184 219144 115040 219473
rect 115208 219144 117156 219473
rect 117324 219144 119180 219473
rect 119348 219144 121296 219473
rect 121464 219144 123320 219473
rect 123488 219144 125436 219473
rect 125604 219144 127460 219473
rect 127628 219144 129576 219473
rect 129744 219144 131692 219473
rect 131860 219144 133716 219473
rect 133884 219144 135832 219473
rect 136000 219144 137856 219473
rect 138024 219144 139972 219473
rect 140140 219144 141996 219473
rect 142164 219144 144112 219473
rect 144280 219144 146136 219473
rect 146304 219144 148252 219473
rect 148420 219144 150368 219473
rect 150536 219144 152392 219473
rect 152560 219144 154508 219473
rect 154676 219144 156532 219473
rect 156700 219144 158648 219473
rect 158816 219144 160672 219473
rect 160840 219144 162788 219473
rect 162956 219144 164812 219473
rect 164980 219144 166928 219473
rect 167096 219144 169044 219473
rect 169212 219144 171068 219473
rect 171236 219144 173184 219473
rect 173352 219144 175208 219473
rect 175376 219144 177324 219473
rect 177492 219144 179348 219473
rect 179516 219144 181464 219473
rect 181632 219144 183488 219473
rect 183656 219144 185604 219473
rect 185772 219144 187720 219473
rect 187888 219144 189744 219473
rect 189912 219144 191860 219473
rect 192028 219144 193884 219473
rect 194052 219144 196000 219473
rect 196168 219144 198024 219473
rect 198192 219144 200140 219473
rect 200308 219144 202164 219473
rect 202332 219144 204280 219473
rect 204448 219144 206396 219473
rect 206564 219144 208420 219473
rect 208588 219144 210536 219473
rect 210704 219144 212560 219473
rect 212728 219144 214676 219473
rect 214844 219144 216700 219473
rect 216868 219144 218816 219473
rect 218984 219144 219478 219473
rect 6 856 219478 219144
rect 6 439 408 856
rect 576 439 1328 856
rect 1496 439 2340 856
rect 2508 439 3260 856
rect 3428 439 4272 856
rect 4440 439 5192 856
rect 5360 439 6204 856
rect 6372 439 7124 856
rect 7292 439 8136 856
rect 8304 439 9056 856
rect 9224 439 10068 856
rect 10236 439 10988 856
rect 11156 439 12000 856
rect 12168 439 12920 856
rect 13088 439 13932 856
rect 14100 439 14852 856
rect 15020 439 15864 856
rect 16032 439 16876 856
rect 17044 439 17796 856
rect 17964 439 18808 856
rect 18976 439 19728 856
rect 19896 439 20740 856
rect 20908 439 21660 856
rect 21828 439 22672 856
rect 22840 439 23592 856
rect 23760 439 24604 856
rect 24772 439 25524 856
rect 25692 439 26536 856
rect 26704 439 27456 856
rect 27624 439 28468 856
rect 28636 439 29388 856
rect 29556 439 30400 856
rect 30568 439 31412 856
rect 31580 439 32332 856
rect 32500 439 33344 856
rect 33512 439 34264 856
rect 34432 439 35276 856
rect 35444 439 36196 856
rect 36364 439 37208 856
rect 37376 439 38128 856
rect 38296 439 39140 856
rect 39308 439 40060 856
rect 40228 439 41072 856
rect 41240 439 41992 856
rect 42160 439 43004 856
rect 43172 439 43924 856
rect 44092 439 44936 856
rect 45104 439 45948 856
rect 46116 439 46868 856
rect 47036 439 47880 856
rect 48048 439 48800 856
rect 48968 439 49812 856
rect 49980 439 50732 856
rect 50900 439 51744 856
rect 51912 439 52664 856
rect 52832 439 53676 856
rect 53844 439 54596 856
rect 54764 439 55608 856
rect 55776 439 56528 856
rect 56696 439 57540 856
rect 57708 439 58460 856
rect 58628 439 59472 856
rect 59640 439 60484 856
rect 60652 439 61404 856
rect 61572 439 62416 856
rect 62584 439 63336 856
rect 63504 439 64348 856
rect 64516 439 65268 856
rect 65436 439 66280 856
rect 66448 439 67200 856
rect 67368 439 68212 856
rect 68380 439 69132 856
rect 69300 439 70144 856
rect 70312 439 71064 856
rect 71232 439 72076 856
rect 72244 439 72996 856
rect 73164 439 74008 856
rect 74176 439 75020 856
rect 75188 439 75940 856
rect 76108 439 76952 856
rect 77120 439 77872 856
rect 78040 439 78884 856
rect 79052 439 79804 856
rect 79972 439 80816 856
rect 80984 439 81736 856
rect 81904 439 82748 856
rect 82916 439 83668 856
rect 83836 439 84680 856
rect 84848 439 85600 856
rect 85768 439 86612 856
rect 86780 439 87532 856
rect 87700 439 88544 856
rect 88712 439 89556 856
rect 89724 439 90476 856
rect 90644 439 91488 856
rect 91656 439 92408 856
rect 92576 439 93420 856
rect 93588 439 94340 856
rect 94508 439 95352 856
rect 95520 439 96272 856
rect 96440 439 97284 856
rect 97452 439 98204 856
rect 98372 439 99216 856
rect 99384 439 100136 856
rect 100304 439 101148 856
rect 101316 439 102068 856
rect 102236 439 103080 856
rect 103248 439 104092 856
rect 104260 439 105012 856
rect 105180 439 106024 856
rect 106192 439 106944 856
rect 107112 439 107956 856
rect 108124 439 108876 856
rect 109044 439 109888 856
rect 110056 439 110808 856
rect 110976 439 111820 856
rect 111988 439 112740 856
rect 112908 439 113752 856
rect 113920 439 114672 856
rect 114840 439 115684 856
rect 115852 439 116604 856
rect 116772 439 117616 856
rect 117784 439 118628 856
rect 118796 439 119548 856
rect 119716 439 120560 856
rect 120728 439 121480 856
rect 121648 439 122492 856
rect 122660 439 123412 856
rect 123580 439 124424 856
rect 124592 439 125344 856
rect 125512 439 126356 856
rect 126524 439 127276 856
rect 127444 439 128288 856
rect 128456 439 129208 856
rect 129376 439 130220 856
rect 130388 439 131140 856
rect 131308 439 132152 856
rect 132320 439 133164 856
rect 133332 439 134084 856
rect 134252 439 135096 856
rect 135264 439 136016 856
rect 136184 439 137028 856
rect 137196 439 137948 856
rect 138116 439 138960 856
rect 139128 439 139880 856
rect 140048 439 140892 856
rect 141060 439 141812 856
rect 141980 439 142824 856
rect 142992 439 143744 856
rect 143912 439 144756 856
rect 144924 439 145676 856
rect 145844 439 146688 856
rect 146856 439 147700 856
rect 147868 439 148620 856
rect 148788 439 149632 856
rect 149800 439 150552 856
rect 150720 439 151564 856
rect 151732 439 152484 856
rect 152652 439 153496 856
rect 153664 439 154416 856
rect 154584 439 155428 856
rect 155596 439 156348 856
rect 156516 439 157360 856
rect 157528 439 158280 856
rect 158448 439 159292 856
rect 159460 439 160212 856
rect 160380 439 161224 856
rect 161392 439 162236 856
rect 162404 439 163156 856
rect 163324 439 164168 856
rect 164336 439 165088 856
rect 165256 439 166100 856
rect 166268 439 167020 856
rect 167188 439 168032 856
rect 168200 439 168952 856
rect 169120 439 169964 856
rect 170132 439 170884 856
rect 171052 439 171896 856
rect 172064 439 172816 856
rect 172984 439 173828 856
rect 173996 439 174748 856
rect 174916 439 175760 856
rect 175928 439 176772 856
rect 176940 439 177692 856
rect 177860 439 178704 856
rect 178872 439 179624 856
rect 179792 439 180636 856
rect 180804 439 181556 856
rect 181724 439 182568 856
rect 182736 439 183488 856
rect 183656 439 184500 856
rect 184668 439 185420 856
rect 185588 439 186432 856
rect 186600 439 187352 856
rect 187520 439 188364 856
rect 188532 439 189284 856
rect 189452 439 190296 856
rect 190464 439 191308 856
rect 191476 439 192228 856
rect 192396 439 193240 856
rect 193408 439 194160 856
rect 194328 439 195172 856
rect 195340 439 196092 856
rect 196260 439 197104 856
rect 197272 439 198024 856
rect 198192 439 199036 856
rect 199204 439 199956 856
rect 200124 439 200968 856
rect 201136 439 201888 856
rect 202056 439 202900 856
rect 203068 439 203820 856
rect 203988 439 204832 856
rect 205000 439 205844 856
rect 206012 439 206764 856
rect 206932 439 207776 856
rect 207944 439 208696 856
rect 208864 439 209708 856
rect 209876 439 210628 856
rect 210796 439 211640 856
rect 211808 439 212560 856
rect 212728 439 213572 856
rect 213740 439 214492 856
rect 214660 439 215504 856
rect 215672 439 216424 856
rect 216592 439 217436 856
rect 217604 439 218356 856
rect 218524 439 219368 856
<< metal3 >>
rect 219186 219376 219986 219496
rect 219186 218424 219986 218544
rect 219186 217336 219986 217456
rect 219186 216384 219986 216504
rect 219186 215296 219986 215416
rect 219186 214344 219986 214464
rect 219186 213392 219986 213512
rect 219186 212304 219986 212424
rect 219186 211352 219986 211472
rect 219186 210264 219986 210384
rect 219186 209312 219986 209432
rect 219186 208224 219986 208344
rect 219186 207272 219986 207392
rect 219186 206320 219986 206440
rect 219186 205232 219986 205352
rect 219186 204280 219986 204400
rect 219186 203192 219986 203312
rect 219186 202240 219986 202360
rect 219186 201152 219986 201272
rect 219186 200200 219986 200320
rect 219186 199248 219986 199368
rect 219186 198160 219986 198280
rect 219186 197208 219986 197328
rect 219186 196120 219986 196240
rect 219186 195168 219986 195288
rect 219186 194216 219986 194336
rect 219186 193128 219986 193248
rect 219186 192176 219986 192296
rect 219186 191088 219986 191208
rect 219186 190136 219986 190256
rect 219186 189048 219986 189168
rect 219186 188096 219986 188216
rect 219186 187144 219986 187264
rect 219186 186056 219986 186176
rect 219186 185104 219986 185224
rect 219186 184016 219986 184136
rect 219186 183064 219986 183184
rect 219186 181976 219986 182096
rect 219186 181024 219986 181144
rect 219186 180072 219986 180192
rect 219186 178984 219986 179104
rect 219186 178032 219986 178152
rect 219186 176944 219986 177064
rect 219186 175992 219986 176112
rect 219186 175040 219986 175160
rect 219186 173952 219986 174072
rect 219186 173000 219986 173120
rect 219186 171912 219986 172032
rect 219186 170960 219986 171080
rect 219186 169872 219986 169992
rect 219186 168920 219986 169040
rect 219186 167968 219986 168088
rect 219186 166880 219986 167000
rect 219186 165928 219986 166048
rect 219186 164840 219986 164960
rect 219186 163888 219986 164008
rect 219186 162800 219986 162920
rect 219186 161848 219986 161968
rect 219186 160896 219986 161016
rect 219186 159808 219986 159928
rect 219186 158856 219986 158976
rect 219186 157768 219986 157888
rect 219186 156816 219986 156936
rect 219186 155728 219986 155848
rect 219186 154776 219986 154896
rect 219186 153824 219986 153944
rect 219186 152736 219986 152856
rect 219186 151784 219986 151904
rect 219186 150696 219986 150816
rect 219186 149744 219986 149864
rect 219186 148792 219986 148912
rect 219186 147704 219986 147824
rect 219186 146752 219986 146872
rect 219186 145664 219986 145784
rect 219186 144712 219986 144832
rect 219186 143624 219986 143744
rect 219186 142672 219986 142792
rect 219186 141720 219986 141840
rect 219186 140632 219986 140752
rect 219186 139680 219986 139800
rect 219186 138592 219986 138712
rect 219186 137640 219986 137760
rect 219186 136552 219986 136672
rect 219186 135600 219986 135720
rect 219186 134648 219986 134768
rect 219186 133560 219986 133680
rect 219186 132608 219986 132728
rect 219186 131520 219986 131640
rect 219186 130568 219986 130688
rect 219186 129616 219986 129736
rect 219186 128528 219986 128648
rect 219186 127576 219986 127696
rect 219186 126488 219986 126608
rect 219186 125536 219986 125656
rect 219186 124448 219986 124568
rect 219186 123496 219986 123616
rect 219186 122544 219986 122664
rect 219186 121456 219986 121576
rect 219186 120504 219986 120624
rect 219186 119416 219986 119536
rect 219186 118464 219986 118584
rect 219186 117376 219986 117496
rect 219186 116424 219986 116544
rect 219186 115472 219986 115592
rect 219186 114384 219986 114504
rect 219186 113432 219986 113552
rect 219186 112344 219986 112464
rect 219186 111392 219986 111512
rect 219186 110440 219986 110560
rect 219186 109352 219986 109472
rect 219186 108400 219986 108520
rect 219186 107312 219986 107432
rect 219186 106360 219986 106480
rect 219186 105272 219986 105392
rect 219186 104320 219986 104440
rect 219186 103368 219986 103488
rect 219186 102280 219986 102400
rect 219186 101328 219986 101448
rect 219186 100240 219986 100360
rect 219186 99288 219986 99408
rect 219186 98200 219986 98320
rect 219186 97248 219986 97368
rect 219186 96296 219986 96416
rect 219186 95208 219986 95328
rect 219186 94256 219986 94376
rect 219186 93168 219986 93288
rect 219186 92216 219986 92336
rect 219186 91128 219986 91248
rect 219186 90176 219986 90296
rect 219186 89224 219986 89344
rect 219186 88136 219986 88256
rect 219186 87184 219986 87304
rect 219186 86096 219986 86216
rect 219186 85144 219986 85264
rect 219186 84192 219986 84312
rect 219186 83104 219986 83224
rect 219186 82152 219986 82272
rect 219186 81064 219986 81184
rect 219186 80112 219986 80232
rect 219186 79024 219986 79144
rect 219186 78072 219986 78192
rect 219186 77120 219986 77240
rect 219186 76032 219986 76152
rect 219186 75080 219986 75200
rect 219186 73992 219986 74112
rect 219186 73040 219986 73160
rect 219186 71952 219986 72072
rect 219186 71000 219986 71120
rect 219186 70048 219986 70168
rect 219186 68960 219986 69080
rect 219186 68008 219986 68128
rect 219186 66920 219986 67040
rect 219186 65968 219986 66088
rect 219186 65016 219986 65136
rect 219186 63928 219986 64048
rect 219186 62976 219986 63096
rect 219186 61888 219986 62008
rect 219186 60936 219986 61056
rect 219186 59848 219986 59968
rect 219186 58896 219986 59016
rect 219186 57944 219986 58064
rect 219186 56856 219986 56976
rect 219186 55904 219986 56024
rect 219186 54816 219986 54936
rect 219186 53864 219986 53984
rect 219186 52776 219986 52896
rect 219186 51824 219986 51944
rect 219186 50872 219986 50992
rect 219186 49784 219986 49904
rect 219186 48832 219986 48952
rect 219186 47744 219986 47864
rect 219186 46792 219986 46912
rect 219186 45704 219986 45824
rect 219186 44752 219986 44872
rect 219186 43800 219986 43920
rect 219186 42712 219986 42832
rect 219186 41760 219986 41880
rect 219186 40672 219986 40792
rect 219186 39720 219986 39840
rect 219186 38768 219986 38888
rect 219186 37680 219986 37800
rect 219186 36728 219986 36848
rect 219186 35640 219986 35760
rect 219186 34688 219986 34808
rect 219186 33600 219986 33720
rect 219186 32648 219986 32768
rect 219186 31696 219986 31816
rect 219186 30608 219986 30728
rect 219186 29656 219986 29776
rect 219186 28568 219986 28688
rect 219186 27616 219986 27736
rect 219186 26528 219986 26648
rect 219186 25576 219986 25696
rect 219186 24624 219986 24744
rect 219186 23536 219986 23656
rect 219186 22584 219986 22704
rect 219186 21496 219986 21616
rect 219186 20544 219986 20664
rect 219186 19592 219986 19712
rect 219186 18504 219986 18624
rect 219186 17552 219986 17672
rect 219186 16464 219986 16584
rect 219186 15512 219986 15632
rect 219186 14424 219986 14544
rect 219186 13472 219986 13592
rect 219186 12520 219986 12640
rect 219186 11432 219986 11552
rect 219186 10480 219986 10600
rect 219186 9392 219986 9512
rect 219186 8440 219986 8560
rect 219186 7352 219986 7472
rect 219186 6400 219986 6520
rect 219186 5448 219986 5568
rect 219186 4360 219986 4480
rect 219186 3408 219986 3528
rect 219186 2320 219986 2440
rect 219186 1368 219986 1488
rect 219186 416 219986 536
<< obsm3 >>
rect 1011 219296 219106 219469
rect 1011 218624 219186 219296
rect 1011 218344 219106 218624
rect 1011 217536 219186 218344
rect 1011 217256 219106 217536
rect 1011 216584 219186 217256
rect 1011 216304 219106 216584
rect 1011 215496 219186 216304
rect 1011 215216 219106 215496
rect 1011 214544 219186 215216
rect 1011 214264 219106 214544
rect 1011 213592 219186 214264
rect 1011 213312 219106 213592
rect 1011 212504 219186 213312
rect 1011 212224 219106 212504
rect 1011 211552 219186 212224
rect 1011 211272 219106 211552
rect 1011 210464 219186 211272
rect 1011 210184 219106 210464
rect 1011 209512 219186 210184
rect 1011 209232 219106 209512
rect 1011 208424 219186 209232
rect 1011 208144 219106 208424
rect 1011 207472 219186 208144
rect 1011 207192 219106 207472
rect 1011 206520 219186 207192
rect 1011 206240 219106 206520
rect 1011 205432 219186 206240
rect 1011 205152 219106 205432
rect 1011 204480 219186 205152
rect 1011 204200 219106 204480
rect 1011 203392 219186 204200
rect 1011 203112 219106 203392
rect 1011 202440 219186 203112
rect 1011 202160 219106 202440
rect 1011 201352 219186 202160
rect 1011 201072 219106 201352
rect 1011 200400 219186 201072
rect 1011 200120 219106 200400
rect 1011 199448 219186 200120
rect 1011 199168 219106 199448
rect 1011 198360 219186 199168
rect 1011 198080 219106 198360
rect 1011 197408 219186 198080
rect 1011 197128 219106 197408
rect 1011 196320 219186 197128
rect 1011 196040 219106 196320
rect 1011 195368 219186 196040
rect 1011 195088 219106 195368
rect 1011 194416 219186 195088
rect 1011 194136 219106 194416
rect 1011 193328 219186 194136
rect 1011 193048 219106 193328
rect 1011 192376 219186 193048
rect 1011 192096 219106 192376
rect 1011 191288 219186 192096
rect 1011 191008 219106 191288
rect 1011 190336 219186 191008
rect 1011 190056 219106 190336
rect 1011 189248 219186 190056
rect 1011 188968 219106 189248
rect 1011 188296 219186 188968
rect 1011 188016 219106 188296
rect 1011 187344 219186 188016
rect 1011 187064 219106 187344
rect 1011 186256 219186 187064
rect 1011 185976 219106 186256
rect 1011 185304 219186 185976
rect 1011 185024 219106 185304
rect 1011 184216 219186 185024
rect 1011 183936 219106 184216
rect 1011 183264 219186 183936
rect 1011 182984 219106 183264
rect 1011 182176 219186 182984
rect 1011 181896 219106 182176
rect 1011 181224 219186 181896
rect 1011 180944 219106 181224
rect 1011 180272 219186 180944
rect 1011 179992 219106 180272
rect 1011 179184 219186 179992
rect 1011 178904 219106 179184
rect 1011 178232 219186 178904
rect 1011 177952 219106 178232
rect 1011 177144 219186 177952
rect 1011 176864 219106 177144
rect 1011 176192 219186 176864
rect 1011 175912 219106 176192
rect 1011 175240 219186 175912
rect 1011 174960 219106 175240
rect 1011 174152 219186 174960
rect 1011 173872 219106 174152
rect 1011 173200 219186 173872
rect 1011 172920 219106 173200
rect 1011 172112 219186 172920
rect 1011 171832 219106 172112
rect 1011 171160 219186 171832
rect 1011 170880 219106 171160
rect 1011 170072 219186 170880
rect 1011 169792 219106 170072
rect 1011 169120 219186 169792
rect 1011 168840 219106 169120
rect 1011 168168 219186 168840
rect 1011 167888 219106 168168
rect 1011 167080 219186 167888
rect 1011 166800 219106 167080
rect 1011 166128 219186 166800
rect 1011 165848 219106 166128
rect 1011 165040 219186 165848
rect 1011 164760 219106 165040
rect 1011 164088 219186 164760
rect 1011 163808 219106 164088
rect 1011 163000 219186 163808
rect 1011 162720 219106 163000
rect 1011 162048 219186 162720
rect 1011 161768 219106 162048
rect 1011 161096 219186 161768
rect 1011 160816 219106 161096
rect 1011 160008 219186 160816
rect 1011 159728 219106 160008
rect 1011 159056 219186 159728
rect 1011 158776 219106 159056
rect 1011 157968 219186 158776
rect 1011 157688 219106 157968
rect 1011 157016 219186 157688
rect 1011 156736 219106 157016
rect 1011 155928 219186 156736
rect 1011 155648 219106 155928
rect 1011 154976 219186 155648
rect 1011 154696 219106 154976
rect 1011 154024 219186 154696
rect 1011 153744 219106 154024
rect 1011 152936 219186 153744
rect 1011 152656 219106 152936
rect 1011 151984 219186 152656
rect 1011 151704 219106 151984
rect 1011 150896 219186 151704
rect 1011 150616 219106 150896
rect 1011 149944 219186 150616
rect 1011 149664 219106 149944
rect 1011 148992 219186 149664
rect 1011 148712 219106 148992
rect 1011 147904 219186 148712
rect 1011 147624 219106 147904
rect 1011 146952 219186 147624
rect 1011 146672 219106 146952
rect 1011 145864 219186 146672
rect 1011 145584 219106 145864
rect 1011 144912 219186 145584
rect 1011 144632 219106 144912
rect 1011 143824 219186 144632
rect 1011 143544 219106 143824
rect 1011 142872 219186 143544
rect 1011 142592 219106 142872
rect 1011 141920 219186 142592
rect 1011 141640 219106 141920
rect 1011 140832 219186 141640
rect 1011 140552 219106 140832
rect 1011 139880 219186 140552
rect 1011 139600 219106 139880
rect 1011 138792 219186 139600
rect 1011 138512 219106 138792
rect 1011 137840 219186 138512
rect 1011 137560 219106 137840
rect 1011 136752 219186 137560
rect 1011 136472 219106 136752
rect 1011 135800 219186 136472
rect 1011 135520 219106 135800
rect 1011 134848 219186 135520
rect 1011 134568 219106 134848
rect 1011 133760 219186 134568
rect 1011 133480 219106 133760
rect 1011 132808 219186 133480
rect 1011 132528 219106 132808
rect 1011 131720 219186 132528
rect 1011 131440 219106 131720
rect 1011 130768 219186 131440
rect 1011 130488 219106 130768
rect 1011 129816 219186 130488
rect 1011 129536 219106 129816
rect 1011 128728 219186 129536
rect 1011 128448 219106 128728
rect 1011 127776 219186 128448
rect 1011 127496 219106 127776
rect 1011 126688 219186 127496
rect 1011 126408 219106 126688
rect 1011 125736 219186 126408
rect 1011 125456 219106 125736
rect 1011 124648 219186 125456
rect 1011 124368 219106 124648
rect 1011 123696 219186 124368
rect 1011 123416 219106 123696
rect 1011 122744 219186 123416
rect 1011 122464 219106 122744
rect 1011 121656 219186 122464
rect 1011 121376 219106 121656
rect 1011 120704 219186 121376
rect 1011 120424 219106 120704
rect 1011 119616 219186 120424
rect 1011 119336 219106 119616
rect 1011 118664 219186 119336
rect 1011 118384 219106 118664
rect 1011 117576 219186 118384
rect 1011 117296 219106 117576
rect 1011 116624 219186 117296
rect 1011 116344 219106 116624
rect 1011 115672 219186 116344
rect 1011 115392 219106 115672
rect 1011 114584 219186 115392
rect 1011 114304 219106 114584
rect 1011 113632 219186 114304
rect 1011 113352 219106 113632
rect 1011 112544 219186 113352
rect 1011 112264 219106 112544
rect 1011 111592 219186 112264
rect 1011 111312 219106 111592
rect 1011 110640 219186 111312
rect 1011 110360 219106 110640
rect 1011 109552 219186 110360
rect 1011 109272 219106 109552
rect 1011 108600 219186 109272
rect 1011 108320 219106 108600
rect 1011 107512 219186 108320
rect 1011 107232 219106 107512
rect 1011 106560 219186 107232
rect 1011 106280 219106 106560
rect 1011 105472 219186 106280
rect 1011 105192 219106 105472
rect 1011 104520 219186 105192
rect 1011 104240 219106 104520
rect 1011 103568 219186 104240
rect 1011 103288 219106 103568
rect 1011 102480 219186 103288
rect 1011 102200 219106 102480
rect 1011 101528 219186 102200
rect 1011 101248 219106 101528
rect 1011 100440 219186 101248
rect 1011 100160 219106 100440
rect 1011 99488 219186 100160
rect 1011 99208 219106 99488
rect 1011 98400 219186 99208
rect 1011 98120 219106 98400
rect 1011 97448 219186 98120
rect 1011 97168 219106 97448
rect 1011 96496 219186 97168
rect 1011 96216 219106 96496
rect 1011 95408 219186 96216
rect 1011 95128 219106 95408
rect 1011 94456 219186 95128
rect 1011 94176 219106 94456
rect 1011 93368 219186 94176
rect 1011 93088 219106 93368
rect 1011 92416 219186 93088
rect 1011 92136 219106 92416
rect 1011 91328 219186 92136
rect 1011 91048 219106 91328
rect 1011 90376 219186 91048
rect 1011 90096 219106 90376
rect 1011 89424 219186 90096
rect 1011 89144 219106 89424
rect 1011 88336 219186 89144
rect 1011 88056 219106 88336
rect 1011 87384 219186 88056
rect 1011 87104 219106 87384
rect 1011 86296 219186 87104
rect 1011 86016 219106 86296
rect 1011 85344 219186 86016
rect 1011 85064 219106 85344
rect 1011 84392 219186 85064
rect 1011 84112 219106 84392
rect 1011 83304 219186 84112
rect 1011 83024 219106 83304
rect 1011 82352 219186 83024
rect 1011 82072 219106 82352
rect 1011 81264 219186 82072
rect 1011 80984 219106 81264
rect 1011 80312 219186 80984
rect 1011 80032 219106 80312
rect 1011 79224 219186 80032
rect 1011 78944 219106 79224
rect 1011 78272 219186 78944
rect 1011 77992 219106 78272
rect 1011 77320 219186 77992
rect 1011 77040 219106 77320
rect 1011 76232 219186 77040
rect 1011 75952 219106 76232
rect 1011 75280 219186 75952
rect 1011 75000 219106 75280
rect 1011 74192 219186 75000
rect 1011 73912 219106 74192
rect 1011 73240 219186 73912
rect 1011 72960 219106 73240
rect 1011 72152 219186 72960
rect 1011 71872 219106 72152
rect 1011 71200 219186 71872
rect 1011 70920 219106 71200
rect 1011 70248 219186 70920
rect 1011 69968 219106 70248
rect 1011 69160 219186 69968
rect 1011 68880 219106 69160
rect 1011 68208 219186 68880
rect 1011 67928 219106 68208
rect 1011 67120 219186 67928
rect 1011 66840 219106 67120
rect 1011 66168 219186 66840
rect 1011 65888 219106 66168
rect 1011 65216 219186 65888
rect 1011 64936 219106 65216
rect 1011 64128 219186 64936
rect 1011 63848 219106 64128
rect 1011 63176 219186 63848
rect 1011 62896 219106 63176
rect 1011 62088 219186 62896
rect 1011 61808 219106 62088
rect 1011 61136 219186 61808
rect 1011 60856 219106 61136
rect 1011 60048 219186 60856
rect 1011 59768 219106 60048
rect 1011 59096 219186 59768
rect 1011 58816 219106 59096
rect 1011 58144 219186 58816
rect 1011 57864 219106 58144
rect 1011 57056 219186 57864
rect 1011 56776 219106 57056
rect 1011 56104 219186 56776
rect 1011 55824 219106 56104
rect 1011 55016 219186 55824
rect 1011 54736 219106 55016
rect 1011 54064 219186 54736
rect 1011 53784 219106 54064
rect 1011 52976 219186 53784
rect 1011 52696 219106 52976
rect 1011 52024 219186 52696
rect 1011 51744 219106 52024
rect 1011 51072 219186 51744
rect 1011 50792 219106 51072
rect 1011 49984 219186 50792
rect 1011 49704 219106 49984
rect 1011 49032 219186 49704
rect 1011 48752 219106 49032
rect 1011 47944 219186 48752
rect 1011 47664 219106 47944
rect 1011 46992 219186 47664
rect 1011 46712 219106 46992
rect 1011 45904 219186 46712
rect 1011 45624 219106 45904
rect 1011 44952 219186 45624
rect 1011 44672 219106 44952
rect 1011 44000 219186 44672
rect 1011 43720 219106 44000
rect 1011 42912 219186 43720
rect 1011 42632 219106 42912
rect 1011 41960 219186 42632
rect 1011 41680 219106 41960
rect 1011 40872 219186 41680
rect 1011 40592 219106 40872
rect 1011 39920 219186 40592
rect 1011 39640 219106 39920
rect 1011 38968 219186 39640
rect 1011 38688 219106 38968
rect 1011 37880 219186 38688
rect 1011 37600 219106 37880
rect 1011 36928 219186 37600
rect 1011 36648 219106 36928
rect 1011 35840 219186 36648
rect 1011 35560 219106 35840
rect 1011 34888 219186 35560
rect 1011 34608 219106 34888
rect 1011 33800 219186 34608
rect 1011 33520 219106 33800
rect 1011 32848 219186 33520
rect 1011 32568 219106 32848
rect 1011 31896 219186 32568
rect 1011 31616 219106 31896
rect 1011 30808 219186 31616
rect 1011 30528 219106 30808
rect 1011 29856 219186 30528
rect 1011 29576 219106 29856
rect 1011 28768 219186 29576
rect 1011 28488 219106 28768
rect 1011 27816 219186 28488
rect 1011 27536 219106 27816
rect 1011 26728 219186 27536
rect 1011 26448 219106 26728
rect 1011 25776 219186 26448
rect 1011 25496 219106 25776
rect 1011 24824 219186 25496
rect 1011 24544 219106 24824
rect 1011 23736 219186 24544
rect 1011 23456 219106 23736
rect 1011 22784 219186 23456
rect 1011 22504 219106 22784
rect 1011 21696 219186 22504
rect 1011 21416 219106 21696
rect 1011 20744 219186 21416
rect 1011 20464 219106 20744
rect 1011 19792 219186 20464
rect 1011 19512 219106 19792
rect 1011 18704 219186 19512
rect 1011 18424 219106 18704
rect 1011 17752 219186 18424
rect 1011 17472 219106 17752
rect 1011 16664 219186 17472
rect 1011 16384 219106 16664
rect 1011 15712 219186 16384
rect 1011 15432 219106 15712
rect 1011 14624 219186 15432
rect 1011 14344 219106 14624
rect 1011 13672 219186 14344
rect 1011 13392 219106 13672
rect 1011 12720 219186 13392
rect 1011 12440 219106 12720
rect 1011 11632 219186 12440
rect 1011 11352 219106 11632
rect 1011 10680 219186 11352
rect 1011 10400 219106 10680
rect 1011 9592 219186 10400
rect 1011 9312 219106 9592
rect 1011 8640 219186 9312
rect 1011 8360 219106 8640
rect 1011 7552 219186 8360
rect 1011 7272 219106 7552
rect 1011 6600 219186 7272
rect 1011 6320 219106 6600
rect 1011 5648 219186 6320
rect 1011 5368 219106 5648
rect 1011 4560 219186 5368
rect 1011 4280 219106 4560
rect 1011 3608 219186 4280
rect 1011 3328 219106 3608
rect 1011 2520 219186 3328
rect 1011 2240 219106 2520
rect 1011 1568 219186 2240
rect 1011 1288 219106 1568
rect 1011 616 219186 1288
rect 1011 443 219106 616
<< metal4 >>
rect 4194 2128 4514 217648
rect 19554 2128 19874 217648
<< obsm4 >>
rect 5013 2128 19474 217648
rect 19954 2128 217783 217648
<< labels >>
rlabel metal3 s 219186 13472 219986 13592 6 cpu_addr_e[0]
port 1 nsew default output
rlabel metal3 s 219186 23536 219986 23656 6 cpu_addr_e[10]
port 2 nsew default output
rlabel metal3 s 219186 24624 219986 24744 6 cpu_addr_e[11]
port 3 nsew default output
rlabel metal3 s 219186 25576 219986 25696 6 cpu_addr_e[12]
port 4 nsew default output
rlabel metal3 s 219186 26528 219986 26648 6 cpu_addr_e[13]
port 5 nsew default output
rlabel metal3 s 219186 27616 219986 27736 6 cpu_addr_e[14]
port 6 nsew default output
rlabel metal3 s 219186 28568 219986 28688 6 cpu_addr_e[15]
port 7 nsew default output
rlabel metal3 s 219186 14424 219986 14544 6 cpu_addr_e[1]
port 8 nsew default output
rlabel metal3 s 219186 15512 219986 15632 6 cpu_addr_e[2]
port 9 nsew default output
rlabel metal3 s 219186 16464 219986 16584 6 cpu_addr_e[3]
port 10 nsew default output
rlabel metal3 s 219186 17552 219986 17672 6 cpu_addr_e[4]
port 11 nsew default output
rlabel metal3 s 219186 18504 219986 18624 6 cpu_addr_e[5]
port 12 nsew default output
rlabel metal3 s 219186 19592 219986 19712 6 cpu_addr_e[6]
port 13 nsew default output
rlabel metal3 s 219186 20544 219986 20664 6 cpu_addr_e[7]
port 14 nsew default output
rlabel metal3 s 219186 21496 219986 21616 6 cpu_addr_e[8]
port 15 nsew default output
rlabel metal3 s 219186 22584 219986 22704 6 cpu_addr_e[9]
port 16 nsew default output
rlabel metal2 s 21716 219200 21772 220000 6 cpu_addr_n[0]
port 17 nsew default output
rlabel metal2 s 42508 219200 42564 220000 6 cpu_addr_n[10]
port 18 nsew default output
rlabel metal2 s 44532 219200 44588 220000 6 cpu_addr_n[11]
port 19 nsew default output
rlabel metal2 s 46648 219200 46704 220000 6 cpu_addr_n[12]
port 20 nsew default output
rlabel metal2 s 48672 219200 48728 220000 6 cpu_addr_n[13]
port 21 nsew default output
rlabel metal2 s 50788 219200 50844 220000 6 cpu_addr_n[14]
port 22 nsew default output
rlabel metal2 s 52812 219200 52868 220000 6 cpu_addr_n[15]
port 23 nsew default output
rlabel metal2 s 23832 219200 23888 220000 6 cpu_addr_n[1]
port 24 nsew default output
rlabel metal2 s 25856 219200 25912 220000 6 cpu_addr_n[2]
port 25 nsew default output
rlabel metal2 s 27972 219200 28028 220000 6 cpu_addr_n[3]
port 26 nsew default output
rlabel metal2 s 29996 219200 30052 220000 6 cpu_addr_n[4]
port 27 nsew default output
rlabel metal2 s 32112 219200 32168 220000 6 cpu_addr_n[5]
port 28 nsew default output
rlabel metal2 s 34136 219200 34192 220000 6 cpu_addr_n[6]
port 29 nsew default output
rlabel metal2 s 36252 219200 36308 220000 6 cpu_addr_n[7]
port 30 nsew default output
rlabel metal2 s 38368 219200 38424 220000 6 cpu_addr_n[8]
port 31 nsew default output
rlabel metal2 s 40392 219200 40448 220000 6 cpu_addr_n[9]
port 32 nsew default output
rlabel metal3 s 219186 45704 219986 45824 6 cpu_dtr_e0[0]
port 33 nsew default input
rlabel metal3 s 219186 55904 219986 56024 6 cpu_dtr_e0[10]
port 34 nsew default input
rlabel metal3 s 219186 56856 219986 56976 6 cpu_dtr_e0[11]
port 35 nsew default input
rlabel metal3 s 219186 57944 219986 58064 6 cpu_dtr_e0[12]
port 36 nsew default input
rlabel metal3 s 219186 58896 219986 59016 6 cpu_dtr_e0[13]
port 37 nsew default input
rlabel metal3 s 219186 59848 219986 59968 6 cpu_dtr_e0[14]
port 38 nsew default input
rlabel metal3 s 219186 60936 219986 61056 6 cpu_dtr_e0[15]
port 39 nsew default input
rlabel metal3 s 219186 61888 219986 62008 6 cpu_dtr_e0[16]
port 40 nsew default input
rlabel metal3 s 219186 62976 219986 63096 6 cpu_dtr_e0[17]
port 41 nsew default input
rlabel metal3 s 219186 63928 219986 64048 6 cpu_dtr_e0[18]
port 42 nsew default input
rlabel metal3 s 219186 65016 219986 65136 6 cpu_dtr_e0[19]
port 43 nsew default input
rlabel metal3 s 219186 46792 219986 46912 6 cpu_dtr_e0[1]
port 44 nsew default input
rlabel metal3 s 219186 65968 219986 66088 6 cpu_dtr_e0[20]
port 45 nsew default input
rlabel metal3 s 219186 66920 219986 67040 6 cpu_dtr_e0[21]
port 46 nsew default input
rlabel metal3 s 219186 68008 219986 68128 6 cpu_dtr_e0[22]
port 47 nsew default input
rlabel metal3 s 219186 68960 219986 69080 6 cpu_dtr_e0[23]
port 48 nsew default input
rlabel metal3 s 219186 70048 219986 70168 6 cpu_dtr_e0[24]
port 49 nsew default input
rlabel metal3 s 219186 71000 219986 71120 6 cpu_dtr_e0[25]
port 50 nsew default input
rlabel metal3 s 219186 71952 219986 72072 6 cpu_dtr_e0[26]
port 51 nsew default input
rlabel metal3 s 219186 73040 219986 73160 6 cpu_dtr_e0[27]
port 52 nsew default input
rlabel metal3 s 219186 73992 219986 74112 6 cpu_dtr_e0[28]
port 53 nsew default input
rlabel metal3 s 219186 75080 219986 75200 6 cpu_dtr_e0[29]
port 54 nsew default input
rlabel metal3 s 219186 47744 219986 47864 6 cpu_dtr_e0[2]
port 55 nsew default input
rlabel metal3 s 219186 76032 219986 76152 6 cpu_dtr_e0[30]
port 56 nsew default input
rlabel metal3 s 219186 77120 219986 77240 6 cpu_dtr_e0[31]
port 57 nsew default input
rlabel metal3 s 219186 48832 219986 48952 6 cpu_dtr_e0[3]
port 58 nsew default input
rlabel metal3 s 219186 49784 219986 49904 6 cpu_dtr_e0[4]
port 59 nsew default input
rlabel metal3 s 219186 50872 219986 50992 6 cpu_dtr_e0[5]
port 60 nsew default input
rlabel metal3 s 219186 51824 219986 51944 6 cpu_dtr_e0[6]
port 61 nsew default input
rlabel metal3 s 219186 52776 219986 52896 6 cpu_dtr_e0[7]
port 62 nsew default input
rlabel metal3 s 219186 53864 219986 53984 6 cpu_dtr_e0[8]
port 63 nsew default input
rlabel metal3 s 219186 54816 219986 54936 6 cpu_dtr_e0[9]
port 64 nsew default input
rlabel metal3 s 219186 78072 219986 78192 6 cpu_dtr_e1[0]
port 65 nsew default input
rlabel metal3 s 219186 88136 219986 88256 6 cpu_dtr_e1[10]
port 66 nsew default input
rlabel metal3 s 219186 89224 219986 89344 6 cpu_dtr_e1[11]
port 67 nsew default input
rlabel metal3 s 219186 90176 219986 90296 6 cpu_dtr_e1[12]
port 68 nsew default input
rlabel metal3 s 219186 91128 219986 91248 6 cpu_dtr_e1[13]
port 69 nsew default input
rlabel metal3 s 219186 92216 219986 92336 6 cpu_dtr_e1[14]
port 70 nsew default input
rlabel metal3 s 219186 93168 219986 93288 6 cpu_dtr_e1[15]
port 71 nsew default input
rlabel metal3 s 219186 94256 219986 94376 6 cpu_dtr_e1[16]
port 72 nsew default input
rlabel metal3 s 219186 95208 219986 95328 6 cpu_dtr_e1[17]
port 73 nsew default input
rlabel metal3 s 219186 96296 219986 96416 6 cpu_dtr_e1[18]
port 74 nsew default input
rlabel metal3 s 219186 97248 219986 97368 6 cpu_dtr_e1[19]
port 75 nsew default input
rlabel metal3 s 219186 79024 219986 79144 6 cpu_dtr_e1[1]
port 76 nsew default input
rlabel metal3 s 219186 98200 219986 98320 6 cpu_dtr_e1[20]
port 77 nsew default input
rlabel metal3 s 219186 99288 219986 99408 6 cpu_dtr_e1[21]
port 78 nsew default input
rlabel metal3 s 219186 100240 219986 100360 6 cpu_dtr_e1[22]
port 79 nsew default input
rlabel metal3 s 219186 101328 219986 101448 6 cpu_dtr_e1[23]
port 80 nsew default input
rlabel metal3 s 219186 102280 219986 102400 6 cpu_dtr_e1[24]
port 81 nsew default input
rlabel metal3 s 219186 103368 219986 103488 6 cpu_dtr_e1[25]
port 82 nsew default input
rlabel metal3 s 219186 104320 219986 104440 6 cpu_dtr_e1[26]
port 83 nsew default input
rlabel metal3 s 219186 105272 219986 105392 6 cpu_dtr_e1[27]
port 84 nsew default input
rlabel metal3 s 219186 106360 219986 106480 6 cpu_dtr_e1[28]
port 85 nsew default input
rlabel metal3 s 219186 107312 219986 107432 6 cpu_dtr_e1[29]
port 86 nsew default input
rlabel metal3 s 219186 80112 219986 80232 6 cpu_dtr_e1[2]
port 87 nsew default input
rlabel metal3 s 219186 108400 219986 108520 6 cpu_dtr_e1[30]
port 88 nsew default input
rlabel metal3 s 219186 109352 219986 109472 6 cpu_dtr_e1[31]
port 89 nsew default input
rlabel metal3 s 219186 81064 219986 81184 6 cpu_dtr_e1[3]
port 90 nsew default input
rlabel metal3 s 219186 82152 219986 82272 6 cpu_dtr_e1[4]
port 91 nsew default input
rlabel metal3 s 219186 83104 219986 83224 6 cpu_dtr_e1[5]
port 92 nsew default input
rlabel metal3 s 219186 84192 219986 84312 6 cpu_dtr_e1[6]
port 93 nsew default input
rlabel metal3 s 219186 85144 219986 85264 6 cpu_dtr_e1[7]
port 94 nsew default input
rlabel metal3 s 219186 86096 219986 86216 6 cpu_dtr_e1[8]
port 95 nsew default input
rlabel metal3 s 219186 87184 219986 87304 6 cpu_dtr_e1[9]
port 96 nsew default input
rlabel metal2 s 88140 219200 88196 220000 6 cpu_dtr_n0[0]
port 97 nsew default input
rlabel metal2 s 108840 219200 108896 220000 6 cpu_dtr_n0[10]
port 98 nsew default input
rlabel metal2 s 110956 219200 111012 220000 6 cpu_dtr_n0[11]
port 99 nsew default input
rlabel metal2 s 113072 219200 113128 220000 6 cpu_dtr_n0[12]
port 100 nsew default input
rlabel metal2 s 115096 219200 115152 220000 6 cpu_dtr_n0[13]
port 101 nsew default input
rlabel metal2 s 117212 219200 117268 220000 6 cpu_dtr_n0[14]
port 102 nsew default input
rlabel metal2 s 119236 219200 119292 220000 6 cpu_dtr_n0[15]
port 103 nsew default input
rlabel metal2 s 121352 219200 121408 220000 6 cpu_dtr_n0[16]
port 104 nsew default input
rlabel metal2 s 123376 219200 123432 220000 6 cpu_dtr_n0[17]
port 105 nsew default input
rlabel metal2 s 125492 219200 125548 220000 6 cpu_dtr_n0[18]
port 106 nsew default input
rlabel metal2 s 127516 219200 127572 220000 6 cpu_dtr_n0[19]
port 107 nsew default input
rlabel metal2 s 90164 219200 90220 220000 6 cpu_dtr_n0[1]
port 108 nsew default input
rlabel metal2 s 129632 219200 129688 220000 6 cpu_dtr_n0[20]
port 109 nsew default input
rlabel metal2 s 131748 219200 131804 220000 6 cpu_dtr_n0[21]
port 110 nsew default input
rlabel metal2 s 133772 219200 133828 220000 6 cpu_dtr_n0[22]
port 111 nsew default input
rlabel metal2 s 135888 219200 135944 220000 6 cpu_dtr_n0[23]
port 112 nsew default input
rlabel metal2 s 137912 219200 137968 220000 6 cpu_dtr_n0[24]
port 113 nsew default input
rlabel metal2 s 140028 219200 140084 220000 6 cpu_dtr_n0[25]
port 114 nsew default input
rlabel metal2 s 142052 219200 142108 220000 6 cpu_dtr_n0[26]
port 115 nsew default input
rlabel metal2 s 144168 219200 144224 220000 6 cpu_dtr_n0[27]
port 116 nsew default input
rlabel metal2 s 146192 219200 146248 220000 6 cpu_dtr_n0[28]
port 117 nsew default input
rlabel metal2 s 148308 219200 148364 220000 6 cpu_dtr_n0[29]
port 118 nsew default input
rlabel metal2 s 92280 219200 92336 220000 6 cpu_dtr_n0[2]
port 119 nsew default input
rlabel metal2 s 150424 219200 150480 220000 6 cpu_dtr_n0[30]
port 120 nsew default input
rlabel metal2 s 152448 219200 152504 220000 6 cpu_dtr_n0[31]
port 121 nsew default input
rlabel metal2 s 94396 219200 94452 220000 6 cpu_dtr_n0[3]
port 122 nsew default input
rlabel metal2 s 96420 219200 96476 220000 6 cpu_dtr_n0[4]
port 123 nsew default input
rlabel metal2 s 98536 219200 98592 220000 6 cpu_dtr_n0[5]
port 124 nsew default input
rlabel metal2 s 100560 219200 100616 220000 6 cpu_dtr_n0[6]
port 125 nsew default input
rlabel metal2 s 102676 219200 102732 220000 6 cpu_dtr_n0[7]
port 126 nsew default input
rlabel metal2 s 104700 219200 104756 220000 6 cpu_dtr_n0[8]
port 127 nsew default input
rlabel metal2 s 106816 219200 106872 220000 6 cpu_dtr_n0[9]
port 128 nsew default input
rlabel metal2 s 154564 219200 154620 220000 6 cpu_dtr_n1[0]
port 129 nsew default input
rlabel metal2 s 175264 219200 175320 220000 6 cpu_dtr_n1[10]
port 130 nsew default input
rlabel metal2 s 177380 219200 177436 220000 6 cpu_dtr_n1[11]
port 131 nsew default input
rlabel metal2 s 179404 219200 179460 220000 6 cpu_dtr_n1[12]
port 132 nsew default input
rlabel metal2 s 181520 219200 181576 220000 6 cpu_dtr_n1[13]
port 133 nsew default input
rlabel metal2 s 183544 219200 183600 220000 6 cpu_dtr_n1[14]
port 134 nsew default input
rlabel metal2 s 185660 219200 185716 220000 6 cpu_dtr_n1[15]
port 135 nsew default input
rlabel metal2 s 187776 219200 187832 220000 6 cpu_dtr_n1[16]
port 136 nsew default input
rlabel metal2 s 189800 219200 189856 220000 6 cpu_dtr_n1[17]
port 137 nsew default input
rlabel metal2 s 191916 219200 191972 220000 6 cpu_dtr_n1[18]
port 138 nsew default input
rlabel metal2 s 193940 219200 193996 220000 6 cpu_dtr_n1[19]
port 139 nsew default input
rlabel metal2 s 156588 219200 156644 220000 6 cpu_dtr_n1[1]
port 140 nsew default input
rlabel metal2 s 196056 219200 196112 220000 6 cpu_dtr_n1[20]
port 141 nsew default input
rlabel metal2 s 198080 219200 198136 220000 6 cpu_dtr_n1[21]
port 142 nsew default input
rlabel metal2 s 200196 219200 200252 220000 6 cpu_dtr_n1[22]
port 143 nsew default input
rlabel metal2 s 202220 219200 202276 220000 6 cpu_dtr_n1[23]
port 144 nsew default input
rlabel metal2 s 204336 219200 204392 220000 6 cpu_dtr_n1[24]
port 145 nsew default input
rlabel metal2 s 206452 219200 206508 220000 6 cpu_dtr_n1[25]
port 146 nsew default input
rlabel metal2 s 208476 219200 208532 220000 6 cpu_dtr_n1[26]
port 147 nsew default input
rlabel metal2 s 210592 219200 210648 220000 6 cpu_dtr_n1[27]
port 148 nsew default input
rlabel metal2 s 212616 219200 212672 220000 6 cpu_dtr_n1[28]
port 149 nsew default input
rlabel metal2 s 214732 219200 214788 220000 6 cpu_dtr_n1[29]
port 150 nsew default input
rlabel metal2 s 158704 219200 158760 220000 6 cpu_dtr_n1[2]
port 151 nsew default input
rlabel metal2 s 216756 219200 216812 220000 6 cpu_dtr_n1[30]
port 152 nsew default input
rlabel metal2 s 218872 219200 218928 220000 6 cpu_dtr_n1[31]
port 153 nsew default input
rlabel metal2 s 160728 219200 160784 220000 6 cpu_dtr_n1[3]
port 154 nsew default input
rlabel metal2 s 162844 219200 162900 220000 6 cpu_dtr_n1[4]
port 155 nsew default input
rlabel metal2 s 164868 219200 164924 220000 6 cpu_dtr_n1[5]
port 156 nsew default input
rlabel metal2 s 166984 219200 167040 220000 6 cpu_dtr_n1[6]
port 157 nsew default input
rlabel metal2 s 169100 219200 169156 220000 6 cpu_dtr_n1[7]
port 158 nsew default input
rlabel metal2 s 171124 219200 171180 220000 6 cpu_dtr_n1[8]
port 159 nsew default input
rlabel metal2 s 173240 219200 173296 220000 6 cpu_dtr_n1[9]
port 160 nsew default input
rlabel metal3 s 219186 29656 219986 29776 6 cpu_dtw_e[0]
port 161 nsew default output
rlabel metal3 s 219186 39720 219986 39840 6 cpu_dtw_e[10]
port 162 nsew default output
rlabel metal3 s 219186 40672 219986 40792 6 cpu_dtw_e[11]
port 163 nsew default output
rlabel metal3 s 219186 41760 219986 41880 6 cpu_dtw_e[12]
port 164 nsew default output
rlabel metal3 s 219186 42712 219986 42832 6 cpu_dtw_e[13]
port 165 nsew default output
rlabel metal3 s 219186 43800 219986 43920 6 cpu_dtw_e[14]
port 166 nsew default output
rlabel metal3 s 219186 44752 219986 44872 6 cpu_dtw_e[15]
port 167 nsew default output
rlabel metal3 s 219186 30608 219986 30728 6 cpu_dtw_e[1]
port 168 nsew default output
rlabel metal3 s 219186 31696 219986 31816 6 cpu_dtw_e[2]
port 169 nsew default output
rlabel metal3 s 219186 32648 219986 32768 6 cpu_dtw_e[3]
port 170 nsew default output
rlabel metal3 s 219186 33600 219986 33720 6 cpu_dtw_e[4]
port 171 nsew default output
rlabel metal3 s 219186 34688 219986 34808 6 cpu_dtw_e[5]
port 172 nsew default output
rlabel metal3 s 219186 35640 219986 35760 6 cpu_dtw_e[6]
port 173 nsew default output
rlabel metal3 s 219186 36728 219986 36848 6 cpu_dtw_e[7]
port 174 nsew default output
rlabel metal3 s 219186 37680 219986 37800 6 cpu_dtw_e[8]
port 175 nsew default output
rlabel metal3 s 219186 38768 219986 38888 6 cpu_dtw_e[9]
port 176 nsew default output
rlabel metal2 s 54928 219200 54984 220000 6 cpu_dtw_n[0]
port 177 nsew default output
rlabel metal2 s 75720 219200 75776 220000 6 cpu_dtw_n[10]
port 178 nsew default output
rlabel metal2 s 77744 219200 77800 220000 6 cpu_dtw_n[11]
port 179 nsew default output
rlabel metal2 s 79860 219200 79916 220000 6 cpu_dtw_n[12]
port 180 nsew default output
rlabel metal2 s 81884 219200 81940 220000 6 cpu_dtw_n[13]
port 181 nsew default output
rlabel metal2 s 84000 219200 84056 220000 6 cpu_dtw_n[14]
port 182 nsew default output
rlabel metal2 s 86024 219200 86080 220000 6 cpu_dtw_n[15]
port 183 nsew default output
rlabel metal2 s 57044 219200 57100 220000 6 cpu_dtw_n[1]
port 184 nsew default output
rlabel metal2 s 59068 219200 59124 220000 6 cpu_dtw_n[2]
port 185 nsew default output
rlabel metal2 s 61184 219200 61240 220000 6 cpu_dtw_n[3]
port 186 nsew default output
rlabel metal2 s 63208 219200 63264 220000 6 cpu_dtw_n[4]
port 187 nsew default output
rlabel metal2 s 65324 219200 65380 220000 6 cpu_dtw_n[5]
port 188 nsew default output
rlabel metal2 s 67348 219200 67404 220000 6 cpu_dtw_n[6]
port 189 nsew default output
rlabel metal2 s 69464 219200 69520 220000 6 cpu_dtw_n[7]
port 190 nsew default output
rlabel metal2 s 71488 219200 71544 220000 6 cpu_dtw_n[8]
port 191 nsew default output
rlabel metal2 s 73604 219200 73660 220000 6 cpu_dtw_n[9]
port 192 nsew default output
rlabel metal3 s 219186 3408 219986 3528 6 cpu_mask_e[0]
port 193 nsew default output
rlabel metal3 s 219186 4360 219986 4480 6 cpu_mask_e[1]
port 194 nsew default output
rlabel metal3 s 219186 5448 219986 5568 6 cpu_mask_e[2]
port 195 nsew default output
rlabel metal3 s 219186 6400 219986 6520 6 cpu_mask_e[3]
port 196 nsew default output
rlabel metal3 s 219186 7352 219986 7472 6 cpu_mask_e[4]
port 197 nsew default output
rlabel metal3 s 219186 8440 219986 8560 6 cpu_mask_e[5]
port 198 nsew default output
rlabel metal3 s 219186 9392 219986 9512 6 cpu_mask_e[6]
port 199 nsew default output
rlabel metal3 s 219186 10480 219986 10600 6 cpu_mask_e[7]
port 200 nsew default output
rlabel metal2 s 1016 219200 1072 220000 6 cpu_mask_n[0]
port 201 nsew default output
rlabel metal2 s 3040 219200 3096 220000 6 cpu_mask_n[1]
port 202 nsew default output
rlabel metal2 s 5156 219200 5212 220000 6 cpu_mask_n[2]
port 203 nsew default output
rlabel metal2 s 7180 219200 7236 220000 6 cpu_mask_n[3]
port 204 nsew default output
rlabel metal2 s 9296 219200 9352 220000 6 cpu_mask_n[4]
port 205 nsew default output
rlabel metal2 s 11320 219200 11376 220000 6 cpu_mask_n[5]
port 206 nsew default output
rlabel metal2 s 13436 219200 13492 220000 6 cpu_mask_n[6]
port 207 nsew default output
rlabel metal2 s 15460 219200 15516 220000 6 cpu_mask_n[7]
port 208 nsew default output
rlabel metal3 s 219186 11432 219986 11552 6 cpu_wen_e[0]
port 209 nsew default output
rlabel metal3 s 219186 12520 219986 12640 6 cpu_wen_e[1]
port 210 nsew default output
rlabel metal2 s 17576 219200 17632 220000 6 cpu_wen_n[0]
port 211 nsew default output
rlabel metal2 s 19692 219200 19748 220000 6 cpu_wen_n[1]
port 212 nsew default output
rlabel metal2 s 109944 0 110000 800 6 io_in[0]
port 213 nsew default input
rlabel metal2 s 139016 0 139072 800 6 io_in[10]
port 214 nsew default input
rlabel metal2 s 141868 0 141924 800 6 io_in[11]
port 215 nsew default input
rlabel metal2 s 144812 0 144868 800 6 io_in[12]
port 216 nsew default input
rlabel metal2 s 147756 0 147812 800 6 io_in[13]
port 217 nsew default input
rlabel metal2 s 150608 0 150664 800 6 io_in[14]
port 218 nsew default input
rlabel metal2 s 153552 0 153608 800 6 io_in[15]
port 219 nsew default input
rlabel metal2 s 156404 0 156460 800 6 io_in[16]
port 220 nsew default input
rlabel metal2 s 159348 0 159404 800 6 io_in[17]
port 221 nsew default input
rlabel metal2 s 162292 0 162348 800 6 io_in[18]
port 222 nsew default input
rlabel metal2 s 165144 0 165200 800 6 io_in[19]
port 223 nsew default input
rlabel metal2 s 112796 0 112852 800 6 io_in[1]
port 224 nsew default input
rlabel metal2 s 168088 0 168144 800 6 io_in[20]
port 225 nsew default input
rlabel metal2 s 170940 0 170996 800 6 io_in[21]
port 226 nsew default input
rlabel metal2 s 173884 0 173940 800 6 io_in[22]
port 227 nsew default input
rlabel metal2 s 176828 0 176884 800 6 io_in[23]
port 228 nsew default input
rlabel metal2 s 179680 0 179736 800 6 io_in[24]
port 229 nsew default input
rlabel metal2 s 182624 0 182680 800 6 io_in[25]
port 230 nsew default input
rlabel metal2 s 185476 0 185532 800 6 io_in[26]
port 231 nsew default input
rlabel metal2 s 188420 0 188476 800 6 io_in[27]
port 232 nsew default input
rlabel metal2 s 191364 0 191420 800 6 io_in[28]
port 233 nsew default input
rlabel metal2 s 194216 0 194272 800 6 io_in[29]
port 234 nsew default input
rlabel metal2 s 115740 0 115796 800 6 io_in[2]
port 235 nsew default input
rlabel metal2 s 197160 0 197216 800 6 io_in[30]
port 236 nsew default input
rlabel metal2 s 200012 0 200068 800 6 io_in[31]
port 237 nsew default input
rlabel metal2 s 202956 0 203012 800 6 io_in[32]
port 238 nsew default input
rlabel metal2 s 205900 0 205956 800 6 io_in[33]
port 239 nsew default input
rlabel metal2 s 208752 0 208808 800 6 io_in[34]
port 240 nsew default input
rlabel metal2 s 211696 0 211752 800 6 io_in[35]
port 241 nsew default input
rlabel metal2 s 214548 0 214604 800 6 io_in[36]
port 242 nsew default input
rlabel metal2 s 217492 0 217548 800 6 io_in[37]
port 243 nsew default input
rlabel metal2 s 118684 0 118740 800 6 io_in[3]
port 244 nsew default input
rlabel metal2 s 121536 0 121592 800 6 io_in[4]
port 245 nsew default input
rlabel metal2 s 124480 0 124536 800 6 io_in[5]
port 246 nsew default input
rlabel metal2 s 127332 0 127388 800 6 io_in[6]
port 247 nsew default input
rlabel metal2 s 130276 0 130332 800 6 io_in[7]
port 248 nsew default input
rlabel metal2 s 133220 0 133276 800 6 io_in[8]
port 249 nsew default input
rlabel metal2 s 136072 0 136128 800 6 io_in[9]
port 250 nsew default input
rlabel metal2 s 110864 0 110920 800 6 io_oeb[0]
port 251 nsew default output
rlabel metal2 s 139936 0 139992 800 6 io_oeb[10]
port 252 nsew default output
rlabel metal2 s 142880 0 142936 800 6 io_oeb[11]
port 253 nsew default output
rlabel metal2 s 145732 0 145788 800 6 io_oeb[12]
port 254 nsew default output
rlabel metal2 s 148676 0 148732 800 6 io_oeb[13]
port 255 nsew default output
rlabel metal2 s 151620 0 151676 800 6 io_oeb[14]
port 256 nsew default output
rlabel metal2 s 154472 0 154528 800 6 io_oeb[15]
port 257 nsew default output
rlabel metal2 s 157416 0 157472 800 6 io_oeb[16]
port 258 nsew default output
rlabel metal2 s 160268 0 160324 800 6 io_oeb[17]
port 259 nsew default output
rlabel metal2 s 163212 0 163268 800 6 io_oeb[18]
port 260 nsew default output
rlabel metal2 s 166156 0 166212 800 6 io_oeb[19]
port 261 nsew default output
rlabel metal2 s 113808 0 113864 800 6 io_oeb[1]
port 262 nsew default output
rlabel metal2 s 169008 0 169064 800 6 io_oeb[20]
port 263 nsew default output
rlabel metal2 s 171952 0 172008 800 6 io_oeb[21]
port 264 nsew default output
rlabel metal2 s 174804 0 174860 800 6 io_oeb[22]
port 265 nsew default output
rlabel metal2 s 177748 0 177804 800 6 io_oeb[23]
port 266 nsew default output
rlabel metal2 s 180692 0 180748 800 6 io_oeb[24]
port 267 nsew default output
rlabel metal2 s 183544 0 183600 800 6 io_oeb[25]
port 268 nsew default output
rlabel metal2 s 186488 0 186544 800 6 io_oeb[26]
port 269 nsew default output
rlabel metal2 s 189340 0 189396 800 6 io_oeb[27]
port 270 nsew default output
rlabel metal2 s 192284 0 192340 800 6 io_oeb[28]
port 271 nsew default output
rlabel metal2 s 195228 0 195284 800 6 io_oeb[29]
port 272 nsew default output
rlabel metal2 s 116660 0 116716 800 6 io_oeb[2]
port 273 nsew default output
rlabel metal2 s 198080 0 198136 800 6 io_oeb[30]
port 274 nsew default output
rlabel metal2 s 201024 0 201080 800 6 io_oeb[31]
port 275 nsew default output
rlabel metal2 s 203876 0 203932 800 6 io_oeb[32]
port 276 nsew default output
rlabel metal2 s 206820 0 206876 800 6 io_oeb[33]
port 277 nsew default output
rlabel metal2 s 209764 0 209820 800 6 io_oeb[34]
port 278 nsew default output
rlabel metal2 s 212616 0 212672 800 6 io_oeb[35]
port 279 nsew default output
rlabel metal2 s 215560 0 215616 800 6 io_oeb[36]
port 280 nsew default output
rlabel metal2 s 218412 0 218468 800 6 io_oeb[37]
port 281 nsew default output
rlabel metal2 s 119604 0 119660 800 6 io_oeb[3]
port 282 nsew default output
rlabel metal2 s 122548 0 122604 800 6 io_oeb[4]
port 283 nsew default output
rlabel metal2 s 125400 0 125456 800 6 io_oeb[5]
port 284 nsew default output
rlabel metal2 s 128344 0 128400 800 6 io_oeb[6]
port 285 nsew default output
rlabel metal2 s 131196 0 131252 800 6 io_oeb[7]
port 286 nsew default output
rlabel metal2 s 134140 0 134196 800 6 io_oeb[8]
port 287 nsew default output
rlabel metal2 s 137084 0 137140 800 6 io_oeb[9]
port 288 nsew default output
rlabel metal2 s 111876 0 111932 800 6 io_out[0]
port 289 nsew default output
rlabel metal2 s 140948 0 141004 800 6 io_out[10]
port 290 nsew default output
rlabel metal2 s 143800 0 143856 800 6 io_out[11]
port 291 nsew default output
rlabel metal2 s 146744 0 146800 800 6 io_out[12]
port 292 nsew default output
rlabel metal2 s 149688 0 149744 800 6 io_out[13]
port 293 nsew default output
rlabel metal2 s 152540 0 152596 800 6 io_out[14]
port 294 nsew default output
rlabel metal2 s 155484 0 155540 800 6 io_out[15]
port 295 nsew default output
rlabel metal2 s 158336 0 158392 800 6 io_out[16]
port 296 nsew default output
rlabel metal2 s 161280 0 161336 800 6 io_out[17]
port 297 nsew default output
rlabel metal2 s 164224 0 164280 800 6 io_out[18]
port 298 nsew default output
rlabel metal2 s 167076 0 167132 800 6 io_out[19]
port 299 nsew default output
rlabel metal2 s 114728 0 114784 800 6 io_out[1]
port 300 nsew default output
rlabel metal2 s 170020 0 170076 800 6 io_out[20]
port 301 nsew default output
rlabel metal2 s 172872 0 172928 800 6 io_out[21]
port 302 nsew default output
rlabel metal2 s 175816 0 175872 800 6 io_out[22]
port 303 nsew default output
rlabel metal2 s 178760 0 178816 800 6 io_out[23]
port 304 nsew default output
rlabel metal2 s 181612 0 181668 800 6 io_out[24]
port 305 nsew default output
rlabel metal2 s 184556 0 184612 800 6 io_out[25]
port 306 nsew default output
rlabel metal2 s 187408 0 187464 800 6 io_out[26]
port 307 nsew default output
rlabel metal2 s 190352 0 190408 800 6 io_out[27]
port 308 nsew default output
rlabel metal2 s 193296 0 193352 800 6 io_out[28]
port 309 nsew default output
rlabel metal2 s 196148 0 196204 800 6 io_out[29]
port 310 nsew default output
rlabel metal2 s 117672 0 117728 800 6 io_out[2]
port 311 nsew default output
rlabel metal2 s 199092 0 199148 800 6 io_out[30]
port 312 nsew default output
rlabel metal2 s 201944 0 202000 800 6 io_out[31]
port 313 nsew default output
rlabel metal2 s 204888 0 204944 800 6 io_out[32]
port 314 nsew default output
rlabel metal2 s 207832 0 207888 800 6 io_out[33]
port 315 nsew default output
rlabel metal2 s 210684 0 210740 800 6 io_out[34]
port 316 nsew default output
rlabel metal2 s 213628 0 213684 800 6 io_out[35]
port 317 nsew default output
rlabel metal2 s 216480 0 216536 800 6 io_out[36]
port 318 nsew default output
rlabel metal2 s 219424 0 219480 800 6 io_out[37]
port 319 nsew default output
rlabel metal2 s 120616 0 120672 800 6 io_out[3]
port 320 nsew default output
rlabel metal2 s 123468 0 123524 800 6 io_out[4]
port 321 nsew default output
rlabel metal2 s 126412 0 126468 800 6 io_out[5]
port 322 nsew default output
rlabel metal2 s 129264 0 129320 800 6 io_out[6]
port 323 nsew default output
rlabel metal2 s 132208 0 132264 800 6 io_out[7]
port 324 nsew default output
rlabel metal2 s 135152 0 135208 800 6 io_out[8]
port 325 nsew default output
rlabel metal2 s 138004 0 138060 800 6 io_out[9]
port 326 nsew default output
rlabel metal2 s 103136 0 103192 800 6 la_data_in[0]
port 327 nsew default input
rlabel metal2 s 106080 0 106136 800 6 la_data_in[1]
port 328 nsew default input
rlabel metal2 s 104148 0 104204 800 6 la_data_out[0]
port 329 nsew default output
rlabel metal2 s 107000 0 107056 800 6 la_data_out[1]
port 330 nsew default output
rlabel metal2 s 108932 0 108988 800 6 la_data_out[2]
port 331 nsew default output
rlabel metal2 s 105068 0 105124 800 6 la_oen[0]
port 332 nsew default input
rlabel metal2 s 108012 0 108068 800 6 la_oen[1]
port 333 nsew default input
rlabel metal3 s 219186 1368 219986 1488 6 one
port 334 nsew default output
rlabel metal3 s 219186 2320 219986 2440 6 ram_ce
port 335 nsew default output
rlabel metal3 s 219186 110440 219986 110560 6 sr0_ce
port 336 nsew default output
rlabel metal3 s 219186 111392 219986 111512 6 sr0_dtr[0]
port 337 nsew default input
rlabel metal3 s 219186 121456 219986 121576 6 sr0_dtr[10]
port 338 nsew default input
rlabel metal3 s 219186 122544 219986 122664 6 sr0_dtr[11]
port 339 nsew default input
rlabel metal3 s 219186 123496 219986 123616 6 sr0_dtr[12]
port 340 nsew default input
rlabel metal3 s 219186 124448 219986 124568 6 sr0_dtr[13]
port 341 nsew default input
rlabel metal3 s 219186 125536 219986 125656 6 sr0_dtr[14]
port 342 nsew default input
rlabel metal3 s 219186 126488 219986 126608 6 sr0_dtr[15]
port 343 nsew default input
rlabel metal3 s 219186 127576 219986 127696 6 sr0_dtr[16]
port 344 nsew default input
rlabel metal3 s 219186 128528 219986 128648 6 sr0_dtr[17]
port 345 nsew default input
rlabel metal3 s 219186 129616 219986 129736 6 sr0_dtr[18]
port 346 nsew default input
rlabel metal3 s 219186 130568 219986 130688 6 sr0_dtr[19]
port 347 nsew default input
rlabel metal3 s 219186 112344 219986 112464 6 sr0_dtr[1]
port 348 nsew default input
rlabel metal3 s 219186 131520 219986 131640 6 sr0_dtr[20]
port 349 nsew default input
rlabel metal3 s 219186 132608 219986 132728 6 sr0_dtr[21]
port 350 nsew default input
rlabel metal3 s 219186 133560 219986 133680 6 sr0_dtr[22]
port 351 nsew default input
rlabel metal3 s 219186 134648 219986 134768 6 sr0_dtr[23]
port 352 nsew default input
rlabel metal3 s 219186 135600 219986 135720 6 sr0_dtr[24]
port 353 nsew default input
rlabel metal3 s 219186 136552 219986 136672 6 sr0_dtr[25]
port 354 nsew default input
rlabel metal3 s 219186 137640 219986 137760 6 sr0_dtr[26]
port 355 nsew default input
rlabel metal3 s 219186 138592 219986 138712 6 sr0_dtr[27]
port 356 nsew default input
rlabel metal3 s 219186 139680 219986 139800 6 sr0_dtr[28]
port 357 nsew default input
rlabel metal3 s 219186 140632 219986 140752 6 sr0_dtr[29]
port 358 nsew default input
rlabel metal3 s 219186 113432 219986 113552 6 sr0_dtr[2]
port 359 nsew default input
rlabel metal3 s 219186 141720 219986 141840 6 sr0_dtr[30]
port 360 nsew default input
rlabel metal3 s 219186 142672 219986 142792 6 sr0_dtr[31]
port 361 nsew default input
rlabel metal3 s 219186 114384 219986 114504 6 sr0_dtr[3]
port 362 nsew default input
rlabel metal3 s 219186 115472 219986 115592 6 sr0_dtr[4]
port 363 nsew default input
rlabel metal3 s 219186 116424 219986 116544 6 sr0_dtr[5]
port 364 nsew default input
rlabel metal3 s 219186 117376 219986 117496 6 sr0_dtr[6]
port 365 nsew default input
rlabel metal3 s 219186 118464 219986 118584 6 sr0_dtr[7]
port 366 nsew default input
rlabel metal3 s 219186 119416 219986 119536 6 sr0_dtr[8]
port 367 nsew default input
rlabel metal3 s 219186 120504 219986 120624 6 sr0_dtr[9]
port 368 nsew default input
rlabel metal3 s 219186 143624 219986 143744 6 sr1_ce
port 369 nsew default output
rlabel metal3 s 219186 144712 219986 144832 6 sr1_dtr[0]
port 370 nsew default input
rlabel metal3 s 219186 154776 219986 154896 6 sr1_dtr[10]
port 371 nsew default input
rlabel metal3 s 219186 155728 219986 155848 6 sr1_dtr[11]
port 372 nsew default input
rlabel metal3 s 219186 156816 219986 156936 6 sr1_dtr[12]
port 373 nsew default input
rlabel metal3 s 219186 157768 219986 157888 6 sr1_dtr[13]
port 374 nsew default input
rlabel metal3 s 219186 158856 219986 158976 6 sr1_dtr[14]
port 375 nsew default input
rlabel metal3 s 219186 159808 219986 159928 6 sr1_dtr[15]
port 376 nsew default input
rlabel metal3 s 219186 160896 219986 161016 6 sr1_dtr[16]
port 377 nsew default input
rlabel metal3 s 219186 161848 219986 161968 6 sr1_dtr[17]
port 378 nsew default input
rlabel metal3 s 219186 162800 219986 162920 6 sr1_dtr[18]
port 379 nsew default input
rlabel metal3 s 219186 163888 219986 164008 6 sr1_dtr[19]
port 380 nsew default input
rlabel metal3 s 219186 145664 219986 145784 6 sr1_dtr[1]
port 381 nsew default input
rlabel metal3 s 219186 164840 219986 164960 6 sr1_dtr[20]
port 382 nsew default input
rlabel metal3 s 219186 165928 219986 166048 6 sr1_dtr[21]
port 383 nsew default input
rlabel metal3 s 219186 166880 219986 167000 6 sr1_dtr[22]
port 384 nsew default input
rlabel metal3 s 219186 167968 219986 168088 6 sr1_dtr[23]
port 385 nsew default input
rlabel metal3 s 219186 168920 219986 169040 6 sr1_dtr[24]
port 386 nsew default input
rlabel metal3 s 219186 169872 219986 169992 6 sr1_dtr[25]
port 387 nsew default input
rlabel metal3 s 219186 170960 219986 171080 6 sr1_dtr[26]
port 388 nsew default input
rlabel metal3 s 219186 171912 219986 172032 6 sr1_dtr[27]
port 389 nsew default input
rlabel metal3 s 219186 173000 219986 173120 6 sr1_dtr[28]
port 390 nsew default input
rlabel metal3 s 219186 173952 219986 174072 6 sr1_dtr[29]
port 391 nsew default input
rlabel metal3 s 219186 146752 219986 146872 6 sr1_dtr[2]
port 392 nsew default input
rlabel metal3 s 219186 175040 219986 175160 6 sr1_dtr[30]
port 393 nsew default input
rlabel metal3 s 219186 175992 219986 176112 6 sr1_dtr[31]
port 394 nsew default input
rlabel metal3 s 219186 147704 219986 147824 6 sr1_dtr[3]
port 395 nsew default input
rlabel metal3 s 219186 148792 219986 148912 6 sr1_dtr[4]
port 396 nsew default input
rlabel metal3 s 219186 149744 219986 149864 6 sr1_dtr[5]
port 397 nsew default input
rlabel metal3 s 219186 150696 219986 150816 6 sr1_dtr[6]
port 398 nsew default input
rlabel metal3 s 219186 151784 219986 151904 6 sr1_dtr[7]
port 399 nsew default input
rlabel metal3 s 219186 152736 219986 152856 6 sr1_dtr[8]
port 400 nsew default input
rlabel metal3 s 219186 153824 219986 153944 6 sr1_dtr[9]
port 401 nsew default input
rlabel metal3 s 219186 178032 219986 178152 6 srx_addr[0]
port 402 nsew default output
rlabel metal3 s 219186 180072 219986 180192 6 srx_addr[1]
port 403 nsew default output
rlabel metal3 s 219186 181976 219986 182096 6 srx_addr[2]
port 404 nsew default output
rlabel metal3 s 219186 184016 219986 184136 6 srx_addr[3]
port 405 nsew default output
rlabel metal3 s 219186 186056 219986 186176 6 srx_addr[4]
port 406 nsew default output
rlabel metal3 s 219186 188096 219986 188216 6 srx_addr[5]
port 407 nsew default output
rlabel metal3 s 219186 190136 219986 190256 6 srx_addr[6]
port 408 nsew default output
rlabel metal3 s 219186 192176 219986 192296 6 srx_addr[7]
port 409 nsew default output
rlabel metal3 s 219186 194216 219986 194336 6 srx_addr[8]
port 410 nsew default output
rlabel metal3 s 219186 196120 219986 196240 6 srx_addr[9]
port 411 nsew default output
rlabel metal3 s 219186 178984 219986 179104 6 srx_dtw[0]
port 412 nsew default output
rlabel metal3 s 219186 198160 219986 198280 6 srx_dtw[10]
port 413 nsew default output
rlabel metal3 s 219186 199248 219986 199368 6 srx_dtw[11]
port 414 nsew default output
rlabel metal3 s 219186 200200 219986 200320 6 srx_dtw[12]
port 415 nsew default output
rlabel metal3 s 219186 201152 219986 201272 6 srx_dtw[13]
port 416 nsew default output
rlabel metal3 s 219186 202240 219986 202360 6 srx_dtw[14]
port 417 nsew default output
rlabel metal3 s 219186 203192 219986 203312 6 srx_dtw[15]
port 418 nsew default output
rlabel metal3 s 219186 204280 219986 204400 6 srx_dtw[16]
port 419 nsew default output
rlabel metal3 s 219186 205232 219986 205352 6 srx_dtw[17]
port 420 nsew default output
rlabel metal3 s 219186 206320 219986 206440 6 srx_dtw[18]
port 421 nsew default output
rlabel metal3 s 219186 207272 219986 207392 6 srx_dtw[19]
port 422 nsew default output
rlabel metal3 s 219186 181024 219986 181144 6 srx_dtw[1]
port 423 nsew default output
rlabel metal3 s 219186 208224 219986 208344 6 srx_dtw[20]
port 424 nsew default output
rlabel metal3 s 219186 209312 219986 209432 6 srx_dtw[21]
port 425 nsew default output
rlabel metal3 s 219186 210264 219986 210384 6 srx_dtw[22]
port 426 nsew default output
rlabel metal3 s 219186 211352 219986 211472 6 srx_dtw[23]
port 427 nsew default output
rlabel metal3 s 219186 212304 219986 212424 6 srx_dtw[24]
port 428 nsew default output
rlabel metal3 s 219186 213392 219986 213512 6 srx_dtw[25]
port 429 nsew default output
rlabel metal3 s 219186 214344 219986 214464 6 srx_dtw[26]
port 430 nsew default output
rlabel metal3 s 219186 215296 219986 215416 6 srx_dtw[27]
port 431 nsew default output
rlabel metal3 s 219186 216384 219986 216504 6 srx_dtw[28]
port 432 nsew default output
rlabel metal3 s 219186 217336 219986 217456 6 srx_dtw[29]
port 433 nsew default output
rlabel metal3 s 219186 183064 219986 183184 6 srx_dtw[2]
port 434 nsew default output
rlabel metal3 s 219186 218424 219986 218544 6 srx_dtw[30]
port 435 nsew default output
rlabel metal3 s 219186 219376 219986 219496 6 srx_dtw[31]
port 436 nsew default output
rlabel metal3 s 219186 185104 219986 185224 6 srx_dtw[3]
port 437 nsew default output
rlabel metal3 s 219186 187144 219986 187264 6 srx_dtw[4]
port 438 nsew default output
rlabel metal3 s 219186 189048 219986 189168 6 srx_dtw[5]
port 439 nsew default output
rlabel metal3 s 219186 191088 219986 191208 6 srx_dtw[6]
port 440 nsew default output
rlabel metal3 s 219186 193128 219986 193248 6 srx_dtw[7]
port 441 nsew default output
rlabel metal3 s 219186 195168 219986 195288 6 srx_dtw[8]
port 442 nsew default output
rlabel metal3 s 219186 197208 219986 197328 6 srx_dtw[9]
port 443 nsew default output
rlabel metal3 s 219186 176944 219986 177064 6 srx_we
port 444 nsew default output
rlabel metal2 s 464 0 520 800 6 wb_clk_i
port 445 nsew default input
rlabel metal2 s 1384 0 1440 800 6 wb_rst_i
port 446 nsew default input
rlabel metal2 s 2396 0 2452 800 6 wbs_ack_o
port 447 nsew default output
rlabel metal2 s 6260 0 6316 800 6 wbs_adr_i[0]
port 448 nsew default input
rlabel metal2 s 39196 0 39252 800 6 wbs_adr_i[10]
port 449 nsew default input
rlabel metal2 s 42048 0 42104 800 6 wbs_adr_i[11]
port 450 nsew default input
rlabel metal2 s 44992 0 45048 800 6 wbs_adr_i[12]
port 451 nsew default input
rlabel metal2 s 47936 0 47992 800 6 wbs_adr_i[13]
port 452 nsew default input
rlabel metal2 s 50788 0 50844 800 6 wbs_adr_i[14]
port 453 nsew default input
rlabel metal2 s 53732 0 53788 800 6 wbs_adr_i[15]
port 454 nsew default input
rlabel metal2 s 56584 0 56640 800 6 wbs_adr_i[16]
port 455 nsew default input
rlabel metal2 s 59528 0 59584 800 6 wbs_adr_i[17]
port 456 nsew default input
rlabel metal2 s 62472 0 62528 800 6 wbs_adr_i[18]
port 457 nsew default input
rlabel metal2 s 65324 0 65380 800 6 wbs_adr_i[19]
port 458 nsew default input
rlabel metal2 s 10124 0 10180 800 6 wbs_adr_i[1]
port 459 nsew default input
rlabel metal2 s 68268 0 68324 800 6 wbs_adr_i[20]
port 460 nsew default input
rlabel metal2 s 71120 0 71176 800 6 wbs_adr_i[21]
port 461 nsew default input
rlabel metal2 s 74064 0 74120 800 6 wbs_adr_i[22]
port 462 nsew default input
rlabel metal2 s 77008 0 77064 800 6 wbs_adr_i[23]
port 463 nsew default input
rlabel metal2 s 79860 0 79916 800 6 wbs_adr_i[24]
port 464 nsew default input
rlabel metal2 s 82804 0 82860 800 6 wbs_adr_i[25]
port 465 nsew default input
rlabel metal2 s 85656 0 85712 800 6 wbs_adr_i[26]
port 466 nsew default input
rlabel metal2 s 88600 0 88656 800 6 wbs_adr_i[27]
port 467 nsew default input
rlabel metal2 s 91544 0 91600 800 6 wbs_adr_i[28]
port 468 nsew default input
rlabel metal2 s 94396 0 94452 800 6 wbs_adr_i[29]
port 469 nsew default input
rlabel metal2 s 13988 0 14044 800 6 wbs_adr_i[2]
port 470 nsew default input
rlabel metal2 s 97340 0 97396 800 6 wbs_adr_i[30]
port 471 nsew default input
rlabel metal2 s 100192 0 100248 800 6 wbs_adr_i[31]
port 472 nsew default input
rlabel metal2 s 17852 0 17908 800 6 wbs_adr_i[3]
port 473 nsew default input
rlabel metal2 s 21716 0 21772 800 6 wbs_adr_i[4]
port 474 nsew default input
rlabel metal2 s 24660 0 24716 800 6 wbs_adr_i[5]
port 475 nsew default input
rlabel metal2 s 27512 0 27568 800 6 wbs_adr_i[6]
port 476 nsew default input
rlabel metal2 s 30456 0 30512 800 6 wbs_adr_i[7]
port 477 nsew default input
rlabel metal2 s 33400 0 33456 800 6 wbs_adr_i[8]
port 478 nsew default input
rlabel metal2 s 36252 0 36308 800 6 wbs_adr_i[9]
port 479 nsew default input
rlabel metal2 s 3316 0 3372 800 6 wbs_cyc_i
port 480 nsew default input
rlabel metal2 s 7180 0 7236 800 6 wbs_dat_i[0]
port 481 nsew default input
rlabel metal2 s 40116 0 40172 800 6 wbs_dat_i[10]
port 482 nsew default input
rlabel metal2 s 43060 0 43116 800 6 wbs_dat_i[11]
port 483 nsew default input
rlabel metal2 s 46004 0 46060 800 6 wbs_dat_i[12]
port 484 nsew default input
rlabel metal2 s 48856 0 48912 800 6 wbs_dat_i[13]
port 485 nsew default input
rlabel metal2 s 51800 0 51856 800 6 wbs_dat_i[14]
port 486 nsew default input
rlabel metal2 s 54652 0 54708 800 6 wbs_dat_i[15]
port 487 nsew default input
rlabel metal2 s 57596 0 57652 800 6 wbs_dat_i[16]
port 488 nsew default input
rlabel metal2 s 60540 0 60596 800 6 wbs_dat_i[17]
port 489 nsew default input
rlabel metal2 s 63392 0 63448 800 6 wbs_dat_i[18]
port 490 nsew default input
rlabel metal2 s 66336 0 66392 800 6 wbs_dat_i[19]
port 491 nsew default input
rlabel metal2 s 11044 0 11100 800 6 wbs_dat_i[1]
port 492 nsew default input
rlabel metal2 s 69188 0 69244 800 6 wbs_dat_i[20]
port 493 nsew default input
rlabel metal2 s 72132 0 72188 800 6 wbs_dat_i[21]
port 494 nsew default input
rlabel metal2 s 75076 0 75132 800 6 wbs_dat_i[22]
port 495 nsew default input
rlabel metal2 s 77928 0 77984 800 6 wbs_dat_i[23]
port 496 nsew default input
rlabel metal2 s 80872 0 80928 800 6 wbs_dat_i[24]
port 497 nsew default input
rlabel metal2 s 83724 0 83780 800 6 wbs_dat_i[25]
port 498 nsew default input
rlabel metal2 s 86668 0 86724 800 6 wbs_dat_i[26]
port 499 nsew default input
rlabel metal2 s 89612 0 89668 800 6 wbs_dat_i[27]
port 500 nsew default input
rlabel metal2 s 92464 0 92520 800 6 wbs_dat_i[28]
port 501 nsew default input
rlabel metal2 s 95408 0 95464 800 6 wbs_dat_i[29]
port 502 nsew default input
rlabel metal2 s 14908 0 14964 800 6 wbs_dat_i[2]
port 503 nsew default input
rlabel metal2 s 98260 0 98316 800 6 wbs_dat_i[30]
port 504 nsew default input
rlabel metal2 s 101204 0 101260 800 6 wbs_dat_i[31]
port 505 nsew default input
rlabel metal2 s 18864 0 18920 800 6 wbs_dat_i[3]
port 506 nsew default input
rlabel metal2 s 22728 0 22784 800 6 wbs_dat_i[4]
port 507 nsew default input
rlabel metal2 s 25580 0 25636 800 6 wbs_dat_i[5]
port 508 nsew default input
rlabel metal2 s 28524 0 28580 800 6 wbs_dat_i[6]
port 509 nsew default input
rlabel metal2 s 31468 0 31524 800 6 wbs_dat_i[7]
port 510 nsew default input
rlabel metal2 s 34320 0 34376 800 6 wbs_dat_i[8]
port 511 nsew default input
rlabel metal2 s 37264 0 37320 800 6 wbs_dat_i[9]
port 512 nsew default input
rlabel metal2 s 8192 0 8248 800 6 wbs_dat_o[0]
port 513 nsew default output
rlabel metal2 s 41128 0 41184 800 6 wbs_dat_o[10]
port 514 nsew default output
rlabel metal2 s 43980 0 44036 800 6 wbs_dat_o[11]
port 515 nsew default output
rlabel metal2 s 46924 0 46980 800 6 wbs_dat_o[12]
port 516 nsew default output
rlabel metal2 s 49868 0 49924 800 6 wbs_dat_o[13]
port 517 nsew default output
rlabel metal2 s 52720 0 52776 800 6 wbs_dat_o[14]
port 518 nsew default output
rlabel metal2 s 55664 0 55720 800 6 wbs_dat_o[15]
port 519 nsew default output
rlabel metal2 s 58516 0 58572 800 6 wbs_dat_o[16]
port 520 nsew default output
rlabel metal2 s 61460 0 61516 800 6 wbs_dat_o[17]
port 521 nsew default output
rlabel metal2 s 64404 0 64460 800 6 wbs_dat_o[18]
port 522 nsew default output
rlabel metal2 s 67256 0 67312 800 6 wbs_dat_o[19]
port 523 nsew default output
rlabel metal2 s 12056 0 12112 800 6 wbs_dat_o[1]
port 524 nsew default output
rlabel metal2 s 70200 0 70256 800 6 wbs_dat_o[20]
port 525 nsew default output
rlabel metal2 s 73052 0 73108 800 6 wbs_dat_o[21]
port 526 nsew default output
rlabel metal2 s 75996 0 76052 800 6 wbs_dat_o[22]
port 527 nsew default output
rlabel metal2 s 78940 0 78996 800 6 wbs_dat_o[23]
port 528 nsew default output
rlabel metal2 s 81792 0 81848 800 6 wbs_dat_o[24]
port 529 nsew default output
rlabel metal2 s 84736 0 84792 800 6 wbs_dat_o[25]
port 530 nsew default output
rlabel metal2 s 87588 0 87644 800 6 wbs_dat_o[26]
port 531 nsew default output
rlabel metal2 s 90532 0 90588 800 6 wbs_dat_o[27]
port 532 nsew default output
rlabel metal2 s 93476 0 93532 800 6 wbs_dat_o[28]
port 533 nsew default output
rlabel metal2 s 96328 0 96384 800 6 wbs_dat_o[29]
port 534 nsew default output
rlabel metal2 s 15920 0 15976 800 6 wbs_dat_o[2]
port 535 nsew default output
rlabel metal2 s 99272 0 99328 800 6 wbs_dat_o[30]
port 536 nsew default output
rlabel metal2 s 102124 0 102180 800 6 wbs_dat_o[31]
port 537 nsew default output
rlabel metal2 s 19784 0 19840 800 6 wbs_dat_o[3]
port 538 nsew default output
rlabel metal2 s 23648 0 23704 800 6 wbs_dat_o[4]
port 539 nsew default output
rlabel metal2 s 26592 0 26648 800 6 wbs_dat_o[5]
port 540 nsew default output
rlabel metal2 s 29444 0 29500 800 6 wbs_dat_o[6]
port 541 nsew default output
rlabel metal2 s 32388 0 32444 800 6 wbs_dat_o[7]
port 542 nsew default output
rlabel metal2 s 35332 0 35388 800 6 wbs_dat_o[8]
port 543 nsew default output
rlabel metal2 s 38184 0 38240 800 6 wbs_dat_o[9]
port 544 nsew default output
rlabel metal2 s 9112 0 9168 800 6 wbs_sel_i[0]
port 545 nsew default input
rlabel metal2 s 12976 0 13032 800 6 wbs_sel_i[1]
port 546 nsew default input
rlabel metal2 s 16932 0 16988 800 6 wbs_sel_i[2]
port 547 nsew default input
rlabel metal2 s 20796 0 20852 800 6 wbs_sel_i[3]
port 548 nsew default input
rlabel metal2 s 4328 0 4384 800 6 wbs_stb_i
port 549 nsew default input
rlabel metal2 s 5248 0 5304 800 6 wbs_we_i
port 550 nsew default input
rlabel metal3 s 219186 416 219986 536 6 zero
port 551 nsew default output
rlabel metal4 s 4194 2128 4514 217648 6 VPWR
port 552 nsew power input
rlabel metal4 s 19554 2128 19874 217648 6 VGND
port 553 nsew ground input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 219986 220000
string LEFview TRUE
<< end >>
