VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 28.980 2924.800 30.180 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2374.980 2924.800 2376.180 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2609.580 2924.800 2610.780 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2844.180 2924.800 2845.380 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3078.780 2924.800 3079.980 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3313.380 2924.800 3314.580 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 263.580 2924.800 264.780 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3482.700 2.400 3483.900 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3195.060 2.400 3196.260 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2908.100 2.400 2909.300 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2620.460 2.400 2621.660 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2333.500 2.400 2334.700 ;
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2045.860 2.400 2047.060 ;
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 498.180 2924.800 499.380 ;
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1758.900 2.400 1760.100 ;
    END
  END analog_io[30]
  PIN analog_io[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 732.780 2924.800 733.980 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 967.380 2924.800 968.580 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1201.980 2924.800 1203.180 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1436.580 2924.800 1437.780 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1671.180 2924.800 1672.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1905.780 2924.800 1906.980 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2140.380 2924.800 2141.580 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 288.950 89.660 289.270 89.720 ;
        RECT 2898.990 89.660 2899.310 89.720 ;
        RECT 288.950 89.520 2899.310 89.660 ;
        RECT 288.950 89.460 289.270 89.520 ;
        RECT 2898.990 89.460 2899.310 89.520 ;
      LAYER via ;
        RECT 288.980 89.460 289.240 89.720 ;
        RECT 2899.020 89.460 2899.280 89.720 ;
      LAYER met2 ;
        RECT 288.970 1005.195 289.250 1005.565 ;
        RECT 289.040 89.750 289.180 1005.195 ;
        RECT 288.980 89.430 289.240 89.750 ;
        RECT 2899.020 89.430 2899.280 89.750 ;
        RECT 2899.080 88.245 2899.220 89.430 ;
        RECT 2899.010 87.875 2899.290 88.245 ;
      LAYER via2 ;
        RECT 288.970 1005.240 289.250 1005.520 ;
        RECT 2899.010 87.920 2899.290 88.200 ;
      LAYER met3 ;
        RECT 288.945 1005.530 289.275 1005.545 ;
        RECT 288.945 1005.400 300.380 1005.530 ;
        RECT 288.945 1005.230 304.000 1005.400 ;
        RECT 288.945 1005.215 289.275 1005.230 ;
        RECT 300.000 1004.800 304.000 1005.230 ;
        RECT 2898.985 88.210 2899.315 88.225 ;
        RECT 2917.600 88.210 2924.800 88.660 ;
        RECT 2898.985 87.910 2924.800 88.210 ;
        RECT 2898.985 87.895 2899.315 87.910 ;
        RECT 2917.600 87.460 2924.800 87.910 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 290.330 2197.660 290.650 2197.720 ;
        RECT 2903.590 2197.660 2903.910 2197.720 ;
        RECT 290.330 2197.520 2903.910 2197.660 ;
        RECT 290.330 2197.460 290.650 2197.520 ;
        RECT 2903.590 2197.460 2903.910 2197.520 ;
      LAYER via ;
        RECT 290.360 2197.460 290.620 2197.720 ;
        RECT 2903.620 2197.460 2903.880 2197.720 ;
      LAYER met2 ;
        RECT 2903.610 2433.875 2903.890 2434.245 ;
        RECT 2903.680 2197.750 2903.820 2433.875 ;
        RECT 290.360 2197.430 290.620 2197.750 ;
        RECT 2903.620 2197.430 2903.880 2197.750 ;
        RECT 290.420 1321.085 290.560 2197.430 ;
        RECT 290.350 1320.715 290.630 1321.085 ;
      LAYER via2 ;
        RECT 2903.610 2433.920 2903.890 2434.200 ;
        RECT 290.350 1320.760 290.630 1321.040 ;
      LAYER met3 ;
        RECT 2903.585 2434.210 2903.915 2434.225 ;
        RECT 2917.600 2434.210 2924.800 2434.660 ;
        RECT 2903.585 2433.910 2924.800 2434.210 ;
        RECT 2903.585 2433.895 2903.915 2433.910 ;
        RECT 2917.600 2433.460 2924.800 2433.910 ;
        RECT 290.325 1321.050 290.655 1321.065 ;
        RECT 290.325 1320.920 300.380 1321.050 ;
        RECT 290.325 1320.750 304.000 1320.920 ;
        RECT 290.325 1320.735 290.655 1320.750 ;
        RECT 300.000 1320.320 304.000 1320.750 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 289.870 2198.000 290.190 2198.060 ;
        RECT 2901.750 2198.000 2902.070 2198.060 ;
        RECT 289.870 2197.860 2902.070 2198.000 ;
        RECT 289.870 2197.800 290.190 2197.860 ;
        RECT 2901.750 2197.800 2902.070 2197.860 ;
      LAYER via ;
        RECT 289.900 2197.800 290.160 2198.060 ;
        RECT 2901.780 2197.800 2902.040 2198.060 ;
      LAYER met2 ;
        RECT 2901.770 2669.155 2902.050 2669.525 ;
        RECT 2901.840 2198.090 2901.980 2669.155 ;
        RECT 289.900 2197.770 290.160 2198.090 ;
        RECT 2901.780 2197.770 2902.040 2198.090 ;
        RECT 289.960 1352.365 290.100 2197.770 ;
        RECT 289.890 1351.995 290.170 1352.365 ;
      LAYER via2 ;
        RECT 2901.770 2669.200 2902.050 2669.480 ;
        RECT 289.890 1352.040 290.170 1352.320 ;
      LAYER met3 ;
        RECT 2901.745 2669.490 2902.075 2669.505 ;
        RECT 2917.600 2669.490 2924.800 2669.940 ;
        RECT 2901.745 2669.190 2924.800 2669.490 ;
        RECT 2901.745 2669.175 2902.075 2669.190 ;
        RECT 2917.600 2668.740 2924.800 2669.190 ;
        RECT 289.865 1352.330 290.195 1352.345 ;
        RECT 289.865 1352.200 300.380 1352.330 ;
        RECT 289.865 1352.030 304.000 1352.200 ;
        RECT 289.865 1352.015 290.195 1352.030 ;
        RECT 300.000 1351.600 304.000 1352.030 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 291.710 2898.400 292.030 2898.460 ;
        RECT 2900.830 2898.400 2901.150 2898.460 ;
        RECT 291.710 2898.260 2901.150 2898.400 ;
        RECT 291.710 2898.200 292.030 2898.260 ;
        RECT 2900.830 2898.200 2901.150 2898.260 ;
      LAYER via ;
        RECT 291.740 2898.200 292.000 2898.460 ;
        RECT 2900.860 2898.200 2901.120 2898.460 ;
      LAYER met2 ;
        RECT 2900.850 2903.755 2901.130 2904.125 ;
        RECT 2900.920 2898.490 2901.060 2903.755 ;
        RECT 291.740 2898.170 292.000 2898.490 ;
        RECT 2900.860 2898.170 2901.120 2898.490 ;
        RECT 291.800 1384.325 291.940 2898.170 ;
        RECT 291.730 1383.955 292.010 1384.325 ;
      LAYER via2 ;
        RECT 2900.850 2903.800 2901.130 2904.080 ;
        RECT 291.730 1384.000 292.010 1384.280 ;
      LAYER met3 ;
        RECT 2900.825 2904.090 2901.155 2904.105 ;
        RECT 2917.600 2904.090 2924.800 2904.540 ;
        RECT 2900.825 2903.790 2924.800 2904.090 ;
        RECT 2900.825 2903.775 2901.155 2903.790 ;
        RECT 2917.600 2903.340 2924.800 2903.790 ;
        RECT 291.705 1384.290 292.035 1384.305 ;
        RECT 291.705 1384.160 300.380 1384.290 ;
        RECT 291.705 1383.990 304.000 1384.160 ;
        RECT 291.705 1383.975 292.035 1383.990 ;
        RECT 300.000 1383.560 304.000 1383.990 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2801.470 3135.040 2801.790 3135.100 ;
        RECT 2825.850 3135.040 2826.170 3135.100 ;
        RECT 2801.470 3134.900 2826.170 3135.040 ;
        RECT 2801.470 3134.840 2801.790 3134.900 ;
        RECT 2825.850 3134.840 2826.170 3134.900 ;
        RECT 1449.070 3134.360 1449.390 3134.420 ;
        RECT 1463.330 3134.360 1463.650 3134.420 ;
        RECT 1449.070 3134.220 1463.650 3134.360 ;
        RECT 1449.070 3134.160 1449.390 3134.220 ;
        RECT 1463.330 3134.160 1463.650 3134.220 ;
        RECT 2125.270 3134.360 2125.590 3134.420 ;
        RECT 2139.530 3134.360 2139.850 3134.420 ;
        RECT 2125.270 3134.220 2139.850 3134.360 ;
        RECT 2125.270 3134.160 2125.590 3134.220 ;
        RECT 2139.530 3134.160 2139.850 3134.220 ;
        RECT 2704.870 3134.360 2705.190 3134.420 ;
        RECT 2743.050 3134.360 2743.370 3134.420 ;
        RECT 2704.870 3134.220 2743.370 3134.360 ;
        RECT 2704.870 3134.160 2705.190 3134.220 ;
        RECT 2743.050 3134.160 2743.370 3134.220 ;
      LAYER via ;
        RECT 2801.500 3134.840 2801.760 3135.100 ;
        RECT 2825.880 3134.840 2826.140 3135.100 ;
        RECT 1449.100 3134.160 1449.360 3134.420 ;
        RECT 1463.360 3134.160 1463.620 3134.420 ;
        RECT 2125.300 3134.160 2125.560 3134.420 ;
        RECT 2139.560 3134.160 2139.820 3134.420 ;
        RECT 2704.900 3134.160 2705.160 3134.420 ;
        RECT 2743.080 3134.160 2743.340 3134.420 ;
      LAYER met2 ;
        RECT 2766.530 3135.210 2766.810 3135.325 ;
        RECT 2767.450 3135.210 2767.730 3135.325 ;
        RECT 2766.530 3135.070 2767.730 3135.210 ;
        RECT 2766.530 3134.955 2766.810 3135.070 ;
        RECT 2767.450 3134.955 2767.730 3135.070 ;
        RECT 2801.490 3134.955 2801.770 3135.325 ;
        RECT 2801.500 3134.810 2801.760 3134.955 ;
        RECT 2825.880 3134.810 2826.140 3135.130 ;
        RECT 2825.940 3134.645 2826.080 3134.810 ;
        RECT 1449.090 3134.275 1449.370 3134.645 ;
        RECT 1449.100 3134.130 1449.360 3134.275 ;
        RECT 1463.360 3134.130 1463.620 3134.450 ;
        RECT 2125.290 3134.275 2125.570 3134.645 ;
        RECT 2125.300 3134.130 2125.560 3134.275 ;
        RECT 2139.560 3134.130 2139.820 3134.450 ;
        RECT 2704.890 3134.275 2705.170 3134.645 ;
        RECT 2704.900 3134.130 2705.160 3134.275 ;
        RECT 2743.080 3134.130 2743.340 3134.450 ;
        RECT 2825.870 3134.275 2826.150 3134.645 ;
        RECT 2863.590 3134.530 2863.870 3134.645 ;
        RECT 2863.200 3134.390 2863.870 3134.530 ;
        RECT 1463.420 3133.285 1463.560 3134.130 ;
        RECT 2139.620 3133.285 2139.760 3134.130 ;
        RECT 2743.140 3133.285 2743.280 3134.130 ;
        RECT 2863.200 3133.965 2863.340 3134.390 ;
        RECT 2863.590 3134.275 2863.870 3134.390 ;
        RECT 2863.130 3133.595 2863.410 3133.965 ;
        RECT 1463.350 3132.915 1463.630 3133.285 ;
        RECT 2139.550 3132.915 2139.830 3133.285 ;
        RECT 2743.070 3132.915 2743.350 3133.285 ;
      LAYER via2 ;
        RECT 2766.530 3135.000 2766.810 3135.280 ;
        RECT 2767.450 3135.000 2767.730 3135.280 ;
        RECT 2801.490 3135.000 2801.770 3135.280 ;
        RECT 1449.090 3134.320 1449.370 3134.600 ;
        RECT 2125.290 3134.320 2125.570 3134.600 ;
        RECT 2704.890 3134.320 2705.170 3134.600 ;
        RECT 2825.870 3134.320 2826.150 3134.600 ;
        RECT 2863.590 3134.320 2863.870 3134.600 ;
        RECT 2863.130 3133.640 2863.410 3133.920 ;
        RECT 1463.350 3132.960 1463.630 3133.240 ;
        RECT 2139.550 3132.960 2139.830 3133.240 ;
        RECT 2743.070 3132.960 2743.350 3133.240 ;
      LAYER met3 ;
        RECT 2917.600 3138.690 2924.800 3139.140 ;
        RECT 2916.710 3138.390 2924.800 3138.690 ;
        RECT 2752.910 3135.290 2753.290 3135.300 ;
        RECT 2766.505 3135.290 2766.835 3135.305 ;
        RECT 2752.910 3134.990 2766.835 3135.290 ;
        RECT 2752.910 3134.980 2753.290 3134.990 ;
        RECT 2766.505 3134.975 2766.835 3134.990 ;
        RECT 2767.425 3135.290 2767.755 3135.305 ;
        RECT 2801.465 3135.290 2801.795 3135.305 ;
        RECT 2767.425 3134.990 2801.795 3135.290 ;
        RECT 2767.425 3134.975 2767.755 3134.990 ;
        RECT 2801.465 3134.975 2801.795 3134.990 ;
        RECT 290.070 3134.610 290.450 3134.620 ;
        RECT 1449.065 3134.610 1449.395 3134.625 ;
        RECT 290.070 3134.310 324.450 3134.610 ;
        RECT 290.070 3134.300 290.450 3134.310 ;
        RECT 324.150 3133.930 324.450 3134.310 ;
        RECT 372.910 3134.310 421.050 3134.610 ;
        RECT 324.150 3133.630 372.290 3133.930 ;
        RECT 371.990 3133.250 372.290 3133.630 ;
        RECT 372.910 3133.250 373.210 3134.310 ;
        RECT 420.750 3133.930 421.050 3134.310 ;
        RECT 469.510 3134.310 517.650 3134.610 ;
        RECT 420.750 3133.630 468.890 3133.930 ;
        RECT 371.990 3132.950 373.210 3133.250 ;
        RECT 468.590 3133.250 468.890 3133.630 ;
        RECT 469.510 3133.250 469.810 3134.310 ;
        RECT 517.350 3133.930 517.650 3134.310 ;
        RECT 566.110 3134.310 614.250 3134.610 ;
        RECT 517.350 3133.630 565.490 3133.930 ;
        RECT 468.590 3132.950 469.810 3133.250 ;
        RECT 565.190 3133.250 565.490 3133.630 ;
        RECT 566.110 3133.250 566.410 3134.310 ;
        RECT 613.950 3133.930 614.250 3134.310 ;
        RECT 662.710 3134.310 710.850 3134.610 ;
        RECT 613.950 3133.630 662.090 3133.930 ;
        RECT 565.190 3132.950 566.410 3133.250 ;
        RECT 661.790 3133.250 662.090 3133.630 ;
        RECT 662.710 3133.250 663.010 3134.310 ;
        RECT 710.550 3133.930 710.850 3134.310 ;
        RECT 759.310 3134.310 807.450 3134.610 ;
        RECT 710.550 3133.630 758.690 3133.930 ;
        RECT 661.790 3132.950 663.010 3133.250 ;
        RECT 758.390 3133.250 758.690 3133.630 ;
        RECT 759.310 3133.250 759.610 3134.310 ;
        RECT 807.150 3133.930 807.450 3134.310 ;
        RECT 855.910 3134.310 904.050 3134.610 ;
        RECT 807.150 3133.630 855.290 3133.930 ;
        RECT 758.390 3132.950 759.610 3133.250 ;
        RECT 854.990 3133.250 855.290 3133.630 ;
        RECT 855.910 3133.250 856.210 3134.310 ;
        RECT 903.750 3133.930 904.050 3134.310 ;
        RECT 952.510 3134.310 1000.650 3134.610 ;
        RECT 903.750 3133.630 951.890 3133.930 ;
        RECT 854.990 3132.950 856.210 3133.250 ;
        RECT 951.590 3133.250 951.890 3133.630 ;
        RECT 952.510 3133.250 952.810 3134.310 ;
        RECT 1000.350 3133.930 1000.650 3134.310 ;
        RECT 1049.110 3134.310 1097.250 3134.610 ;
        RECT 1000.350 3133.630 1048.490 3133.930 ;
        RECT 951.590 3132.950 952.810 3133.250 ;
        RECT 1048.190 3133.250 1048.490 3133.630 ;
        RECT 1049.110 3133.250 1049.410 3134.310 ;
        RECT 1096.950 3133.930 1097.250 3134.310 ;
        RECT 1145.710 3134.310 1193.850 3134.610 ;
        RECT 1096.950 3133.630 1145.090 3133.930 ;
        RECT 1048.190 3132.950 1049.410 3133.250 ;
        RECT 1144.790 3133.250 1145.090 3133.630 ;
        RECT 1145.710 3133.250 1146.010 3134.310 ;
        RECT 1193.550 3133.930 1193.850 3134.310 ;
        RECT 1242.310 3134.310 1290.450 3134.610 ;
        RECT 1193.550 3133.630 1241.690 3133.930 ;
        RECT 1144.790 3132.950 1146.010 3133.250 ;
        RECT 1241.390 3133.250 1241.690 3133.630 ;
        RECT 1242.310 3133.250 1242.610 3134.310 ;
        RECT 1290.150 3133.930 1290.450 3134.310 ;
        RECT 1338.910 3134.310 1387.050 3134.610 ;
        RECT 1290.150 3133.630 1338.290 3133.930 ;
        RECT 1241.390 3132.950 1242.610 3133.250 ;
        RECT 1337.990 3133.250 1338.290 3133.630 ;
        RECT 1338.910 3133.250 1339.210 3134.310 ;
        RECT 1386.750 3133.930 1387.050 3134.310 ;
        RECT 1435.510 3134.310 1449.395 3134.610 ;
        RECT 1386.750 3133.630 1434.890 3133.930 ;
        RECT 1337.990 3132.950 1339.210 3133.250 ;
        RECT 1434.590 3133.250 1434.890 3133.630 ;
        RECT 1435.510 3133.250 1435.810 3134.310 ;
        RECT 1449.065 3134.295 1449.395 3134.310 ;
        RECT 1497.110 3134.610 1497.490 3134.620 ;
        RECT 2125.265 3134.610 2125.595 3134.625 ;
        RECT 1497.110 3134.310 1580.250 3134.610 ;
        RECT 1497.110 3134.300 1497.490 3134.310 ;
        RECT 1579.950 3133.930 1580.250 3134.310 ;
        RECT 1628.710 3134.310 1676.850 3134.610 ;
        RECT 1579.950 3133.630 1628.090 3133.930 ;
        RECT 1434.590 3132.950 1435.810 3133.250 ;
        RECT 1463.325 3133.250 1463.655 3133.265 ;
        RECT 1497.110 3133.250 1497.490 3133.260 ;
        RECT 1463.325 3132.950 1497.490 3133.250 ;
        RECT 1627.790 3133.250 1628.090 3133.630 ;
        RECT 1628.710 3133.250 1629.010 3134.310 ;
        RECT 1676.550 3133.930 1676.850 3134.310 ;
        RECT 1725.310 3134.310 1773.450 3134.610 ;
        RECT 1676.550 3133.630 1724.690 3133.930 ;
        RECT 1627.790 3132.950 1629.010 3133.250 ;
        RECT 1724.390 3133.250 1724.690 3133.630 ;
        RECT 1725.310 3133.250 1725.610 3134.310 ;
        RECT 1773.150 3133.930 1773.450 3134.310 ;
        RECT 1821.910 3134.310 1870.050 3134.610 ;
        RECT 1773.150 3133.630 1821.290 3133.930 ;
        RECT 1724.390 3132.950 1725.610 3133.250 ;
        RECT 1820.990 3133.250 1821.290 3133.630 ;
        RECT 1821.910 3133.250 1822.210 3134.310 ;
        RECT 1869.750 3133.930 1870.050 3134.310 ;
        RECT 1918.510 3134.310 1966.650 3134.610 ;
        RECT 1869.750 3133.630 1917.890 3133.930 ;
        RECT 1820.990 3132.950 1822.210 3133.250 ;
        RECT 1917.590 3133.250 1917.890 3133.630 ;
        RECT 1918.510 3133.250 1918.810 3134.310 ;
        RECT 1966.350 3133.930 1966.650 3134.310 ;
        RECT 2015.110 3134.310 2063.250 3134.610 ;
        RECT 1966.350 3133.630 2014.490 3133.930 ;
        RECT 1917.590 3132.950 1918.810 3133.250 ;
        RECT 2014.190 3133.250 2014.490 3133.630 ;
        RECT 2015.110 3133.250 2015.410 3134.310 ;
        RECT 2062.950 3133.930 2063.250 3134.310 ;
        RECT 2111.710 3134.310 2125.595 3134.610 ;
        RECT 2062.950 3133.630 2111.090 3133.930 ;
        RECT 2014.190 3132.950 2015.410 3133.250 ;
        RECT 2110.790 3133.250 2111.090 3133.630 ;
        RECT 2111.710 3133.250 2112.010 3134.310 ;
        RECT 2125.265 3134.295 2125.595 3134.310 ;
        RECT 2173.310 3134.610 2173.690 3134.620 ;
        RECT 2704.865 3134.610 2705.195 3134.625 ;
        RECT 2173.310 3134.310 2256.450 3134.610 ;
        RECT 2173.310 3134.300 2173.690 3134.310 ;
        RECT 2256.150 3133.930 2256.450 3134.310 ;
        RECT 2304.910 3134.310 2353.050 3134.610 ;
        RECT 2256.150 3133.630 2304.290 3133.930 ;
        RECT 2110.790 3132.950 2112.010 3133.250 ;
        RECT 2139.525 3133.250 2139.855 3133.265 ;
        RECT 2173.310 3133.250 2173.690 3133.260 ;
        RECT 2139.525 3132.950 2173.690 3133.250 ;
        RECT 2303.990 3133.250 2304.290 3133.630 ;
        RECT 2304.910 3133.250 2305.210 3134.310 ;
        RECT 2352.750 3133.930 2353.050 3134.310 ;
        RECT 2401.510 3134.310 2449.650 3134.610 ;
        RECT 2352.750 3133.630 2400.890 3133.930 ;
        RECT 2303.990 3132.950 2305.210 3133.250 ;
        RECT 2400.590 3133.250 2400.890 3133.630 ;
        RECT 2401.510 3133.250 2401.810 3134.310 ;
        RECT 2449.350 3133.930 2449.650 3134.310 ;
        RECT 2498.110 3134.310 2546.250 3134.610 ;
        RECT 2449.350 3133.630 2497.490 3133.930 ;
        RECT 2400.590 3132.950 2401.810 3133.250 ;
        RECT 2497.190 3133.250 2497.490 3133.630 ;
        RECT 2498.110 3133.250 2498.410 3134.310 ;
        RECT 2545.950 3133.930 2546.250 3134.310 ;
        RECT 2594.710 3134.310 2642.850 3134.610 ;
        RECT 2545.950 3133.630 2594.090 3133.930 ;
        RECT 2497.190 3132.950 2498.410 3133.250 ;
        RECT 2593.790 3133.250 2594.090 3133.630 ;
        RECT 2594.710 3133.250 2595.010 3134.310 ;
        RECT 2642.550 3133.930 2642.850 3134.310 ;
        RECT 2691.310 3134.310 2705.195 3134.610 ;
        RECT 2642.550 3133.630 2690.690 3133.930 ;
        RECT 2593.790 3132.950 2595.010 3133.250 ;
        RECT 2690.390 3133.250 2690.690 3133.630 ;
        RECT 2691.310 3133.250 2691.610 3134.310 ;
        RECT 2704.865 3134.295 2705.195 3134.310 ;
        RECT 2825.845 3134.610 2826.175 3134.625 ;
        RECT 2863.565 3134.610 2863.895 3134.625 ;
        RECT 2825.845 3134.310 2849.850 3134.610 ;
        RECT 2825.845 3134.295 2826.175 3134.310 ;
        RECT 2849.550 3133.930 2849.850 3134.310 ;
        RECT 2863.565 3134.310 2884.810 3134.610 ;
        RECT 2863.565 3134.295 2863.895 3134.310 ;
        RECT 2863.105 3133.930 2863.435 3133.945 ;
        RECT 2849.550 3133.630 2863.435 3133.930 ;
        RECT 2884.510 3133.930 2884.810 3134.310 ;
        RECT 2916.710 3133.930 2917.010 3138.390 ;
        RECT 2917.600 3137.940 2924.800 3138.390 ;
        RECT 2884.510 3133.630 2917.010 3133.930 ;
        RECT 2863.105 3133.615 2863.435 3133.630 ;
        RECT 2690.390 3132.950 2691.610 3133.250 ;
        RECT 2743.045 3133.250 2743.375 3133.265 ;
        RECT 2752.910 3133.250 2753.290 3133.260 ;
        RECT 2743.045 3132.950 2753.290 3133.250 ;
        RECT 1463.325 3132.935 1463.655 3132.950 ;
        RECT 1497.110 3132.940 1497.490 3132.950 ;
        RECT 2139.525 3132.935 2139.855 3132.950 ;
        RECT 2173.310 3132.940 2173.690 3132.950 ;
        RECT 2743.045 3132.935 2743.375 3132.950 ;
        RECT 2752.910 3132.940 2753.290 3132.950 ;
        RECT 290.070 1415.570 290.450 1415.580 ;
        RECT 290.070 1415.440 300.380 1415.570 ;
        RECT 290.070 1415.270 304.000 1415.440 ;
        RECT 290.070 1415.260 290.450 1415.270 ;
        RECT 300.000 1414.840 304.000 1415.270 ;
      LAYER via3 ;
        RECT 2752.940 3134.980 2753.260 3135.300 ;
        RECT 290.100 3134.300 290.420 3134.620 ;
        RECT 1497.140 3134.300 1497.460 3134.620 ;
        RECT 1497.140 3132.940 1497.460 3133.260 ;
        RECT 2173.340 3134.300 2173.660 3134.620 ;
        RECT 2173.340 3132.940 2173.660 3133.260 ;
        RECT 2752.940 3132.940 2753.260 3133.260 ;
        RECT 290.100 1415.260 290.420 1415.580 ;
      LAYER met4 ;
        RECT 2752.935 3134.975 2753.265 3135.305 ;
        RECT 290.095 3134.295 290.425 3134.625 ;
        RECT 1497.135 3134.295 1497.465 3134.625 ;
        RECT 2173.335 3134.295 2173.665 3134.625 ;
        RECT 290.110 1415.585 290.410 3134.295 ;
        RECT 1497.150 3133.265 1497.450 3134.295 ;
        RECT 2173.350 3133.265 2173.650 3134.295 ;
        RECT 2752.950 3133.265 2753.250 3134.975 ;
        RECT 1497.135 3132.935 1497.465 3133.265 ;
        RECT 2173.335 3132.935 2173.665 3133.265 ;
        RECT 2752.935 3132.935 2753.265 3133.265 ;
        RECT 290.095 1415.255 290.425 1415.585 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2801.470 3369.640 2801.790 3369.700 ;
        RECT 2825.850 3369.640 2826.170 3369.700 ;
        RECT 2801.470 3369.500 2826.170 3369.640 ;
        RECT 2801.470 3369.440 2801.790 3369.500 ;
        RECT 2825.850 3369.440 2826.170 3369.500 ;
        RECT 1449.070 3368.960 1449.390 3369.020 ;
        RECT 1463.330 3368.960 1463.650 3369.020 ;
        RECT 1449.070 3368.820 1463.650 3368.960 ;
        RECT 1449.070 3368.760 1449.390 3368.820 ;
        RECT 1463.330 3368.760 1463.650 3368.820 ;
        RECT 2704.870 3368.960 2705.190 3369.020 ;
        RECT 2743.050 3368.960 2743.370 3369.020 ;
        RECT 2704.870 3368.820 2743.370 3368.960 ;
        RECT 2704.870 3368.760 2705.190 3368.820 ;
        RECT 2743.050 3368.760 2743.370 3368.820 ;
      LAYER via ;
        RECT 2801.500 3369.440 2801.760 3369.700 ;
        RECT 2825.880 3369.440 2826.140 3369.700 ;
        RECT 1449.100 3368.760 1449.360 3369.020 ;
        RECT 1463.360 3368.760 1463.620 3369.020 ;
        RECT 2704.900 3368.760 2705.160 3369.020 ;
        RECT 2743.080 3368.760 2743.340 3369.020 ;
      LAYER met2 ;
        RECT 2766.530 3369.810 2766.810 3369.925 ;
        RECT 2767.450 3369.810 2767.730 3369.925 ;
        RECT 2766.530 3369.670 2767.730 3369.810 ;
        RECT 2766.530 3369.555 2766.810 3369.670 ;
        RECT 2767.450 3369.555 2767.730 3369.670 ;
        RECT 2801.490 3369.555 2801.770 3369.925 ;
        RECT 2801.500 3369.410 2801.760 3369.555 ;
        RECT 2825.880 3369.410 2826.140 3369.730 ;
        RECT 2825.940 3369.245 2826.080 3369.410 ;
        RECT 1449.090 3368.875 1449.370 3369.245 ;
        RECT 1449.100 3368.730 1449.360 3368.875 ;
        RECT 1463.360 3368.730 1463.620 3369.050 ;
        RECT 2704.890 3368.875 2705.170 3369.245 ;
        RECT 2704.900 3368.730 2705.160 3368.875 ;
        RECT 2743.080 3368.730 2743.340 3369.050 ;
        RECT 2825.870 3368.875 2826.150 3369.245 ;
        RECT 2863.590 3369.130 2863.870 3369.245 ;
        RECT 2863.200 3368.990 2863.870 3369.130 ;
        RECT 1463.420 3367.885 1463.560 3368.730 ;
        RECT 2743.140 3367.885 2743.280 3368.730 ;
        RECT 2863.200 3368.565 2863.340 3368.990 ;
        RECT 2863.590 3368.875 2863.870 3368.990 ;
        RECT 2863.130 3368.195 2863.410 3368.565 ;
        RECT 1463.350 3367.515 1463.630 3367.885 ;
        RECT 2743.070 3367.515 2743.350 3367.885 ;
      LAYER via2 ;
        RECT 2766.530 3369.600 2766.810 3369.880 ;
        RECT 2767.450 3369.600 2767.730 3369.880 ;
        RECT 2801.490 3369.600 2801.770 3369.880 ;
        RECT 1449.090 3368.920 1449.370 3369.200 ;
        RECT 2704.890 3368.920 2705.170 3369.200 ;
        RECT 2825.870 3368.920 2826.150 3369.200 ;
        RECT 2863.590 3368.920 2863.870 3369.200 ;
        RECT 2863.130 3368.240 2863.410 3368.520 ;
        RECT 1463.350 3367.560 1463.630 3367.840 ;
        RECT 2743.070 3367.560 2743.350 3367.840 ;
      LAYER met3 ;
        RECT 2917.600 3373.290 2924.800 3373.740 ;
        RECT 2916.710 3372.990 2924.800 3373.290 ;
        RECT 2752.910 3369.890 2753.290 3369.900 ;
        RECT 2766.505 3369.890 2766.835 3369.905 ;
        RECT 2752.910 3369.590 2766.835 3369.890 ;
        RECT 2752.910 3369.580 2753.290 3369.590 ;
        RECT 2766.505 3369.575 2766.835 3369.590 ;
        RECT 2767.425 3369.890 2767.755 3369.905 ;
        RECT 2801.465 3369.890 2801.795 3369.905 ;
        RECT 2767.425 3369.590 2801.795 3369.890 ;
        RECT 2767.425 3369.575 2767.755 3369.590 ;
        RECT 2801.465 3369.575 2801.795 3369.590 ;
        RECT 286.390 3369.210 286.770 3369.220 ;
        RECT 1449.065 3369.210 1449.395 3369.225 ;
        RECT 286.390 3368.910 324.450 3369.210 ;
        RECT 286.390 3368.900 286.770 3368.910 ;
        RECT 324.150 3368.530 324.450 3368.910 ;
        RECT 372.910 3368.910 421.050 3369.210 ;
        RECT 324.150 3368.230 372.290 3368.530 ;
        RECT 371.990 3367.850 372.290 3368.230 ;
        RECT 372.910 3367.850 373.210 3368.910 ;
        RECT 420.750 3368.530 421.050 3368.910 ;
        RECT 469.510 3368.910 517.650 3369.210 ;
        RECT 420.750 3368.230 468.890 3368.530 ;
        RECT 371.990 3367.550 373.210 3367.850 ;
        RECT 468.590 3367.850 468.890 3368.230 ;
        RECT 469.510 3367.850 469.810 3368.910 ;
        RECT 517.350 3368.530 517.650 3368.910 ;
        RECT 566.110 3368.910 614.250 3369.210 ;
        RECT 517.350 3368.230 565.490 3368.530 ;
        RECT 468.590 3367.550 469.810 3367.850 ;
        RECT 565.190 3367.850 565.490 3368.230 ;
        RECT 566.110 3367.850 566.410 3368.910 ;
        RECT 613.950 3368.530 614.250 3368.910 ;
        RECT 662.710 3368.910 710.850 3369.210 ;
        RECT 613.950 3368.230 662.090 3368.530 ;
        RECT 565.190 3367.550 566.410 3367.850 ;
        RECT 661.790 3367.850 662.090 3368.230 ;
        RECT 662.710 3367.850 663.010 3368.910 ;
        RECT 710.550 3368.530 710.850 3368.910 ;
        RECT 759.310 3368.910 807.450 3369.210 ;
        RECT 710.550 3368.230 758.690 3368.530 ;
        RECT 661.790 3367.550 663.010 3367.850 ;
        RECT 758.390 3367.850 758.690 3368.230 ;
        RECT 759.310 3367.850 759.610 3368.910 ;
        RECT 807.150 3368.530 807.450 3368.910 ;
        RECT 855.910 3368.910 904.050 3369.210 ;
        RECT 807.150 3368.230 855.290 3368.530 ;
        RECT 758.390 3367.550 759.610 3367.850 ;
        RECT 854.990 3367.850 855.290 3368.230 ;
        RECT 855.910 3367.850 856.210 3368.910 ;
        RECT 903.750 3368.530 904.050 3368.910 ;
        RECT 952.510 3368.910 1000.650 3369.210 ;
        RECT 903.750 3368.230 951.890 3368.530 ;
        RECT 854.990 3367.550 856.210 3367.850 ;
        RECT 951.590 3367.850 951.890 3368.230 ;
        RECT 952.510 3367.850 952.810 3368.910 ;
        RECT 1000.350 3368.530 1000.650 3368.910 ;
        RECT 1049.110 3368.910 1097.250 3369.210 ;
        RECT 1000.350 3368.230 1048.490 3368.530 ;
        RECT 951.590 3367.550 952.810 3367.850 ;
        RECT 1048.190 3367.850 1048.490 3368.230 ;
        RECT 1049.110 3367.850 1049.410 3368.910 ;
        RECT 1096.950 3368.530 1097.250 3368.910 ;
        RECT 1145.710 3368.910 1193.850 3369.210 ;
        RECT 1096.950 3368.230 1145.090 3368.530 ;
        RECT 1048.190 3367.550 1049.410 3367.850 ;
        RECT 1144.790 3367.850 1145.090 3368.230 ;
        RECT 1145.710 3367.850 1146.010 3368.910 ;
        RECT 1193.550 3368.530 1193.850 3368.910 ;
        RECT 1242.310 3368.910 1290.450 3369.210 ;
        RECT 1193.550 3368.230 1241.690 3368.530 ;
        RECT 1144.790 3367.550 1146.010 3367.850 ;
        RECT 1241.390 3367.850 1241.690 3368.230 ;
        RECT 1242.310 3367.850 1242.610 3368.910 ;
        RECT 1290.150 3368.530 1290.450 3368.910 ;
        RECT 1338.910 3368.910 1387.050 3369.210 ;
        RECT 1290.150 3368.230 1338.290 3368.530 ;
        RECT 1241.390 3367.550 1242.610 3367.850 ;
        RECT 1337.990 3367.850 1338.290 3368.230 ;
        RECT 1338.910 3367.850 1339.210 3368.910 ;
        RECT 1386.750 3368.530 1387.050 3368.910 ;
        RECT 1435.510 3368.910 1449.395 3369.210 ;
        RECT 1386.750 3368.230 1434.890 3368.530 ;
        RECT 1337.990 3367.550 1339.210 3367.850 ;
        RECT 1434.590 3367.850 1434.890 3368.230 ;
        RECT 1435.510 3367.850 1435.810 3368.910 ;
        RECT 1449.065 3368.895 1449.395 3368.910 ;
        RECT 1497.110 3369.210 1497.490 3369.220 ;
        RECT 2704.865 3369.210 2705.195 3369.225 ;
        RECT 1497.110 3368.910 1580.250 3369.210 ;
        RECT 1497.110 3368.900 1497.490 3368.910 ;
        RECT 1579.950 3368.530 1580.250 3368.910 ;
        RECT 1628.710 3368.910 1676.850 3369.210 ;
        RECT 1579.950 3368.230 1628.090 3368.530 ;
        RECT 1434.590 3367.550 1435.810 3367.850 ;
        RECT 1463.325 3367.850 1463.655 3367.865 ;
        RECT 1497.110 3367.850 1497.490 3367.860 ;
        RECT 1463.325 3367.550 1497.490 3367.850 ;
        RECT 1627.790 3367.850 1628.090 3368.230 ;
        RECT 1628.710 3367.850 1629.010 3368.910 ;
        RECT 1676.550 3368.530 1676.850 3368.910 ;
        RECT 1725.310 3368.910 1773.450 3369.210 ;
        RECT 1676.550 3368.230 1724.690 3368.530 ;
        RECT 1627.790 3367.550 1629.010 3367.850 ;
        RECT 1724.390 3367.850 1724.690 3368.230 ;
        RECT 1725.310 3367.850 1725.610 3368.910 ;
        RECT 1773.150 3368.530 1773.450 3368.910 ;
        RECT 1821.910 3368.910 1870.050 3369.210 ;
        RECT 1773.150 3368.230 1821.290 3368.530 ;
        RECT 1724.390 3367.550 1725.610 3367.850 ;
        RECT 1820.990 3367.850 1821.290 3368.230 ;
        RECT 1821.910 3367.850 1822.210 3368.910 ;
        RECT 1869.750 3368.530 1870.050 3368.910 ;
        RECT 1918.510 3368.910 1966.650 3369.210 ;
        RECT 1869.750 3368.230 1917.890 3368.530 ;
        RECT 1820.990 3367.550 1822.210 3367.850 ;
        RECT 1917.590 3367.850 1917.890 3368.230 ;
        RECT 1918.510 3367.850 1918.810 3368.910 ;
        RECT 1966.350 3368.530 1966.650 3368.910 ;
        RECT 2015.110 3368.910 2063.250 3369.210 ;
        RECT 1966.350 3368.230 2014.490 3368.530 ;
        RECT 1917.590 3367.550 1918.810 3367.850 ;
        RECT 2014.190 3367.850 2014.490 3368.230 ;
        RECT 2015.110 3367.850 2015.410 3368.910 ;
        RECT 2062.950 3368.530 2063.250 3368.910 ;
        RECT 2159.550 3368.910 2207.690 3369.210 ;
        RECT 2062.950 3368.230 2111.090 3368.530 ;
        RECT 2014.190 3367.550 2015.410 3367.850 ;
        RECT 2110.790 3367.850 2111.090 3368.230 ;
        RECT 2159.550 3367.850 2159.850 3368.910 ;
        RECT 2110.790 3367.550 2159.850 3367.850 ;
        RECT 2207.390 3367.850 2207.690 3368.910 ;
        RECT 2208.310 3368.910 2256.450 3369.210 ;
        RECT 2208.310 3367.850 2208.610 3368.910 ;
        RECT 2256.150 3368.530 2256.450 3368.910 ;
        RECT 2304.910 3368.910 2353.050 3369.210 ;
        RECT 2256.150 3368.230 2304.290 3368.530 ;
        RECT 2207.390 3367.550 2208.610 3367.850 ;
        RECT 2303.990 3367.850 2304.290 3368.230 ;
        RECT 2304.910 3367.850 2305.210 3368.910 ;
        RECT 2352.750 3368.530 2353.050 3368.910 ;
        RECT 2401.510 3368.910 2449.650 3369.210 ;
        RECT 2352.750 3368.230 2400.890 3368.530 ;
        RECT 2303.990 3367.550 2305.210 3367.850 ;
        RECT 2400.590 3367.850 2400.890 3368.230 ;
        RECT 2401.510 3367.850 2401.810 3368.910 ;
        RECT 2449.350 3368.530 2449.650 3368.910 ;
        RECT 2498.110 3368.910 2546.250 3369.210 ;
        RECT 2449.350 3368.230 2497.490 3368.530 ;
        RECT 2400.590 3367.550 2401.810 3367.850 ;
        RECT 2497.190 3367.850 2497.490 3368.230 ;
        RECT 2498.110 3367.850 2498.410 3368.910 ;
        RECT 2545.950 3368.530 2546.250 3368.910 ;
        RECT 2594.710 3368.910 2642.850 3369.210 ;
        RECT 2545.950 3368.230 2594.090 3368.530 ;
        RECT 2497.190 3367.550 2498.410 3367.850 ;
        RECT 2593.790 3367.850 2594.090 3368.230 ;
        RECT 2594.710 3367.850 2595.010 3368.910 ;
        RECT 2642.550 3368.530 2642.850 3368.910 ;
        RECT 2691.310 3368.910 2705.195 3369.210 ;
        RECT 2642.550 3368.230 2690.690 3368.530 ;
        RECT 2593.790 3367.550 2595.010 3367.850 ;
        RECT 2690.390 3367.850 2690.690 3368.230 ;
        RECT 2691.310 3367.850 2691.610 3368.910 ;
        RECT 2704.865 3368.895 2705.195 3368.910 ;
        RECT 2825.845 3369.210 2826.175 3369.225 ;
        RECT 2863.565 3369.210 2863.895 3369.225 ;
        RECT 2825.845 3368.910 2849.850 3369.210 ;
        RECT 2825.845 3368.895 2826.175 3368.910 ;
        RECT 2849.550 3368.530 2849.850 3368.910 ;
        RECT 2863.565 3368.910 2884.810 3369.210 ;
        RECT 2863.565 3368.895 2863.895 3368.910 ;
        RECT 2863.105 3368.530 2863.435 3368.545 ;
        RECT 2849.550 3368.230 2863.435 3368.530 ;
        RECT 2884.510 3368.530 2884.810 3368.910 ;
        RECT 2916.710 3368.530 2917.010 3372.990 ;
        RECT 2917.600 3372.540 2924.800 3372.990 ;
        RECT 2884.510 3368.230 2917.010 3368.530 ;
        RECT 2863.105 3368.215 2863.435 3368.230 ;
        RECT 2690.390 3367.550 2691.610 3367.850 ;
        RECT 2743.045 3367.850 2743.375 3367.865 ;
        RECT 2752.910 3367.850 2753.290 3367.860 ;
        RECT 2743.045 3367.550 2753.290 3367.850 ;
        RECT 1463.325 3367.535 1463.655 3367.550 ;
        RECT 1497.110 3367.540 1497.490 3367.550 ;
        RECT 2743.045 3367.535 2743.375 3367.550 ;
        RECT 2752.910 3367.540 2753.290 3367.550 ;
        RECT 286.390 1447.530 286.770 1447.540 ;
        RECT 286.390 1447.400 300.380 1447.530 ;
        RECT 286.390 1447.230 304.000 1447.400 ;
        RECT 286.390 1447.220 286.770 1447.230 ;
        RECT 300.000 1446.800 304.000 1447.230 ;
      LAYER via3 ;
        RECT 2752.940 3369.580 2753.260 3369.900 ;
        RECT 286.420 3368.900 286.740 3369.220 ;
        RECT 1497.140 3368.900 1497.460 3369.220 ;
        RECT 1497.140 3367.540 1497.460 3367.860 ;
        RECT 2752.940 3367.540 2753.260 3367.860 ;
        RECT 286.420 1447.220 286.740 1447.540 ;
      LAYER met4 ;
        RECT 2752.935 3369.575 2753.265 3369.905 ;
        RECT 286.415 3368.895 286.745 3369.225 ;
        RECT 1497.135 3368.895 1497.465 3369.225 ;
        RECT 286.430 1447.545 286.730 3368.895 ;
        RECT 1497.150 3367.865 1497.450 3368.895 ;
        RECT 2752.950 3367.865 2753.250 3369.575 ;
        RECT 1497.135 3367.535 1497.465 3367.865 ;
        RECT 2752.935 3367.535 2753.265 3367.865 ;
        RECT 286.415 1447.215 286.745 1447.545 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2795.490 3443.080 2795.810 3443.140 ;
        RECT 2798.250 3443.080 2798.570 3443.140 ;
        RECT 2795.490 3442.940 2798.570 3443.080 ;
        RECT 2795.490 3442.880 2795.810 3442.940 ;
        RECT 2798.250 3442.880 2798.570 3442.940 ;
        RECT 2795.030 3422.340 2795.350 3422.400 ;
        RECT 2795.490 3422.340 2795.810 3422.400 ;
        RECT 2795.030 3422.200 2795.810 3422.340 ;
        RECT 2795.030 3422.140 2795.350 3422.200 ;
        RECT 2795.490 3422.140 2795.810 3422.200 ;
        RECT 2795.490 3394.940 2795.810 3395.200 ;
        RECT 2795.580 3394.520 2795.720 3394.940 ;
        RECT 2795.490 3394.260 2795.810 3394.520 ;
        RECT 2795.490 3332.920 2795.810 3332.980 ;
        RECT 2796.870 3332.920 2797.190 3332.980 ;
        RECT 2795.490 3332.780 2797.190 3332.920 ;
        RECT 2795.490 3332.720 2795.810 3332.780 ;
        RECT 2796.870 3332.720 2797.190 3332.780 ;
        RECT 2795.490 3308.780 2795.810 3308.840 ;
        RECT 2796.870 3308.780 2797.190 3308.840 ;
        RECT 2795.490 3308.640 2797.190 3308.780 ;
        RECT 2795.490 3308.580 2795.810 3308.640 ;
        RECT 2796.870 3308.580 2797.190 3308.640 ;
        RECT 2795.490 3284.640 2795.810 3284.700 ;
        RECT 2795.950 3284.640 2796.270 3284.700 ;
        RECT 2795.490 3284.500 2796.270 3284.640 ;
        RECT 2795.490 3284.440 2795.810 3284.500 ;
        RECT 2795.950 3284.440 2796.270 3284.500 ;
        RECT 2795.490 3236.360 2795.810 3236.420 ;
        RECT 2795.950 3236.360 2796.270 3236.420 ;
        RECT 2795.490 3236.220 2796.270 3236.360 ;
        RECT 2795.490 3236.160 2795.810 3236.220 ;
        RECT 2795.950 3236.160 2796.270 3236.220 ;
        RECT 2795.490 3202.020 2795.810 3202.080 ;
        RECT 2795.950 3202.020 2796.270 3202.080 ;
        RECT 2795.490 3201.880 2796.270 3202.020 ;
        RECT 2795.490 3201.820 2795.810 3201.880 ;
        RECT 2795.950 3201.820 2796.270 3201.880 ;
        RECT 2795.030 3153.400 2795.350 3153.460 ;
        RECT 2795.950 3153.400 2796.270 3153.460 ;
        RECT 2795.030 3153.260 2796.270 3153.400 ;
        RECT 2795.030 3153.200 2795.350 3153.260 ;
        RECT 2795.950 3153.200 2796.270 3153.260 ;
        RECT 2795.950 3091.180 2796.270 3091.240 ;
        RECT 2796.870 3091.180 2797.190 3091.240 ;
        RECT 2795.950 3091.040 2797.190 3091.180 ;
        RECT 2795.950 3090.980 2796.270 3091.040 ;
        RECT 2796.870 3090.980 2797.190 3091.040 ;
        RECT 2795.490 3042.900 2795.810 3042.960 ;
        RECT 2797.330 3042.900 2797.650 3042.960 ;
        RECT 2795.490 3042.760 2797.650 3042.900 ;
        RECT 2795.490 3042.700 2795.810 3042.760 ;
        RECT 2797.330 3042.700 2797.650 3042.760 ;
        RECT 2795.950 2987.820 2796.270 2987.880 ;
        RECT 2796.870 2987.820 2797.190 2987.880 ;
        RECT 2795.950 2987.680 2797.190 2987.820 ;
        RECT 2795.950 2987.620 2796.270 2987.680 ;
        RECT 2796.870 2987.620 2797.190 2987.680 ;
        RECT 2795.950 2946.680 2796.270 2946.740 ;
        RECT 2796.870 2946.680 2797.190 2946.740 ;
        RECT 2795.950 2946.540 2797.190 2946.680 ;
        RECT 2795.950 2946.480 2796.270 2946.540 ;
        RECT 2796.870 2946.480 2797.190 2946.540 ;
        RECT 2796.870 2912.340 2797.190 2912.400 ;
        RECT 2796.500 2912.200 2797.190 2912.340 ;
        RECT 2796.500 2911.720 2796.640 2912.200 ;
        RECT 2796.870 2912.140 2797.190 2912.200 ;
        RECT 2796.410 2911.460 2796.730 2911.720 ;
        RECT 2795.030 2815.580 2795.350 2815.840 ;
        RECT 2795.120 2815.160 2795.260 2815.580 ;
        RECT 2795.030 2814.900 2795.350 2815.160 ;
        RECT 2794.570 2767.160 2794.890 2767.220 ;
        RECT 2794.570 2767.020 2795.260 2767.160 ;
        RECT 2794.570 2766.960 2794.890 2767.020 ;
        RECT 2795.120 2766.880 2795.260 2767.020 ;
        RECT 2795.030 2766.620 2795.350 2766.880 ;
        RECT 2794.570 2753.220 2794.890 2753.280 ;
        RECT 2795.030 2753.220 2795.350 2753.280 ;
        RECT 2794.570 2753.080 2795.350 2753.220 ;
        RECT 2794.570 2753.020 2794.890 2753.080 ;
        RECT 2795.030 2753.020 2795.350 2753.080 ;
        RECT 2794.570 2718.680 2794.890 2718.940 ;
        RECT 2794.660 2718.200 2794.800 2718.680 ;
        RECT 2795.030 2718.200 2795.350 2718.260 ;
        RECT 2794.660 2718.060 2795.350 2718.200 ;
        RECT 2795.030 2718.000 2795.350 2718.060 ;
        RECT 2795.030 2670.260 2795.350 2670.320 ;
        RECT 2795.950 2670.260 2796.270 2670.320 ;
        RECT 2795.030 2670.120 2796.270 2670.260 ;
        RECT 2795.030 2670.060 2795.350 2670.120 ;
        RECT 2795.950 2670.060 2796.270 2670.120 ;
        RECT 2795.950 2622.120 2796.270 2622.380 ;
        RECT 2796.040 2621.980 2796.180 2622.120 ;
        RECT 2796.410 2621.980 2796.730 2622.040 ;
        RECT 2796.040 2621.840 2796.730 2621.980 ;
        RECT 2796.410 2621.780 2796.730 2621.840 ;
        RECT 2795.490 2560.100 2795.810 2560.160 ;
        RECT 2796.870 2560.100 2797.190 2560.160 ;
        RECT 2795.490 2559.960 2797.190 2560.100 ;
        RECT 2795.490 2559.900 2795.810 2559.960 ;
        RECT 2796.870 2559.900 2797.190 2559.960 ;
        RECT 2795.950 2511.820 2796.270 2511.880 ;
        RECT 2796.870 2511.820 2797.190 2511.880 ;
        RECT 2795.950 2511.680 2797.190 2511.820 ;
        RECT 2795.950 2511.620 2796.270 2511.680 ;
        RECT 2796.870 2511.620 2797.190 2511.680 ;
        RECT 2795.490 2463.200 2795.810 2463.260 ;
        RECT 2795.950 2463.200 2796.270 2463.260 ;
        RECT 2795.490 2463.060 2796.270 2463.200 ;
        RECT 2795.490 2463.000 2795.810 2463.060 ;
        RECT 2795.950 2463.000 2796.270 2463.060 ;
        RECT 2795.490 2428.860 2795.810 2428.920 ;
        RECT 2795.950 2428.860 2796.270 2428.920 ;
        RECT 2795.490 2428.720 2796.270 2428.860 ;
        RECT 2795.490 2428.660 2795.810 2428.720 ;
        RECT 2795.950 2428.660 2796.270 2428.720 ;
        RECT 2795.030 2380.580 2795.350 2380.640 ;
        RECT 2795.950 2380.580 2796.270 2380.640 ;
        RECT 2795.030 2380.440 2796.270 2380.580 ;
        RECT 2795.030 2380.380 2795.350 2380.440 ;
        RECT 2795.950 2380.380 2796.270 2380.440 ;
        RECT 2795.490 2366.640 2795.810 2366.700 ;
        RECT 2795.950 2366.640 2796.270 2366.700 ;
        RECT 2795.490 2366.500 2796.270 2366.640 ;
        RECT 2795.490 2366.440 2795.810 2366.500 ;
        RECT 2795.950 2366.440 2796.270 2366.500 ;
        RECT 2795.950 2332.300 2796.270 2332.360 ;
        RECT 2795.580 2332.160 2796.270 2332.300 ;
        RECT 2795.580 2332.020 2795.720 2332.160 ;
        RECT 2795.950 2332.100 2796.270 2332.160 ;
        RECT 2795.490 2331.760 2795.810 2332.020 ;
        RECT 2795.030 2284.020 2795.350 2284.080 ;
        RECT 2795.950 2284.020 2796.270 2284.080 ;
        RECT 2795.030 2283.880 2796.270 2284.020 ;
        RECT 2795.030 2283.820 2795.350 2283.880 ;
        RECT 2795.950 2283.820 2796.270 2283.880 ;
        RECT 2795.950 2235.880 2796.270 2236.140 ;
        RECT 2796.040 2235.460 2796.180 2235.880 ;
        RECT 2795.950 2235.200 2796.270 2235.460 ;
        RECT 2795.490 2222.140 2795.810 2222.200 ;
        RECT 2795.950 2222.140 2796.270 2222.200 ;
        RECT 2795.490 2222.000 2796.270 2222.140 ;
        RECT 2795.490 2221.940 2795.810 2222.000 ;
        RECT 2795.950 2221.940 2796.270 2222.000 ;
      LAYER via ;
        RECT 2795.520 3442.880 2795.780 3443.140 ;
        RECT 2798.280 3442.880 2798.540 3443.140 ;
        RECT 2795.060 3422.140 2795.320 3422.400 ;
        RECT 2795.520 3422.140 2795.780 3422.400 ;
        RECT 2795.520 3394.940 2795.780 3395.200 ;
        RECT 2795.520 3394.260 2795.780 3394.520 ;
        RECT 2795.520 3332.720 2795.780 3332.980 ;
        RECT 2796.900 3332.720 2797.160 3332.980 ;
        RECT 2795.520 3308.580 2795.780 3308.840 ;
        RECT 2796.900 3308.580 2797.160 3308.840 ;
        RECT 2795.520 3284.440 2795.780 3284.700 ;
        RECT 2795.980 3284.440 2796.240 3284.700 ;
        RECT 2795.520 3236.160 2795.780 3236.420 ;
        RECT 2795.980 3236.160 2796.240 3236.420 ;
        RECT 2795.520 3201.820 2795.780 3202.080 ;
        RECT 2795.980 3201.820 2796.240 3202.080 ;
        RECT 2795.060 3153.200 2795.320 3153.460 ;
        RECT 2795.980 3153.200 2796.240 3153.460 ;
        RECT 2795.980 3090.980 2796.240 3091.240 ;
        RECT 2796.900 3090.980 2797.160 3091.240 ;
        RECT 2795.520 3042.700 2795.780 3042.960 ;
        RECT 2797.360 3042.700 2797.620 3042.960 ;
        RECT 2795.980 2987.620 2796.240 2987.880 ;
        RECT 2796.900 2987.620 2797.160 2987.880 ;
        RECT 2795.980 2946.480 2796.240 2946.740 ;
        RECT 2796.900 2946.480 2797.160 2946.740 ;
        RECT 2796.900 2912.140 2797.160 2912.400 ;
        RECT 2796.440 2911.460 2796.700 2911.720 ;
        RECT 2795.060 2815.580 2795.320 2815.840 ;
        RECT 2795.060 2814.900 2795.320 2815.160 ;
        RECT 2794.600 2766.960 2794.860 2767.220 ;
        RECT 2795.060 2766.620 2795.320 2766.880 ;
        RECT 2794.600 2753.020 2794.860 2753.280 ;
        RECT 2795.060 2753.020 2795.320 2753.280 ;
        RECT 2794.600 2718.680 2794.860 2718.940 ;
        RECT 2795.060 2718.000 2795.320 2718.260 ;
        RECT 2795.060 2670.060 2795.320 2670.320 ;
        RECT 2795.980 2670.060 2796.240 2670.320 ;
        RECT 2795.980 2622.120 2796.240 2622.380 ;
        RECT 2796.440 2621.780 2796.700 2622.040 ;
        RECT 2795.520 2559.900 2795.780 2560.160 ;
        RECT 2796.900 2559.900 2797.160 2560.160 ;
        RECT 2795.980 2511.620 2796.240 2511.880 ;
        RECT 2796.900 2511.620 2797.160 2511.880 ;
        RECT 2795.520 2463.000 2795.780 2463.260 ;
        RECT 2795.980 2463.000 2796.240 2463.260 ;
        RECT 2795.520 2428.660 2795.780 2428.920 ;
        RECT 2795.980 2428.660 2796.240 2428.920 ;
        RECT 2795.060 2380.380 2795.320 2380.640 ;
        RECT 2795.980 2380.380 2796.240 2380.640 ;
        RECT 2795.520 2366.440 2795.780 2366.700 ;
        RECT 2795.980 2366.440 2796.240 2366.700 ;
        RECT 2795.980 2332.100 2796.240 2332.360 ;
        RECT 2795.520 2331.760 2795.780 2332.020 ;
        RECT 2795.060 2283.820 2795.320 2284.080 ;
        RECT 2795.980 2283.820 2796.240 2284.080 ;
        RECT 2795.980 2235.880 2796.240 2236.140 ;
        RECT 2795.980 2235.200 2796.240 2235.460 ;
        RECT 2795.520 2221.940 2795.780 2222.200 ;
        RECT 2795.980 2221.940 2796.240 2222.200 ;
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
        RECT 2798.340 3443.170 2798.480 3517.600 ;
        RECT 2795.520 3442.850 2795.780 3443.170 ;
        RECT 2798.280 3442.850 2798.540 3443.170 ;
        RECT 2795.580 3429.650 2795.720 3442.850 ;
        RECT 2795.120 3429.510 2795.720 3429.650 ;
        RECT 2795.120 3422.430 2795.260 3429.510 ;
        RECT 2795.060 3422.110 2795.320 3422.430 ;
        RECT 2795.520 3422.110 2795.780 3422.430 ;
        RECT 2795.580 3395.230 2795.720 3422.110 ;
        RECT 2795.520 3394.910 2795.780 3395.230 ;
        RECT 2795.520 3394.230 2795.780 3394.550 ;
        RECT 2795.580 3333.010 2795.720 3394.230 ;
        RECT 2795.520 3332.690 2795.780 3333.010 ;
        RECT 2796.900 3332.690 2797.160 3333.010 ;
        RECT 2796.960 3308.870 2797.100 3332.690 ;
        RECT 2795.520 3308.550 2795.780 3308.870 ;
        RECT 2796.900 3308.550 2797.160 3308.870 ;
        RECT 2795.580 3284.730 2795.720 3308.550 ;
        RECT 2795.520 3284.410 2795.780 3284.730 ;
        RECT 2795.980 3284.410 2796.240 3284.730 ;
        RECT 2796.040 3236.450 2796.180 3284.410 ;
        RECT 2795.520 3236.130 2795.780 3236.450 ;
        RECT 2795.980 3236.130 2796.240 3236.450 ;
        RECT 2795.580 3202.110 2795.720 3236.130 ;
        RECT 2795.520 3201.790 2795.780 3202.110 ;
        RECT 2795.980 3201.790 2796.240 3202.110 ;
        RECT 2796.040 3153.490 2796.180 3201.790 ;
        RECT 2795.060 3153.170 2795.320 3153.490 ;
        RECT 2795.980 3153.170 2796.240 3153.490 ;
        RECT 2795.120 3152.890 2795.260 3153.170 ;
        RECT 2795.120 3152.750 2795.720 3152.890 ;
        RECT 2795.580 3105.290 2795.720 3152.750 ;
        RECT 2795.580 3105.150 2796.180 3105.290 ;
        RECT 2796.040 3091.270 2796.180 3105.150 ;
        RECT 2795.980 3090.950 2796.240 3091.270 ;
        RECT 2796.900 3090.950 2797.160 3091.270 ;
        RECT 2796.960 3043.525 2797.100 3090.950 ;
        RECT 2795.510 3043.155 2795.790 3043.525 ;
        RECT 2796.890 3043.155 2797.170 3043.525 ;
        RECT 2795.580 3042.990 2795.720 3043.155 ;
        RECT 2795.520 3042.670 2795.780 3042.990 ;
        RECT 2797.360 3042.670 2797.620 3042.990 ;
        RECT 2797.420 3035.930 2797.560 3042.670 ;
        RECT 2796.960 3035.790 2797.560 3035.930 ;
        RECT 2796.960 2987.910 2797.100 3035.790 ;
        RECT 2795.980 2987.590 2796.240 2987.910 ;
        RECT 2796.900 2987.590 2797.160 2987.910 ;
        RECT 2796.040 2946.770 2796.180 2987.590 ;
        RECT 2795.980 2946.450 2796.240 2946.770 ;
        RECT 2796.900 2946.450 2797.160 2946.770 ;
        RECT 2796.960 2912.430 2797.100 2946.450 ;
        RECT 2796.900 2912.110 2797.160 2912.430 ;
        RECT 2796.440 2911.430 2796.700 2911.750 ;
        RECT 2796.500 2863.210 2796.640 2911.430 ;
        RECT 2795.580 2863.070 2796.640 2863.210 ;
        RECT 2795.580 2849.610 2795.720 2863.070 ;
        RECT 2795.120 2849.470 2795.720 2849.610 ;
        RECT 2795.120 2815.870 2795.260 2849.470 ;
        RECT 2795.060 2815.550 2795.320 2815.870 ;
        RECT 2795.060 2814.870 2795.320 2815.190 ;
        RECT 2795.120 2801.330 2795.260 2814.870 ;
        RECT 2794.660 2801.190 2795.260 2801.330 ;
        RECT 2794.660 2767.250 2794.800 2801.190 ;
        RECT 2794.600 2766.930 2794.860 2767.250 ;
        RECT 2795.060 2766.590 2795.320 2766.910 ;
        RECT 2795.120 2753.310 2795.260 2766.590 ;
        RECT 2794.600 2752.990 2794.860 2753.310 ;
        RECT 2795.060 2752.990 2795.320 2753.310 ;
        RECT 2794.660 2718.970 2794.800 2752.990 ;
        RECT 2794.600 2718.650 2794.860 2718.970 ;
        RECT 2795.060 2717.970 2795.320 2718.290 ;
        RECT 2795.120 2670.350 2795.260 2717.970 ;
        RECT 2795.060 2670.030 2795.320 2670.350 ;
        RECT 2795.980 2670.030 2796.240 2670.350 ;
        RECT 2796.040 2622.410 2796.180 2670.030 ;
        RECT 2795.980 2622.090 2796.240 2622.410 ;
        RECT 2796.440 2621.750 2796.700 2622.070 ;
        RECT 2796.500 2608.325 2796.640 2621.750 ;
        RECT 2795.510 2607.955 2795.790 2608.325 ;
        RECT 2796.430 2607.955 2796.710 2608.325 ;
        RECT 2795.580 2560.190 2795.720 2607.955 ;
        RECT 2795.520 2559.870 2795.780 2560.190 ;
        RECT 2796.900 2559.870 2797.160 2560.190 ;
        RECT 2796.960 2511.910 2797.100 2559.870 ;
        RECT 2795.980 2511.590 2796.240 2511.910 ;
        RECT 2796.900 2511.590 2797.160 2511.910 ;
        RECT 2796.040 2464.165 2796.180 2511.590 ;
        RECT 2795.970 2463.795 2796.250 2464.165 ;
        RECT 2795.510 2463.115 2795.790 2463.485 ;
        RECT 2795.520 2462.970 2795.780 2463.115 ;
        RECT 2795.980 2462.970 2796.240 2463.290 ;
        RECT 2796.040 2428.950 2796.180 2462.970 ;
        RECT 2795.520 2428.630 2795.780 2428.950 ;
        RECT 2795.980 2428.630 2796.240 2428.950 ;
        RECT 2795.580 2415.090 2795.720 2428.630 ;
        RECT 2795.580 2414.950 2796.180 2415.090 ;
        RECT 2796.040 2380.670 2796.180 2414.950 ;
        RECT 2795.060 2380.410 2795.320 2380.670 ;
        RECT 2795.060 2380.350 2795.720 2380.410 ;
        RECT 2795.980 2380.350 2796.240 2380.670 ;
        RECT 2795.120 2380.270 2795.720 2380.350 ;
        RECT 2795.580 2366.730 2795.720 2380.270 ;
        RECT 2795.520 2366.410 2795.780 2366.730 ;
        RECT 2795.980 2366.410 2796.240 2366.730 ;
        RECT 2796.040 2332.390 2796.180 2366.410 ;
        RECT 2795.980 2332.070 2796.240 2332.390 ;
        RECT 2795.520 2331.730 2795.780 2332.050 ;
        RECT 2795.580 2318.530 2795.720 2331.730 ;
        RECT 2795.580 2318.390 2796.180 2318.530 ;
        RECT 2796.040 2284.110 2796.180 2318.390 ;
        RECT 2795.060 2283.850 2795.320 2284.110 ;
        RECT 2795.980 2283.850 2796.240 2284.110 ;
        RECT 2795.060 2283.790 2796.240 2283.850 ;
        RECT 2795.120 2283.710 2796.180 2283.790 ;
        RECT 2796.040 2236.170 2796.180 2283.710 ;
        RECT 2795.980 2235.850 2796.240 2236.170 ;
        RECT 2795.980 2235.170 2796.240 2235.490 ;
        RECT 2796.040 2222.230 2796.180 2235.170 ;
        RECT 2795.520 2221.910 2795.780 2222.230 ;
        RECT 2795.980 2221.910 2796.240 2222.230 ;
        RECT 2795.580 2198.285 2795.720 2221.910 ;
        RECT 2795.510 2197.915 2795.790 2198.285 ;
      LAYER via2 ;
        RECT 2795.510 3043.200 2795.790 3043.480 ;
        RECT 2796.890 3043.200 2797.170 3043.480 ;
        RECT 2795.510 2608.000 2795.790 2608.280 ;
        RECT 2796.430 2608.000 2796.710 2608.280 ;
        RECT 2795.970 2463.840 2796.250 2464.120 ;
        RECT 2795.510 2463.160 2795.790 2463.440 ;
        RECT 2795.510 2197.960 2795.790 2198.240 ;
      LAYER met3 ;
        RECT 2795.485 3043.490 2795.815 3043.505 ;
        RECT 2796.865 3043.490 2797.195 3043.505 ;
        RECT 2795.485 3043.190 2797.195 3043.490 ;
        RECT 2795.485 3043.175 2795.815 3043.190 ;
        RECT 2796.865 3043.175 2797.195 3043.190 ;
        RECT 2795.485 2608.290 2795.815 2608.305 ;
        RECT 2796.405 2608.290 2796.735 2608.305 ;
        RECT 2795.485 2607.990 2796.735 2608.290 ;
        RECT 2795.485 2607.975 2795.815 2607.990 ;
        RECT 2796.405 2607.975 2796.735 2607.990 ;
        RECT 2795.945 2464.130 2796.275 2464.145 ;
        RECT 2795.270 2463.830 2796.275 2464.130 ;
        RECT 2795.270 2463.465 2795.570 2463.830 ;
        RECT 2795.945 2463.815 2796.275 2463.830 ;
        RECT 2795.270 2463.150 2795.815 2463.465 ;
        RECT 2795.485 2463.135 2795.815 2463.150 ;
        RECT 284.550 2198.250 284.930 2198.260 ;
        RECT 2795.485 2198.250 2795.815 2198.265 ;
        RECT 284.550 2197.950 2795.815 2198.250 ;
        RECT 284.550 2197.940 284.930 2197.950 ;
        RECT 2795.485 2197.935 2795.815 2197.950 ;
        RECT 284.550 1478.810 284.930 1478.820 ;
        RECT 284.550 1478.680 300.380 1478.810 ;
        RECT 284.550 1478.510 304.000 1478.680 ;
        RECT 284.550 1478.500 284.930 1478.510 ;
        RECT 300.000 1478.080 304.000 1478.510 ;
      LAYER via3 ;
        RECT 284.580 2197.940 284.900 2198.260 ;
        RECT 284.580 1478.500 284.900 1478.820 ;
      LAYER met4 ;
        RECT 284.575 2197.935 284.905 2198.265 ;
        RECT 284.590 1478.825 284.890 2197.935 ;
        RECT 284.575 1478.495 284.905 1478.825 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
        RECT 2474.040 3503.205 2474.180 3517.600 ;
        RECT 2473.970 3502.835 2474.250 3503.205 ;
      LAYER via2 ;
        RECT 2473.970 3502.880 2474.250 3503.160 ;
      LAYER met3 ;
        RECT 288.230 3503.170 288.610 3503.180 ;
        RECT 2473.945 3503.170 2474.275 3503.185 ;
        RECT 288.230 3502.870 2474.275 3503.170 ;
        RECT 288.230 3502.860 288.610 3502.870 ;
        RECT 2473.945 3502.855 2474.275 3502.870 ;
        RECT 288.230 1510.770 288.610 1510.780 ;
        RECT 288.230 1510.640 300.380 1510.770 ;
        RECT 288.230 1510.470 304.000 1510.640 ;
        RECT 288.230 1510.460 288.610 1510.470 ;
        RECT 300.000 1510.040 304.000 1510.470 ;
      LAYER via3 ;
        RECT 288.260 3502.860 288.580 3503.180 ;
        RECT 288.260 1510.460 288.580 1510.780 ;
      LAYER met4 ;
        RECT 288.255 3502.855 288.585 3503.185 ;
        RECT 288.270 1510.785 288.570 3502.855 ;
        RECT 288.255 1510.455 288.585 1510.785 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2145.970 3464.160 2146.290 3464.220 ;
        RECT 2149.650 3464.160 2149.970 3464.220 ;
        RECT 2145.970 3464.020 2149.970 3464.160 ;
        RECT 2145.970 3463.960 2146.290 3464.020 ;
        RECT 2149.650 3463.960 2149.970 3464.020 ;
        RECT 2145.970 3367.260 2146.290 3367.320 ;
        RECT 2147.350 3367.260 2147.670 3367.320 ;
        RECT 2145.970 3367.120 2147.670 3367.260 ;
        RECT 2145.970 3367.060 2146.290 3367.120 ;
        RECT 2147.350 3367.060 2147.670 3367.120 ;
        RECT 2146.890 3236.360 2147.210 3236.420 ;
        RECT 2147.350 3236.360 2147.670 3236.420 ;
        RECT 2146.890 3236.220 2147.670 3236.360 ;
        RECT 2146.890 3236.160 2147.210 3236.220 ;
        RECT 2147.350 3236.160 2147.670 3236.220 ;
        RECT 2146.890 3202.020 2147.210 3202.080 ;
        RECT 2147.350 3202.020 2147.670 3202.080 ;
        RECT 2146.890 3201.880 2147.670 3202.020 ;
        RECT 2146.890 3201.820 2147.210 3201.880 ;
        RECT 2147.350 3201.820 2147.670 3201.880 ;
        RECT 2146.430 3153.400 2146.750 3153.460 ;
        RECT 2147.350 3153.400 2147.670 3153.460 ;
        RECT 2146.430 3153.260 2147.670 3153.400 ;
        RECT 2146.430 3153.200 2146.750 3153.260 ;
        RECT 2147.350 3153.200 2147.670 3153.260 ;
        RECT 2147.350 3091.180 2147.670 3091.240 ;
        RECT 2148.270 3091.180 2148.590 3091.240 ;
        RECT 2147.350 3091.040 2148.590 3091.180 ;
        RECT 2147.350 3090.980 2147.670 3091.040 ;
        RECT 2148.270 3090.980 2148.590 3091.040 ;
        RECT 2146.430 3043.240 2146.750 3043.300 ;
        RECT 2148.270 3043.240 2148.590 3043.300 ;
        RECT 2146.430 3043.100 2148.590 3043.240 ;
        RECT 2146.430 3043.040 2146.750 3043.100 ;
        RECT 2148.270 3043.040 2148.590 3043.100 ;
        RECT 2145.970 3042.560 2146.290 3042.620 ;
        RECT 2146.430 3042.560 2146.750 3042.620 ;
        RECT 2145.970 3042.420 2146.750 3042.560 ;
        RECT 2145.970 3042.360 2146.290 3042.420 ;
        RECT 2146.430 3042.360 2146.750 3042.420 ;
        RECT 2145.970 2994.960 2146.290 2995.020 ;
        RECT 2146.890 2994.960 2147.210 2995.020 ;
        RECT 2145.970 2994.820 2147.210 2994.960 ;
        RECT 2145.970 2994.760 2146.290 2994.820 ;
        RECT 2146.890 2994.760 2147.210 2994.820 ;
        RECT 2145.970 2994.280 2146.290 2994.340 ;
        RECT 2146.890 2994.280 2147.210 2994.340 ;
        RECT 2145.970 2994.140 2147.210 2994.280 ;
        RECT 2145.970 2994.080 2146.290 2994.140 ;
        RECT 2146.890 2994.080 2147.210 2994.140 ;
        RECT 2145.970 2946.680 2146.290 2946.740 ;
        RECT 2147.350 2946.680 2147.670 2946.740 ;
        RECT 2145.970 2946.540 2147.670 2946.680 ;
        RECT 2145.970 2946.480 2146.290 2946.540 ;
        RECT 2147.350 2946.480 2147.670 2946.540 ;
        RECT 2146.890 2898.060 2147.210 2898.120 ;
        RECT 2147.810 2898.060 2148.130 2898.120 ;
        RECT 2146.890 2897.920 2148.130 2898.060 ;
        RECT 2146.890 2897.860 2147.210 2897.920 ;
        RECT 2147.810 2897.860 2148.130 2897.920 ;
        RECT 2146.890 2849.780 2147.210 2849.840 ;
        RECT 2148.270 2849.780 2148.590 2849.840 ;
        RECT 2146.890 2849.640 2148.590 2849.780 ;
        RECT 2146.890 2849.580 2147.210 2849.640 ;
        RECT 2148.270 2849.580 2148.590 2849.640 ;
        RECT 2147.350 2818.840 2147.670 2818.900 ;
        RECT 2148.270 2818.840 2148.590 2818.900 ;
        RECT 2147.350 2818.700 2148.590 2818.840 ;
        RECT 2147.350 2818.640 2147.670 2818.700 ;
        RECT 2148.270 2818.640 2148.590 2818.700 ;
        RECT 2146.430 2801.160 2146.750 2801.220 ;
        RECT 2147.350 2801.160 2147.670 2801.220 ;
        RECT 2146.430 2801.020 2147.670 2801.160 ;
        RECT 2146.430 2800.960 2146.750 2801.020 ;
        RECT 2147.350 2800.960 2147.670 2801.020 ;
        RECT 2146.430 2753.220 2146.750 2753.280 ;
        RECT 2147.810 2753.220 2148.130 2753.280 ;
        RECT 2146.430 2753.080 2148.130 2753.220 ;
        RECT 2146.430 2753.020 2146.750 2753.080 ;
        RECT 2147.810 2753.020 2148.130 2753.080 ;
        RECT 2145.970 2656.660 2146.290 2656.720 ;
        RECT 2147.350 2656.660 2147.670 2656.720 ;
        RECT 2145.970 2656.520 2147.670 2656.660 ;
        RECT 2145.970 2656.460 2146.290 2656.520 ;
        RECT 2147.350 2656.460 2147.670 2656.520 ;
        RECT 2147.350 2622.120 2147.670 2622.380 ;
        RECT 2147.440 2621.980 2147.580 2622.120 ;
        RECT 2147.810 2621.980 2148.130 2622.040 ;
        RECT 2147.440 2621.840 2148.130 2621.980 ;
        RECT 2147.810 2621.780 2148.130 2621.840 ;
        RECT 2146.890 2560.100 2147.210 2560.160 ;
        RECT 2148.270 2560.100 2148.590 2560.160 ;
        RECT 2146.890 2559.960 2148.590 2560.100 ;
        RECT 2146.890 2559.900 2147.210 2559.960 ;
        RECT 2148.270 2559.900 2148.590 2559.960 ;
        RECT 2147.350 2511.820 2147.670 2511.880 ;
        RECT 2148.270 2511.820 2148.590 2511.880 ;
        RECT 2147.350 2511.680 2148.590 2511.820 ;
        RECT 2147.350 2511.620 2147.670 2511.680 ;
        RECT 2148.270 2511.620 2148.590 2511.680 ;
        RECT 2147.350 2429.000 2147.670 2429.260 ;
        RECT 2147.440 2428.860 2147.580 2429.000 ;
        RECT 2147.810 2428.860 2148.130 2428.920 ;
        RECT 2147.440 2428.720 2148.130 2428.860 ;
        RECT 2147.810 2428.660 2148.130 2428.720 ;
        RECT 2147.810 2414.920 2148.130 2414.980 ;
        RECT 2148.270 2414.920 2148.590 2414.980 ;
        RECT 2147.810 2414.780 2148.590 2414.920 ;
        RECT 2147.810 2414.720 2148.130 2414.780 ;
        RECT 2148.270 2414.720 2148.590 2414.780 ;
        RECT 2148.270 2380.580 2148.590 2380.640 ;
        RECT 2147.900 2380.440 2148.590 2380.580 ;
        RECT 2147.900 2380.300 2148.040 2380.440 ;
        RECT 2148.270 2380.380 2148.590 2380.440 ;
        RECT 2147.810 2380.040 2148.130 2380.300 ;
        RECT 2147.350 2235.880 2147.670 2236.140 ;
        RECT 2147.440 2235.460 2147.580 2235.880 ;
        RECT 2147.350 2235.200 2147.670 2235.460 ;
        RECT 2146.890 2222.140 2147.210 2222.200 ;
        RECT 2147.350 2222.140 2147.670 2222.200 ;
        RECT 2146.890 2222.000 2147.670 2222.140 ;
        RECT 2146.890 2221.940 2147.210 2222.000 ;
        RECT 2147.350 2221.940 2147.670 2222.000 ;
        RECT 285.270 2198.340 285.590 2198.400 ;
        RECT 2146.890 2198.340 2147.210 2198.400 ;
        RECT 285.270 2198.200 2147.210 2198.340 ;
        RECT 285.270 2198.140 285.590 2198.200 ;
        RECT 2146.890 2198.140 2147.210 2198.200 ;
      LAYER via ;
        RECT 2146.000 3463.960 2146.260 3464.220 ;
        RECT 2149.680 3463.960 2149.940 3464.220 ;
        RECT 2146.000 3367.060 2146.260 3367.320 ;
        RECT 2147.380 3367.060 2147.640 3367.320 ;
        RECT 2146.920 3236.160 2147.180 3236.420 ;
        RECT 2147.380 3236.160 2147.640 3236.420 ;
        RECT 2146.920 3201.820 2147.180 3202.080 ;
        RECT 2147.380 3201.820 2147.640 3202.080 ;
        RECT 2146.460 3153.200 2146.720 3153.460 ;
        RECT 2147.380 3153.200 2147.640 3153.460 ;
        RECT 2147.380 3090.980 2147.640 3091.240 ;
        RECT 2148.300 3090.980 2148.560 3091.240 ;
        RECT 2146.460 3043.040 2146.720 3043.300 ;
        RECT 2148.300 3043.040 2148.560 3043.300 ;
        RECT 2146.000 3042.360 2146.260 3042.620 ;
        RECT 2146.460 3042.360 2146.720 3042.620 ;
        RECT 2146.000 2994.760 2146.260 2995.020 ;
        RECT 2146.920 2994.760 2147.180 2995.020 ;
        RECT 2146.000 2994.080 2146.260 2994.340 ;
        RECT 2146.920 2994.080 2147.180 2994.340 ;
        RECT 2146.000 2946.480 2146.260 2946.740 ;
        RECT 2147.380 2946.480 2147.640 2946.740 ;
        RECT 2146.920 2897.860 2147.180 2898.120 ;
        RECT 2147.840 2897.860 2148.100 2898.120 ;
        RECT 2146.920 2849.580 2147.180 2849.840 ;
        RECT 2148.300 2849.580 2148.560 2849.840 ;
        RECT 2147.380 2818.640 2147.640 2818.900 ;
        RECT 2148.300 2818.640 2148.560 2818.900 ;
        RECT 2146.460 2800.960 2146.720 2801.220 ;
        RECT 2147.380 2800.960 2147.640 2801.220 ;
        RECT 2146.460 2753.020 2146.720 2753.280 ;
        RECT 2147.840 2753.020 2148.100 2753.280 ;
        RECT 2146.000 2656.460 2146.260 2656.720 ;
        RECT 2147.380 2656.460 2147.640 2656.720 ;
        RECT 2147.380 2622.120 2147.640 2622.380 ;
        RECT 2147.840 2621.780 2148.100 2622.040 ;
        RECT 2146.920 2559.900 2147.180 2560.160 ;
        RECT 2148.300 2559.900 2148.560 2560.160 ;
        RECT 2147.380 2511.620 2147.640 2511.880 ;
        RECT 2148.300 2511.620 2148.560 2511.880 ;
        RECT 2147.380 2429.000 2147.640 2429.260 ;
        RECT 2147.840 2428.660 2148.100 2428.920 ;
        RECT 2147.840 2414.720 2148.100 2414.980 ;
        RECT 2148.300 2414.720 2148.560 2414.980 ;
        RECT 2148.300 2380.380 2148.560 2380.640 ;
        RECT 2147.840 2380.040 2148.100 2380.300 ;
        RECT 2147.380 2235.880 2147.640 2236.140 ;
        RECT 2147.380 2235.200 2147.640 2235.460 ;
        RECT 2146.920 2221.940 2147.180 2222.200 ;
        RECT 2147.380 2221.940 2147.640 2222.200 ;
        RECT 285.300 2198.140 285.560 2198.400 ;
        RECT 2146.920 2198.140 2147.180 2198.400 ;
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
        RECT 2149.280 3517.370 2149.420 3517.600 ;
        RECT 2149.280 3517.230 2149.880 3517.370 ;
        RECT 2149.740 3464.250 2149.880 3517.230 ;
        RECT 2146.000 3463.930 2146.260 3464.250 ;
        RECT 2149.680 3463.930 2149.940 3464.250 ;
        RECT 2146.060 3367.350 2146.200 3463.930 ;
        RECT 2146.000 3367.030 2146.260 3367.350 ;
        RECT 2147.380 3367.030 2147.640 3367.350 ;
        RECT 2147.440 3236.450 2147.580 3367.030 ;
        RECT 2146.920 3236.130 2147.180 3236.450 ;
        RECT 2147.380 3236.130 2147.640 3236.450 ;
        RECT 2146.980 3202.110 2147.120 3236.130 ;
        RECT 2146.920 3201.790 2147.180 3202.110 ;
        RECT 2147.380 3201.790 2147.640 3202.110 ;
        RECT 2147.440 3153.490 2147.580 3201.790 ;
        RECT 2146.460 3153.170 2146.720 3153.490 ;
        RECT 2147.380 3153.170 2147.640 3153.490 ;
        RECT 2146.520 3152.890 2146.660 3153.170 ;
        RECT 2146.520 3152.750 2147.120 3152.890 ;
        RECT 2146.980 3105.290 2147.120 3152.750 ;
        RECT 2146.980 3105.150 2147.580 3105.290 ;
        RECT 2147.440 3091.270 2147.580 3105.150 ;
        RECT 2147.380 3090.950 2147.640 3091.270 ;
        RECT 2148.300 3090.950 2148.560 3091.270 ;
        RECT 2148.360 3043.330 2148.500 3090.950 ;
        RECT 2146.460 3043.010 2146.720 3043.330 ;
        RECT 2148.300 3043.010 2148.560 3043.330 ;
        RECT 2146.520 3042.650 2146.660 3043.010 ;
        RECT 2146.000 3042.330 2146.260 3042.650 ;
        RECT 2146.460 3042.330 2146.720 3042.650 ;
        RECT 2146.060 2995.050 2146.200 3042.330 ;
        RECT 2146.000 2994.730 2146.260 2995.050 ;
        RECT 2146.920 2994.730 2147.180 2995.050 ;
        RECT 2146.980 2994.370 2147.120 2994.730 ;
        RECT 2146.000 2994.050 2146.260 2994.370 ;
        RECT 2146.920 2994.050 2147.180 2994.370 ;
        RECT 2146.060 2946.770 2146.200 2994.050 ;
        RECT 2146.000 2946.450 2146.260 2946.770 ;
        RECT 2147.380 2946.450 2147.640 2946.770 ;
        RECT 2147.440 2912.170 2147.580 2946.450 ;
        RECT 2147.440 2912.030 2148.040 2912.170 ;
        RECT 2147.900 2898.150 2148.040 2912.030 ;
        RECT 2146.920 2897.830 2147.180 2898.150 ;
        RECT 2147.840 2897.830 2148.100 2898.150 ;
        RECT 2146.980 2849.870 2147.120 2897.830 ;
        RECT 2146.920 2849.550 2147.180 2849.870 ;
        RECT 2148.300 2849.550 2148.560 2849.870 ;
        RECT 2148.360 2818.930 2148.500 2849.550 ;
        RECT 2147.380 2818.610 2147.640 2818.930 ;
        RECT 2148.300 2818.610 2148.560 2818.930 ;
        RECT 2147.440 2801.250 2147.580 2818.610 ;
        RECT 2146.460 2800.930 2146.720 2801.250 ;
        RECT 2147.380 2800.930 2147.640 2801.250 ;
        RECT 2146.520 2753.310 2146.660 2800.930 ;
        RECT 2146.460 2752.990 2146.720 2753.310 ;
        RECT 2147.840 2752.990 2148.100 2753.310 ;
        RECT 2147.900 2719.165 2148.040 2752.990 ;
        RECT 2147.830 2718.795 2148.110 2719.165 ;
        RECT 2146.910 2718.115 2147.190 2718.485 ;
        RECT 2146.980 2704.885 2147.120 2718.115 ;
        RECT 2145.990 2704.515 2146.270 2704.885 ;
        RECT 2146.910 2704.515 2147.190 2704.885 ;
        RECT 2146.060 2656.750 2146.200 2704.515 ;
        RECT 2146.000 2656.430 2146.260 2656.750 ;
        RECT 2147.380 2656.430 2147.640 2656.750 ;
        RECT 2147.440 2622.410 2147.580 2656.430 ;
        RECT 2147.380 2622.090 2147.640 2622.410 ;
        RECT 2147.840 2621.750 2148.100 2622.070 ;
        RECT 2147.900 2608.325 2148.040 2621.750 ;
        RECT 2146.910 2607.955 2147.190 2608.325 ;
        RECT 2147.830 2607.955 2148.110 2608.325 ;
        RECT 2146.980 2560.190 2147.120 2607.955 ;
        RECT 2146.920 2559.870 2147.180 2560.190 ;
        RECT 2148.300 2559.870 2148.560 2560.190 ;
        RECT 2148.360 2511.910 2148.500 2559.870 ;
        RECT 2147.380 2511.590 2147.640 2511.910 ;
        RECT 2148.300 2511.590 2148.560 2511.910 ;
        RECT 2147.440 2429.290 2147.580 2511.590 ;
        RECT 2147.380 2428.970 2147.640 2429.290 ;
        RECT 2147.840 2428.630 2148.100 2428.950 ;
        RECT 2147.900 2415.010 2148.040 2428.630 ;
        RECT 2147.840 2414.690 2148.100 2415.010 ;
        RECT 2148.300 2414.690 2148.560 2415.010 ;
        RECT 2148.360 2380.670 2148.500 2414.690 ;
        RECT 2148.300 2380.350 2148.560 2380.670 ;
        RECT 2147.840 2380.010 2148.100 2380.330 ;
        RECT 2147.900 2366.810 2148.040 2380.010 ;
        RECT 2147.900 2366.670 2148.500 2366.810 ;
        RECT 2148.360 2318.645 2148.500 2366.670 ;
        RECT 2147.370 2318.275 2147.650 2318.645 ;
        RECT 2148.290 2318.275 2148.570 2318.645 ;
        RECT 2147.440 2236.170 2147.580 2318.275 ;
        RECT 2147.380 2235.850 2147.640 2236.170 ;
        RECT 2147.380 2235.170 2147.640 2235.490 ;
        RECT 2147.440 2222.230 2147.580 2235.170 ;
        RECT 2146.920 2221.910 2147.180 2222.230 ;
        RECT 2147.380 2221.910 2147.640 2222.230 ;
        RECT 2146.980 2198.430 2147.120 2221.910 ;
        RECT 285.300 2198.110 285.560 2198.430 ;
        RECT 2146.920 2198.110 2147.180 2198.430 ;
        RECT 285.360 1542.085 285.500 2198.110 ;
        RECT 285.290 1541.715 285.570 1542.085 ;
      LAYER via2 ;
        RECT 2147.830 2718.840 2148.110 2719.120 ;
        RECT 2146.910 2718.160 2147.190 2718.440 ;
        RECT 2145.990 2704.560 2146.270 2704.840 ;
        RECT 2146.910 2704.560 2147.190 2704.840 ;
        RECT 2146.910 2608.000 2147.190 2608.280 ;
        RECT 2147.830 2608.000 2148.110 2608.280 ;
        RECT 2147.370 2318.320 2147.650 2318.600 ;
        RECT 2148.290 2318.320 2148.570 2318.600 ;
        RECT 285.290 1541.760 285.570 1542.040 ;
      LAYER met3 ;
        RECT 2147.805 2719.130 2148.135 2719.145 ;
        RECT 2147.590 2718.815 2148.135 2719.130 ;
        RECT 2146.885 2718.450 2147.215 2718.465 ;
        RECT 2147.590 2718.450 2147.890 2718.815 ;
        RECT 2146.885 2718.150 2147.890 2718.450 ;
        RECT 2146.885 2718.135 2147.215 2718.150 ;
        RECT 2145.965 2704.850 2146.295 2704.865 ;
        RECT 2146.885 2704.850 2147.215 2704.865 ;
        RECT 2145.965 2704.550 2147.215 2704.850 ;
        RECT 2145.965 2704.535 2146.295 2704.550 ;
        RECT 2146.885 2704.535 2147.215 2704.550 ;
        RECT 2146.885 2608.290 2147.215 2608.305 ;
        RECT 2147.805 2608.290 2148.135 2608.305 ;
        RECT 2146.885 2607.990 2148.135 2608.290 ;
        RECT 2146.885 2607.975 2147.215 2607.990 ;
        RECT 2147.805 2607.975 2148.135 2607.990 ;
        RECT 2147.345 2318.610 2147.675 2318.625 ;
        RECT 2148.265 2318.610 2148.595 2318.625 ;
        RECT 2147.345 2318.310 2148.595 2318.610 ;
        RECT 2147.345 2318.295 2147.675 2318.310 ;
        RECT 2148.265 2318.295 2148.595 2318.310 ;
        RECT 285.265 1542.050 285.595 1542.065 ;
        RECT 285.265 1541.920 300.380 1542.050 ;
        RECT 285.265 1541.750 304.000 1541.920 ;
        RECT 285.265 1541.735 285.595 1541.750 ;
        RECT 300.000 1541.320 304.000 1541.750 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 681.790 3503.260 682.110 3503.320 ;
        RECT 1824.890 3503.260 1825.210 3503.320 ;
        RECT 681.790 3503.120 1825.210 3503.260 ;
        RECT 681.790 3503.060 682.110 3503.120 ;
        RECT 1824.890 3503.060 1825.210 3503.120 ;
        RECT 284.810 2199.360 285.130 2199.420 ;
        RECT 681.790 2199.360 682.110 2199.420 ;
        RECT 284.810 2199.220 682.110 2199.360 ;
        RECT 284.810 2199.160 285.130 2199.220 ;
        RECT 681.790 2199.160 682.110 2199.220 ;
      LAYER via ;
        RECT 681.820 3503.060 682.080 3503.320 ;
        RECT 1824.920 3503.060 1825.180 3503.320 ;
        RECT 284.840 2199.160 285.100 2199.420 ;
        RECT 681.820 2199.160 682.080 2199.420 ;
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
        RECT 1824.980 3503.350 1825.120 3517.600 ;
        RECT 681.820 3503.030 682.080 3503.350 ;
        RECT 1824.920 3503.030 1825.180 3503.350 ;
        RECT 681.880 2199.450 682.020 3503.030 ;
        RECT 284.840 2199.130 285.100 2199.450 ;
        RECT 681.820 2199.130 682.080 2199.450 ;
        RECT 284.900 1574.045 285.040 2199.130 ;
        RECT 284.830 1573.675 285.110 1574.045 ;
      LAYER via2 ;
        RECT 284.830 1573.720 285.110 1574.000 ;
      LAYER met3 ;
        RECT 284.805 1574.010 285.135 1574.025 ;
        RECT 284.805 1573.880 300.380 1574.010 ;
        RECT 284.805 1573.710 304.000 1573.880 ;
        RECT 284.805 1573.695 285.135 1573.710 ;
        RECT 300.000 1573.280 304.000 1573.710 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1498.290 3443.080 1498.610 3443.140 ;
        RECT 1500.590 3443.080 1500.910 3443.140 ;
        RECT 1498.290 3442.940 1500.910 3443.080 ;
        RECT 1498.290 3442.880 1498.610 3442.940 ;
        RECT 1500.590 3442.880 1500.910 3442.940 ;
        RECT 1497.830 3422.340 1498.150 3422.400 ;
        RECT 1498.290 3422.340 1498.610 3422.400 ;
        RECT 1497.830 3422.200 1498.610 3422.340 ;
        RECT 1497.830 3422.140 1498.150 3422.200 ;
        RECT 1498.290 3422.140 1498.610 3422.200 ;
        RECT 1498.290 3394.940 1498.610 3395.200 ;
        RECT 1498.380 3394.520 1498.520 3394.940 ;
        RECT 1498.290 3394.260 1498.610 3394.520 ;
        RECT 1498.290 3332.920 1498.610 3332.980 ;
        RECT 1499.670 3332.920 1499.990 3332.980 ;
        RECT 1498.290 3332.780 1499.990 3332.920 ;
        RECT 1498.290 3332.720 1498.610 3332.780 ;
        RECT 1499.670 3332.720 1499.990 3332.780 ;
        RECT 1498.290 3308.780 1498.610 3308.840 ;
        RECT 1499.670 3308.780 1499.990 3308.840 ;
        RECT 1498.290 3308.640 1499.990 3308.780 ;
        RECT 1498.290 3308.580 1498.610 3308.640 ;
        RECT 1499.670 3308.580 1499.990 3308.640 ;
        RECT 1498.290 3284.640 1498.610 3284.700 ;
        RECT 1498.750 3284.640 1499.070 3284.700 ;
        RECT 1498.290 3284.500 1499.070 3284.640 ;
        RECT 1498.290 3284.440 1498.610 3284.500 ;
        RECT 1498.750 3284.440 1499.070 3284.500 ;
        RECT 1498.290 3236.360 1498.610 3236.420 ;
        RECT 1498.750 3236.360 1499.070 3236.420 ;
        RECT 1498.290 3236.220 1499.070 3236.360 ;
        RECT 1498.290 3236.160 1498.610 3236.220 ;
        RECT 1498.750 3236.160 1499.070 3236.220 ;
        RECT 1498.290 3202.020 1498.610 3202.080 ;
        RECT 1498.750 3202.020 1499.070 3202.080 ;
        RECT 1498.290 3201.880 1499.070 3202.020 ;
        RECT 1498.290 3201.820 1498.610 3201.880 ;
        RECT 1498.750 3201.820 1499.070 3201.880 ;
        RECT 1497.830 3153.400 1498.150 3153.460 ;
        RECT 1498.750 3153.400 1499.070 3153.460 ;
        RECT 1497.830 3153.260 1499.070 3153.400 ;
        RECT 1497.830 3153.200 1498.150 3153.260 ;
        RECT 1498.750 3153.200 1499.070 3153.260 ;
        RECT 1497.830 3056.840 1498.150 3056.900 ;
        RECT 1498.750 3056.840 1499.070 3056.900 ;
        RECT 1497.830 3056.700 1499.070 3056.840 ;
        RECT 1497.830 3056.640 1498.150 3056.700 ;
        RECT 1498.750 3056.640 1499.070 3056.700 ;
        RECT 1498.290 2995.300 1498.610 2995.360 ;
        RECT 1499.210 2995.300 1499.530 2995.360 ;
        RECT 1498.290 2995.160 1499.530 2995.300 ;
        RECT 1498.290 2995.100 1498.610 2995.160 ;
        RECT 1499.210 2995.100 1499.530 2995.160 ;
        RECT 1498.290 2994.620 1498.610 2994.680 ;
        RECT 1499.210 2994.620 1499.530 2994.680 ;
        RECT 1498.290 2994.480 1499.530 2994.620 ;
        RECT 1498.290 2994.420 1498.610 2994.480 ;
        RECT 1499.210 2994.420 1499.530 2994.480 ;
        RECT 1498.290 2946.680 1498.610 2946.740 ;
        RECT 1499.670 2946.680 1499.990 2946.740 ;
        RECT 1498.290 2946.540 1499.990 2946.680 ;
        RECT 1498.290 2946.480 1498.610 2946.540 ;
        RECT 1499.670 2946.480 1499.990 2946.540 ;
        RECT 1499.670 2912.340 1499.990 2912.400 ;
        RECT 1499.300 2912.200 1499.990 2912.340 ;
        RECT 1499.300 2911.720 1499.440 2912.200 ;
        RECT 1499.670 2912.140 1499.990 2912.200 ;
        RECT 1499.210 2911.460 1499.530 2911.720 ;
        RECT 1497.830 2815.580 1498.150 2815.840 ;
        RECT 1497.920 2815.160 1498.060 2815.580 ;
        RECT 1497.830 2814.900 1498.150 2815.160 ;
        RECT 1497.830 2767.500 1498.150 2767.560 ;
        RECT 1497.460 2767.360 1498.150 2767.500 ;
        RECT 1497.460 2766.880 1497.600 2767.360 ;
        RECT 1497.830 2767.300 1498.150 2767.360 ;
        RECT 1497.370 2766.620 1497.690 2766.880 ;
        RECT 1497.370 2746.080 1497.690 2746.140 ;
        RECT 1497.830 2746.080 1498.150 2746.140 ;
        RECT 1497.370 2745.940 1498.150 2746.080 ;
        RECT 1497.370 2745.880 1497.690 2745.940 ;
        RECT 1497.830 2745.880 1498.150 2745.940 ;
        RECT 1497.830 2718.680 1498.150 2718.940 ;
        RECT 1497.920 2718.260 1498.060 2718.680 ;
        RECT 1497.830 2718.000 1498.150 2718.260 ;
        RECT 1497.830 2656.660 1498.150 2656.720 ;
        RECT 1498.290 2656.660 1498.610 2656.720 ;
        RECT 1497.830 2656.520 1498.610 2656.660 ;
        RECT 1497.830 2656.460 1498.150 2656.520 ;
        RECT 1498.290 2656.460 1498.610 2656.520 ;
        RECT 1497.370 2608.380 1497.690 2608.440 ;
        RECT 1498.750 2608.380 1499.070 2608.440 ;
        RECT 1497.370 2608.240 1499.070 2608.380 ;
        RECT 1497.370 2608.180 1497.690 2608.240 ;
        RECT 1498.750 2608.180 1499.070 2608.240 ;
        RECT 1497.370 2511.820 1497.690 2511.880 ;
        RECT 1498.750 2511.820 1499.070 2511.880 ;
        RECT 1497.370 2511.680 1499.070 2511.820 ;
        RECT 1497.370 2511.620 1497.690 2511.680 ;
        RECT 1498.750 2511.620 1499.070 2511.680 ;
        RECT 1497.370 2463.200 1497.690 2463.260 ;
        RECT 1498.290 2463.200 1498.610 2463.260 ;
        RECT 1497.370 2463.060 1498.610 2463.200 ;
        RECT 1497.370 2463.000 1497.690 2463.060 ;
        RECT 1498.290 2463.000 1498.610 2463.060 ;
        RECT 1498.290 2332.100 1498.610 2332.360 ;
        RECT 1498.380 2331.960 1498.520 2332.100 ;
        RECT 1498.750 2331.960 1499.070 2332.020 ;
        RECT 1498.380 2331.820 1499.070 2331.960 ;
        RECT 1498.750 2331.760 1499.070 2331.820 ;
        RECT 1498.750 2318.360 1499.070 2318.420 ;
        RECT 1499.210 2318.360 1499.530 2318.420 ;
        RECT 1498.750 2318.220 1499.530 2318.360 ;
        RECT 1498.750 2318.160 1499.070 2318.220 ;
        RECT 1499.210 2318.160 1499.530 2318.220 ;
        RECT 1499.210 2284.020 1499.530 2284.080 ;
        RECT 1498.840 2283.880 1499.530 2284.020 ;
        RECT 1498.840 2283.740 1498.980 2283.880 ;
        RECT 1499.210 2283.820 1499.530 2283.880 ;
        RECT 1498.750 2283.480 1499.070 2283.740 ;
        RECT 1498.290 2222.140 1498.610 2222.200 ;
        RECT 1499.210 2222.140 1499.530 2222.200 ;
        RECT 1498.290 2222.000 1499.530 2222.140 ;
        RECT 1498.290 2221.940 1498.610 2222.000 ;
        RECT 1499.210 2221.940 1499.530 2222.000 ;
        RECT 284.350 2198.680 284.670 2198.740 ;
        RECT 1498.290 2198.680 1498.610 2198.740 ;
        RECT 284.350 2198.540 1498.610 2198.680 ;
        RECT 284.350 2198.480 284.670 2198.540 ;
        RECT 1498.290 2198.480 1498.610 2198.540 ;
      LAYER via ;
        RECT 1498.320 3442.880 1498.580 3443.140 ;
        RECT 1500.620 3442.880 1500.880 3443.140 ;
        RECT 1497.860 3422.140 1498.120 3422.400 ;
        RECT 1498.320 3422.140 1498.580 3422.400 ;
        RECT 1498.320 3394.940 1498.580 3395.200 ;
        RECT 1498.320 3394.260 1498.580 3394.520 ;
        RECT 1498.320 3332.720 1498.580 3332.980 ;
        RECT 1499.700 3332.720 1499.960 3332.980 ;
        RECT 1498.320 3308.580 1498.580 3308.840 ;
        RECT 1499.700 3308.580 1499.960 3308.840 ;
        RECT 1498.320 3284.440 1498.580 3284.700 ;
        RECT 1498.780 3284.440 1499.040 3284.700 ;
        RECT 1498.320 3236.160 1498.580 3236.420 ;
        RECT 1498.780 3236.160 1499.040 3236.420 ;
        RECT 1498.320 3201.820 1498.580 3202.080 ;
        RECT 1498.780 3201.820 1499.040 3202.080 ;
        RECT 1497.860 3153.200 1498.120 3153.460 ;
        RECT 1498.780 3153.200 1499.040 3153.460 ;
        RECT 1497.860 3056.640 1498.120 3056.900 ;
        RECT 1498.780 3056.640 1499.040 3056.900 ;
        RECT 1498.320 2995.100 1498.580 2995.360 ;
        RECT 1499.240 2995.100 1499.500 2995.360 ;
        RECT 1498.320 2994.420 1498.580 2994.680 ;
        RECT 1499.240 2994.420 1499.500 2994.680 ;
        RECT 1498.320 2946.480 1498.580 2946.740 ;
        RECT 1499.700 2946.480 1499.960 2946.740 ;
        RECT 1499.700 2912.140 1499.960 2912.400 ;
        RECT 1499.240 2911.460 1499.500 2911.720 ;
        RECT 1497.860 2815.580 1498.120 2815.840 ;
        RECT 1497.860 2814.900 1498.120 2815.160 ;
        RECT 1497.860 2767.300 1498.120 2767.560 ;
        RECT 1497.400 2766.620 1497.660 2766.880 ;
        RECT 1497.400 2745.880 1497.660 2746.140 ;
        RECT 1497.860 2745.880 1498.120 2746.140 ;
        RECT 1497.860 2718.680 1498.120 2718.940 ;
        RECT 1497.860 2718.000 1498.120 2718.260 ;
        RECT 1497.860 2656.460 1498.120 2656.720 ;
        RECT 1498.320 2656.460 1498.580 2656.720 ;
        RECT 1497.400 2608.180 1497.660 2608.440 ;
        RECT 1498.780 2608.180 1499.040 2608.440 ;
        RECT 1497.400 2511.620 1497.660 2511.880 ;
        RECT 1498.780 2511.620 1499.040 2511.880 ;
        RECT 1497.400 2463.000 1497.660 2463.260 ;
        RECT 1498.320 2463.000 1498.580 2463.260 ;
        RECT 1498.320 2332.100 1498.580 2332.360 ;
        RECT 1498.780 2331.760 1499.040 2332.020 ;
        RECT 1498.780 2318.160 1499.040 2318.420 ;
        RECT 1499.240 2318.160 1499.500 2318.420 ;
        RECT 1499.240 2283.820 1499.500 2284.080 ;
        RECT 1498.780 2283.480 1499.040 2283.740 ;
        RECT 1498.320 2221.940 1498.580 2222.200 ;
        RECT 1499.240 2221.940 1499.500 2222.200 ;
        RECT 284.380 2198.480 284.640 2198.740 ;
        RECT 1498.320 2198.480 1498.580 2198.740 ;
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
        RECT 1500.680 3443.170 1500.820 3517.600 ;
        RECT 1498.320 3442.850 1498.580 3443.170 ;
        RECT 1500.620 3442.850 1500.880 3443.170 ;
        RECT 1498.380 3429.650 1498.520 3442.850 ;
        RECT 1497.920 3429.510 1498.520 3429.650 ;
        RECT 1497.920 3422.430 1498.060 3429.510 ;
        RECT 1497.860 3422.110 1498.120 3422.430 ;
        RECT 1498.320 3422.110 1498.580 3422.430 ;
        RECT 1498.380 3395.230 1498.520 3422.110 ;
        RECT 1498.320 3394.910 1498.580 3395.230 ;
        RECT 1498.320 3394.230 1498.580 3394.550 ;
        RECT 1498.380 3333.010 1498.520 3394.230 ;
        RECT 1498.320 3332.690 1498.580 3333.010 ;
        RECT 1499.700 3332.690 1499.960 3333.010 ;
        RECT 1499.760 3308.870 1499.900 3332.690 ;
        RECT 1498.320 3308.550 1498.580 3308.870 ;
        RECT 1499.700 3308.550 1499.960 3308.870 ;
        RECT 1498.380 3284.730 1498.520 3308.550 ;
        RECT 1498.320 3284.410 1498.580 3284.730 ;
        RECT 1498.780 3284.410 1499.040 3284.730 ;
        RECT 1498.840 3236.450 1498.980 3284.410 ;
        RECT 1498.320 3236.130 1498.580 3236.450 ;
        RECT 1498.780 3236.130 1499.040 3236.450 ;
        RECT 1498.380 3202.110 1498.520 3236.130 ;
        RECT 1498.320 3201.790 1498.580 3202.110 ;
        RECT 1498.780 3201.790 1499.040 3202.110 ;
        RECT 1498.840 3153.490 1498.980 3201.790 ;
        RECT 1497.860 3153.170 1498.120 3153.490 ;
        RECT 1498.780 3153.170 1499.040 3153.490 ;
        RECT 1497.920 3152.890 1498.060 3153.170 ;
        RECT 1497.920 3152.750 1498.520 3152.890 ;
        RECT 1498.380 3105.290 1498.520 3152.750 ;
        RECT 1498.380 3105.150 1498.980 3105.290 ;
        RECT 1498.840 3056.930 1498.980 3105.150 ;
        RECT 1497.860 3056.610 1498.120 3056.930 ;
        RECT 1498.780 3056.610 1499.040 3056.930 ;
        RECT 1497.920 3056.330 1498.060 3056.610 ;
        RECT 1497.920 3056.190 1498.520 3056.330 ;
        RECT 1498.380 2995.390 1498.520 3056.190 ;
        RECT 1498.320 2995.070 1498.580 2995.390 ;
        RECT 1499.240 2995.070 1499.500 2995.390 ;
        RECT 1499.300 2994.710 1499.440 2995.070 ;
        RECT 1498.320 2994.390 1498.580 2994.710 ;
        RECT 1499.240 2994.390 1499.500 2994.710 ;
        RECT 1498.380 2946.770 1498.520 2994.390 ;
        RECT 1498.320 2946.450 1498.580 2946.770 ;
        RECT 1499.700 2946.450 1499.960 2946.770 ;
        RECT 1499.760 2912.430 1499.900 2946.450 ;
        RECT 1499.700 2912.110 1499.960 2912.430 ;
        RECT 1499.240 2911.430 1499.500 2911.750 ;
        RECT 1499.300 2863.210 1499.440 2911.430 ;
        RECT 1498.380 2863.070 1499.440 2863.210 ;
        RECT 1498.380 2849.610 1498.520 2863.070 ;
        RECT 1497.920 2849.470 1498.520 2849.610 ;
        RECT 1497.920 2815.870 1498.060 2849.470 ;
        RECT 1497.860 2815.550 1498.120 2815.870 ;
        RECT 1497.860 2814.870 1498.120 2815.190 ;
        RECT 1497.920 2767.590 1498.060 2814.870 ;
        RECT 1497.860 2767.270 1498.120 2767.590 ;
        RECT 1497.400 2766.590 1497.660 2766.910 ;
        RECT 1497.460 2746.170 1497.600 2766.590 ;
        RECT 1497.400 2745.850 1497.660 2746.170 ;
        RECT 1497.860 2745.850 1498.120 2746.170 ;
        RECT 1497.920 2718.970 1498.060 2745.850 ;
        RECT 1497.860 2718.650 1498.120 2718.970 ;
        RECT 1497.860 2717.970 1498.120 2718.290 ;
        RECT 1497.920 2656.750 1498.060 2717.970 ;
        RECT 1497.390 2656.235 1497.670 2656.605 ;
        RECT 1497.860 2656.430 1498.120 2656.750 ;
        RECT 1498.320 2656.605 1498.580 2656.750 ;
        RECT 1498.310 2656.235 1498.590 2656.605 ;
        RECT 1497.460 2608.470 1497.600 2656.235 ;
        RECT 1497.400 2608.150 1497.660 2608.470 ;
        RECT 1498.780 2608.150 1499.040 2608.470 ;
        RECT 1498.840 2573.530 1498.980 2608.150 ;
        RECT 1498.380 2573.390 1498.980 2573.530 ;
        RECT 1498.380 2560.045 1498.520 2573.390 ;
        RECT 1497.390 2559.675 1497.670 2560.045 ;
        RECT 1498.310 2559.675 1498.590 2560.045 ;
        RECT 1497.460 2511.910 1497.600 2559.675 ;
        RECT 1497.400 2511.590 1497.660 2511.910 ;
        RECT 1498.780 2511.590 1499.040 2511.910 ;
        RECT 1498.840 2476.970 1498.980 2511.590 ;
        RECT 1498.380 2476.830 1498.980 2476.970 ;
        RECT 1498.380 2463.290 1498.520 2476.830 ;
        RECT 1497.400 2462.970 1497.660 2463.290 ;
        RECT 1498.320 2462.970 1498.580 2463.290 ;
        RECT 1497.460 2415.205 1497.600 2462.970 ;
        RECT 1497.390 2414.835 1497.670 2415.205 ;
        RECT 1498.770 2414.835 1499.050 2415.205 ;
        RECT 1498.840 2380.410 1498.980 2414.835 ;
        RECT 1498.380 2380.270 1498.980 2380.410 ;
        RECT 1498.380 2332.390 1498.520 2380.270 ;
        RECT 1498.320 2332.070 1498.580 2332.390 ;
        RECT 1498.780 2331.730 1499.040 2332.050 ;
        RECT 1498.840 2318.450 1498.980 2331.730 ;
        RECT 1498.780 2318.130 1499.040 2318.450 ;
        RECT 1499.240 2318.130 1499.500 2318.450 ;
        RECT 1499.300 2284.110 1499.440 2318.130 ;
        RECT 1499.240 2283.790 1499.500 2284.110 ;
        RECT 1498.780 2283.450 1499.040 2283.770 ;
        RECT 1498.840 2270.250 1498.980 2283.450 ;
        RECT 1498.840 2270.110 1499.440 2270.250 ;
        RECT 1499.300 2222.230 1499.440 2270.110 ;
        RECT 1498.320 2221.910 1498.580 2222.230 ;
        RECT 1499.240 2221.910 1499.500 2222.230 ;
        RECT 1498.380 2198.770 1498.520 2221.910 ;
        RECT 284.380 2198.450 284.640 2198.770 ;
        RECT 1498.320 2198.450 1498.580 2198.770 ;
        RECT 284.440 1605.325 284.580 2198.450 ;
        RECT 284.370 1604.955 284.650 1605.325 ;
      LAYER via2 ;
        RECT 1497.390 2656.280 1497.670 2656.560 ;
        RECT 1498.310 2656.280 1498.590 2656.560 ;
        RECT 1497.390 2559.720 1497.670 2560.000 ;
        RECT 1498.310 2559.720 1498.590 2560.000 ;
        RECT 1497.390 2414.880 1497.670 2415.160 ;
        RECT 1498.770 2414.880 1499.050 2415.160 ;
        RECT 284.370 1605.000 284.650 1605.280 ;
      LAYER met3 ;
        RECT 1497.365 2656.570 1497.695 2656.585 ;
        RECT 1498.285 2656.570 1498.615 2656.585 ;
        RECT 1497.365 2656.270 1498.615 2656.570 ;
        RECT 1497.365 2656.255 1497.695 2656.270 ;
        RECT 1498.285 2656.255 1498.615 2656.270 ;
        RECT 1497.365 2560.010 1497.695 2560.025 ;
        RECT 1498.285 2560.010 1498.615 2560.025 ;
        RECT 1497.365 2559.710 1498.615 2560.010 ;
        RECT 1497.365 2559.695 1497.695 2559.710 ;
        RECT 1498.285 2559.695 1498.615 2559.710 ;
        RECT 1497.365 2415.170 1497.695 2415.185 ;
        RECT 1498.745 2415.170 1499.075 2415.185 ;
        RECT 1497.365 2414.870 1499.075 2415.170 ;
        RECT 1497.365 2414.855 1497.695 2414.870 ;
        RECT 1498.745 2414.855 1499.075 2414.870 ;
        RECT 284.345 1605.290 284.675 1605.305 ;
        RECT 284.345 1605.160 300.380 1605.290 ;
        RECT 284.345 1604.990 304.000 1605.160 ;
        RECT 284.345 1604.975 284.675 1604.990 ;
        RECT 300.000 1604.560 304.000 1604.990 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 444.430 319.500 444.750 319.560 ;
        RECT 482.610 319.500 482.930 319.560 ;
        RECT 444.430 319.360 482.930 319.500 ;
        RECT 444.430 319.300 444.750 319.360 ;
        RECT 482.610 319.300 482.930 319.360 ;
        RECT 737.910 318.820 738.230 318.880 ;
        RECT 772.410 318.820 772.730 318.880 ;
        RECT 737.910 318.680 772.730 318.820 ;
        RECT 737.910 318.620 738.230 318.680 ;
        RECT 772.410 318.620 772.730 318.680 ;
        RECT 580.130 318.140 580.450 318.200 ;
        RECT 593.930 318.140 594.250 318.200 ;
        RECT 580.130 318.000 594.250 318.140 ;
        RECT 580.130 317.940 580.450 318.000 ;
        RECT 593.930 317.940 594.250 318.000 ;
      LAYER via ;
        RECT 444.460 319.300 444.720 319.560 ;
        RECT 482.640 319.300 482.900 319.560 ;
        RECT 737.940 318.620 738.200 318.880 ;
        RECT 772.440 318.620 772.700 318.880 ;
        RECT 580.160 317.940 580.420 318.200 ;
        RECT 593.960 317.940 594.220 318.200 ;
      LAYER met2 ;
        RECT 675.830 320.435 676.110 320.805 ;
        RECT 444.460 319.445 444.720 319.590 ;
        RECT 482.640 319.445 482.900 319.590 ;
        RECT 444.450 319.075 444.730 319.445 ;
        RECT 482.630 319.075 482.910 319.445 ;
        RECT 593.950 319.075 594.230 319.445 ;
        RECT 594.020 318.230 594.160 319.075 ;
        RECT 675.900 318.765 676.040 320.435 ;
        RECT 700.210 319.755 700.490 320.125 ;
        RECT 675.830 318.395 676.110 318.765 ;
        RECT 580.160 318.085 580.420 318.230 ;
        RECT 580.150 317.715 580.430 318.085 ;
        RECT 593.960 317.910 594.220 318.230 ;
        RECT 700.280 318.085 700.420 319.755 ;
        RECT 772.430 319.075 772.710 319.445 ;
        RECT 772.500 318.910 772.640 319.075 ;
        RECT 737.940 318.765 738.200 318.910 ;
        RECT 737.930 318.395 738.210 318.765 ;
        RECT 772.440 318.590 772.700 318.910 ;
        RECT 700.210 317.715 700.490 318.085 ;
      LAYER via2 ;
        RECT 675.830 320.480 676.110 320.760 ;
        RECT 444.450 319.120 444.730 319.400 ;
        RECT 482.630 319.120 482.910 319.400 ;
        RECT 593.950 319.120 594.230 319.400 ;
        RECT 700.210 319.800 700.490 320.080 ;
        RECT 675.830 318.440 676.110 318.720 ;
        RECT 580.150 317.760 580.430 318.040 ;
        RECT 772.430 319.120 772.710 319.400 ;
        RECT 737.930 318.440 738.210 318.720 ;
        RECT 700.210 317.760 700.490 318.040 ;
      LAYER met3 ;
        RECT 287.310 1036.810 287.690 1036.820 ;
        RECT 287.310 1036.680 300.380 1036.810 ;
        RECT 287.310 1036.510 304.000 1036.680 ;
        RECT 287.310 1036.500 287.690 1036.510 ;
        RECT 300.000 1036.080 304.000 1036.510 ;
        RECT 2917.600 322.810 2924.800 323.260 ;
        RECT 2916.710 322.510 2924.800 322.810 ;
        RECT 627.710 320.770 628.090 320.780 ;
        RECT 675.805 320.770 676.135 320.785 ;
        RECT 627.710 320.470 676.135 320.770 ;
        RECT 627.710 320.460 628.090 320.470 ;
        RECT 675.805 320.455 676.135 320.470 ;
        RECT 578.950 320.090 579.330 320.100 ;
        RECT 700.185 320.090 700.515 320.105 ;
        RECT 544.030 319.790 579.330 320.090 ;
        RECT 287.310 319.410 287.690 319.420 ;
        RECT 444.425 319.410 444.755 319.425 ;
        RECT 287.310 319.110 324.450 319.410 ;
        RECT 287.310 319.100 287.690 319.110 ;
        RECT 324.150 318.730 324.450 319.110 ;
        RECT 372.910 319.110 444.755 319.410 ;
        RECT 324.150 318.430 372.290 318.730 ;
        RECT 371.990 318.050 372.290 318.430 ;
        RECT 372.910 318.050 373.210 319.110 ;
        RECT 444.425 319.095 444.755 319.110 ;
        RECT 482.605 319.410 482.935 319.425 ;
        RECT 482.605 319.110 496.490 319.410 ;
        RECT 482.605 319.095 482.935 319.110 ;
        RECT 371.990 317.750 373.210 318.050 ;
        RECT 496.190 318.050 496.490 319.110 ;
        RECT 544.030 318.730 544.330 319.790 ;
        RECT 578.950 319.780 579.330 319.790 ;
        RECT 676.510 319.790 700.515 320.090 ;
        RECT 593.925 319.410 594.255 319.425 ;
        RECT 627.710 319.410 628.090 319.420 ;
        RECT 593.925 319.110 628.090 319.410 ;
        RECT 593.925 319.095 594.255 319.110 ;
        RECT 627.710 319.100 628.090 319.110 ;
        RECT 497.110 318.430 544.330 318.730 ;
        RECT 675.805 318.730 676.135 318.745 ;
        RECT 676.510 318.730 676.810 319.790 ;
        RECT 700.185 319.775 700.515 319.790 ;
        RECT 772.405 319.410 772.735 319.425 ;
        RECT 772.405 319.110 807.450 319.410 ;
        RECT 772.405 319.095 772.735 319.110 ;
        RECT 737.905 318.730 738.235 318.745 ;
        RECT 675.805 318.430 676.810 318.730 ;
        RECT 724.350 318.430 738.235 318.730 ;
        RECT 807.150 318.730 807.450 319.110 ;
        RECT 855.910 319.110 904.050 319.410 ;
        RECT 807.150 318.430 855.290 318.730 ;
        RECT 497.110 318.050 497.410 318.430 ;
        RECT 675.805 318.415 676.135 318.430 ;
        RECT 496.190 317.750 497.410 318.050 ;
        RECT 578.950 318.050 579.330 318.060 ;
        RECT 580.125 318.050 580.455 318.065 ;
        RECT 578.950 317.750 580.455 318.050 ;
        RECT 578.950 317.740 579.330 317.750 ;
        RECT 580.125 317.735 580.455 317.750 ;
        RECT 700.185 318.050 700.515 318.065 ;
        RECT 724.350 318.050 724.650 318.430 ;
        RECT 737.905 318.415 738.235 318.430 ;
        RECT 700.185 317.750 724.650 318.050 ;
        RECT 854.990 318.050 855.290 318.430 ;
        RECT 855.910 318.050 856.210 319.110 ;
        RECT 903.750 318.730 904.050 319.110 ;
        RECT 952.510 319.110 1000.650 319.410 ;
        RECT 903.750 318.430 951.890 318.730 ;
        RECT 854.990 317.750 856.210 318.050 ;
        RECT 951.590 318.050 951.890 318.430 ;
        RECT 952.510 318.050 952.810 319.110 ;
        RECT 1000.350 318.730 1000.650 319.110 ;
        RECT 1049.110 319.110 1097.250 319.410 ;
        RECT 1000.350 318.430 1048.490 318.730 ;
        RECT 951.590 317.750 952.810 318.050 ;
        RECT 1048.190 318.050 1048.490 318.430 ;
        RECT 1049.110 318.050 1049.410 319.110 ;
        RECT 1096.950 318.730 1097.250 319.110 ;
        RECT 1145.710 319.110 1193.850 319.410 ;
        RECT 1096.950 318.430 1145.090 318.730 ;
        RECT 1048.190 317.750 1049.410 318.050 ;
        RECT 1144.790 318.050 1145.090 318.430 ;
        RECT 1145.710 318.050 1146.010 319.110 ;
        RECT 1193.550 318.730 1193.850 319.110 ;
        RECT 1242.310 319.110 1290.450 319.410 ;
        RECT 1193.550 318.430 1241.690 318.730 ;
        RECT 1144.790 317.750 1146.010 318.050 ;
        RECT 1241.390 318.050 1241.690 318.430 ;
        RECT 1242.310 318.050 1242.610 319.110 ;
        RECT 1290.150 318.730 1290.450 319.110 ;
        RECT 1338.910 319.110 1387.050 319.410 ;
        RECT 1290.150 318.430 1338.290 318.730 ;
        RECT 1241.390 317.750 1242.610 318.050 ;
        RECT 1337.990 318.050 1338.290 318.430 ;
        RECT 1338.910 318.050 1339.210 319.110 ;
        RECT 1386.750 318.730 1387.050 319.110 ;
        RECT 1435.510 319.110 1483.650 319.410 ;
        RECT 1386.750 318.430 1434.890 318.730 ;
        RECT 1337.990 317.750 1339.210 318.050 ;
        RECT 1434.590 318.050 1434.890 318.430 ;
        RECT 1435.510 318.050 1435.810 319.110 ;
        RECT 1483.350 318.730 1483.650 319.110 ;
        RECT 1532.110 319.110 1580.250 319.410 ;
        RECT 1483.350 318.430 1531.490 318.730 ;
        RECT 1434.590 317.750 1435.810 318.050 ;
        RECT 1531.190 318.050 1531.490 318.430 ;
        RECT 1532.110 318.050 1532.410 319.110 ;
        RECT 1579.950 318.730 1580.250 319.110 ;
        RECT 1628.710 319.110 1676.850 319.410 ;
        RECT 1579.950 318.430 1628.090 318.730 ;
        RECT 1531.190 317.750 1532.410 318.050 ;
        RECT 1627.790 318.050 1628.090 318.430 ;
        RECT 1628.710 318.050 1629.010 319.110 ;
        RECT 1676.550 318.730 1676.850 319.110 ;
        RECT 1725.310 319.110 1773.450 319.410 ;
        RECT 1676.550 318.430 1724.690 318.730 ;
        RECT 1627.790 317.750 1629.010 318.050 ;
        RECT 1724.390 318.050 1724.690 318.430 ;
        RECT 1725.310 318.050 1725.610 319.110 ;
        RECT 1773.150 318.730 1773.450 319.110 ;
        RECT 1821.910 319.110 1870.050 319.410 ;
        RECT 1773.150 318.430 1821.290 318.730 ;
        RECT 1724.390 317.750 1725.610 318.050 ;
        RECT 1820.990 318.050 1821.290 318.430 ;
        RECT 1821.910 318.050 1822.210 319.110 ;
        RECT 1869.750 318.730 1870.050 319.110 ;
        RECT 1918.510 319.110 1966.650 319.410 ;
        RECT 1869.750 318.430 1917.890 318.730 ;
        RECT 1820.990 317.750 1822.210 318.050 ;
        RECT 1917.590 318.050 1917.890 318.430 ;
        RECT 1918.510 318.050 1918.810 319.110 ;
        RECT 1966.350 318.730 1966.650 319.110 ;
        RECT 2015.110 319.110 2063.250 319.410 ;
        RECT 1966.350 318.430 2014.490 318.730 ;
        RECT 1917.590 317.750 1918.810 318.050 ;
        RECT 2014.190 318.050 2014.490 318.430 ;
        RECT 2015.110 318.050 2015.410 319.110 ;
        RECT 2062.950 318.730 2063.250 319.110 ;
        RECT 2111.710 319.110 2159.850 319.410 ;
        RECT 2062.950 318.430 2111.090 318.730 ;
        RECT 2014.190 317.750 2015.410 318.050 ;
        RECT 2110.790 318.050 2111.090 318.430 ;
        RECT 2111.710 318.050 2112.010 319.110 ;
        RECT 2159.550 318.730 2159.850 319.110 ;
        RECT 2208.310 319.110 2256.450 319.410 ;
        RECT 2159.550 318.430 2207.690 318.730 ;
        RECT 2110.790 317.750 2112.010 318.050 ;
        RECT 2207.390 318.050 2207.690 318.430 ;
        RECT 2208.310 318.050 2208.610 319.110 ;
        RECT 2256.150 318.730 2256.450 319.110 ;
        RECT 2304.910 319.110 2353.050 319.410 ;
        RECT 2256.150 318.430 2304.290 318.730 ;
        RECT 2207.390 317.750 2208.610 318.050 ;
        RECT 2303.990 318.050 2304.290 318.430 ;
        RECT 2304.910 318.050 2305.210 319.110 ;
        RECT 2352.750 318.730 2353.050 319.110 ;
        RECT 2401.510 319.110 2449.650 319.410 ;
        RECT 2352.750 318.430 2400.890 318.730 ;
        RECT 2303.990 317.750 2305.210 318.050 ;
        RECT 2400.590 318.050 2400.890 318.430 ;
        RECT 2401.510 318.050 2401.810 319.110 ;
        RECT 2449.350 318.730 2449.650 319.110 ;
        RECT 2498.110 319.110 2546.250 319.410 ;
        RECT 2449.350 318.430 2497.490 318.730 ;
        RECT 2400.590 317.750 2401.810 318.050 ;
        RECT 2497.190 318.050 2497.490 318.430 ;
        RECT 2498.110 318.050 2498.410 319.110 ;
        RECT 2545.950 318.730 2546.250 319.110 ;
        RECT 2594.710 319.110 2642.850 319.410 ;
        RECT 2545.950 318.430 2594.090 318.730 ;
        RECT 2497.190 317.750 2498.410 318.050 ;
        RECT 2593.790 318.050 2594.090 318.430 ;
        RECT 2594.710 318.050 2595.010 319.110 ;
        RECT 2642.550 318.730 2642.850 319.110 ;
        RECT 2691.310 319.110 2739.450 319.410 ;
        RECT 2642.550 318.430 2690.690 318.730 ;
        RECT 2593.790 317.750 2595.010 318.050 ;
        RECT 2690.390 318.050 2690.690 318.430 ;
        RECT 2691.310 318.050 2691.610 319.110 ;
        RECT 2739.150 318.730 2739.450 319.110 ;
        RECT 2787.910 319.110 2836.050 319.410 ;
        RECT 2739.150 318.430 2787.290 318.730 ;
        RECT 2690.390 317.750 2691.610 318.050 ;
        RECT 2786.990 318.050 2787.290 318.430 ;
        RECT 2787.910 318.050 2788.210 319.110 ;
        RECT 2835.750 318.730 2836.050 319.110 ;
        RECT 2916.710 318.730 2917.010 322.510 ;
        RECT 2917.600 322.060 2924.800 322.510 ;
        RECT 2835.750 318.430 2883.890 318.730 ;
        RECT 2786.990 317.750 2788.210 318.050 ;
        RECT 2883.590 318.050 2883.890 318.430 ;
        RECT 2884.510 318.430 2917.010 318.730 ;
        RECT 2884.510 318.050 2884.810 318.430 ;
        RECT 2883.590 317.750 2884.810 318.050 ;
        RECT 700.185 317.735 700.515 317.750 ;
      LAYER via3 ;
        RECT 287.340 1036.500 287.660 1036.820 ;
        RECT 627.740 320.460 628.060 320.780 ;
        RECT 287.340 319.100 287.660 319.420 ;
        RECT 578.980 319.780 579.300 320.100 ;
        RECT 627.740 319.100 628.060 319.420 ;
        RECT 578.980 317.740 579.300 318.060 ;
      LAYER met4 ;
        RECT 287.335 1036.495 287.665 1036.825 ;
        RECT 287.350 319.425 287.650 1036.495 ;
        RECT 627.735 320.455 628.065 320.785 ;
        RECT 578.975 319.775 579.305 320.105 ;
        RECT 287.335 319.095 287.665 319.425 ;
        RECT 578.990 318.065 579.290 319.775 ;
        RECT 627.750 319.425 628.050 320.455 ;
        RECT 627.735 319.095 628.065 319.425 ;
        RECT 578.975 317.735 579.305 318.065 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 682.250 3501.220 682.570 3501.280 ;
        RECT 1175.830 3501.220 1176.150 3501.280 ;
        RECT 682.250 3501.080 1176.150 3501.220 ;
        RECT 682.250 3501.020 682.570 3501.080 ;
        RECT 1175.830 3501.020 1176.150 3501.080 ;
        RECT 283.890 2199.020 284.210 2199.080 ;
        RECT 682.250 2199.020 682.570 2199.080 ;
        RECT 283.890 2198.880 682.570 2199.020 ;
        RECT 283.890 2198.820 284.210 2198.880 ;
        RECT 682.250 2198.820 682.570 2198.880 ;
      LAYER via ;
        RECT 682.280 3501.020 682.540 3501.280 ;
        RECT 1175.860 3501.020 1176.120 3501.280 ;
        RECT 283.920 2198.820 284.180 2199.080 ;
        RECT 682.280 2198.820 682.540 2199.080 ;
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
        RECT 1175.920 3501.310 1176.060 3517.600 ;
        RECT 682.280 3500.990 682.540 3501.310 ;
        RECT 1175.860 3500.990 1176.120 3501.310 ;
        RECT 682.340 2199.110 682.480 3500.990 ;
        RECT 283.920 2198.790 284.180 2199.110 ;
        RECT 682.280 2198.790 682.540 2199.110 ;
        RECT 283.980 1636.605 284.120 2198.790 ;
        RECT 283.910 1636.235 284.190 1636.605 ;
      LAYER via2 ;
        RECT 283.910 1636.280 284.190 1636.560 ;
      LAYER met3 ;
        RECT 283.885 1636.570 284.215 1636.585 ;
        RECT 283.885 1636.440 300.380 1636.570 ;
        RECT 283.885 1636.270 304.000 1636.440 ;
        RECT 283.885 1636.255 284.215 1636.270 ;
        RECT 300.000 1635.840 304.000 1636.270 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 288.490 3504.960 288.810 3505.020 ;
        RECT 851.530 3504.960 851.850 3505.020 ;
        RECT 288.490 3504.820 851.850 3504.960 ;
        RECT 288.490 3504.760 288.810 3504.820 ;
        RECT 851.530 3504.760 851.850 3504.820 ;
      LAYER via ;
        RECT 288.520 3504.760 288.780 3505.020 ;
        RECT 851.560 3504.760 851.820 3505.020 ;
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
        RECT 851.620 3505.050 851.760 3517.600 ;
        RECT 288.520 3504.730 288.780 3505.050 ;
        RECT 851.560 3504.730 851.820 3505.050 ;
        RECT 288.580 1668.565 288.720 3504.730 ;
        RECT 288.510 1668.195 288.790 1668.565 ;
      LAYER via2 ;
        RECT 288.510 1668.240 288.790 1668.520 ;
      LAYER met3 ;
        RECT 288.485 1668.530 288.815 1668.545 ;
        RECT 288.485 1668.400 300.380 1668.530 ;
        RECT 288.485 1668.230 304.000 1668.400 ;
        RECT 288.485 1668.215 288.815 1668.230 ;
        RECT 300.000 1667.800 304.000 1668.230 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 297.690 3503.260 298.010 3503.320 ;
        RECT 527.230 3503.260 527.550 3503.320 ;
        RECT 297.690 3503.120 527.550 3503.260 ;
        RECT 297.690 3503.060 298.010 3503.120 ;
        RECT 527.230 3503.060 527.550 3503.120 ;
      LAYER via ;
        RECT 297.720 3503.060 297.980 3503.320 ;
        RECT 527.260 3503.060 527.520 3503.320 ;
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
        RECT 527.320 3503.350 527.460 3517.600 ;
        RECT 297.720 3503.030 297.980 3503.350 ;
        RECT 527.260 3503.030 527.520 3503.350 ;
        RECT 297.780 1699.845 297.920 3503.030 ;
        RECT 297.710 1699.475 297.990 1699.845 ;
      LAYER via2 ;
        RECT 297.710 1699.520 297.990 1699.800 ;
      LAYER met3 ;
        RECT 297.685 1699.810 298.015 1699.825 ;
        RECT 297.685 1699.680 300.380 1699.810 ;
        RECT 297.685 1699.510 304.000 1699.680 ;
        RECT 297.685 1699.495 298.015 1699.510 ;
        RECT 300.000 1699.080 304.000 1699.510 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 202.470 3499.860 202.790 3499.920 ;
        RECT 210.290 3499.860 210.610 3499.920 ;
        RECT 202.470 3499.720 210.610 3499.860 ;
        RECT 202.470 3499.660 202.790 3499.720 ;
        RECT 210.290 3499.660 210.610 3499.720 ;
        RECT 210.290 1731.860 210.610 1731.920 ;
        RECT 282.970 1731.860 283.290 1731.920 ;
        RECT 210.290 1731.720 283.290 1731.860 ;
        RECT 210.290 1731.660 210.610 1731.720 ;
        RECT 282.970 1731.660 283.290 1731.720 ;
      LAYER via ;
        RECT 202.500 3499.660 202.760 3499.920 ;
        RECT 210.320 3499.660 210.580 3499.920 ;
        RECT 210.320 1731.660 210.580 1731.920 ;
        RECT 283.000 1731.660 283.260 1731.920 ;
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
        RECT 202.560 3499.950 202.700 3517.600 ;
        RECT 202.500 3499.630 202.760 3499.950 ;
        RECT 210.320 3499.630 210.580 3499.950 ;
        RECT 210.380 1731.950 210.520 3499.630 ;
        RECT 210.320 1731.630 210.580 1731.950 ;
        RECT 283.000 1731.805 283.260 1731.950 ;
        RECT 282.990 1731.435 283.270 1731.805 ;
      LAYER via2 ;
        RECT 282.990 1731.480 283.270 1731.760 ;
      LAYER met3 ;
        RECT 282.965 1731.770 283.295 1731.785 ;
        RECT 282.965 1731.640 300.380 1731.770 ;
        RECT 282.965 1731.470 304.000 1731.640 ;
        RECT 282.965 1731.455 283.295 1731.470 ;
        RECT 300.000 1731.040 304.000 1731.470 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 23.990 1766.200 24.310 1766.260 ;
        RECT 282.970 1766.200 283.290 1766.260 ;
        RECT 23.990 1766.060 283.290 1766.200 ;
        RECT 23.990 1766.000 24.310 1766.060 ;
        RECT 282.970 1766.000 283.290 1766.060 ;
      LAYER via ;
        RECT 24.020 1766.000 24.280 1766.260 ;
        RECT 283.000 1766.000 283.260 1766.260 ;
      LAYER met2 ;
        RECT 24.010 3411.035 24.290 3411.405 ;
        RECT 24.080 1766.290 24.220 3411.035 ;
        RECT 24.020 1765.970 24.280 1766.290 ;
        RECT 283.000 1765.970 283.260 1766.290 ;
        RECT 283.060 1763.085 283.200 1765.970 ;
        RECT 282.990 1762.715 283.270 1763.085 ;
      LAYER via2 ;
        RECT 24.010 3411.080 24.290 3411.360 ;
        RECT 282.990 1762.760 283.270 1763.040 ;
      LAYER met3 ;
        RECT -4.800 3411.370 2.400 3411.820 ;
        RECT 23.985 3411.370 24.315 3411.385 ;
        RECT -4.800 3411.070 24.315 3411.370 ;
        RECT -4.800 3410.620 2.400 3411.070 ;
        RECT 23.985 3411.055 24.315 3411.070 ;
        RECT 282.965 1763.050 283.295 1763.065 ;
        RECT 282.965 1762.920 300.380 1763.050 ;
        RECT 282.965 1762.750 304.000 1762.920 ;
        RECT 282.965 1762.735 283.295 1762.750 ;
        RECT 300.000 1762.320 304.000 1762.750 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 20.310 3119.060 20.630 3119.120 ;
        RECT 24.910 3119.060 25.230 3119.120 ;
        RECT 20.310 3118.920 25.230 3119.060 ;
        RECT 20.310 3118.860 20.630 3118.920 ;
        RECT 24.910 3118.860 25.230 3118.920 ;
        RECT 24.910 1800.880 25.230 1800.940 ;
        RECT 282.970 1800.880 283.290 1800.940 ;
        RECT 24.910 1800.740 283.290 1800.880 ;
        RECT 24.910 1800.680 25.230 1800.740 ;
        RECT 282.970 1800.680 283.290 1800.740 ;
      LAYER via ;
        RECT 20.340 3118.860 20.600 3119.120 ;
        RECT 24.940 3118.860 25.200 3119.120 ;
        RECT 24.940 1800.680 25.200 1800.940 ;
        RECT 283.000 1800.680 283.260 1800.940 ;
      LAYER met2 ;
        RECT 20.330 3124.075 20.610 3124.445 ;
        RECT 20.400 3119.150 20.540 3124.075 ;
        RECT 20.340 3118.830 20.600 3119.150 ;
        RECT 24.940 3118.830 25.200 3119.150 ;
        RECT 25.000 1800.970 25.140 3118.830 ;
        RECT 24.940 1800.650 25.200 1800.970 ;
        RECT 283.000 1800.650 283.260 1800.970 ;
        RECT 283.060 1795.045 283.200 1800.650 ;
        RECT 282.990 1794.675 283.270 1795.045 ;
      LAYER via2 ;
        RECT 20.330 3124.120 20.610 3124.400 ;
        RECT 282.990 1794.720 283.270 1795.000 ;
      LAYER met3 ;
        RECT -4.800 3124.410 2.400 3124.860 ;
        RECT 20.305 3124.410 20.635 3124.425 ;
        RECT -4.800 3124.110 20.635 3124.410 ;
        RECT -4.800 3123.660 2.400 3124.110 ;
        RECT 20.305 3124.095 20.635 3124.110 ;
        RECT 282.965 1795.010 283.295 1795.025 ;
        RECT 282.965 1794.880 300.380 1795.010 ;
        RECT 282.965 1794.710 304.000 1794.880 ;
        RECT 282.965 1794.695 283.295 1794.710 ;
        RECT 300.000 1794.280 304.000 1794.710 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 1828.420 17.410 1828.480 ;
        RECT 282.970 1828.420 283.290 1828.480 ;
        RECT 17.090 1828.280 283.290 1828.420 ;
        RECT 17.090 1828.220 17.410 1828.280 ;
        RECT 282.970 1828.220 283.290 1828.280 ;
      LAYER via ;
        RECT 17.120 1828.220 17.380 1828.480 ;
        RECT 283.000 1828.220 283.260 1828.480 ;
      LAYER met2 ;
        RECT 17.110 2836.435 17.390 2836.805 ;
        RECT 17.180 1828.510 17.320 2836.435 ;
        RECT 17.120 1828.190 17.380 1828.510 ;
        RECT 283.000 1828.190 283.260 1828.510 ;
        RECT 283.060 1826.325 283.200 1828.190 ;
        RECT 282.990 1825.955 283.270 1826.325 ;
      LAYER via2 ;
        RECT 17.110 2836.480 17.390 2836.760 ;
        RECT 282.990 1826.000 283.270 1826.280 ;
      LAYER met3 ;
        RECT -4.800 2836.770 2.400 2837.220 ;
        RECT 17.085 2836.770 17.415 2836.785 ;
        RECT -4.800 2836.470 17.415 2836.770 ;
        RECT -4.800 2836.020 2.400 2836.470 ;
        RECT 17.085 2836.455 17.415 2836.470 ;
        RECT 282.965 1826.290 283.295 1826.305 ;
        RECT 282.965 1826.160 300.380 1826.290 ;
        RECT 282.965 1825.990 304.000 1826.160 ;
        RECT 282.965 1825.975 283.295 1825.990 ;
        RECT 300.000 1825.560 304.000 1825.990 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 18.470 1862.760 18.790 1862.820 ;
        RECT 282.970 1862.760 283.290 1862.820 ;
        RECT 18.470 1862.620 283.290 1862.760 ;
        RECT 18.470 1862.560 18.790 1862.620 ;
        RECT 282.970 1862.560 283.290 1862.620 ;
      LAYER via ;
        RECT 18.500 1862.560 18.760 1862.820 ;
        RECT 283.000 1862.560 283.260 1862.820 ;
      LAYER met2 ;
        RECT 18.490 2549.475 18.770 2549.845 ;
        RECT 18.560 1862.850 18.700 2549.475 ;
        RECT 18.500 1862.530 18.760 1862.850 ;
        RECT 283.000 1862.530 283.260 1862.850 ;
        RECT 283.060 1858.285 283.200 1862.530 ;
        RECT 282.990 1857.915 283.270 1858.285 ;
      LAYER via2 ;
        RECT 18.490 2549.520 18.770 2549.800 ;
        RECT 282.990 1857.960 283.270 1858.240 ;
      LAYER met3 ;
        RECT -4.800 2549.810 2.400 2550.260 ;
        RECT 18.465 2549.810 18.795 2549.825 ;
        RECT -4.800 2549.510 18.795 2549.810 ;
        RECT -4.800 2549.060 2.400 2549.510 ;
        RECT 18.465 2549.495 18.795 2549.510 ;
        RECT 282.965 1858.250 283.295 1858.265 ;
        RECT 282.965 1858.120 300.380 1858.250 ;
        RECT 282.965 1857.950 304.000 1858.120 ;
        RECT 282.965 1857.935 283.295 1857.950 ;
        RECT 300.000 1857.520 304.000 1857.950 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 19.850 1890.640 20.170 1890.700 ;
        RECT 282.970 1890.640 283.290 1890.700 ;
        RECT 19.850 1890.500 283.290 1890.640 ;
        RECT 19.850 1890.440 20.170 1890.500 ;
        RECT 282.970 1890.440 283.290 1890.500 ;
      LAYER via ;
        RECT 19.880 1890.440 20.140 1890.700 ;
        RECT 283.000 1890.440 283.260 1890.700 ;
      LAYER met2 ;
        RECT 19.870 2261.835 20.150 2262.205 ;
        RECT 19.940 1890.730 20.080 2261.835 ;
        RECT 19.880 1890.410 20.140 1890.730 ;
        RECT 283.000 1890.410 283.260 1890.730 ;
        RECT 283.060 1889.565 283.200 1890.410 ;
        RECT 282.990 1889.195 283.270 1889.565 ;
      LAYER via2 ;
        RECT 19.870 2261.880 20.150 2262.160 ;
        RECT 282.990 1889.240 283.270 1889.520 ;
      LAYER met3 ;
        RECT -4.800 2262.170 2.400 2262.620 ;
        RECT 19.845 2262.170 20.175 2262.185 ;
        RECT -4.800 2261.870 20.175 2262.170 ;
        RECT -4.800 2261.420 2.400 2261.870 ;
        RECT 19.845 2261.855 20.175 2261.870 ;
        RECT 282.965 1889.530 283.295 1889.545 ;
        RECT 282.965 1889.400 300.380 1889.530 ;
        RECT 282.965 1889.230 304.000 1889.400 ;
        RECT 282.965 1889.215 283.295 1889.230 ;
        RECT 300.000 1888.800 304.000 1889.230 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 13.870 1973.940 14.190 1974.000 ;
        RECT 26.750 1973.940 27.070 1974.000 ;
        RECT 13.870 1973.800 27.070 1973.940 ;
        RECT 13.870 1973.740 14.190 1973.800 ;
        RECT 26.750 1973.740 27.070 1973.800 ;
        RECT 110.470 1924.640 110.790 1924.700 ;
        RECT 193.270 1924.640 193.590 1924.700 ;
        RECT 110.470 1924.500 193.590 1924.640 ;
        RECT 110.470 1924.440 110.790 1924.500 ;
        RECT 193.270 1924.440 193.590 1924.500 ;
        RECT 214.430 1924.640 214.750 1924.700 ;
        RECT 214.430 1924.500 255.140 1924.640 ;
        RECT 214.430 1924.440 214.750 1924.500 ;
        RECT 26.750 1924.300 27.070 1924.360 ;
        RECT 96.670 1924.300 96.990 1924.360 ;
        RECT 26.750 1924.160 96.990 1924.300 ;
        RECT 26.750 1924.100 27.070 1924.160 ;
        RECT 96.670 1924.100 96.990 1924.160 ;
        RECT 255.000 1923.960 255.140 1924.500 ;
        RECT 282.970 1923.960 283.290 1924.020 ;
        RECT 255.000 1923.820 283.290 1923.960 ;
        RECT 282.970 1923.760 283.290 1923.820 ;
      LAYER via ;
        RECT 13.900 1973.740 14.160 1974.000 ;
        RECT 26.780 1973.740 27.040 1974.000 ;
        RECT 110.500 1924.440 110.760 1924.700 ;
        RECT 193.300 1924.440 193.560 1924.700 ;
        RECT 214.460 1924.440 214.720 1924.700 ;
        RECT 26.780 1924.100 27.040 1924.360 ;
        RECT 96.700 1924.100 96.960 1924.360 ;
        RECT 283.000 1923.760 283.260 1924.020 ;
      LAYER met2 ;
        RECT 13.890 1974.875 14.170 1975.245 ;
        RECT 13.960 1974.030 14.100 1974.875 ;
        RECT 13.900 1973.710 14.160 1974.030 ;
        RECT 26.780 1973.710 27.040 1974.030 ;
        RECT 26.840 1924.390 26.980 1973.710 ;
        RECT 110.500 1924.410 110.760 1924.730 ;
        RECT 193.290 1924.555 193.570 1924.925 ;
        RECT 214.450 1924.555 214.730 1924.925 ;
        RECT 193.300 1924.410 193.560 1924.555 ;
        RECT 214.460 1924.410 214.720 1924.555 ;
        RECT 26.780 1924.070 27.040 1924.390 ;
        RECT 96.700 1924.245 96.960 1924.390 ;
        RECT 110.560 1924.245 110.700 1924.410 ;
        RECT 96.690 1923.875 96.970 1924.245 ;
        RECT 110.490 1923.875 110.770 1924.245 ;
        RECT 283.000 1923.730 283.260 1924.050 ;
        RECT 283.060 1920.845 283.200 1923.730 ;
        RECT 282.990 1920.475 283.270 1920.845 ;
      LAYER via2 ;
        RECT 13.890 1974.920 14.170 1975.200 ;
        RECT 193.290 1924.600 193.570 1924.880 ;
        RECT 214.450 1924.600 214.730 1924.880 ;
        RECT 96.690 1923.920 96.970 1924.200 ;
        RECT 110.490 1923.920 110.770 1924.200 ;
        RECT 282.990 1920.520 283.270 1920.800 ;
      LAYER met3 ;
        RECT -4.800 1975.210 2.400 1975.660 ;
        RECT 13.865 1975.210 14.195 1975.225 ;
        RECT -4.800 1974.910 14.195 1975.210 ;
        RECT -4.800 1974.460 2.400 1974.910 ;
        RECT 13.865 1974.895 14.195 1974.910 ;
        RECT 193.265 1924.890 193.595 1924.905 ;
        RECT 214.425 1924.890 214.755 1924.905 ;
        RECT 193.265 1924.590 214.755 1924.890 ;
        RECT 193.265 1924.575 193.595 1924.590 ;
        RECT 214.425 1924.575 214.755 1924.590 ;
        RECT 96.665 1924.210 96.995 1924.225 ;
        RECT 110.465 1924.210 110.795 1924.225 ;
        RECT 96.665 1923.910 110.795 1924.210 ;
        RECT 96.665 1923.895 96.995 1923.910 ;
        RECT 110.465 1923.895 110.795 1923.910 ;
        RECT 282.965 1920.810 283.295 1920.825 ;
        RECT 282.965 1920.680 300.380 1920.810 ;
        RECT 282.965 1920.510 304.000 1920.680 ;
        RECT 282.965 1920.495 283.295 1920.510 ;
        RECT 300.000 1920.080 304.000 1920.510 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 448.110 554.100 448.430 554.160 ;
        RECT 482.610 554.100 482.930 554.160 ;
        RECT 448.110 553.960 482.930 554.100 ;
        RECT 448.110 553.900 448.430 553.960 ;
        RECT 482.610 553.900 482.930 553.960 ;
        RECT 737.910 553.420 738.230 553.480 ;
        RECT 772.410 553.420 772.730 553.480 ;
        RECT 737.910 553.280 772.730 553.420 ;
        RECT 737.910 553.220 738.230 553.280 ;
        RECT 772.410 553.220 772.730 553.280 ;
        RECT 580.130 552.740 580.450 552.800 ;
        RECT 593.930 552.740 594.250 552.800 ;
        RECT 580.130 552.600 594.250 552.740 ;
        RECT 580.130 552.540 580.450 552.600 ;
        RECT 593.930 552.540 594.250 552.600 ;
      LAYER via ;
        RECT 448.140 553.900 448.400 554.160 ;
        RECT 482.640 553.900 482.900 554.160 ;
        RECT 737.940 553.220 738.200 553.480 ;
        RECT 772.440 553.220 772.700 553.480 ;
        RECT 580.160 552.540 580.420 552.800 ;
        RECT 593.960 552.540 594.220 552.800 ;
      LAYER met2 ;
        RECT 675.830 555.035 676.110 555.405 ;
        RECT 448.140 554.045 448.400 554.190 ;
        RECT 482.640 554.045 482.900 554.190 ;
        RECT 448.130 553.675 448.410 554.045 ;
        RECT 482.630 553.675 482.910 554.045 ;
        RECT 593.950 553.675 594.230 554.045 ;
        RECT 594.020 552.830 594.160 553.675 ;
        RECT 675.900 553.365 676.040 555.035 ;
        RECT 700.210 554.355 700.490 554.725 ;
        RECT 675.830 552.995 676.110 553.365 ;
        RECT 580.160 552.685 580.420 552.830 ;
        RECT 580.150 552.315 580.430 552.685 ;
        RECT 593.960 552.510 594.220 552.830 ;
        RECT 700.280 552.685 700.420 554.355 ;
        RECT 772.430 553.675 772.710 554.045 ;
        RECT 772.500 553.510 772.640 553.675 ;
        RECT 737.940 553.365 738.200 553.510 ;
        RECT 737.930 552.995 738.210 553.365 ;
        RECT 772.440 553.190 772.700 553.510 ;
        RECT 700.210 552.315 700.490 552.685 ;
      LAYER via2 ;
        RECT 675.830 555.080 676.110 555.360 ;
        RECT 448.130 553.720 448.410 554.000 ;
        RECT 482.630 553.720 482.910 554.000 ;
        RECT 593.950 553.720 594.230 554.000 ;
        RECT 700.210 554.400 700.490 554.680 ;
        RECT 675.830 553.040 676.110 553.320 ;
        RECT 580.150 552.360 580.430 552.640 ;
        RECT 772.430 553.720 772.710 554.000 ;
        RECT 737.930 553.040 738.210 553.320 ;
        RECT 700.210 552.360 700.490 552.640 ;
      LAYER met3 ;
        RECT 284.550 1068.090 284.930 1068.100 ;
        RECT 284.550 1067.960 300.380 1068.090 ;
        RECT 284.550 1067.790 304.000 1067.960 ;
        RECT 284.550 1067.780 284.930 1067.790 ;
        RECT 300.000 1067.360 304.000 1067.790 ;
        RECT 2917.600 557.410 2924.800 557.860 ;
        RECT 2916.710 557.110 2924.800 557.410 ;
        RECT 627.710 555.370 628.090 555.380 ;
        RECT 675.805 555.370 676.135 555.385 ;
        RECT 627.710 555.070 676.135 555.370 ;
        RECT 627.710 555.060 628.090 555.070 ;
        RECT 675.805 555.055 676.135 555.070 ;
        RECT 578.950 554.690 579.330 554.700 ;
        RECT 700.185 554.690 700.515 554.705 ;
        RECT 544.030 554.390 579.330 554.690 ;
        RECT 284.550 554.010 284.930 554.020 ;
        RECT 448.105 554.010 448.435 554.025 ;
        RECT 284.550 553.710 324.450 554.010 ;
        RECT 284.550 553.700 284.930 553.710 ;
        RECT 324.150 553.330 324.450 553.710 ;
        RECT 372.910 553.710 448.435 554.010 ;
        RECT 324.150 553.030 372.290 553.330 ;
        RECT 371.990 552.650 372.290 553.030 ;
        RECT 372.910 552.650 373.210 553.710 ;
        RECT 448.105 553.695 448.435 553.710 ;
        RECT 482.605 554.010 482.935 554.025 ;
        RECT 482.605 553.710 496.490 554.010 ;
        RECT 482.605 553.695 482.935 553.710 ;
        RECT 371.990 552.350 373.210 552.650 ;
        RECT 496.190 552.650 496.490 553.710 ;
        RECT 544.030 553.330 544.330 554.390 ;
        RECT 578.950 554.380 579.330 554.390 ;
        RECT 676.510 554.390 700.515 554.690 ;
        RECT 593.925 554.010 594.255 554.025 ;
        RECT 627.710 554.010 628.090 554.020 ;
        RECT 593.925 553.710 628.090 554.010 ;
        RECT 593.925 553.695 594.255 553.710 ;
        RECT 627.710 553.700 628.090 553.710 ;
        RECT 497.110 553.030 544.330 553.330 ;
        RECT 675.805 553.330 676.135 553.345 ;
        RECT 676.510 553.330 676.810 554.390 ;
        RECT 700.185 554.375 700.515 554.390 ;
        RECT 772.405 554.010 772.735 554.025 ;
        RECT 772.405 553.710 807.450 554.010 ;
        RECT 772.405 553.695 772.735 553.710 ;
        RECT 737.905 553.330 738.235 553.345 ;
        RECT 675.805 553.030 676.810 553.330 ;
        RECT 724.350 553.030 738.235 553.330 ;
        RECT 807.150 553.330 807.450 553.710 ;
        RECT 855.910 553.710 904.050 554.010 ;
        RECT 807.150 553.030 855.290 553.330 ;
        RECT 497.110 552.650 497.410 553.030 ;
        RECT 675.805 553.015 676.135 553.030 ;
        RECT 496.190 552.350 497.410 552.650 ;
        RECT 578.950 552.650 579.330 552.660 ;
        RECT 580.125 552.650 580.455 552.665 ;
        RECT 578.950 552.350 580.455 552.650 ;
        RECT 578.950 552.340 579.330 552.350 ;
        RECT 580.125 552.335 580.455 552.350 ;
        RECT 700.185 552.650 700.515 552.665 ;
        RECT 724.350 552.650 724.650 553.030 ;
        RECT 737.905 553.015 738.235 553.030 ;
        RECT 700.185 552.350 724.650 552.650 ;
        RECT 854.990 552.650 855.290 553.030 ;
        RECT 855.910 552.650 856.210 553.710 ;
        RECT 903.750 553.330 904.050 553.710 ;
        RECT 952.510 553.710 1000.650 554.010 ;
        RECT 903.750 553.030 951.890 553.330 ;
        RECT 854.990 552.350 856.210 552.650 ;
        RECT 951.590 552.650 951.890 553.030 ;
        RECT 952.510 552.650 952.810 553.710 ;
        RECT 1000.350 553.330 1000.650 553.710 ;
        RECT 1049.110 553.710 1097.250 554.010 ;
        RECT 1000.350 553.030 1048.490 553.330 ;
        RECT 951.590 552.350 952.810 552.650 ;
        RECT 1048.190 552.650 1048.490 553.030 ;
        RECT 1049.110 552.650 1049.410 553.710 ;
        RECT 1096.950 553.330 1097.250 553.710 ;
        RECT 1145.710 553.710 1193.850 554.010 ;
        RECT 1096.950 553.030 1145.090 553.330 ;
        RECT 1048.190 552.350 1049.410 552.650 ;
        RECT 1144.790 552.650 1145.090 553.030 ;
        RECT 1145.710 552.650 1146.010 553.710 ;
        RECT 1193.550 553.330 1193.850 553.710 ;
        RECT 1242.310 553.710 1290.450 554.010 ;
        RECT 1193.550 553.030 1241.690 553.330 ;
        RECT 1144.790 552.350 1146.010 552.650 ;
        RECT 1241.390 552.650 1241.690 553.030 ;
        RECT 1242.310 552.650 1242.610 553.710 ;
        RECT 1290.150 553.330 1290.450 553.710 ;
        RECT 1338.910 553.710 1387.050 554.010 ;
        RECT 1290.150 553.030 1338.290 553.330 ;
        RECT 1241.390 552.350 1242.610 552.650 ;
        RECT 1337.990 552.650 1338.290 553.030 ;
        RECT 1338.910 552.650 1339.210 553.710 ;
        RECT 1386.750 553.330 1387.050 553.710 ;
        RECT 1435.510 553.710 1483.650 554.010 ;
        RECT 1386.750 553.030 1434.890 553.330 ;
        RECT 1337.990 552.350 1339.210 552.650 ;
        RECT 1434.590 552.650 1434.890 553.030 ;
        RECT 1435.510 552.650 1435.810 553.710 ;
        RECT 1483.350 553.330 1483.650 553.710 ;
        RECT 1532.110 553.710 1580.250 554.010 ;
        RECT 1483.350 553.030 1531.490 553.330 ;
        RECT 1434.590 552.350 1435.810 552.650 ;
        RECT 1531.190 552.650 1531.490 553.030 ;
        RECT 1532.110 552.650 1532.410 553.710 ;
        RECT 1579.950 553.330 1580.250 553.710 ;
        RECT 1628.710 553.710 1676.850 554.010 ;
        RECT 1579.950 553.030 1628.090 553.330 ;
        RECT 1531.190 552.350 1532.410 552.650 ;
        RECT 1627.790 552.650 1628.090 553.030 ;
        RECT 1628.710 552.650 1629.010 553.710 ;
        RECT 1676.550 553.330 1676.850 553.710 ;
        RECT 1725.310 553.710 1773.450 554.010 ;
        RECT 1676.550 553.030 1724.690 553.330 ;
        RECT 1627.790 552.350 1629.010 552.650 ;
        RECT 1724.390 552.650 1724.690 553.030 ;
        RECT 1725.310 552.650 1725.610 553.710 ;
        RECT 1773.150 553.330 1773.450 553.710 ;
        RECT 1821.910 553.710 1870.050 554.010 ;
        RECT 1773.150 553.030 1821.290 553.330 ;
        RECT 1724.390 552.350 1725.610 552.650 ;
        RECT 1820.990 552.650 1821.290 553.030 ;
        RECT 1821.910 552.650 1822.210 553.710 ;
        RECT 1869.750 553.330 1870.050 553.710 ;
        RECT 1918.510 553.710 1966.650 554.010 ;
        RECT 1869.750 553.030 1917.890 553.330 ;
        RECT 1820.990 552.350 1822.210 552.650 ;
        RECT 1917.590 552.650 1917.890 553.030 ;
        RECT 1918.510 552.650 1918.810 553.710 ;
        RECT 1966.350 553.330 1966.650 553.710 ;
        RECT 2015.110 553.710 2063.250 554.010 ;
        RECT 1966.350 553.030 2014.490 553.330 ;
        RECT 1917.590 552.350 1918.810 552.650 ;
        RECT 2014.190 552.650 2014.490 553.030 ;
        RECT 2015.110 552.650 2015.410 553.710 ;
        RECT 2062.950 553.330 2063.250 553.710 ;
        RECT 2111.710 553.710 2159.850 554.010 ;
        RECT 2062.950 553.030 2111.090 553.330 ;
        RECT 2014.190 552.350 2015.410 552.650 ;
        RECT 2110.790 552.650 2111.090 553.030 ;
        RECT 2111.710 552.650 2112.010 553.710 ;
        RECT 2159.550 553.330 2159.850 553.710 ;
        RECT 2208.310 553.710 2256.450 554.010 ;
        RECT 2159.550 553.030 2207.690 553.330 ;
        RECT 2110.790 552.350 2112.010 552.650 ;
        RECT 2207.390 552.650 2207.690 553.030 ;
        RECT 2208.310 552.650 2208.610 553.710 ;
        RECT 2256.150 553.330 2256.450 553.710 ;
        RECT 2304.910 553.710 2353.050 554.010 ;
        RECT 2256.150 553.030 2304.290 553.330 ;
        RECT 2207.390 552.350 2208.610 552.650 ;
        RECT 2303.990 552.650 2304.290 553.030 ;
        RECT 2304.910 552.650 2305.210 553.710 ;
        RECT 2352.750 553.330 2353.050 553.710 ;
        RECT 2401.510 553.710 2449.650 554.010 ;
        RECT 2352.750 553.030 2400.890 553.330 ;
        RECT 2303.990 552.350 2305.210 552.650 ;
        RECT 2400.590 552.650 2400.890 553.030 ;
        RECT 2401.510 552.650 2401.810 553.710 ;
        RECT 2449.350 553.330 2449.650 553.710 ;
        RECT 2498.110 553.710 2546.250 554.010 ;
        RECT 2449.350 553.030 2497.490 553.330 ;
        RECT 2400.590 552.350 2401.810 552.650 ;
        RECT 2497.190 552.650 2497.490 553.030 ;
        RECT 2498.110 552.650 2498.410 553.710 ;
        RECT 2545.950 553.330 2546.250 553.710 ;
        RECT 2594.710 553.710 2642.850 554.010 ;
        RECT 2545.950 553.030 2594.090 553.330 ;
        RECT 2497.190 552.350 2498.410 552.650 ;
        RECT 2593.790 552.650 2594.090 553.030 ;
        RECT 2594.710 552.650 2595.010 553.710 ;
        RECT 2642.550 553.330 2642.850 553.710 ;
        RECT 2691.310 553.710 2739.450 554.010 ;
        RECT 2642.550 553.030 2690.690 553.330 ;
        RECT 2593.790 552.350 2595.010 552.650 ;
        RECT 2690.390 552.650 2690.690 553.030 ;
        RECT 2691.310 552.650 2691.610 553.710 ;
        RECT 2739.150 553.330 2739.450 553.710 ;
        RECT 2787.910 553.710 2836.050 554.010 ;
        RECT 2739.150 553.030 2787.290 553.330 ;
        RECT 2690.390 552.350 2691.610 552.650 ;
        RECT 2786.990 552.650 2787.290 553.030 ;
        RECT 2787.910 552.650 2788.210 553.710 ;
        RECT 2835.750 553.330 2836.050 553.710 ;
        RECT 2916.710 553.330 2917.010 557.110 ;
        RECT 2917.600 556.660 2924.800 557.110 ;
        RECT 2835.750 553.030 2883.890 553.330 ;
        RECT 2786.990 552.350 2788.210 552.650 ;
        RECT 2883.590 552.650 2883.890 553.030 ;
        RECT 2884.510 553.030 2917.010 553.330 ;
        RECT 2884.510 552.650 2884.810 553.030 ;
        RECT 2883.590 552.350 2884.810 552.650 ;
        RECT 700.185 552.335 700.515 552.350 ;
      LAYER via3 ;
        RECT 284.580 1067.780 284.900 1068.100 ;
        RECT 627.740 555.060 628.060 555.380 ;
        RECT 284.580 553.700 284.900 554.020 ;
        RECT 578.980 554.380 579.300 554.700 ;
        RECT 627.740 553.700 628.060 554.020 ;
        RECT 578.980 552.340 579.300 552.660 ;
      LAYER met4 ;
        RECT 284.575 1067.775 284.905 1068.105 ;
        RECT 284.590 554.025 284.890 1067.775 ;
        RECT 627.735 555.055 628.065 555.385 ;
        RECT 578.975 554.375 579.305 554.705 ;
        RECT 284.575 553.695 284.905 554.025 ;
        RECT 578.990 552.665 579.290 554.375 ;
        RECT 627.750 554.025 628.050 555.055 ;
        RECT 627.735 553.695 628.065 554.025 ;
        RECT 578.975 552.335 579.305 552.665 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 16.170 1946.060 16.490 1946.120 ;
        RECT 282.970 1946.060 283.290 1946.120 ;
        RECT 16.170 1945.920 283.290 1946.060 ;
        RECT 16.170 1945.860 16.490 1945.920 ;
        RECT 282.970 1945.860 283.290 1945.920 ;
      LAYER via ;
        RECT 16.200 1945.860 16.460 1946.120 ;
        RECT 283.000 1945.860 283.260 1946.120 ;
      LAYER met2 ;
        RECT 282.990 1952.435 283.270 1952.805 ;
        RECT 283.060 1946.150 283.200 1952.435 ;
        RECT 16.200 1945.830 16.460 1946.150 ;
        RECT 283.000 1945.830 283.260 1946.150 ;
        RECT 16.260 1687.605 16.400 1945.830 ;
        RECT 16.190 1687.235 16.470 1687.605 ;
      LAYER via2 ;
        RECT 282.990 1952.480 283.270 1952.760 ;
        RECT 16.190 1687.280 16.470 1687.560 ;
      LAYER met3 ;
        RECT 282.965 1952.770 283.295 1952.785 ;
        RECT 282.965 1952.640 300.380 1952.770 ;
        RECT 282.965 1952.470 304.000 1952.640 ;
        RECT 282.965 1952.455 283.295 1952.470 ;
        RECT 300.000 1952.040 304.000 1952.470 ;
        RECT -4.800 1687.570 2.400 1688.020 ;
        RECT 16.165 1687.570 16.495 1687.585 ;
        RECT -4.800 1687.270 16.495 1687.570 ;
        RECT -4.800 1686.820 2.400 1687.270 ;
        RECT 16.165 1687.255 16.495 1687.270 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 15.250 1476.520 15.570 1476.580 ;
        RECT 283.430 1476.520 283.750 1476.580 ;
        RECT 15.250 1476.380 283.750 1476.520 ;
        RECT 15.250 1476.320 15.570 1476.380 ;
        RECT 283.430 1476.320 283.750 1476.380 ;
      LAYER via ;
        RECT 15.280 1476.320 15.540 1476.580 ;
        RECT 283.460 1476.320 283.720 1476.580 ;
      LAYER met2 ;
        RECT 283.450 1983.715 283.730 1984.085 ;
        RECT 283.520 1476.610 283.660 1983.715 ;
        RECT 15.280 1476.290 15.540 1476.610 ;
        RECT 283.460 1476.290 283.720 1476.610 ;
        RECT 15.340 1472.045 15.480 1476.290 ;
        RECT 15.270 1471.675 15.550 1472.045 ;
      LAYER via2 ;
        RECT 283.450 1983.760 283.730 1984.040 ;
        RECT 15.270 1471.720 15.550 1472.000 ;
      LAYER met3 ;
        RECT 283.425 1984.050 283.755 1984.065 ;
        RECT 283.425 1983.920 300.380 1984.050 ;
        RECT 283.425 1983.750 304.000 1983.920 ;
        RECT 283.425 1983.735 283.755 1983.750 ;
        RECT 300.000 1983.320 304.000 1983.750 ;
        RECT -4.800 1472.010 2.400 1472.460 ;
        RECT 15.245 1472.010 15.575 1472.025 ;
        RECT -4.800 1471.710 15.575 1472.010 ;
        RECT -4.800 1471.260 2.400 1471.710 ;
        RECT 15.245 1471.695 15.575 1471.710 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 1262.660 17.410 1262.720 ;
        RECT 285.730 1262.660 286.050 1262.720 ;
        RECT 17.090 1262.520 286.050 1262.660 ;
        RECT 17.090 1262.460 17.410 1262.520 ;
        RECT 285.730 1262.460 286.050 1262.520 ;
      LAYER via ;
        RECT 17.120 1262.460 17.380 1262.720 ;
        RECT 285.760 1262.460 286.020 1262.720 ;
      LAYER met2 ;
        RECT 285.750 2015.675 286.030 2016.045 ;
        RECT 285.820 1262.750 285.960 2015.675 ;
        RECT 17.120 1262.430 17.380 1262.750 ;
        RECT 285.760 1262.430 286.020 1262.750 ;
        RECT 17.180 1256.485 17.320 1262.430 ;
        RECT 17.110 1256.115 17.390 1256.485 ;
      LAYER via2 ;
        RECT 285.750 2015.720 286.030 2016.000 ;
        RECT 17.110 1256.160 17.390 1256.440 ;
      LAYER met3 ;
        RECT 285.725 2016.010 286.055 2016.025 ;
        RECT 285.725 2015.880 300.380 2016.010 ;
        RECT 285.725 2015.710 304.000 2015.880 ;
        RECT 285.725 2015.695 286.055 2015.710 ;
        RECT 300.000 2015.280 304.000 2015.710 ;
        RECT -4.800 1256.450 2.400 1256.900 ;
        RECT 17.085 1256.450 17.415 1256.465 ;
        RECT -4.800 1256.150 17.415 1256.450 ;
        RECT -4.800 1255.700 2.400 1256.150 ;
        RECT 17.085 1256.135 17.415 1256.150 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.550 2042.620 17.870 2042.680 ;
        RECT 285.730 2042.620 286.050 2042.680 ;
        RECT 17.550 2042.480 286.050 2042.620 ;
        RECT 17.550 2042.420 17.870 2042.480 ;
        RECT 285.730 2042.420 286.050 2042.480 ;
      LAYER via ;
        RECT 17.580 2042.420 17.840 2042.680 ;
        RECT 285.760 2042.420 286.020 2042.680 ;
      LAYER met2 ;
        RECT 285.750 2046.955 286.030 2047.325 ;
        RECT 285.820 2042.710 285.960 2046.955 ;
        RECT 17.580 2042.390 17.840 2042.710 ;
        RECT 285.760 2042.390 286.020 2042.710 ;
        RECT 17.640 1040.925 17.780 2042.390 ;
        RECT 17.570 1040.555 17.850 1040.925 ;
      LAYER via2 ;
        RECT 285.750 2047.000 286.030 2047.280 ;
        RECT 17.570 1040.600 17.850 1040.880 ;
      LAYER met3 ;
        RECT 285.725 2047.290 286.055 2047.305 ;
        RECT 285.725 2047.160 300.380 2047.290 ;
        RECT 285.725 2046.990 304.000 2047.160 ;
        RECT 285.725 2046.975 286.055 2046.990 ;
        RECT 300.000 2046.560 304.000 2046.990 ;
        RECT -4.800 1040.890 2.400 1041.340 ;
        RECT 17.545 1040.890 17.875 1040.905 ;
        RECT -4.800 1040.590 17.875 1040.890 ;
        RECT -4.800 1040.140 2.400 1040.590 ;
        RECT 17.545 1040.575 17.875 1040.590 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 25.370 2077.300 25.690 2077.360 ;
        RECT 285.730 2077.300 286.050 2077.360 ;
        RECT 25.370 2077.160 286.050 2077.300 ;
        RECT 25.370 2077.100 25.690 2077.160 ;
        RECT 285.730 2077.100 286.050 2077.160 ;
        RECT 13.870 827.460 14.190 827.520 ;
        RECT 25.370 827.460 25.690 827.520 ;
        RECT 13.870 827.320 25.690 827.460 ;
        RECT 13.870 827.260 14.190 827.320 ;
        RECT 25.370 827.260 25.690 827.320 ;
      LAYER via ;
        RECT 25.400 2077.100 25.660 2077.360 ;
        RECT 285.760 2077.100 286.020 2077.360 ;
        RECT 13.900 827.260 14.160 827.520 ;
        RECT 25.400 827.260 25.660 827.520 ;
      LAYER met2 ;
        RECT 285.750 2078.915 286.030 2079.285 ;
        RECT 285.820 2077.390 285.960 2078.915 ;
        RECT 25.400 2077.070 25.660 2077.390 ;
        RECT 285.760 2077.070 286.020 2077.390 ;
        RECT 25.460 827.550 25.600 2077.070 ;
        RECT 13.900 827.230 14.160 827.550 ;
        RECT 25.400 827.230 25.660 827.550 ;
        RECT 13.960 825.365 14.100 827.230 ;
        RECT 13.890 824.995 14.170 825.365 ;
      LAYER via2 ;
        RECT 285.750 2078.960 286.030 2079.240 ;
        RECT 13.890 825.040 14.170 825.320 ;
      LAYER met3 ;
        RECT 285.725 2079.250 286.055 2079.265 ;
        RECT 285.725 2079.120 300.380 2079.250 ;
        RECT 285.725 2078.950 304.000 2079.120 ;
        RECT 285.725 2078.935 286.055 2078.950 ;
        RECT 300.000 2078.520 304.000 2078.950 ;
        RECT -4.800 825.330 2.400 825.780 ;
        RECT 13.865 825.330 14.195 825.345 ;
        RECT -4.800 825.030 14.195 825.330 ;
        RECT -4.800 824.580 2.400 825.030 ;
        RECT 13.865 825.015 14.195 825.030 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 24.450 2104.840 24.770 2104.900 ;
        RECT 285.730 2104.840 286.050 2104.900 ;
        RECT 24.450 2104.700 286.050 2104.840 ;
        RECT 24.450 2104.640 24.770 2104.700 ;
        RECT 285.730 2104.640 286.050 2104.700 ;
        RECT 13.870 611.900 14.190 611.960 ;
        RECT 24.450 611.900 24.770 611.960 ;
        RECT 13.870 611.760 24.770 611.900 ;
        RECT 13.870 611.700 14.190 611.760 ;
        RECT 24.450 611.700 24.770 611.760 ;
      LAYER via ;
        RECT 24.480 2104.640 24.740 2104.900 ;
        RECT 285.760 2104.640 286.020 2104.900 ;
        RECT 13.900 611.700 14.160 611.960 ;
        RECT 24.480 611.700 24.740 611.960 ;
      LAYER met2 ;
        RECT 285.750 2110.195 286.030 2110.565 ;
        RECT 285.820 2104.930 285.960 2110.195 ;
        RECT 24.480 2104.610 24.740 2104.930 ;
        RECT 285.760 2104.610 286.020 2104.930 ;
        RECT 24.540 611.990 24.680 2104.610 ;
        RECT 13.900 611.670 14.160 611.990 ;
        RECT 24.480 611.670 24.740 611.990 ;
        RECT 13.960 610.485 14.100 611.670 ;
        RECT 13.890 610.115 14.170 610.485 ;
      LAYER via2 ;
        RECT 285.750 2110.240 286.030 2110.520 ;
        RECT 13.890 610.160 14.170 610.440 ;
      LAYER met3 ;
        RECT 285.725 2110.530 286.055 2110.545 ;
        RECT 285.725 2110.400 300.380 2110.530 ;
        RECT 285.725 2110.230 304.000 2110.400 ;
        RECT 285.725 2110.215 286.055 2110.230 ;
        RECT 300.000 2109.800 304.000 2110.230 ;
        RECT -4.800 610.450 2.400 610.900 ;
        RECT 13.865 610.450 14.195 610.465 ;
        RECT -4.800 610.150 14.195 610.450 ;
        RECT -4.800 609.700 2.400 610.150 ;
        RECT 13.865 610.135 14.195 610.150 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 51.590 2139.180 51.910 2139.240 ;
        RECT 285.730 2139.180 286.050 2139.240 ;
        RECT 51.590 2139.040 286.050 2139.180 ;
        RECT 51.590 2138.980 51.910 2139.040 ;
        RECT 285.730 2138.980 286.050 2139.040 ;
        RECT 17.090 400.080 17.410 400.140 ;
        RECT 51.590 400.080 51.910 400.140 ;
        RECT 17.090 399.940 51.910 400.080 ;
        RECT 17.090 399.880 17.410 399.940 ;
        RECT 51.590 399.880 51.910 399.940 ;
      LAYER via ;
        RECT 51.620 2138.980 51.880 2139.240 ;
        RECT 285.760 2138.980 286.020 2139.240 ;
        RECT 17.120 399.880 17.380 400.140 ;
        RECT 51.620 399.880 51.880 400.140 ;
      LAYER met2 ;
        RECT 285.750 2142.155 286.030 2142.525 ;
        RECT 285.820 2139.270 285.960 2142.155 ;
        RECT 51.620 2138.950 51.880 2139.270 ;
        RECT 285.760 2138.950 286.020 2139.270 ;
        RECT 51.680 400.170 51.820 2138.950 ;
        RECT 17.120 399.850 17.380 400.170 ;
        RECT 51.620 399.850 51.880 400.170 ;
        RECT 17.180 394.925 17.320 399.850 ;
        RECT 17.110 394.555 17.390 394.925 ;
      LAYER via2 ;
        RECT 285.750 2142.200 286.030 2142.480 ;
        RECT 17.110 394.600 17.390 394.880 ;
      LAYER met3 ;
        RECT 285.725 2142.490 286.055 2142.505 ;
        RECT 285.725 2142.360 300.380 2142.490 ;
        RECT 285.725 2142.190 304.000 2142.360 ;
        RECT 285.725 2142.175 286.055 2142.190 ;
        RECT 300.000 2141.760 304.000 2142.190 ;
        RECT -4.800 394.890 2.400 395.340 ;
        RECT 17.085 394.890 17.415 394.905 ;
        RECT -4.800 394.590 17.415 394.890 ;
        RECT -4.800 394.140 2.400 394.590 ;
        RECT 17.085 394.575 17.415 394.590 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 79.190 2173.860 79.510 2173.920 ;
        RECT 283.430 2173.860 283.750 2173.920 ;
        RECT 79.190 2173.720 283.750 2173.860 ;
        RECT 79.190 2173.660 79.510 2173.720 ;
        RECT 283.430 2173.660 283.750 2173.720 ;
        RECT 17.090 179.420 17.410 179.480 ;
        RECT 79.190 179.420 79.510 179.480 ;
        RECT 17.090 179.280 79.510 179.420 ;
        RECT 17.090 179.220 17.410 179.280 ;
        RECT 79.190 179.220 79.510 179.280 ;
      LAYER via ;
        RECT 79.220 2173.660 79.480 2173.920 ;
        RECT 283.460 2173.660 283.720 2173.920 ;
        RECT 17.120 179.220 17.380 179.480 ;
        RECT 79.220 179.220 79.480 179.480 ;
      LAYER met2 ;
        RECT 79.220 2173.630 79.480 2173.950 ;
        RECT 283.460 2173.805 283.720 2173.950 ;
        RECT 79.280 179.510 79.420 2173.630 ;
        RECT 283.450 2173.435 283.730 2173.805 ;
        RECT 17.120 179.365 17.380 179.510 ;
        RECT 17.110 178.995 17.390 179.365 ;
        RECT 79.220 179.190 79.480 179.510 ;
      LAYER via2 ;
        RECT 283.450 2173.480 283.730 2173.760 ;
        RECT 17.110 179.040 17.390 179.320 ;
      LAYER met3 ;
        RECT 283.425 2173.770 283.755 2173.785 ;
        RECT 283.425 2173.640 300.380 2173.770 ;
        RECT 283.425 2173.470 304.000 2173.640 ;
        RECT 283.425 2173.455 283.755 2173.470 ;
        RECT 300.000 2173.040 304.000 2173.470 ;
        RECT -4.800 179.330 2.400 179.780 ;
        RECT 17.085 179.330 17.415 179.345 ;
        RECT -4.800 179.030 17.415 179.330 ;
        RECT -4.800 178.580 2.400 179.030 ;
        RECT 17.085 179.015 17.415 179.030 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 283.890 793.460 284.210 793.520 ;
        RECT 2898.990 793.460 2899.310 793.520 ;
        RECT 283.890 793.320 2899.310 793.460 ;
        RECT 283.890 793.260 284.210 793.320 ;
        RECT 2898.990 793.260 2899.310 793.320 ;
      LAYER via ;
        RECT 283.920 793.260 284.180 793.520 ;
        RECT 2899.020 793.260 2899.280 793.520 ;
      LAYER met2 ;
        RECT 283.910 1099.715 284.190 1100.085 ;
        RECT 283.980 793.550 284.120 1099.715 ;
        RECT 283.920 793.230 284.180 793.550 ;
        RECT 2899.020 793.230 2899.280 793.550 ;
        RECT 2899.080 792.045 2899.220 793.230 ;
        RECT 2899.010 791.675 2899.290 792.045 ;
      LAYER via2 ;
        RECT 283.910 1099.760 284.190 1100.040 ;
        RECT 2899.010 791.720 2899.290 792.000 ;
      LAYER met3 ;
        RECT 283.885 1100.050 284.215 1100.065 ;
        RECT 283.885 1099.920 300.380 1100.050 ;
        RECT 283.885 1099.750 304.000 1099.920 ;
        RECT 283.885 1099.735 284.215 1099.750 ;
        RECT 300.000 1099.320 304.000 1099.750 ;
        RECT 2898.985 792.010 2899.315 792.025 ;
        RECT 2917.600 792.010 2924.800 792.460 ;
        RECT 2898.985 791.710 2924.800 792.010 ;
        RECT 2898.985 791.695 2899.315 791.710 ;
        RECT 2917.600 791.260 2924.800 791.710 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 287.570 1008.000 287.890 1008.060 ;
        RECT 287.200 1007.860 287.890 1008.000 ;
        RECT 285.730 1007.320 286.050 1007.380 ;
        RECT 287.200 1007.320 287.340 1007.860 ;
        RECT 287.570 1007.800 287.890 1007.860 ;
        RECT 285.730 1007.180 287.340 1007.320 ;
        RECT 285.730 1007.120 286.050 1007.180 ;
        RECT 285.730 1003.240 286.050 1003.300 ;
        RECT 2900.830 1003.240 2901.150 1003.300 ;
        RECT 285.730 1003.100 2901.150 1003.240 ;
        RECT 285.730 1003.040 286.050 1003.100 ;
        RECT 2900.830 1003.040 2901.150 1003.100 ;
      LAYER via ;
        RECT 285.760 1007.120 286.020 1007.380 ;
        RECT 287.600 1007.800 287.860 1008.060 ;
        RECT 285.760 1003.040 286.020 1003.300 ;
        RECT 2900.860 1003.040 2901.120 1003.300 ;
      LAYER met2 ;
        RECT 287.590 1130.995 287.870 1131.365 ;
        RECT 287.660 1008.090 287.800 1130.995 ;
        RECT 2900.850 1026.275 2901.130 1026.645 ;
        RECT 287.600 1007.770 287.860 1008.090 ;
        RECT 285.760 1007.090 286.020 1007.410 ;
        RECT 285.820 1003.330 285.960 1007.090 ;
        RECT 2900.920 1003.330 2901.060 1026.275 ;
        RECT 285.760 1003.010 286.020 1003.330 ;
        RECT 2900.860 1003.010 2901.120 1003.330 ;
      LAYER via2 ;
        RECT 287.590 1131.040 287.870 1131.320 ;
        RECT 2900.850 1026.320 2901.130 1026.600 ;
      LAYER met3 ;
        RECT 287.565 1131.330 287.895 1131.345 ;
        RECT 287.565 1131.200 300.380 1131.330 ;
        RECT 287.565 1131.030 304.000 1131.200 ;
        RECT 287.565 1131.015 287.895 1131.030 ;
        RECT 300.000 1130.600 304.000 1131.030 ;
        RECT 2900.825 1026.610 2901.155 1026.625 ;
        RECT 2917.600 1026.610 2924.800 1027.060 ;
        RECT 2900.825 1026.310 2924.800 1026.610 ;
        RECT 2900.825 1026.295 2901.155 1026.310 ;
        RECT 2917.600 1025.860 2924.800 1026.310 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 284.810 1027.720 285.130 1027.780 ;
        RECT 284.810 1027.580 285.960 1027.720 ;
        RECT 284.810 1027.520 285.130 1027.580 ;
        RECT 285.820 1026.080 285.960 1027.580 ;
        RECT 2899.450 1027.040 2899.770 1027.100 ;
        RECT 2900.830 1027.040 2901.150 1027.100 ;
        RECT 2899.450 1026.900 2901.150 1027.040 ;
        RECT 2899.450 1026.840 2899.770 1026.900 ;
        RECT 2900.830 1026.840 2901.150 1026.900 ;
        RECT 285.730 1025.820 286.050 1026.080 ;
        RECT 285.730 1008.000 286.050 1008.060 ;
        RECT 285.360 1007.860 286.050 1008.000 ;
        RECT 285.360 1006.980 285.500 1007.860 ;
        RECT 285.730 1007.800 286.050 1007.860 ;
        RECT 289.870 1006.980 290.190 1007.040 ;
        RECT 285.360 1006.840 290.190 1006.980 ;
        RECT 289.870 1006.780 290.190 1006.840 ;
        RECT 289.870 1002.560 290.190 1002.620 ;
        RECT 2899.450 1002.560 2899.770 1002.620 ;
        RECT 289.870 1002.420 2899.770 1002.560 ;
        RECT 289.870 1002.360 290.190 1002.420 ;
        RECT 2899.450 1002.360 2899.770 1002.420 ;
      LAYER via ;
        RECT 284.840 1027.520 285.100 1027.780 ;
        RECT 2899.480 1026.840 2899.740 1027.100 ;
        RECT 2900.860 1026.840 2901.120 1027.100 ;
        RECT 285.760 1025.820 286.020 1026.080 ;
        RECT 285.760 1007.800 286.020 1008.060 ;
        RECT 289.900 1006.780 290.160 1007.040 ;
        RECT 289.900 1002.360 290.160 1002.620 ;
        RECT 2899.480 1002.360 2899.740 1002.620 ;
      LAYER met2 ;
        RECT 2900.850 1260.875 2901.130 1261.245 ;
        RECT 284.830 1162.955 285.110 1163.325 ;
        RECT 284.900 1027.810 285.040 1162.955 ;
        RECT 284.840 1027.490 285.100 1027.810 ;
        RECT 2900.920 1027.130 2901.060 1260.875 ;
        RECT 2899.480 1026.810 2899.740 1027.130 ;
        RECT 2900.860 1026.810 2901.120 1027.130 ;
        RECT 285.760 1025.790 286.020 1026.110 ;
        RECT 285.820 1008.090 285.960 1025.790 ;
        RECT 285.760 1007.770 286.020 1008.090 ;
        RECT 289.900 1006.750 290.160 1007.070 ;
        RECT 289.960 1002.650 290.100 1006.750 ;
        RECT 2899.540 1002.650 2899.680 1026.810 ;
        RECT 289.900 1002.330 290.160 1002.650 ;
        RECT 2899.480 1002.330 2899.740 1002.650 ;
      LAYER via2 ;
        RECT 2900.850 1260.920 2901.130 1261.200 ;
        RECT 284.830 1163.000 285.110 1163.280 ;
      LAYER met3 ;
        RECT 2900.825 1261.210 2901.155 1261.225 ;
        RECT 2917.600 1261.210 2924.800 1261.660 ;
        RECT 2900.825 1260.910 2924.800 1261.210 ;
        RECT 2900.825 1260.895 2901.155 1260.910 ;
        RECT 2917.600 1260.460 2924.800 1260.910 ;
        RECT 284.805 1163.290 285.135 1163.305 ;
        RECT 284.805 1163.160 300.380 1163.290 ;
        RECT 284.805 1162.990 304.000 1163.160 ;
        RECT 284.805 1162.975 285.135 1162.990 ;
        RECT 300.000 1162.560 304.000 1162.990 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 286.190 1000.520 286.510 1000.580 ;
        RECT 2903.590 1000.520 2903.910 1000.580 ;
        RECT 286.190 1000.380 2903.910 1000.520 ;
        RECT 286.190 1000.320 286.510 1000.380 ;
        RECT 2903.590 1000.320 2903.910 1000.380 ;
      LAYER via ;
        RECT 286.220 1000.320 286.480 1000.580 ;
        RECT 2903.620 1000.320 2903.880 1000.580 ;
      LAYER met2 ;
        RECT 2903.610 1495.475 2903.890 1495.845 ;
        RECT 286.210 1194.235 286.490 1194.605 ;
        RECT 286.280 1000.610 286.420 1194.235 ;
        RECT 2903.680 1000.610 2903.820 1495.475 ;
        RECT 286.220 1000.290 286.480 1000.610 ;
        RECT 2903.620 1000.290 2903.880 1000.610 ;
      LAYER via2 ;
        RECT 2903.610 1495.520 2903.890 1495.800 ;
        RECT 286.210 1194.280 286.490 1194.560 ;
      LAYER met3 ;
        RECT 2903.585 1495.810 2903.915 1495.825 ;
        RECT 2917.600 1495.810 2924.800 1496.260 ;
        RECT 2903.585 1495.510 2924.800 1495.810 ;
        RECT 2903.585 1495.495 2903.915 1495.510 ;
        RECT 2917.600 1495.060 2924.800 1495.510 ;
        RECT 286.185 1194.570 286.515 1194.585 ;
        RECT 286.185 1194.440 300.380 1194.570 ;
        RECT 286.185 1194.270 304.000 1194.440 ;
        RECT 286.185 1194.255 286.515 1194.270 ;
        RECT 300.000 1193.840 304.000 1194.270 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 289.410 999.500 289.730 999.560 ;
        RECT 2902.210 999.500 2902.530 999.560 ;
        RECT 289.410 999.360 2902.530 999.500 ;
        RECT 289.410 999.300 289.730 999.360 ;
        RECT 2902.210 999.300 2902.530 999.360 ;
      LAYER via ;
        RECT 289.440 999.300 289.700 999.560 ;
        RECT 2902.240 999.300 2902.500 999.560 ;
      LAYER met2 ;
        RECT 2902.230 1730.075 2902.510 1730.445 ;
        RECT 289.430 1226.195 289.710 1226.565 ;
        RECT 289.500 999.590 289.640 1226.195 ;
        RECT 2902.300 999.590 2902.440 1730.075 ;
        RECT 289.440 999.270 289.700 999.590 ;
        RECT 2902.240 999.270 2902.500 999.590 ;
      LAYER via2 ;
        RECT 2902.230 1730.120 2902.510 1730.400 ;
        RECT 289.430 1226.240 289.710 1226.520 ;
      LAYER met3 ;
        RECT 2902.205 1730.410 2902.535 1730.425 ;
        RECT 2917.600 1730.410 2924.800 1730.860 ;
        RECT 2902.205 1730.110 2924.800 1730.410 ;
        RECT 2902.205 1730.095 2902.535 1730.110 ;
        RECT 2917.600 1729.660 2924.800 1730.110 ;
        RECT 289.405 1226.530 289.735 1226.545 ;
        RECT 289.405 1226.400 300.380 1226.530 ;
        RECT 289.405 1226.230 304.000 1226.400 ;
        RECT 289.405 1226.215 289.735 1226.230 ;
        RECT 300.000 1225.800 304.000 1226.230 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 287.570 2194.600 287.890 2194.660 ;
        RECT 2903.130 2194.600 2903.450 2194.660 ;
        RECT 287.570 2194.460 2903.450 2194.600 ;
        RECT 287.570 2194.400 287.890 2194.460 ;
        RECT 2903.130 2194.400 2903.450 2194.460 ;
      LAYER via ;
        RECT 287.600 2194.400 287.860 2194.660 ;
        RECT 2903.160 2194.400 2903.420 2194.660 ;
      LAYER met2 ;
        RECT 287.600 2194.370 287.860 2194.690 ;
        RECT 2903.160 2194.370 2903.420 2194.690 ;
        RECT 287.660 1257.845 287.800 2194.370 ;
        RECT 2903.220 1965.045 2903.360 2194.370 ;
        RECT 2903.150 1964.675 2903.430 1965.045 ;
        RECT 287.590 1257.475 287.870 1257.845 ;
      LAYER via2 ;
        RECT 2903.150 1964.720 2903.430 1965.000 ;
        RECT 287.590 1257.520 287.870 1257.800 ;
      LAYER met3 ;
        RECT 2903.125 1965.010 2903.455 1965.025 ;
        RECT 2917.600 1965.010 2924.800 1965.460 ;
        RECT 2903.125 1964.710 2924.800 1965.010 ;
        RECT 2903.125 1964.695 2903.455 1964.710 ;
        RECT 2917.600 1964.260 2924.800 1964.710 ;
        RECT 287.565 1257.810 287.895 1257.825 ;
        RECT 287.565 1257.680 300.380 1257.810 ;
        RECT 287.565 1257.510 304.000 1257.680 ;
        RECT 287.565 1257.495 287.895 1257.510 ;
        RECT 300.000 1257.080 304.000 1257.510 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 290.790 2194.940 291.110 2195.000 ;
        RECT 2900.370 2194.940 2900.690 2195.000 ;
        RECT 290.790 2194.800 2900.690 2194.940 ;
        RECT 290.790 2194.740 291.110 2194.800 ;
        RECT 2900.370 2194.740 2900.690 2194.800 ;
      LAYER via ;
        RECT 290.820 2194.740 291.080 2195.000 ;
        RECT 2900.400 2194.740 2900.660 2195.000 ;
      LAYER met2 ;
        RECT 2900.390 2199.275 2900.670 2199.645 ;
        RECT 2900.460 2195.030 2900.600 2199.275 ;
        RECT 290.820 2194.710 291.080 2195.030 ;
        RECT 2900.400 2194.710 2900.660 2195.030 ;
        RECT 290.880 1289.805 291.020 2194.710 ;
        RECT 290.810 1289.435 291.090 1289.805 ;
      LAYER via2 ;
        RECT 2900.390 2199.320 2900.670 2199.600 ;
        RECT 290.810 1289.480 291.090 1289.760 ;
      LAYER met3 ;
        RECT 2900.365 2199.610 2900.695 2199.625 ;
        RECT 2917.600 2199.610 2924.800 2200.060 ;
        RECT 2900.365 2199.310 2924.800 2199.610 ;
        RECT 2900.365 2199.295 2900.695 2199.310 ;
        RECT 2917.600 2198.860 2924.800 2199.310 ;
        RECT 290.785 1289.770 291.115 1289.785 ;
        RECT 290.785 1289.640 300.380 1289.770 ;
        RECT 290.785 1289.470 304.000 1289.640 ;
        RECT 290.785 1289.455 291.115 1289.470 ;
        RECT 300.000 1289.040 304.000 1289.470 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 444.430 201.860 444.750 201.920 ;
        RECT 482.610 201.860 482.930 201.920 ;
        RECT 444.430 201.720 482.930 201.860 ;
        RECT 444.430 201.660 444.750 201.720 ;
        RECT 482.610 201.660 482.930 201.720 ;
        RECT 737.910 201.180 738.230 201.240 ;
        RECT 772.410 201.180 772.730 201.240 ;
        RECT 737.910 201.040 772.730 201.180 ;
        RECT 737.910 200.980 738.230 201.040 ;
        RECT 772.410 200.980 772.730 201.040 ;
        RECT 580.130 200.500 580.450 200.560 ;
        RECT 593.930 200.500 594.250 200.560 ;
        RECT 580.130 200.360 594.250 200.500 ;
        RECT 580.130 200.300 580.450 200.360 ;
        RECT 593.930 200.300 594.250 200.360 ;
      LAYER via ;
        RECT 444.460 201.660 444.720 201.920 ;
        RECT 482.640 201.660 482.900 201.920 ;
        RECT 737.940 200.980 738.200 201.240 ;
        RECT 772.440 200.980 772.700 201.240 ;
        RECT 580.160 200.300 580.420 200.560 ;
        RECT 593.960 200.300 594.220 200.560 ;
      LAYER met2 ;
        RECT 675.830 202.795 676.110 203.165 ;
        RECT 444.460 201.805 444.720 201.950 ;
        RECT 482.640 201.805 482.900 201.950 ;
        RECT 444.450 201.435 444.730 201.805 ;
        RECT 482.630 201.435 482.910 201.805 ;
        RECT 593.950 201.435 594.230 201.805 ;
        RECT 594.020 200.590 594.160 201.435 ;
        RECT 675.900 201.125 676.040 202.795 ;
        RECT 700.210 202.115 700.490 202.485 ;
        RECT 675.830 200.755 676.110 201.125 ;
        RECT 580.160 200.445 580.420 200.590 ;
        RECT 580.150 200.075 580.430 200.445 ;
        RECT 593.960 200.270 594.220 200.590 ;
        RECT 700.280 200.445 700.420 202.115 ;
        RECT 772.430 201.435 772.710 201.805 ;
        RECT 772.500 201.270 772.640 201.435 ;
        RECT 737.940 201.125 738.200 201.270 ;
        RECT 737.930 200.755 738.210 201.125 ;
        RECT 772.440 200.950 772.700 201.270 ;
        RECT 700.210 200.075 700.490 200.445 ;
      LAYER via2 ;
        RECT 675.830 202.840 676.110 203.120 ;
        RECT 444.450 201.480 444.730 201.760 ;
        RECT 482.630 201.480 482.910 201.760 ;
        RECT 593.950 201.480 594.230 201.760 ;
        RECT 700.210 202.160 700.490 202.440 ;
        RECT 675.830 200.800 676.110 201.080 ;
        RECT 580.150 200.120 580.430 200.400 ;
        RECT 772.430 201.480 772.710 201.760 ;
        RECT 737.930 200.800 738.210 201.080 ;
        RECT 700.210 200.120 700.490 200.400 ;
      LAYER met3 ;
        RECT 288.230 1015.730 288.610 1015.740 ;
        RECT 288.230 1015.600 300.380 1015.730 ;
        RECT 288.230 1015.430 304.000 1015.600 ;
        RECT 288.230 1015.420 288.610 1015.430 ;
        RECT 300.000 1015.000 304.000 1015.430 ;
        RECT 2917.600 205.170 2924.800 205.620 ;
        RECT 2916.710 204.870 2924.800 205.170 ;
        RECT 627.710 203.130 628.090 203.140 ;
        RECT 675.805 203.130 676.135 203.145 ;
        RECT 627.710 202.830 676.135 203.130 ;
        RECT 627.710 202.820 628.090 202.830 ;
        RECT 675.805 202.815 676.135 202.830 ;
        RECT 578.950 202.450 579.330 202.460 ;
        RECT 700.185 202.450 700.515 202.465 ;
        RECT 544.030 202.150 579.330 202.450 ;
        RECT 288.230 201.770 288.610 201.780 ;
        RECT 444.425 201.770 444.755 201.785 ;
        RECT 288.230 201.470 324.450 201.770 ;
        RECT 288.230 201.460 288.610 201.470 ;
        RECT 324.150 201.090 324.450 201.470 ;
        RECT 372.910 201.470 444.755 201.770 ;
        RECT 324.150 200.790 372.290 201.090 ;
        RECT 371.990 200.410 372.290 200.790 ;
        RECT 372.910 200.410 373.210 201.470 ;
        RECT 444.425 201.455 444.755 201.470 ;
        RECT 482.605 201.770 482.935 201.785 ;
        RECT 482.605 201.470 496.490 201.770 ;
        RECT 482.605 201.455 482.935 201.470 ;
        RECT 371.990 200.110 373.210 200.410 ;
        RECT 496.190 200.410 496.490 201.470 ;
        RECT 544.030 201.090 544.330 202.150 ;
        RECT 578.950 202.140 579.330 202.150 ;
        RECT 676.510 202.150 700.515 202.450 ;
        RECT 593.925 201.770 594.255 201.785 ;
        RECT 627.710 201.770 628.090 201.780 ;
        RECT 593.925 201.470 628.090 201.770 ;
        RECT 593.925 201.455 594.255 201.470 ;
        RECT 627.710 201.460 628.090 201.470 ;
        RECT 497.110 200.790 544.330 201.090 ;
        RECT 675.805 201.090 676.135 201.105 ;
        RECT 676.510 201.090 676.810 202.150 ;
        RECT 700.185 202.135 700.515 202.150 ;
        RECT 772.405 201.770 772.735 201.785 ;
        RECT 772.405 201.470 807.450 201.770 ;
        RECT 772.405 201.455 772.735 201.470 ;
        RECT 737.905 201.090 738.235 201.105 ;
        RECT 675.805 200.790 676.810 201.090 ;
        RECT 724.350 200.790 738.235 201.090 ;
        RECT 807.150 201.090 807.450 201.470 ;
        RECT 855.910 201.470 904.050 201.770 ;
        RECT 807.150 200.790 855.290 201.090 ;
        RECT 497.110 200.410 497.410 200.790 ;
        RECT 675.805 200.775 676.135 200.790 ;
        RECT 496.190 200.110 497.410 200.410 ;
        RECT 578.950 200.410 579.330 200.420 ;
        RECT 580.125 200.410 580.455 200.425 ;
        RECT 578.950 200.110 580.455 200.410 ;
        RECT 578.950 200.100 579.330 200.110 ;
        RECT 580.125 200.095 580.455 200.110 ;
        RECT 700.185 200.410 700.515 200.425 ;
        RECT 724.350 200.410 724.650 200.790 ;
        RECT 737.905 200.775 738.235 200.790 ;
        RECT 700.185 200.110 724.650 200.410 ;
        RECT 854.990 200.410 855.290 200.790 ;
        RECT 855.910 200.410 856.210 201.470 ;
        RECT 903.750 201.090 904.050 201.470 ;
        RECT 952.510 201.470 1000.650 201.770 ;
        RECT 903.750 200.790 951.890 201.090 ;
        RECT 854.990 200.110 856.210 200.410 ;
        RECT 951.590 200.410 951.890 200.790 ;
        RECT 952.510 200.410 952.810 201.470 ;
        RECT 1000.350 201.090 1000.650 201.470 ;
        RECT 1049.110 201.470 1097.250 201.770 ;
        RECT 1000.350 200.790 1048.490 201.090 ;
        RECT 951.590 200.110 952.810 200.410 ;
        RECT 1048.190 200.410 1048.490 200.790 ;
        RECT 1049.110 200.410 1049.410 201.470 ;
        RECT 1096.950 201.090 1097.250 201.470 ;
        RECT 1145.710 201.470 1193.850 201.770 ;
        RECT 1096.950 200.790 1145.090 201.090 ;
        RECT 1048.190 200.110 1049.410 200.410 ;
        RECT 1144.790 200.410 1145.090 200.790 ;
        RECT 1145.710 200.410 1146.010 201.470 ;
        RECT 1193.550 201.090 1193.850 201.470 ;
        RECT 1242.310 201.470 1290.450 201.770 ;
        RECT 1193.550 200.790 1241.690 201.090 ;
        RECT 1144.790 200.110 1146.010 200.410 ;
        RECT 1241.390 200.410 1241.690 200.790 ;
        RECT 1242.310 200.410 1242.610 201.470 ;
        RECT 1290.150 201.090 1290.450 201.470 ;
        RECT 1338.910 201.470 1387.050 201.770 ;
        RECT 1290.150 200.790 1338.290 201.090 ;
        RECT 1241.390 200.110 1242.610 200.410 ;
        RECT 1337.990 200.410 1338.290 200.790 ;
        RECT 1338.910 200.410 1339.210 201.470 ;
        RECT 1386.750 201.090 1387.050 201.470 ;
        RECT 1435.510 201.470 1483.650 201.770 ;
        RECT 1386.750 200.790 1434.890 201.090 ;
        RECT 1337.990 200.110 1339.210 200.410 ;
        RECT 1434.590 200.410 1434.890 200.790 ;
        RECT 1435.510 200.410 1435.810 201.470 ;
        RECT 1483.350 201.090 1483.650 201.470 ;
        RECT 1532.110 201.470 1580.250 201.770 ;
        RECT 1483.350 200.790 1531.490 201.090 ;
        RECT 1434.590 200.110 1435.810 200.410 ;
        RECT 1531.190 200.410 1531.490 200.790 ;
        RECT 1532.110 200.410 1532.410 201.470 ;
        RECT 1579.950 201.090 1580.250 201.470 ;
        RECT 1628.710 201.470 1676.850 201.770 ;
        RECT 1579.950 200.790 1628.090 201.090 ;
        RECT 1531.190 200.110 1532.410 200.410 ;
        RECT 1627.790 200.410 1628.090 200.790 ;
        RECT 1628.710 200.410 1629.010 201.470 ;
        RECT 1676.550 201.090 1676.850 201.470 ;
        RECT 1725.310 201.470 1773.450 201.770 ;
        RECT 1676.550 200.790 1724.690 201.090 ;
        RECT 1627.790 200.110 1629.010 200.410 ;
        RECT 1724.390 200.410 1724.690 200.790 ;
        RECT 1725.310 200.410 1725.610 201.470 ;
        RECT 1773.150 201.090 1773.450 201.470 ;
        RECT 1821.910 201.470 1870.050 201.770 ;
        RECT 1773.150 200.790 1821.290 201.090 ;
        RECT 1724.390 200.110 1725.610 200.410 ;
        RECT 1820.990 200.410 1821.290 200.790 ;
        RECT 1821.910 200.410 1822.210 201.470 ;
        RECT 1869.750 201.090 1870.050 201.470 ;
        RECT 1918.510 201.470 1966.650 201.770 ;
        RECT 1869.750 200.790 1917.890 201.090 ;
        RECT 1820.990 200.110 1822.210 200.410 ;
        RECT 1917.590 200.410 1917.890 200.790 ;
        RECT 1918.510 200.410 1918.810 201.470 ;
        RECT 1966.350 201.090 1966.650 201.470 ;
        RECT 2015.110 201.470 2063.250 201.770 ;
        RECT 1966.350 200.790 2014.490 201.090 ;
        RECT 1917.590 200.110 1918.810 200.410 ;
        RECT 2014.190 200.410 2014.490 200.790 ;
        RECT 2015.110 200.410 2015.410 201.470 ;
        RECT 2062.950 201.090 2063.250 201.470 ;
        RECT 2111.710 201.470 2159.850 201.770 ;
        RECT 2062.950 200.790 2111.090 201.090 ;
        RECT 2014.190 200.110 2015.410 200.410 ;
        RECT 2110.790 200.410 2111.090 200.790 ;
        RECT 2111.710 200.410 2112.010 201.470 ;
        RECT 2159.550 201.090 2159.850 201.470 ;
        RECT 2208.310 201.470 2256.450 201.770 ;
        RECT 2159.550 200.790 2207.690 201.090 ;
        RECT 2110.790 200.110 2112.010 200.410 ;
        RECT 2207.390 200.410 2207.690 200.790 ;
        RECT 2208.310 200.410 2208.610 201.470 ;
        RECT 2256.150 201.090 2256.450 201.470 ;
        RECT 2304.910 201.470 2353.050 201.770 ;
        RECT 2256.150 200.790 2304.290 201.090 ;
        RECT 2207.390 200.110 2208.610 200.410 ;
        RECT 2303.990 200.410 2304.290 200.790 ;
        RECT 2304.910 200.410 2305.210 201.470 ;
        RECT 2352.750 201.090 2353.050 201.470 ;
        RECT 2401.510 201.470 2449.650 201.770 ;
        RECT 2352.750 200.790 2400.890 201.090 ;
        RECT 2303.990 200.110 2305.210 200.410 ;
        RECT 2400.590 200.410 2400.890 200.790 ;
        RECT 2401.510 200.410 2401.810 201.470 ;
        RECT 2449.350 201.090 2449.650 201.470 ;
        RECT 2498.110 201.470 2546.250 201.770 ;
        RECT 2449.350 200.790 2497.490 201.090 ;
        RECT 2400.590 200.110 2401.810 200.410 ;
        RECT 2497.190 200.410 2497.490 200.790 ;
        RECT 2498.110 200.410 2498.410 201.470 ;
        RECT 2545.950 201.090 2546.250 201.470 ;
        RECT 2594.710 201.470 2642.850 201.770 ;
        RECT 2545.950 200.790 2594.090 201.090 ;
        RECT 2497.190 200.110 2498.410 200.410 ;
        RECT 2593.790 200.410 2594.090 200.790 ;
        RECT 2594.710 200.410 2595.010 201.470 ;
        RECT 2642.550 201.090 2642.850 201.470 ;
        RECT 2691.310 201.470 2739.450 201.770 ;
        RECT 2642.550 200.790 2690.690 201.090 ;
        RECT 2593.790 200.110 2595.010 200.410 ;
        RECT 2690.390 200.410 2690.690 200.790 ;
        RECT 2691.310 200.410 2691.610 201.470 ;
        RECT 2739.150 201.090 2739.450 201.470 ;
        RECT 2787.910 201.470 2836.050 201.770 ;
        RECT 2739.150 200.790 2787.290 201.090 ;
        RECT 2690.390 200.110 2691.610 200.410 ;
        RECT 2786.990 200.410 2787.290 200.790 ;
        RECT 2787.910 200.410 2788.210 201.470 ;
        RECT 2835.750 201.090 2836.050 201.470 ;
        RECT 2916.710 201.090 2917.010 204.870 ;
        RECT 2917.600 204.420 2924.800 204.870 ;
        RECT 2835.750 200.790 2883.890 201.090 ;
        RECT 2786.990 200.110 2788.210 200.410 ;
        RECT 2883.590 200.410 2883.890 200.790 ;
        RECT 2884.510 200.790 2917.010 201.090 ;
        RECT 2884.510 200.410 2884.810 200.790 ;
        RECT 2883.590 200.110 2884.810 200.410 ;
        RECT 700.185 200.095 700.515 200.110 ;
      LAYER via3 ;
        RECT 288.260 1015.420 288.580 1015.740 ;
        RECT 627.740 202.820 628.060 203.140 ;
        RECT 288.260 201.460 288.580 201.780 ;
        RECT 578.980 202.140 579.300 202.460 ;
        RECT 627.740 201.460 628.060 201.780 ;
        RECT 578.980 200.100 579.300 200.420 ;
      LAYER met4 ;
        RECT 288.255 1015.415 288.585 1015.745 ;
        RECT 288.270 201.785 288.570 1015.415 ;
        RECT 627.735 202.815 628.065 203.145 ;
        RECT 578.975 202.135 579.305 202.465 ;
        RECT 288.255 201.455 288.585 201.785 ;
        RECT 578.990 200.425 579.290 202.135 ;
        RECT 627.750 201.785 628.050 202.815 ;
        RECT 627.735 201.455 628.065 201.785 ;
        RECT 578.975 200.095 579.305 200.425 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2902.230 2551.515 2902.510 2551.885 ;
        RECT 2902.300 2197.605 2902.440 2551.515 ;
        RECT 2902.230 2197.235 2902.510 2197.605 ;
      LAYER via2 ;
        RECT 2902.230 2551.560 2902.510 2551.840 ;
        RECT 2902.230 2197.280 2902.510 2197.560 ;
      LAYER met3 ;
        RECT 2902.205 2551.850 2902.535 2551.865 ;
        RECT 2917.600 2551.850 2924.800 2552.300 ;
        RECT 2902.205 2551.550 2924.800 2551.850 ;
        RECT 2902.205 2551.535 2902.535 2551.550 ;
        RECT 2917.600 2551.100 2924.800 2551.550 ;
        RECT 285.470 2197.570 285.850 2197.580 ;
        RECT 2902.205 2197.570 2902.535 2197.585 ;
        RECT 285.470 2197.270 2902.535 2197.570 ;
        RECT 285.470 2197.260 285.850 2197.270 ;
        RECT 2902.205 2197.255 2902.535 2197.270 ;
        RECT 285.470 1331.250 285.850 1331.260 ;
        RECT 285.470 1331.120 300.380 1331.250 ;
        RECT 285.470 1330.950 304.000 1331.120 ;
        RECT 285.470 1330.940 285.850 1330.950 ;
        RECT 300.000 1330.520 304.000 1330.950 ;
      LAYER via3 ;
        RECT 285.500 2197.260 285.820 2197.580 ;
        RECT 285.500 1330.940 285.820 1331.260 ;
      LAYER met4 ;
        RECT 285.495 2197.255 285.825 2197.585 ;
        RECT 285.510 1331.265 285.810 2197.255 ;
        RECT 285.495 1330.935 285.825 1331.265 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 291.250 2781.100 291.570 2781.160 ;
        RECT 2900.830 2781.100 2901.150 2781.160 ;
        RECT 291.250 2780.960 2901.150 2781.100 ;
        RECT 291.250 2780.900 291.570 2780.960 ;
        RECT 2900.830 2780.900 2901.150 2780.960 ;
      LAYER via ;
        RECT 291.280 2780.900 291.540 2781.160 ;
        RECT 2900.860 2780.900 2901.120 2781.160 ;
      LAYER met2 ;
        RECT 2900.850 2786.115 2901.130 2786.485 ;
        RECT 2900.920 2781.190 2901.060 2786.115 ;
        RECT 291.280 2780.870 291.540 2781.190 ;
        RECT 2900.860 2780.870 2901.120 2781.190 ;
        RECT 291.340 1363.245 291.480 2780.870 ;
        RECT 291.270 1362.875 291.550 1363.245 ;
      LAYER via2 ;
        RECT 2900.850 2786.160 2901.130 2786.440 ;
        RECT 291.270 1362.920 291.550 1363.200 ;
      LAYER met3 ;
        RECT 2900.825 2786.450 2901.155 2786.465 ;
        RECT 2917.600 2786.450 2924.800 2786.900 ;
        RECT 2900.825 2786.150 2924.800 2786.450 ;
        RECT 2900.825 2786.135 2901.155 2786.150 ;
        RECT 2917.600 2785.700 2924.800 2786.150 ;
        RECT 291.245 1363.210 291.575 1363.225 ;
        RECT 291.245 1363.080 300.380 1363.210 ;
        RECT 291.245 1362.910 304.000 1363.080 ;
        RECT 291.245 1362.895 291.575 1362.910 ;
        RECT 300.000 1362.480 304.000 1362.910 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2801.470 3017.400 2801.790 3017.460 ;
        RECT 2825.850 3017.400 2826.170 3017.460 ;
        RECT 2801.470 3017.260 2826.170 3017.400 ;
        RECT 2801.470 3017.200 2801.790 3017.260 ;
        RECT 2825.850 3017.200 2826.170 3017.260 ;
        RECT 1449.070 3016.720 1449.390 3016.780 ;
        RECT 1463.330 3016.720 1463.650 3016.780 ;
        RECT 1449.070 3016.580 1463.650 3016.720 ;
        RECT 1449.070 3016.520 1449.390 3016.580 ;
        RECT 1463.330 3016.520 1463.650 3016.580 ;
        RECT 2125.270 3016.720 2125.590 3016.780 ;
        RECT 2149.650 3016.720 2149.970 3016.780 ;
        RECT 2125.270 3016.580 2149.970 3016.720 ;
        RECT 2125.270 3016.520 2125.590 3016.580 ;
        RECT 2149.650 3016.520 2149.970 3016.580 ;
        RECT 2704.870 3016.720 2705.190 3016.780 ;
        RECT 2743.050 3016.720 2743.370 3016.780 ;
        RECT 2704.870 3016.580 2743.370 3016.720 ;
        RECT 2704.870 3016.520 2705.190 3016.580 ;
        RECT 2743.050 3016.520 2743.370 3016.580 ;
      LAYER via ;
        RECT 2801.500 3017.200 2801.760 3017.460 ;
        RECT 2825.880 3017.200 2826.140 3017.460 ;
        RECT 1449.100 3016.520 1449.360 3016.780 ;
        RECT 1463.360 3016.520 1463.620 3016.780 ;
        RECT 2125.300 3016.520 2125.560 3016.780 ;
        RECT 2149.680 3016.520 2149.940 3016.780 ;
        RECT 2704.900 3016.520 2705.160 3016.780 ;
        RECT 2743.080 3016.520 2743.340 3016.780 ;
      LAYER met2 ;
        RECT 2766.990 3017.315 2767.270 3017.685 ;
        RECT 2801.490 3017.315 2801.770 3017.685 ;
        RECT 298.630 3016.635 298.910 3017.005 ;
        RECT 1449.090 3016.635 1449.370 3017.005 ;
        RECT 298.700 2981.645 298.840 3016.635 ;
        RECT 1449.100 3016.490 1449.360 3016.635 ;
        RECT 1463.360 3016.490 1463.620 3016.810 ;
        RECT 2125.290 3016.635 2125.570 3017.005 ;
        RECT 2125.300 3016.490 2125.560 3016.635 ;
        RECT 2149.680 3016.490 2149.940 3016.810 ;
        RECT 2207.630 3016.635 2207.910 3017.005 ;
        RECT 2704.890 3016.635 2705.170 3017.005 ;
        RECT 1463.420 3015.645 1463.560 3016.490 ;
        RECT 2149.740 3016.325 2149.880 3016.490 ;
        RECT 2149.670 3015.955 2149.950 3016.325 ;
        RECT 1463.350 3015.275 1463.630 3015.645 ;
        RECT 2207.700 3014.965 2207.840 3016.635 ;
        RECT 2704.900 3016.490 2705.160 3016.635 ;
        RECT 2743.080 3016.490 2743.340 3016.810 ;
        RECT 2743.140 3015.645 2743.280 3016.490 ;
        RECT 2743.070 3015.275 2743.350 3015.645 ;
        RECT 2766.530 3015.530 2766.810 3015.645 ;
        RECT 2767.060 3015.530 2767.200 3017.315 ;
        RECT 2801.500 3017.170 2801.760 3017.315 ;
        RECT 2825.880 3017.170 2826.140 3017.490 ;
        RECT 2825.940 3017.005 2826.080 3017.170 ;
        RECT 2825.870 3016.635 2826.150 3017.005 ;
        RECT 2863.590 3016.890 2863.870 3017.005 ;
        RECT 2863.200 3016.750 2863.870 3016.890 ;
        RECT 2863.200 3016.325 2863.340 3016.750 ;
        RECT 2863.590 3016.635 2863.870 3016.750 ;
        RECT 2863.130 3015.955 2863.410 3016.325 ;
        RECT 2766.530 3015.390 2767.200 3015.530 ;
        RECT 2766.530 3015.275 2766.810 3015.390 ;
        RECT 2207.630 3014.595 2207.910 3014.965 ;
        RECT 298.630 2981.275 298.910 2981.645 ;
      LAYER via2 ;
        RECT 2766.990 3017.360 2767.270 3017.640 ;
        RECT 2801.490 3017.360 2801.770 3017.640 ;
        RECT 298.630 3016.680 298.910 3016.960 ;
        RECT 1449.090 3016.680 1449.370 3016.960 ;
        RECT 2125.290 3016.680 2125.570 3016.960 ;
        RECT 2207.630 3016.680 2207.910 3016.960 ;
        RECT 2704.890 3016.680 2705.170 3016.960 ;
        RECT 2149.670 3016.000 2149.950 3016.280 ;
        RECT 1463.350 3015.320 1463.630 3015.600 ;
        RECT 2743.070 3015.320 2743.350 3015.600 ;
        RECT 2766.530 3015.320 2766.810 3015.600 ;
        RECT 2825.870 3016.680 2826.150 3016.960 ;
        RECT 2863.590 3016.680 2863.870 3016.960 ;
        RECT 2863.130 3016.000 2863.410 3016.280 ;
        RECT 2207.630 3014.640 2207.910 3014.920 ;
        RECT 298.630 2981.320 298.910 2981.600 ;
      LAYER met3 ;
        RECT 2917.600 3021.050 2924.800 3021.500 ;
        RECT 2916.710 3020.750 2924.800 3021.050 ;
        RECT 2766.965 3017.650 2767.295 3017.665 ;
        RECT 2801.465 3017.650 2801.795 3017.665 ;
        RECT 2766.965 3017.350 2801.795 3017.650 ;
        RECT 2766.965 3017.335 2767.295 3017.350 ;
        RECT 2801.465 3017.335 2801.795 3017.350 ;
        RECT 298.605 3016.970 298.935 3016.985 ;
        RECT 1449.065 3016.970 1449.395 3016.985 ;
        RECT 298.605 3016.670 324.450 3016.970 ;
        RECT 298.605 3016.655 298.935 3016.670 ;
        RECT 324.150 3016.290 324.450 3016.670 ;
        RECT 372.910 3016.670 421.050 3016.970 ;
        RECT 324.150 3015.990 372.290 3016.290 ;
        RECT 371.990 3015.610 372.290 3015.990 ;
        RECT 372.910 3015.610 373.210 3016.670 ;
        RECT 420.750 3016.290 421.050 3016.670 ;
        RECT 469.510 3016.670 517.650 3016.970 ;
        RECT 420.750 3015.990 468.890 3016.290 ;
        RECT 371.990 3015.310 373.210 3015.610 ;
        RECT 468.590 3015.610 468.890 3015.990 ;
        RECT 469.510 3015.610 469.810 3016.670 ;
        RECT 517.350 3016.290 517.650 3016.670 ;
        RECT 566.110 3016.670 614.250 3016.970 ;
        RECT 517.350 3015.990 565.490 3016.290 ;
        RECT 468.590 3015.310 469.810 3015.610 ;
        RECT 565.190 3015.610 565.490 3015.990 ;
        RECT 566.110 3015.610 566.410 3016.670 ;
        RECT 613.950 3016.290 614.250 3016.670 ;
        RECT 662.710 3016.670 710.850 3016.970 ;
        RECT 613.950 3015.990 662.090 3016.290 ;
        RECT 565.190 3015.310 566.410 3015.610 ;
        RECT 661.790 3015.610 662.090 3015.990 ;
        RECT 662.710 3015.610 663.010 3016.670 ;
        RECT 710.550 3016.290 710.850 3016.670 ;
        RECT 759.310 3016.670 807.450 3016.970 ;
        RECT 710.550 3015.990 758.690 3016.290 ;
        RECT 661.790 3015.310 663.010 3015.610 ;
        RECT 758.390 3015.610 758.690 3015.990 ;
        RECT 759.310 3015.610 759.610 3016.670 ;
        RECT 807.150 3016.290 807.450 3016.670 ;
        RECT 855.910 3016.670 904.050 3016.970 ;
        RECT 807.150 3015.990 855.290 3016.290 ;
        RECT 758.390 3015.310 759.610 3015.610 ;
        RECT 854.990 3015.610 855.290 3015.990 ;
        RECT 855.910 3015.610 856.210 3016.670 ;
        RECT 903.750 3016.290 904.050 3016.670 ;
        RECT 952.510 3016.670 1000.650 3016.970 ;
        RECT 903.750 3015.990 951.890 3016.290 ;
        RECT 854.990 3015.310 856.210 3015.610 ;
        RECT 951.590 3015.610 951.890 3015.990 ;
        RECT 952.510 3015.610 952.810 3016.670 ;
        RECT 1000.350 3016.290 1000.650 3016.670 ;
        RECT 1049.110 3016.670 1097.250 3016.970 ;
        RECT 1000.350 3015.990 1048.490 3016.290 ;
        RECT 951.590 3015.310 952.810 3015.610 ;
        RECT 1048.190 3015.610 1048.490 3015.990 ;
        RECT 1049.110 3015.610 1049.410 3016.670 ;
        RECT 1096.950 3016.290 1097.250 3016.670 ;
        RECT 1145.710 3016.670 1193.850 3016.970 ;
        RECT 1096.950 3015.990 1145.090 3016.290 ;
        RECT 1048.190 3015.310 1049.410 3015.610 ;
        RECT 1144.790 3015.610 1145.090 3015.990 ;
        RECT 1145.710 3015.610 1146.010 3016.670 ;
        RECT 1193.550 3016.290 1193.850 3016.670 ;
        RECT 1242.310 3016.670 1290.450 3016.970 ;
        RECT 1193.550 3015.990 1241.690 3016.290 ;
        RECT 1144.790 3015.310 1146.010 3015.610 ;
        RECT 1241.390 3015.610 1241.690 3015.990 ;
        RECT 1242.310 3015.610 1242.610 3016.670 ;
        RECT 1290.150 3016.290 1290.450 3016.670 ;
        RECT 1338.910 3016.670 1387.050 3016.970 ;
        RECT 1290.150 3015.990 1338.290 3016.290 ;
        RECT 1241.390 3015.310 1242.610 3015.610 ;
        RECT 1337.990 3015.610 1338.290 3015.990 ;
        RECT 1338.910 3015.610 1339.210 3016.670 ;
        RECT 1386.750 3016.290 1387.050 3016.670 ;
        RECT 1435.510 3016.670 1449.395 3016.970 ;
        RECT 1386.750 3015.990 1434.890 3016.290 ;
        RECT 1337.990 3015.310 1339.210 3015.610 ;
        RECT 1434.590 3015.610 1434.890 3015.990 ;
        RECT 1435.510 3015.610 1435.810 3016.670 ;
        RECT 1449.065 3016.655 1449.395 3016.670 ;
        RECT 1497.110 3016.970 1497.490 3016.980 ;
        RECT 2125.265 3016.970 2125.595 3016.985 ;
        RECT 1497.110 3016.670 1580.250 3016.970 ;
        RECT 1497.110 3016.660 1497.490 3016.670 ;
        RECT 1579.950 3016.290 1580.250 3016.670 ;
        RECT 1628.710 3016.670 1676.850 3016.970 ;
        RECT 1579.950 3015.990 1628.090 3016.290 ;
        RECT 1434.590 3015.310 1435.810 3015.610 ;
        RECT 1463.325 3015.610 1463.655 3015.625 ;
        RECT 1497.110 3015.610 1497.490 3015.620 ;
        RECT 1463.325 3015.310 1497.490 3015.610 ;
        RECT 1627.790 3015.610 1628.090 3015.990 ;
        RECT 1628.710 3015.610 1629.010 3016.670 ;
        RECT 1676.550 3016.290 1676.850 3016.670 ;
        RECT 1725.310 3016.670 1773.450 3016.970 ;
        RECT 1676.550 3015.990 1724.690 3016.290 ;
        RECT 1627.790 3015.310 1629.010 3015.610 ;
        RECT 1724.390 3015.610 1724.690 3015.990 ;
        RECT 1725.310 3015.610 1725.610 3016.670 ;
        RECT 1773.150 3016.290 1773.450 3016.670 ;
        RECT 1821.910 3016.670 1870.050 3016.970 ;
        RECT 1773.150 3015.990 1821.290 3016.290 ;
        RECT 1724.390 3015.310 1725.610 3015.610 ;
        RECT 1820.990 3015.610 1821.290 3015.990 ;
        RECT 1821.910 3015.610 1822.210 3016.670 ;
        RECT 1869.750 3016.290 1870.050 3016.670 ;
        RECT 1918.510 3016.670 1966.650 3016.970 ;
        RECT 1869.750 3015.990 1917.890 3016.290 ;
        RECT 1820.990 3015.310 1822.210 3015.610 ;
        RECT 1917.590 3015.610 1917.890 3015.990 ;
        RECT 1918.510 3015.610 1918.810 3016.670 ;
        RECT 1966.350 3016.290 1966.650 3016.670 ;
        RECT 2015.110 3016.670 2125.595 3016.970 ;
        RECT 1966.350 3015.990 2014.490 3016.290 ;
        RECT 1917.590 3015.310 1918.810 3015.610 ;
        RECT 2014.190 3015.610 2014.490 3015.990 ;
        RECT 2015.110 3015.610 2015.410 3016.670 ;
        RECT 2125.265 3016.655 2125.595 3016.670 ;
        RECT 2207.605 3016.970 2207.935 3016.985 ;
        RECT 2704.865 3016.970 2705.195 3016.985 ;
        RECT 2207.605 3016.670 2256.450 3016.970 ;
        RECT 2207.605 3016.655 2207.935 3016.670 ;
        RECT 2149.645 3016.290 2149.975 3016.305 ;
        RECT 2173.310 3016.290 2173.690 3016.300 ;
        RECT 2149.645 3015.990 2173.690 3016.290 ;
        RECT 2256.150 3016.290 2256.450 3016.670 ;
        RECT 2304.910 3016.670 2353.050 3016.970 ;
        RECT 2256.150 3015.990 2304.290 3016.290 ;
        RECT 2149.645 3015.975 2149.975 3015.990 ;
        RECT 2173.310 3015.980 2173.690 3015.990 ;
        RECT 2014.190 3015.310 2015.410 3015.610 ;
        RECT 2303.990 3015.610 2304.290 3015.990 ;
        RECT 2304.910 3015.610 2305.210 3016.670 ;
        RECT 2352.750 3016.290 2353.050 3016.670 ;
        RECT 2401.510 3016.670 2449.650 3016.970 ;
        RECT 2352.750 3015.990 2400.890 3016.290 ;
        RECT 2303.990 3015.310 2305.210 3015.610 ;
        RECT 2400.590 3015.610 2400.890 3015.990 ;
        RECT 2401.510 3015.610 2401.810 3016.670 ;
        RECT 2449.350 3016.290 2449.650 3016.670 ;
        RECT 2498.110 3016.670 2546.250 3016.970 ;
        RECT 2449.350 3015.990 2497.490 3016.290 ;
        RECT 2400.590 3015.310 2401.810 3015.610 ;
        RECT 2497.190 3015.610 2497.490 3015.990 ;
        RECT 2498.110 3015.610 2498.410 3016.670 ;
        RECT 2545.950 3016.290 2546.250 3016.670 ;
        RECT 2594.710 3016.670 2642.850 3016.970 ;
        RECT 2545.950 3015.990 2594.090 3016.290 ;
        RECT 2497.190 3015.310 2498.410 3015.610 ;
        RECT 2593.790 3015.610 2594.090 3015.990 ;
        RECT 2594.710 3015.610 2595.010 3016.670 ;
        RECT 2642.550 3016.290 2642.850 3016.670 ;
        RECT 2691.310 3016.670 2705.195 3016.970 ;
        RECT 2642.550 3015.990 2690.690 3016.290 ;
        RECT 2593.790 3015.310 2595.010 3015.610 ;
        RECT 2690.390 3015.610 2690.690 3015.990 ;
        RECT 2691.310 3015.610 2691.610 3016.670 ;
        RECT 2704.865 3016.655 2705.195 3016.670 ;
        RECT 2825.845 3016.970 2826.175 3016.985 ;
        RECT 2863.565 3016.970 2863.895 3016.985 ;
        RECT 2825.845 3016.670 2849.850 3016.970 ;
        RECT 2825.845 3016.655 2826.175 3016.670 ;
        RECT 2849.550 3016.290 2849.850 3016.670 ;
        RECT 2863.565 3016.670 2884.810 3016.970 ;
        RECT 2863.565 3016.655 2863.895 3016.670 ;
        RECT 2863.105 3016.290 2863.435 3016.305 ;
        RECT 2849.550 3015.990 2863.435 3016.290 ;
        RECT 2884.510 3016.290 2884.810 3016.670 ;
        RECT 2916.710 3016.290 2917.010 3020.750 ;
        RECT 2917.600 3020.300 2924.800 3020.750 ;
        RECT 2884.510 3015.990 2917.010 3016.290 ;
        RECT 2863.105 3015.975 2863.435 3015.990 ;
        RECT 2690.390 3015.310 2691.610 3015.610 ;
        RECT 2743.045 3015.610 2743.375 3015.625 ;
        RECT 2766.505 3015.610 2766.835 3015.625 ;
        RECT 2743.045 3015.310 2766.835 3015.610 ;
        RECT 1463.325 3015.295 1463.655 3015.310 ;
        RECT 1497.110 3015.300 1497.490 3015.310 ;
        RECT 2743.045 3015.295 2743.375 3015.310 ;
        RECT 2766.505 3015.295 2766.835 3015.310 ;
        RECT 2173.310 3014.930 2173.690 3014.940 ;
        RECT 2207.605 3014.930 2207.935 3014.945 ;
        RECT 2173.310 3014.630 2207.935 3014.930 ;
        RECT 2173.310 3014.620 2173.690 3014.630 ;
        RECT 2207.605 3014.615 2207.935 3014.630 ;
        RECT 298.605 2981.610 298.935 2981.625 ;
        RECT 295.630 2981.310 298.935 2981.610 ;
        RECT 295.630 2980.930 295.930 2981.310 ;
        RECT 298.605 2981.295 298.935 2981.310 ;
        RECT 297.430 2980.930 297.810 2980.940 ;
        RECT 295.630 2980.630 297.810 2980.930 ;
        RECT 297.430 2980.620 297.810 2980.630 ;
        RECT 294.670 1394.490 295.050 1394.500 ;
        RECT 294.670 1394.360 300.380 1394.490 ;
        RECT 294.670 1394.190 304.000 1394.360 ;
        RECT 294.670 1394.180 295.050 1394.190 ;
        RECT 300.000 1393.760 304.000 1394.190 ;
      LAYER via3 ;
        RECT 1497.140 3016.660 1497.460 3016.980 ;
        RECT 1497.140 3015.300 1497.460 3015.620 ;
        RECT 2173.340 3015.980 2173.660 3016.300 ;
        RECT 2173.340 3014.620 2173.660 3014.940 ;
        RECT 297.460 2980.620 297.780 2980.940 ;
        RECT 294.700 1394.180 295.020 1394.500 ;
      LAYER met4 ;
        RECT 1497.135 3016.655 1497.465 3016.985 ;
        RECT 1497.150 3015.625 1497.450 3016.655 ;
        RECT 2173.335 3015.975 2173.665 3016.305 ;
        RECT 1497.135 3015.295 1497.465 3015.625 ;
        RECT 2173.350 3014.945 2173.650 3015.975 ;
        RECT 2173.335 3014.615 2173.665 3014.945 ;
        RECT 297.455 2980.615 297.785 2980.945 ;
        RECT 297.470 2888.450 297.770 2980.615 ;
        RECT 296.550 2888.150 297.770 2888.450 ;
        RECT 296.550 2864.650 296.850 2888.150 ;
        RECT 295.630 2864.350 296.850 2864.650 ;
        RECT 295.630 2766.050 295.930 2864.350 ;
        RECT 294.710 2765.750 295.930 2766.050 ;
        RECT 294.710 2286.650 295.010 2765.750 ;
        RECT 294.710 2286.350 295.930 2286.650 ;
        RECT 295.630 2198.250 295.930 2286.350 ;
        RECT 294.710 2197.950 295.930 2198.250 ;
        RECT 294.710 1394.505 295.010 2197.950 ;
        RECT 294.695 1394.175 295.025 1394.505 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2801.470 3252.000 2801.790 3252.060 ;
        RECT 2825.850 3252.000 2826.170 3252.060 ;
        RECT 2801.470 3251.860 2826.170 3252.000 ;
        RECT 2801.470 3251.800 2801.790 3251.860 ;
        RECT 2825.850 3251.800 2826.170 3251.860 ;
        RECT 2125.270 3251.320 2125.590 3251.380 ;
        RECT 2172.650 3251.320 2172.970 3251.380 ;
        RECT 2125.270 3251.180 2172.970 3251.320 ;
        RECT 2125.270 3251.120 2125.590 3251.180 ;
        RECT 2172.650 3251.120 2172.970 3251.180 ;
        RECT 2704.870 3251.320 2705.190 3251.380 ;
        RECT 2743.050 3251.320 2743.370 3251.380 ;
        RECT 2704.870 3251.180 2743.370 3251.320 ;
        RECT 2704.870 3251.120 2705.190 3251.180 ;
        RECT 2743.050 3251.120 2743.370 3251.180 ;
      LAYER via ;
        RECT 2801.500 3251.800 2801.760 3252.060 ;
        RECT 2825.880 3251.800 2826.140 3252.060 ;
        RECT 2125.300 3251.120 2125.560 3251.380 ;
        RECT 2172.680 3251.120 2172.940 3251.380 ;
        RECT 2704.900 3251.120 2705.160 3251.380 ;
        RECT 2743.080 3251.120 2743.340 3251.380 ;
      LAYER met2 ;
        RECT 2766.530 3252.170 2766.810 3252.285 ;
        RECT 2767.450 3252.170 2767.730 3252.285 ;
        RECT 2766.530 3252.030 2767.730 3252.170 ;
        RECT 2766.530 3251.915 2766.810 3252.030 ;
        RECT 2767.450 3251.915 2767.730 3252.030 ;
        RECT 2801.490 3251.915 2801.770 3252.285 ;
        RECT 2801.500 3251.770 2801.760 3251.915 ;
        RECT 2825.880 3251.770 2826.140 3252.090 ;
        RECT 2825.940 3251.605 2826.080 3251.770 ;
        RECT 2125.290 3251.235 2125.570 3251.605 ;
        RECT 2125.300 3251.090 2125.560 3251.235 ;
        RECT 2172.680 3251.090 2172.940 3251.410 ;
        RECT 2704.890 3251.235 2705.170 3251.605 ;
        RECT 2704.900 3251.090 2705.160 3251.235 ;
        RECT 2743.080 3251.090 2743.340 3251.410 ;
        RECT 2825.870 3251.235 2826.150 3251.605 ;
        RECT 2863.590 3251.490 2863.870 3251.605 ;
        RECT 2863.200 3251.350 2863.870 3251.490 ;
        RECT 2172.740 3250.925 2172.880 3251.090 ;
        RECT 2172.670 3250.555 2172.950 3250.925 ;
        RECT 2743.140 3250.245 2743.280 3251.090 ;
        RECT 2863.200 3250.925 2863.340 3251.350 ;
        RECT 2863.590 3251.235 2863.870 3251.350 ;
        RECT 2863.130 3250.555 2863.410 3250.925 ;
        RECT 2743.070 3249.875 2743.350 3250.245 ;
      LAYER via2 ;
        RECT 2766.530 3251.960 2766.810 3252.240 ;
        RECT 2767.450 3251.960 2767.730 3252.240 ;
        RECT 2801.490 3251.960 2801.770 3252.240 ;
        RECT 2125.290 3251.280 2125.570 3251.560 ;
        RECT 2704.890 3251.280 2705.170 3251.560 ;
        RECT 2825.870 3251.280 2826.150 3251.560 ;
        RECT 2172.670 3250.600 2172.950 3250.880 ;
        RECT 2863.590 3251.280 2863.870 3251.560 ;
        RECT 2863.130 3250.600 2863.410 3250.880 ;
        RECT 2743.070 3249.920 2743.350 3250.200 ;
      LAYER met3 ;
        RECT 2917.600 3255.650 2924.800 3256.100 ;
        RECT 2916.710 3255.350 2924.800 3255.650 ;
        RECT 2752.910 3252.250 2753.290 3252.260 ;
        RECT 2766.505 3252.250 2766.835 3252.265 ;
        RECT 2752.910 3251.950 2766.835 3252.250 ;
        RECT 2752.910 3251.940 2753.290 3251.950 ;
        RECT 2766.505 3251.935 2766.835 3251.950 ;
        RECT 2767.425 3252.250 2767.755 3252.265 ;
        RECT 2801.465 3252.250 2801.795 3252.265 ;
        RECT 2767.425 3251.950 2801.795 3252.250 ;
        RECT 2767.425 3251.935 2767.755 3251.950 ;
        RECT 2801.465 3251.935 2801.795 3251.950 ;
        RECT 290.990 3251.570 291.370 3251.580 ;
        RECT 1497.110 3251.570 1497.490 3251.580 ;
        RECT 2125.265 3251.570 2125.595 3251.585 ;
        RECT 2704.865 3251.570 2705.195 3251.585 ;
        RECT 290.990 3251.270 324.450 3251.570 ;
        RECT 290.990 3251.260 291.370 3251.270 ;
        RECT 324.150 3250.890 324.450 3251.270 ;
        RECT 372.910 3251.270 421.050 3251.570 ;
        RECT 324.150 3250.590 372.290 3250.890 ;
        RECT 371.990 3250.210 372.290 3250.590 ;
        RECT 372.910 3250.210 373.210 3251.270 ;
        RECT 420.750 3250.890 421.050 3251.270 ;
        RECT 469.510 3251.270 517.650 3251.570 ;
        RECT 420.750 3250.590 468.890 3250.890 ;
        RECT 371.990 3249.910 373.210 3250.210 ;
        RECT 468.590 3250.210 468.890 3250.590 ;
        RECT 469.510 3250.210 469.810 3251.270 ;
        RECT 517.350 3250.890 517.650 3251.270 ;
        RECT 566.110 3251.270 614.250 3251.570 ;
        RECT 517.350 3250.590 565.490 3250.890 ;
        RECT 468.590 3249.910 469.810 3250.210 ;
        RECT 565.190 3250.210 565.490 3250.590 ;
        RECT 566.110 3250.210 566.410 3251.270 ;
        RECT 613.950 3250.890 614.250 3251.270 ;
        RECT 662.710 3251.270 710.850 3251.570 ;
        RECT 613.950 3250.590 662.090 3250.890 ;
        RECT 565.190 3249.910 566.410 3250.210 ;
        RECT 661.790 3250.210 662.090 3250.590 ;
        RECT 662.710 3250.210 663.010 3251.270 ;
        RECT 710.550 3250.890 710.850 3251.270 ;
        RECT 759.310 3251.270 807.450 3251.570 ;
        RECT 710.550 3250.590 758.690 3250.890 ;
        RECT 661.790 3249.910 663.010 3250.210 ;
        RECT 758.390 3250.210 758.690 3250.590 ;
        RECT 759.310 3250.210 759.610 3251.270 ;
        RECT 807.150 3250.890 807.450 3251.270 ;
        RECT 855.910 3251.270 904.050 3251.570 ;
        RECT 807.150 3250.590 855.290 3250.890 ;
        RECT 758.390 3249.910 759.610 3250.210 ;
        RECT 854.990 3250.210 855.290 3250.590 ;
        RECT 855.910 3250.210 856.210 3251.270 ;
        RECT 903.750 3250.890 904.050 3251.270 ;
        RECT 952.510 3251.270 1000.650 3251.570 ;
        RECT 903.750 3250.590 951.890 3250.890 ;
        RECT 854.990 3249.910 856.210 3250.210 ;
        RECT 951.590 3250.210 951.890 3250.590 ;
        RECT 952.510 3250.210 952.810 3251.270 ;
        RECT 1000.350 3250.890 1000.650 3251.270 ;
        RECT 1049.110 3251.270 1097.250 3251.570 ;
        RECT 1000.350 3250.590 1048.490 3250.890 ;
        RECT 951.590 3249.910 952.810 3250.210 ;
        RECT 1048.190 3250.210 1048.490 3250.590 ;
        RECT 1049.110 3250.210 1049.410 3251.270 ;
        RECT 1096.950 3250.890 1097.250 3251.270 ;
        RECT 1145.710 3251.270 1193.850 3251.570 ;
        RECT 1096.950 3250.590 1145.090 3250.890 ;
        RECT 1048.190 3249.910 1049.410 3250.210 ;
        RECT 1144.790 3250.210 1145.090 3250.590 ;
        RECT 1145.710 3250.210 1146.010 3251.270 ;
        RECT 1193.550 3250.890 1193.850 3251.270 ;
        RECT 1242.310 3251.270 1290.450 3251.570 ;
        RECT 1193.550 3250.590 1241.690 3250.890 ;
        RECT 1144.790 3249.910 1146.010 3250.210 ;
        RECT 1241.390 3250.210 1241.690 3250.590 ;
        RECT 1242.310 3250.210 1242.610 3251.270 ;
        RECT 1290.150 3250.890 1290.450 3251.270 ;
        RECT 1338.910 3251.270 1387.050 3251.570 ;
        RECT 1290.150 3250.590 1338.290 3250.890 ;
        RECT 1241.390 3249.910 1242.610 3250.210 ;
        RECT 1337.990 3250.210 1338.290 3250.590 ;
        RECT 1338.910 3250.210 1339.210 3251.270 ;
        RECT 1386.750 3250.890 1387.050 3251.270 ;
        RECT 1435.510 3251.270 1463.410 3251.570 ;
        RECT 1386.750 3250.590 1434.890 3250.890 ;
        RECT 1337.990 3249.910 1339.210 3250.210 ;
        RECT 1434.590 3250.210 1434.890 3250.590 ;
        RECT 1435.510 3250.210 1435.810 3251.270 ;
        RECT 1434.590 3249.910 1435.810 3250.210 ;
        RECT 1463.110 3250.210 1463.410 3251.270 ;
        RECT 1497.110 3251.270 1580.250 3251.570 ;
        RECT 1497.110 3251.260 1497.490 3251.270 ;
        RECT 1579.950 3250.890 1580.250 3251.270 ;
        RECT 1628.710 3251.270 1676.850 3251.570 ;
        RECT 1579.950 3250.590 1628.090 3250.890 ;
        RECT 1497.110 3250.210 1497.490 3250.220 ;
        RECT 1463.110 3249.910 1497.490 3250.210 ;
        RECT 1627.790 3250.210 1628.090 3250.590 ;
        RECT 1628.710 3250.210 1629.010 3251.270 ;
        RECT 1676.550 3250.890 1676.850 3251.270 ;
        RECT 1725.310 3251.270 1773.450 3251.570 ;
        RECT 1676.550 3250.590 1724.690 3250.890 ;
        RECT 1627.790 3249.910 1629.010 3250.210 ;
        RECT 1724.390 3250.210 1724.690 3250.590 ;
        RECT 1725.310 3250.210 1725.610 3251.270 ;
        RECT 1773.150 3250.890 1773.450 3251.270 ;
        RECT 1821.910 3251.270 1870.050 3251.570 ;
        RECT 1773.150 3250.590 1821.290 3250.890 ;
        RECT 1724.390 3249.910 1725.610 3250.210 ;
        RECT 1820.990 3250.210 1821.290 3250.590 ;
        RECT 1821.910 3250.210 1822.210 3251.270 ;
        RECT 1869.750 3250.890 1870.050 3251.270 ;
        RECT 1918.510 3251.270 1966.650 3251.570 ;
        RECT 1869.750 3250.590 1917.890 3250.890 ;
        RECT 1820.990 3249.910 1822.210 3250.210 ;
        RECT 1917.590 3250.210 1917.890 3250.590 ;
        RECT 1918.510 3250.210 1918.810 3251.270 ;
        RECT 1966.350 3250.890 1966.650 3251.270 ;
        RECT 2015.110 3251.270 2063.250 3251.570 ;
        RECT 1966.350 3250.590 2014.490 3250.890 ;
        RECT 1917.590 3249.910 1918.810 3250.210 ;
        RECT 2014.190 3250.210 2014.490 3250.590 ;
        RECT 2015.110 3250.210 2015.410 3251.270 ;
        RECT 2062.950 3250.890 2063.250 3251.270 ;
        RECT 2111.710 3251.270 2125.595 3251.570 ;
        RECT 2062.950 3250.590 2111.090 3250.890 ;
        RECT 2014.190 3249.910 2015.410 3250.210 ;
        RECT 2110.790 3250.210 2111.090 3250.590 ;
        RECT 2111.710 3250.210 2112.010 3251.270 ;
        RECT 2125.265 3251.255 2125.595 3251.270 ;
        RECT 2186.230 3251.270 2256.450 3251.570 ;
        RECT 2172.645 3250.890 2172.975 3250.905 ;
        RECT 2186.230 3250.890 2186.530 3251.270 ;
        RECT 2172.645 3250.590 2186.530 3250.890 ;
        RECT 2256.150 3250.890 2256.450 3251.270 ;
        RECT 2304.910 3251.270 2353.050 3251.570 ;
        RECT 2256.150 3250.590 2304.290 3250.890 ;
        RECT 2172.645 3250.575 2172.975 3250.590 ;
        RECT 2110.790 3249.910 2112.010 3250.210 ;
        RECT 2303.990 3250.210 2304.290 3250.590 ;
        RECT 2304.910 3250.210 2305.210 3251.270 ;
        RECT 2352.750 3250.890 2353.050 3251.270 ;
        RECT 2401.510 3251.270 2449.650 3251.570 ;
        RECT 2352.750 3250.590 2400.890 3250.890 ;
        RECT 2303.990 3249.910 2305.210 3250.210 ;
        RECT 2400.590 3250.210 2400.890 3250.590 ;
        RECT 2401.510 3250.210 2401.810 3251.270 ;
        RECT 2449.350 3250.890 2449.650 3251.270 ;
        RECT 2498.110 3251.270 2546.250 3251.570 ;
        RECT 2449.350 3250.590 2497.490 3250.890 ;
        RECT 2400.590 3249.910 2401.810 3250.210 ;
        RECT 2497.190 3250.210 2497.490 3250.590 ;
        RECT 2498.110 3250.210 2498.410 3251.270 ;
        RECT 2545.950 3250.890 2546.250 3251.270 ;
        RECT 2594.710 3251.270 2642.850 3251.570 ;
        RECT 2545.950 3250.590 2594.090 3250.890 ;
        RECT 2497.190 3249.910 2498.410 3250.210 ;
        RECT 2593.790 3250.210 2594.090 3250.590 ;
        RECT 2594.710 3250.210 2595.010 3251.270 ;
        RECT 2642.550 3250.890 2642.850 3251.270 ;
        RECT 2691.310 3251.270 2705.195 3251.570 ;
        RECT 2642.550 3250.590 2690.690 3250.890 ;
        RECT 2593.790 3249.910 2595.010 3250.210 ;
        RECT 2690.390 3250.210 2690.690 3250.590 ;
        RECT 2691.310 3250.210 2691.610 3251.270 ;
        RECT 2704.865 3251.255 2705.195 3251.270 ;
        RECT 2825.845 3251.570 2826.175 3251.585 ;
        RECT 2863.565 3251.570 2863.895 3251.585 ;
        RECT 2825.845 3251.270 2849.850 3251.570 ;
        RECT 2825.845 3251.255 2826.175 3251.270 ;
        RECT 2849.550 3250.890 2849.850 3251.270 ;
        RECT 2863.565 3251.270 2884.810 3251.570 ;
        RECT 2863.565 3251.255 2863.895 3251.270 ;
        RECT 2863.105 3250.890 2863.435 3250.905 ;
        RECT 2849.550 3250.590 2863.435 3250.890 ;
        RECT 2884.510 3250.890 2884.810 3251.270 ;
        RECT 2916.710 3250.890 2917.010 3255.350 ;
        RECT 2917.600 3254.900 2924.800 3255.350 ;
        RECT 2884.510 3250.590 2917.010 3250.890 ;
        RECT 2863.105 3250.575 2863.435 3250.590 ;
        RECT 2690.390 3249.910 2691.610 3250.210 ;
        RECT 2743.045 3250.210 2743.375 3250.225 ;
        RECT 2752.910 3250.210 2753.290 3250.220 ;
        RECT 2743.045 3249.910 2753.290 3250.210 ;
        RECT 1497.110 3249.900 1497.490 3249.910 ;
        RECT 2743.045 3249.895 2743.375 3249.910 ;
        RECT 2752.910 3249.900 2753.290 3249.910 ;
        RECT 290.990 1426.450 291.370 1426.460 ;
        RECT 290.990 1426.320 300.380 1426.450 ;
        RECT 290.990 1426.150 304.000 1426.320 ;
        RECT 290.990 1426.140 291.370 1426.150 ;
        RECT 300.000 1425.720 304.000 1426.150 ;
      LAYER via3 ;
        RECT 2752.940 3251.940 2753.260 3252.260 ;
        RECT 291.020 3251.260 291.340 3251.580 ;
        RECT 1497.140 3251.260 1497.460 3251.580 ;
        RECT 1497.140 3249.900 1497.460 3250.220 ;
        RECT 2752.940 3249.900 2753.260 3250.220 ;
        RECT 291.020 1426.140 291.340 1426.460 ;
      LAYER met4 ;
        RECT 2752.935 3251.935 2753.265 3252.265 ;
        RECT 291.015 3251.255 291.345 3251.585 ;
        RECT 1497.135 3251.255 1497.465 3251.585 ;
        RECT 291.030 1426.465 291.330 3251.255 ;
        RECT 1497.150 3250.225 1497.450 3251.255 ;
        RECT 2752.950 3250.225 2753.250 3251.935 ;
        RECT 1497.135 3249.895 1497.465 3250.225 ;
        RECT 2752.935 3249.895 2753.265 3250.225 ;
        RECT 291.015 1426.135 291.345 1426.465 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 290.790 3484.900 291.110 3484.960 ;
        RECT 2900.830 3484.900 2901.150 3484.960 ;
        RECT 290.790 3484.760 2901.150 3484.900 ;
        RECT 290.790 3484.700 291.110 3484.760 ;
        RECT 2900.830 3484.700 2901.150 3484.760 ;
      LAYER via ;
        RECT 290.820 3484.700 291.080 3484.960 ;
        RECT 2900.860 3484.700 2901.120 3484.960 ;
      LAYER met2 ;
        RECT 2900.850 3489.915 2901.130 3490.285 ;
        RECT 2900.920 3484.990 2901.060 3489.915 ;
        RECT 290.820 3484.670 291.080 3484.990 ;
        RECT 2900.860 3484.670 2901.120 3484.990 ;
        RECT 290.880 2196.925 291.020 3484.670 ;
        RECT 290.810 2196.555 291.090 2196.925 ;
      LAYER via2 ;
        RECT 2900.850 3489.960 2901.130 3490.240 ;
        RECT 290.810 2196.600 291.090 2196.880 ;
      LAYER met3 ;
        RECT 2900.825 3490.250 2901.155 3490.265 ;
        RECT 2917.600 3490.250 2924.800 3490.700 ;
        RECT 2900.825 3489.950 2924.800 3490.250 ;
        RECT 2900.825 3489.935 2901.155 3489.950 ;
        RECT 2917.600 3489.500 2924.800 3489.950 ;
        RECT 290.785 2196.890 291.115 2196.905 ;
        RECT 293.750 2196.890 294.130 2196.900 ;
        RECT 290.785 2196.590 294.130 2196.890 ;
        RECT 290.785 2196.575 291.115 2196.590 ;
        RECT 293.750 2196.580 294.130 2196.590 ;
        RECT 293.750 1457.730 294.130 1457.740 ;
        RECT 293.750 1457.600 300.380 1457.730 ;
        RECT 293.750 1457.430 304.000 1457.600 ;
        RECT 293.750 1457.420 294.130 1457.430 ;
        RECT 300.000 1457.000 304.000 1457.430 ;
      LAYER via3 ;
        RECT 293.780 2196.580 294.100 2196.900 ;
        RECT 293.780 1457.420 294.100 1457.740 ;
      LAYER met4 ;
        RECT 293.775 2196.575 294.105 2196.905 ;
        RECT 293.790 1457.745 294.090 2196.575 ;
        RECT 293.775 1457.415 294.105 1457.745 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
        RECT 2635.960 3502.525 2636.100 3517.600 ;
        RECT 2635.890 3502.155 2636.170 3502.525 ;
        RECT 299.090 2897.635 299.370 2898.005 ;
        RECT 299.160 2851.085 299.300 2897.635 ;
        RECT 299.090 2850.715 299.370 2851.085 ;
      LAYER via2 ;
        RECT 2635.890 3502.200 2636.170 3502.480 ;
        RECT 299.090 2897.680 299.370 2897.960 ;
        RECT 299.090 2850.760 299.370 2851.040 ;
      LAYER met3 ;
        RECT 295.590 3502.490 295.970 3502.500 ;
        RECT 2635.865 3502.490 2636.195 3502.505 ;
        RECT 295.590 3502.190 2636.195 3502.490 ;
        RECT 295.590 3502.180 295.970 3502.190 ;
        RECT 2635.865 3502.175 2636.195 3502.190 ;
        RECT 296.510 2908.170 296.890 2908.180 ;
        RECT 299.270 2908.170 299.650 2908.180 ;
        RECT 296.510 2907.870 299.650 2908.170 ;
        RECT 296.510 2907.860 296.890 2907.870 ;
        RECT 299.270 2907.860 299.650 2907.870 ;
        RECT 299.065 2897.980 299.395 2897.985 ;
        RECT 299.065 2897.970 299.650 2897.980 ;
        RECT 298.840 2897.670 299.650 2897.970 ;
        RECT 299.065 2897.660 299.650 2897.670 ;
        RECT 299.065 2897.655 299.395 2897.660 ;
        RECT 299.065 2851.050 299.395 2851.065 ;
        RECT 298.390 2850.750 299.395 2851.050 ;
        RECT 298.390 2850.380 298.690 2850.750 ;
        RECT 299.065 2850.735 299.395 2850.750 ;
        RECT 298.350 2850.060 298.730 2850.380 ;
        RECT 298.350 2816.370 298.730 2816.380 ;
        RECT 297.470 2816.070 298.730 2816.370 ;
        RECT 297.470 2815.020 297.770 2816.070 ;
        RECT 298.350 2816.060 298.730 2816.070 ;
        RECT 297.430 2814.700 297.810 2815.020 ;
        RECT 295.590 1489.690 295.970 1489.700 ;
        RECT 295.590 1489.560 300.380 1489.690 ;
        RECT 295.590 1489.390 304.000 1489.560 ;
        RECT 295.590 1489.380 295.970 1489.390 ;
        RECT 300.000 1488.960 304.000 1489.390 ;
      LAYER via3 ;
        RECT 295.620 3502.180 295.940 3502.500 ;
        RECT 296.540 2907.860 296.860 2908.180 ;
        RECT 299.300 2907.860 299.620 2908.180 ;
        RECT 299.300 2897.660 299.620 2897.980 ;
        RECT 298.380 2850.060 298.700 2850.380 ;
        RECT 298.380 2816.060 298.700 2816.380 ;
        RECT 297.460 2814.700 297.780 2815.020 ;
        RECT 295.620 1489.380 295.940 1489.700 ;
      LAYER met4 ;
        RECT 295.615 3502.175 295.945 3502.505 ;
        RECT 295.630 2983.650 295.930 3502.175 ;
        RECT 295.630 2983.350 296.850 2983.650 ;
        RECT 296.550 2908.185 296.850 2983.350 ;
        RECT 296.535 2907.855 296.865 2908.185 ;
        RECT 299.295 2907.855 299.625 2908.185 ;
        RECT 299.310 2897.985 299.610 2907.855 ;
        RECT 299.295 2897.655 299.625 2897.985 ;
        RECT 298.375 2850.055 298.705 2850.385 ;
        RECT 298.390 2816.385 298.690 2850.055 ;
        RECT 298.375 2816.055 298.705 2816.385 ;
        RECT 297.455 2814.695 297.785 2815.025 ;
        RECT 297.470 2766.050 297.770 2814.695 ;
        RECT 296.550 2765.750 297.770 2766.050 ;
        RECT 296.550 2762.650 296.850 2765.750 ;
        RECT 295.630 2762.350 296.850 2762.650 ;
        RECT 295.630 2290.050 295.930 2762.350 ;
        RECT 295.630 2289.750 296.850 2290.050 ;
        RECT 296.550 2194.850 296.850 2289.750 ;
        RECT 295.630 2194.550 296.850 2194.850 ;
        RECT 295.630 1489.705 295.930 2194.550 ;
        RECT 295.615 1489.375 295.945 1489.705 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 296.310 3501.560 296.630 3501.620 ;
        RECT 2311.570 3501.560 2311.890 3501.620 ;
        RECT 296.310 3501.420 2311.890 3501.560 ;
        RECT 296.310 3501.360 296.630 3501.420 ;
        RECT 2311.570 3501.360 2311.890 3501.420 ;
      LAYER via ;
        RECT 296.340 3501.360 296.600 3501.620 ;
        RECT 2311.600 3501.360 2311.860 3501.620 ;
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
        RECT 2311.660 3501.650 2311.800 3517.600 ;
        RECT 296.340 3501.330 296.600 3501.650 ;
        RECT 2311.600 3501.330 2311.860 3501.650 ;
        RECT 296.400 1521.005 296.540 3501.330 ;
        RECT 296.330 1520.635 296.610 1521.005 ;
      LAYER via2 ;
        RECT 296.330 1520.680 296.610 1520.960 ;
      LAYER met3 ;
        RECT 296.305 1520.970 296.635 1520.985 ;
        RECT 296.305 1520.840 300.380 1520.970 ;
        RECT 296.305 1520.670 304.000 1520.840 ;
        RECT 296.305 1520.655 296.635 1520.670 ;
        RECT 300.000 1520.240 304.000 1520.670 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 295.850 3502.240 296.170 3502.300 ;
        RECT 1987.270 3502.240 1987.590 3502.300 ;
        RECT 295.850 3502.100 1987.590 3502.240 ;
        RECT 295.850 3502.040 296.170 3502.100 ;
        RECT 1987.270 3502.040 1987.590 3502.100 ;
      LAYER via ;
        RECT 295.880 3502.040 296.140 3502.300 ;
        RECT 1987.300 3502.040 1987.560 3502.300 ;
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
        RECT 1987.360 3502.330 1987.500 3517.600 ;
        RECT 295.880 3502.010 296.140 3502.330 ;
        RECT 1987.300 3502.010 1987.560 3502.330 ;
        RECT 295.940 1552.965 296.080 3502.010 ;
        RECT 295.870 1552.595 296.150 1552.965 ;
      LAYER via2 ;
        RECT 295.870 1552.640 296.150 1552.920 ;
      LAYER met3 ;
        RECT 295.845 1552.930 296.175 1552.945 ;
        RECT 295.845 1552.800 300.380 1552.930 ;
        RECT 295.845 1552.630 304.000 1552.800 ;
        RECT 295.845 1552.615 296.175 1552.630 ;
        RECT 300.000 1552.200 304.000 1552.630 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 294.930 3502.920 295.250 3502.980 ;
        RECT 1662.510 3502.920 1662.830 3502.980 ;
        RECT 294.930 3502.780 1662.830 3502.920 ;
        RECT 294.930 3502.720 295.250 3502.780 ;
        RECT 1662.510 3502.720 1662.830 3502.780 ;
      LAYER via ;
        RECT 294.960 3502.720 295.220 3502.980 ;
        RECT 1662.540 3502.720 1662.800 3502.980 ;
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
        RECT 1662.600 3503.010 1662.740 3517.600 ;
        RECT 294.960 3502.690 295.220 3503.010 ;
        RECT 1662.540 3502.690 1662.800 3503.010 ;
        RECT 295.020 1584.245 295.160 3502.690 ;
        RECT 294.950 1583.875 295.230 1584.245 ;
      LAYER via2 ;
        RECT 294.950 1583.920 295.230 1584.200 ;
      LAYER met3 ;
        RECT 294.925 1584.210 295.255 1584.225 ;
        RECT 294.925 1584.080 300.380 1584.210 ;
        RECT 294.925 1583.910 304.000 1584.080 ;
        RECT 294.925 1583.895 295.255 1583.910 ;
        RECT 300.000 1583.480 304.000 1583.910 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 294.470 3503.940 294.790 3504.000 ;
        RECT 1338.210 3503.940 1338.530 3504.000 ;
        RECT 294.470 3503.800 1338.530 3503.940 ;
        RECT 294.470 3503.740 294.790 3503.800 ;
        RECT 1338.210 3503.740 1338.530 3503.800 ;
      LAYER via ;
        RECT 294.500 3503.740 294.760 3504.000 ;
        RECT 1338.240 3503.740 1338.500 3504.000 ;
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
        RECT 1338.300 3504.030 1338.440 3517.600 ;
        RECT 294.500 3503.710 294.760 3504.030 ;
        RECT 1338.240 3503.710 1338.500 3504.030 ;
        RECT 294.560 1615.525 294.700 3503.710 ;
        RECT 294.490 1615.155 294.770 1615.525 ;
      LAYER via2 ;
        RECT 294.490 1615.200 294.770 1615.480 ;
      LAYER met3 ;
        RECT 294.465 1615.490 294.795 1615.505 ;
        RECT 294.465 1615.360 300.380 1615.490 ;
        RECT 294.465 1615.190 304.000 1615.360 ;
        RECT 294.465 1615.175 294.795 1615.190 ;
        RECT 300.000 1614.760 304.000 1615.190 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 448.110 436.460 448.430 436.520 ;
        RECT 482.610 436.460 482.930 436.520 ;
        RECT 448.110 436.320 482.930 436.460 ;
        RECT 448.110 436.260 448.430 436.320 ;
        RECT 482.610 436.260 482.930 436.320 ;
        RECT 727.790 435.780 728.110 435.840 ;
        RECT 772.410 435.780 772.730 435.840 ;
        RECT 727.790 435.640 772.730 435.780 ;
        RECT 727.790 435.580 728.110 435.640 ;
        RECT 772.410 435.580 772.730 435.640 ;
        RECT 580.130 435.100 580.450 435.160 ;
        RECT 604.050 435.100 604.370 435.160 ;
        RECT 580.130 434.960 604.370 435.100 ;
        RECT 580.130 434.900 580.450 434.960 ;
        RECT 604.050 434.900 604.370 434.960 ;
      LAYER via ;
        RECT 448.140 436.260 448.400 436.520 ;
        RECT 482.640 436.260 482.900 436.520 ;
        RECT 727.820 435.580 728.080 435.840 ;
        RECT 772.440 435.580 772.700 435.840 ;
        RECT 580.160 434.900 580.420 435.160 ;
        RECT 604.080 434.900 604.340 435.160 ;
      LAYER met2 ;
        RECT 717.230 436.715 717.510 437.085 ;
        RECT 448.140 436.405 448.400 436.550 ;
        RECT 482.640 436.405 482.900 436.550 ;
        RECT 448.130 436.035 448.410 436.405 ;
        RECT 482.630 436.035 482.910 436.405 ;
        RECT 604.070 436.035 604.350 436.405 ;
        RECT 640.870 436.290 641.150 436.405 ;
        RECT 641.790 436.290 642.070 436.405 ;
        RECT 640.870 436.150 642.070 436.290 ;
        RECT 640.870 436.035 641.150 436.150 ;
        RECT 641.790 436.035 642.070 436.150 ;
        RECT 604.140 435.190 604.280 436.035 ;
        RECT 580.160 435.045 580.420 435.190 ;
        RECT 580.150 434.675 580.430 435.045 ;
        RECT 604.080 434.870 604.340 435.190 ;
        RECT 717.300 435.045 717.440 436.715 ;
        RECT 772.430 436.035 772.710 436.405 ;
        RECT 772.500 435.870 772.640 436.035 ;
        RECT 727.820 435.550 728.080 435.870 ;
        RECT 772.440 435.550 772.700 435.870 ;
        RECT 727.880 435.045 728.020 435.550 ;
        RECT 717.230 434.675 717.510 435.045 ;
        RECT 727.810 434.675 728.090 435.045 ;
      LAYER via2 ;
        RECT 717.230 436.760 717.510 437.040 ;
        RECT 448.130 436.080 448.410 436.360 ;
        RECT 482.630 436.080 482.910 436.360 ;
        RECT 604.070 436.080 604.350 436.360 ;
        RECT 640.870 436.080 641.150 436.360 ;
        RECT 641.790 436.080 642.070 436.360 ;
        RECT 580.150 434.720 580.430 435.000 ;
        RECT 772.430 436.080 772.710 436.360 ;
        RECT 717.230 434.720 717.510 435.000 ;
        RECT 727.810 434.720 728.090 435.000 ;
      LAYER met3 ;
        RECT 285.470 1047.010 285.850 1047.020 ;
        RECT 285.470 1046.880 300.380 1047.010 ;
        RECT 285.470 1046.710 304.000 1046.880 ;
        RECT 285.470 1046.700 285.850 1046.710 ;
        RECT 300.000 1046.280 304.000 1046.710 ;
        RECT 2917.600 439.770 2924.800 440.220 ;
        RECT 2916.710 439.470 2924.800 439.770 ;
        RECT 578.950 437.050 579.330 437.060 ;
        RECT 544.030 436.750 579.330 437.050 ;
        RECT 285.470 436.370 285.850 436.380 ;
        RECT 448.105 436.370 448.435 436.385 ;
        RECT 285.470 436.070 324.450 436.370 ;
        RECT 285.470 436.060 285.850 436.070 ;
        RECT 324.150 435.690 324.450 436.070 ;
        RECT 372.910 436.070 448.435 436.370 ;
        RECT 324.150 435.390 372.290 435.690 ;
        RECT 371.990 435.010 372.290 435.390 ;
        RECT 372.910 435.010 373.210 436.070 ;
        RECT 448.105 436.055 448.435 436.070 ;
        RECT 482.605 436.370 482.935 436.385 ;
        RECT 482.605 436.070 496.490 436.370 ;
        RECT 482.605 436.055 482.935 436.070 ;
        RECT 371.990 434.710 373.210 435.010 ;
        RECT 496.190 435.010 496.490 436.070 ;
        RECT 544.030 435.690 544.330 436.750 ;
        RECT 578.950 436.740 579.330 436.750 ;
        RECT 669.110 437.050 669.490 437.060 ;
        RECT 717.205 437.050 717.535 437.065 ;
        RECT 669.110 436.750 717.535 437.050 ;
        RECT 669.110 436.740 669.490 436.750 ;
        RECT 717.205 436.735 717.535 436.750 ;
        RECT 604.045 436.370 604.375 436.385 ;
        RECT 640.845 436.370 641.175 436.385 ;
        RECT 604.045 436.070 641.175 436.370 ;
        RECT 604.045 436.055 604.375 436.070 ;
        RECT 640.845 436.055 641.175 436.070 ;
        RECT 641.765 436.370 642.095 436.385 ;
        RECT 772.405 436.370 772.735 436.385 ;
        RECT 641.765 436.070 651.970 436.370 ;
        RECT 641.765 436.055 642.095 436.070 ;
        RECT 497.110 435.390 544.330 435.690 ;
        RECT 651.670 435.690 651.970 436.070 ;
        RECT 772.405 436.070 807.450 436.370 ;
        RECT 772.405 436.055 772.735 436.070 ;
        RECT 669.110 435.690 669.490 435.700 ;
        RECT 651.670 435.390 669.490 435.690 ;
        RECT 807.150 435.690 807.450 436.070 ;
        RECT 855.910 436.070 904.050 436.370 ;
        RECT 807.150 435.390 855.290 435.690 ;
        RECT 497.110 435.010 497.410 435.390 ;
        RECT 669.110 435.380 669.490 435.390 ;
        RECT 496.190 434.710 497.410 435.010 ;
        RECT 578.950 435.010 579.330 435.020 ;
        RECT 580.125 435.010 580.455 435.025 ;
        RECT 578.950 434.710 580.455 435.010 ;
        RECT 578.950 434.700 579.330 434.710 ;
        RECT 580.125 434.695 580.455 434.710 ;
        RECT 717.205 435.010 717.535 435.025 ;
        RECT 727.785 435.010 728.115 435.025 ;
        RECT 717.205 434.710 728.115 435.010 ;
        RECT 854.990 435.010 855.290 435.390 ;
        RECT 855.910 435.010 856.210 436.070 ;
        RECT 903.750 435.690 904.050 436.070 ;
        RECT 952.510 436.070 1000.650 436.370 ;
        RECT 903.750 435.390 951.890 435.690 ;
        RECT 854.990 434.710 856.210 435.010 ;
        RECT 951.590 435.010 951.890 435.390 ;
        RECT 952.510 435.010 952.810 436.070 ;
        RECT 1000.350 435.690 1000.650 436.070 ;
        RECT 1049.110 436.070 1097.250 436.370 ;
        RECT 1000.350 435.390 1048.490 435.690 ;
        RECT 951.590 434.710 952.810 435.010 ;
        RECT 1048.190 435.010 1048.490 435.390 ;
        RECT 1049.110 435.010 1049.410 436.070 ;
        RECT 1096.950 435.690 1097.250 436.070 ;
        RECT 1145.710 436.070 1193.850 436.370 ;
        RECT 1096.950 435.390 1145.090 435.690 ;
        RECT 1048.190 434.710 1049.410 435.010 ;
        RECT 1144.790 435.010 1145.090 435.390 ;
        RECT 1145.710 435.010 1146.010 436.070 ;
        RECT 1193.550 435.690 1193.850 436.070 ;
        RECT 1242.310 436.070 1290.450 436.370 ;
        RECT 1193.550 435.390 1241.690 435.690 ;
        RECT 1144.790 434.710 1146.010 435.010 ;
        RECT 1241.390 435.010 1241.690 435.390 ;
        RECT 1242.310 435.010 1242.610 436.070 ;
        RECT 1290.150 435.690 1290.450 436.070 ;
        RECT 1338.910 436.070 1387.050 436.370 ;
        RECT 1290.150 435.390 1338.290 435.690 ;
        RECT 1241.390 434.710 1242.610 435.010 ;
        RECT 1337.990 435.010 1338.290 435.390 ;
        RECT 1338.910 435.010 1339.210 436.070 ;
        RECT 1386.750 435.690 1387.050 436.070 ;
        RECT 1435.510 436.070 1483.650 436.370 ;
        RECT 1386.750 435.390 1434.890 435.690 ;
        RECT 1337.990 434.710 1339.210 435.010 ;
        RECT 1434.590 435.010 1434.890 435.390 ;
        RECT 1435.510 435.010 1435.810 436.070 ;
        RECT 1483.350 435.690 1483.650 436.070 ;
        RECT 1532.110 436.070 1580.250 436.370 ;
        RECT 1483.350 435.390 1531.490 435.690 ;
        RECT 1434.590 434.710 1435.810 435.010 ;
        RECT 1531.190 435.010 1531.490 435.390 ;
        RECT 1532.110 435.010 1532.410 436.070 ;
        RECT 1579.950 435.690 1580.250 436.070 ;
        RECT 1628.710 436.070 1676.850 436.370 ;
        RECT 1579.950 435.390 1628.090 435.690 ;
        RECT 1531.190 434.710 1532.410 435.010 ;
        RECT 1627.790 435.010 1628.090 435.390 ;
        RECT 1628.710 435.010 1629.010 436.070 ;
        RECT 1676.550 435.690 1676.850 436.070 ;
        RECT 1725.310 436.070 1773.450 436.370 ;
        RECT 1676.550 435.390 1724.690 435.690 ;
        RECT 1627.790 434.710 1629.010 435.010 ;
        RECT 1724.390 435.010 1724.690 435.390 ;
        RECT 1725.310 435.010 1725.610 436.070 ;
        RECT 1773.150 435.690 1773.450 436.070 ;
        RECT 1821.910 436.070 1870.050 436.370 ;
        RECT 1773.150 435.390 1821.290 435.690 ;
        RECT 1724.390 434.710 1725.610 435.010 ;
        RECT 1820.990 435.010 1821.290 435.390 ;
        RECT 1821.910 435.010 1822.210 436.070 ;
        RECT 1869.750 435.690 1870.050 436.070 ;
        RECT 1918.510 436.070 1966.650 436.370 ;
        RECT 1869.750 435.390 1917.890 435.690 ;
        RECT 1820.990 434.710 1822.210 435.010 ;
        RECT 1917.590 435.010 1917.890 435.390 ;
        RECT 1918.510 435.010 1918.810 436.070 ;
        RECT 1966.350 435.690 1966.650 436.070 ;
        RECT 2015.110 436.070 2063.250 436.370 ;
        RECT 1966.350 435.390 2014.490 435.690 ;
        RECT 1917.590 434.710 1918.810 435.010 ;
        RECT 2014.190 435.010 2014.490 435.390 ;
        RECT 2015.110 435.010 2015.410 436.070 ;
        RECT 2062.950 435.690 2063.250 436.070 ;
        RECT 2111.710 436.070 2159.850 436.370 ;
        RECT 2062.950 435.390 2111.090 435.690 ;
        RECT 2014.190 434.710 2015.410 435.010 ;
        RECT 2110.790 435.010 2111.090 435.390 ;
        RECT 2111.710 435.010 2112.010 436.070 ;
        RECT 2159.550 435.690 2159.850 436.070 ;
        RECT 2208.310 436.070 2256.450 436.370 ;
        RECT 2159.550 435.390 2207.690 435.690 ;
        RECT 2110.790 434.710 2112.010 435.010 ;
        RECT 2207.390 435.010 2207.690 435.390 ;
        RECT 2208.310 435.010 2208.610 436.070 ;
        RECT 2256.150 435.690 2256.450 436.070 ;
        RECT 2304.910 436.070 2353.050 436.370 ;
        RECT 2256.150 435.390 2304.290 435.690 ;
        RECT 2207.390 434.710 2208.610 435.010 ;
        RECT 2303.990 435.010 2304.290 435.390 ;
        RECT 2304.910 435.010 2305.210 436.070 ;
        RECT 2352.750 435.690 2353.050 436.070 ;
        RECT 2401.510 436.070 2449.650 436.370 ;
        RECT 2352.750 435.390 2400.890 435.690 ;
        RECT 2303.990 434.710 2305.210 435.010 ;
        RECT 2400.590 435.010 2400.890 435.390 ;
        RECT 2401.510 435.010 2401.810 436.070 ;
        RECT 2449.350 435.690 2449.650 436.070 ;
        RECT 2498.110 436.070 2546.250 436.370 ;
        RECT 2449.350 435.390 2497.490 435.690 ;
        RECT 2400.590 434.710 2401.810 435.010 ;
        RECT 2497.190 435.010 2497.490 435.390 ;
        RECT 2498.110 435.010 2498.410 436.070 ;
        RECT 2545.950 435.690 2546.250 436.070 ;
        RECT 2594.710 436.070 2642.850 436.370 ;
        RECT 2545.950 435.390 2594.090 435.690 ;
        RECT 2497.190 434.710 2498.410 435.010 ;
        RECT 2593.790 435.010 2594.090 435.390 ;
        RECT 2594.710 435.010 2595.010 436.070 ;
        RECT 2642.550 435.690 2642.850 436.070 ;
        RECT 2691.310 436.070 2739.450 436.370 ;
        RECT 2642.550 435.390 2690.690 435.690 ;
        RECT 2593.790 434.710 2595.010 435.010 ;
        RECT 2690.390 435.010 2690.690 435.390 ;
        RECT 2691.310 435.010 2691.610 436.070 ;
        RECT 2739.150 435.690 2739.450 436.070 ;
        RECT 2787.910 436.070 2836.050 436.370 ;
        RECT 2739.150 435.390 2787.290 435.690 ;
        RECT 2690.390 434.710 2691.610 435.010 ;
        RECT 2786.990 435.010 2787.290 435.390 ;
        RECT 2787.910 435.010 2788.210 436.070 ;
        RECT 2835.750 435.690 2836.050 436.070 ;
        RECT 2916.710 435.690 2917.010 439.470 ;
        RECT 2917.600 439.020 2924.800 439.470 ;
        RECT 2835.750 435.390 2883.890 435.690 ;
        RECT 2786.990 434.710 2788.210 435.010 ;
        RECT 2883.590 435.010 2883.890 435.390 ;
        RECT 2884.510 435.390 2917.010 435.690 ;
        RECT 2884.510 435.010 2884.810 435.390 ;
        RECT 2883.590 434.710 2884.810 435.010 ;
        RECT 717.205 434.695 717.535 434.710 ;
        RECT 727.785 434.695 728.115 434.710 ;
      LAYER via3 ;
        RECT 285.500 1046.700 285.820 1047.020 ;
        RECT 285.500 436.060 285.820 436.380 ;
        RECT 578.980 436.740 579.300 437.060 ;
        RECT 669.140 436.740 669.460 437.060 ;
        RECT 669.140 435.380 669.460 435.700 ;
        RECT 578.980 434.700 579.300 435.020 ;
      LAYER met4 ;
        RECT 285.495 1046.695 285.825 1047.025 ;
        RECT 285.510 436.385 285.810 1046.695 ;
        RECT 578.975 436.735 579.305 437.065 ;
        RECT 669.135 436.735 669.465 437.065 ;
        RECT 285.495 436.055 285.825 436.385 ;
        RECT 578.990 435.025 579.290 436.735 ;
        RECT 669.150 435.705 669.450 436.735 ;
        RECT 669.135 435.375 669.465 435.705 ;
        RECT 578.975 434.695 579.305 435.025 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 294.010 3504.620 294.330 3504.680 ;
        RECT 1013.910 3504.620 1014.230 3504.680 ;
        RECT 294.010 3504.480 1014.230 3504.620 ;
        RECT 294.010 3504.420 294.330 3504.480 ;
        RECT 1013.910 3504.420 1014.230 3504.480 ;
      LAYER via ;
        RECT 294.040 3504.420 294.300 3504.680 ;
        RECT 1013.940 3504.420 1014.200 3504.680 ;
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
        RECT 1014.000 3504.710 1014.140 3517.600 ;
        RECT 294.040 3504.390 294.300 3504.710 ;
        RECT 1013.940 3504.390 1014.200 3504.710 ;
        RECT 294.100 1647.485 294.240 3504.390 ;
        RECT 294.030 1647.115 294.310 1647.485 ;
      LAYER via2 ;
        RECT 294.030 1647.160 294.310 1647.440 ;
      LAYER met3 ;
        RECT 294.005 1647.450 294.335 1647.465 ;
        RECT 294.005 1647.320 300.380 1647.450 ;
        RECT 294.005 1647.150 304.000 1647.320 ;
        RECT 294.005 1647.135 294.335 1647.150 ;
        RECT 300.000 1646.720 304.000 1647.150 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 293.550 3500.540 293.870 3500.600 ;
        RECT 689.150 3500.540 689.470 3500.600 ;
        RECT 293.550 3500.400 689.470 3500.540 ;
        RECT 293.550 3500.340 293.870 3500.400 ;
        RECT 689.150 3500.340 689.470 3500.400 ;
      LAYER via ;
        RECT 293.580 3500.340 293.840 3500.600 ;
        RECT 689.180 3500.340 689.440 3500.600 ;
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
        RECT 689.240 3500.630 689.380 3517.600 ;
        RECT 293.580 3500.310 293.840 3500.630 ;
        RECT 689.180 3500.310 689.440 3500.630 ;
        RECT 293.640 1678.765 293.780 3500.310 ;
        RECT 293.570 1678.395 293.850 1678.765 ;
      LAYER via2 ;
        RECT 293.570 1678.440 293.850 1678.720 ;
      LAYER met3 ;
        RECT 293.545 1678.730 293.875 1678.745 ;
        RECT 293.545 1678.600 300.380 1678.730 ;
        RECT 293.545 1678.430 304.000 1678.600 ;
        RECT 293.545 1678.415 293.875 1678.430 ;
        RECT 300.000 1678.000 304.000 1678.430 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 292.630 3500.200 292.950 3500.260 ;
        RECT 364.850 3500.200 365.170 3500.260 ;
        RECT 292.630 3500.060 365.170 3500.200 ;
        RECT 292.630 3500.000 292.950 3500.060 ;
        RECT 364.850 3500.000 365.170 3500.060 ;
      LAYER via ;
        RECT 292.660 3500.000 292.920 3500.260 ;
        RECT 364.880 3500.000 365.140 3500.260 ;
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
        RECT 364.940 3500.290 365.080 3517.600 ;
        RECT 292.660 3499.970 292.920 3500.290 ;
        RECT 364.880 3499.970 365.140 3500.290 ;
        RECT 292.720 1710.725 292.860 3499.970 ;
        RECT 292.650 1710.355 292.930 1710.725 ;
      LAYER via2 ;
        RECT 292.650 1710.400 292.930 1710.680 ;
      LAYER met3 ;
        RECT 292.625 1710.690 292.955 1710.705 ;
        RECT 292.625 1710.560 300.380 1710.690 ;
        RECT 292.625 1710.390 304.000 1710.560 ;
        RECT 292.625 1710.375 292.955 1710.390 ;
        RECT 300.000 1709.960 304.000 1710.390 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 40.550 3501.900 40.870 3501.960 ;
        RECT 65.390 3501.900 65.710 3501.960 ;
        RECT 40.550 3501.760 65.710 3501.900 ;
        RECT 40.550 3501.700 40.870 3501.760 ;
        RECT 65.390 3501.700 65.710 3501.760 ;
        RECT 65.390 1745.460 65.710 1745.520 ;
        RECT 282.970 1745.460 283.290 1745.520 ;
        RECT 65.390 1745.320 283.290 1745.460 ;
        RECT 65.390 1745.260 65.710 1745.320 ;
        RECT 282.970 1745.260 283.290 1745.320 ;
      LAYER via ;
        RECT 40.580 3501.700 40.840 3501.960 ;
        RECT 65.420 3501.700 65.680 3501.960 ;
        RECT 65.420 1745.260 65.680 1745.520 ;
        RECT 283.000 1745.260 283.260 1745.520 ;
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
        RECT 40.640 3501.990 40.780 3517.600 ;
        RECT 40.580 3501.670 40.840 3501.990 ;
        RECT 65.420 3501.670 65.680 3501.990 ;
        RECT 65.480 1745.550 65.620 3501.670 ;
        RECT 65.420 1745.230 65.680 1745.550 ;
        RECT 283.000 1745.230 283.260 1745.550 ;
        RECT 283.060 1742.005 283.200 1745.230 ;
        RECT 282.990 1741.635 283.270 1742.005 ;
      LAYER via2 ;
        RECT 282.990 1741.680 283.270 1741.960 ;
      LAYER met3 ;
        RECT 282.965 1741.970 283.295 1741.985 ;
        RECT 282.965 1741.840 300.380 1741.970 ;
        RECT 282.965 1741.670 304.000 1741.840 ;
        RECT 282.965 1741.655 283.295 1741.670 ;
        RECT 300.000 1741.240 304.000 1741.670 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.250 3263.900 15.570 3263.960 ;
        RECT 72.290 3263.900 72.610 3263.960 ;
        RECT 15.250 3263.760 72.610 3263.900 ;
        RECT 15.250 3263.700 15.570 3263.760 ;
        RECT 72.290 3263.700 72.610 3263.760 ;
        RECT 72.290 1780.140 72.610 1780.200 ;
        RECT 282.970 1780.140 283.290 1780.200 ;
        RECT 72.290 1780.000 283.290 1780.140 ;
        RECT 72.290 1779.940 72.610 1780.000 ;
        RECT 282.970 1779.940 283.290 1780.000 ;
      LAYER via ;
        RECT 15.280 3263.700 15.540 3263.960 ;
        RECT 72.320 3263.700 72.580 3263.960 ;
        RECT 72.320 1779.940 72.580 1780.200 ;
        RECT 283.000 1779.940 283.260 1780.200 ;
      LAYER met2 ;
        RECT 15.270 3267.555 15.550 3267.925 ;
        RECT 15.340 3263.990 15.480 3267.555 ;
        RECT 15.280 3263.670 15.540 3263.990 ;
        RECT 72.320 3263.670 72.580 3263.990 ;
        RECT 72.380 1780.230 72.520 3263.670 ;
        RECT 72.320 1779.910 72.580 1780.230 ;
        RECT 283.000 1779.910 283.260 1780.230 ;
        RECT 283.060 1773.965 283.200 1779.910 ;
        RECT 282.990 1773.595 283.270 1773.965 ;
      LAYER via2 ;
        RECT 15.270 3267.600 15.550 3267.880 ;
        RECT 282.990 1773.640 283.270 1773.920 ;
      LAYER met3 ;
        RECT -4.800 3267.890 2.400 3268.340 ;
        RECT 15.245 3267.890 15.575 3267.905 ;
        RECT -4.800 3267.590 15.575 3267.890 ;
        RECT -4.800 3267.140 2.400 3267.590 ;
        RECT 15.245 3267.575 15.575 3267.590 ;
        RECT 282.965 1773.930 283.295 1773.945 ;
        RECT 282.965 1773.800 300.380 1773.930 ;
        RECT 282.965 1773.630 304.000 1773.800 ;
        RECT 282.965 1773.615 283.295 1773.630 ;
        RECT 300.000 1773.200 304.000 1773.630 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.170 2974.220 16.490 2974.280 ;
        RECT 86.550 2974.220 86.870 2974.280 ;
        RECT 16.170 2974.080 86.870 2974.220 ;
        RECT 16.170 2974.020 16.490 2974.080 ;
        RECT 86.550 2974.020 86.870 2974.080 ;
        RECT 86.550 1807.680 86.870 1807.740 ;
        RECT 282.970 1807.680 283.290 1807.740 ;
        RECT 86.550 1807.540 283.290 1807.680 ;
        RECT 86.550 1807.480 86.870 1807.540 ;
        RECT 282.970 1807.480 283.290 1807.540 ;
      LAYER via ;
        RECT 16.200 2974.020 16.460 2974.280 ;
        RECT 86.580 2974.020 86.840 2974.280 ;
        RECT 86.580 1807.480 86.840 1807.740 ;
        RECT 283.000 1807.480 283.260 1807.740 ;
      LAYER met2 ;
        RECT 16.190 2979.915 16.470 2980.285 ;
        RECT 16.260 2974.310 16.400 2979.915 ;
        RECT 16.200 2973.990 16.460 2974.310 ;
        RECT 86.580 2973.990 86.840 2974.310 ;
        RECT 86.640 1807.770 86.780 2973.990 ;
        RECT 86.580 1807.450 86.840 1807.770 ;
        RECT 283.000 1807.450 283.260 1807.770 ;
        RECT 283.060 1805.245 283.200 1807.450 ;
        RECT 282.990 1804.875 283.270 1805.245 ;
      LAYER via2 ;
        RECT 16.190 2979.960 16.470 2980.240 ;
        RECT 282.990 1804.920 283.270 1805.200 ;
      LAYER met3 ;
        RECT -4.800 2980.250 2.400 2980.700 ;
        RECT 16.165 2980.250 16.495 2980.265 ;
        RECT -4.800 2979.950 16.495 2980.250 ;
        RECT -4.800 2979.500 2.400 2979.950 ;
        RECT 16.165 2979.935 16.495 2979.950 ;
        RECT 282.965 1805.210 283.295 1805.225 ;
        RECT 282.965 1805.080 300.380 1805.210 ;
        RECT 282.965 1804.910 304.000 1805.080 ;
        RECT 282.965 1804.895 283.295 1804.910 ;
        RECT 300.000 1804.480 304.000 1804.910 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.010 1842.360 18.330 1842.420 ;
        RECT 282.970 1842.360 283.290 1842.420 ;
        RECT 18.010 1842.220 283.290 1842.360 ;
        RECT 18.010 1842.160 18.330 1842.220 ;
        RECT 282.970 1842.160 283.290 1842.220 ;
      LAYER via ;
        RECT 18.040 1842.160 18.300 1842.420 ;
        RECT 283.000 1842.160 283.260 1842.420 ;
      LAYER met2 ;
        RECT 18.030 2692.955 18.310 2693.325 ;
        RECT 18.100 1842.450 18.240 2692.955 ;
        RECT 18.040 1842.130 18.300 1842.450 ;
        RECT 283.000 1842.130 283.260 1842.450 ;
        RECT 283.060 1837.205 283.200 1842.130 ;
        RECT 282.990 1836.835 283.270 1837.205 ;
      LAYER via2 ;
        RECT 18.030 2693.000 18.310 2693.280 ;
        RECT 282.990 1836.880 283.270 1837.160 ;
      LAYER met3 ;
        RECT -4.800 2693.290 2.400 2693.740 ;
        RECT 18.005 2693.290 18.335 2693.305 ;
        RECT -4.800 2692.990 18.335 2693.290 ;
        RECT -4.800 2692.540 2.400 2692.990 ;
        RECT 18.005 2692.975 18.335 2692.990 ;
        RECT 282.965 1837.170 283.295 1837.185 ;
        RECT 282.965 1837.040 300.380 1837.170 ;
        RECT 282.965 1836.870 304.000 1837.040 ;
        RECT 282.965 1836.855 283.295 1836.870 ;
        RECT 300.000 1836.440 304.000 1836.870 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 14.790 2401.320 15.110 2401.380 ;
        RECT 100.350 2401.320 100.670 2401.380 ;
        RECT 14.790 2401.180 100.670 2401.320 ;
        RECT 14.790 2401.120 15.110 2401.180 ;
        RECT 100.350 2401.120 100.670 2401.180 ;
        RECT 100.350 1869.900 100.670 1869.960 ;
        RECT 282.970 1869.900 283.290 1869.960 ;
        RECT 100.350 1869.760 283.290 1869.900 ;
        RECT 100.350 1869.700 100.670 1869.760 ;
        RECT 282.970 1869.700 283.290 1869.760 ;
      LAYER via ;
        RECT 14.820 2401.120 15.080 2401.380 ;
        RECT 100.380 2401.120 100.640 2401.380 ;
        RECT 100.380 1869.700 100.640 1869.960 ;
        RECT 283.000 1869.700 283.260 1869.960 ;
      LAYER met2 ;
        RECT 14.810 2405.315 15.090 2405.685 ;
        RECT 14.880 2401.410 15.020 2405.315 ;
        RECT 14.820 2401.090 15.080 2401.410 ;
        RECT 100.380 2401.090 100.640 2401.410 ;
        RECT 100.440 1869.990 100.580 2401.090 ;
        RECT 100.380 1869.670 100.640 1869.990 ;
        RECT 283.000 1869.670 283.260 1869.990 ;
        RECT 283.060 1868.485 283.200 1869.670 ;
        RECT 282.990 1868.115 283.270 1868.485 ;
      LAYER via2 ;
        RECT 14.810 2405.360 15.090 2405.640 ;
        RECT 282.990 1868.160 283.270 1868.440 ;
      LAYER met3 ;
        RECT -4.800 2405.650 2.400 2406.100 ;
        RECT 14.785 2405.650 15.115 2405.665 ;
        RECT -4.800 2405.350 15.115 2405.650 ;
        RECT -4.800 2404.900 2.400 2405.350 ;
        RECT 14.785 2405.335 15.115 2405.350 ;
        RECT 282.965 1868.450 283.295 1868.465 ;
        RECT 282.965 1868.320 300.380 1868.450 ;
        RECT 282.965 1868.150 304.000 1868.320 ;
        RECT 282.965 1868.135 283.295 1868.150 ;
        RECT 300.000 1867.720 304.000 1868.150 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 1903.220 16.030 1903.280 ;
        RECT 282.970 1903.220 283.290 1903.280 ;
        RECT 15.710 1903.080 283.290 1903.220 ;
        RECT 15.710 1903.020 16.030 1903.080 ;
        RECT 282.970 1903.020 283.290 1903.080 ;
      LAYER via ;
        RECT 15.740 1903.020 16.000 1903.280 ;
        RECT 283.000 1903.020 283.260 1903.280 ;
      LAYER met2 ;
        RECT 15.730 2118.355 16.010 2118.725 ;
        RECT 15.800 1903.310 15.940 2118.355 ;
        RECT 15.740 1902.990 16.000 1903.310 ;
        RECT 283.000 1902.990 283.260 1903.310 ;
        RECT 283.060 1900.445 283.200 1902.990 ;
        RECT 282.990 1900.075 283.270 1900.445 ;
      LAYER via2 ;
        RECT 15.730 2118.400 16.010 2118.680 ;
        RECT 282.990 1900.120 283.270 1900.400 ;
      LAYER met3 ;
        RECT -4.800 2118.690 2.400 2119.140 ;
        RECT 15.705 2118.690 16.035 2118.705 ;
        RECT -4.800 2118.390 16.035 2118.690 ;
        RECT -4.800 2117.940 2.400 2118.390 ;
        RECT 15.705 2118.375 16.035 2118.390 ;
        RECT 282.965 1900.410 283.295 1900.425 ;
        RECT 282.965 1900.280 300.380 1900.410 ;
        RECT 282.965 1900.110 304.000 1900.280 ;
        RECT 282.965 1900.095 283.295 1900.110 ;
        RECT 300.000 1899.680 304.000 1900.110 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.250 1925.320 15.570 1925.380 ;
        RECT 282.970 1925.320 283.290 1925.380 ;
        RECT 15.250 1925.180 283.290 1925.320 ;
        RECT 15.250 1925.120 15.570 1925.180 ;
        RECT 282.970 1925.120 283.290 1925.180 ;
      LAYER via ;
        RECT 15.280 1925.120 15.540 1925.380 ;
        RECT 283.000 1925.120 283.260 1925.380 ;
      LAYER met2 ;
        RECT 282.990 1931.355 283.270 1931.725 ;
        RECT 283.060 1925.410 283.200 1931.355 ;
        RECT 15.280 1925.090 15.540 1925.410 ;
        RECT 283.000 1925.090 283.260 1925.410 ;
        RECT 15.340 1831.085 15.480 1925.090 ;
        RECT 15.270 1830.715 15.550 1831.085 ;
      LAYER via2 ;
        RECT 282.990 1931.400 283.270 1931.680 ;
        RECT 15.270 1830.760 15.550 1831.040 ;
      LAYER met3 ;
        RECT 282.965 1931.690 283.295 1931.705 ;
        RECT 282.965 1931.560 300.380 1931.690 ;
        RECT 282.965 1931.390 304.000 1931.560 ;
        RECT 282.965 1931.375 283.295 1931.390 ;
        RECT 300.000 1930.960 304.000 1931.390 ;
        RECT -4.800 1831.050 2.400 1831.500 ;
        RECT 15.245 1831.050 15.575 1831.065 ;
        RECT -4.800 1830.750 15.575 1831.050 ;
        RECT -4.800 1830.300 2.400 1830.750 ;
        RECT 15.245 1830.735 15.575 1830.750 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 282.970 676.160 283.290 676.220 ;
        RECT 2900.830 676.160 2901.150 676.220 ;
        RECT 282.970 676.020 2901.150 676.160 ;
        RECT 282.970 675.960 283.290 676.020 ;
        RECT 2900.830 675.960 2901.150 676.020 ;
      LAYER via ;
        RECT 283.000 675.960 283.260 676.220 ;
        RECT 2900.860 675.960 2901.120 676.220 ;
      LAYER met2 ;
        RECT 282.990 1078.635 283.270 1079.005 ;
        RECT 283.060 676.250 283.200 1078.635 ;
        RECT 283.000 675.930 283.260 676.250 ;
        RECT 2900.860 675.930 2901.120 676.250 ;
        RECT 2900.920 674.405 2901.060 675.930 ;
        RECT 2900.850 674.035 2901.130 674.405 ;
      LAYER via2 ;
        RECT 282.990 1078.680 283.270 1078.960 ;
        RECT 2900.850 674.080 2901.130 674.360 ;
      LAYER met3 ;
        RECT 282.965 1078.970 283.295 1078.985 ;
        RECT 282.965 1078.840 300.380 1078.970 ;
        RECT 282.965 1078.670 304.000 1078.840 ;
        RECT 282.965 1078.655 283.295 1078.670 ;
        RECT 300.000 1078.240 304.000 1078.670 ;
        RECT 2900.825 674.370 2901.155 674.385 ;
        RECT 2917.600 674.370 2924.800 674.820 ;
        RECT 2900.825 674.070 2924.800 674.370 ;
        RECT 2900.825 674.055 2901.155 674.070 ;
        RECT 2917.600 673.620 2924.800 674.070 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 19.390 1960.000 19.710 1960.060 ;
        RECT 282.970 1960.000 283.290 1960.060 ;
        RECT 19.390 1959.860 283.290 1960.000 ;
        RECT 19.390 1959.800 19.710 1959.860 ;
        RECT 282.970 1959.800 283.290 1959.860 ;
      LAYER via ;
        RECT 19.420 1959.800 19.680 1960.060 ;
        RECT 283.000 1959.800 283.260 1960.060 ;
      LAYER met2 ;
        RECT 282.990 1962.635 283.270 1963.005 ;
        RECT 283.060 1960.090 283.200 1962.635 ;
        RECT 19.420 1959.770 19.680 1960.090 ;
        RECT 283.000 1959.770 283.260 1960.090 ;
        RECT 19.480 1544.125 19.620 1959.770 ;
        RECT 19.410 1543.755 19.690 1544.125 ;
      LAYER via2 ;
        RECT 282.990 1962.680 283.270 1962.960 ;
        RECT 19.410 1543.800 19.690 1544.080 ;
      LAYER met3 ;
        RECT 282.965 1962.970 283.295 1962.985 ;
        RECT 282.965 1962.840 300.380 1962.970 ;
        RECT 282.965 1962.670 304.000 1962.840 ;
        RECT 282.965 1962.655 283.295 1962.670 ;
        RECT 300.000 1962.240 304.000 1962.670 ;
        RECT -4.800 1544.090 2.400 1544.540 ;
        RECT 19.385 1544.090 19.715 1544.105 ;
        RECT -4.800 1543.790 19.715 1544.090 ;
        RECT -4.800 1543.340 2.400 1543.790 ;
        RECT 19.385 1543.775 19.715 1543.790 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 26.290 1994.340 26.610 1994.400 ;
        RECT 283.430 1994.340 283.750 1994.400 ;
        RECT 26.290 1994.200 283.750 1994.340 ;
        RECT 26.290 1994.140 26.610 1994.200 ;
        RECT 283.430 1994.140 283.750 1994.200 ;
        RECT 13.870 1331.340 14.190 1331.400 ;
        RECT 26.290 1331.340 26.610 1331.400 ;
        RECT 13.870 1331.200 26.610 1331.340 ;
        RECT 13.870 1331.140 14.190 1331.200 ;
        RECT 26.290 1331.140 26.610 1331.200 ;
      LAYER via ;
        RECT 26.320 1994.140 26.580 1994.400 ;
        RECT 283.460 1994.140 283.720 1994.400 ;
        RECT 13.900 1331.140 14.160 1331.400 ;
        RECT 26.320 1331.140 26.580 1331.400 ;
      LAYER met2 ;
        RECT 283.450 1994.595 283.730 1994.965 ;
        RECT 283.520 1994.430 283.660 1994.595 ;
        RECT 26.320 1994.110 26.580 1994.430 ;
        RECT 283.460 1994.110 283.720 1994.430 ;
        RECT 26.380 1331.430 26.520 1994.110 ;
        RECT 13.900 1331.110 14.160 1331.430 ;
        RECT 26.320 1331.110 26.580 1331.430 ;
        RECT 13.960 1328.565 14.100 1331.110 ;
        RECT 13.890 1328.195 14.170 1328.565 ;
      LAYER via2 ;
        RECT 283.450 1994.640 283.730 1994.920 ;
        RECT 13.890 1328.240 14.170 1328.520 ;
      LAYER met3 ;
        RECT 283.425 1994.930 283.755 1994.945 ;
        RECT 283.425 1994.800 300.380 1994.930 ;
        RECT 283.425 1994.630 304.000 1994.800 ;
        RECT 283.425 1994.615 283.755 1994.630 ;
        RECT 300.000 1994.200 304.000 1994.630 ;
        RECT -4.800 1328.530 2.400 1328.980 ;
        RECT 13.865 1328.530 14.195 1328.545 ;
        RECT -4.800 1328.230 14.195 1328.530 ;
        RECT -4.800 1327.780 2.400 1328.230 ;
        RECT 13.865 1328.215 14.195 1328.230 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 25.830 2021.880 26.150 2021.940 ;
        RECT 285.730 2021.880 286.050 2021.940 ;
        RECT 25.830 2021.740 286.050 2021.880 ;
        RECT 25.830 2021.680 26.150 2021.740 ;
        RECT 285.730 2021.680 286.050 2021.740 ;
        RECT 13.870 1115.440 14.190 1115.500 ;
        RECT 25.830 1115.440 26.150 1115.500 ;
        RECT 13.870 1115.300 26.150 1115.440 ;
        RECT 13.870 1115.240 14.190 1115.300 ;
        RECT 25.830 1115.240 26.150 1115.300 ;
      LAYER via ;
        RECT 25.860 2021.680 26.120 2021.940 ;
        RECT 285.760 2021.680 286.020 2021.940 ;
        RECT 13.900 1115.240 14.160 1115.500 ;
        RECT 25.860 1115.240 26.120 1115.500 ;
      LAYER met2 ;
        RECT 285.750 2025.875 286.030 2026.245 ;
        RECT 285.820 2021.970 285.960 2025.875 ;
        RECT 25.860 2021.650 26.120 2021.970 ;
        RECT 285.760 2021.650 286.020 2021.970 ;
        RECT 25.920 1115.530 26.060 2021.650 ;
        RECT 13.900 1115.210 14.160 1115.530 ;
        RECT 25.860 1115.210 26.120 1115.530 ;
        RECT 13.960 1113.005 14.100 1115.210 ;
        RECT 13.890 1112.635 14.170 1113.005 ;
      LAYER via2 ;
        RECT 285.750 2025.920 286.030 2026.200 ;
        RECT 13.890 1112.680 14.170 1112.960 ;
      LAYER met3 ;
        RECT 285.725 2026.210 286.055 2026.225 ;
        RECT 285.725 2026.080 300.380 2026.210 ;
        RECT 285.725 2025.910 304.000 2026.080 ;
        RECT 285.725 2025.895 286.055 2025.910 ;
        RECT 300.000 2025.480 304.000 2025.910 ;
        RECT -4.800 1112.970 2.400 1113.420 ;
        RECT 13.865 1112.970 14.195 1112.985 ;
        RECT -4.800 1112.670 14.195 1112.970 ;
        RECT -4.800 1112.220 2.400 1112.670 ;
        RECT 13.865 1112.655 14.195 1112.670 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 155.090 2056.560 155.410 2056.620 ;
        RECT 285.730 2056.560 286.050 2056.620 ;
        RECT 155.090 2056.420 286.050 2056.560 ;
        RECT 155.090 2056.360 155.410 2056.420 ;
        RECT 285.730 2056.360 286.050 2056.420 ;
        RECT 16.170 903.960 16.490 904.020 ;
        RECT 155.090 903.960 155.410 904.020 ;
        RECT 16.170 903.820 155.410 903.960 ;
        RECT 16.170 903.760 16.490 903.820 ;
        RECT 155.090 903.760 155.410 903.820 ;
      LAYER via ;
        RECT 155.120 2056.360 155.380 2056.620 ;
        RECT 285.760 2056.360 286.020 2056.620 ;
        RECT 16.200 903.760 16.460 904.020 ;
        RECT 155.120 903.760 155.380 904.020 ;
      LAYER met2 ;
        RECT 285.750 2057.835 286.030 2058.205 ;
        RECT 285.820 2056.650 285.960 2057.835 ;
        RECT 155.120 2056.330 155.380 2056.650 ;
        RECT 285.760 2056.330 286.020 2056.650 ;
        RECT 155.180 904.050 155.320 2056.330 ;
        RECT 16.200 903.730 16.460 904.050 ;
        RECT 155.120 903.730 155.380 904.050 ;
        RECT 16.260 897.445 16.400 903.730 ;
        RECT 16.190 897.075 16.470 897.445 ;
      LAYER via2 ;
        RECT 285.750 2057.880 286.030 2058.160 ;
        RECT 16.190 897.120 16.470 897.400 ;
      LAYER met3 ;
        RECT 285.725 2058.170 286.055 2058.185 ;
        RECT 285.725 2058.040 300.380 2058.170 ;
        RECT 285.725 2057.870 304.000 2058.040 ;
        RECT 285.725 2057.855 286.055 2057.870 ;
        RECT 300.000 2057.440 304.000 2057.870 ;
        RECT -4.800 897.410 2.400 897.860 ;
        RECT 16.165 897.410 16.495 897.425 ;
        RECT -4.800 897.110 16.495 897.410 ;
        RECT -4.800 896.660 2.400 897.110 ;
        RECT 16.165 897.095 16.495 897.110 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 168.890 2084.100 169.210 2084.160 ;
        RECT 285.730 2084.100 286.050 2084.160 ;
        RECT 168.890 2083.960 286.050 2084.100 ;
        RECT 168.890 2083.900 169.210 2083.960 ;
        RECT 285.730 2083.900 286.050 2083.960 ;
        RECT 16.170 682.960 16.490 683.020 ;
        RECT 168.890 682.960 169.210 683.020 ;
        RECT 16.170 682.820 169.210 682.960 ;
        RECT 16.170 682.760 16.490 682.820 ;
        RECT 168.890 682.760 169.210 682.820 ;
      LAYER via ;
        RECT 168.920 2083.900 169.180 2084.160 ;
        RECT 285.760 2083.900 286.020 2084.160 ;
        RECT 16.200 682.760 16.460 683.020 ;
        RECT 168.920 682.760 169.180 683.020 ;
      LAYER met2 ;
        RECT 285.750 2089.115 286.030 2089.485 ;
        RECT 285.820 2084.190 285.960 2089.115 ;
        RECT 168.920 2083.870 169.180 2084.190 ;
        RECT 285.760 2083.870 286.020 2084.190 ;
        RECT 168.980 683.050 169.120 2083.870 ;
        RECT 16.200 682.730 16.460 683.050 ;
        RECT 168.920 682.730 169.180 683.050 ;
        RECT 16.260 681.885 16.400 682.730 ;
        RECT 16.190 681.515 16.470 681.885 ;
      LAYER via2 ;
        RECT 285.750 2089.160 286.030 2089.440 ;
        RECT 16.190 681.560 16.470 681.840 ;
      LAYER met3 ;
        RECT 285.725 2089.450 286.055 2089.465 ;
        RECT 285.725 2089.320 300.380 2089.450 ;
        RECT 285.725 2089.150 304.000 2089.320 ;
        RECT 285.725 2089.135 286.055 2089.150 ;
        RECT 300.000 2088.720 304.000 2089.150 ;
        RECT -4.800 681.850 2.400 682.300 ;
        RECT 16.165 681.850 16.495 681.865 ;
        RECT -4.800 681.550 16.495 681.850 ;
        RECT -4.800 681.100 2.400 681.550 ;
        RECT 16.165 681.535 16.495 681.550 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 217.190 2118.440 217.510 2118.500 ;
        RECT 285.730 2118.440 286.050 2118.500 ;
        RECT 217.190 2118.300 286.050 2118.440 ;
        RECT 217.190 2118.240 217.510 2118.300 ;
        RECT 285.730 2118.240 286.050 2118.300 ;
        RECT 17.090 469.100 17.410 469.160 ;
        RECT 217.190 469.100 217.510 469.160 ;
        RECT 17.090 468.960 217.510 469.100 ;
        RECT 17.090 468.900 17.410 468.960 ;
        RECT 217.190 468.900 217.510 468.960 ;
      LAYER via ;
        RECT 217.220 2118.240 217.480 2118.500 ;
        RECT 285.760 2118.240 286.020 2118.500 ;
        RECT 17.120 468.900 17.380 469.160 ;
        RECT 217.220 468.900 217.480 469.160 ;
      LAYER met2 ;
        RECT 285.750 2121.075 286.030 2121.445 ;
        RECT 285.820 2118.530 285.960 2121.075 ;
        RECT 217.220 2118.210 217.480 2118.530 ;
        RECT 285.760 2118.210 286.020 2118.530 ;
        RECT 217.280 469.190 217.420 2118.210 ;
        RECT 17.120 468.870 17.380 469.190 ;
        RECT 217.220 468.870 217.480 469.190 ;
        RECT 17.180 466.325 17.320 468.870 ;
        RECT 17.110 465.955 17.390 466.325 ;
      LAYER via2 ;
        RECT 285.750 2121.120 286.030 2121.400 ;
        RECT 17.110 466.000 17.390 466.280 ;
      LAYER met3 ;
        RECT 285.725 2121.410 286.055 2121.425 ;
        RECT 285.725 2121.280 300.380 2121.410 ;
        RECT 285.725 2121.110 304.000 2121.280 ;
        RECT 285.725 2121.095 286.055 2121.110 ;
        RECT 300.000 2120.680 304.000 2121.110 ;
        RECT -4.800 466.290 2.400 466.740 ;
        RECT 17.085 466.290 17.415 466.305 ;
        RECT -4.800 465.990 17.415 466.290 ;
        RECT -4.800 465.540 2.400 465.990 ;
        RECT 17.085 465.975 17.415 465.990 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 230.990 2145.980 231.310 2146.040 ;
        RECT 285.730 2145.980 286.050 2146.040 ;
        RECT 230.990 2145.840 286.050 2145.980 ;
        RECT 230.990 2145.780 231.310 2145.840 ;
        RECT 285.730 2145.780 286.050 2145.840 ;
        RECT 17.090 255.240 17.410 255.300 ;
        RECT 230.990 255.240 231.310 255.300 ;
        RECT 17.090 255.100 231.310 255.240 ;
        RECT 17.090 255.040 17.410 255.100 ;
        RECT 230.990 255.040 231.310 255.100 ;
      LAYER via ;
        RECT 231.020 2145.780 231.280 2146.040 ;
        RECT 285.760 2145.780 286.020 2146.040 ;
        RECT 17.120 255.040 17.380 255.300 ;
        RECT 231.020 255.040 231.280 255.300 ;
      LAYER met2 ;
        RECT 285.750 2152.355 286.030 2152.725 ;
        RECT 285.820 2146.070 285.960 2152.355 ;
        RECT 231.020 2145.750 231.280 2146.070 ;
        RECT 285.760 2145.750 286.020 2146.070 ;
        RECT 231.080 255.330 231.220 2145.750 ;
        RECT 17.120 255.010 17.380 255.330 ;
        RECT 231.020 255.010 231.280 255.330 ;
        RECT 17.180 250.765 17.320 255.010 ;
        RECT 17.110 250.395 17.390 250.765 ;
      LAYER via2 ;
        RECT 285.750 2152.400 286.030 2152.680 ;
        RECT 17.110 250.440 17.390 250.720 ;
      LAYER met3 ;
        RECT 285.725 2152.690 286.055 2152.705 ;
        RECT 285.725 2152.560 300.380 2152.690 ;
        RECT 285.725 2152.390 304.000 2152.560 ;
        RECT 285.725 2152.375 286.055 2152.390 ;
        RECT 300.000 2151.960 304.000 2152.390 ;
        RECT -4.800 250.730 2.400 251.180 ;
        RECT 17.085 250.730 17.415 250.745 ;
        RECT -4.800 250.430 17.415 250.730 ;
        RECT -4.800 249.980 2.400 250.430 ;
        RECT 17.085 250.415 17.415 250.430 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 258.590 2180.660 258.910 2180.720 ;
        RECT 282.970 2180.660 283.290 2180.720 ;
        RECT 258.590 2180.520 283.290 2180.660 ;
        RECT 258.590 2180.460 258.910 2180.520 ;
        RECT 282.970 2180.460 283.290 2180.520 ;
        RECT 17.090 41.380 17.410 41.440 ;
        RECT 258.590 41.380 258.910 41.440 ;
        RECT 17.090 41.240 258.910 41.380 ;
        RECT 17.090 41.180 17.410 41.240 ;
        RECT 258.590 41.180 258.910 41.240 ;
      LAYER via ;
        RECT 258.620 2180.460 258.880 2180.720 ;
        RECT 283.000 2180.460 283.260 2180.720 ;
        RECT 17.120 41.180 17.380 41.440 ;
        RECT 258.620 41.180 258.880 41.440 ;
      LAYER met2 ;
        RECT 258.620 2180.430 258.880 2180.750 ;
        RECT 283.000 2180.605 283.260 2180.750 ;
        RECT 258.680 41.470 258.820 2180.430 ;
        RECT 282.990 2180.235 283.270 2180.605 ;
        RECT 17.120 41.150 17.380 41.470 ;
        RECT 258.620 41.150 258.880 41.470 ;
        RECT 17.180 35.885 17.320 41.150 ;
        RECT 17.110 35.515 17.390 35.885 ;
      LAYER via2 ;
        RECT 282.990 2180.280 283.270 2180.560 ;
        RECT 17.110 35.560 17.390 35.840 ;
      LAYER met3 ;
        RECT 300.000 2183.920 304.000 2184.520 ;
        RECT 282.965 2180.570 283.295 2180.585 ;
        RECT 300.230 2180.570 300.530 2183.920 ;
        RECT 282.965 2180.270 300.530 2180.570 ;
        RECT 282.965 2180.255 283.295 2180.270 ;
        RECT -4.800 35.850 2.400 36.300 ;
        RECT 17.085 35.850 17.415 35.865 ;
        RECT -4.800 35.550 17.415 35.850 ;
        RECT -4.800 35.100 2.400 35.550 ;
        RECT 17.085 35.535 17.415 35.550 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 286.650 910.760 286.970 910.820 ;
        RECT 2900.830 910.760 2901.150 910.820 ;
        RECT 286.650 910.620 2901.150 910.760 ;
        RECT 286.650 910.560 286.970 910.620 ;
        RECT 2900.830 910.560 2901.150 910.620 ;
      LAYER via ;
        RECT 286.680 910.560 286.940 910.820 ;
        RECT 2900.860 910.560 2901.120 910.820 ;
      LAYER met2 ;
        RECT 286.670 1109.915 286.950 1110.285 ;
        RECT 286.740 910.850 286.880 1109.915 ;
        RECT 286.680 910.530 286.940 910.850 ;
        RECT 2900.860 910.530 2901.120 910.850 ;
        RECT 2900.920 909.685 2901.060 910.530 ;
        RECT 2900.850 909.315 2901.130 909.685 ;
      LAYER via2 ;
        RECT 286.670 1109.960 286.950 1110.240 ;
        RECT 2900.850 909.360 2901.130 909.640 ;
      LAYER met3 ;
        RECT 286.645 1110.250 286.975 1110.265 ;
        RECT 286.645 1110.120 300.380 1110.250 ;
        RECT 286.645 1109.950 304.000 1110.120 ;
        RECT 286.645 1109.935 286.975 1109.950 ;
        RECT 300.000 1109.520 304.000 1109.950 ;
        RECT 2900.825 909.650 2901.155 909.665 ;
        RECT 2917.600 909.650 2924.800 910.100 ;
        RECT 2900.825 909.350 2924.800 909.650 ;
        RECT 2900.825 909.335 2901.155 909.350 ;
        RECT 2917.600 908.900 2924.800 909.350 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 287.570 1007.320 287.890 1007.380 ;
        RECT 288.950 1007.320 289.270 1007.380 ;
        RECT 287.570 1007.180 289.270 1007.320 ;
        RECT 287.570 1007.120 287.890 1007.180 ;
        RECT 288.950 1007.120 289.270 1007.180 ;
        RECT 287.570 1002.900 287.890 1002.960 ;
        RECT 2900.370 1002.900 2900.690 1002.960 ;
        RECT 287.570 1002.760 2900.690 1002.900 ;
        RECT 287.570 1002.700 287.890 1002.760 ;
        RECT 2900.370 1002.700 2900.690 1002.760 ;
      LAYER via ;
        RECT 287.600 1007.120 287.860 1007.380 ;
        RECT 288.980 1007.120 289.240 1007.380 ;
        RECT 287.600 1002.700 287.860 1002.960 ;
        RECT 2900.400 1002.700 2900.660 1002.960 ;
      LAYER met2 ;
        RECT 2900.390 1143.915 2900.670 1144.285 ;
        RECT 288.970 1141.875 289.250 1142.245 ;
        RECT 289.040 1007.410 289.180 1141.875 ;
        RECT 287.600 1007.090 287.860 1007.410 ;
        RECT 288.980 1007.090 289.240 1007.410 ;
        RECT 287.660 1002.990 287.800 1007.090 ;
        RECT 2900.460 1002.990 2900.600 1143.915 ;
        RECT 287.600 1002.670 287.860 1002.990 ;
        RECT 2900.400 1002.670 2900.660 1002.990 ;
      LAYER via2 ;
        RECT 2900.390 1143.960 2900.670 1144.240 ;
        RECT 288.970 1141.920 289.250 1142.200 ;
      LAYER met3 ;
        RECT 2900.365 1144.250 2900.695 1144.265 ;
        RECT 2917.600 1144.250 2924.800 1144.700 ;
        RECT 2900.365 1143.950 2924.800 1144.250 ;
        RECT 2900.365 1143.935 2900.695 1143.950 ;
        RECT 2917.600 1143.500 2924.800 1143.950 ;
        RECT 288.945 1142.210 289.275 1142.225 ;
        RECT 288.945 1142.080 300.380 1142.210 ;
        RECT 288.945 1141.910 304.000 1142.080 ;
        RECT 288.945 1141.895 289.275 1141.910 ;
        RECT 300.000 1141.480 304.000 1141.910 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 285.270 1004.260 285.590 1004.320 ;
        RECT 2904.050 1004.260 2904.370 1004.320 ;
        RECT 285.270 1004.120 2904.370 1004.260 ;
        RECT 285.270 1004.060 285.590 1004.120 ;
        RECT 2904.050 1004.060 2904.370 1004.120 ;
      LAYER via ;
        RECT 285.300 1004.060 285.560 1004.320 ;
        RECT 2904.080 1004.060 2904.340 1004.320 ;
      LAYER met2 ;
        RECT 2904.070 1378.515 2904.350 1378.885 ;
        RECT 285.750 1173.155 286.030 1173.525 ;
        RECT 285.820 1026.530 285.960 1173.155 ;
        RECT 285.360 1026.390 285.960 1026.530 ;
        RECT 285.360 1004.350 285.500 1026.390 ;
        RECT 2904.140 1004.350 2904.280 1378.515 ;
        RECT 285.300 1004.030 285.560 1004.350 ;
        RECT 2904.080 1004.030 2904.340 1004.350 ;
      LAYER via2 ;
        RECT 2904.070 1378.560 2904.350 1378.840 ;
        RECT 285.750 1173.200 286.030 1173.480 ;
      LAYER met3 ;
        RECT 2904.045 1378.850 2904.375 1378.865 ;
        RECT 2917.600 1378.850 2924.800 1379.300 ;
        RECT 2904.045 1378.550 2924.800 1378.850 ;
        RECT 2904.045 1378.535 2904.375 1378.550 ;
        RECT 2917.600 1378.100 2924.800 1378.550 ;
        RECT 285.725 1173.490 286.055 1173.505 ;
        RECT 285.725 1173.360 300.380 1173.490 ;
        RECT 285.725 1173.190 304.000 1173.360 ;
        RECT 285.725 1173.175 286.055 1173.190 ;
        RECT 300.000 1172.760 304.000 1173.190 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 288.490 1003.580 288.810 1003.640 ;
        RECT 2902.670 1003.580 2902.990 1003.640 ;
        RECT 288.490 1003.440 2902.990 1003.580 ;
        RECT 288.490 1003.380 288.810 1003.440 ;
        RECT 2902.670 1003.380 2902.990 1003.440 ;
      LAYER via ;
        RECT 288.520 1003.380 288.780 1003.640 ;
        RECT 2902.700 1003.380 2902.960 1003.640 ;
      LAYER met2 ;
        RECT 2902.690 1613.115 2902.970 1613.485 ;
        RECT 288.510 1205.115 288.790 1205.485 ;
        RECT 288.580 1003.670 288.720 1205.115 ;
        RECT 2902.760 1003.670 2902.900 1613.115 ;
        RECT 288.520 1003.350 288.780 1003.670 ;
        RECT 2902.700 1003.350 2902.960 1003.670 ;
      LAYER via2 ;
        RECT 2902.690 1613.160 2902.970 1613.440 ;
        RECT 288.510 1205.160 288.790 1205.440 ;
      LAYER met3 ;
        RECT 2902.665 1613.450 2902.995 1613.465 ;
        RECT 2917.600 1613.450 2924.800 1613.900 ;
        RECT 2902.665 1613.150 2924.800 1613.450 ;
        RECT 2902.665 1613.135 2902.995 1613.150 ;
        RECT 2917.600 1612.700 2924.800 1613.150 ;
        RECT 288.485 1205.450 288.815 1205.465 ;
        RECT 288.485 1205.320 300.380 1205.450 ;
        RECT 288.485 1205.150 304.000 1205.320 ;
        RECT 288.485 1205.135 288.815 1205.150 ;
        RECT 300.000 1204.720 304.000 1205.150 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2901.310 1847.715 2901.590 1848.085 ;
        RECT 2901.380 1003.525 2901.520 1847.715 ;
        RECT 2901.310 1003.155 2901.590 1003.525 ;
      LAYER via2 ;
        RECT 2901.310 1847.760 2901.590 1848.040 ;
        RECT 2901.310 1003.200 2901.590 1003.480 ;
      LAYER met3 ;
        RECT 2901.285 1848.050 2901.615 1848.065 ;
        RECT 2917.600 1848.050 2924.800 1848.500 ;
        RECT 2901.285 1847.750 2924.800 1848.050 ;
        RECT 2901.285 1847.735 2901.615 1847.750 ;
        RECT 2917.600 1847.300 2924.800 1847.750 ;
        RECT 289.150 1236.730 289.530 1236.740 ;
        RECT 289.150 1236.600 300.380 1236.730 ;
        RECT 289.150 1236.430 304.000 1236.600 ;
        RECT 289.150 1236.420 289.530 1236.430 ;
        RECT 300.000 1236.000 304.000 1236.430 ;
        RECT 289.150 1003.490 289.530 1003.500 ;
        RECT 2901.285 1003.490 2901.615 1003.505 ;
        RECT 289.150 1003.190 2901.615 1003.490 ;
        RECT 289.150 1003.180 289.530 1003.190 ;
        RECT 2901.285 1003.175 2901.615 1003.190 ;
      LAYER via3 ;
        RECT 289.180 1236.420 289.500 1236.740 ;
        RECT 289.180 1003.180 289.500 1003.500 ;
      LAYER met4 ;
        RECT 289.175 1236.415 289.505 1236.745 ;
        RECT 289.190 1003.505 289.490 1236.415 ;
        RECT 289.175 1003.175 289.505 1003.505 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 287.110 2189.840 287.430 2189.900 ;
        RECT 2902.210 2189.840 2902.530 2189.900 ;
        RECT 287.110 2189.700 2902.530 2189.840 ;
        RECT 287.110 2189.640 287.430 2189.700 ;
        RECT 2902.210 2189.640 2902.530 2189.700 ;
      LAYER via ;
        RECT 287.140 2189.640 287.400 2189.900 ;
        RECT 2902.240 2189.640 2902.500 2189.900 ;
      LAYER met2 ;
        RECT 287.140 2189.610 287.400 2189.930 ;
        RECT 2902.240 2189.610 2902.500 2189.930 ;
        RECT 287.200 1268.725 287.340 2189.610 ;
        RECT 2902.300 2082.685 2902.440 2189.610 ;
        RECT 2902.230 2082.315 2902.510 2082.685 ;
        RECT 287.130 1268.355 287.410 1268.725 ;
      LAYER via2 ;
        RECT 2902.230 2082.360 2902.510 2082.640 ;
        RECT 287.130 1268.400 287.410 1268.680 ;
      LAYER met3 ;
        RECT 2902.205 2082.650 2902.535 2082.665 ;
        RECT 2917.600 2082.650 2924.800 2083.100 ;
        RECT 2902.205 2082.350 2924.800 2082.650 ;
        RECT 2902.205 2082.335 2902.535 2082.350 ;
        RECT 2917.600 2081.900 2924.800 2082.350 ;
        RECT 287.105 1268.690 287.435 1268.705 ;
        RECT 287.105 1268.560 300.380 1268.690 ;
        RECT 287.105 1268.390 304.000 1268.560 ;
        RECT 287.105 1268.375 287.435 1268.390 ;
        RECT 300.000 1267.960 304.000 1268.390 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 286.650 2191.200 286.970 2191.260 ;
        RECT 2904.050 2191.200 2904.370 2191.260 ;
        RECT 286.650 2191.060 2904.370 2191.200 ;
        RECT 286.650 2191.000 286.970 2191.060 ;
        RECT 2904.050 2191.000 2904.370 2191.060 ;
      LAYER via ;
        RECT 286.680 2191.000 286.940 2191.260 ;
        RECT 2904.080 2191.000 2904.340 2191.260 ;
      LAYER met2 ;
        RECT 2904.070 2316.915 2904.350 2317.285 ;
        RECT 2904.140 2191.290 2904.280 2316.915 ;
        RECT 286.680 2190.970 286.940 2191.290 ;
        RECT 2904.080 2190.970 2904.340 2191.290 ;
        RECT 286.740 1300.005 286.880 2190.970 ;
        RECT 286.670 1299.635 286.950 1300.005 ;
      LAYER via2 ;
        RECT 2904.070 2316.960 2904.350 2317.240 ;
        RECT 286.670 1299.680 286.950 1299.960 ;
      LAYER met3 ;
        RECT 2904.045 2317.250 2904.375 2317.265 ;
        RECT 2917.600 2317.250 2924.800 2317.700 ;
        RECT 2904.045 2316.950 2924.800 2317.250 ;
        RECT 2904.045 2316.935 2904.375 2316.950 ;
        RECT 2917.600 2316.500 2924.800 2316.950 ;
        RECT 286.645 1299.970 286.975 1299.985 ;
        RECT 286.645 1299.840 300.380 1299.970 ;
        RECT 286.645 1299.670 304.000 1299.840 ;
        RECT 286.645 1299.655 286.975 1299.670 ;
        RECT 300.000 1299.240 304.000 1299.670 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 448.110 146.780 448.430 146.840 ;
        RECT 482.610 146.780 482.930 146.840 ;
        RECT 448.110 146.640 482.930 146.780 ;
        RECT 448.110 146.580 448.430 146.640 ;
        RECT 482.610 146.580 482.930 146.640 ;
        RECT 580.130 145.420 580.450 145.480 ;
        RECT 604.050 145.420 604.370 145.480 ;
        RECT 580.130 145.280 604.370 145.420 ;
        RECT 580.130 145.220 580.450 145.280 ;
        RECT 604.050 145.220 604.370 145.280 ;
        RECT 725.030 145.420 725.350 145.480 ;
        RECT 772.410 145.420 772.730 145.480 ;
        RECT 725.030 145.280 772.730 145.420 ;
        RECT 725.030 145.220 725.350 145.280 ;
        RECT 772.410 145.220 772.730 145.280 ;
      LAYER via ;
        RECT 448.140 146.580 448.400 146.840 ;
        RECT 482.640 146.580 482.900 146.840 ;
        RECT 580.160 145.220 580.420 145.480 ;
        RECT 604.080 145.220 604.340 145.480 ;
        RECT 725.060 145.220 725.320 145.480 ;
        RECT 772.440 145.220 772.700 145.480 ;
      LAYER met2 ;
        RECT 717.230 147.035 717.510 147.405 ;
        RECT 448.140 146.725 448.400 146.870 ;
        RECT 482.640 146.725 482.900 146.870 ;
        RECT 448.130 146.355 448.410 146.725 ;
        RECT 482.630 146.355 482.910 146.725 ;
        RECT 604.070 146.355 604.350 146.725 ;
        RECT 640.870 146.610 641.150 146.725 ;
        RECT 641.790 146.610 642.070 146.725 ;
        RECT 640.870 146.470 642.070 146.610 ;
        RECT 640.870 146.355 641.150 146.470 ;
        RECT 641.790 146.355 642.070 146.470 ;
        RECT 604.140 145.510 604.280 146.355 ;
        RECT 580.160 145.365 580.420 145.510 ;
        RECT 580.150 144.995 580.430 145.365 ;
        RECT 604.080 145.190 604.340 145.510 ;
        RECT 717.300 145.365 717.440 147.035 ;
        RECT 772.430 146.355 772.710 146.725 ;
        RECT 772.500 145.510 772.640 146.355 ;
        RECT 725.060 145.365 725.320 145.510 ;
        RECT 717.230 144.995 717.510 145.365 ;
        RECT 725.050 144.995 725.330 145.365 ;
        RECT 772.440 145.190 772.700 145.510 ;
      LAYER via2 ;
        RECT 717.230 147.080 717.510 147.360 ;
        RECT 448.130 146.400 448.410 146.680 ;
        RECT 482.630 146.400 482.910 146.680 ;
        RECT 604.070 146.400 604.350 146.680 ;
        RECT 640.870 146.400 641.150 146.680 ;
        RECT 641.790 146.400 642.070 146.680 ;
        RECT 580.150 145.040 580.430 145.320 ;
        RECT 772.430 146.400 772.710 146.680 ;
        RECT 717.230 145.040 717.510 145.320 ;
        RECT 725.050 145.040 725.330 145.320 ;
      LAYER met3 ;
        RECT 283.630 1025.930 284.010 1025.940 ;
        RECT 283.630 1025.800 300.380 1025.930 ;
        RECT 283.630 1025.630 304.000 1025.800 ;
        RECT 283.630 1025.620 284.010 1025.630 ;
        RECT 300.000 1025.200 304.000 1025.630 ;
        RECT 578.950 147.370 579.330 147.380 ;
        RECT 544.030 147.070 579.330 147.370 ;
        RECT 283.630 146.690 284.010 146.700 ;
        RECT 448.105 146.690 448.435 146.705 ;
        RECT 283.630 146.390 324.450 146.690 ;
        RECT 283.630 146.380 284.010 146.390 ;
        RECT 324.150 146.010 324.450 146.390 ;
        RECT 372.910 146.390 448.435 146.690 ;
        RECT 324.150 145.710 372.290 146.010 ;
        RECT 371.990 145.330 372.290 145.710 ;
        RECT 372.910 145.330 373.210 146.390 ;
        RECT 448.105 146.375 448.435 146.390 ;
        RECT 482.605 146.690 482.935 146.705 ;
        RECT 482.605 146.390 496.490 146.690 ;
        RECT 482.605 146.375 482.935 146.390 ;
        RECT 371.990 145.030 373.210 145.330 ;
        RECT 496.190 145.330 496.490 146.390 ;
        RECT 544.030 146.010 544.330 147.070 ;
        RECT 578.950 147.060 579.330 147.070 ;
        RECT 669.110 147.370 669.490 147.380 ;
        RECT 717.205 147.370 717.535 147.385 ;
        RECT 669.110 147.070 717.535 147.370 ;
        RECT 669.110 147.060 669.490 147.070 ;
        RECT 717.205 147.055 717.535 147.070 ;
        RECT 604.045 146.690 604.375 146.705 ;
        RECT 640.845 146.690 641.175 146.705 ;
        RECT 604.045 146.390 641.175 146.690 ;
        RECT 604.045 146.375 604.375 146.390 ;
        RECT 640.845 146.375 641.175 146.390 ;
        RECT 641.765 146.690 642.095 146.705 ;
        RECT 772.405 146.690 772.735 146.705 ;
        RECT 2917.600 146.690 2924.800 147.140 ;
        RECT 641.765 146.390 651.970 146.690 ;
        RECT 641.765 146.375 642.095 146.390 ;
        RECT 497.110 145.710 544.330 146.010 ;
        RECT 651.670 146.010 651.970 146.390 ;
        RECT 772.405 146.390 807.450 146.690 ;
        RECT 772.405 146.375 772.735 146.390 ;
        RECT 669.110 146.010 669.490 146.020 ;
        RECT 651.670 145.710 669.490 146.010 ;
        RECT 807.150 146.010 807.450 146.390 ;
        RECT 855.910 146.390 904.050 146.690 ;
        RECT 807.150 145.710 855.290 146.010 ;
        RECT 497.110 145.330 497.410 145.710 ;
        RECT 669.110 145.700 669.490 145.710 ;
        RECT 496.190 145.030 497.410 145.330 ;
        RECT 578.950 145.330 579.330 145.340 ;
        RECT 580.125 145.330 580.455 145.345 ;
        RECT 578.950 145.030 580.455 145.330 ;
        RECT 578.950 145.020 579.330 145.030 ;
        RECT 580.125 145.015 580.455 145.030 ;
        RECT 717.205 145.330 717.535 145.345 ;
        RECT 725.025 145.330 725.355 145.345 ;
        RECT 717.205 145.030 725.355 145.330 ;
        RECT 854.990 145.330 855.290 145.710 ;
        RECT 855.910 145.330 856.210 146.390 ;
        RECT 903.750 146.010 904.050 146.390 ;
        RECT 952.510 146.390 1000.650 146.690 ;
        RECT 903.750 145.710 951.890 146.010 ;
        RECT 854.990 145.030 856.210 145.330 ;
        RECT 951.590 145.330 951.890 145.710 ;
        RECT 952.510 145.330 952.810 146.390 ;
        RECT 1000.350 146.010 1000.650 146.390 ;
        RECT 1049.110 146.390 1097.250 146.690 ;
        RECT 1000.350 145.710 1048.490 146.010 ;
        RECT 951.590 145.030 952.810 145.330 ;
        RECT 1048.190 145.330 1048.490 145.710 ;
        RECT 1049.110 145.330 1049.410 146.390 ;
        RECT 1096.950 146.010 1097.250 146.390 ;
        RECT 1145.710 146.390 1193.850 146.690 ;
        RECT 1096.950 145.710 1145.090 146.010 ;
        RECT 1048.190 145.030 1049.410 145.330 ;
        RECT 1144.790 145.330 1145.090 145.710 ;
        RECT 1145.710 145.330 1146.010 146.390 ;
        RECT 1193.550 146.010 1193.850 146.390 ;
        RECT 1242.310 146.390 1290.450 146.690 ;
        RECT 1193.550 145.710 1241.690 146.010 ;
        RECT 1144.790 145.030 1146.010 145.330 ;
        RECT 1241.390 145.330 1241.690 145.710 ;
        RECT 1242.310 145.330 1242.610 146.390 ;
        RECT 1290.150 146.010 1290.450 146.390 ;
        RECT 1338.910 146.390 1387.050 146.690 ;
        RECT 1290.150 145.710 1338.290 146.010 ;
        RECT 1241.390 145.030 1242.610 145.330 ;
        RECT 1337.990 145.330 1338.290 145.710 ;
        RECT 1338.910 145.330 1339.210 146.390 ;
        RECT 1386.750 146.010 1387.050 146.390 ;
        RECT 1435.510 146.390 1483.650 146.690 ;
        RECT 1386.750 145.710 1434.890 146.010 ;
        RECT 1337.990 145.030 1339.210 145.330 ;
        RECT 1434.590 145.330 1434.890 145.710 ;
        RECT 1435.510 145.330 1435.810 146.390 ;
        RECT 1483.350 146.010 1483.650 146.390 ;
        RECT 1532.110 146.390 1580.250 146.690 ;
        RECT 1483.350 145.710 1531.490 146.010 ;
        RECT 1434.590 145.030 1435.810 145.330 ;
        RECT 1531.190 145.330 1531.490 145.710 ;
        RECT 1532.110 145.330 1532.410 146.390 ;
        RECT 1579.950 146.010 1580.250 146.390 ;
        RECT 1628.710 146.390 1676.850 146.690 ;
        RECT 1579.950 145.710 1628.090 146.010 ;
        RECT 1531.190 145.030 1532.410 145.330 ;
        RECT 1627.790 145.330 1628.090 145.710 ;
        RECT 1628.710 145.330 1629.010 146.390 ;
        RECT 1676.550 146.010 1676.850 146.390 ;
        RECT 1725.310 146.390 1773.450 146.690 ;
        RECT 1676.550 145.710 1724.690 146.010 ;
        RECT 1627.790 145.030 1629.010 145.330 ;
        RECT 1724.390 145.330 1724.690 145.710 ;
        RECT 1725.310 145.330 1725.610 146.390 ;
        RECT 1773.150 146.010 1773.450 146.390 ;
        RECT 1821.910 146.390 1870.050 146.690 ;
        RECT 1773.150 145.710 1821.290 146.010 ;
        RECT 1724.390 145.030 1725.610 145.330 ;
        RECT 1820.990 145.330 1821.290 145.710 ;
        RECT 1821.910 145.330 1822.210 146.390 ;
        RECT 1869.750 146.010 1870.050 146.390 ;
        RECT 1918.510 146.390 1966.650 146.690 ;
        RECT 1869.750 145.710 1917.890 146.010 ;
        RECT 1820.990 145.030 1822.210 145.330 ;
        RECT 1917.590 145.330 1917.890 145.710 ;
        RECT 1918.510 145.330 1918.810 146.390 ;
        RECT 1966.350 146.010 1966.650 146.390 ;
        RECT 2015.110 146.390 2063.250 146.690 ;
        RECT 1966.350 145.710 2014.490 146.010 ;
        RECT 1917.590 145.030 1918.810 145.330 ;
        RECT 2014.190 145.330 2014.490 145.710 ;
        RECT 2015.110 145.330 2015.410 146.390 ;
        RECT 2062.950 146.010 2063.250 146.390 ;
        RECT 2111.710 146.390 2159.850 146.690 ;
        RECT 2062.950 145.710 2111.090 146.010 ;
        RECT 2014.190 145.030 2015.410 145.330 ;
        RECT 2110.790 145.330 2111.090 145.710 ;
        RECT 2111.710 145.330 2112.010 146.390 ;
        RECT 2159.550 146.010 2159.850 146.390 ;
        RECT 2208.310 146.390 2256.450 146.690 ;
        RECT 2159.550 145.710 2207.690 146.010 ;
        RECT 2110.790 145.030 2112.010 145.330 ;
        RECT 2207.390 145.330 2207.690 145.710 ;
        RECT 2208.310 145.330 2208.610 146.390 ;
        RECT 2256.150 146.010 2256.450 146.390 ;
        RECT 2304.910 146.390 2353.050 146.690 ;
        RECT 2256.150 145.710 2304.290 146.010 ;
        RECT 2207.390 145.030 2208.610 145.330 ;
        RECT 2303.990 145.330 2304.290 145.710 ;
        RECT 2304.910 145.330 2305.210 146.390 ;
        RECT 2352.750 146.010 2353.050 146.390 ;
        RECT 2401.510 146.390 2449.650 146.690 ;
        RECT 2352.750 145.710 2400.890 146.010 ;
        RECT 2303.990 145.030 2305.210 145.330 ;
        RECT 2400.590 145.330 2400.890 145.710 ;
        RECT 2401.510 145.330 2401.810 146.390 ;
        RECT 2449.350 146.010 2449.650 146.390 ;
        RECT 2498.110 146.390 2546.250 146.690 ;
        RECT 2449.350 145.710 2497.490 146.010 ;
        RECT 2400.590 145.030 2401.810 145.330 ;
        RECT 2497.190 145.330 2497.490 145.710 ;
        RECT 2498.110 145.330 2498.410 146.390 ;
        RECT 2545.950 146.010 2546.250 146.390 ;
        RECT 2594.710 146.390 2642.850 146.690 ;
        RECT 2545.950 145.710 2594.090 146.010 ;
        RECT 2497.190 145.030 2498.410 145.330 ;
        RECT 2593.790 145.330 2594.090 145.710 ;
        RECT 2594.710 145.330 2595.010 146.390 ;
        RECT 2642.550 146.010 2642.850 146.390 ;
        RECT 2691.310 146.390 2739.450 146.690 ;
        RECT 2642.550 145.710 2690.690 146.010 ;
        RECT 2593.790 145.030 2595.010 145.330 ;
        RECT 2690.390 145.330 2690.690 145.710 ;
        RECT 2691.310 145.330 2691.610 146.390 ;
        RECT 2739.150 146.010 2739.450 146.390 ;
        RECT 2787.910 146.390 2836.050 146.690 ;
        RECT 2739.150 145.710 2787.290 146.010 ;
        RECT 2690.390 145.030 2691.610 145.330 ;
        RECT 2786.990 145.330 2787.290 145.710 ;
        RECT 2787.910 145.330 2788.210 146.390 ;
        RECT 2835.750 146.010 2836.050 146.390 ;
        RECT 2916.710 146.390 2924.800 146.690 ;
        RECT 2916.710 146.010 2917.010 146.390 ;
        RECT 2835.750 145.710 2883.890 146.010 ;
        RECT 2786.990 145.030 2788.210 145.330 ;
        RECT 2883.590 145.330 2883.890 145.710 ;
        RECT 2884.510 145.710 2917.010 146.010 ;
        RECT 2917.600 145.940 2924.800 146.390 ;
        RECT 2884.510 145.330 2884.810 145.710 ;
        RECT 2883.590 145.030 2884.810 145.330 ;
        RECT 717.205 145.015 717.535 145.030 ;
        RECT 725.025 145.015 725.355 145.030 ;
      LAYER via3 ;
        RECT 283.660 1025.620 283.980 1025.940 ;
        RECT 283.660 146.380 283.980 146.700 ;
        RECT 578.980 147.060 579.300 147.380 ;
        RECT 669.140 147.060 669.460 147.380 ;
        RECT 669.140 145.700 669.460 146.020 ;
        RECT 578.980 145.020 579.300 145.340 ;
      LAYER met4 ;
        RECT 283.655 1025.615 283.985 1025.945 ;
        RECT 283.670 146.705 283.970 1025.615 ;
        RECT 578.975 147.055 579.305 147.385 ;
        RECT 669.135 147.055 669.465 147.385 ;
        RECT 283.655 146.375 283.985 146.705 ;
        RECT 578.990 145.345 579.290 147.055 ;
        RECT 669.150 146.025 669.450 147.055 ;
        RECT 669.135 145.695 669.465 146.025 ;
        RECT 578.975 145.015 579.305 145.345 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 286.190 2191.540 286.510 2191.600 ;
        RECT 2902.670 2191.540 2902.990 2191.600 ;
        RECT 286.190 2191.400 2902.990 2191.540 ;
        RECT 286.190 2191.340 286.510 2191.400 ;
        RECT 2902.670 2191.340 2902.990 2191.400 ;
      LAYER via ;
        RECT 286.220 2191.340 286.480 2191.600 ;
        RECT 2902.700 2191.340 2902.960 2191.600 ;
      LAYER met2 ;
        RECT 2902.690 2493.035 2902.970 2493.405 ;
        RECT 2902.760 2191.630 2902.900 2493.035 ;
        RECT 286.220 2191.310 286.480 2191.630 ;
        RECT 2902.700 2191.310 2902.960 2191.630 ;
        RECT 286.280 1342.165 286.420 2191.310 ;
        RECT 286.210 1341.795 286.490 1342.165 ;
      LAYER via2 ;
        RECT 2902.690 2493.080 2902.970 2493.360 ;
        RECT 286.210 1341.840 286.490 1342.120 ;
      LAYER met3 ;
        RECT 2902.665 2493.370 2902.995 2493.385 ;
        RECT 2917.600 2493.370 2924.800 2493.820 ;
        RECT 2902.665 2493.070 2924.800 2493.370 ;
        RECT 2902.665 2493.055 2902.995 2493.070 ;
        RECT 2917.600 2492.620 2924.800 2493.070 ;
        RECT 286.185 1342.130 286.515 1342.145 ;
        RECT 286.185 1342.000 300.380 1342.130 ;
        RECT 286.185 1341.830 304.000 1342.000 ;
        RECT 286.185 1341.815 286.515 1341.830 ;
        RECT 300.000 1341.400 304.000 1341.830 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 283.430 2190.860 283.750 2190.920 ;
        RECT 2901.290 2190.860 2901.610 2190.920 ;
        RECT 283.430 2190.720 2901.610 2190.860 ;
        RECT 283.430 2190.660 283.750 2190.720 ;
        RECT 2901.290 2190.660 2901.610 2190.720 ;
      LAYER via ;
        RECT 283.460 2190.660 283.720 2190.920 ;
        RECT 2901.320 2190.660 2901.580 2190.920 ;
      LAYER met2 ;
        RECT 2901.310 2727.635 2901.590 2728.005 ;
        RECT 2901.380 2190.950 2901.520 2727.635 ;
        RECT 283.460 2190.630 283.720 2190.950 ;
        RECT 2901.320 2190.630 2901.580 2190.950 ;
        RECT 283.520 2179.810 283.660 2190.630 ;
        RECT 283.060 2179.670 283.660 2179.810 ;
        RECT 283.060 1963.570 283.200 2179.670 ;
        RECT 282.600 1963.430 283.200 1963.570 ;
        RECT 282.600 1959.490 282.740 1963.430 ;
        RECT 282.600 1959.350 283.200 1959.490 ;
        RECT 283.060 1953.370 283.200 1959.350 ;
        RECT 282.600 1953.230 283.200 1953.370 ;
        RECT 282.600 1945.210 282.740 1953.230 ;
        RECT 282.600 1945.070 283.200 1945.210 ;
        RECT 283.060 1939.205 283.200 1945.070 ;
        RECT 282.990 1938.835 283.270 1939.205 ;
      LAYER via2 ;
        RECT 2901.310 2727.680 2901.590 2727.960 ;
        RECT 282.990 1938.880 283.270 1939.160 ;
      LAYER met3 ;
        RECT 2901.285 2727.970 2901.615 2727.985 ;
        RECT 2917.600 2727.970 2924.800 2728.420 ;
        RECT 2901.285 2727.670 2924.800 2727.970 ;
        RECT 2901.285 2727.655 2901.615 2727.670 ;
        RECT 2917.600 2727.220 2924.800 2727.670 ;
        RECT 282.965 1939.170 283.295 1939.185 ;
        RECT 283.630 1939.170 284.010 1939.180 ;
        RECT 282.965 1938.870 284.010 1939.170 ;
        RECT 282.965 1938.855 283.295 1938.870 ;
        RECT 283.630 1938.860 284.010 1938.870 ;
        RECT 283.630 1373.410 284.010 1373.420 ;
        RECT 283.630 1373.280 300.380 1373.410 ;
        RECT 283.630 1373.110 304.000 1373.280 ;
        RECT 283.630 1373.100 284.010 1373.110 ;
        RECT 300.000 1372.680 304.000 1373.110 ;
      LAYER via3 ;
        RECT 283.660 1938.860 283.980 1939.180 ;
        RECT 283.660 1373.100 283.980 1373.420 ;
      LAYER met4 ;
        RECT 283.655 1938.855 283.985 1939.185 ;
        RECT 283.670 1373.425 283.970 1938.855 ;
        RECT 283.655 1373.095 283.985 1373.425 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 298.610 2960.280 298.930 2960.340 ;
        RECT 2900.830 2960.280 2901.150 2960.340 ;
        RECT 298.610 2960.140 2901.150 2960.280 ;
        RECT 298.610 2960.080 298.930 2960.140 ;
        RECT 2900.830 2960.080 2901.150 2960.140 ;
      LAYER via ;
        RECT 298.640 2960.080 298.900 2960.340 ;
        RECT 2900.860 2960.080 2901.120 2960.340 ;
      LAYER met2 ;
        RECT 2900.850 2962.235 2901.130 2962.605 ;
        RECT 2900.920 2960.370 2901.060 2962.235 ;
        RECT 298.640 2960.050 298.900 2960.370 ;
        RECT 2900.860 2960.050 2901.120 2960.370 ;
        RECT 298.700 1405.405 298.840 2960.050 ;
        RECT 298.630 1405.035 298.910 1405.405 ;
      LAYER via2 ;
        RECT 2900.850 2962.280 2901.130 2962.560 ;
        RECT 298.630 1405.080 298.910 1405.360 ;
      LAYER met3 ;
        RECT 2900.825 2962.570 2901.155 2962.585 ;
        RECT 2917.600 2962.570 2924.800 2963.020 ;
        RECT 2900.825 2962.270 2924.800 2962.570 ;
        RECT 2900.825 2962.255 2901.155 2962.270 ;
        RECT 2917.600 2961.820 2924.800 2962.270 ;
        RECT 298.605 1405.370 298.935 1405.385 ;
        RECT 298.605 1405.240 300.380 1405.370 ;
        RECT 298.605 1405.070 304.000 1405.240 ;
        RECT 298.605 1405.055 298.935 1405.070 ;
        RECT 300.000 1404.640 304.000 1405.070 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 298.150 3194.880 298.470 3194.940 ;
        RECT 2900.830 3194.880 2901.150 3194.940 ;
        RECT 298.150 3194.740 2901.150 3194.880 ;
        RECT 298.150 3194.680 298.470 3194.740 ;
        RECT 2900.830 3194.680 2901.150 3194.740 ;
      LAYER via ;
        RECT 298.180 3194.680 298.440 3194.940 ;
        RECT 2900.860 3194.680 2901.120 3194.940 ;
      LAYER met2 ;
        RECT 2900.850 3196.835 2901.130 3197.205 ;
        RECT 2900.920 3194.970 2901.060 3196.835 ;
        RECT 298.180 3194.650 298.440 3194.970 ;
        RECT 2900.860 3194.650 2901.120 3194.970 ;
        RECT 298.240 1436.685 298.380 3194.650 ;
        RECT 298.170 1436.315 298.450 1436.685 ;
      LAYER via2 ;
        RECT 2900.850 3196.880 2901.130 3197.160 ;
        RECT 298.170 1436.360 298.450 1436.640 ;
      LAYER met3 ;
        RECT 2900.825 3197.170 2901.155 3197.185 ;
        RECT 2917.600 3197.170 2924.800 3197.620 ;
        RECT 2900.825 3196.870 2924.800 3197.170 ;
        RECT 2900.825 3196.855 2901.155 3196.870 ;
        RECT 2917.600 3196.420 2924.800 3196.870 ;
        RECT 298.145 1436.650 298.475 1436.665 ;
        RECT 298.145 1436.520 300.380 1436.650 ;
        RECT 298.145 1436.350 304.000 1436.520 ;
        RECT 298.145 1436.335 298.475 1436.350 ;
        RECT 300.000 1435.920 304.000 1436.350 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1497.460 3429.680 1506.340 3429.820 ;
        RECT 296.770 3429.480 297.090 3429.540 ;
        RECT 1497.460 3429.480 1497.600 3429.680 ;
        RECT 296.770 3429.340 1497.600 3429.480 ;
        RECT 1506.200 3429.480 1506.340 3429.680 ;
        RECT 2762.920 3429.680 2798.940 3429.820 ;
        RECT 2762.920 3429.480 2763.060 3429.680 ;
        RECT 1506.200 3429.340 2763.060 3429.480 ;
        RECT 2798.800 3429.480 2798.940 3429.680 ;
        RECT 2900.830 3429.480 2901.150 3429.540 ;
        RECT 2798.800 3429.340 2901.150 3429.480 ;
        RECT 296.770 3429.280 297.090 3429.340 ;
        RECT 2900.830 3429.280 2901.150 3429.340 ;
      LAYER via ;
        RECT 296.800 3429.280 297.060 3429.540 ;
        RECT 2900.860 3429.280 2901.120 3429.540 ;
      LAYER met2 ;
        RECT 2900.850 3431.435 2901.130 3431.805 ;
        RECT 2900.920 3429.570 2901.060 3431.435 ;
        RECT 296.800 3429.250 297.060 3429.570 ;
        RECT 2900.860 3429.250 2901.120 3429.570 ;
        RECT 296.860 1468.645 297.000 3429.250 ;
        RECT 296.790 1468.275 297.070 1468.645 ;
      LAYER via2 ;
        RECT 2900.850 3431.480 2901.130 3431.760 ;
        RECT 296.790 1468.320 297.070 1468.600 ;
      LAYER met3 ;
        RECT 2900.825 3431.770 2901.155 3431.785 ;
        RECT 2917.600 3431.770 2924.800 3432.220 ;
        RECT 2900.825 3431.470 2924.800 3431.770 ;
        RECT 2900.825 3431.455 2901.155 3431.470 ;
        RECT 2917.600 3431.020 2924.800 3431.470 ;
        RECT 296.765 1468.610 297.095 1468.625 ;
        RECT 296.765 1468.480 300.380 1468.610 ;
        RECT 296.765 1468.310 304.000 1468.480 ;
        RECT 296.765 1468.295 297.095 1468.310 ;
        RECT 300.000 1467.880 304.000 1468.310 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
        RECT 2717.380 3501.845 2717.520 3517.600 ;
        RECT 2717.310 3501.475 2717.590 3501.845 ;
      LAYER via2 ;
        RECT 2717.310 3501.520 2717.590 3501.800 ;
      LAYER met3 ;
        RECT 289.150 3501.810 289.530 3501.820 ;
        RECT 2717.285 3501.810 2717.615 3501.825 ;
        RECT 289.150 3501.510 2717.615 3501.810 ;
        RECT 289.150 3501.500 289.530 3501.510 ;
        RECT 2717.285 3501.495 2717.615 3501.510 ;
        RECT 289.150 1499.890 289.530 1499.900 ;
        RECT 289.150 1499.760 300.380 1499.890 ;
        RECT 289.150 1499.590 304.000 1499.760 ;
        RECT 289.150 1499.580 289.530 1499.590 ;
        RECT 300.000 1499.160 304.000 1499.590 ;
      LAYER via3 ;
        RECT 289.180 3501.500 289.500 3501.820 ;
        RECT 289.180 1499.580 289.500 1499.900 ;
      LAYER met4 ;
        RECT 289.175 3501.495 289.505 3501.825 ;
        RECT 289.190 1499.905 289.490 3501.495 ;
        RECT 289.175 1499.575 289.505 1499.905 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
        RECT 2392.620 3503.885 2392.760 3517.600 ;
        RECT 2392.550 3503.515 2392.830 3503.885 ;
      LAYER via2 ;
        RECT 2392.550 3503.560 2392.830 3503.840 ;
      LAYER met3 ;
        RECT 287.310 3503.850 287.690 3503.860 ;
        RECT 2392.525 3503.850 2392.855 3503.865 ;
        RECT 287.310 3503.550 2392.855 3503.850 ;
        RECT 287.310 3503.540 287.690 3503.550 ;
        RECT 2392.525 3503.535 2392.855 3503.550 ;
        RECT 287.310 1531.850 287.690 1531.860 ;
        RECT 287.310 1531.720 300.380 1531.850 ;
        RECT 287.310 1531.550 304.000 1531.720 ;
        RECT 287.310 1531.540 287.690 1531.550 ;
        RECT 300.000 1531.120 304.000 1531.550 ;
      LAYER via3 ;
        RECT 287.340 3503.540 287.660 3503.860 ;
        RECT 287.340 1531.540 287.660 1531.860 ;
      LAYER met4 ;
        RECT 287.335 3503.535 287.665 3503.865 ;
        RECT 287.350 1531.865 287.650 3503.535 ;
        RECT 287.335 1531.535 287.665 1531.865 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 295.390 3501.900 295.710 3501.960 ;
        RECT 2068.230 3501.900 2068.550 3501.960 ;
        RECT 295.390 3501.760 2068.550 3501.900 ;
        RECT 295.390 3501.700 295.710 3501.760 ;
        RECT 2068.230 3501.700 2068.550 3501.760 ;
      LAYER via ;
        RECT 295.420 3501.700 295.680 3501.960 ;
        RECT 2068.260 3501.700 2068.520 3501.960 ;
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
        RECT 2068.320 3501.990 2068.460 3517.600 ;
        RECT 295.420 3501.670 295.680 3501.990 ;
        RECT 2068.260 3501.670 2068.520 3501.990 ;
        RECT 295.480 1563.165 295.620 3501.670 ;
        RECT 295.410 1562.795 295.690 1563.165 ;
      LAYER via2 ;
        RECT 295.410 1562.840 295.690 1563.120 ;
      LAYER met3 ;
        RECT 295.385 1563.130 295.715 1563.145 ;
        RECT 295.385 1563.000 300.380 1563.130 ;
        RECT 295.385 1562.830 304.000 1563.000 ;
        RECT 295.385 1562.815 295.715 1562.830 ;
        RECT 300.000 1562.400 304.000 1562.830 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 289.410 3502.580 289.730 3502.640 ;
        RECT 1743.930 3502.580 1744.250 3502.640 ;
        RECT 289.410 3502.440 1744.250 3502.580 ;
        RECT 289.410 3502.380 289.730 3502.440 ;
        RECT 1743.930 3502.380 1744.250 3502.440 ;
      LAYER via ;
        RECT 289.440 3502.380 289.700 3502.640 ;
        RECT 1743.960 3502.380 1744.220 3502.640 ;
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
        RECT 1744.020 3502.670 1744.160 3517.600 ;
        RECT 289.440 3502.350 289.700 3502.670 ;
        RECT 1743.960 3502.350 1744.220 3502.670 ;
        RECT 289.500 1595.125 289.640 3502.350 ;
        RECT 289.430 1594.755 289.710 1595.125 ;
      LAYER via2 ;
        RECT 289.430 1594.800 289.710 1595.080 ;
      LAYER met3 ;
        RECT 289.405 1595.090 289.735 1595.105 ;
        RECT 289.405 1594.960 300.380 1595.090 ;
        RECT 289.405 1594.790 304.000 1594.960 ;
        RECT 289.405 1594.775 289.735 1594.790 ;
        RECT 300.000 1594.360 304.000 1594.790 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 297.230 3503.600 297.550 3503.660 ;
        RECT 1419.170 3503.600 1419.490 3503.660 ;
        RECT 297.230 3503.460 1419.490 3503.600 ;
        RECT 297.230 3503.400 297.550 3503.460 ;
        RECT 1419.170 3503.400 1419.490 3503.460 ;
      LAYER via ;
        RECT 297.260 3503.400 297.520 3503.660 ;
        RECT 1419.200 3503.400 1419.460 3503.660 ;
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
        RECT 1419.260 3503.690 1419.400 3517.600 ;
        RECT 297.260 3503.370 297.520 3503.690 ;
        RECT 1419.200 3503.370 1419.460 3503.690 ;
        RECT 297.320 1626.405 297.460 3503.370 ;
        RECT 297.250 1626.035 297.530 1626.405 ;
      LAYER via2 ;
        RECT 297.250 1626.080 297.530 1626.360 ;
      LAYER met3 ;
        RECT 297.225 1626.370 297.555 1626.385 ;
        RECT 297.225 1626.240 300.380 1626.370 ;
        RECT 297.225 1626.070 304.000 1626.240 ;
        RECT 297.225 1626.055 297.555 1626.070 ;
        RECT 300.000 1625.640 304.000 1626.070 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 448.110 381.380 448.430 381.440 ;
        RECT 482.610 381.380 482.930 381.440 ;
        RECT 448.110 381.240 482.930 381.380 ;
        RECT 448.110 381.180 448.430 381.240 ;
        RECT 482.610 381.180 482.930 381.240 ;
        RECT 737.910 380.700 738.230 380.760 ;
        RECT 772.410 380.700 772.730 380.760 ;
        RECT 737.910 380.560 772.730 380.700 ;
        RECT 737.910 380.500 738.230 380.560 ;
        RECT 772.410 380.500 772.730 380.560 ;
        RECT 580.130 380.020 580.450 380.080 ;
        RECT 593.930 380.020 594.250 380.080 ;
        RECT 580.130 379.880 594.250 380.020 ;
        RECT 580.130 379.820 580.450 379.880 ;
        RECT 593.930 379.820 594.250 379.880 ;
      LAYER via ;
        RECT 448.140 381.180 448.400 381.440 ;
        RECT 482.640 381.180 482.900 381.440 ;
        RECT 737.940 380.500 738.200 380.760 ;
        RECT 772.440 380.500 772.700 380.760 ;
        RECT 580.160 379.820 580.420 380.080 ;
        RECT 593.960 379.820 594.220 380.080 ;
      LAYER met2 ;
        RECT 675.830 382.315 676.110 382.685 ;
        RECT 448.140 381.325 448.400 381.470 ;
        RECT 482.640 381.325 482.900 381.470 ;
        RECT 448.130 380.955 448.410 381.325 ;
        RECT 482.630 380.955 482.910 381.325 ;
        RECT 593.950 380.955 594.230 381.325 ;
        RECT 594.020 380.110 594.160 380.955 ;
        RECT 675.900 380.645 676.040 382.315 ;
        RECT 700.210 381.635 700.490 382.005 ;
        RECT 675.830 380.275 676.110 380.645 ;
        RECT 580.160 379.965 580.420 380.110 ;
        RECT 580.150 379.595 580.430 379.965 ;
        RECT 593.960 379.790 594.220 380.110 ;
        RECT 700.280 379.965 700.420 381.635 ;
        RECT 772.430 380.955 772.710 381.325 ;
        RECT 772.500 380.790 772.640 380.955 ;
        RECT 737.940 380.645 738.200 380.790 ;
        RECT 737.930 380.275 738.210 380.645 ;
        RECT 772.440 380.470 772.700 380.790 ;
        RECT 700.210 379.595 700.490 379.965 ;
      LAYER via2 ;
        RECT 675.830 382.360 676.110 382.640 ;
        RECT 448.130 381.000 448.410 381.280 ;
        RECT 482.630 381.000 482.910 381.280 ;
        RECT 593.950 381.000 594.230 381.280 ;
        RECT 700.210 381.680 700.490 381.960 ;
        RECT 675.830 380.320 676.110 380.600 ;
        RECT 580.150 379.640 580.430 379.920 ;
        RECT 772.430 381.000 772.710 381.280 ;
        RECT 737.930 380.320 738.210 380.600 ;
        RECT 700.210 379.640 700.490 379.920 ;
      LAYER met3 ;
        RECT 286.390 1057.890 286.770 1057.900 ;
        RECT 286.390 1057.760 300.380 1057.890 ;
        RECT 286.390 1057.590 304.000 1057.760 ;
        RECT 286.390 1057.580 286.770 1057.590 ;
        RECT 300.000 1057.160 304.000 1057.590 ;
        RECT 627.710 382.650 628.090 382.660 ;
        RECT 675.805 382.650 676.135 382.665 ;
        RECT 627.710 382.350 676.135 382.650 ;
        RECT 627.710 382.340 628.090 382.350 ;
        RECT 675.805 382.335 676.135 382.350 ;
        RECT 578.950 381.970 579.330 381.980 ;
        RECT 700.185 381.970 700.515 381.985 ;
        RECT 544.030 381.670 579.330 381.970 ;
        RECT 286.390 381.290 286.770 381.300 ;
        RECT 448.105 381.290 448.435 381.305 ;
        RECT 286.390 380.990 324.450 381.290 ;
        RECT 286.390 380.980 286.770 380.990 ;
        RECT 324.150 380.610 324.450 380.990 ;
        RECT 372.910 380.990 448.435 381.290 ;
        RECT 324.150 380.310 372.290 380.610 ;
        RECT 371.990 379.930 372.290 380.310 ;
        RECT 372.910 379.930 373.210 380.990 ;
        RECT 448.105 380.975 448.435 380.990 ;
        RECT 482.605 381.290 482.935 381.305 ;
        RECT 482.605 380.990 496.490 381.290 ;
        RECT 482.605 380.975 482.935 380.990 ;
        RECT 371.990 379.630 373.210 379.930 ;
        RECT 496.190 379.930 496.490 380.990 ;
        RECT 544.030 380.610 544.330 381.670 ;
        RECT 578.950 381.660 579.330 381.670 ;
        RECT 676.510 381.670 700.515 381.970 ;
        RECT 593.925 381.290 594.255 381.305 ;
        RECT 627.710 381.290 628.090 381.300 ;
        RECT 593.925 380.990 628.090 381.290 ;
        RECT 593.925 380.975 594.255 380.990 ;
        RECT 627.710 380.980 628.090 380.990 ;
        RECT 497.110 380.310 544.330 380.610 ;
        RECT 675.805 380.610 676.135 380.625 ;
        RECT 676.510 380.610 676.810 381.670 ;
        RECT 700.185 381.655 700.515 381.670 ;
        RECT 772.405 381.290 772.735 381.305 ;
        RECT 2917.600 381.290 2924.800 381.740 ;
        RECT 772.405 380.990 807.450 381.290 ;
        RECT 772.405 380.975 772.735 380.990 ;
        RECT 737.905 380.610 738.235 380.625 ;
        RECT 675.805 380.310 676.810 380.610 ;
        RECT 724.350 380.310 738.235 380.610 ;
        RECT 807.150 380.610 807.450 380.990 ;
        RECT 855.910 380.990 904.050 381.290 ;
        RECT 807.150 380.310 855.290 380.610 ;
        RECT 497.110 379.930 497.410 380.310 ;
        RECT 675.805 380.295 676.135 380.310 ;
        RECT 496.190 379.630 497.410 379.930 ;
        RECT 578.950 379.930 579.330 379.940 ;
        RECT 580.125 379.930 580.455 379.945 ;
        RECT 578.950 379.630 580.455 379.930 ;
        RECT 578.950 379.620 579.330 379.630 ;
        RECT 580.125 379.615 580.455 379.630 ;
        RECT 700.185 379.930 700.515 379.945 ;
        RECT 724.350 379.930 724.650 380.310 ;
        RECT 737.905 380.295 738.235 380.310 ;
        RECT 700.185 379.630 724.650 379.930 ;
        RECT 854.990 379.930 855.290 380.310 ;
        RECT 855.910 379.930 856.210 380.990 ;
        RECT 903.750 380.610 904.050 380.990 ;
        RECT 952.510 380.990 1000.650 381.290 ;
        RECT 903.750 380.310 951.890 380.610 ;
        RECT 854.990 379.630 856.210 379.930 ;
        RECT 951.590 379.930 951.890 380.310 ;
        RECT 952.510 379.930 952.810 380.990 ;
        RECT 1000.350 380.610 1000.650 380.990 ;
        RECT 1049.110 380.990 1097.250 381.290 ;
        RECT 1000.350 380.310 1048.490 380.610 ;
        RECT 951.590 379.630 952.810 379.930 ;
        RECT 1048.190 379.930 1048.490 380.310 ;
        RECT 1049.110 379.930 1049.410 380.990 ;
        RECT 1096.950 380.610 1097.250 380.990 ;
        RECT 1145.710 380.990 1193.850 381.290 ;
        RECT 1096.950 380.310 1145.090 380.610 ;
        RECT 1048.190 379.630 1049.410 379.930 ;
        RECT 1144.790 379.930 1145.090 380.310 ;
        RECT 1145.710 379.930 1146.010 380.990 ;
        RECT 1193.550 380.610 1193.850 380.990 ;
        RECT 1242.310 380.990 1290.450 381.290 ;
        RECT 1193.550 380.310 1241.690 380.610 ;
        RECT 1144.790 379.630 1146.010 379.930 ;
        RECT 1241.390 379.930 1241.690 380.310 ;
        RECT 1242.310 379.930 1242.610 380.990 ;
        RECT 1290.150 380.610 1290.450 380.990 ;
        RECT 1338.910 380.990 1387.050 381.290 ;
        RECT 1290.150 380.310 1338.290 380.610 ;
        RECT 1241.390 379.630 1242.610 379.930 ;
        RECT 1337.990 379.930 1338.290 380.310 ;
        RECT 1338.910 379.930 1339.210 380.990 ;
        RECT 1386.750 380.610 1387.050 380.990 ;
        RECT 1435.510 380.990 1483.650 381.290 ;
        RECT 1386.750 380.310 1434.890 380.610 ;
        RECT 1337.990 379.630 1339.210 379.930 ;
        RECT 1434.590 379.930 1434.890 380.310 ;
        RECT 1435.510 379.930 1435.810 380.990 ;
        RECT 1483.350 380.610 1483.650 380.990 ;
        RECT 1532.110 380.990 1580.250 381.290 ;
        RECT 1483.350 380.310 1531.490 380.610 ;
        RECT 1434.590 379.630 1435.810 379.930 ;
        RECT 1531.190 379.930 1531.490 380.310 ;
        RECT 1532.110 379.930 1532.410 380.990 ;
        RECT 1579.950 380.610 1580.250 380.990 ;
        RECT 1628.710 380.990 1676.850 381.290 ;
        RECT 1579.950 380.310 1628.090 380.610 ;
        RECT 1531.190 379.630 1532.410 379.930 ;
        RECT 1627.790 379.930 1628.090 380.310 ;
        RECT 1628.710 379.930 1629.010 380.990 ;
        RECT 1676.550 380.610 1676.850 380.990 ;
        RECT 1725.310 380.990 1773.450 381.290 ;
        RECT 1676.550 380.310 1724.690 380.610 ;
        RECT 1627.790 379.630 1629.010 379.930 ;
        RECT 1724.390 379.930 1724.690 380.310 ;
        RECT 1725.310 379.930 1725.610 380.990 ;
        RECT 1773.150 380.610 1773.450 380.990 ;
        RECT 1821.910 380.990 1870.050 381.290 ;
        RECT 1773.150 380.310 1821.290 380.610 ;
        RECT 1724.390 379.630 1725.610 379.930 ;
        RECT 1820.990 379.930 1821.290 380.310 ;
        RECT 1821.910 379.930 1822.210 380.990 ;
        RECT 1869.750 380.610 1870.050 380.990 ;
        RECT 1918.510 380.990 1966.650 381.290 ;
        RECT 1869.750 380.310 1917.890 380.610 ;
        RECT 1820.990 379.630 1822.210 379.930 ;
        RECT 1917.590 379.930 1917.890 380.310 ;
        RECT 1918.510 379.930 1918.810 380.990 ;
        RECT 1966.350 380.610 1966.650 380.990 ;
        RECT 2015.110 380.990 2063.250 381.290 ;
        RECT 1966.350 380.310 2014.490 380.610 ;
        RECT 1917.590 379.630 1918.810 379.930 ;
        RECT 2014.190 379.930 2014.490 380.310 ;
        RECT 2015.110 379.930 2015.410 380.990 ;
        RECT 2062.950 380.610 2063.250 380.990 ;
        RECT 2111.710 380.990 2159.850 381.290 ;
        RECT 2062.950 380.310 2111.090 380.610 ;
        RECT 2014.190 379.630 2015.410 379.930 ;
        RECT 2110.790 379.930 2111.090 380.310 ;
        RECT 2111.710 379.930 2112.010 380.990 ;
        RECT 2159.550 380.610 2159.850 380.990 ;
        RECT 2208.310 380.990 2256.450 381.290 ;
        RECT 2159.550 380.310 2207.690 380.610 ;
        RECT 2110.790 379.630 2112.010 379.930 ;
        RECT 2207.390 379.930 2207.690 380.310 ;
        RECT 2208.310 379.930 2208.610 380.990 ;
        RECT 2256.150 380.610 2256.450 380.990 ;
        RECT 2304.910 380.990 2353.050 381.290 ;
        RECT 2256.150 380.310 2304.290 380.610 ;
        RECT 2207.390 379.630 2208.610 379.930 ;
        RECT 2303.990 379.930 2304.290 380.310 ;
        RECT 2304.910 379.930 2305.210 380.990 ;
        RECT 2352.750 380.610 2353.050 380.990 ;
        RECT 2401.510 380.990 2449.650 381.290 ;
        RECT 2352.750 380.310 2400.890 380.610 ;
        RECT 2303.990 379.630 2305.210 379.930 ;
        RECT 2400.590 379.930 2400.890 380.310 ;
        RECT 2401.510 379.930 2401.810 380.990 ;
        RECT 2449.350 380.610 2449.650 380.990 ;
        RECT 2498.110 380.990 2546.250 381.290 ;
        RECT 2449.350 380.310 2497.490 380.610 ;
        RECT 2400.590 379.630 2401.810 379.930 ;
        RECT 2497.190 379.930 2497.490 380.310 ;
        RECT 2498.110 379.930 2498.410 380.990 ;
        RECT 2545.950 380.610 2546.250 380.990 ;
        RECT 2594.710 380.990 2642.850 381.290 ;
        RECT 2545.950 380.310 2594.090 380.610 ;
        RECT 2497.190 379.630 2498.410 379.930 ;
        RECT 2593.790 379.930 2594.090 380.310 ;
        RECT 2594.710 379.930 2595.010 380.990 ;
        RECT 2642.550 380.610 2642.850 380.990 ;
        RECT 2691.310 380.990 2739.450 381.290 ;
        RECT 2642.550 380.310 2690.690 380.610 ;
        RECT 2593.790 379.630 2595.010 379.930 ;
        RECT 2690.390 379.930 2690.690 380.310 ;
        RECT 2691.310 379.930 2691.610 380.990 ;
        RECT 2739.150 380.610 2739.450 380.990 ;
        RECT 2787.910 380.990 2836.050 381.290 ;
        RECT 2739.150 380.310 2787.290 380.610 ;
        RECT 2690.390 379.630 2691.610 379.930 ;
        RECT 2786.990 379.930 2787.290 380.310 ;
        RECT 2787.910 379.930 2788.210 380.990 ;
        RECT 2835.750 380.610 2836.050 380.990 ;
        RECT 2916.710 380.990 2924.800 381.290 ;
        RECT 2916.710 380.610 2917.010 380.990 ;
        RECT 2835.750 380.310 2883.890 380.610 ;
        RECT 2786.990 379.630 2788.210 379.930 ;
        RECT 2883.590 379.930 2883.890 380.310 ;
        RECT 2884.510 380.310 2917.010 380.610 ;
        RECT 2917.600 380.540 2924.800 380.990 ;
        RECT 2884.510 379.930 2884.810 380.310 ;
        RECT 2883.590 379.630 2884.810 379.930 ;
        RECT 700.185 379.615 700.515 379.630 ;
      LAYER via3 ;
        RECT 286.420 1057.580 286.740 1057.900 ;
        RECT 627.740 382.340 628.060 382.660 ;
        RECT 286.420 380.980 286.740 381.300 ;
        RECT 578.980 381.660 579.300 381.980 ;
        RECT 627.740 380.980 628.060 381.300 ;
        RECT 578.980 379.620 579.300 379.940 ;
      LAYER met4 ;
        RECT 286.415 1057.575 286.745 1057.905 ;
        RECT 286.430 381.305 286.730 1057.575 ;
        RECT 627.735 382.335 628.065 382.665 ;
        RECT 578.975 381.655 579.305 381.985 ;
        RECT 286.415 380.975 286.745 381.305 ;
        RECT 578.990 379.945 579.290 381.655 ;
        RECT 627.750 381.305 628.050 382.335 ;
        RECT 627.735 380.975 628.065 381.305 ;
        RECT 578.975 379.615 579.305 379.945 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 288.950 3504.280 289.270 3504.340 ;
        RECT 1094.870 3504.280 1095.190 3504.340 ;
        RECT 288.950 3504.140 1095.190 3504.280 ;
        RECT 288.950 3504.080 289.270 3504.140 ;
        RECT 1094.870 3504.080 1095.190 3504.140 ;
      LAYER via ;
        RECT 288.980 3504.080 289.240 3504.340 ;
        RECT 1094.900 3504.080 1095.160 3504.340 ;
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
        RECT 1094.960 3504.370 1095.100 3517.600 ;
        RECT 288.980 3504.050 289.240 3504.370 ;
        RECT 1094.900 3504.050 1095.160 3504.370 ;
        RECT 289.040 1657.685 289.180 3504.050 ;
        RECT 288.970 1657.315 289.250 1657.685 ;
      LAYER via2 ;
        RECT 288.970 1657.360 289.250 1657.640 ;
      LAYER met3 ;
        RECT 288.945 1657.650 289.275 1657.665 ;
        RECT 288.945 1657.520 300.380 1657.650 ;
        RECT 288.945 1657.350 304.000 1657.520 ;
        RECT 288.945 1657.335 289.275 1657.350 ;
        RECT 300.000 1656.920 304.000 1657.350 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 293.090 3500.880 293.410 3500.940 ;
        RECT 770.570 3500.880 770.890 3500.940 ;
        RECT 293.090 3500.740 770.890 3500.880 ;
        RECT 293.090 3500.680 293.410 3500.740 ;
        RECT 770.570 3500.680 770.890 3500.740 ;
      LAYER via ;
        RECT 293.120 3500.680 293.380 3500.940 ;
        RECT 770.600 3500.680 770.860 3500.940 ;
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
        RECT 770.660 3500.970 770.800 3517.600 ;
        RECT 293.120 3500.650 293.380 3500.970 ;
        RECT 770.600 3500.650 770.860 3500.970 ;
        RECT 293.180 1689.645 293.320 3500.650 ;
        RECT 293.110 1689.275 293.390 1689.645 ;
      LAYER via2 ;
        RECT 293.110 1689.320 293.390 1689.600 ;
      LAYER met3 ;
        RECT 293.085 1689.610 293.415 1689.625 ;
        RECT 293.085 1689.480 300.380 1689.610 ;
        RECT 293.085 1689.310 304.000 1689.480 ;
        RECT 293.085 1689.295 293.415 1689.310 ;
        RECT 300.000 1688.880 304.000 1689.310 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 292.170 3501.220 292.490 3501.280 ;
        RECT 445.810 3501.220 446.130 3501.280 ;
        RECT 292.170 3501.080 446.130 3501.220 ;
        RECT 292.170 3501.020 292.490 3501.080 ;
        RECT 445.810 3501.020 446.130 3501.080 ;
      LAYER via ;
        RECT 292.200 3501.020 292.460 3501.280 ;
        RECT 445.840 3501.020 446.100 3501.280 ;
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
        RECT 445.900 3501.310 446.040 3517.600 ;
        RECT 292.200 3500.990 292.460 3501.310 ;
        RECT 445.840 3500.990 446.100 3501.310 ;
        RECT 292.260 1720.925 292.400 3500.990 ;
        RECT 292.190 1720.555 292.470 1720.925 ;
      LAYER via2 ;
        RECT 292.190 1720.600 292.470 1720.880 ;
      LAYER met3 ;
        RECT 292.165 1720.890 292.495 1720.905 ;
        RECT 292.165 1720.760 300.380 1720.890 ;
        RECT 292.165 1720.590 304.000 1720.760 ;
        RECT 292.165 1720.575 292.495 1720.590 ;
        RECT 300.000 1720.160 304.000 1720.590 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 121.510 3498.500 121.830 3498.560 ;
        RECT 123.810 3498.500 124.130 3498.560 ;
        RECT 121.510 3498.360 124.130 3498.500 ;
        RECT 121.510 3498.300 121.830 3498.360 ;
        RECT 123.810 3498.300 124.130 3498.360 ;
        RECT 123.810 1759.400 124.130 1759.460 ;
        RECT 282.970 1759.400 283.290 1759.460 ;
        RECT 123.810 1759.260 283.290 1759.400 ;
        RECT 123.810 1759.200 124.130 1759.260 ;
        RECT 282.970 1759.200 283.290 1759.260 ;
      LAYER via ;
        RECT 121.540 3498.300 121.800 3498.560 ;
        RECT 123.840 3498.300 124.100 3498.560 ;
        RECT 123.840 1759.200 124.100 1759.460 ;
        RECT 283.000 1759.200 283.260 1759.460 ;
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
        RECT 121.600 3498.590 121.740 3517.600 ;
        RECT 121.540 3498.270 121.800 3498.590 ;
        RECT 123.840 3498.270 124.100 3498.590 ;
        RECT 123.900 1759.490 124.040 3498.270 ;
        RECT 123.840 1759.170 124.100 1759.490 ;
        RECT 283.000 1759.170 283.260 1759.490 ;
        RECT 283.060 1752.885 283.200 1759.170 ;
        RECT 282.990 1752.515 283.270 1752.885 ;
      LAYER via2 ;
        RECT 282.990 1752.560 283.270 1752.840 ;
      LAYER met3 ;
        RECT 282.965 1752.850 283.295 1752.865 ;
        RECT 282.965 1752.720 300.380 1752.850 ;
        RECT 282.965 1752.550 304.000 1752.720 ;
        RECT 282.965 1752.535 283.295 1752.550 ;
        RECT 300.000 1752.120 304.000 1752.550 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 3339.720 17.410 3339.780 ;
        RECT 106.790 3339.720 107.110 3339.780 ;
        RECT 17.090 3339.580 107.110 3339.720 ;
        RECT 17.090 3339.520 17.410 3339.580 ;
        RECT 106.790 3339.520 107.110 3339.580 ;
        RECT 106.790 1786.940 107.110 1787.000 ;
        RECT 282.970 1786.940 283.290 1787.000 ;
        RECT 106.790 1786.800 283.290 1786.940 ;
        RECT 106.790 1786.740 107.110 1786.800 ;
        RECT 282.970 1786.740 283.290 1786.800 ;
      LAYER via ;
        RECT 17.120 3339.520 17.380 3339.780 ;
        RECT 106.820 3339.520 107.080 3339.780 ;
        RECT 106.820 1786.740 107.080 1787.000 ;
        RECT 283.000 1786.740 283.260 1787.000 ;
      LAYER met2 ;
        RECT 17.110 3339.635 17.390 3340.005 ;
        RECT 17.120 3339.490 17.380 3339.635 ;
        RECT 106.820 3339.490 107.080 3339.810 ;
        RECT 106.880 1787.030 107.020 3339.490 ;
        RECT 106.820 1786.710 107.080 1787.030 ;
        RECT 283.000 1786.710 283.260 1787.030 ;
        RECT 283.060 1784.165 283.200 1786.710 ;
        RECT 282.990 1783.795 283.270 1784.165 ;
      LAYER via2 ;
        RECT 17.110 3339.680 17.390 3339.960 ;
        RECT 282.990 1783.840 283.270 1784.120 ;
      LAYER met3 ;
        RECT -4.800 3339.970 2.400 3340.420 ;
        RECT 17.085 3339.970 17.415 3339.985 ;
        RECT -4.800 3339.670 17.415 3339.970 ;
        RECT -4.800 3339.220 2.400 3339.670 ;
        RECT 17.085 3339.655 17.415 3339.670 ;
        RECT 282.965 1784.130 283.295 1784.145 ;
        RECT 282.965 1784.000 300.380 1784.130 ;
        RECT 282.965 1783.830 304.000 1784.000 ;
        RECT 282.965 1783.815 283.295 1783.830 ;
        RECT 300.000 1783.400 304.000 1783.830 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 3050.040 17.410 3050.100 ;
        RECT 141.290 3050.040 141.610 3050.100 ;
        RECT 17.090 3049.900 141.610 3050.040 ;
        RECT 17.090 3049.840 17.410 3049.900 ;
        RECT 141.290 3049.840 141.610 3049.900 ;
        RECT 141.290 1821.620 141.610 1821.680 ;
        RECT 282.970 1821.620 283.290 1821.680 ;
        RECT 141.290 1821.480 283.290 1821.620 ;
        RECT 141.290 1821.420 141.610 1821.480 ;
        RECT 282.970 1821.420 283.290 1821.480 ;
      LAYER via ;
        RECT 17.120 3049.840 17.380 3050.100 ;
        RECT 141.320 3049.840 141.580 3050.100 ;
        RECT 141.320 1821.420 141.580 1821.680 ;
        RECT 283.000 1821.420 283.260 1821.680 ;
      LAYER met2 ;
        RECT 17.110 3051.995 17.390 3052.365 ;
        RECT 17.180 3050.130 17.320 3051.995 ;
        RECT 17.120 3049.810 17.380 3050.130 ;
        RECT 141.320 3049.810 141.580 3050.130 ;
        RECT 141.380 1821.710 141.520 3049.810 ;
        RECT 141.320 1821.390 141.580 1821.710 ;
        RECT 283.000 1821.390 283.260 1821.710 ;
        RECT 283.060 1816.125 283.200 1821.390 ;
        RECT 282.990 1815.755 283.270 1816.125 ;
      LAYER via2 ;
        RECT 17.110 3052.040 17.390 3052.320 ;
        RECT 282.990 1815.800 283.270 1816.080 ;
      LAYER met3 ;
        RECT -4.800 3052.330 2.400 3052.780 ;
        RECT 17.085 3052.330 17.415 3052.345 ;
        RECT -4.800 3052.030 17.415 3052.330 ;
        RECT -4.800 3051.580 2.400 3052.030 ;
        RECT 17.085 3052.015 17.415 3052.030 ;
        RECT 282.965 1816.090 283.295 1816.105 ;
        RECT 282.965 1815.960 300.380 1816.090 ;
        RECT 282.965 1815.790 304.000 1815.960 ;
        RECT 282.965 1815.775 283.295 1815.790 ;
        RECT 300.000 1815.360 304.000 1815.790 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 2760.360 16.030 2760.420 ;
        RECT 161.990 2760.360 162.310 2760.420 ;
        RECT 15.710 2760.220 162.310 2760.360 ;
        RECT 15.710 2760.160 16.030 2760.220 ;
        RECT 161.990 2760.160 162.310 2760.220 ;
        RECT 161.990 1849.160 162.310 1849.220 ;
        RECT 282.970 1849.160 283.290 1849.220 ;
        RECT 161.990 1849.020 283.290 1849.160 ;
        RECT 161.990 1848.960 162.310 1849.020 ;
        RECT 282.970 1848.960 283.290 1849.020 ;
      LAYER via ;
        RECT 15.740 2760.160 16.000 2760.420 ;
        RECT 162.020 2760.160 162.280 2760.420 ;
        RECT 162.020 1848.960 162.280 1849.220 ;
        RECT 283.000 1848.960 283.260 1849.220 ;
      LAYER met2 ;
        RECT 15.730 2765.035 16.010 2765.405 ;
        RECT 15.800 2760.450 15.940 2765.035 ;
        RECT 15.740 2760.130 16.000 2760.450 ;
        RECT 162.020 2760.130 162.280 2760.450 ;
        RECT 162.080 1849.250 162.220 2760.130 ;
        RECT 162.020 1848.930 162.280 1849.250 ;
        RECT 283.000 1848.930 283.260 1849.250 ;
        RECT 283.060 1847.405 283.200 1848.930 ;
        RECT 282.990 1847.035 283.270 1847.405 ;
      LAYER via2 ;
        RECT 15.730 2765.080 16.010 2765.360 ;
        RECT 282.990 1847.080 283.270 1847.360 ;
      LAYER met3 ;
        RECT -4.800 2765.370 2.400 2765.820 ;
        RECT 15.705 2765.370 16.035 2765.385 ;
        RECT -4.800 2765.070 16.035 2765.370 ;
        RECT -4.800 2764.620 2.400 2765.070 ;
        RECT 15.705 2765.055 16.035 2765.070 ;
        RECT 282.965 1847.370 283.295 1847.385 ;
        RECT 282.965 1847.240 300.380 1847.370 ;
        RECT 282.965 1847.070 304.000 1847.240 ;
        RECT 282.965 1847.055 283.295 1847.070 ;
        RECT 300.000 1846.640 304.000 1847.070 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.930 1883.500 19.250 1883.560 ;
        RECT 282.970 1883.500 283.290 1883.560 ;
        RECT 18.930 1883.360 283.290 1883.500 ;
        RECT 18.930 1883.300 19.250 1883.360 ;
        RECT 282.970 1883.300 283.290 1883.360 ;
      LAYER via ;
        RECT 18.960 1883.300 19.220 1883.560 ;
        RECT 283.000 1883.300 283.260 1883.560 ;
      LAYER met2 ;
        RECT 18.950 2477.395 19.230 2477.765 ;
        RECT 19.020 1883.590 19.160 2477.395 ;
        RECT 18.960 1883.270 19.220 1883.590 ;
        RECT 283.000 1883.270 283.260 1883.590 ;
        RECT 283.060 1879.365 283.200 1883.270 ;
        RECT 282.990 1878.995 283.270 1879.365 ;
      LAYER via2 ;
        RECT 18.950 2477.440 19.230 2477.720 ;
        RECT 282.990 1879.040 283.270 1879.320 ;
      LAYER met3 ;
        RECT -4.800 2477.730 2.400 2478.180 ;
        RECT 18.925 2477.730 19.255 2477.745 ;
        RECT -4.800 2477.430 19.255 2477.730 ;
        RECT -4.800 2476.980 2.400 2477.430 ;
        RECT 18.925 2477.415 19.255 2477.430 ;
        RECT 282.965 1879.330 283.295 1879.345 ;
        RECT 282.965 1879.200 300.380 1879.330 ;
        RECT 282.965 1879.030 304.000 1879.200 ;
        RECT 282.965 1879.015 283.295 1879.030 ;
        RECT 300.000 1878.600 304.000 1879.030 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 1911.040 16.950 1911.100 ;
        RECT 282.970 1911.040 283.290 1911.100 ;
        RECT 16.630 1910.900 283.290 1911.040 ;
        RECT 16.630 1910.840 16.950 1910.900 ;
        RECT 282.970 1910.840 283.290 1910.900 ;
      LAYER via ;
        RECT 16.660 1910.840 16.920 1911.100 ;
        RECT 283.000 1910.840 283.260 1911.100 ;
      LAYER met2 ;
        RECT 16.650 2189.755 16.930 2190.125 ;
        RECT 16.720 1911.130 16.860 2189.755 ;
        RECT 16.660 1910.810 16.920 1911.130 ;
        RECT 283.000 1910.810 283.260 1911.130 ;
        RECT 283.060 1910.645 283.200 1910.810 ;
        RECT 282.990 1910.275 283.270 1910.645 ;
      LAYER via2 ;
        RECT 16.650 2189.800 16.930 2190.080 ;
        RECT 282.990 1910.320 283.270 1910.600 ;
      LAYER met3 ;
        RECT -4.800 2190.090 2.400 2190.540 ;
        RECT 16.625 2190.090 16.955 2190.105 ;
        RECT -4.800 2189.790 16.955 2190.090 ;
        RECT -4.800 2189.340 2.400 2189.790 ;
        RECT 16.625 2189.775 16.955 2189.790 ;
        RECT 282.965 1910.610 283.295 1910.625 ;
        RECT 282.965 1910.480 300.380 1910.610 ;
        RECT 282.965 1910.310 304.000 1910.480 ;
        RECT 282.965 1910.295 283.295 1910.310 ;
        RECT 300.000 1909.880 304.000 1910.310 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 1903.900 16.950 1903.960 ;
        RECT 282.970 1903.900 283.290 1903.960 ;
        RECT 16.630 1903.760 283.290 1903.900 ;
        RECT 16.630 1903.700 16.950 1903.760 ;
        RECT 282.970 1903.700 283.290 1903.760 ;
      LAYER via ;
        RECT 16.660 1903.700 16.920 1903.960 ;
        RECT 283.000 1903.700 283.260 1903.960 ;
      LAYER met2 ;
        RECT 282.990 1938.155 283.270 1938.525 ;
        RECT 283.060 1932.290 283.200 1938.155 ;
        RECT 282.600 1932.150 283.200 1932.290 ;
        RECT 282.600 1920.050 282.740 1932.150 ;
        RECT 282.600 1919.910 283.200 1920.050 ;
        RECT 283.060 1911.890 283.200 1919.910 ;
        RECT 282.600 1911.750 283.200 1911.890 ;
        RECT 282.600 1909.850 282.740 1911.750 ;
        RECT 282.600 1909.710 283.200 1909.850 ;
        RECT 283.060 1903.990 283.200 1909.710 ;
        RECT 16.660 1903.670 16.920 1903.990 ;
        RECT 283.000 1903.670 283.260 1903.990 ;
        RECT 16.720 1903.165 16.860 1903.670 ;
        RECT 16.650 1902.795 16.930 1903.165 ;
      LAYER via2 ;
        RECT 282.990 1938.200 283.270 1938.480 ;
        RECT 16.650 1902.840 16.930 1903.120 ;
      LAYER met3 ;
        RECT 300.000 1941.160 304.000 1941.760 ;
        RECT 300.230 1939.170 300.530 1941.160 ;
        RECT 284.590 1938.870 300.530 1939.170 ;
        RECT 282.965 1938.490 283.295 1938.505 ;
        RECT 284.590 1938.490 284.890 1938.870 ;
        RECT 282.965 1938.190 284.890 1938.490 ;
        RECT 282.965 1938.175 283.295 1938.190 ;
        RECT -4.800 1903.130 2.400 1903.580 ;
        RECT 16.625 1903.130 16.955 1903.145 ;
        RECT -4.800 1902.830 16.955 1903.130 ;
        RECT -4.800 1902.380 2.400 1902.830 ;
        RECT 16.625 1902.815 16.955 1902.830 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 283.430 620.740 283.750 620.800 ;
        RECT 2900.830 620.740 2901.150 620.800 ;
        RECT 283.430 620.600 2901.150 620.740 ;
        RECT 283.430 620.540 283.750 620.600 ;
        RECT 2900.830 620.540 2901.150 620.600 ;
      LAYER via ;
        RECT 283.460 620.540 283.720 620.800 ;
        RECT 2900.860 620.540 2901.120 620.800 ;
      LAYER met2 ;
        RECT 283.450 1088.835 283.730 1089.205 ;
        RECT 283.520 620.830 283.660 1088.835 ;
        RECT 283.460 620.510 283.720 620.830 ;
        RECT 2900.860 620.510 2901.120 620.830 ;
        RECT 2900.920 615.925 2901.060 620.510 ;
        RECT 2900.850 615.555 2901.130 615.925 ;
      LAYER via2 ;
        RECT 283.450 1088.880 283.730 1089.160 ;
        RECT 2900.850 615.600 2901.130 615.880 ;
      LAYER met3 ;
        RECT 283.425 1089.170 283.755 1089.185 ;
        RECT 283.425 1089.040 300.380 1089.170 ;
        RECT 283.425 1088.870 304.000 1089.040 ;
        RECT 283.425 1088.855 283.755 1088.870 ;
        RECT 300.000 1088.440 304.000 1088.870 ;
        RECT 2900.825 615.890 2901.155 615.905 ;
        RECT 2917.600 615.890 2924.800 616.340 ;
        RECT 2900.825 615.590 2924.800 615.890 ;
        RECT 2900.825 615.575 2901.155 615.590 ;
        RECT 2917.600 615.140 2924.800 615.590 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 20.310 1973.600 20.630 1973.660 ;
        RECT 282.510 1973.600 282.830 1973.660 ;
        RECT 20.310 1973.460 282.830 1973.600 ;
        RECT 20.310 1973.400 20.630 1973.460 ;
        RECT 282.510 1973.400 282.830 1973.460 ;
      LAYER via ;
        RECT 20.340 1973.400 20.600 1973.660 ;
        RECT 282.540 1973.400 282.800 1973.660 ;
      LAYER met2 ;
        RECT 20.340 1973.370 20.600 1973.690 ;
        RECT 282.530 1973.515 282.810 1973.885 ;
        RECT 282.540 1973.370 282.800 1973.515 ;
        RECT 20.400 1615.525 20.540 1973.370 ;
        RECT 20.330 1615.155 20.610 1615.525 ;
      LAYER via2 ;
        RECT 282.530 1973.560 282.810 1973.840 ;
        RECT 20.330 1615.200 20.610 1615.480 ;
      LAYER met3 ;
        RECT 282.505 1973.850 282.835 1973.865 ;
        RECT 282.505 1973.720 300.380 1973.850 ;
        RECT 282.505 1973.550 304.000 1973.720 ;
        RECT 282.505 1973.535 282.835 1973.550 ;
        RECT 300.000 1973.120 304.000 1973.550 ;
        RECT -4.800 1615.490 2.400 1615.940 ;
        RECT 20.305 1615.490 20.635 1615.505 ;
        RECT -4.800 1615.190 20.635 1615.490 ;
        RECT -4.800 1614.740 2.400 1615.190 ;
        RECT 20.305 1615.175 20.635 1615.190 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 175.790 2001.140 176.110 2001.200 ;
        RECT 283.430 2001.140 283.750 2001.200 ;
        RECT 175.790 2001.000 283.750 2001.140 ;
        RECT 175.790 2000.940 176.110 2001.000 ;
        RECT 283.430 2000.940 283.750 2001.000 ;
        RECT 17.090 1400.700 17.410 1400.760 ;
        RECT 175.790 1400.700 176.110 1400.760 ;
        RECT 17.090 1400.560 176.110 1400.700 ;
        RECT 17.090 1400.500 17.410 1400.560 ;
        RECT 175.790 1400.500 176.110 1400.560 ;
      LAYER via ;
        RECT 175.820 2000.940 176.080 2001.200 ;
        RECT 283.460 2000.940 283.720 2001.200 ;
        RECT 17.120 1400.500 17.380 1400.760 ;
        RECT 175.820 1400.500 176.080 1400.760 ;
      LAYER met2 ;
        RECT 283.450 2004.795 283.730 2005.165 ;
        RECT 283.520 2001.230 283.660 2004.795 ;
        RECT 175.820 2000.910 176.080 2001.230 ;
        RECT 283.460 2000.910 283.720 2001.230 ;
        RECT 175.880 1400.790 176.020 2000.910 ;
        RECT 17.120 1400.645 17.380 1400.790 ;
        RECT 17.110 1400.275 17.390 1400.645 ;
        RECT 175.820 1400.470 176.080 1400.790 ;
      LAYER via2 ;
        RECT 283.450 2004.840 283.730 2005.120 ;
        RECT 17.110 1400.320 17.390 1400.600 ;
      LAYER met3 ;
        RECT 283.425 2005.130 283.755 2005.145 ;
        RECT 283.425 2005.000 300.380 2005.130 ;
        RECT 283.425 2004.830 304.000 2005.000 ;
        RECT 283.425 2004.815 283.755 2004.830 ;
        RECT 300.000 2004.400 304.000 2004.830 ;
        RECT -4.800 1400.610 2.400 1401.060 ;
        RECT 17.085 1400.610 17.415 1400.625 ;
        RECT -4.800 1400.310 17.415 1400.610 ;
        RECT -4.800 1399.860 2.400 1400.310 ;
        RECT 17.085 1400.295 17.415 1400.310 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 189.590 2035.820 189.910 2035.880 ;
        RECT 285.730 2035.820 286.050 2035.880 ;
        RECT 189.590 2035.680 286.050 2035.820 ;
        RECT 189.590 2035.620 189.910 2035.680 ;
        RECT 285.730 2035.620 286.050 2035.680 ;
        RECT 17.090 1186.840 17.410 1186.900 ;
        RECT 189.590 1186.840 189.910 1186.900 ;
        RECT 17.090 1186.700 189.910 1186.840 ;
        RECT 17.090 1186.640 17.410 1186.700 ;
        RECT 189.590 1186.640 189.910 1186.700 ;
      LAYER via ;
        RECT 189.620 2035.620 189.880 2035.880 ;
        RECT 285.760 2035.620 286.020 2035.880 ;
        RECT 17.120 1186.640 17.380 1186.900 ;
        RECT 189.620 1186.640 189.880 1186.900 ;
      LAYER met2 ;
        RECT 285.750 2036.755 286.030 2037.125 ;
        RECT 285.820 2035.910 285.960 2036.755 ;
        RECT 189.620 2035.590 189.880 2035.910 ;
        RECT 285.760 2035.590 286.020 2035.910 ;
        RECT 189.680 1186.930 189.820 2035.590 ;
        RECT 17.120 1186.610 17.380 1186.930 ;
        RECT 189.620 1186.610 189.880 1186.930 ;
        RECT 17.180 1185.085 17.320 1186.610 ;
        RECT 17.110 1184.715 17.390 1185.085 ;
      LAYER via2 ;
        RECT 285.750 2036.800 286.030 2037.080 ;
        RECT 17.110 1184.760 17.390 1185.040 ;
      LAYER met3 ;
        RECT 285.725 2037.090 286.055 2037.105 ;
        RECT 285.725 2036.960 300.380 2037.090 ;
        RECT 285.725 2036.790 304.000 2036.960 ;
        RECT 285.725 2036.775 286.055 2036.790 ;
        RECT 300.000 2036.360 304.000 2036.790 ;
        RECT -4.800 1185.050 2.400 1185.500 ;
        RECT 17.085 1185.050 17.415 1185.065 ;
        RECT -4.800 1184.750 17.415 1185.050 ;
        RECT -4.800 1184.300 2.400 1184.750 ;
        RECT 17.085 1184.735 17.415 1184.750 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 265.490 2063.360 265.810 2063.420 ;
        RECT 285.730 2063.360 286.050 2063.420 ;
        RECT 265.490 2063.220 286.050 2063.360 ;
        RECT 265.490 2063.160 265.810 2063.220 ;
        RECT 285.730 2063.160 286.050 2063.220 ;
        RECT 15.710 972.640 16.030 972.700 ;
        RECT 265.490 972.640 265.810 972.700 ;
        RECT 15.710 972.500 265.810 972.640 ;
        RECT 15.710 972.440 16.030 972.500 ;
        RECT 265.490 972.440 265.810 972.500 ;
      LAYER via ;
        RECT 265.520 2063.160 265.780 2063.420 ;
        RECT 285.760 2063.160 286.020 2063.420 ;
        RECT 15.740 972.440 16.000 972.700 ;
        RECT 265.520 972.440 265.780 972.700 ;
      LAYER met2 ;
        RECT 285.750 2068.035 286.030 2068.405 ;
        RECT 285.820 2063.450 285.960 2068.035 ;
        RECT 265.520 2063.130 265.780 2063.450 ;
        RECT 285.760 2063.130 286.020 2063.450 ;
        RECT 265.580 972.730 265.720 2063.130 ;
        RECT 15.740 972.410 16.000 972.730 ;
        RECT 265.520 972.410 265.780 972.730 ;
        RECT 15.800 969.525 15.940 972.410 ;
        RECT 15.730 969.155 16.010 969.525 ;
      LAYER via2 ;
        RECT 285.750 2068.080 286.030 2068.360 ;
        RECT 15.730 969.200 16.010 969.480 ;
      LAYER met3 ;
        RECT 285.725 2068.370 286.055 2068.385 ;
        RECT 285.725 2068.240 300.380 2068.370 ;
        RECT 285.725 2068.070 304.000 2068.240 ;
        RECT 285.725 2068.055 286.055 2068.070 ;
        RECT 300.000 2067.640 304.000 2068.070 ;
        RECT -4.800 969.490 2.400 969.940 ;
        RECT 15.705 969.490 16.035 969.505 ;
        RECT -4.800 969.190 16.035 969.490 ;
        RECT -4.800 968.740 2.400 969.190 ;
        RECT 15.705 969.175 16.035 969.190 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 99.890 2097.700 100.210 2097.760 ;
        RECT 285.730 2097.700 286.050 2097.760 ;
        RECT 99.890 2097.560 286.050 2097.700 ;
        RECT 99.890 2097.500 100.210 2097.560 ;
        RECT 285.730 2097.500 286.050 2097.560 ;
        RECT 15.710 758.780 16.030 758.840 ;
        RECT 99.890 758.780 100.210 758.840 ;
        RECT 15.710 758.640 100.210 758.780 ;
        RECT 15.710 758.580 16.030 758.640 ;
        RECT 99.890 758.580 100.210 758.640 ;
      LAYER via ;
        RECT 99.920 2097.500 100.180 2097.760 ;
        RECT 285.760 2097.500 286.020 2097.760 ;
        RECT 15.740 758.580 16.000 758.840 ;
        RECT 99.920 758.580 100.180 758.840 ;
      LAYER met2 ;
        RECT 285.750 2099.995 286.030 2100.365 ;
        RECT 285.820 2097.790 285.960 2099.995 ;
        RECT 99.920 2097.470 100.180 2097.790 ;
        RECT 285.760 2097.470 286.020 2097.790 ;
        RECT 99.980 758.870 100.120 2097.470 ;
        RECT 15.740 758.550 16.000 758.870 ;
        RECT 99.920 758.550 100.180 758.870 ;
        RECT 15.800 753.965 15.940 758.550 ;
        RECT 15.730 753.595 16.010 753.965 ;
      LAYER via2 ;
        RECT 285.750 2100.040 286.030 2100.320 ;
        RECT 15.730 753.640 16.010 753.920 ;
      LAYER met3 ;
        RECT 285.725 2100.330 286.055 2100.345 ;
        RECT 285.725 2100.200 300.380 2100.330 ;
        RECT 285.725 2100.030 304.000 2100.200 ;
        RECT 285.725 2100.015 286.055 2100.030 ;
        RECT 300.000 2099.600 304.000 2100.030 ;
        RECT -4.800 753.930 2.400 754.380 ;
        RECT 15.705 753.930 16.035 753.945 ;
        RECT -4.800 753.630 16.035 753.930 ;
        RECT -4.800 753.180 2.400 753.630 ;
        RECT 15.705 753.615 16.035 753.630 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 86.090 2125.580 86.410 2125.640 ;
        RECT 285.730 2125.580 286.050 2125.640 ;
        RECT 86.090 2125.440 286.050 2125.580 ;
        RECT 86.090 2125.380 86.410 2125.440 ;
        RECT 285.730 2125.380 286.050 2125.440 ;
        RECT 16.170 544.920 16.490 544.980 ;
        RECT 86.090 544.920 86.410 544.980 ;
        RECT 16.170 544.780 86.410 544.920 ;
        RECT 16.170 544.720 16.490 544.780 ;
        RECT 86.090 544.720 86.410 544.780 ;
      LAYER via ;
        RECT 86.120 2125.380 86.380 2125.640 ;
        RECT 285.760 2125.380 286.020 2125.640 ;
        RECT 16.200 544.720 16.460 544.980 ;
        RECT 86.120 544.720 86.380 544.980 ;
      LAYER met2 ;
        RECT 285.750 2131.275 286.030 2131.645 ;
        RECT 285.820 2125.670 285.960 2131.275 ;
        RECT 86.120 2125.350 86.380 2125.670 ;
        RECT 285.760 2125.350 286.020 2125.670 ;
        RECT 86.180 545.010 86.320 2125.350 ;
        RECT 16.200 544.690 16.460 545.010 ;
        RECT 86.120 544.690 86.380 545.010 ;
        RECT 16.260 538.405 16.400 544.690 ;
        RECT 16.190 538.035 16.470 538.405 ;
      LAYER via2 ;
        RECT 285.750 2131.320 286.030 2131.600 ;
        RECT 16.190 538.080 16.470 538.360 ;
      LAYER met3 ;
        RECT 285.725 2131.610 286.055 2131.625 ;
        RECT 285.725 2131.480 300.380 2131.610 ;
        RECT 285.725 2131.310 304.000 2131.480 ;
        RECT 285.725 2131.295 286.055 2131.310 ;
        RECT 300.000 2130.880 304.000 2131.310 ;
        RECT -4.800 538.370 2.400 538.820 ;
        RECT 16.165 538.370 16.495 538.385 ;
        RECT -4.800 538.070 16.495 538.370 ;
        RECT -4.800 537.620 2.400 538.070 ;
        RECT 16.165 538.055 16.495 538.070 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 196.490 2159.920 196.810 2159.980 ;
        RECT 283.430 2159.920 283.750 2159.980 ;
        RECT 196.490 2159.780 283.750 2159.920 ;
        RECT 196.490 2159.720 196.810 2159.780 ;
        RECT 283.430 2159.720 283.750 2159.780 ;
        RECT 16.630 324.260 16.950 324.320 ;
        RECT 196.490 324.260 196.810 324.320 ;
        RECT 16.630 324.120 196.810 324.260 ;
        RECT 16.630 324.060 16.950 324.120 ;
        RECT 196.490 324.060 196.810 324.120 ;
      LAYER via ;
        RECT 196.520 2159.720 196.780 2159.980 ;
        RECT 283.460 2159.720 283.720 2159.980 ;
        RECT 16.660 324.060 16.920 324.320 ;
        RECT 196.520 324.060 196.780 324.320 ;
      LAYER met2 ;
        RECT 196.520 2159.690 196.780 2160.010 ;
        RECT 283.450 2159.835 283.730 2160.205 ;
        RECT 283.460 2159.690 283.720 2159.835 ;
        RECT 196.580 324.350 196.720 2159.690 ;
        RECT 16.660 324.030 16.920 324.350 ;
        RECT 196.520 324.030 196.780 324.350 ;
        RECT 16.720 322.845 16.860 324.030 ;
        RECT 16.650 322.475 16.930 322.845 ;
      LAYER via2 ;
        RECT 283.450 2159.880 283.730 2160.160 ;
        RECT 16.650 322.520 16.930 322.800 ;
      LAYER met3 ;
        RECT 300.000 2162.840 304.000 2163.440 ;
        RECT 283.425 2160.170 283.755 2160.185 ;
        RECT 300.230 2160.170 300.530 2162.840 ;
        RECT 283.425 2159.870 300.530 2160.170 ;
        RECT 283.425 2159.855 283.755 2159.870 ;
        RECT -4.800 322.810 2.400 323.260 ;
        RECT 16.625 322.810 16.955 322.825 ;
        RECT -4.800 322.510 16.955 322.810 ;
        RECT -4.800 322.060 2.400 322.510 ;
        RECT 16.625 322.495 16.955 322.510 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 244.790 2194.600 245.110 2194.660 ;
        RECT 282.970 2194.600 283.290 2194.660 ;
        RECT 244.790 2194.460 283.290 2194.600 ;
        RECT 244.790 2194.400 245.110 2194.460 ;
        RECT 282.970 2194.400 283.290 2194.460 ;
        RECT 15.710 110.400 16.030 110.460 ;
        RECT 244.790 110.400 245.110 110.460 ;
        RECT 15.710 110.260 245.110 110.400 ;
        RECT 15.710 110.200 16.030 110.260 ;
        RECT 244.790 110.200 245.110 110.260 ;
      LAYER via ;
        RECT 244.820 2194.400 245.080 2194.660 ;
        RECT 283.000 2194.400 283.260 2194.660 ;
        RECT 15.740 110.200 16.000 110.460 ;
        RECT 244.820 110.200 245.080 110.460 ;
      LAYER met2 ;
        RECT 244.820 2194.370 245.080 2194.690 ;
        RECT 282.990 2194.515 283.270 2194.885 ;
        RECT 283.000 2194.370 283.260 2194.515 ;
        RECT 244.880 110.490 245.020 2194.370 ;
        RECT 15.740 110.170 16.000 110.490 ;
        RECT 244.820 110.170 245.080 110.490 ;
        RECT 15.800 107.285 15.940 110.170 ;
        RECT 15.730 106.915 16.010 107.285 ;
      LAYER via2 ;
        RECT 282.990 2194.560 283.270 2194.840 ;
        RECT 15.730 106.960 16.010 107.240 ;
      LAYER met3 ;
        RECT 282.965 2194.850 283.295 2194.865 ;
        RECT 282.965 2194.720 300.380 2194.850 ;
        RECT 282.965 2194.550 304.000 2194.720 ;
        RECT 282.965 2194.535 283.295 2194.550 ;
        RECT 300.000 2194.120 304.000 2194.550 ;
        RECT -4.800 107.250 2.400 107.700 ;
        RECT 15.705 107.250 16.035 107.265 ;
        RECT -4.800 106.950 16.035 107.250 ;
        RECT -4.800 106.500 2.400 106.950 ;
        RECT 15.705 106.935 16.035 106.950 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 287.110 855.340 287.430 855.400 ;
        RECT 2900.830 855.340 2901.150 855.400 ;
        RECT 287.110 855.200 2901.150 855.340 ;
        RECT 287.110 855.140 287.430 855.200 ;
        RECT 2900.830 855.140 2901.150 855.200 ;
      LAYER via ;
        RECT 287.140 855.140 287.400 855.400 ;
        RECT 2900.860 855.140 2901.120 855.400 ;
      LAYER met2 ;
        RECT 287.130 1120.795 287.410 1121.165 ;
        RECT 287.200 855.430 287.340 1120.795 ;
        RECT 287.140 855.110 287.400 855.430 ;
        RECT 2900.860 855.110 2901.120 855.430 ;
        RECT 2900.920 850.525 2901.060 855.110 ;
        RECT 2900.850 850.155 2901.130 850.525 ;
      LAYER via2 ;
        RECT 287.130 1120.840 287.410 1121.120 ;
        RECT 2900.850 850.200 2901.130 850.480 ;
      LAYER met3 ;
        RECT 287.105 1121.130 287.435 1121.145 ;
        RECT 287.105 1121.000 300.380 1121.130 ;
        RECT 287.105 1120.830 304.000 1121.000 ;
        RECT 287.105 1120.815 287.435 1120.830 ;
        RECT 300.000 1120.400 304.000 1120.830 ;
        RECT 2900.825 850.490 2901.155 850.505 ;
        RECT 2917.600 850.490 2924.800 850.940 ;
        RECT 2900.825 850.190 2924.800 850.490 ;
        RECT 2900.825 850.175 2901.155 850.190 ;
        RECT 2917.600 849.740 2924.800 850.190 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 284.810 1003.920 285.130 1003.980 ;
        RECT 2899.910 1003.920 2900.230 1003.980 ;
        RECT 284.810 1003.780 2900.230 1003.920 ;
        RECT 284.810 1003.720 285.130 1003.780 ;
        RECT 2899.910 1003.720 2900.230 1003.780 ;
      LAYER via ;
        RECT 284.840 1003.720 285.100 1003.980 ;
        RECT 2899.940 1003.720 2900.200 1003.980 ;
      LAYER met2 ;
        RECT 285.290 1152.075 285.570 1152.445 ;
        RECT 285.360 1027.210 285.500 1152.075 ;
        RECT 2899.930 1084.755 2900.210 1085.125 ;
        RECT 284.900 1027.070 285.500 1027.210 ;
        RECT 284.900 1004.010 285.040 1027.070 ;
        RECT 2900.000 1004.010 2900.140 1084.755 ;
        RECT 284.840 1003.690 285.100 1004.010 ;
        RECT 2899.940 1003.690 2900.200 1004.010 ;
      LAYER via2 ;
        RECT 285.290 1152.120 285.570 1152.400 ;
        RECT 2899.930 1084.800 2900.210 1085.080 ;
      LAYER met3 ;
        RECT 285.265 1152.410 285.595 1152.425 ;
        RECT 285.265 1152.280 300.380 1152.410 ;
        RECT 285.265 1152.110 304.000 1152.280 ;
        RECT 285.265 1152.095 285.595 1152.110 ;
        RECT 300.000 1151.680 304.000 1152.110 ;
        RECT 2899.905 1085.090 2900.235 1085.105 ;
        RECT 2917.600 1085.090 2924.800 1085.540 ;
        RECT 2899.905 1084.790 2924.800 1085.090 ;
        RECT 2899.905 1084.775 2900.235 1084.790 ;
        RECT 2917.600 1084.340 2924.800 1084.790 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 288.030 1000.180 288.350 1000.240 ;
        RECT 2904.510 1000.180 2904.830 1000.240 ;
        RECT 288.030 1000.040 2904.830 1000.180 ;
        RECT 288.030 999.980 288.350 1000.040 ;
        RECT 2904.510 999.980 2904.830 1000.040 ;
      LAYER via ;
        RECT 288.060 999.980 288.320 1000.240 ;
        RECT 2904.540 999.980 2904.800 1000.240 ;
      LAYER met2 ;
        RECT 2904.530 1319.355 2904.810 1319.725 ;
        RECT 288.050 1184.035 288.330 1184.405 ;
        RECT 288.120 1000.270 288.260 1184.035 ;
        RECT 2904.600 1000.270 2904.740 1319.355 ;
        RECT 288.060 999.950 288.320 1000.270 ;
        RECT 2904.540 999.950 2904.800 1000.270 ;
      LAYER via2 ;
        RECT 2904.530 1319.400 2904.810 1319.680 ;
        RECT 288.050 1184.080 288.330 1184.360 ;
      LAYER met3 ;
        RECT 2904.505 1319.690 2904.835 1319.705 ;
        RECT 2917.600 1319.690 2924.800 1320.140 ;
        RECT 2904.505 1319.390 2924.800 1319.690 ;
        RECT 2904.505 1319.375 2904.835 1319.390 ;
        RECT 2917.600 1318.940 2924.800 1319.390 ;
        RECT 288.025 1184.370 288.355 1184.385 ;
        RECT 288.025 1184.240 300.380 1184.370 ;
        RECT 288.025 1184.070 304.000 1184.240 ;
        RECT 288.025 1184.055 288.355 1184.070 ;
        RECT 300.000 1183.640 304.000 1184.070 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 284.350 999.840 284.670 999.900 ;
        RECT 2903.130 999.840 2903.450 999.900 ;
        RECT 284.350 999.700 2903.450 999.840 ;
        RECT 284.350 999.640 284.670 999.700 ;
        RECT 2903.130 999.640 2903.450 999.700 ;
      LAYER via ;
        RECT 284.380 999.640 284.640 999.900 ;
        RECT 2903.160 999.640 2903.420 999.900 ;
      LAYER met2 ;
        RECT 2903.150 1553.955 2903.430 1554.325 ;
        RECT 284.370 1215.315 284.650 1215.685 ;
        RECT 284.440 999.930 284.580 1215.315 ;
        RECT 2903.220 999.930 2903.360 1553.955 ;
        RECT 284.380 999.610 284.640 999.930 ;
        RECT 2903.160 999.610 2903.420 999.930 ;
      LAYER via2 ;
        RECT 2903.150 1554.000 2903.430 1554.280 ;
        RECT 284.370 1215.360 284.650 1215.640 ;
      LAYER met3 ;
        RECT 2903.125 1554.290 2903.455 1554.305 ;
        RECT 2917.600 1554.290 2924.800 1554.740 ;
        RECT 2903.125 1553.990 2924.800 1554.290 ;
        RECT 2903.125 1553.975 2903.455 1553.990 ;
        RECT 2917.600 1553.540 2924.800 1553.990 ;
        RECT 284.345 1215.650 284.675 1215.665 ;
        RECT 284.345 1215.520 300.380 1215.650 ;
        RECT 284.345 1215.350 304.000 1215.520 ;
        RECT 284.345 1215.335 284.675 1215.350 ;
        RECT 300.000 1214.920 304.000 1215.350 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 299.070 1002.220 299.390 1002.280 ;
        RECT 2901.750 1002.220 2902.070 1002.280 ;
        RECT 299.070 1002.080 2902.070 1002.220 ;
        RECT 299.070 1002.020 299.390 1002.080 ;
        RECT 2901.750 1002.020 2902.070 1002.080 ;
      LAYER via ;
        RECT 299.100 1002.020 299.360 1002.280 ;
        RECT 2901.780 1002.020 2902.040 1002.280 ;
      LAYER met2 ;
        RECT 2901.770 1789.235 2902.050 1789.605 ;
        RECT 299.090 1024.915 299.370 1025.285 ;
        RECT 299.160 1002.310 299.300 1024.915 ;
        RECT 2901.840 1002.310 2901.980 1789.235 ;
        RECT 299.100 1001.990 299.360 1002.310 ;
        RECT 2901.780 1001.990 2902.040 1002.310 ;
      LAYER via2 ;
        RECT 2901.770 1789.280 2902.050 1789.560 ;
        RECT 299.090 1024.960 299.370 1025.240 ;
      LAYER met3 ;
        RECT 2901.745 1789.570 2902.075 1789.585 ;
        RECT 2917.600 1789.570 2924.800 1790.020 ;
        RECT 2901.745 1789.270 2924.800 1789.570 ;
        RECT 2901.745 1789.255 2902.075 1789.270 ;
        RECT 2917.600 1788.820 2924.800 1789.270 ;
        RECT 288.230 1247.610 288.610 1247.620 ;
        RECT 288.230 1247.480 300.380 1247.610 ;
        RECT 288.230 1247.310 304.000 1247.480 ;
        RECT 288.230 1247.300 288.610 1247.310 ;
        RECT 300.000 1246.880 304.000 1247.310 ;
        RECT 288.230 1025.250 288.610 1025.260 ;
        RECT 299.065 1025.250 299.395 1025.265 ;
        RECT 288.230 1024.950 299.395 1025.250 ;
        RECT 288.230 1024.940 288.610 1024.950 ;
        RECT 299.065 1024.935 299.395 1024.950 ;
      LAYER via3 ;
        RECT 288.260 1247.300 288.580 1247.620 ;
        RECT 288.260 1024.940 288.580 1025.260 ;
      LAYER met4 ;
        RECT 288.255 1247.295 288.585 1247.625 ;
        RECT 288.270 1025.265 288.570 1247.295 ;
        RECT 288.255 1024.935 288.585 1025.265 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 299.990 2190.180 300.310 2190.240 ;
        RECT 2901.750 2190.180 2902.070 2190.240 ;
        RECT 299.990 2190.040 2902.070 2190.180 ;
        RECT 299.990 2189.980 300.310 2190.040 ;
        RECT 2901.750 2189.980 2902.070 2190.040 ;
        RECT 288.950 1597.560 289.270 1597.620 ;
        RECT 299.990 1597.560 300.310 1597.620 ;
        RECT 288.950 1597.420 300.310 1597.560 ;
        RECT 288.950 1597.360 289.270 1597.420 ;
        RECT 299.990 1597.360 300.310 1597.420 ;
      LAYER via ;
        RECT 300.020 2189.980 300.280 2190.240 ;
        RECT 2901.780 2189.980 2902.040 2190.240 ;
        RECT 288.980 1597.360 289.240 1597.620 ;
        RECT 300.020 1597.360 300.280 1597.620 ;
      LAYER met2 ;
        RECT 300.020 2189.950 300.280 2190.270 ;
        RECT 2901.780 2189.950 2902.040 2190.270 ;
        RECT 300.080 1597.650 300.220 2189.950 ;
        RECT 2901.840 2024.205 2901.980 2189.950 ;
        RECT 2901.770 2023.835 2902.050 2024.205 ;
        RECT 288.980 1597.330 289.240 1597.650 ;
        RECT 300.020 1597.330 300.280 1597.650 ;
        RECT 289.040 1278.925 289.180 1597.330 ;
        RECT 288.970 1278.555 289.250 1278.925 ;
      LAYER via2 ;
        RECT 2901.770 2023.880 2902.050 2024.160 ;
        RECT 288.970 1278.600 289.250 1278.880 ;
      LAYER met3 ;
        RECT 2901.745 2024.170 2902.075 2024.185 ;
        RECT 2917.600 2024.170 2924.800 2024.620 ;
        RECT 2901.745 2023.870 2924.800 2024.170 ;
        RECT 2901.745 2023.855 2902.075 2023.870 ;
        RECT 2917.600 2023.420 2924.800 2023.870 ;
        RECT 288.945 1278.890 289.275 1278.905 ;
        RECT 288.945 1278.760 300.380 1278.890 ;
        RECT 288.945 1278.590 304.000 1278.760 ;
        RECT 288.945 1278.575 289.275 1278.590 ;
        RECT 300.000 1278.160 304.000 1278.590 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 288.030 2256.480 288.350 2256.540 ;
        RECT 2900.830 2256.480 2901.150 2256.540 ;
        RECT 288.030 2256.340 2901.150 2256.480 ;
        RECT 288.030 2256.280 288.350 2256.340 ;
        RECT 2900.830 2256.280 2901.150 2256.340 ;
      LAYER via ;
        RECT 288.060 2256.280 288.320 2256.540 ;
        RECT 2900.860 2256.280 2901.120 2256.540 ;
      LAYER met2 ;
        RECT 2900.850 2258.435 2901.130 2258.805 ;
        RECT 2900.920 2256.570 2901.060 2258.435 ;
        RECT 288.060 2256.250 288.320 2256.570 ;
        RECT 2900.860 2256.250 2901.120 2256.570 ;
        RECT 288.120 1310.205 288.260 2256.250 ;
        RECT 288.050 1309.835 288.330 1310.205 ;
      LAYER via2 ;
        RECT 2900.850 2258.480 2901.130 2258.760 ;
        RECT 288.050 1309.880 288.330 1310.160 ;
      LAYER met3 ;
        RECT 2900.825 2258.770 2901.155 2258.785 ;
        RECT 2917.600 2258.770 2924.800 2259.220 ;
        RECT 2900.825 2258.470 2924.800 2258.770 ;
        RECT 2900.825 2258.455 2901.155 2258.470 ;
        RECT 2917.600 2258.020 2924.800 2258.470 ;
        RECT 288.025 1310.170 288.355 1310.185 ;
        RECT 288.025 1310.040 300.380 1310.170 ;
        RECT 288.025 1309.870 304.000 1310.040 ;
        RECT 288.025 1309.855 288.355 1309.870 ;
        RECT 300.000 1309.440 304.000 1309.870 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 633.030 26.080 633.350 26.140 ;
        RECT 1428.370 26.080 1428.690 26.140 ;
        RECT 633.030 25.940 1428.690 26.080 ;
        RECT 633.030 25.880 633.350 25.940 ;
        RECT 1428.370 25.880 1428.690 25.940 ;
      LAYER via ;
        RECT 633.060 25.880 633.320 26.140 ;
        RECT 1428.400 25.880 1428.660 26.140 ;
      LAYER met2 ;
        RECT 1430.770 1000.690 1431.050 1004.000 ;
        RECT 1428.460 1000.550 1431.050 1000.690 ;
        RECT 1428.460 26.170 1428.600 1000.550 ;
        RECT 1430.770 1000.000 1431.050 1000.550 ;
        RECT 633.060 25.850 633.320 26.170 ;
        RECT 1428.400 25.850 1428.660 26.170 ;
        RECT 633.120 2.400 633.260 25.850 ;
        RECT 632.910 -4.800 633.470 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2417.250 -4.800 2417.810 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2434.730 -4.800 2435.290 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2452.670 -4.800 2453.230 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2470.610 -4.800 2471.170 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2488.550 -4.800 2489.110 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2506.030 -4.800 2506.590 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2523.970 -4.800 2524.530 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2541.910 -4.800 2542.470 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2559.850 -4.800 2560.410 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2577.790 -4.800 2578.350 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 811.390 -4.800 811.950 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2595.270 -4.800 2595.830 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2613.210 -4.800 2613.770 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2631.150 -4.800 2631.710 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2649.090 -4.800 2649.650 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2667.030 -4.800 2667.590 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2684.510 -4.800 2685.070 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2702.450 -4.800 2703.010 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2720.390 -4.800 2720.950 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2738.330 -4.800 2738.890 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2755.810 -4.800 2756.370 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 829.330 -4.800 829.890 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2773.750 -4.800 2774.310 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2791.690 -4.800 2792.250 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2809.630 -4.800 2810.190 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2827.570 -4.800 2828.130 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2845.050 -4.800 2845.610 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2862.990 -4.800 2863.550 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2880.930 -4.800 2881.490 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 846.810 -4.800 847.370 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 864.750 -4.800 865.310 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 882.690 -4.800 883.250 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 900.630 -4.800 901.190 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 918.570 -4.800 919.130 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 936.050 -4.800 936.610 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1455.970 25.400 1456.290 25.460 ;
        RECT 652.440 25.260 1456.290 25.400 ;
        RECT 650.970 25.060 651.290 25.120 ;
        RECT 652.440 25.060 652.580 25.260 ;
        RECT 1455.970 25.200 1456.290 25.260 ;
        RECT 650.970 24.920 652.580 25.060 ;
        RECT 650.970 24.860 651.290 24.920 ;
      LAYER via ;
        RECT 651.000 24.860 651.260 25.120 ;
        RECT 1456.000 25.200 1456.260 25.460 ;
      LAYER met2 ;
        RECT 1462.510 1000.690 1462.790 1004.000 ;
        RECT 1456.060 1000.550 1462.790 1000.690 ;
        RECT 1456.060 25.490 1456.200 1000.550 ;
        RECT 1462.510 1000.000 1462.790 1000.550 ;
        RECT 1456.000 25.170 1456.260 25.490 ;
        RECT 651.000 24.830 651.260 25.150 ;
        RECT 651.060 2.400 651.200 24.830 ;
        RECT 650.850 -4.800 651.410 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 989.870 -4.800 990.430 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1043.230 -4.800 1043.790 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1061.170 -4.800 1061.730 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1079.110 -4.800 1079.670 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1096.590 -4.800 1097.150 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1114.530 -4.800 1115.090 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1132.470 -4.800 1133.030 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1150.410 -4.800 1150.970 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 668.790 -4.800 669.350 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1168.350 -4.800 1168.910 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1185.830 -4.800 1186.390 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1203.770 -4.800 1204.330 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1221.710 -4.800 1222.270 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1239.650 -4.800 1240.210 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 -4.800 1257.690 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1275.070 -4.800 1275.630 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1293.010 -4.800 1293.570 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1310.950 -4.800 1311.510 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1328.890 -4.800 1329.450 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 686.270 -4.800 686.830 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1346.370 -4.800 1346.930 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1364.310 -4.800 1364.870 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1382.250 -4.800 1382.810 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1400.190 -4.800 1400.750 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1418.130 -4.800 1418.690 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1435.610 -4.800 1436.170 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1453.550 -4.800 1454.110 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1471.490 -4.800 1472.050 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1489.430 -4.800 1489.990 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1506.910 -4.800 1507.470 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 704.210 -4.800 704.770 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1524.850 -4.800 1525.410 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1542.790 -4.800 1543.350 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1560.730 -4.800 1561.290 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1578.670 -4.800 1579.230 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1596.150 -4.800 1596.710 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1614.090 -4.800 1614.650 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1632.030 -4.800 1632.590 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1649.970 -4.800 1650.530 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1667.910 -4.800 1668.470 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1685.390 -4.800 1685.950 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 722.150 -4.800 722.710 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1703.330 -4.800 1703.890 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1721.270 -4.800 1721.830 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1739.210 -4.800 1739.770 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1756.690 -4.800 1757.250 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1774.630 -4.800 1775.190 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1792.570 -4.800 1793.130 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1810.510 -4.800 1811.070 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1828.450 -4.800 1829.010 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1845.930 -4.800 1846.490 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1863.870 -4.800 1864.430 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 740.090 -4.800 740.650 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1881.810 -4.800 1882.370 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1935.170 -4.800 1935.730 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1988.990 -4.800 1989.550 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2024.410 -4.800 2024.970 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2042.350 -4.800 2042.910 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 757.570 -4.800 758.130 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2060.290 -4.800 2060.850 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2078.230 -4.800 2078.790 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2095.710 -4.800 2096.270 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2113.650 -4.800 2114.210 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2131.590 -4.800 2132.150 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2149.530 -4.800 2150.090 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2167.470 -4.800 2168.030 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2184.950 -4.800 2185.510 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2202.890 -4.800 2203.450 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2220.830 -4.800 2221.390 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 775.510 -4.800 776.070 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2238.770 -4.800 2239.330 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2256.250 -4.800 2256.810 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2274.190 -4.800 2274.750 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2292.130 -4.800 2292.690 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2310.070 -4.800 2310.630 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2328.010 -4.800 2328.570 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2345.490 -4.800 2346.050 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2363.430 -4.800 2363.990 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2381.370 -4.800 2381.930 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2399.310 -4.800 2399.870 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 793.450 -4.800 794.010 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 639.010 25.740 639.330 25.800 ;
        RECT 1435.270 25.740 1435.590 25.800 ;
        RECT 639.010 25.600 1435.590 25.740 ;
        RECT 639.010 25.540 639.330 25.600 ;
        RECT 1435.270 25.540 1435.590 25.600 ;
      LAYER via ;
        RECT 639.040 25.540 639.300 25.800 ;
        RECT 1435.300 25.540 1435.560 25.800 ;
      LAYER met2 ;
        RECT 1441.350 1000.690 1441.630 1004.000 ;
        RECT 1435.360 1000.550 1441.630 1000.690 ;
        RECT 1435.360 25.830 1435.500 1000.550 ;
        RECT 1441.350 1000.000 1441.630 1000.550 ;
        RECT 639.040 25.510 639.300 25.830 ;
        RECT 1435.300 25.510 1435.560 25.830 ;
        RECT 639.100 2.400 639.240 25.510 ;
        RECT 638.890 -4.800 639.450 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2422.770 -4.800 2423.330 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2440.710 -4.800 2441.270 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2458.650 -4.800 2459.210 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2476.590 -4.800 2477.150 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2494.530 -4.800 2495.090 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2512.010 -4.800 2512.570 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2529.950 -4.800 2530.510 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2547.890 -4.800 2548.450 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2565.830 -4.800 2566.390 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2583.770 -4.800 2584.330 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 817.370 -4.800 817.930 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2601.250 -4.800 2601.810 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2619.190 -4.800 2619.750 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2637.130 -4.800 2637.690 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2655.070 -4.800 2655.630 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2672.550 -4.800 2673.110 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2690.490 -4.800 2691.050 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2708.430 -4.800 2708.990 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2726.370 -4.800 2726.930 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2744.310 -4.800 2744.870 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2761.790 -4.800 2762.350 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 835.310 -4.800 835.870 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2779.730 -4.800 2780.290 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2797.670 -4.800 2798.230 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2815.610 -4.800 2816.170 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2833.550 -4.800 2834.110 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2851.030 -4.800 2851.590 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2868.970 -4.800 2869.530 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 852.790 -4.800 853.350 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 870.730 -4.800 871.290 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 888.670 -4.800 889.230 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 906.610 -4.800 907.170 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 924.090 -4.800 924.650 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 942.030 -4.800 942.590 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 977.910 -4.800 978.470 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 656.950 24.720 657.270 24.780 ;
        RECT 1469.770 24.720 1470.090 24.780 ;
        RECT 656.950 24.580 1470.090 24.720 ;
        RECT 656.950 24.520 657.270 24.580 ;
        RECT 1469.770 24.520 1470.090 24.580 ;
      LAYER via ;
        RECT 656.980 24.520 657.240 24.780 ;
        RECT 1469.800 24.520 1470.060 24.780 ;
      LAYER met2 ;
        RECT 1473.090 1000.690 1473.370 1004.000 ;
        RECT 1469.860 1000.550 1473.370 1000.690 ;
        RECT 1469.860 24.810 1470.000 1000.550 ;
        RECT 1473.090 1000.000 1473.370 1000.550 ;
        RECT 656.980 24.490 657.240 24.810 ;
        RECT 1469.800 24.490 1470.060 24.810 ;
        RECT 657.040 2.400 657.180 24.490 ;
        RECT 656.830 -4.800 657.390 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 995.850 -4.800 996.410 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1031.270 -4.800 1031.830 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1049.210 -4.800 1049.770 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1067.150 -4.800 1067.710 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1085.090 -4.800 1085.650 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1102.570 -4.800 1103.130 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1120.510 -4.800 1121.070 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1138.450 -4.800 1139.010 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1156.390 -4.800 1156.950 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 674.430 24.380 674.750 24.440 ;
        RECT 1490.470 24.380 1490.790 24.440 ;
        RECT 674.430 24.240 1490.790 24.380 ;
        RECT 674.430 24.180 674.750 24.240 ;
        RECT 1490.470 24.180 1490.790 24.240 ;
      LAYER via ;
        RECT 674.460 24.180 674.720 24.440 ;
        RECT 1490.500 24.180 1490.760 24.440 ;
      LAYER met2 ;
        RECT 1494.250 1000.690 1494.530 1004.000 ;
        RECT 1490.560 1000.550 1494.530 1000.690 ;
        RECT 1490.560 24.470 1490.700 1000.550 ;
        RECT 1494.250 1000.000 1494.530 1000.550 ;
        RECT 674.460 24.150 674.720 24.470 ;
        RECT 1490.500 24.150 1490.760 24.470 ;
        RECT 674.520 2.400 674.660 24.150 ;
        RECT 674.310 -4.800 674.870 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1173.870 -4.800 1174.430 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1191.810 -4.800 1192.370 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1209.750 -4.800 1210.310 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1227.690 -4.800 1228.250 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1245.630 -4.800 1246.190 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1263.110 -4.800 1263.670 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1281.050 -4.800 1281.610 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1298.990 -4.800 1299.550 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1316.930 -4.800 1317.490 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1334.870 -4.800 1335.430 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 692.250 -4.800 692.810 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1352.350 -4.800 1352.910 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1370.290 -4.800 1370.850 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1388.230 -4.800 1388.790 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1406.170 -4.800 1406.730 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1423.650 -4.800 1424.210 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1441.590 -4.800 1442.150 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1459.530 -4.800 1460.090 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1477.470 -4.800 1478.030 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1495.410 -4.800 1495.970 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1512.890 -4.800 1513.450 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 710.190 -4.800 710.750 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1530.830 -4.800 1531.390 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1548.770 -4.800 1549.330 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1566.710 -4.800 1567.270 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1584.650 -4.800 1585.210 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1602.130 -4.800 1602.690 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1620.070 -4.800 1620.630 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1638.010 -4.800 1638.570 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1655.950 -4.800 1656.510 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1673.430 -4.800 1673.990 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1691.370 -4.800 1691.930 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 728.130 -4.800 728.690 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1709.310 -4.800 1709.870 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1727.250 -4.800 1727.810 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1745.190 -4.800 1745.750 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1762.670 -4.800 1763.230 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1780.610 -4.800 1781.170 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1798.550 -4.800 1799.110 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1816.490 -4.800 1817.050 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1834.430 -4.800 1834.990 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1851.910 -4.800 1852.470 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1869.850 -4.800 1870.410 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 746.070 -4.800 746.630 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1887.790 -4.800 1888.350 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1923.210 -4.800 1923.770 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1977.030 -4.800 1977.590 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1994.970 -4.800 1995.530 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2030.390 -4.800 2030.950 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2048.330 -4.800 2048.890 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 763.550 -4.800 764.110 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2066.270 -4.800 2066.830 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2084.210 -4.800 2084.770 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2101.690 -4.800 2102.250 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2119.630 -4.800 2120.190 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2137.570 -4.800 2138.130 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2155.510 -4.800 2156.070 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2172.990 -4.800 2173.550 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2190.930 -4.800 2191.490 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2208.870 -4.800 2209.430 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2226.810 -4.800 2227.370 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 781.490 -4.800 782.050 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2244.750 -4.800 2245.310 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2262.230 -4.800 2262.790 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2280.170 -4.800 2280.730 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2298.110 -4.800 2298.670 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2316.050 -4.800 2316.610 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2333.990 -4.800 2334.550 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2351.470 -4.800 2352.030 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2369.410 -4.800 2369.970 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2387.350 -4.800 2387.910 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2405.290 -4.800 2405.850 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 799.430 -4.800 799.990 2.400 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1449.070 25.060 1449.390 25.120 ;
        RECT 652.900 24.920 1449.390 25.060 ;
        RECT 644.990 24.720 645.310 24.780 ;
        RECT 652.900 24.720 653.040 24.920 ;
        RECT 1449.070 24.860 1449.390 24.920 ;
        RECT 644.990 24.580 653.040 24.720 ;
        RECT 644.990 24.520 645.310 24.580 ;
      LAYER via ;
        RECT 645.020 24.520 645.280 24.780 ;
        RECT 1449.100 24.860 1449.360 25.120 ;
      LAYER met2 ;
        RECT 1451.930 1000.690 1452.210 1004.000 ;
        RECT 1449.160 1000.550 1452.210 1000.690 ;
        RECT 1449.160 25.150 1449.300 1000.550 ;
        RECT 1451.930 1000.000 1452.210 1000.550 ;
        RECT 1449.100 24.830 1449.360 25.150 ;
        RECT 645.020 24.490 645.280 24.810 ;
        RECT 645.080 2.400 645.220 24.490 ;
        RECT 644.870 -4.800 645.430 2.400 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2428.750 -4.800 2429.310 2.400 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2446.690 -4.800 2447.250 2.400 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2464.630 -4.800 2465.190 2.400 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2482.570 -4.800 2483.130 2.400 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2500.510 -4.800 2501.070 2.400 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2517.990 -4.800 2518.550 2.400 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2535.930 -4.800 2536.490 2.400 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2553.870 -4.800 2554.430 2.400 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2571.810 -4.800 2572.370 2.400 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2589.290 -4.800 2589.850 2.400 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 823.350 -4.800 823.910 2.400 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2607.230 -4.800 2607.790 2.400 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2625.170 -4.800 2625.730 2.400 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2643.110 -4.800 2643.670 2.400 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2661.050 -4.800 2661.610 2.400 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2678.530 -4.800 2679.090 2.400 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2696.470 -4.800 2697.030 2.400 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2714.410 -4.800 2714.970 2.400 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2732.350 -4.800 2732.910 2.400 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2750.290 -4.800 2750.850 2.400 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2767.770 -4.800 2768.330 2.400 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 840.830 -4.800 841.390 2.400 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2785.710 -4.800 2786.270 2.400 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2803.650 -4.800 2804.210 2.400 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2821.590 -4.800 2822.150 2.400 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2839.070 -4.800 2839.630 2.400 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2857.010 -4.800 2857.570 2.400 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2874.950 -4.800 2875.510 2.400 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 858.770 -4.800 859.330 2.400 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 876.710 -4.800 877.270 2.400 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 894.650 -4.800 895.210 2.400 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 912.590 -4.800 913.150 2.400 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 930.070 -4.800 930.630 2.400 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 948.010 -4.800 948.570 2.400 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 983.890 -4.800 984.450 2.400 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 662.930 24.040 663.250 24.100 ;
        RECT 1483.570 24.040 1483.890 24.100 ;
        RECT 662.930 23.900 1483.890 24.040 ;
        RECT 662.930 23.840 663.250 23.900 ;
        RECT 1483.570 23.840 1483.890 23.900 ;
      LAYER via ;
        RECT 662.960 23.840 663.220 24.100 ;
        RECT 1483.600 23.840 1483.860 24.100 ;
      LAYER met2 ;
        RECT 1483.670 1000.620 1483.950 1004.000 ;
        RECT 1483.660 1000.000 1483.950 1000.620 ;
        RECT 1483.660 24.130 1483.800 1000.000 ;
        RECT 662.960 23.810 663.220 24.130 ;
        RECT 1483.600 23.810 1483.860 24.130 ;
        RECT 663.020 2.400 663.160 23.810 ;
        RECT 662.810 -4.800 663.370 2.400 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1001.830 -4.800 1002.390 2.400 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1037.250 -4.800 1037.810 2.400 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1055.190 -4.800 1055.750 2.400 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1073.130 -4.800 1073.690 2.400 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1090.610 -4.800 1091.170 2.400 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1108.550 -4.800 1109.110 2.400 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1126.490 -4.800 1127.050 2.400 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1144.430 -4.800 1144.990 2.400 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1162.370 -4.800 1162.930 2.400 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 680.290 -4.800 680.850 2.400 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1179.850 -4.800 1180.410 2.400 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1197.790 -4.800 1198.350 2.400 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1215.730 -4.800 1216.290 2.400 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1233.670 -4.800 1234.230 2.400 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1251.610 -4.800 1252.170 2.400 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1269.090 -4.800 1269.650 2.400 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1287.030 -4.800 1287.590 2.400 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1304.970 -4.800 1305.530 2.400 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1322.910 -4.800 1323.470 2.400 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1340.390 -4.800 1340.950 2.400 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 698.230 -4.800 698.790 2.400 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1358.330 -4.800 1358.890 2.400 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1376.270 -4.800 1376.830 2.400 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1394.210 -4.800 1394.770 2.400 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1412.150 -4.800 1412.710 2.400 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1429.630 -4.800 1430.190 2.400 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1447.570 -4.800 1448.130 2.400 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1465.510 -4.800 1466.070 2.400 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1483.450 -4.800 1484.010 2.400 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1501.390 -4.800 1501.950 2.400 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1518.870 -4.800 1519.430 2.400 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 716.170 -4.800 716.730 2.400 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1536.810 -4.800 1537.370 2.400 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1554.750 -4.800 1555.310 2.400 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1572.690 -4.800 1573.250 2.400 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1590.170 -4.800 1590.730 2.400 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1608.110 -4.800 1608.670 2.400 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1626.050 -4.800 1626.610 2.400 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1643.990 -4.800 1644.550 2.400 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1661.930 -4.800 1662.490 2.400 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1679.410 -4.800 1679.970 2.400 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1697.350 -4.800 1697.910 2.400 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 734.110 -4.800 734.670 2.400 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1715.290 -4.800 1715.850 2.400 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1733.230 -4.800 1733.790 2.400 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1751.170 -4.800 1751.730 2.400 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1768.650 -4.800 1769.210 2.400 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1786.590 -4.800 1787.150 2.400 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1804.530 -4.800 1805.090 2.400 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1822.470 -4.800 1823.030 2.400 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1839.950 -4.800 1840.510 2.400 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1857.890 -4.800 1858.450 2.400 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1875.830 -4.800 1876.390 2.400 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 752.050 -4.800 752.610 2.400 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1893.770 -4.800 1894.330 2.400 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1929.190 -4.800 1929.750 2.400 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1983.010 -4.800 1983.570 2.400 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2000.950 -4.800 2001.510 2.400 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2018.430 -4.800 2018.990 2.400 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2036.370 -4.800 2036.930 2.400 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2054.310 -4.800 2054.870 2.400 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 769.530 -4.800 770.090 2.400 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2072.250 -4.800 2072.810 2.400 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2089.730 -4.800 2090.290 2.400 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2107.670 -4.800 2108.230 2.400 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2125.610 -4.800 2126.170 2.400 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2143.550 -4.800 2144.110 2.400 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2161.490 -4.800 2162.050 2.400 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2178.970 -4.800 2179.530 2.400 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2196.910 -4.800 2197.470 2.400 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2214.850 -4.800 2215.410 2.400 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2232.790 -4.800 2233.350 2.400 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 787.470 -4.800 788.030 2.400 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2250.730 -4.800 2251.290 2.400 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2268.210 -4.800 2268.770 2.400 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2286.150 -4.800 2286.710 2.400 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2304.090 -4.800 2304.650 2.400 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2322.030 -4.800 2322.590 2.400 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2339.510 -4.800 2340.070 2.400 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2357.450 -4.800 2358.010 2.400 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2375.390 -4.800 2375.950 2.400 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2393.330 -4.800 2393.890 2.400 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2411.270 -4.800 2411.830 2.400 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 805.410 -4.800 805.970 2.400 ;
    END
  END la_oen[9]
  PIN user_clock2
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 303.670 2287.420 303.990 2287.480 ;
        RECT 318.390 2287.420 318.710 2287.480 ;
        RECT 969.290 2287.420 969.610 2287.480 ;
        RECT 1568.670 2287.420 1568.990 2287.480 ;
        RECT 2214.970 2287.420 2215.290 2287.480 ;
        RECT 303.670 2287.280 2215.290 2287.420 ;
        RECT 303.670 2287.220 303.990 2287.280 ;
        RECT 318.390 2287.220 318.710 2287.280 ;
        RECT 969.290 2287.220 969.610 2287.280 ;
        RECT 1568.670 2287.220 1568.990 2287.280 ;
        RECT 2214.970 2287.220 2215.290 2287.280 ;
        RECT 2.830 15.540 3.150 15.600 ;
        RECT 303.670 15.540 303.990 15.600 ;
        RECT 2.830 15.400 303.990 15.540 ;
        RECT 2.830 15.340 3.150 15.400 ;
        RECT 303.670 15.340 303.990 15.400 ;
      LAYER via ;
        RECT 303.700 2287.220 303.960 2287.480 ;
        RECT 318.420 2287.220 318.680 2287.480 ;
        RECT 969.320 2287.220 969.580 2287.480 ;
        RECT 1568.700 2287.220 1568.960 2287.480 ;
        RECT 2215.000 2287.220 2215.260 2287.480 ;
        RECT 2.860 15.340 3.120 15.600 ;
        RECT 303.700 15.340 303.960 15.600 ;
      LAYER met2 ;
        RECT 969.310 2290.395 969.590 2290.765 ;
        RECT 1568.690 2290.395 1568.970 2290.765 ;
        RECT 318.410 2287.675 318.690 2288.045 ;
        RECT 318.480 2287.510 318.620 2287.675 ;
        RECT 969.380 2287.510 969.520 2290.395 ;
        RECT 1568.760 2287.510 1568.900 2290.395 ;
        RECT 2214.990 2289.715 2215.270 2290.085 ;
        RECT 2215.060 2287.510 2215.200 2289.715 ;
        RECT 303.700 2287.190 303.960 2287.510 ;
        RECT 318.420 2287.190 318.680 2287.510 ;
        RECT 969.320 2287.190 969.580 2287.510 ;
        RECT 1568.700 2287.190 1568.960 2287.510 ;
        RECT 2215.000 2287.190 2215.260 2287.510 ;
        RECT 303.760 1003.410 303.900 2287.190 ;
        RECT 305.150 1003.410 305.430 1004.000 ;
        RECT 303.760 1003.270 305.430 1003.410 ;
        RECT 303.760 15.630 303.900 1003.270 ;
        RECT 305.150 1000.000 305.430 1003.270 ;
        RECT 2.860 15.310 3.120 15.630 ;
        RECT 303.700 15.310 303.960 15.630 ;
        RECT 2.920 2.400 3.060 15.310 ;
        RECT 2.710 -4.800 3.270 2.400 ;
      LAYER via2 ;
        RECT 969.310 2290.440 969.590 2290.720 ;
        RECT 1568.690 2290.440 1568.970 2290.720 ;
        RECT 318.410 2287.720 318.690 2288.000 ;
        RECT 2214.990 2289.760 2215.270 2290.040 ;
      LAYER met3 ;
        RECT 969.285 2290.740 969.615 2290.745 ;
        RECT 969.030 2290.730 969.615 2290.740 ;
        RECT 968.830 2290.430 969.615 2290.730 ;
        RECT 969.030 2290.420 969.615 2290.430 ;
        RECT 969.285 2290.415 969.615 2290.420 ;
        RECT 1568.665 2290.740 1568.995 2290.745 ;
        RECT 1568.665 2290.730 1569.250 2290.740 ;
        RECT 1568.665 2290.430 1569.450 2290.730 ;
        RECT 1568.665 2290.420 1569.250 2290.430 ;
        RECT 1568.665 2290.415 1568.995 2290.420 ;
        RECT 2214.965 2290.050 2215.295 2290.065 ;
        RECT 2215.630 2290.050 2216.010 2290.060 ;
        RECT 2214.965 2289.750 2216.010 2290.050 ;
        RECT 2214.965 2289.735 2215.295 2289.750 ;
        RECT 2215.630 2289.740 2216.010 2289.750 ;
        RECT 318.385 2288.020 318.715 2288.025 ;
        RECT 318.385 2288.010 318.970 2288.020 ;
        RECT 318.385 2287.710 319.170 2288.010 ;
        RECT 318.385 2287.700 318.970 2287.710 ;
        RECT 318.385 2287.695 318.715 2287.700 ;
      LAYER via3 ;
        RECT 969.060 2290.420 969.380 2290.740 ;
        RECT 1568.900 2290.420 1569.220 2290.740 ;
        RECT 2215.660 2289.740 2215.980 2290.060 ;
        RECT 318.620 2287.700 318.940 2288.020 ;
      LAYER met4 ;
        RECT 319.015 2296.850 319.315 2304.600 ;
        RECT 318.630 2296.550 319.315 2296.850 ;
        RECT 969.015 2296.850 969.315 2304.600 ;
        RECT 1569.015 2296.850 1569.315 2304.600 ;
        RECT 2219.015 2301.950 2219.315 2304.600 ;
        RECT 969.015 2296.550 969.370 2296.850 ;
        RECT 318.630 2288.025 318.930 2296.550 ;
        RECT 969.070 2290.745 969.370 2296.550 ;
        RECT 1568.910 2296.550 1569.315 2296.850 ;
        RECT 2215.670 2301.650 2219.315 2301.950 ;
        RECT 1568.910 2290.745 1569.210 2296.550 ;
        RECT 969.055 2290.415 969.385 2290.745 ;
        RECT 1568.895 2290.415 1569.225 2290.745 ;
        RECT 2215.670 2290.065 2215.970 2301.650 ;
        RECT 2219.015 2300.000 2219.315 2301.650 ;
        RECT 2215.655 2289.735 2215.985 2290.065 ;
        RECT 318.615 2287.695 318.945 2288.025 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 311.030 15.540 311.350 15.600 ;
        RECT 305.600 15.400 311.350 15.540 ;
        RECT 8.350 15.200 8.670 15.260 ;
        RECT 305.600 15.200 305.740 15.400 ;
        RECT 311.030 15.340 311.350 15.400 ;
        RECT 8.350 15.060 305.740 15.200 ;
        RECT 8.350 15.000 8.670 15.060 ;
      LAYER via ;
        RECT 8.380 15.000 8.640 15.260 ;
        RECT 311.060 15.340 311.320 15.600 ;
      LAYER met2 ;
        RECT 315.730 1000.690 316.010 1004.000 ;
        RECT 311.120 1000.550 316.010 1000.690 ;
        RECT 311.120 15.630 311.260 1000.550 ;
        RECT 315.730 1000.000 316.010 1000.550 ;
        RECT 311.060 15.310 311.320 15.630 ;
        RECT 8.380 14.970 8.640 15.290 ;
        RECT 8.440 2.400 8.580 14.970 ;
        RECT 8.230 -4.800 8.790 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 14.330 15.880 14.650 15.940 ;
        RECT 324.830 15.880 325.150 15.940 ;
        RECT 14.330 15.740 325.150 15.880 ;
        RECT 14.330 15.680 14.650 15.740 ;
        RECT 324.830 15.680 325.150 15.740 ;
      LAYER via ;
        RECT 14.360 15.680 14.620 15.940 ;
        RECT 324.860 15.680 325.120 15.940 ;
      LAYER met2 ;
        RECT 326.310 1000.690 326.590 1004.000 ;
        RECT 324.920 1000.550 326.590 1000.690 ;
        RECT 324.920 15.970 325.060 1000.550 ;
        RECT 326.310 1000.000 326.590 1000.550 ;
        RECT 14.360 15.650 14.620 15.970 ;
        RECT 324.860 15.650 325.120 15.970 ;
        RECT 14.420 2.400 14.560 15.650 ;
        RECT 14.210 -4.800 14.770 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 38.250 16.900 38.570 16.960 ;
        RECT 325.750 16.900 326.070 16.960 ;
        RECT 38.250 16.760 326.070 16.900 ;
        RECT 38.250 16.700 38.570 16.760 ;
        RECT 325.750 16.700 326.070 16.760 ;
        RECT 325.750 16.220 326.070 16.280 ;
        RECT 365.770 16.220 366.090 16.280 ;
        RECT 325.750 16.080 366.090 16.220 ;
        RECT 325.750 16.020 326.070 16.080 ;
        RECT 365.770 16.020 366.090 16.080 ;
      LAYER via ;
        RECT 38.280 16.700 38.540 16.960 ;
        RECT 325.780 16.700 326.040 16.960 ;
        RECT 325.780 16.020 326.040 16.280 ;
        RECT 365.800 16.020 366.060 16.280 ;
      LAYER met2 ;
        RECT 368.630 1000.690 368.910 1004.000 ;
        RECT 365.860 1000.550 368.910 1000.690 ;
        RECT 38.280 16.670 38.540 16.990 ;
        RECT 325.780 16.670 326.040 16.990 ;
        RECT 38.340 2.400 38.480 16.670 ;
        RECT 325.840 16.310 325.980 16.670 ;
        RECT 365.860 16.310 366.000 1000.550 ;
        RECT 368.630 1000.000 368.910 1000.550 ;
        RECT 325.780 15.990 326.040 16.310 ;
        RECT 365.800 15.990 366.060 16.310 ;
        RECT 38.130 -4.800 38.690 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 241.110 21.320 241.430 21.380 ;
        RECT 724.570 21.320 724.890 21.380 ;
        RECT 241.110 21.180 724.890 21.320 ;
        RECT 241.110 21.120 241.430 21.180 ;
        RECT 724.570 21.120 724.890 21.180 ;
      LAYER via ;
        RECT 241.140 21.120 241.400 21.380 ;
        RECT 724.600 21.120 724.860 21.380 ;
      LAYER met2 ;
        RECT 729.730 1000.690 730.010 1004.000 ;
        RECT 724.660 1000.550 730.010 1000.690 ;
        RECT 724.660 21.410 724.800 1000.550 ;
        RECT 729.730 1000.000 730.010 1000.550 ;
        RECT 241.140 21.090 241.400 21.410 ;
        RECT 724.600 21.090 724.860 21.410 ;
        RECT 241.200 10.610 241.340 21.090 ;
        RECT 240.740 10.470 241.340 10.610 ;
        RECT 240.740 2.400 240.880 10.470 ;
        RECT 240.530 -4.800 241.090 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 258.130 21.660 258.450 21.720 ;
        RECT 759.070 21.660 759.390 21.720 ;
        RECT 258.130 21.520 759.390 21.660 ;
        RECT 258.130 21.460 258.450 21.520 ;
        RECT 759.070 21.460 759.390 21.520 ;
      LAYER via ;
        RECT 258.160 21.460 258.420 21.720 ;
        RECT 759.100 21.460 759.360 21.720 ;
      LAYER met2 ;
        RECT 761.470 1000.690 761.750 1004.000 ;
        RECT 759.160 1000.550 761.750 1000.690 ;
        RECT 759.160 21.750 759.300 1000.550 ;
        RECT 761.470 1000.000 761.750 1000.550 ;
        RECT 258.160 21.430 258.420 21.750 ;
        RECT 759.100 21.430 759.360 21.750 ;
        RECT 258.220 2.400 258.360 21.430 ;
        RECT 258.010 -4.800 258.570 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 276.070 22.000 276.390 22.060 ;
        RECT 793.570 22.000 793.890 22.060 ;
        RECT 276.070 21.860 793.890 22.000 ;
        RECT 276.070 21.800 276.390 21.860 ;
        RECT 793.570 21.800 793.890 21.860 ;
      LAYER via ;
        RECT 276.100 21.800 276.360 22.060 ;
        RECT 793.600 21.800 793.860 22.060 ;
      LAYER met2 ;
        RECT 793.670 1000.620 793.950 1004.000 ;
        RECT 793.660 1000.000 793.950 1000.620 ;
        RECT 793.660 22.090 793.800 1000.000 ;
        RECT 276.100 21.770 276.360 22.090 ;
        RECT 793.600 21.770 793.860 22.090 ;
        RECT 276.160 2.400 276.300 21.770 ;
        RECT 275.950 -4.800 276.510 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 294.010 22.340 294.330 22.400 ;
        RECT 821.170 22.340 821.490 22.400 ;
        RECT 294.010 22.200 821.490 22.340 ;
        RECT 294.010 22.140 294.330 22.200 ;
        RECT 821.170 22.140 821.490 22.200 ;
      LAYER via ;
        RECT 294.040 22.140 294.300 22.400 ;
        RECT 821.200 22.140 821.460 22.400 ;
      LAYER met2 ;
        RECT 825.410 1000.690 825.690 1004.000 ;
        RECT 821.260 1000.550 825.690 1000.690 ;
        RECT 821.260 22.430 821.400 1000.550 ;
        RECT 825.410 1000.000 825.690 1000.550 ;
        RECT 294.040 22.110 294.300 22.430 ;
        RECT 821.200 22.110 821.460 22.430 ;
        RECT 294.100 2.400 294.240 22.110 ;
        RECT 293.890 -4.800 294.450 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 311.950 22.680 312.270 22.740 ;
        RECT 855.670 22.680 855.990 22.740 ;
        RECT 311.950 22.540 855.990 22.680 ;
        RECT 311.950 22.480 312.270 22.540 ;
        RECT 855.670 22.480 855.990 22.540 ;
      LAYER via ;
        RECT 311.980 22.480 312.240 22.740 ;
        RECT 855.700 22.480 855.960 22.740 ;
      LAYER met2 ;
        RECT 857.150 1000.690 857.430 1004.000 ;
        RECT 855.760 1000.550 857.430 1000.690 ;
        RECT 855.760 22.770 855.900 1000.550 ;
        RECT 857.150 1000.000 857.430 1000.550 ;
        RECT 311.980 22.450 312.240 22.770 ;
        RECT 855.700 22.450 855.960 22.770 ;
        RECT 312.040 2.400 312.180 22.450 ;
        RECT 311.830 -4.800 312.390 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 329.890 23.020 330.210 23.080 ;
        RECT 883.270 23.020 883.590 23.080 ;
        RECT 329.890 22.880 883.590 23.020 ;
        RECT 329.890 22.820 330.210 22.880 ;
        RECT 883.270 22.820 883.590 22.880 ;
      LAYER via ;
        RECT 329.920 22.820 330.180 23.080 ;
        RECT 883.300 22.820 883.560 23.080 ;
      LAYER met2 ;
        RECT 888.890 1000.690 889.170 1004.000 ;
        RECT 883.360 1000.550 889.170 1000.690 ;
        RECT 883.360 23.110 883.500 1000.550 ;
        RECT 888.890 1000.000 889.170 1000.550 ;
        RECT 329.920 22.790 330.180 23.110 ;
        RECT 883.300 22.790 883.560 23.110 ;
        RECT 329.980 2.400 330.120 22.790 ;
        RECT 329.770 -4.800 330.330 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 347.370 23.360 347.690 23.420 ;
        RECT 917.770 23.360 918.090 23.420 ;
        RECT 347.370 23.220 918.090 23.360 ;
        RECT 347.370 23.160 347.690 23.220 ;
        RECT 917.770 23.160 918.090 23.220 ;
      LAYER via ;
        RECT 347.400 23.160 347.660 23.420 ;
        RECT 917.800 23.160 918.060 23.420 ;
      LAYER met2 ;
        RECT 921.090 1000.690 921.370 1004.000 ;
        RECT 917.860 1000.550 921.370 1000.690 ;
        RECT 917.860 23.450 918.000 1000.550 ;
        RECT 921.090 1000.000 921.370 1000.550 ;
        RECT 347.400 23.130 347.660 23.450 ;
        RECT 917.800 23.130 918.060 23.450 ;
        RECT 347.460 2.400 347.600 23.130 ;
        RECT 347.250 -4.800 347.810 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 365.310 23.700 365.630 23.760 ;
        RECT 952.270 23.700 952.590 23.760 ;
        RECT 365.310 23.560 952.590 23.700 ;
        RECT 365.310 23.500 365.630 23.560 ;
        RECT 952.270 23.500 952.590 23.560 ;
      LAYER via ;
        RECT 365.340 23.500 365.600 23.760 ;
        RECT 952.300 23.500 952.560 23.760 ;
      LAYER met2 ;
        RECT 952.830 1000.690 953.110 1004.000 ;
        RECT 952.360 1000.550 953.110 1000.690 ;
        RECT 952.360 23.790 952.500 1000.550 ;
        RECT 952.830 1000.000 953.110 1000.550 ;
        RECT 365.340 23.470 365.600 23.790 ;
        RECT 952.300 23.470 952.560 23.790 ;
        RECT 365.400 2.400 365.540 23.470 ;
        RECT 365.190 -4.800 365.750 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 383.250 27.440 383.570 27.500 ;
        RECT 979.870 27.440 980.190 27.500 ;
        RECT 383.250 27.300 980.190 27.440 ;
        RECT 383.250 27.240 383.570 27.300 ;
        RECT 979.870 27.240 980.190 27.300 ;
      LAYER via ;
        RECT 383.280 27.240 383.540 27.500 ;
        RECT 979.900 27.240 980.160 27.500 ;
      LAYER met2 ;
        RECT 984.570 1000.690 984.850 1004.000 ;
        RECT 979.960 1000.550 984.850 1000.690 ;
        RECT 979.960 27.530 980.100 1000.550 ;
        RECT 984.570 1000.000 984.850 1000.550 ;
        RECT 383.280 27.210 383.540 27.530 ;
        RECT 979.900 27.210 980.160 27.530 ;
        RECT 383.340 2.400 383.480 27.210 ;
        RECT 383.130 -4.800 383.690 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1016.310 1000.690 1016.590 1004.000 ;
        RECT 1014.460 1000.550 1016.590 1000.690 ;
        RECT 1014.460 26.365 1014.600 1000.550 ;
        RECT 1016.310 1000.000 1016.590 1000.550 ;
        RECT 401.210 25.995 401.490 26.365 ;
        RECT 1014.390 25.995 1014.670 26.365 ;
        RECT 401.280 2.400 401.420 25.995 ;
        RECT 401.070 -4.800 401.630 2.400 ;
      LAYER via2 ;
        RECT 401.210 26.040 401.490 26.320 ;
        RECT 1014.390 26.040 1014.670 26.320 ;
      LAYER met3 ;
        RECT 401.185 26.330 401.515 26.345 ;
        RECT 1014.365 26.330 1014.695 26.345 ;
        RECT 401.185 26.030 1014.695 26.330 ;
        RECT 401.185 26.015 401.515 26.030 ;
        RECT 1014.365 26.015 1014.695 26.030 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 62.170 27.100 62.490 27.160 ;
        RECT 407.170 27.100 407.490 27.160 ;
        RECT 62.170 26.960 407.490 27.100 ;
        RECT 62.170 26.900 62.490 26.960 ;
        RECT 407.170 26.900 407.490 26.960 ;
      LAYER via ;
        RECT 62.200 26.900 62.460 27.160 ;
        RECT 407.200 26.900 407.460 27.160 ;
      LAYER met2 ;
        RECT 410.950 1000.690 411.230 1004.000 ;
        RECT 407.260 1000.550 411.230 1000.690 ;
        RECT 407.260 27.190 407.400 1000.550 ;
        RECT 410.950 1000.000 411.230 1000.550 ;
        RECT 62.200 26.870 62.460 27.190 ;
        RECT 407.200 26.870 407.460 27.190 ;
        RECT 62.260 2.400 62.400 26.870 ;
        RECT 62.050 -4.800 62.610 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 419.130 27.100 419.450 27.160 ;
        RECT 1041.970 27.100 1042.290 27.160 ;
        RECT 419.130 26.960 1042.290 27.100 ;
        RECT 419.130 26.900 419.450 26.960 ;
        RECT 1041.970 26.900 1042.290 26.960 ;
      LAYER via ;
        RECT 419.160 26.900 419.420 27.160 ;
        RECT 1042.000 26.900 1042.260 27.160 ;
      LAYER met2 ;
        RECT 1048.510 1000.690 1048.790 1004.000 ;
        RECT 1042.060 1000.550 1048.790 1000.690 ;
        RECT 1042.060 27.190 1042.200 1000.550 ;
        RECT 1048.510 1000.000 1048.790 1000.550 ;
        RECT 419.160 26.870 419.420 27.190 ;
        RECT 1042.000 26.870 1042.260 27.190 ;
        RECT 419.220 2.400 419.360 26.870 ;
        RECT 419.010 -4.800 419.570 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1080.250 1000.690 1080.530 1004.000 ;
        RECT 1076.560 1000.550 1080.530 1000.690 ;
        RECT 1076.560 25.685 1076.700 1000.550 ;
        RECT 1080.250 1000.000 1080.530 1000.550 ;
        RECT 436.630 25.315 436.910 25.685 ;
        RECT 1076.490 25.315 1076.770 25.685 ;
        RECT 436.700 2.400 436.840 25.315 ;
        RECT 436.490 -4.800 437.050 2.400 ;
      LAYER via2 ;
        RECT 436.630 25.360 436.910 25.640 ;
        RECT 1076.490 25.360 1076.770 25.640 ;
      LAYER met3 ;
        RECT 436.605 25.650 436.935 25.665 ;
        RECT 1076.465 25.650 1076.795 25.665 ;
        RECT 436.605 25.350 1076.795 25.650 ;
        RECT 436.605 25.335 436.935 25.350 ;
        RECT 1076.465 25.335 1076.795 25.350 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 455.930 26.760 456.250 26.820 ;
        RECT 1110.970 26.760 1111.290 26.820 ;
        RECT 455.930 26.620 1111.290 26.760 ;
        RECT 455.930 26.560 456.250 26.620 ;
        RECT 1110.970 26.560 1111.290 26.620 ;
      LAYER via ;
        RECT 455.960 26.560 456.220 26.820 ;
        RECT 1111.000 26.560 1111.260 26.820 ;
      LAYER met2 ;
        RECT 1111.990 1000.690 1112.270 1004.000 ;
        RECT 1111.060 1000.550 1112.270 1000.690 ;
        RECT 1111.060 26.850 1111.200 1000.550 ;
        RECT 1111.990 1000.000 1112.270 1000.550 ;
        RECT 455.960 26.530 456.220 26.850 ;
        RECT 1111.000 26.530 1111.260 26.850 ;
        RECT 456.020 26.250 456.160 26.530 ;
        RECT 454.640 26.110 456.160 26.250 ;
        RECT 454.640 2.400 454.780 26.110 ;
        RECT 454.430 -4.800 454.990 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1143.730 1000.690 1144.010 1004.000 ;
        RECT 1138.660 1000.550 1144.010 1000.690 ;
        RECT 1138.660 25.005 1138.800 1000.550 ;
        RECT 1143.730 1000.000 1144.010 1000.550 ;
        RECT 472.510 24.635 472.790 25.005 ;
        RECT 1138.590 24.635 1138.870 25.005 ;
        RECT 472.580 2.400 472.720 24.635 ;
        RECT 472.370 -4.800 472.930 2.400 ;
      LAYER via2 ;
        RECT 472.510 24.680 472.790 24.960 ;
        RECT 1138.590 24.680 1138.870 24.960 ;
      LAYER met3 ;
        RECT 472.485 24.970 472.815 24.985 ;
        RECT 1138.565 24.970 1138.895 24.985 ;
        RECT 472.485 24.670 1138.895 24.970 ;
        RECT 472.485 24.655 472.815 24.670 ;
        RECT 1138.565 24.655 1138.895 24.670 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 532.290 26.420 532.610 26.480 ;
        RECT 1173.070 26.420 1173.390 26.480 ;
        RECT 532.290 26.280 1173.390 26.420 ;
        RECT 532.290 26.220 532.610 26.280 ;
        RECT 1173.070 26.220 1173.390 26.280 ;
        RECT 494.110 26.080 494.430 26.140 ;
        RECT 494.110 25.940 531.600 26.080 ;
        RECT 494.110 25.880 494.430 25.940 ;
        RECT 531.460 25.800 531.600 25.940 ;
        RECT 531.370 25.540 531.690 25.800 ;
      LAYER via ;
        RECT 532.320 26.220 532.580 26.480 ;
        RECT 1173.100 26.220 1173.360 26.480 ;
        RECT 494.140 25.880 494.400 26.140 ;
        RECT 531.400 25.540 531.660 25.800 ;
      LAYER met2 ;
        RECT 1175.930 1000.690 1176.210 1004.000 ;
        RECT 1173.160 1000.550 1176.210 1000.690 ;
        RECT 1173.160 26.510 1173.300 1000.550 ;
        RECT 1175.930 1000.000 1176.210 1000.550 ;
        RECT 532.320 26.190 532.580 26.510 ;
        RECT 1173.100 26.190 1173.360 26.510 ;
        RECT 494.140 25.850 494.400 26.170 ;
        RECT 494.200 13.330 494.340 25.850 ;
        RECT 531.400 25.740 531.660 25.830 ;
        RECT 532.380 25.740 532.520 26.190 ;
        RECT 531.400 25.600 532.520 25.740 ;
        RECT 531.400 25.510 531.660 25.600 ;
        RECT 490.520 13.190 494.340 13.330 ;
        RECT 490.520 2.400 490.660 13.190 ;
        RECT 490.310 -4.800 490.870 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 507.910 32.540 508.230 32.600 ;
        RECT 1207.570 32.540 1207.890 32.600 ;
        RECT 507.910 32.400 1207.890 32.540 ;
        RECT 507.910 32.340 508.230 32.400 ;
        RECT 1207.570 32.340 1207.890 32.400 ;
      LAYER via ;
        RECT 507.940 32.340 508.200 32.600 ;
        RECT 1207.600 32.340 1207.860 32.600 ;
      LAYER met2 ;
        RECT 1207.670 1000.620 1207.950 1004.000 ;
        RECT 1207.660 1000.000 1207.950 1000.620 ;
        RECT 1207.660 32.630 1207.800 1000.000 ;
        RECT 507.940 32.310 508.200 32.630 ;
        RECT 1207.600 32.310 1207.860 32.630 ;
        RECT 508.000 2.400 508.140 32.310 ;
        RECT 507.790 -4.800 508.350 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1239.410 1000.690 1239.690 1004.000 ;
        RECT 1235.260 1000.550 1239.690 1000.690 ;
        RECT 1235.260 24.325 1235.400 1000.550 ;
        RECT 1239.410 1000.000 1239.690 1000.550 ;
        RECT 525.870 23.955 526.150 24.325 ;
        RECT 1235.190 23.955 1235.470 24.325 ;
        RECT 525.940 2.400 526.080 23.955 ;
        RECT 525.730 -4.800 526.290 2.400 ;
      LAYER via2 ;
        RECT 525.870 24.000 526.150 24.280 ;
        RECT 1235.190 24.000 1235.470 24.280 ;
      LAYER met3 ;
        RECT 525.845 24.290 526.175 24.305 ;
        RECT 1235.165 24.290 1235.495 24.305 ;
        RECT 525.845 23.990 1235.495 24.290 ;
        RECT 525.845 23.975 526.175 23.990 ;
        RECT 1235.165 23.975 1235.495 23.990 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 543.790 32.200 544.110 32.260 ;
        RECT 1269.670 32.200 1269.990 32.260 ;
        RECT 543.790 32.060 1269.990 32.200 ;
        RECT 543.790 32.000 544.110 32.060 ;
        RECT 1269.670 32.000 1269.990 32.060 ;
      LAYER via ;
        RECT 543.820 32.000 544.080 32.260 ;
        RECT 1269.700 32.000 1269.960 32.260 ;
      LAYER met2 ;
        RECT 1271.610 1000.690 1271.890 1004.000 ;
        RECT 1269.760 1000.550 1271.890 1000.690 ;
        RECT 1269.760 32.290 1269.900 1000.550 ;
        RECT 1271.610 1000.000 1271.890 1000.550 ;
        RECT 543.820 31.970 544.080 32.290 ;
        RECT 1269.700 31.970 1269.960 32.290 ;
        RECT 543.880 2.400 544.020 31.970 ;
        RECT 543.670 -4.800 544.230 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 561.730 31.860 562.050 31.920 ;
        RECT 1297.270 31.860 1297.590 31.920 ;
        RECT 561.730 31.720 1297.590 31.860 ;
        RECT 561.730 31.660 562.050 31.720 ;
        RECT 1297.270 31.660 1297.590 31.720 ;
      LAYER via ;
        RECT 561.760 31.660 562.020 31.920 ;
        RECT 1297.300 31.660 1297.560 31.920 ;
      LAYER met2 ;
        RECT 1303.350 1000.690 1303.630 1004.000 ;
        RECT 1297.360 1000.550 1303.630 1000.690 ;
        RECT 1297.360 31.950 1297.500 1000.550 ;
        RECT 1303.350 1000.000 1303.630 1000.550 ;
        RECT 561.760 31.630 562.020 31.950 ;
        RECT 1297.300 31.630 1297.560 31.950 ;
        RECT 561.820 2.400 561.960 31.630 ;
        RECT 561.610 -4.800 562.170 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 580.590 31.520 580.910 31.580 ;
        RECT 1331.770 31.520 1332.090 31.580 ;
        RECT 580.590 31.380 1332.090 31.520 ;
        RECT 580.590 31.320 580.910 31.380 ;
        RECT 1331.770 31.320 1332.090 31.380 ;
      LAYER via ;
        RECT 580.620 31.320 580.880 31.580 ;
        RECT 1331.800 31.320 1332.060 31.580 ;
      LAYER met2 ;
        RECT 1335.090 1000.690 1335.370 1004.000 ;
        RECT 1331.860 1000.550 1335.370 1000.690 ;
        RECT 1331.860 31.610 1332.000 1000.550 ;
        RECT 1335.090 1000.000 1335.370 1000.550 ;
        RECT 580.620 31.290 580.880 31.610 ;
        RECT 1331.800 31.290 1332.060 31.610 ;
        RECT 580.680 17.410 580.820 31.290 ;
        RECT 579.760 17.270 580.820 17.410 ;
        RECT 579.760 2.400 579.900 17.270 ;
        RECT 579.550 -4.800 580.110 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 86.090 26.420 86.410 26.480 ;
        RECT 448.570 26.420 448.890 26.480 ;
        RECT 86.090 26.280 448.890 26.420 ;
        RECT 86.090 26.220 86.410 26.280 ;
        RECT 448.570 26.220 448.890 26.280 ;
      LAYER via ;
        RECT 86.120 26.220 86.380 26.480 ;
        RECT 448.600 26.220 448.860 26.480 ;
      LAYER met2 ;
        RECT 453.730 1000.690 454.010 1004.000 ;
        RECT 448.660 1000.550 454.010 1000.690 ;
        RECT 448.660 26.510 448.800 1000.550 ;
        RECT 453.730 1000.000 454.010 1000.550 ;
        RECT 86.120 26.190 86.380 26.510 ;
        RECT 448.600 26.190 448.860 26.510 ;
        RECT 86.180 2.400 86.320 26.190 ;
        RECT 85.970 -4.800 86.530 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 597.150 31.180 597.470 31.240 ;
        RECT 1366.270 31.180 1366.590 31.240 ;
        RECT 597.150 31.040 1366.590 31.180 ;
        RECT 597.150 30.980 597.470 31.040 ;
        RECT 1366.270 30.980 1366.590 31.040 ;
      LAYER via ;
        RECT 597.180 30.980 597.440 31.240 ;
        RECT 1366.300 30.980 1366.560 31.240 ;
      LAYER met2 ;
        RECT 1366.830 1000.690 1367.110 1004.000 ;
        RECT 1366.360 1000.550 1367.110 1000.690 ;
        RECT 1366.360 31.270 1366.500 1000.550 ;
        RECT 1366.830 1000.000 1367.110 1000.550 ;
        RECT 597.180 30.950 597.440 31.270 ;
        RECT 1366.300 30.950 1366.560 31.270 ;
        RECT 597.240 2.400 597.380 30.950 ;
        RECT 597.030 -4.800 597.590 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 615.090 30.840 615.410 30.900 ;
        RECT 1393.870 30.840 1394.190 30.900 ;
        RECT 615.090 30.700 1394.190 30.840 ;
        RECT 615.090 30.640 615.410 30.700 ;
        RECT 1393.870 30.640 1394.190 30.700 ;
      LAYER via ;
        RECT 615.120 30.640 615.380 30.900 ;
        RECT 1393.900 30.640 1394.160 30.900 ;
      LAYER met2 ;
        RECT 1399.030 1000.690 1399.310 1004.000 ;
        RECT 1393.960 1000.550 1399.310 1000.690 ;
        RECT 1393.960 30.930 1394.100 1000.550 ;
        RECT 1399.030 1000.000 1399.310 1000.550 ;
        RECT 615.120 30.610 615.380 30.930 ;
        RECT 1393.900 30.610 1394.160 30.930 ;
        RECT 615.180 2.400 615.320 30.610 ;
        RECT 614.970 -4.800 615.530 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 110.010 26.080 110.330 26.140 ;
        RECT 489.970 26.080 490.290 26.140 ;
        RECT 110.010 25.940 490.290 26.080 ;
        RECT 110.010 25.880 110.330 25.940 ;
        RECT 489.970 25.880 490.290 25.940 ;
      LAYER via ;
        RECT 110.040 25.880 110.300 26.140 ;
        RECT 490.000 25.880 490.260 26.140 ;
      LAYER met2 ;
        RECT 496.050 1000.690 496.330 1004.000 ;
        RECT 490.060 1000.550 496.330 1000.690 ;
        RECT 490.060 26.170 490.200 1000.550 ;
        RECT 496.050 1000.000 496.330 1000.550 ;
        RECT 110.040 25.850 110.300 26.170 ;
        RECT 490.000 25.850 490.260 26.170 ;
        RECT 110.100 13.330 110.240 25.850 ;
        RECT 109.640 13.190 110.240 13.330 ;
        RECT 109.640 2.400 109.780 13.190 ;
        RECT 109.430 -4.800 109.990 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 521.250 26.420 521.570 26.480 ;
        RECT 521.250 26.280 532.060 26.420 ;
        RECT 521.250 26.220 521.570 26.280 ;
        RECT 531.920 26.080 532.060 26.280 ;
        RECT 538.270 26.080 538.590 26.140 ;
        RECT 531.920 25.940 538.590 26.080 ;
        RECT 538.270 25.880 538.590 25.940 ;
        RECT 133.470 25.740 133.790 25.800 ;
        RECT 520.330 25.740 520.650 25.800 ;
        RECT 133.470 25.600 520.650 25.740 ;
        RECT 133.470 25.540 133.790 25.600 ;
        RECT 520.330 25.540 520.650 25.600 ;
      LAYER via ;
        RECT 521.280 26.220 521.540 26.480 ;
        RECT 538.300 25.880 538.560 26.140 ;
        RECT 133.500 25.540 133.760 25.800 ;
        RECT 520.360 25.540 520.620 25.800 ;
      LAYER met2 ;
        RECT 538.370 1000.620 538.650 1004.000 ;
        RECT 538.360 1000.000 538.650 1000.620 ;
        RECT 520.420 26.790 521.480 26.930 ;
        RECT 520.420 25.830 520.560 26.790 ;
        RECT 521.340 26.510 521.480 26.790 ;
        RECT 521.280 26.190 521.540 26.510 ;
        RECT 538.360 26.170 538.500 1000.000 ;
        RECT 538.300 25.850 538.560 26.170 ;
        RECT 133.500 25.510 133.760 25.830 ;
        RECT 520.360 25.510 520.620 25.830 ;
        RECT 133.560 2.400 133.700 25.510 ;
        RECT 133.350 -4.800 133.910 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 151.410 25.060 151.730 25.120 ;
        RECT 565.870 25.060 566.190 25.120 ;
        RECT 151.410 24.920 566.190 25.060 ;
        RECT 151.410 24.860 151.730 24.920 ;
        RECT 565.870 24.860 566.190 24.920 ;
      LAYER via ;
        RECT 151.440 24.860 151.700 25.120 ;
        RECT 565.900 24.860 566.160 25.120 ;
      LAYER met2 ;
        RECT 570.570 1000.690 570.850 1004.000 ;
        RECT 565.960 1000.550 570.850 1000.690 ;
        RECT 565.960 25.150 566.100 1000.550 ;
        RECT 570.570 1000.000 570.850 1000.550 ;
        RECT 151.440 24.830 151.700 25.150 ;
        RECT 565.900 24.830 566.160 25.150 ;
        RECT 151.500 2.400 151.640 24.830 ;
        RECT 151.290 -4.800 151.850 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 169.350 24.720 169.670 24.780 ;
        RECT 600.370 24.720 600.690 24.780 ;
        RECT 169.350 24.580 600.690 24.720 ;
        RECT 169.350 24.520 169.670 24.580 ;
        RECT 600.370 24.520 600.690 24.580 ;
      LAYER via ;
        RECT 169.380 24.520 169.640 24.780 ;
        RECT 600.400 24.520 600.660 24.780 ;
      LAYER met2 ;
        RECT 602.310 1000.690 602.590 1004.000 ;
        RECT 600.460 1000.550 602.590 1000.690 ;
        RECT 600.460 24.810 600.600 1000.550 ;
        RECT 602.310 1000.000 602.590 1000.550 ;
        RECT 169.380 24.490 169.640 24.810 ;
        RECT 600.400 24.490 600.660 24.810 ;
        RECT 169.440 2.400 169.580 24.490 ;
        RECT 169.230 -4.800 169.790 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 186.830 24.380 187.150 24.440 ;
        RECT 627.970 24.380 628.290 24.440 ;
        RECT 186.830 24.240 628.290 24.380 ;
        RECT 186.830 24.180 187.150 24.240 ;
        RECT 627.970 24.180 628.290 24.240 ;
      LAYER via ;
        RECT 186.860 24.180 187.120 24.440 ;
        RECT 628.000 24.180 628.260 24.440 ;
      LAYER met2 ;
        RECT 634.050 1000.690 634.330 1004.000 ;
        RECT 628.060 1000.550 634.330 1000.690 ;
        RECT 628.060 24.470 628.200 1000.550 ;
        RECT 634.050 1000.000 634.330 1000.550 ;
        RECT 186.860 24.150 187.120 24.470 ;
        RECT 628.000 24.150 628.260 24.470 ;
        RECT 186.920 2.400 187.060 24.150 ;
        RECT 186.710 -4.800 187.270 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 204.770 24.040 205.090 24.100 ;
        RECT 662.470 24.040 662.790 24.100 ;
        RECT 204.770 23.900 662.790 24.040 ;
        RECT 204.770 23.840 205.090 23.900 ;
        RECT 662.470 23.840 662.790 23.900 ;
      LAYER via ;
        RECT 204.800 23.840 205.060 24.100 ;
        RECT 662.500 23.840 662.760 24.100 ;
      LAYER met2 ;
        RECT 666.250 1000.690 666.530 1004.000 ;
        RECT 662.560 1000.550 666.530 1000.690 ;
        RECT 662.560 24.130 662.700 1000.550 ;
        RECT 666.250 1000.000 666.530 1000.550 ;
        RECT 204.800 23.810 205.060 24.130 ;
        RECT 662.500 23.810 662.760 24.130 ;
        RECT 204.860 2.400 205.000 23.810 ;
        RECT 204.650 -4.800 205.210 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 222.710 20.980 223.030 21.040 ;
        RECT 696.970 20.980 697.290 21.040 ;
        RECT 222.710 20.840 697.290 20.980 ;
        RECT 222.710 20.780 223.030 20.840 ;
        RECT 696.970 20.780 697.290 20.840 ;
      LAYER via ;
        RECT 222.740 20.780 223.000 21.040 ;
        RECT 697.000 20.780 697.260 21.040 ;
      LAYER met2 ;
        RECT 697.990 1000.690 698.270 1004.000 ;
        RECT 697.060 1000.550 698.270 1000.690 ;
        RECT 697.060 21.070 697.200 1000.550 ;
        RECT 697.990 1000.000 698.270 1000.550 ;
        RECT 222.740 20.750 223.000 21.070 ;
        RECT 697.000 20.750 697.260 21.070 ;
        RECT 222.800 2.400 222.940 20.750 ;
        RECT 222.590 -4.800 223.150 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 20.310 16.220 20.630 16.280 ;
        RECT 20.310 16.080 325.520 16.220 ;
        RECT 20.310 16.020 20.630 16.080 ;
        RECT 325.380 15.880 325.520 16.080 ;
        RECT 331.270 15.880 331.590 15.940 ;
        RECT 325.380 15.740 331.590 15.880 ;
        RECT 331.270 15.680 331.590 15.740 ;
      LAYER via ;
        RECT 20.340 16.020 20.600 16.280 ;
        RECT 331.300 15.680 331.560 15.940 ;
      LAYER met2 ;
        RECT 336.890 1000.690 337.170 1004.000 ;
        RECT 331.360 1000.550 337.170 1000.690 ;
        RECT 20.340 15.990 20.600 16.310 ;
        RECT 20.400 2.400 20.540 15.990 ;
        RECT 331.360 15.970 331.500 1000.550 ;
        RECT 336.890 1000.000 337.170 1000.550 ;
        RECT 331.300 15.650 331.560 15.970 ;
        RECT 20.190 -4.800 20.750 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 44.230 20.640 44.550 20.700 ;
        RECT 328.050 20.640 328.370 20.700 ;
        RECT 44.230 20.500 328.370 20.640 ;
        RECT 44.230 20.440 44.550 20.500 ;
        RECT 328.050 20.440 328.370 20.500 ;
        RECT 328.050 16.560 328.370 16.620 ;
        RECT 372.670 16.560 372.990 16.620 ;
        RECT 328.050 16.420 372.990 16.560 ;
        RECT 328.050 16.360 328.370 16.420 ;
        RECT 372.670 16.360 372.990 16.420 ;
      LAYER via ;
        RECT 44.260 20.440 44.520 20.700 ;
        RECT 328.080 20.440 328.340 20.700 ;
        RECT 328.080 16.360 328.340 16.620 ;
        RECT 372.700 16.360 372.960 16.620 ;
      LAYER met2 ;
        RECT 379.210 1000.690 379.490 1004.000 ;
        RECT 372.760 1000.550 379.490 1000.690 ;
        RECT 44.260 20.410 44.520 20.730 ;
        RECT 328.080 20.410 328.340 20.730 ;
        RECT 44.320 2.400 44.460 20.410 ;
        RECT 328.140 16.650 328.280 20.410 ;
        RECT 372.760 16.650 372.900 1000.550 ;
        RECT 379.210 1000.000 379.490 1000.550 ;
        RECT 328.080 16.330 328.340 16.650 ;
        RECT 372.700 16.330 372.960 16.650 ;
        RECT 44.110 -4.800 44.670 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 651.890 987.260 652.210 987.320 ;
        RECT 740.210 987.260 740.530 987.320 ;
        RECT 651.890 987.120 740.530 987.260 ;
        RECT 651.890 987.060 652.210 987.120 ;
        RECT 740.210 987.060 740.530 987.120 ;
        RECT 246.630 25.400 246.950 25.460 ;
        RECT 592.550 25.400 592.870 25.460 ;
        RECT 246.630 25.260 592.870 25.400 ;
        RECT 246.630 25.200 246.950 25.260 ;
        RECT 592.550 25.200 592.870 25.260 ;
        RECT 593.930 25.400 594.250 25.460 ;
        RECT 651.890 25.400 652.210 25.460 ;
        RECT 593.930 25.260 652.210 25.400 ;
        RECT 593.930 25.200 594.250 25.260 ;
        RECT 651.890 25.200 652.210 25.260 ;
      LAYER via ;
        RECT 651.920 987.060 652.180 987.320 ;
        RECT 740.240 987.060 740.500 987.320 ;
        RECT 246.660 25.200 246.920 25.460 ;
        RECT 592.580 25.200 592.840 25.460 ;
        RECT 593.960 25.200 594.220 25.460 ;
        RECT 651.920 25.200 652.180 25.460 ;
      LAYER met2 ;
        RECT 740.310 1000.620 740.590 1004.000 ;
        RECT 740.300 1000.000 740.590 1000.620 ;
        RECT 740.300 987.350 740.440 1000.000 ;
        RECT 651.920 987.030 652.180 987.350 ;
        RECT 740.240 987.030 740.500 987.350 ;
        RECT 592.640 26.110 594.160 26.250 ;
        RECT 592.640 25.490 592.780 26.110 ;
        RECT 594.020 25.490 594.160 26.110 ;
        RECT 651.980 25.490 652.120 987.030 ;
        RECT 246.660 25.170 246.920 25.490 ;
        RECT 592.580 25.170 592.840 25.490 ;
        RECT 593.960 25.170 594.220 25.490 ;
        RECT 651.920 25.170 652.180 25.490 ;
        RECT 246.720 2.400 246.860 25.170 ;
        RECT 246.510 -4.800 247.070 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 264.110 33.560 264.430 33.620 ;
        RECT 765.970 33.560 766.290 33.620 ;
        RECT 264.110 33.420 766.290 33.560 ;
        RECT 264.110 33.360 264.430 33.420 ;
        RECT 765.970 33.360 766.290 33.420 ;
      LAYER via ;
        RECT 264.140 33.360 264.400 33.620 ;
        RECT 766.000 33.360 766.260 33.620 ;
      LAYER met2 ;
        RECT 772.050 1000.690 772.330 1004.000 ;
        RECT 766.060 1000.550 772.330 1000.690 ;
        RECT 766.060 33.650 766.200 1000.550 ;
        RECT 772.050 1000.000 772.330 1000.550 ;
        RECT 264.140 33.330 264.400 33.650 ;
        RECT 766.000 33.330 766.260 33.650 ;
        RECT 264.200 2.400 264.340 33.330 ;
        RECT 263.990 -4.800 264.550 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 638.090 986.920 638.410 986.980 ;
        RECT 804.150 986.920 804.470 986.980 ;
        RECT 638.090 986.780 804.470 986.920 ;
        RECT 638.090 986.720 638.410 986.780 ;
        RECT 804.150 986.720 804.470 986.780 ;
        RECT 400.270 27.780 400.590 27.840 ;
        RECT 382.880 27.640 400.590 27.780 ;
        RECT 327.590 27.440 327.910 27.500 ;
        RECT 382.880 27.440 383.020 27.640 ;
        RECT 400.270 27.580 400.590 27.640 ;
        RECT 519.870 27.780 520.190 27.840 ;
        RECT 547.010 27.780 547.330 27.840 ;
        RECT 519.870 27.640 547.330 27.780 ;
        RECT 519.870 27.580 520.190 27.640 ;
        RECT 547.010 27.580 547.330 27.640 ;
        RECT 327.590 27.300 383.020 27.440 ;
        RECT 327.590 27.240 327.910 27.300 ;
        RECT 400.270 26.760 400.590 26.820 ;
        RECT 400.270 26.620 455.700 26.760 ;
        RECT 400.270 26.560 400.590 26.620 ;
        RECT 455.560 26.420 455.700 26.620 ;
        RECT 519.870 26.420 520.190 26.480 ;
        RECT 455.560 26.280 520.190 26.420 ;
        RECT 519.870 26.220 520.190 26.280 ;
        RECT 547.010 25.740 547.330 25.800 ;
        RECT 593.010 25.740 593.330 25.800 ;
        RECT 547.010 25.600 593.330 25.740 ;
        RECT 547.010 25.540 547.330 25.600 ;
        RECT 593.010 25.540 593.330 25.600 ;
        RECT 594.390 25.060 594.710 25.120 ;
        RECT 638.090 25.060 638.410 25.120 ;
        RECT 594.390 24.920 638.410 25.060 ;
        RECT 594.390 24.860 594.710 24.920 ;
        RECT 638.090 24.860 638.410 24.920 ;
        RECT 282.050 23.700 282.370 23.760 ;
        RECT 327.590 23.700 327.910 23.760 ;
        RECT 282.050 23.560 327.910 23.700 ;
        RECT 282.050 23.500 282.370 23.560 ;
        RECT 327.590 23.500 327.910 23.560 ;
      LAYER via ;
        RECT 638.120 986.720 638.380 986.980 ;
        RECT 804.180 986.720 804.440 986.980 ;
        RECT 327.620 27.240 327.880 27.500 ;
        RECT 400.300 27.580 400.560 27.840 ;
        RECT 519.900 27.580 520.160 27.840 ;
        RECT 547.040 27.580 547.300 27.840 ;
        RECT 400.300 26.560 400.560 26.820 ;
        RECT 519.900 26.220 520.160 26.480 ;
        RECT 547.040 25.540 547.300 25.800 ;
        RECT 593.040 25.540 593.300 25.800 ;
        RECT 594.420 24.860 594.680 25.120 ;
        RECT 638.120 24.860 638.380 25.120 ;
        RECT 282.080 23.500 282.340 23.760 ;
        RECT 327.620 23.500 327.880 23.760 ;
      LAYER met2 ;
        RECT 804.250 1000.620 804.530 1004.000 ;
        RECT 804.240 1000.000 804.530 1000.620 ;
        RECT 804.240 987.010 804.380 1000.000 ;
        RECT 638.120 986.690 638.380 987.010 ;
        RECT 804.180 986.690 804.440 987.010 ;
        RECT 400.300 27.550 400.560 27.870 ;
        RECT 519.900 27.550 520.160 27.870 ;
        RECT 547.040 27.550 547.300 27.870 ;
        RECT 327.620 27.210 327.880 27.530 ;
        RECT 327.680 23.790 327.820 27.210 ;
        RECT 400.360 26.850 400.500 27.550 ;
        RECT 400.300 26.530 400.560 26.850 ;
        RECT 519.960 26.510 520.100 27.550 ;
        RECT 519.900 26.190 520.160 26.510 ;
        RECT 547.100 25.830 547.240 27.550 ;
        RECT 547.040 25.510 547.300 25.830 ;
        RECT 593.040 25.510 593.300 25.830 ;
        RECT 593.100 24.890 593.240 25.510 ;
        RECT 638.180 25.150 638.320 986.690 ;
        RECT 594.420 24.890 594.680 25.150 ;
        RECT 593.100 24.830 594.680 24.890 ;
        RECT 638.120 24.830 638.380 25.150 ;
        RECT 593.100 24.750 594.620 24.830 ;
        RECT 282.080 23.470 282.340 23.790 ;
        RECT 327.620 23.470 327.880 23.790 ;
        RECT 282.140 2.400 282.280 23.470 ;
        RECT 281.930 -4.800 282.490 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 299.990 33.220 300.310 33.280 ;
        RECT 834.970 33.220 835.290 33.280 ;
        RECT 299.990 33.080 835.290 33.220 ;
        RECT 299.990 33.020 300.310 33.080 ;
        RECT 834.970 33.020 835.290 33.080 ;
      LAYER via ;
        RECT 300.020 33.020 300.280 33.280 ;
        RECT 835.000 33.020 835.260 33.280 ;
      LAYER met2 ;
        RECT 835.990 1000.690 836.270 1004.000 ;
        RECT 835.060 1000.550 836.270 1000.690 ;
        RECT 835.060 33.310 835.200 1000.550 ;
        RECT 835.990 1000.000 836.270 1000.550 ;
        RECT 300.020 32.990 300.280 33.310 ;
        RECT 835.000 32.990 835.260 33.310 ;
        RECT 300.080 2.400 300.220 32.990 ;
        RECT 299.870 -4.800 300.430 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 317.930 32.880 318.250 32.940 ;
        RECT 862.570 32.880 862.890 32.940 ;
        RECT 317.930 32.740 862.890 32.880 ;
        RECT 317.930 32.680 318.250 32.740 ;
        RECT 862.570 32.680 862.890 32.740 ;
      LAYER via ;
        RECT 317.960 32.680 318.220 32.940 ;
        RECT 862.600 32.680 862.860 32.940 ;
      LAYER met2 ;
        RECT 867.730 1000.690 868.010 1004.000 ;
        RECT 862.660 1000.550 868.010 1000.690 ;
        RECT 862.660 32.970 862.800 1000.550 ;
        RECT 867.730 1000.000 868.010 1000.550 ;
        RECT 317.960 32.650 318.220 32.970 ;
        RECT 862.600 32.650 862.860 32.970 ;
        RECT 318.020 2.400 318.160 32.650 ;
        RECT 317.810 -4.800 318.370 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 335.870 15.540 336.190 15.600 ;
        RECT 897.070 15.540 897.390 15.600 ;
        RECT 335.870 15.400 897.390 15.540 ;
        RECT 335.870 15.340 336.190 15.400 ;
        RECT 897.070 15.340 897.390 15.400 ;
      LAYER via ;
        RECT 335.900 15.340 336.160 15.600 ;
        RECT 897.100 15.340 897.360 15.600 ;
      LAYER met2 ;
        RECT 899.470 1000.690 899.750 1004.000 ;
        RECT 897.160 1000.550 899.750 1000.690 ;
        RECT 897.160 15.630 897.300 1000.550 ;
        RECT 899.470 1000.000 899.750 1000.550 ;
        RECT 335.900 15.310 336.160 15.630 ;
        RECT 897.100 15.310 897.360 15.630 ;
        RECT 335.960 2.400 336.100 15.310 ;
        RECT 335.750 -4.800 336.310 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 358.410 993.380 358.730 993.440 ;
        RECT 931.570 993.380 931.890 993.440 ;
        RECT 358.410 993.240 931.890 993.380 ;
        RECT 358.410 993.180 358.730 993.240 ;
        RECT 931.570 993.180 931.890 993.240 ;
        RECT 353.350 16.900 353.670 16.960 ;
        RECT 358.410 16.900 358.730 16.960 ;
        RECT 353.350 16.760 358.730 16.900 ;
        RECT 353.350 16.700 353.670 16.760 ;
        RECT 358.410 16.700 358.730 16.760 ;
      LAYER via ;
        RECT 358.440 993.180 358.700 993.440 ;
        RECT 931.600 993.180 931.860 993.440 ;
        RECT 353.380 16.700 353.640 16.960 ;
        RECT 358.440 16.700 358.700 16.960 ;
      LAYER met2 ;
        RECT 931.670 1000.620 931.950 1004.000 ;
        RECT 931.660 1000.000 931.950 1000.620 ;
        RECT 931.660 993.470 931.800 1000.000 ;
        RECT 358.440 993.150 358.700 993.470 ;
        RECT 931.600 993.150 931.860 993.470 ;
        RECT 358.500 16.990 358.640 993.150 ;
        RECT 353.380 16.670 353.640 16.990 ;
        RECT 358.440 16.670 358.700 16.990 ;
        RECT 353.440 2.400 353.580 16.670 ;
        RECT 353.230 -4.800 353.790 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 371.290 16.220 371.610 16.280 ;
        RECT 959.170 16.220 959.490 16.280 ;
        RECT 371.290 16.080 959.490 16.220 ;
        RECT 371.290 16.020 371.610 16.080 ;
        RECT 959.170 16.020 959.490 16.080 ;
      LAYER via ;
        RECT 371.320 16.020 371.580 16.280 ;
        RECT 959.200 16.020 959.460 16.280 ;
      LAYER met2 ;
        RECT 963.410 1000.690 963.690 1004.000 ;
        RECT 959.260 1000.550 963.690 1000.690 ;
        RECT 959.260 16.310 959.400 1000.550 ;
        RECT 963.410 1000.000 963.690 1000.550 ;
        RECT 371.320 15.990 371.580 16.310 ;
        RECT 959.200 15.990 959.460 16.310 ;
        RECT 371.380 2.400 371.520 15.990 ;
        RECT 371.170 -4.800 371.730 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 392.910 992.700 393.230 992.760 ;
        RECT 995.050 992.700 995.370 992.760 ;
        RECT 392.910 992.560 995.370 992.700 ;
        RECT 392.910 992.500 393.230 992.560 ;
        RECT 995.050 992.500 995.370 992.560 ;
        RECT 389.230 16.900 389.550 16.960 ;
        RECT 392.910 16.900 393.230 16.960 ;
        RECT 389.230 16.760 393.230 16.900 ;
        RECT 389.230 16.700 389.550 16.760 ;
        RECT 392.910 16.700 393.230 16.760 ;
      LAYER via ;
        RECT 392.940 992.500 393.200 992.760 ;
        RECT 995.080 992.500 995.340 992.760 ;
        RECT 389.260 16.700 389.520 16.960 ;
        RECT 392.940 16.700 393.200 16.960 ;
      LAYER met2 ;
        RECT 995.150 1000.620 995.430 1004.000 ;
        RECT 995.140 1000.000 995.430 1000.620 ;
        RECT 995.140 992.790 995.280 1000.000 ;
        RECT 392.940 992.470 393.200 992.790 ;
        RECT 995.080 992.470 995.340 992.790 ;
        RECT 393.000 16.990 393.140 992.470 ;
        RECT 389.260 16.670 389.520 16.990 ;
        RECT 392.940 16.670 393.200 16.990 ;
        RECT 389.320 2.400 389.460 16.670 ;
        RECT 389.110 -4.800 389.670 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 407.170 16.900 407.490 16.960 ;
        RECT 1021.270 16.900 1021.590 16.960 ;
        RECT 407.170 16.760 1021.590 16.900 ;
        RECT 407.170 16.700 407.490 16.760 ;
        RECT 1021.270 16.700 1021.590 16.760 ;
      LAYER via ;
        RECT 407.200 16.700 407.460 16.960 ;
        RECT 1021.300 16.700 1021.560 16.960 ;
      LAYER met2 ;
        RECT 1027.350 1000.690 1027.630 1004.000 ;
        RECT 1021.360 1000.550 1027.630 1000.690 ;
        RECT 1021.360 16.990 1021.500 1000.550 ;
        RECT 1027.350 1000.000 1027.630 1000.550 ;
        RECT 407.200 16.670 407.460 16.990 ;
        RECT 1021.300 16.670 1021.560 16.990 ;
        RECT 407.260 2.400 407.400 16.670 ;
        RECT 407.050 -4.800 407.610 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 420.970 20.640 421.290 20.700 ;
        RECT 396.680 20.500 421.290 20.640 ;
        RECT 68.150 20.300 68.470 20.360 ;
        RECT 396.680 20.300 396.820 20.500 ;
        RECT 420.970 20.440 421.290 20.500 ;
        RECT 68.150 20.160 396.820 20.300 ;
        RECT 68.150 20.100 68.470 20.160 ;
      LAYER via ;
        RECT 68.180 20.100 68.440 20.360 ;
        RECT 421.000 20.440 421.260 20.700 ;
      LAYER met2 ;
        RECT 421.530 1000.690 421.810 1004.000 ;
        RECT 421.060 1000.550 421.810 1000.690 ;
        RECT 421.060 20.730 421.200 1000.550 ;
        RECT 421.530 1000.000 421.810 1000.550 ;
        RECT 421.000 20.410 421.260 20.730 ;
        RECT 68.180 20.070 68.440 20.390 ;
        RECT 68.240 2.400 68.380 20.070 ;
        RECT 68.030 -4.800 68.590 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 427.410 992.360 427.730 992.420 ;
        RECT 1058.990 992.360 1059.310 992.420 ;
        RECT 427.410 992.220 1059.310 992.360 ;
        RECT 427.410 992.160 427.730 992.220 ;
        RECT 1058.990 992.160 1059.310 992.220 ;
        RECT 424.650 20.640 424.970 20.700 ;
        RECT 427.410 20.640 427.730 20.700 ;
        RECT 424.650 20.500 427.730 20.640 ;
        RECT 424.650 20.440 424.970 20.500 ;
        RECT 427.410 20.440 427.730 20.500 ;
      LAYER via ;
        RECT 427.440 992.160 427.700 992.420 ;
        RECT 1059.020 992.160 1059.280 992.420 ;
        RECT 424.680 20.440 424.940 20.700 ;
        RECT 427.440 20.440 427.700 20.700 ;
      LAYER met2 ;
        RECT 1059.090 1000.620 1059.370 1004.000 ;
        RECT 1059.080 1000.000 1059.370 1000.620 ;
        RECT 1059.080 992.450 1059.220 1000.000 ;
        RECT 427.440 992.130 427.700 992.450 ;
        RECT 1059.020 992.130 1059.280 992.450 ;
        RECT 427.500 20.730 427.640 992.130 ;
        RECT 424.680 20.410 424.940 20.730 ;
        RECT 427.440 20.410 427.700 20.730 ;
        RECT 424.740 2.400 424.880 20.410 ;
        RECT 424.530 -4.800 425.090 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1090.270 20.300 1090.590 20.360 ;
        RECT 472.580 20.160 1090.590 20.300 ;
        RECT 442.590 19.960 442.910 20.020 ;
        RECT 472.580 19.960 472.720 20.160 ;
        RECT 1090.270 20.100 1090.590 20.160 ;
        RECT 442.590 19.820 472.720 19.960 ;
        RECT 442.590 19.760 442.910 19.820 ;
      LAYER via ;
        RECT 442.620 19.760 442.880 20.020 ;
        RECT 1090.300 20.100 1090.560 20.360 ;
      LAYER met2 ;
        RECT 1090.830 1000.690 1091.110 1004.000 ;
        RECT 1090.360 1000.550 1091.110 1000.690 ;
        RECT 1090.360 20.390 1090.500 1000.550 ;
        RECT 1090.830 1000.000 1091.110 1000.550 ;
        RECT 1090.300 20.070 1090.560 20.390 ;
        RECT 442.620 19.730 442.880 20.050 ;
        RECT 442.680 2.400 442.820 19.730 ;
        RECT 442.470 -4.800 443.030 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 461.910 991.680 462.230 991.740 ;
        RECT 1122.470 991.680 1122.790 991.740 ;
        RECT 461.910 991.540 1122.790 991.680 ;
        RECT 461.910 991.480 462.230 991.540 ;
        RECT 1122.470 991.480 1122.790 991.540 ;
        RECT 460.990 917.900 461.310 917.960 ;
        RECT 461.910 917.900 462.230 917.960 ;
        RECT 460.990 917.760 462.230 917.900 ;
        RECT 460.990 917.700 461.310 917.760 ;
        RECT 461.910 917.700 462.230 917.760 ;
        RECT 460.990 772.720 461.310 772.780 ;
        RECT 461.910 772.720 462.230 772.780 ;
        RECT 460.990 772.580 462.230 772.720 ;
        RECT 460.990 772.520 461.310 772.580 ;
        RECT 461.910 772.520 462.230 772.580 ;
        RECT 460.530 675.820 460.850 675.880 ;
        RECT 461.910 675.820 462.230 675.880 ;
        RECT 460.530 675.680 462.230 675.820 ;
        RECT 460.530 675.620 460.850 675.680 ;
        RECT 461.910 675.620 462.230 675.680 ;
        RECT 460.990 579.600 461.310 579.660 ;
        RECT 461.910 579.600 462.230 579.660 ;
        RECT 460.990 579.460 462.230 579.600 ;
        RECT 460.990 579.400 461.310 579.460 ;
        RECT 461.910 579.400 462.230 579.460 ;
        RECT 460.990 531.660 461.310 531.720 ;
        RECT 461.910 531.660 462.230 531.720 ;
        RECT 460.990 531.520 462.230 531.660 ;
        RECT 460.990 531.460 461.310 531.520 ;
        RECT 461.910 531.460 462.230 531.520 ;
        RECT 461.910 483.040 462.230 483.100 ;
        RECT 462.830 483.040 463.150 483.100 ;
        RECT 461.910 482.900 463.150 483.040 ;
        RECT 461.910 482.840 462.230 482.900 ;
        RECT 462.830 482.840 463.150 482.900 ;
        RECT 461.910 435.100 462.230 435.160 ;
        RECT 462.830 435.100 463.150 435.160 ;
        RECT 461.910 434.960 463.150 435.100 ;
        RECT 461.910 434.900 462.230 434.960 ;
        RECT 462.830 434.900 463.150 434.960 ;
        RECT 460.990 289.580 461.310 289.640 ;
        RECT 461.910 289.580 462.230 289.640 ;
        RECT 460.990 289.440 462.230 289.580 ;
        RECT 460.990 289.380 461.310 289.440 ;
        RECT 461.910 289.380 462.230 289.440 ;
        RECT 460.990 241.640 461.310 241.700 ;
        RECT 461.910 241.640 462.230 241.700 ;
        RECT 460.990 241.500 462.230 241.640 ;
        RECT 460.990 241.440 461.310 241.500 ;
        RECT 461.910 241.440 462.230 241.500 ;
        RECT 460.990 193.020 461.310 193.080 ;
        RECT 461.910 193.020 462.230 193.080 ;
        RECT 460.990 192.880 462.230 193.020 ;
        RECT 460.990 192.820 461.310 192.880 ;
        RECT 461.910 192.820 462.230 192.880 ;
        RECT 460.990 145.080 461.310 145.140 ;
        RECT 461.910 145.080 462.230 145.140 ;
        RECT 460.990 144.940 462.230 145.080 ;
        RECT 460.990 144.880 461.310 144.940 ;
        RECT 461.910 144.880 462.230 144.940 ;
        RECT 460.990 96.460 461.310 96.520 ;
        RECT 461.910 96.460 462.230 96.520 ;
        RECT 460.990 96.320 462.230 96.460 ;
        RECT 460.990 96.260 461.310 96.320 ;
        RECT 461.910 96.260 462.230 96.320 ;
        RECT 460.990 48.520 461.310 48.580 ;
        RECT 461.910 48.520 462.230 48.580 ;
        RECT 460.990 48.380 462.230 48.520 ;
        RECT 460.990 48.320 461.310 48.380 ;
        RECT 461.910 48.320 462.230 48.380 ;
        RECT 460.530 2.960 460.850 3.020 ;
        RECT 462.370 2.960 462.690 3.020 ;
        RECT 460.530 2.820 462.690 2.960 ;
        RECT 460.530 2.760 460.850 2.820 ;
        RECT 462.370 2.760 462.690 2.820 ;
      LAYER via ;
        RECT 461.940 991.480 462.200 991.740 ;
        RECT 1122.500 991.480 1122.760 991.740 ;
        RECT 461.020 917.700 461.280 917.960 ;
        RECT 461.940 917.700 462.200 917.960 ;
        RECT 461.020 772.520 461.280 772.780 ;
        RECT 461.940 772.520 462.200 772.780 ;
        RECT 460.560 675.620 460.820 675.880 ;
        RECT 461.940 675.620 462.200 675.880 ;
        RECT 461.020 579.400 461.280 579.660 ;
        RECT 461.940 579.400 462.200 579.660 ;
        RECT 461.020 531.460 461.280 531.720 ;
        RECT 461.940 531.460 462.200 531.720 ;
        RECT 461.940 482.840 462.200 483.100 ;
        RECT 462.860 482.840 463.120 483.100 ;
        RECT 461.940 434.900 462.200 435.160 ;
        RECT 462.860 434.900 463.120 435.160 ;
        RECT 461.020 289.380 461.280 289.640 ;
        RECT 461.940 289.380 462.200 289.640 ;
        RECT 461.020 241.440 461.280 241.700 ;
        RECT 461.940 241.440 462.200 241.700 ;
        RECT 461.020 192.820 461.280 193.080 ;
        RECT 461.940 192.820 462.200 193.080 ;
        RECT 461.020 144.880 461.280 145.140 ;
        RECT 461.940 144.880 462.200 145.140 ;
        RECT 461.020 96.260 461.280 96.520 ;
        RECT 461.940 96.260 462.200 96.520 ;
        RECT 461.020 48.320 461.280 48.580 ;
        RECT 461.940 48.320 462.200 48.580 ;
        RECT 460.560 2.760 460.820 3.020 ;
        RECT 462.400 2.760 462.660 3.020 ;
      LAYER met2 ;
        RECT 1122.570 1000.620 1122.850 1004.000 ;
        RECT 1122.560 1000.000 1122.850 1000.620 ;
        RECT 1122.560 991.770 1122.700 1000.000 ;
        RECT 461.940 991.450 462.200 991.770 ;
        RECT 1122.500 991.450 1122.760 991.770 ;
        RECT 462.000 966.125 462.140 991.450 ;
        RECT 461.010 965.755 461.290 966.125 ;
        RECT 461.930 965.755 462.210 966.125 ;
        RECT 461.080 917.990 461.220 965.755 ;
        RECT 461.020 917.670 461.280 917.990 ;
        RECT 461.940 917.670 462.200 917.990 ;
        RECT 462.000 869.565 462.140 917.670 ;
        RECT 461.010 869.195 461.290 869.565 ;
        RECT 461.930 869.195 462.210 869.565 ;
        RECT 461.080 821.285 461.220 869.195 ;
        RECT 461.010 820.915 461.290 821.285 ;
        RECT 461.930 820.915 462.210 821.285 ;
        RECT 462.000 772.810 462.140 820.915 ;
        RECT 461.020 772.490 461.280 772.810 ;
        RECT 461.940 772.490 462.200 772.810 ;
        RECT 461.080 724.725 461.220 772.490 ;
        RECT 461.010 724.355 461.290 724.725 ;
        RECT 461.930 724.355 462.210 724.725 ;
        RECT 462.000 675.910 462.140 724.355 ;
        RECT 460.560 675.590 460.820 675.910 ;
        RECT 461.940 675.590 462.200 675.910 ;
        RECT 460.620 628.165 460.760 675.590 ;
        RECT 460.550 627.795 460.830 628.165 ;
        RECT 461.930 627.795 462.210 628.165 ;
        RECT 462.000 579.690 462.140 627.795 ;
        RECT 461.020 579.370 461.280 579.690 ;
        RECT 461.940 579.370 462.200 579.690 ;
        RECT 461.080 531.750 461.220 579.370 ;
        RECT 461.020 531.430 461.280 531.750 ;
        RECT 461.940 531.430 462.200 531.750 ;
        RECT 462.000 483.130 462.140 531.430 ;
        RECT 461.940 482.810 462.200 483.130 ;
        RECT 462.860 482.810 463.120 483.130 ;
        RECT 462.920 435.190 463.060 482.810 ;
        RECT 461.940 434.870 462.200 435.190 ;
        RECT 462.860 434.870 463.120 435.190 ;
        RECT 462.000 289.670 462.140 434.870 ;
        RECT 461.020 289.350 461.280 289.670 ;
        RECT 461.940 289.350 462.200 289.670 ;
        RECT 461.080 241.730 461.220 289.350 ;
        RECT 461.020 241.410 461.280 241.730 ;
        RECT 461.940 241.410 462.200 241.730 ;
        RECT 462.000 193.110 462.140 241.410 ;
        RECT 461.020 192.790 461.280 193.110 ;
        RECT 461.940 192.790 462.200 193.110 ;
        RECT 461.080 145.170 461.220 192.790 ;
        RECT 461.020 144.850 461.280 145.170 ;
        RECT 461.940 144.850 462.200 145.170 ;
        RECT 462.000 96.550 462.140 144.850 ;
        RECT 461.020 96.230 461.280 96.550 ;
        RECT 461.940 96.230 462.200 96.550 ;
        RECT 461.080 48.610 461.220 96.230 ;
        RECT 461.020 48.290 461.280 48.610 ;
        RECT 461.940 48.290 462.200 48.610 ;
        RECT 462.000 16.050 462.140 48.290 ;
        RECT 462.000 15.910 462.600 16.050 ;
        RECT 462.460 3.050 462.600 15.910 ;
        RECT 460.560 2.730 460.820 3.050 ;
        RECT 462.400 2.730 462.660 3.050 ;
        RECT 460.620 2.400 460.760 2.730 ;
        RECT 460.410 -4.800 460.970 2.400 ;
      LAYER via2 ;
        RECT 461.010 965.800 461.290 966.080 ;
        RECT 461.930 965.800 462.210 966.080 ;
        RECT 461.010 869.240 461.290 869.520 ;
        RECT 461.930 869.240 462.210 869.520 ;
        RECT 461.010 820.960 461.290 821.240 ;
        RECT 461.930 820.960 462.210 821.240 ;
        RECT 461.010 724.400 461.290 724.680 ;
        RECT 461.930 724.400 462.210 724.680 ;
        RECT 460.550 627.840 460.830 628.120 ;
        RECT 461.930 627.840 462.210 628.120 ;
      LAYER met3 ;
        RECT 460.985 966.090 461.315 966.105 ;
        RECT 461.905 966.090 462.235 966.105 ;
        RECT 460.985 965.790 462.235 966.090 ;
        RECT 460.985 965.775 461.315 965.790 ;
        RECT 461.905 965.775 462.235 965.790 ;
        RECT 460.985 869.530 461.315 869.545 ;
        RECT 461.905 869.530 462.235 869.545 ;
        RECT 460.985 869.230 462.235 869.530 ;
        RECT 460.985 869.215 461.315 869.230 ;
        RECT 461.905 869.215 462.235 869.230 ;
        RECT 460.985 821.250 461.315 821.265 ;
        RECT 461.905 821.250 462.235 821.265 ;
        RECT 460.985 820.950 462.235 821.250 ;
        RECT 460.985 820.935 461.315 820.950 ;
        RECT 461.905 820.935 462.235 820.950 ;
        RECT 460.985 724.690 461.315 724.705 ;
        RECT 461.905 724.690 462.235 724.705 ;
        RECT 460.985 724.390 462.235 724.690 ;
        RECT 460.985 724.375 461.315 724.390 ;
        RECT 461.905 724.375 462.235 724.390 ;
        RECT 460.525 628.130 460.855 628.145 ;
        RECT 461.905 628.130 462.235 628.145 ;
        RECT 460.525 627.830 462.235 628.130 ;
        RECT 460.525 627.815 460.855 627.830 ;
        RECT 461.905 627.815 462.235 627.830 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 478.470 19.960 478.790 20.020 ;
        RECT 1152.370 19.960 1152.690 20.020 ;
        RECT 478.470 19.820 1152.690 19.960 ;
        RECT 478.470 19.760 478.790 19.820 ;
        RECT 1152.370 19.760 1152.690 19.820 ;
      LAYER via ;
        RECT 478.500 19.760 478.760 20.020 ;
        RECT 1152.400 19.760 1152.660 20.020 ;
      LAYER met2 ;
        RECT 1154.770 1000.690 1155.050 1004.000 ;
        RECT 1152.460 1000.550 1155.050 1000.690 ;
        RECT 1152.460 20.050 1152.600 1000.550 ;
        RECT 1154.770 1000.000 1155.050 1000.550 ;
        RECT 478.500 19.730 478.760 20.050 ;
        RECT 1152.400 19.730 1152.660 20.050 ;
        RECT 478.560 2.400 478.700 19.730 ;
        RECT 478.350 -4.800 478.910 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 495.950 991.000 496.270 991.060 ;
        RECT 1186.410 991.000 1186.730 991.060 ;
        RECT 495.950 990.860 1186.730 991.000 ;
        RECT 495.950 990.800 496.270 990.860 ;
        RECT 1186.410 990.800 1186.730 990.860 ;
      LAYER via ;
        RECT 495.980 990.800 496.240 991.060 ;
        RECT 1186.440 990.800 1186.700 991.060 ;
      LAYER met2 ;
        RECT 1186.510 1000.620 1186.790 1004.000 ;
        RECT 1186.500 1000.000 1186.790 1000.620 ;
        RECT 1186.500 991.090 1186.640 1000.000 ;
        RECT 495.980 990.770 496.240 991.090 ;
        RECT 1186.440 990.770 1186.700 991.090 ;
        RECT 496.040 3.130 496.180 990.770 ;
        RECT 496.040 2.990 496.640 3.130 ;
        RECT 496.500 2.400 496.640 2.990 ;
        RECT 496.290 -4.800 496.850 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 513.890 19.620 514.210 19.680 ;
        RECT 531.370 19.620 531.690 19.680 ;
        RECT 513.890 19.480 531.690 19.620 ;
        RECT 513.890 19.420 514.210 19.480 ;
        RECT 531.370 19.420 531.690 19.480 ;
        RECT 578.290 19.620 578.610 19.680 ;
        RECT 1214.470 19.620 1214.790 19.680 ;
        RECT 578.290 19.480 1214.790 19.620 ;
        RECT 578.290 19.420 578.610 19.480 ;
        RECT 1214.470 19.420 1214.790 19.480 ;
      LAYER via ;
        RECT 513.920 19.420 514.180 19.680 ;
        RECT 531.400 19.420 531.660 19.680 ;
        RECT 578.320 19.420 578.580 19.680 ;
        RECT 1214.500 19.420 1214.760 19.680 ;
      LAYER met2 ;
        RECT 1218.250 1000.690 1218.530 1004.000 ;
        RECT 1214.560 1000.550 1218.530 1000.690 ;
        RECT 531.390 19.875 531.670 20.245 ;
        RECT 578.310 19.875 578.590 20.245 ;
        RECT 531.460 19.710 531.600 19.875 ;
        RECT 578.380 19.710 578.520 19.875 ;
        RECT 1214.560 19.710 1214.700 1000.550 ;
        RECT 1218.250 1000.000 1218.530 1000.550 ;
        RECT 513.920 19.390 514.180 19.710 ;
        RECT 531.400 19.390 531.660 19.710 ;
        RECT 578.320 19.390 578.580 19.710 ;
        RECT 1214.500 19.390 1214.760 19.710 ;
        RECT 513.980 2.400 514.120 19.390 ;
        RECT 513.770 -4.800 514.330 2.400 ;
      LAYER via2 ;
        RECT 531.390 19.920 531.670 20.200 ;
        RECT 578.310 19.920 578.590 20.200 ;
      LAYER met3 ;
        RECT 531.365 20.210 531.695 20.225 ;
        RECT 578.285 20.210 578.615 20.225 ;
        RECT 531.365 19.910 578.615 20.210 ;
        RECT 531.365 19.895 531.695 19.910 ;
        RECT 578.285 19.895 578.615 19.910 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 537.810 990.320 538.130 990.380 ;
        RECT 1249.890 990.320 1250.210 990.380 ;
        RECT 537.810 990.180 1250.210 990.320 ;
        RECT 537.810 990.120 538.130 990.180 ;
        RECT 1249.890 990.120 1250.210 990.180 ;
        RECT 531.830 19.620 532.150 19.680 ;
        RECT 537.810 19.620 538.130 19.680 ;
        RECT 531.830 19.480 538.130 19.620 ;
        RECT 531.830 19.420 532.150 19.480 ;
        RECT 537.810 19.420 538.130 19.480 ;
      LAYER via ;
        RECT 537.840 990.120 538.100 990.380 ;
        RECT 1249.920 990.120 1250.180 990.380 ;
        RECT 531.860 19.420 532.120 19.680 ;
        RECT 537.840 19.420 538.100 19.680 ;
      LAYER met2 ;
        RECT 1249.990 1000.620 1250.270 1004.000 ;
        RECT 1249.980 1000.000 1250.270 1000.620 ;
        RECT 1249.980 990.410 1250.120 1000.000 ;
        RECT 537.840 990.090 538.100 990.410 ;
        RECT 1249.920 990.090 1250.180 990.410 ;
        RECT 537.900 19.710 538.040 990.090 ;
        RECT 531.860 19.390 532.120 19.710 ;
        RECT 537.840 19.390 538.100 19.710 ;
        RECT 531.920 2.400 532.060 19.390 ;
        RECT 531.710 -4.800 532.270 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 579.210 18.940 579.530 19.000 ;
        RECT 1276.570 18.940 1276.890 19.000 ;
        RECT 579.210 18.800 1276.890 18.940 ;
        RECT 579.210 18.740 579.530 18.800 ;
        RECT 1276.570 18.740 1276.890 18.800 ;
        RECT 549.770 9.760 550.090 9.820 ;
        RECT 579.210 9.760 579.530 9.820 ;
        RECT 549.770 9.620 579.530 9.760 ;
        RECT 549.770 9.560 550.090 9.620 ;
        RECT 579.210 9.560 579.530 9.620 ;
      LAYER via ;
        RECT 579.240 18.740 579.500 19.000 ;
        RECT 1276.600 18.740 1276.860 19.000 ;
        RECT 549.800 9.560 550.060 9.820 ;
        RECT 579.240 9.560 579.500 9.820 ;
      LAYER met2 ;
        RECT 1282.190 1000.690 1282.470 1004.000 ;
        RECT 1276.660 1000.550 1282.470 1000.690 ;
        RECT 1276.660 19.030 1276.800 1000.550 ;
        RECT 1282.190 1000.000 1282.470 1000.550 ;
        RECT 579.240 18.710 579.500 19.030 ;
        RECT 1276.600 18.710 1276.860 19.030 ;
        RECT 579.300 9.850 579.440 18.710 ;
        RECT 549.800 9.530 550.060 9.850 ;
        RECT 579.240 9.530 579.500 9.850 ;
        RECT 549.860 2.400 550.000 9.530 ;
        RECT 549.650 -4.800 550.210 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 567.710 18.600 568.030 18.660 ;
        RECT 1311.070 18.600 1311.390 18.660 ;
        RECT 567.710 18.460 1311.390 18.600 ;
        RECT 567.710 18.400 568.030 18.460 ;
        RECT 1311.070 18.400 1311.390 18.460 ;
      LAYER via ;
        RECT 567.740 18.400 568.000 18.660 ;
        RECT 1311.100 18.400 1311.360 18.660 ;
      LAYER met2 ;
        RECT 1313.930 1000.690 1314.210 1004.000 ;
        RECT 1311.160 1000.550 1314.210 1000.690 ;
        RECT 1311.160 18.690 1311.300 1000.550 ;
        RECT 1313.930 1000.000 1314.210 1000.550 ;
        RECT 567.740 18.370 568.000 18.690 ;
        RECT 1311.100 18.370 1311.360 18.690 ;
        RECT 567.800 2.400 567.940 18.370 ;
        RECT 567.590 -4.800 568.150 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1345.670 1000.620 1345.950 1004.000 ;
        RECT 1345.660 1000.000 1345.950 1000.620 ;
        RECT 1345.660 989.925 1345.800 1000.000 ;
        RECT 586.130 989.555 586.410 989.925 ;
        RECT 1345.590 989.555 1345.870 989.925 ;
        RECT 586.200 3.130 586.340 989.555 ;
        RECT 585.740 2.990 586.340 3.130 ;
        RECT 585.740 2.400 585.880 2.990 ;
        RECT 585.530 -4.800 586.090 2.400 ;
      LAYER via2 ;
        RECT 586.130 989.600 586.410 989.880 ;
        RECT 1345.590 989.600 1345.870 989.880 ;
      LAYER met3 ;
        RECT 586.105 989.890 586.435 989.905 ;
        RECT 1345.565 989.890 1345.895 989.905 ;
        RECT 586.105 989.590 1345.895 989.890 ;
        RECT 586.105 989.575 586.435 989.590 ;
        RECT 1345.565 989.575 1345.895 989.590 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 462.370 20.300 462.690 20.360 ;
        RECT 412.780 20.160 462.690 20.300 ;
        RECT 91.610 19.960 91.930 20.020 ;
        RECT 412.780 19.960 412.920 20.160 ;
        RECT 462.370 20.100 462.690 20.160 ;
        RECT 91.610 19.820 412.920 19.960 ;
        RECT 91.610 19.760 91.930 19.820 ;
      LAYER via ;
        RECT 91.640 19.760 91.900 20.020 ;
        RECT 462.400 20.100 462.660 20.360 ;
      LAYER met2 ;
        RECT 464.310 1000.690 464.590 1004.000 ;
        RECT 462.460 1000.550 464.590 1000.690 ;
        RECT 462.460 20.390 462.600 1000.550 ;
        RECT 464.310 1000.000 464.590 1000.550 ;
        RECT 462.400 20.070 462.660 20.390 ;
        RECT 91.640 19.730 91.900 20.050 ;
        RECT 91.700 2.400 91.840 19.730 ;
        RECT 91.490 -4.800 92.050 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 603.130 17.920 603.450 17.980 ;
        RECT 1373.170 17.920 1373.490 17.980 ;
        RECT 603.130 17.780 1373.490 17.920 ;
        RECT 603.130 17.720 603.450 17.780 ;
        RECT 1373.170 17.720 1373.490 17.780 ;
      LAYER via ;
        RECT 603.160 17.720 603.420 17.980 ;
        RECT 1373.200 17.720 1373.460 17.980 ;
      LAYER met2 ;
        RECT 1377.410 1000.690 1377.690 1004.000 ;
        RECT 1373.260 1000.550 1377.690 1000.690 ;
        RECT 1373.260 18.010 1373.400 1000.550 ;
        RECT 1377.410 1000.000 1377.690 1000.550 ;
        RECT 603.160 17.690 603.420 18.010 ;
        RECT 1373.200 17.690 1373.460 18.010 ;
        RECT 603.220 2.400 603.360 17.690 ;
        RECT 603.010 -4.800 603.570 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 621.070 17.240 621.390 17.300 ;
        RECT 1407.670 17.240 1407.990 17.300 ;
        RECT 621.070 17.100 1407.990 17.240 ;
        RECT 621.070 17.040 621.390 17.100 ;
        RECT 1407.670 17.040 1407.990 17.100 ;
      LAYER via ;
        RECT 621.100 17.040 621.360 17.300 ;
        RECT 1407.700 17.040 1407.960 17.300 ;
      LAYER met2 ;
        RECT 1409.610 1000.690 1409.890 1004.000 ;
        RECT 1407.760 1000.550 1409.890 1000.690 ;
        RECT 1407.760 17.330 1407.900 1000.550 ;
        RECT 1409.610 1000.000 1409.890 1000.550 ;
        RECT 621.100 17.010 621.360 17.330 ;
        RECT 1407.700 17.010 1407.960 17.330 ;
        RECT 621.160 2.400 621.300 17.010 ;
        RECT 620.950 -4.800 621.510 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 503.770 19.280 504.090 19.340 ;
        RECT 138.160 19.140 504.090 19.280 ;
        RECT 115.530 18.940 115.850 19.000 ;
        RECT 138.160 18.940 138.300 19.140 ;
        RECT 503.770 19.080 504.090 19.140 ;
        RECT 115.530 18.800 138.300 18.940 ;
        RECT 115.530 18.740 115.850 18.800 ;
      LAYER via ;
        RECT 115.560 18.740 115.820 19.000 ;
        RECT 503.800 19.080 504.060 19.340 ;
      LAYER met2 ;
        RECT 506.630 1000.690 506.910 1004.000 ;
        RECT 503.860 1000.550 506.910 1000.690 ;
        RECT 503.860 19.370 504.000 1000.550 ;
        RECT 506.630 1000.000 506.910 1000.550 ;
        RECT 503.800 19.050 504.060 19.370 ;
        RECT 115.560 18.710 115.820 19.030 ;
        RECT 115.620 2.400 115.760 18.710 ;
        RECT 115.410 -4.800 115.970 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 139.450 18.940 139.770 19.000 ;
        RECT 545.170 18.940 545.490 19.000 ;
        RECT 139.450 18.800 545.490 18.940 ;
        RECT 139.450 18.740 139.770 18.800 ;
        RECT 545.170 18.740 545.490 18.800 ;
      LAYER via ;
        RECT 139.480 18.740 139.740 19.000 ;
        RECT 545.200 18.740 545.460 19.000 ;
      LAYER met2 ;
        RECT 549.410 1000.690 549.690 1004.000 ;
        RECT 545.260 1000.550 549.690 1000.690 ;
        RECT 545.260 19.030 545.400 1000.550 ;
        RECT 549.410 1000.000 549.690 1000.550 ;
        RECT 139.480 18.710 139.740 19.030 ;
        RECT 545.200 18.710 545.460 19.030 ;
        RECT 139.540 2.400 139.680 18.710 ;
        RECT 139.330 -4.800 139.890 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 157.390 18.260 157.710 18.320 ;
        RECT 157.390 18.120 555.520 18.260 ;
        RECT 157.390 18.060 157.710 18.120 ;
        RECT 555.380 17.920 555.520 18.120 ;
        RECT 579.670 17.920 579.990 17.980 ;
        RECT 555.380 17.780 579.990 17.920 ;
        RECT 579.670 17.720 579.990 17.780 ;
      LAYER via ;
        RECT 157.420 18.060 157.680 18.320 ;
        RECT 579.700 17.720 579.960 17.980 ;
      LAYER met2 ;
        RECT 581.150 1000.690 581.430 1004.000 ;
        RECT 579.760 1000.550 581.430 1000.690 ;
        RECT 157.420 18.030 157.680 18.350 ;
        RECT 157.480 2.400 157.620 18.030 ;
        RECT 579.760 18.010 579.900 1000.550 ;
        RECT 581.150 1000.000 581.430 1000.550 ;
        RECT 579.700 17.690 579.960 18.010 ;
        RECT 157.270 -4.800 157.830 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 174.870 17.580 175.190 17.640 ;
        RECT 607.270 17.580 607.590 17.640 ;
        RECT 174.870 17.440 607.590 17.580 ;
        RECT 174.870 17.380 175.190 17.440 ;
        RECT 607.270 17.380 607.590 17.440 ;
      LAYER via ;
        RECT 174.900 17.380 175.160 17.640 ;
        RECT 607.300 17.380 607.560 17.640 ;
      LAYER met2 ;
        RECT 612.890 1000.690 613.170 1004.000 ;
        RECT 607.360 1000.550 613.170 1000.690 ;
        RECT 607.360 17.670 607.500 1000.550 ;
        RECT 612.890 1000.000 613.170 1000.550 ;
        RECT 174.900 17.350 175.160 17.670 ;
        RECT 607.300 17.350 607.560 17.670 ;
        RECT 174.960 2.400 175.100 17.350 ;
        RECT 174.750 -4.800 175.310 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 192.810 14.180 193.130 14.240 ;
        RECT 642.230 14.180 642.550 14.240 ;
        RECT 192.810 14.040 642.550 14.180 ;
        RECT 192.810 13.980 193.130 14.040 ;
        RECT 642.230 13.980 642.550 14.040 ;
      LAYER via ;
        RECT 192.840 13.980 193.100 14.240 ;
        RECT 642.260 13.980 642.520 14.240 ;
      LAYER met2 ;
        RECT 644.630 1000.690 644.910 1004.000 ;
        RECT 642.320 1000.550 644.910 1000.690 ;
        RECT 642.320 14.270 642.460 1000.550 ;
        RECT 644.630 1000.000 644.910 1000.550 ;
        RECT 192.840 13.950 193.100 14.270 ;
        RECT 642.260 13.950 642.520 14.270 ;
        RECT 192.900 2.400 193.040 13.950 ;
        RECT 192.690 -4.800 193.250 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 213.510 987.600 213.830 987.660 ;
        RECT 676.730 987.600 677.050 987.660 ;
        RECT 213.510 987.460 677.050 987.600 ;
        RECT 213.510 987.400 213.830 987.460 ;
        RECT 676.730 987.400 677.050 987.460 ;
        RECT 210.750 17.240 211.070 17.300 ;
        RECT 213.510 17.240 213.830 17.300 ;
        RECT 210.750 17.100 213.830 17.240 ;
        RECT 210.750 17.040 211.070 17.100 ;
        RECT 213.510 17.040 213.830 17.100 ;
      LAYER via ;
        RECT 213.540 987.400 213.800 987.660 ;
        RECT 676.760 987.400 677.020 987.660 ;
        RECT 210.780 17.040 211.040 17.300 ;
        RECT 213.540 17.040 213.800 17.300 ;
      LAYER met2 ;
        RECT 676.830 1000.620 677.110 1004.000 ;
        RECT 676.820 1000.000 677.110 1000.620 ;
        RECT 676.820 987.690 676.960 1000.000 ;
        RECT 213.540 987.370 213.800 987.690 ;
        RECT 676.760 987.370 677.020 987.690 ;
        RECT 213.600 17.330 213.740 987.370 ;
        RECT 210.780 17.010 211.040 17.330 ;
        RECT 213.540 17.010 213.800 17.330 ;
        RECT 210.840 2.400 210.980 17.010 ;
        RECT 210.630 -4.800 211.190 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 275.610 14.860 275.930 14.920 ;
        RECT 703.870 14.860 704.190 14.920 ;
        RECT 275.610 14.720 704.190 14.860 ;
        RECT 275.610 14.660 275.930 14.720 ;
        RECT 703.870 14.660 704.190 14.720 ;
        RECT 228.690 13.840 229.010 13.900 ;
        RECT 275.610 13.840 275.930 13.900 ;
        RECT 228.690 13.700 275.930 13.840 ;
        RECT 228.690 13.640 229.010 13.700 ;
        RECT 275.610 13.640 275.930 13.700 ;
      LAYER via ;
        RECT 275.640 14.660 275.900 14.920 ;
        RECT 703.900 14.660 704.160 14.920 ;
        RECT 228.720 13.640 228.980 13.900 ;
        RECT 275.640 13.640 275.900 13.900 ;
      LAYER met2 ;
        RECT 708.570 1000.690 708.850 1004.000 ;
        RECT 703.960 1000.550 708.850 1000.690 ;
        RECT 703.960 14.950 704.100 1000.550 ;
        RECT 708.570 1000.000 708.850 1000.550 ;
        RECT 275.640 14.630 275.900 14.950 ;
        RECT 703.900 14.630 704.160 14.950 ;
        RECT 275.700 13.930 275.840 14.630 ;
        RECT 228.720 13.610 228.980 13.930 ;
        RECT 275.640 13.610 275.900 13.930 ;
        RECT 228.780 2.400 228.920 13.610 ;
        RECT 228.570 -4.800 229.130 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 54.810 992.020 55.130 992.080 ;
        RECT 389.690 992.020 390.010 992.080 ;
        RECT 54.810 991.880 390.010 992.020 ;
        RECT 54.810 991.820 55.130 991.880 ;
        RECT 389.690 991.820 390.010 991.880 ;
        RECT 50.210 17.580 50.530 17.640 ;
        RECT 54.810 17.580 55.130 17.640 ;
        RECT 50.210 17.440 55.130 17.580 ;
        RECT 50.210 17.380 50.530 17.440 ;
        RECT 54.810 17.380 55.130 17.440 ;
      LAYER via ;
        RECT 54.840 991.820 55.100 992.080 ;
        RECT 389.720 991.820 389.980 992.080 ;
        RECT 50.240 17.380 50.500 17.640 ;
        RECT 54.840 17.380 55.100 17.640 ;
      LAYER met2 ;
        RECT 389.790 1000.620 390.070 1004.000 ;
        RECT 389.780 1000.000 390.070 1000.620 ;
        RECT 389.780 992.110 389.920 1000.000 ;
        RECT 54.840 991.790 55.100 992.110 ;
        RECT 389.720 991.790 389.980 992.110 ;
        RECT 54.900 17.670 55.040 991.790 ;
        RECT 50.240 17.350 50.500 17.670 ;
        RECT 54.840 17.350 55.100 17.670 ;
        RECT 50.300 2.400 50.440 17.350 ;
        RECT 50.090 -4.800 50.650 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 254.910 988.280 255.230 988.340 ;
        RECT 750.790 988.280 751.110 988.340 ;
        RECT 254.910 988.140 751.110 988.280 ;
        RECT 254.910 988.080 255.230 988.140 ;
        RECT 750.790 988.080 751.110 988.140 ;
        RECT 252.610 14.860 252.930 14.920 ;
        RECT 254.910 14.860 255.230 14.920 ;
        RECT 252.610 14.720 255.230 14.860 ;
        RECT 252.610 14.660 252.930 14.720 ;
        RECT 254.910 14.660 255.230 14.720 ;
      LAYER via ;
        RECT 254.940 988.080 255.200 988.340 ;
        RECT 750.820 988.080 751.080 988.340 ;
        RECT 252.640 14.660 252.900 14.920 ;
        RECT 254.940 14.660 255.200 14.920 ;
      LAYER met2 ;
        RECT 750.890 1000.620 751.170 1004.000 ;
        RECT 750.880 1000.000 751.170 1000.620 ;
        RECT 750.880 988.370 751.020 1000.000 ;
        RECT 254.940 988.050 255.200 988.370 ;
        RECT 750.820 988.050 751.080 988.370 ;
        RECT 255.000 14.950 255.140 988.050 ;
        RECT 252.640 14.630 252.900 14.950 ;
        RECT 254.940 14.630 255.200 14.950 ;
        RECT 252.700 2.400 252.840 14.630 ;
        RECT 252.490 -4.800 253.050 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 275.610 988.620 275.930 988.680 ;
        RECT 782.530 988.620 782.850 988.680 ;
        RECT 275.610 988.480 782.850 988.620 ;
        RECT 275.610 988.420 275.930 988.480 ;
        RECT 782.530 988.420 782.850 988.480 ;
        RECT 270.090 14.860 270.410 14.920 ;
        RECT 275.150 14.860 275.470 14.920 ;
        RECT 270.090 14.720 275.470 14.860 ;
        RECT 270.090 14.660 270.410 14.720 ;
        RECT 275.150 14.660 275.470 14.720 ;
      LAYER via ;
        RECT 275.640 988.420 275.900 988.680 ;
        RECT 782.560 988.420 782.820 988.680 ;
        RECT 270.120 14.660 270.380 14.920 ;
        RECT 275.180 14.660 275.440 14.920 ;
      LAYER met2 ;
        RECT 782.630 1000.620 782.910 1004.000 ;
        RECT 782.620 1000.000 782.910 1000.620 ;
        RECT 782.620 988.710 782.760 1000.000 ;
        RECT 275.640 988.390 275.900 988.710 ;
        RECT 782.560 988.390 782.820 988.710 ;
        RECT 275.700 15.370 275.840 988.390 ;
        RECT 275.240 15.230 275.840 15.370 ;
        RECT 275.240 14.950 275.380 15.230 ;
        RECT 270.120 14.630 270.380 14.950 ;
        RECT 275.180 14.630 275.440 14.950 ;
        RECT 270.180 2.400 270.320 14.630 ;
        RECT 269.970 -4.800 270.530 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 289.410 988.960 289.730 989.020 ;
        RECT 814.730 988.960 815.050 989.020 ;
        RECT 289.410 988.820 815.050 988.960 ;
        RECT 289.410 988.760 289.730 988.820 ;
        RECT 814.730 988.760 815.050 988.820 ;
      LAYER via ;
        RECT 289.440 988.760 289.700 989.020 ;
        RECT 814.760 988.760 815.020 989.020 ;
      LAYER met2 ;
        RECT 814.830 1000.620 815.110 1004.000 ;
        RECT 814.820 1000.000 815.110 1000.620 ;
        RECT 814.820 989.050 814.960 1000.000 ;
        RECT 289.440 988.730 289.700 989.050 ;
        RECT 814.760 988.730 815.020 989.050 ;
        RECT 289.500 16.730 289.640 988.730 ;
        RECT 288.120 16.590 289.640 16.730 ;
        RECT 288.120 2.400 288.260 16.590 ;
        RECT 287.910 -4.800 288.470 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 305.970 15.200 306.290 15.260 ;
        RECT 841.870 15.200 842.190 15.260 ;
        RECT 305.970 15.060 842.190 15.200 ;
        RECT 305.970 15.000 306.290 15.060 ;
        RECT 841.870 15.000 842.190 15.060 ;
      LAYER via ;
        RECT 306.000 15.000 306.260 15.260 ;
        RECT 841.900 15.000 842.160 15.260 ;
      LAYER met2 ;
        RECT 846.570 1000.690 846.850 1004.000 ;
        RECT 841.960 1000.550 846.850 1000.690 ;
        RECT 841.960 15.290 842.100 1000.550 ;
        RECT 846.570 1000.000 846.850 1000.550 ;
        RECT 306.000 14.970 306.260 15.290 ;
        RECT 841.900 14.970 842.160 15.290 ;
        RECT 306.060 2.400 306.200 14.970 ;
        RECT 305.850 -4.800 306.410 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 323.910 989.300 324.230 989.360 ;
        RECT 878.210 989.300 878.530 989.360 ;
        RECT 323.910 989.160 878.530 989.300 ;
        RECT 323.910 989.100 324.230 989.160 ;
        RECT 878.210 989.100 878.530 989.160 ;
      LAYER via ;
        RECT 323.940 989.100 324.200 989.360 ;
        RECT 878.240 989.100 878.500 989.360 ;
      LAYER met2 ;
        RECT 878.310 1000.620 878.590 1004.000 ;
        RECT 878.300 1000.000 878.590 1000.620 ;
        RECT 878.300 989.390 878.440 1000.000 ;
        RECT 323.940 989.070 324.200 989.390 ;
        RECT 878.240 989.070 878.500 989.390 ;
        RECT 324.000 2.400 324.140 989.070 ;
        RECT 323.790 -4.800 324.350 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 341.390 15.880 341.710 15.940 ;
        RECT 903.970 15.880 904.290 15.940 ;
        RECT 341.390 15.740 904.290 15.880 ;
        RECT 341.390 15.680 341.710 15.740 ;
        RECT 903.970 15.680 904.290 15.740 ;
      LAYER via ;
        RECT 341.420 15.680 341.680 15.940 ;
        RECT 904.000 15.680 904.260 15.940 ;
      LAYER met2 ;
        RECT 910.510 1000.690 910.790 1004.000 ;
        RECT 904.060 1000.550 910.790 1000.690 ;
        RECT 904.060 15.970 904.200 1000.550 ;
        RECT 910.510 1000.000 910.790 1000.550 ;
        RECT 341.420 15.650 341.680 15.970 ;
        RECT 904.000 15.650 904.260 15.970 ;
        RECT 341.480 2.400 341.620 15.650 ;
        RECT 341.270 -4.800 341.830 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 364.850 989.640 365.170 989.700 ;
        RECT 942.150 989.640 942.470 989.700 ;
        RECT 364.850 989.500 942.470 989.640 ;
        RECT 364.850 989.440 365.170 989.500 ;
        RECT 942.150 989.440 942.470 989.500 ;
        RECT 359.330 16.900 359.650 16.960 ;
        RECT 364.850 16.900 365.170 16.960 ;
        RECT 359.330 16.760 365.170 16.900 ;
        RECT 359.330 16.700 359.650 16.760 ;
        RECT 364.850 16.700 365.170 16.760 ;
      LAYER via ;
        RECT 364.880 989.440 365.140 989.700 ;
        RECT 942.180 989.440 942.440 989.700 ;
        RECT 359.360 16.700 359.620 16.960 ;
        RECT 364.880 16.700 365.140 16.960 ;
      LAYER met2 ;
        RECT 942.250 1000.620 942.530 1004.000 ;
        RECT 942.240 1000.000 942.530 1000.620 ;
        RECT 942.240 989.730 942.380 1000.000 ;
        RECT 364.880 989.410 365.140 989.730 ;
        RECT 942.180 989.410 942.440 989.730 ;
        RECT 364.940 16.990 365.080 989.410 ;
        RECT 359.360 16.670 359.620 16.990 ;
        RECT 364.880 16.670 365.140 16.990 ;
        RECT 359.420 2.400 359.560 16.670 ;
        RECT 359.210 -4.800 359.770 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 377.270 16.560 377.590 16.620 ;
        RECT 972.970 16.560 973.290 16.620 ;
        RECT 377.270 16.420 973.290 16.560 ;
        RECT 377.270 16.360 377.590 16.420 ;
        RECT 972.970 16.360 973.290 16.420 ;
      LAYER via ;
        RECT 377.300 16.360 377.560 16.620 ;
        RECT 973.000 16.360 973.260 16.620 ;
      LAYER met2 ;
        RECT 973.990 1000.690 974.270 1004.000 ;
        RECT 973.060 1000.550 974.270 1000.690 ;
        RECT 973.060 16.650 973.200 1000.550 ;
        RECT 973.990 1000.000 974.270 1000.550 ;
        RECT 377.300 16.330 377.560 16.650 ;
        RECT 973.000 16.330 973.260 16.650 ;
        RECT 377.360 2.400 377.500 16.330 ;
        RECT 377.150 -4.800 377.710 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 399.810 993.040 400.130 993.100 ;
        RECT 1005.630 993.040 1005.950 993.100 ;
        RECT 399.810 992.900 1005.950 993.040 ;
        RECT 399.810 992.840 400.130 992.900 ;
        RECT 1005.630 992.840 1005.950 992.900 ;
        RECT 395.210 16.900 395.530 16.960 ;
        RECT 399.810 16.900 400.130 16.960 ;
        RECT 395.210 16.760 400.130 16.900 ;
        RECT 395.210 16.700 395.530 16.760 ;
        RECT 399.810 16.700 400.130 16.760 ;
      LAYER via ;
        RECT 399.840 992.840 400.100 993.100 ;
        RECT 1005.660 992.840 1005.920 993.100 ;
        RECT 395.240 16.700 395.500 16.960 ;
        RECT 399.840 16.700 400.100 16.960 ;
      LAYER met2 ;
        RECT 1005.730 1000.620 1006.010 1004.000 ;
        RECT 1005.720 1000.000 1006.010 1000.620 ;
        RECT 1005.720 993.130 1005.860 1000.000 ;
        RECT 399.840 992.810 400.100 993.130 ;
        RECT 1005.660 992.810 1005.920 993.130 ;
        RECT 399.900 16.990 400.040 992.810 ;
        RECT 395.240 16.670 395.500 16.990 ;
        RECT 399.840 16.670 400.100 16.990 ;
        RECT 395.300 2.400 395.440 16.670 ;
        RECT 395.090 -4.800 395.650 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 434.770 20.640 435.090 20.700 ;
        RECT 1035.070 20.640 1035.390 20.700 ;
        RECT 434.770 20.500 1035.390 20.640 ;
        RECT 434.770 20.440 435.090 20.500 ;
        RECT 1035.070 20.440 1035.390 20.500 ;
        RECT 413.150 19.960 413.470 20.020 ;
        RECT 434.770 19.960 435.090 20.020 ;
        RECT 413.150 19.820 435.090 19.960 ;
        RECT 413.150 19.760 413.470 19.820 ;
        RECT 434.770 19.760 435.090 19.820 ;
      LAYER via ;
        RECT 434.800 20.440 435.060 20.700 ;
        RECT 1035.100 20.440 1035.360 20.700 ;
        RECT 413.180 19.760 413.440 20.020 ;
        RECT 434.800 19.760 435.060 20.020 ;
      LAYER met2 ;
        RECT 1037.930 1000.690 1038.210 1004.000 ;
        RECT 1035.160 1000.550 1038.210 1000.690 ;
        RECT 1035.160 20.730 1035.300 1000.550 ;
        RECT 1037.930 1000.000 1038.210 1000.550 ;
        RECT 434.800 20.410 435.060 20.730 ;
        RECT 1035.100 20.410 1035.360 20.730 ;
        RECT 434.860 20.050 435.000 20.410 ;
        RECT 413.180 19.730 413.440 20.050 ;
        RECT 434.800 19.730 435.060 20.050 ;
        RECT 413.240 2.400 413.380 19.730 ;
        RECT 413.030 -4.800 413.590 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 75.510 991.340 75.830 991.400 ;
        RECT 432.470 991.340 432.790 991.400 ;
        RECT 75.510 991.200 432.790 991.340 ;
        RECT 75.510 991.140 75.830 991.200 ;
        RECT 432.470 991.140 432.790 991.200 ;
      LAYER via ;
        RECT 75.540 991.140 75.800 991.400 ;
        RECT 432.500 991.140 432.760 991.400 ;
      LAYER met2 ;
        RECT 432.570 1000.620 432.850 1004.000 ;
        RECT 432.560 1000.000 432.850 1000.620 ;
        RECT 432.560 991.430 432.700 1000.000 ;
        RECT 75.540 991.110 75.800 991.430 ;
        RECT 432.500 991.110 432.760 991.430 ;
        RECT 75.600 17.410 75.740 991.110 ;
        RECT 74.220 17.270 75.740 17.410 ;
        RECT 74.220 2.400 74.360 17.270 ;
        RECT 74.010 -4.800 74.570 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 434.310 992.020 434.630 992.080 ;
        RECT 1069.570 992.020 1069.890 992.080 ;
        RECT 434.310 991.880 1069.890 992.020 ;
        RECT 434.310 991.820 434.630 991.880 ;
        RECT 1069.570 991.820 1069.890 991.880 ;
        RECT 430.630 20.640 430.950 20.700 ;
        RECT 434.310 20.640 434.630 20.700 ;
        RECT 430.630 20.500 434.630 20.640 ;
        RECT 430.630 20.440 430.950 20.500 ;
        RECT 434.310 20.440 434.630 20.500 ;
      LAYER via ;
        RECT 434.340 991.820 434.600 992.080 ;
        RECT 1069.600 991.820 1069.860 992.080 ;
        RECT 430.660 20.440 430.920 20.700 ;
        RECT 434.340 20.440 434.600 20.700 ;
      LAYER met2 ;
        RECT 1069.670 1000.620 1069.950 1004.000 ;
        RECT 1069.660 1000.000 1069.950 1000.620 ;
        RECT 1069.660 992.110 1069.800 1000.000 ;
        RECT 434.340 991.790 434.600 992.110 ;
        RECT 1069.600 991.790 1069.860 992.110 ;
        RECT 434.400 20.730 434.540 991.790 ;
        RECT 430.660 20.410 430.920 20.730 ;
        RECT 434.340 20.410 434.600 20.730 ;
        RECT 430.720 2.400 430.860 20.410 ;
        RECT 430.510 -4.800 431.070 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1101.410 1000.690 1101.690 1004.000 ;
        RECT 1097.260 1000.550 1101.690 1000.690 ;
        RECT 1097.260 18.885 1097.400 1000.550 ;
        RECT 1101.410 1000.000 1101.690 1000.550 ;
        RECT 448.590 18.515 448.870 18.885 ;
        RECT 1097.190 18.515 1097.470 18.885 ;
        RECT 448.660 2.400 448.800 18.515 ;
        RECT 448.450 -4.800 449.010 2.400 ;
      LAYER via2 ;
        RECT 448.590 18.560 448.870 18.840 ;
        RECT 1097.190 18.560 1097.470 18.840 ;
      LAYER met3 ;
        RECT 448.565 18.850 448.895 18.865 ;
        RECT 1097.165 18.850 1097.495 18.865 ;
        RECT 448.565 18.550 1097.495 18.850 ;
        RECT 448.565 18.535 448.895 18.550 ;
        RECT 1097.165 18.535 1097.495 18.550 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 468.810 991.340 469.130 991.400 ;
        RECT 1133.050 991.340 1133.370 991.400 ;
        RECT 468.810 991.200 1133.370 991.340 ;
        RECT 468.810 991.140 469.130 991.200 ;
        RECT 1133.050 991.140 1133.370 991.200 ;
        RECT 466.510 20.300 466.830 20.360 ;
        RECT 468.810 20.300 469.130 20.360 ;
        RECT 466.510 20.160 469.130 20.300 ;
        RECT 466.510 20.100 466.830 20.160 ;
        RECT 468.810 20.100 469.130 20.160 ;
      LAYER via ;
        RECT 468.840 991.140 469.100 991.400 ;
        RECT 1133.080 991.140 1133.340 991.400 ;
        RECT 466.540 20.100 466.800 20.360 ;
        RECT 468.840 20.100 469.100 20.360 ;
      LAYER met2 ;
        RECT 1133.150 1000.620 1133.430 1004.000 ;
        RECT 1133.140 1000.000 1133.430 1000.620 ;
        RECT 1133.140 991.430 1133.280 1000.000 ;
        RECT 468.840 991.110 469.100 991.430 ;
        RECT 1133.080 991.110 1133.340 991.430 ;
        RECT 468.900 20.390 469.040 991.110 ;
        RECT 466.540 20.070 466.800 20.390 ;
        RECT 468.840 20.070 469.100 20.390 ;
        RECT 466.600 2.400 466.740 20.070 ;
        RECT 466.390 -4.800 466.950 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1165.350 1000.690 1165.630 1004.000 ;
        RECT 1159.360 1000.550 1165.630 1000.690 ;
        RECT 1159.360 18.205 1159.500 1000.550 ;
        RECT 1165.350 1000.000 1165.630 1000.550 ;
        RECT 484.470 17.835 484.750 18.205 ;
        RECT 1159.290 17.835 1159.570 18.205 ;
        RECT 484.540 2.400 484.680 17.835 ;
        RECT 484.330 -4.800 484.890 2.400 ;
      LAYER via2 ;
        RECT 484.470 17.880 484.750 18.160 ;
        RECT 1159.290 17.880 1159.570 18.160 ;
      LAYER met3 ;
        RECT 484.445 18.170 484.775 18.185 ;
        RECT 1159.265 18.170 1159.595 18.185 ;
        RECT 484.445 17.870 1159.595 18.170 ;
        RECT 484.445 17.855 484.775 17.870 ;
        RECT 1159.265 17.855 1159.595 17.870 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 503.310 990.660 503.630 990.720 ;
        RECT 1196.990 990.660 1197.310 990.720 ;
        RECT 503.310 990.520 1197.310 990.660 ;
        RECT 503.310 990.460 503.630 990.520 ;
        RECT 1196.990 990.460 1197.310 990.520 ;
      LAYER via ;
        RECT 503.340 990.460 503.600 990.720 ;
        RECT 1197.020 990.460 1197.280 990.720 ;
      LAYER met2 ;
        RECT 1197.090 1000.620 1197.370 1004.000 ;
        RECT 1197.080 1000.000 1197.370 1000.620 ;
        RECT 1197.080 990.750 1197.220 1000.000 ;
        RECT 503.340 990.430 503.600 990.750 ;
        RECT 1197.020 990.430 1197.280 990.750 ;
        RECT 503.400 3.130 503.540 990.430 ;
        RECT 502.480 2.990 503.540 3.130 ;
        RECT 502.480 2.400 502.620 2.990 ;
        RECT 502.270 -4.800 502.830 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 519.870 19.280 520.190 19.340 ;
        RECT 1228.270 19.280 1228.590 19.340 ;
        RECT 519.870 19.140 573.920 19.280 ;
        RECT 519.870 19.080 520.190 19.140 ;
        RECT 573.780 18.940 573.920 19.140 ;
        RECT 578.380 19.140 1228.590 19.280 ;
        RECT 578.380 18.940 578.520 19.140 ;
        RECT 1228.270 19.080 1228.590 19.140 ;
        RECT 573.780 18.800 578.520 18.940 ;
      LAYER via ;
        RECT 519.900 19.080 520.160 19.340 ;
        RECT 1228.300 19.080 1228.560 19.340 ;
      LAYER met2 ;
        RECT 1228.830 1000.690 1229.110 1004.000 ;
        RECT 1228.360 1000.550 1229.110 1000.690 ;
        RECT 1228.360 19.370 1228.500 1000.550 ;
        RECT 1228.830 1000.000 1229.110 1000.550 ;
        RECT 519.900 19.050 520.160 19.370 ;
        RECT 1228.300 19.050 1228.560 19.370 ;
        RECT 519.960 2.400 520.100 19.050 ;
        RECT 519.750 -4.800 520.310 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 537.350 989.980 537.670 990.040 ;
        RECT 1260.470 989.980 1260.790 990.040 ;
        RECT 537.350 989.840 1260.790 989.980 ;
        RECT 537.350 989.780 537.670 989.840 ;
        RECT 1260.470 989.780 1260.790 989.840 ;
      LAYER via ;
        RECT 537.380 989.780 537.640 990.040 ;
        RECT 1260.500 989.780 1260.760 990.040 ;
      LAYER met2 ;
        RECT 1260.570 1000.620 1260.850 1004.000 ;
        RECT 1260.560 1000.000 1260.850 1000.620 ;
        RECT 1260.560 990.070 1260.700 1000.000 ;
        RECT 537.380 989.750 537.640 990.070 ;
        RECT 1260.500 989.750 1260.760 990.070 ;
        RECT 537.440 18.940 537.580 989.750 ;
        RECT 537.440 18.800 538.040 18.940 ;
        RECT 537.900 2.400 538.040 18.800 ;
        RECT 537.690 -4.800 538.250 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1292.770 1000.690 1293.050 1004.000 ;
        RECT 1290.460 1000.550 1293.050 1000.690 ;
        RECT 1290.460 17.525 1290.600 1000.550 ;
        RECT 1292.770 1000.000 1293.050 1000.550 ;
        RECT 555.770 17.155 556.050 17.525 ;
        RECT 1290.390 17.155 1290.670 17.525 ;
        RECT 555.840 2.400 555.980 17.155 ;
        RECT 555.630 -4.800 556.190 2.400 ;
      LAYER via2 ;
        RECT 555.770 17.200 556.050 17.480 ;
        RECT 1290.390 17.200 1290.670 17.480 ;
      LAYER met3 ;
        RECT 555.745 17.490 556.075 17.505 ;
        RECT 1290.365 17.490 1290.695 17.505 ;
        RECT 555.745 17.190 1290.695 17.490 ;
        RECT 555.745 17.175 556.075 17.190 ;
        RECT 1290.365 17.175 1290.695 17.190 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 573.690 25.060 574.010 25.120 ;
        RECT 579.210 25.060 579.530 25.120 ;
        RECT 573.690 24.920 579.530 25.060 ;
        RECT 573.690 24.860 574.010 24.920 ;
        RECT 579.210 24.860 579.530 24.920 ;
      LAYER via ;
        RECT 573.720 24.860 573.980 25.120 ;
        RECT 579.240 24.860 579.500 25.120 ;
      LAYER met2 ;
        RECT 1324.510 1000.620 1324.790 1004.000 ;
        RECT 1324.500 1000.000 1324.790 1000.620 ;
        RECT 1324.500 990.605 1324.640 1000.000 ;
        RECT 579.230 990.235 579.510 990.605 ;
        RECT 1324.430 990.235 1324.710 990.605 ;
        RECT 579.300 25.150 579.440 990.235 ;
        RECT 573.720 24.830 573.980 25.150 ;
        RECT 579.240 24.830 579.500 25.150 ;
        RECT 573.780 2.400 573.920 24.830 ;
        RECT 573.570 -4.800 574.130 2.400 ;
      LAYER via2 ;
        RECT 579.230 990.280 579.510 990.560 ;
        RECT 1324.430 990.280 1324.710 990.560 ;
      LAYER met3 ;
        RECT 579.205 990.570 579.535 990.585 ;
        RECT 1324.405 990.570 1324.735 990.585 ;
        RECT 579.205 990.270 1324.735 990.570 ;
        RECT 579.205 990.255 579.535 990.270 ;
        RECT 1324.405 990.255 1324.735 990.270 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 591.170 18.260 591.490 18.320 ;
        RECT 1352.470 18.260 1352.790 18.320 ;
        RECT 591.170 18.120 1352.790 18.260 ;
        RECT 591.170 18.060 591.490 18.120 ;
        RECT 1352.470 18.060 1352.790 18.120 ;
      LAYER via ;
        RECT 591.200 18.060 591.460 18.320 ;
        RECT 1352.500 18.060 1352.760 18.320 ;
      LAYER met2 ;
        RECT 1356.250 1000.690 1356.530 1004.000 ;
        RECT 1352.560 1000.550 1356.530 1000.690 ;
        RECT 1352.560 18.350 1352.700 1000.550 ;
        RECT 1356.250 1000.000 1356.530 1000.550 ;
        RECT 591.200 18.030 591.460 18.350 ;
        RECT 1352.500 18.030 1352.760 18.350 ;
        RECT 591.260 2.400 591.400 18.030 ;
        RECT 591.050 -4.800 591.610 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 103.110 990.660 103.430 990.720 ;
        RECT 474.790 990.660 475.110 990.720 ;
        RECT 103.110 990.520 475.110 990.660 ;
        RECT 103.110 990.460 103.430 990.520 ;
        RECT 474.790 990.460 475.110 990.520 ;
        RECT 97.590 17.580 97.910 17.640 ;
        RECT 103.110 17.580 103.430 17.640 ;
        RECT 97.590 17.440 103.430 17.580 ;
        RECT 97.590 17.380 97.910 17.440 ;
        RECT 103.110 17.380 103.430 17.440 ;
      LAYER via ;
        RECT 103.140 990.460 103.400 990.720 ;
        RECT 474.820 990.460 475.080 990.720 ;
        RECT 97.620 17.380 97.880 17.640 ;
        RECT 103.140 17.380 103.400 17.640 ;
      LAYER met2 ;
        RECT 474.890 1000.620 475.170 1004.000 ;
        RECT 474.880 1000.000 475.170 1000.620 ;
        RECT 474.880 990.750 475.020 1000.000 ;
        RECT 103.140 990.430 103.400 990.750 ;
        RECT 474.820 990.430 475.080 990.750 ;
        RECT 103.200 17.670 103.340 990.430 ;
        RECT 97.620 17.350 97.880 17.670 ;
        RECT 103.140 17.350 103.400 17.670 ;
        RECT 97.680 2.400 97.820 17.350 ;
        RECT 97.470 -4.800 98.030 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 609.110 17.580 609.430 17.640 ;
        RECT 1386.970 17.580 1387.290 17.640 ;
        RECT 609.110 17.440 1387.290 17.580 ;
        RECT 609.110 17.380 609.430 17.440 ;
        RECT 1386.970 17.380 1387.290 17.440 ;
      LAYER via ;
        RECT 609.140 17.380 609.400 17.640 ;
        RECT 1387.000 17.380 1387.260 17.640 ;
      LAYER met2 ;
        RECT 1388.450 1000.690 1388.730 1004.000 ;
        RECT 1387.060 1000.550 1388.730 1000.690 ;
        RECT 1387.060 17.670 1387.200 1000.550 ;
        RECT 1388.450 1000.000 1388.730 1000.550 ;
        RECT 609.140 17.350 609.400 17.670 ;
        RECT 1387.000 17.350 1387.260 17.670 ;
        RECT 609.200 2.400 609.340 17.350 ;
        RECT 608.990 -4.800 609.550 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1420.190 1000.690 1420.470 1004.000 ;
        RECT 1414.660 1000.550 1420.470 1000.690 ;
        RECT 1414.660 16.845 1414.800 1000.550 ;
        RECT 1420.190 1000.000 1420.470 1000.550 ;
        RECT 627.070 16.475 627.350 16.845 ;
        RECT 1414.590 16.475 1414.870 16.845 ;
        RECT 627.140 2.400 627.280 16.475 ;
        RECT 626.930 -4.800 627.490 2.400 ;
      LAYER via2 ;
        RECT 627.070 16.520 627.350 16.800 ;
        RECT 1414.590 16.520 1414.870 16.800 ;
      LAYER met3 ;
        RECT 627.045 16.810 627.375 16.825 ;
        RECT 1414.565 16.810 1414.895 16.825 ;
        RECT 627.045 16.510 1414.895 16.810 ;
        RECT 627.045 16.495 627.375 16.510 ;
        RECT 1414.565 16.495 1414.895 16.510 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 510.670 19.620 510.990 19.680 ;
        RECT 137.700 19.480 510.990 19.620 ;
        RECT 121.510 19.280 121.830 19.340 ;
        RECT 137.700 19.280 137.840 19.480 ;
        RECT 510.670 19.420 510.990 19.480 ;
        RECT 121.510 19.140 137.840 19.280 ;
        RECT 121.510 19.080 121.830 19.140 ;
      LAYER via ;
        RECT 121.540 19.080 121.800 19.340 ;
        RECT 510.700 19.420 510.960 19.680 ;
      LAYER met2 ;
        RECT 517.210 1000.690 517.490 1004.000 ;
        RECT 510.760 1000.550 517.490 1000.690 ;
        RECT 510.760 19.710 510.900 1000.550 ;
        RECT 517.210 1000.000 517.490 1000.550 ;
        RECT 510.700 19.390 510.960 19.710 ;
        RECT 121.540 19.050 121.800 19.370 ;
        RECT 121.600 2.400 121.740 19.050 ;
        RECT 121.390 -4.800 121.950 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 145.430 18.600 145.750 18.660 ;
        RECT 558.970 18.600 559.290 18.660 ;
        RECT 145.430 18.460 559.290 18.600 ;
        RECT 145.430 18.400 145.750 18.460 ;
        RECT 558.970 18.400 559.290 18.460 ;
      LAYER via ;
        RECT 145.460 18.400 145.720 18.660 ;
        RECT 559.000 18.400 559.260 18.660 ;
      LAYER met2 ;
        RECT 559.990 1000.690 560.270 1004.000 ;
        RECT 559.060 1000.550 560.270 1000.690 ;
        RECT 559.060 18.690 559.200 1000.550 ;
        RECT 559.990 1000.000 560.270 1000.550 ;
        RECT 145.460 18.370 145.720 18.690 ;
        RECT 559.000 18.370 559.260 18.690 ;
        RECT 145.520 2.400 145.660 18.370 ;
        RECT 145.310 -4.800 145.870 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 548.850 18.940 549.170 19.000 ;
        RECT 573.230 18.940 573.550 19.000 ;
        RECT 548.850 18.800 573.550 18.940 ;
        RECT 548.850 18.740 549.170 18.800 ;
        RECT 573.230 18.740 573.550 18.800 ;
        RECT 163.370 17.920 163.690 17.980 ;
        RECT 548.850 17.920 549.170 17.980 ;
        RECT 163.370 17.780 549.170 17.920 ;
        RECT 163.370 17.720 163.690 17.780 ;
        RECT 548.850 17.720 549.170 17.780 ;
      LAYER via ;
        RECT 548.880 18.740 549.140 19.000 ;
        RECT 573.260 18.740 573.520 19.000 ;
        RECT 163.400 17.720 163.660 17.980 ;
        RECT 548.880 17.720 549.140 17.980 ;
      LAYER met2 ;
        RECT 591.730 1000.690 592.010 1004.000 ;
        RECT 586.660 1000.550 592.010 1000.690 ;
        RECT 586.660 19.565 586.800 1000.550 ;
        RECT 591.730 1000.000 592.010 1000.550 ;
        RECT 573.250 19.195 573.530 19.565 ;
        RECT 586.590 19.195 586.870 19.565 ;
        RECT 573.320 19.030 573.460 19.195 ;
        RECT 548.880 18.710 549.140 19.030 ;
        RECT 573.260 18.710 573.520 19.030 ;
        RECT 548.940 18.010 549.080 18.710 ;
        RECT 163.400 17.690 163.660 18.010 ;
        RECT 548.880 17.690 549.140 18.010 ;
        RECT 163.460 2.400 163.600 17.690 ;
        RECT 163.250 -4.800 163.810 2.400 ;
      LAYER via2 ;
        RECT 573.250 19.240 573.530 19.520 ;
        RECT 586.590 19.240 586.870 19.520 ;
      LAYER met3 ;
        RECT 573.225 19.530 573.555 19.545 ;
        RECT 586.565 19.530 586.895 19.545 ;
        RECT 573.225 19.230 586.895 19.530 ;
        RECT 573.225 19.215 573.555 19.230 ;
        RECT 586.565 19.215 586.895 19.230 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 213.970 17.240 214.290 17.300 ;
        RECT 620.610 17.240 620.930 17.300 ;
        RECT 213.970 17.100 620.930 17.240 ;
        RECT 213.970 17.040 214.290 17.100 ;
        RECT 620.610 17.040 620.930 17.100 ;
        RECT 180.850 14.860 181.170 14.920 ;
        RECT 213.970 14.860 214.290 14.920 ;
        RECT 180.850 14.720 214.290 14.860 ;
        RECT 180.850 14.660 181.170 14.720 ;
        RECT 213.970 14.660 214.290 14.720 ;
      LAYER via ;
        RECT 214.000 17.040 214.260 17.300 ;
        RECT 620.640 17.040 620.900 17.300 ;
        RECT 180.880 14.660 181.140 14.920 ;
        RECT 214.000 14.660 214.260 14.920 ;
      LAYER met2 ;
        RECT 623.470 1000.690 623.750 1004.000 ;
        RECT 621.160 1000.550 623.750 1000.690 ;
        RECT 621.160 18.090 621.300 1000.550 ;
        RECT 623.470 1000.000 623.750 1000.550 ;
        RECT 620.700 17.950 621.300 18.090 ;
        RECT 620.700 17.330 620.840 17.950 ;
        RECT 214.000 17.010 214.260 17.330 ;
        RECT 620.640 17.010 620.900 17.330 ;
        RECT 214.060 14.950 214.200 17.010 ;
        RECT 180.880 14.630 181.140 14.950 ;
        RECT 214.000 14.630 214.260 14.950 ;
        RECT 180.940 2.400 181.080 14.630 ;
        RECT 180.730 -4.800 181.290 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 199.710 987.260 200.030 987.320 ;
        RECT 651.430 987.260 651.750 987.320 ;
        RECT 199.710 987.120 651.750 987.260 ;
        RECT 199.710 987.060 200.030 987.120 ;
        RECT 651.430 987.060 651.750 987.120 ;
      LAYER via ;
        RECT 199.740 987.060 200.000 987.320 ;
        RECT 651.460 987.060 651.720 987.320 ;
      LAYER met2 ;
        RECT 655.210 1000.690 655.490 1004.000 ;
        RECT 651.520 1000.550 655.490 1000.690 ;
        RECT 651.520 987.350 651.660 1000.550 ;
        RECT 655.210 1000.000 655.490 1000.550 ;
        RECT 199.740 987.030 200.000 987.350 ;
        RECT 651.460 987.030 651.720 987.350 ;
        RECT 199.800 17.410 199.940 987.030 ;
        RECT 198.880 17.270 199.940 17.410 ;
        RECT 198.880 2.400 199.020 17.270 ;
        RECT 198.670 -4.800 199.230 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 216.730 14.860 217.050 14.920 ;
        RECT 216.730 14.720 234.440 14.860 ;
        RECT 216.730 14.660 217.050 14.720 ;
        RECT 234.300 14.520 234.440 14.720 ;
        RECT 683.170 14.520 683.490 14.580 ;
        RECT 234.300 14.380 683.490 14.520 ;
        RECT 683.170 14.320 683.490 14.380 ;
      LAYER via ;
        RECT 216.760 14.660 217.020 14.920 ;
        RECT 683.200 14.320 683.460 14.580 ;
      LAYER met2 ;
        RECT 687.410 1000.690 687.690 1004.000 ;
        RECT 683.260 1000.550 687.690 1000.690 ;
        RECT 216.760 14.630 217.020 14.950 ;
        RECT 216.820 2.400 216.960 14.630 ;
        RECT 683.260 14.610 683.400 1000.550 ;
        RECT 687.410 1000.000 687.690 1000.550 ;
        RECT 683.200 14.290 683.460 14.610 ;
        RECT 216.610 -4.800 217.170 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 240.650 987.940 240.970 988.000 ;
        RECT 719.050 987.940 719.370 988.000 ;
        RECT 240.650 987.800 719.370 987.940 ;
        RECT 240.650 987.740 240.970 987.800 ;
        RECT 719.050 987.740 719.370 987.800 ;
        RECT 234.670 14.860 234.990 14.920 ;
        RECT 240.650 14.860 240.970 14.920 ;
        RECT 234.670 14.720 240.970 14.860 ;
        RECT 234.670 14.660 234.990 14.720 ;
        RECT 240.650 14.660 240.970 14.720 ;
      LAYER via ;
        RECT 240.680 987.740 240.940 988.000 ;
        RECT 719.080 987.740 719.340 988.000 ;
        RECT 234.700 14.660 234.960 14.920 ;
        RECT 240.680 14.660 240.940 14.920 ;
      LAYER met2 ;
        RECT 719.150 1000.620 719.430 1004.000 ;
        RECT 719.140 1000.000 719.430 1000.620 ;
        RECT 719.140 988.030 719.280 1000.000 ;
        RECT 240.680 987.710 240.940 988.030 ;
        RECT 719.080 987.710 719.340 988.030 ;
        RECT 240.740 14.950 240.880 987.710 ;
        RECT 234.700 14.630 234.960 14.950 ;
        RECT 240.680 14.630 240.940 14.950 ;
        RECT 234.760 2.400 234.900 14.630 ;
        RECT 234.550 -4.800 235.110 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 61.710 991.680 62.030 991.740 ;
        RECT 400.270 991.680 400.590 991.740 ;
        RECT 61.710 991.540 400.590 991.680 ;
        RECT 61.710 991.480 62.030 991.540 ;
        RECT 400.270 991.480 400.590 991.540 ;
        RECT 56.190 17.580 56.510 17.640 ;
        RECT 61.710 17.580 62.030 17.640 ;
        RECT 56.190 17.440 62.030 17.580 ;
        RECT 56.190 17.380 56.510 17.440 ;
        RECT 61.710 17.380 62.030 17.440 ;
      LAYER via ;
        RECT 61.740 991.480 62.000 991.740 ;
        RECT 400.300 991.480 400.560 991.740 ;
        RECT 56.220 17.380 56.480 17.640 ;
        RECT 61.740 17.380 62.000 17.640 ;
      LAYER met2 ;
        RECT 400.370 1000.620 400.650 1004.000 ;
        RECT 400.360 1000.000 400.650 1000.620 ;
        RECT 400.360 991.770 400.500 1000.000 ;
        RECT 61.740 991.450 62.000 991.770 ;
        RECT 400.300 991.450 400.560 991.770 ;
        RECT 61.800 17.670 61.940 991.450 ;
        RECT 56.220 17.350 56.480 17.670 ;
        RECT 61.740 17.350 62.000 17.670 ;
        RECT 56.280 2.400 56.420 17.350 ;
        RECT 56.070 -4.800 56.630 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 82.410 991.000 82.730 991.060 ;
        RECT 443.050 991.000 443.370 991.060 ;
        RECT 82.410 990.860 443.370 991.000 ;
        RECT 82.410 990.800 82.730 990.860 ;
        RECT 443.050 990.800 443.370 990.860 ;
        RECT 80.110 17.580 80.430 17.640 ;
        RECT 82.410 17.580 82.730 17.640 ;
        RECT 80.110 17.440 82.730 17.580 ;
        RECT 80.110 17.380 80.430 17.440 ;
        RECT 82.410 17.380 82.730 17.440 ;
      LAYER via ;
        RECT 82.440 990.800 82.700 991.060 ;
        RECT 443.080 990.800 443.340 991.060 ;
        RECT 80.140 17.380 80.400 17.640 ;
        RECT 82.440 17.380 82.700 17.640 ;
      LAYER met2 ;
        RECT 443.150 1000.620 443.430 1004.000 ;
        RECT 443.140 1000.000 443.430 1000.620 ;
        RECT 443.140 991.090 443.280 1000.000 ;
        RECT 82.440 990.770 82.700 991.090 ;
        RECT 443.080 990.770 443.340 991.090 ;
        RECT 82.500 17.670 82.640 990.770 ;
        RECT 80.140 17.350 80.400 17.670 ;
        RECT 82.440 17.350 82.700 17.670 ;
        RECT 80.200 2.400 80.340 17.350 ;
        RECT 79.990 -4.800 80.550 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 109.550 990.320 109.870 990.380 ;
        RECT 485.370 990.320 485.690 990.380 ;
        RECT 109.550 990.180 485.690 990.320 ;
        RECT 109.550 990.120 109.870 990.180 ;
        RECT 485.370 990.120 485.690 990.180 ;
        RECT 103.570 17.580 103.890 17.640 ;
        RECT 109.550 17.580 109.870 17.640 ;
        RECT 103.570 17.440 109.870 17.580 ;
        RECT 103.570 17.380 103.890 17.440 ;
        RECT 109.550 17.380 109.870 17.440 ;
      LAYER via ;
        RECT 109.580 990.120 109.840 990.380 ;
        RECT 485.400 990.120 485.660 990.380 ;
        RECT 103.600 17.380 103.860 17.640 ;
        RECT 109.580 17.380 109.840 17.640 ;
      LAYER met2 ;
        RECT 485.470 1000.620 485.750 1004.000 ;
        RECT 485.460 1000.000 485.750 1000.620 ;
        RECT 485.460 990.410 485.600 1000.000 ;
        RECT 109.580 990.090 109.840 990.410 ;
        RECT 485.400 990.090 485.660 990.410 ;
        RECT 109.640 17.670 109.780 990.090 ;
        RECT 103.600 17.350 103.860 17.670 ;
        RECT 109.580 17.350 109.840 17.670 ;
        RECT 103.660 2.400 103.800 17.350 ;
        RECT 103.450 -4.800 104.010 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 130.710 989.980 131.030 990.040 ;
        RECT 527.690 989.980 528.010 990.040 ;
        RECT 130.710 989.840 528.010 989.980 ;
        RECT 130.710 989.780 131.030 989.840 ;
        RECT 527.690 989.780 528.010 989.840 ;
        RECT 127.490 17.580 127.810 17.640 ;
        RECT 130.710 17.580 131.030 17.640 ;
        RECT 127.490 17.440 131.030 17.580 ;
        RECT 127.490 17.380 127.810 17.440 ;
        RECT 130.710 17.380 131.030 17.440 ;
      LAYER via ;
        RECT 130.740 989.780 131.000 990.040 ;
        RECT 527.720 989.780 527.980 990.040 ;
        RECT 127.520 17.380 127.780 17.640 ;
        RECT 130.740 17.380 131.000 17.640 ;
      LAYER met2 ;
        RECT 527.790 1000.620 528.070 1004.000 ;
        RECT 527.780 1000.000 528.070 1000.620 ;
        RECT 527.780 990.070 527.920 1000.000 ;
        RECT 130.740 989.750 131.000 990.070 ;
        RECT 527.720 989.750 527.980 990.070 ;
        RECT 130.800 17.670 130.940 989.750 ;
        RECT 127.520 17.350 127.780 17.670 ;
        RECT 130.740 17.350 131.000 17.670 ;
        RECT 127.580 2.400 127.720 17.350 ;
        RECT 127.370 -4.800 127.930 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 161.990 992.360 162.310 992.420 ;
        RECT 347.370 992.360 347.690 992.420 ;
        RECT 161.990 992.220 347.690 992.360 ;
        RECT 161.990 992.160 162.310 992.220 ;
        RECT 347.370 992.160 347.690 992.220 ;
        RECT 26.290 17.240 26.610 17.300 ;
        RECT 161.990 17.240 162.310 17.300 ;
        RECT 26.290 17.100 162.310 17.240 ;
        RECT 26.290 17.040 26.610 17.100 ;
        RECT 161.990 17.040 162.310 17.100 ;
      LAYER via ;
        RECT 162.020 992.160 162.280 992.420 ;
        RECT 347.400 992.160 347.660 992.420 ;
        RECT 26.320 17.040 26.580 17.300 ;
        RECT 162.020 17.040 162.280 17.300 ;
      LAYER met2 ;
        RECT 347.470 1000.620 347.750 1004.000 ;
        RECT 347.460 1000.000 347.750 1000.620 ;
        RECT 347.460 992.450 347.600 1000.000 ;
        RECT 162.020 992.130 162.280 992.450 ;
        RECT 347.400 992.130 347.660 992.450 ;
        RECT 162.080 17.330 162.220 992.130 ;
        RECT 26.320 17.010 26.580 17.330 ;
        RECT 162.020 17.010 162.280 17.330 ;
        RECT 26.380 2.400 26.520 17.010 ;
        RECT 26.170 -4.800 26.730 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 352.430 16.900 352.750 16.960 ;
        RECT 327.680 16.760 352.750 16.900 ;
        RECT 32.270 16.560 32.590 16.620 ;
        RECT 327.680 16.560 327.820 16.760 ;
        RECT 352.430 16.700 352.750 16.760 ;
        RECT 32.270 16.420 327.820 16.560 ;
        RECT 32.270 16.360 32.590 16.420 ;
      LAYER via ;
        RECT 32.300 16.360 32.560 16.620 ;
        RECT 352.460 16.700 352.720 16.960 ;
      LAYER met2 ;
        RECT 358.050 1000.690 358.330 1004.000 ;
        RECT 352.520 1000.550 358.330 1000.690 ;
        RECT 352.520 16.990 352.660 1000.550 ;
        RECT 358.050 1000.000 358.330 1000.550 ;
        RECT 352.460 16.670 352.720 16.990 ;
        RECT 32.300 16.330 32.560 16.650 ;
        RECT 32.360 2.400 32.500 16.330 ;
        RECT 32.150 -4.800 32.710 2.400 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 681.480 2743.600 684.050 2744.660 ;
        RECT 1331.480 2743.600 1334.050 2744.660 ;
        RECT 1931.480 2743.600 1934.050 2744.660 ;
        RECT 2581.480 2743.600 2584.050 2744.660 ;
      LAYER via3 ;
        RECT 682.500 2743.620 684.020 2744.630 ;
        RECT 1332.500 2743.620 1334.020 2744.630 ;
        RECT 1932.500 2743.620 1934.020 2744.630 ;
        RECT 2582.500 2743.620 2584.020 2744.630 ;
      LAYER met4 ;
        RECT -38.180 -32.820 -35.180 3552.500 ;
        RECT -28.780 -23.420 -25.780 3543.100 ;
        RECT -19.380 -14.020 -16.380 3533.700 ;
        RECT -9.980 -4.620 -6.980 3524.300 ;
        RECT 4.020 -9.320 7.020 3529.000 ;
        RECT 22.020 -18.720 25.020 3538.400 ;
        RECT 40.020 -28.120 43.020 3547.800 ;
        RECT 58.020 -37.520 61.020 3557.200 ;
        RECT 184.020 -9.320 187.020 3529.000 ;
        RECT 202.020 -18.720 205.020 3538.400 ;
        RECT 220.020 -28.120 223.020 3547.800 ;
        RECT 238.020 -37.520 241.020 3557.200 ;
        RECT 364.020 2771.235 367.020 3529.000 ;
        RECT 382.020 2771.235 385.020 3538.400 ;
        RECT 400.020 2771.235 403.020 3547.800 ;
        RECT 418.020 2771.235 421.020 3557.200 ;
        RECT 544.020 2771.235 547.020 3529.000 ;
        RECT 562.020 2771.235 565.020 3538.400 ;
        RECT 580.020 2771.235 583.020 3547.800 ;
        RECT 598.020 2771.235 601.020 3557.200 ;
        RECT 682.470 2303.670 684.070 2744.680 ;
        RECT 418.020 2215.000 421.020 2285.000 ;
        RECT 598.020 2215.000 601.020 2285.000 ;
        RECT 724.020 2215.000 727.020 3529.000 ;
        RECT 742.020 2215.000 745.020 3538.400 ;
        RECT 760.020 2215.000 763.020 3547.800 ;
        RECT 778.020 2215.000 781.020 3557.200 ;
        RECT 904.020 2215.000 907.020 3529.000 ;
        RECT 922.020 2215.000 925.020 3538.400 ;
        RECT 940.020 2771.235 943.020 3547.800 ;
        RECT 958.020 2771.235 961.020 3557.200 ;
        RECT 1084.020 2771.235 1087.020 3529.000 ;
        RECT 1102.020 2771.235 1105.020 3538.400 ;
        RECT 1120.020 2771.235 1123.020 3547.800 ;
        RECT 1138.020 2771.235 1141.020 3557.200 ;
        RECT 1264.020 2771.235 1267.020 3529.000 ;
        RECT 1282.020 2771.235 1285.020 3538.400 ;
        RECT 1300.020 2771.235 1303.020 3547.800 ;
        RECT 1318.020 2771.235 1321.020 3557.200 ;
        RECT 1332.470 2303.670 1334.070 2744.680 ;
        RECT 958.020 2215.000 961.020 2285.000 ;
        RECT 1138.020 2215.000 1141.020 2285.000 ;
        RECT 1318.020 2215.000 1321.020 2285.000 ;
        RECT 1444.020 2215.000 1447.020 3529.000 ;
        RECT 1462.020 2215.000 1465.020 3538.400 ;
        RECT 1480.020 2215.000 1483.020 3547.800 ;
        RECT 1498.020 2215.000 1501.020 3557.200 ;
        RECT 1624.020 2771.235 1627.020 3529.000 ;
        RECT 1642.020 2771.235 1645.020 3538.400 ;
        RECT 1660.020 2771.235 1663.020 3547.800 ;
        RECT 1678.020 2771.235 1681.020 3557.200 ;
        RECT 1804.020 2771.235 1807.020 3529.000 ;
        RECT 1822.020 2771.235 1825.020 3538.400 ;
        RECT 1840.020 2771.235 1843.020 3547.800 ;
        RECT 1858.020 2771.235 1861.020 3557.200 ;
        RECT 1932.470 2303.670 1934.070 2744.680 ;
        RECT 321.040 1010.640 322.640 2188.880 ;
        RECT 364.020 -9.320 367.020 985.000 ;
        RECT 382.020 -18.720 385.020 985.000 ;
        RECT 400.020 -28.120 403.020 985.000 ;
        RECT 418.020 -37.520 421.020 985.000 ;
        RECT 544.020 -9.320 547.020 985.000 ;
        RECT 562.020 -18.720 565.020 985.000 ;
        RECT 580.020 -28.120 583.020 985.000 ;
        RECT 598.020 -37.520 601.020 985.000 ;
        RECT 724.020 -9.320 727.020 985.000 ;
        RECT 742.020 -18.720 745.020 985.000 ;
        RECT 760.020 -28.120 763.020 985.000 ;
        RECT 778.020 -37.520 781.020 985.000 ;
        RECT 904.020 -9.320 907.020 985.000 ;
        RECT 922.020 -18.720 925.020 985.000 ;
        RECT 940.020 -28.120 943.020 985.000 ;
        RECT 958.020 -37.520 961.020 985.000 ;
        RECT 1084.020 -9.320 1087.020 985.000 ;
        RECT 1102.020 -18.720 1105.020 985.000 ;
        RECT 1120.020 -28.120 1123.020 985.000 ;
        RECT 1138.020 -37.520 1141.020 985.000 ;
        RECT 1264.020 -9.320 1267.020 985.000 ;
        RECT 1282.020 -18.720 1285.020 985.000 ;
        RECT 1300.020 -28.120 1303.020 985.000 ;
        RECT 1318.020 -37.520 1321.020 985.000 ;
        RECT 1444.020 -9.320 1447.020 985.000 ;
        RECT 1462.020 -18.720 1465.020 985.000 ;
        RECT 1480.020 -28.120 1483.020 985.000 ;
        RECT 1498.020 -37.520 1501.020 985.000 ;
        RECT 1624.020 -9.320 1627.020 2285.000 ;
        RECT 1642.020 -18.720 1645.020 2285.000 ;
        RECT 1660.020 -28.120 1663.020 2285.000 ;
        RECT 1678.020 -37.520 1681.020 2285.000 ;
        RECT 1804.020 -9.320 1807.020 2285.000 ;
        RECT 1822.020 -18.720 1825.020 2285.000 ;
        RECT 1840.020 -28.120 1843.020 2285.000 ;
        RECT 1858.020 -37.520 1861.020 2285.000 ;
        RECT 1984.020 -9.320 1987.020 3529.000 ;
        RECT 2002.020 -18.720 2005.020 3538.400 ;
        RECT 2020.020 -28.120 2023.020 3547.800 ;
        RECT 2038.020 -37.520 2041.020 3557.200 ;
        RECT 2164.020 -9.320 2167.020 3529.000 ;
        RECT 2182.020 2771.235 2185.020 3538.400 ;
        RECT 2200.020 2771.235 2203.020 3547.800 ;
        RECT 2218.020 2771.235 2221.020 3557.200 ;
        RECT 2344.020 2771.235 2347.020 3529.000 ;
        RECT 2362.020 2771.235 2365.020 3538.400 ;
        RECT 2380.020 2771.235 2383.020 3547.800 ;
        RECT 2398.020 2771.235 2401.020 3557.200 ;
        RECT 2524.020 2771.235 2527.020 3529.000 ;
        RECT 2542.020 2771.235 2545.020 3538.400 ;
        RECT 2560.020 2771.235 2563.020 3547.800 ;
        RECT 2578.020 2771.235 2581.020 3557.200 ;
        RECT 2582.470 2303.670 2584.070 2744.680 ;
        RECT 2182.020 -18.720 2185.020 2285.000 ;
        RECT 2200.020 -28.120 2203.020 2285.000 ;
        RECT 2218.020 -37.520 2221.020 2285.000 ;
        RECT 2344.020 -9.320 2347.020 2285.000 ;
        RECT 2362.020 -18.720 2365.020 2285.000 ;
        RECT 2380.020 -28.120 2383.020 2285.000 ;
        RECT 2398.020 -37.520 2401.020 2285.000 ;
        RECT 2524.020 -9.320 2527.020 2285.000 ;
        RECT 2542.020 -18.720 2545.020 2285.000 ;
        RECT 2560.020 -28.120 2563.020 2285.000 ;
        RECT 2578.020 -37.520 2581.020 2285.000 ;
        RECT 2704.020 -9.320 2707.020 3529.000 ;
        RECT 2722.020 -18.720 2725.020 3538.400 ;
        RECT 2740.020 -28.120 2743.020 3547.800 ;
        RECT 2758.020 -37.520 2761.020 3557.200 ;
        RECT 2884.020 -9.320 2887.020 3529.000 ;
        RECT 2902.020 -18.720 2905.020 3538.400 ;
        RECT 2926.600 -4.620 2929.600 3524.300 ;
        RECT 2936.000 -14.020 2939.000 3533.700 ;
        RECT 2945.400 -23.420 2948.400 3543.100 ;
        RECT 2954.800 -32.820 2957.800 3552.500 ;
      LAYER via4 ;
        RECT -37.270 3551.210 -36.090 3552.390 ;
        RECT -37.270 3549.610 -36.090 3550.790 ;
        RECT 58.930 3551.210 60.110 3552.390 ;
        RECT 58.930 3549.610 60.110 3550.790 ;
        RECT -37.270 3485.090 -36.090 3486.270 ;
        RECT -37.270 3483.490 -36.090 3484.670 ;
        RECT -37.270 3305.090 -36.090 3306.270 ;
        RECT -37.270 3303.490 -36.090 3304.670 ;
        RECT -37.270 3125.090 -36.090 3126.270 ;
        RECT -37.270 3123.490 -36.090 3124.670 ;
        RECT -37.270 2945.090 -36.090 2946.270 ;
        RECT -37.270 2943.490 -36.090 2944.670 ;
        RECT -37.270 2765.090 -36.090 2766.270 ;
        RECT -37.270 2763.490 -36.090 2764.670 ;
        RECT -37.270 2585.090 -36.090 2586.270 ;
        RECT -37.270 2583.490 -36.090 2584.670 ;
        RECT -37.270 2405.090 -36.090 2406.270 ;
        RECT -37.270 2403.490 -36.090 2404.670 ;
        RECT -37.270 2225.090 -36.090 2226.270 ;
        RECT -37.270 2223.490 -36.090 2224.670 ;
        RECT -37.270 2045.090 -36.090 2046.270 ;
        RECT -37.270 2043.490 -36.090 2044.670 ;
        RECT -37.270 1865.090 -36.090 1866.270 ;
        RECT -37.270 1863.490 -36.090 1864.670 ;
        RECT -37.270 1685.090 -36.090 1686.270 ;
        RECT -37.270 1683.490 -36.090 1684.670 ;
        RECT -37.270 1505.090 -36.090 1506.270 ;
        RECT -37.270 1503.490 -36.090 1504.670 ;
        RECT -37.270 1325.090 -36.090 1326.270 ;
        RECT -37.270 1323.490 -36.090 1324.670 ;
        RECT -37.270 1145.090 -36.090 1146.270 ;
        RECT -37.270 1143.490 -36.090 1144.670 ;
        RECT -37.270 965.090 -36.090 966.270 ;
        RECT -37.270 963.490 -36.090 964.670 ;
        RECT -37.270 785.090 -36.090 786.270 ;
        RECT -37.270 783.490 -36.090 784.670 ;
        RECT -37.270 605.090 -36.090 606.270 ;
        RECT -37.270 603.490 -36.090 604.670 ;
        RECT -37.270 425.090 -36.090 426.270 ;
        RECT -37.270 423.490 -36.090 424.670 ;
        RECT -37.270 245.090 -36.090 246.270 ;
        RECT -37.270 243.490 -36.090 244.670 ;
        RECT -37.270 65.090 -36.090 66.270 ;
        RECT -37.270 63.490 -36.090 64.670 ;
        RECT -27.870 3541.810 -26.690 3542.990 ;
        RECT -27.870 3540.210 -26.690 3541.390 ;
        RECT 40.930 3541.810 42.110 3542.990 ;
        RECT 40.930 3540.210 42.110 3541.390 ;
        RECT -27.870 3467.090 -26.690 3468.270 ;
        RECT -27.870 3465.490 -26.690 3466.670 ;
        RECT -27.870 3287.090 -26.690 3288.270 ;
        RECT -27.870 3285.490 -26.690 3286.670 ;
        RECT -27.870 3107.090 -26.690 3108.270 ;
        RECT -27.870 3105.490 -26.690 3106.670 ;
        RECT -27.870 2927.090 -26.690 2928.270 ;
        RECT -27.870 2925.490 -26.690 2926.670 ;
        RECT -27.870 2747.090 -26.690 2748.270 ;
        RECT -27.870 2745.490 -26.690 2746.670 ;
        RECT -27.870 2567.090 -26.690 2568.270 ;
        RECT -27.870 2565.490 -26.690 2566.670 ;
        RECT -27.870 2387.090 -26.690 2388.270 ;
        RECT -27.870 2385.490 -26.690 2386.670 ;
        RECT -27.870 2207.090 -26.690 2208.270 ;
        RECT -27.870 2205.490 -26.690 2206.670 ;
        RECT -27.870 2027.090 -26.690 2028.270 ;
        RECT -27.870 2025.490 -26.690 2026.670 ;
        RECT -27.870 1847.090 -26.690 1848.270 ;
        RECT -27.870 1845.490 -26.690 1846.670 ;
        RECT -27.870 1667.090 -26.690 1668.270 ;
        RECT -27.870 1665.490 -26.690 1666.670 ;
        RECT -27.870 1487.090 -26.690 1488.270 ;
        RECT -27.870 1485.490 -26.690 1486.670 ;
        RECT -27.870 1307.090 -26.690 1308.270 ;
        RECT -27.870 1305.490 -26.690 1306.670 ;
        RECT -27.870 1127.090 -26.690 1128.270 ;
        RECT -27.870 1125.490 -26.690 1126.670 ;
        RECT -27.870 947.090 -26.690 948.270 ;
        RECT -27.870 945.490 -26.690 946.670 ;
        RECT -27.870 767.090 -26.690 768.270 ;
        RECT -27.870 765.490 -26.690 766.670 ;
        RECT -27.870 587.090 -26.690 588.270 ;
        RECT -27.870 585.490 -26.690 586.670 ;
        RECT -27.870 407.090 -26.690 408.270 ;
        RECT -27.870 405.490 -26.690 406.670 ;
        RECT -27.870 227.090 -26.690 228.270 ;
        RECT -27.870 225.490 -26.690 226.670 ;
        RECT -27.870 47.090 -26.690 48.270 ;
        RECT -27.870 45.490 -26.690 46.670 ;
        RECT -18.470 3532.410 -17.290 3533.590 ;
        RECT -18.470 3530.810 -17.290 3531.990 ;
        RECT 22.930 3532.410 24.110 3533.590 ;
        RECT 22.930 3530.810 24.110 3531.990 ;
        RECT -18.470 3449.090 -17.290 3450.270 ;
        RECT -18.470 3447.490 -17.290 3448.670 ;
        RECT -18.470 3269.090 -17.290 3270.270 ;
        RECT -18.470 3267.490 -17.290 3268.670 ;
        RECT -18.470 3089.090 -17.290 3090.270 ;
        RECT -18.470 3087.490 -17.290 3088.670 ;
        RECT -18.470 2909.090 -17.290 2910.270 ;
        RECT -18.470 2907.490 -17.290 2908.670 ;
        RECT -18.470 2729.090 -17.290 2730.270 ;
        RECT -18.470 2727.490 -17.290 2728.670 ;
        RECT -18.470 2549.090 -17.290 2550.270 ;
        RECT -18.470 2547.490 -17.290 2548.670 ;
        RECT -18.470 2369.090 -17.290 2370.270 ;
        RECT -18.470 2367.490 -17.290 2368.670 ;
        RECT -18.470 2189.090 -17.290 2190.270 ;
        RECT -18.470 2187.490 -17.290 2188.670 ;
        RECT -18.470 2009.090 -17.290 2010.270 ;
        RECT -18.470 2007.490 -17.290 2008.670 ;
        RECT -18.470 1829.090 -17.290 1830.270 ;
        RECT -18.470 1827.490 -17.290 1828.670 ;
        RECT -18.470 1649.090 -17.290 1650.270 ;
        RECT -18.470 1647.490 -17.290 1648.670 ;
        RECT -18.470 1469.090 -17.290 1470.270 ;
        RECT -18.470 1467.490 -17.290 1468.670 ;
        RECT -18.470 1289.090 -17.290 1290.270 ;
        RECT -18.470 1287.490 -17.290 1288.670 ;
        RECT -18.470 1109.090 -17.290 1110.270 ;
        RECT -18.470 1107.490 -17.290 1108.670 ;
        RECT -18.470 929.090 -17.290 930.270 ;
        RECT -18.470 927.490 -17.290 928.670 ;
        RECT -18.470 749.090 -17.290 750.270 ;
        RECT -18.470 747.490 -17.290 748.670 ;
        RECT -18.470 569.090 -17.290 570.270 ;
        RECT -18.470 567.490 -17.290 568.670 ;
        RECT -18.470 389.090 -17.290 390.270 ;
        RECT -18.470 387.490 -17.290 388.670 ;
        RECT -18.470 209.090 -17.290 210.270 ;
        RECT -18.470 207.490 -17.290 208.670 ;
        RECT -18.470 29.090 -17.290 30.270 ;
        RECT -18.470 27.490 -17.290 28.670 ;
        RECT -9.070 3523.010 -7.890 3524.190 ;
        RECT -9.070 3521.410 -7.890 3522.590 ;
        RECT -9.070 3431.090 -7.890 3432.270 ;
        RECT -9.070 3429.490 -7.890 3430.670 ;
        RECT -9.070 3251.090 -7.890 3252.270 ;
        RECT -9.070 3249.490 -7.890 3250.670 ;
        RECT -9.070 3071.090 -7.890 3072.270 ;
        RECT -9.070 3069.490 -7.890 3070.670 ;
        RECT -9.070 2891.090 -7.890 2892.270 ;
        RECT -9.070 2889.490 -7.890 2890.670 ;
        RECT -9.070 2711.090 -7.890 2712.270 ;
        RECT -9.070 2709.490 -7.890 2710.670 ;
        RECT -9.070 2531.090 -7.890 2532.270 ;
        RECT -9.070 2529.490 -7.890 2530.670 ;
        RECT -9.070 2351.090 -7.890 2352.270 ;
        RECT -9.070 2349.490 -7.890 2350.670 ;
        RECT -9.070 2171.090 -7.890 2172.270 ;
        RECT -9.070 2169.490 -7.890 2170.670 ;
        RECT -9.070 1991.090 -7.890 1992.270 ;
        RECT -9.070 1989.490 -7.890 1990.670 ;
        RECT -9.070 1811.090 -7.890 1812.270 ;
        RECT -9.070 1809.490 -7.890 1810.670 ;
        RECT -9.070 1631.090 -7.890 1632.270 ;
        RECT -9.070 1629.490 -7.890 1630.670 ;
        RECT -9.070 1451.090 -7.890 1452.270 ;
        RECT -9.070 1449.490 -7.890 1450.670 ;
        RECT -9.070 1271.090 -7.890 1272.270 ;
        RECT -9.070 1269.490 -7.890 1270.670 ;
        RECT -9.070 1091.090 -7.890 1092.270 ;
        RECT -9.070 1089.490 -7.890 1090.670 ;
        RECT -9.070 911.090 -7.890 912.270 ;
        RECT -9.070 909.490 -7.890 910.670 ;
        RECT -9.070 731.090 -7.890 732.270 ;
        RECT -9.070 729.490 -7.890 730.670 ;
        RECT -9.070 551.090 -7.890 552.270 ;
        RECT -9.070 549.490 -7.890 550.670 ;
        RECT -9.070 371.090 -7.890 372.270 ;
        RECT -9.070 369.490 -7.890 370.670 ;
        RECT -9.070 191.090 -7.890 192.270 ;
        RECT -9.070 189.490 -7.890 190.670 ;
        RECT -9.070 11.090 -7.890 12.270 ;
        RECT -9.070 9.490 -7.890 10.670 ;
        RECT -9.070 -2.910 -7.890 -1.730 ;
        RECT -9.070 -4.510 -7.890 -3.330 ;
        RECT 4.930 3523.010 6.110 3524.190 ;
        RECT 4.930 3521.410 6.110 3522.590 ;
        RECT 4.930 3431.090 6.110 3432.270 ;
        RECT 4.930 3429.490 6.110 3430.670 ;
        RECT 4.930 3251.090 6.110 3252.270 ;
        RECT 4.930 3249.490 6.110 3250.670 ;
        RECT 4.930 3071.090 6.110 3072.270 ;
        RECT 4.930 3069.490 6.110 3070.670 ;
        RECT 4.930 2891.090 6.110 2892.270 ;
        RECT 4.930 2889.490 6.110 2890.670 ;
        RECT 4.930 2711.090 6.110 2712.270 ;
        RECT 4.930 2709.490 6.110 2710.670 ;
        RECT 4.930 2531.090 6.110 2532.270 ;
        RECT 4.930 2529.490 6.110 2530.670 ;
        RECT 4.930 2351.090 6.110 2352.270 ;
        RECT 4.930 2349.490 6.110 2350.670 ;
        RECT 4.930 2171.090 6.110 2172.270 ;
        RECT 4.930 2169.490 6.110 2170.670 ;
        RECT 4.930 1991.090 6.110 1992.270 ;
        RECT 4.930 1989.490 6.110 1990.670 ;
        RECT 4.930 1811.090 6.110 1812.270 ;
        RECT 4.930 1809.490 6.110 1810.670 ;
        RECT 4.930 1631.090 6.110 1632.270 ;
        RECT 4.930 1629.490 6.110 1630.670 ;
        RECT 4.930 1451.090 6.110 1452.270 ;
        RECT 4.930 1449.490 6.110 1450.670 ;
        RECT 4.930 1271.090 6.110 1272.270 ;
        RECT 4.930 1269.490 6.110 1270.670 ;
        RECT 4.930 1091.090 6.110 1092.270 ;
        RECT 4.930 1089.490 6.110 1090.670 ;
        RECT 4.930 911.090 6.110 912.270 ;
        RECT 4.930 909.490 6.110 910.670 ;
        RECT 4.930 731.090 6.110 732.270 ;
        RECT 4.930 729.490 6.110 730.670 ;
        RECT 4.930 551.090 6.110 552.270 ;
        RECT 4.930 549.490 6.110 550.670 ;
        RECT 4.930 371.090 6.110 372.270 ;
        RECT 4.930 369.490 6.110 370.670 ;
        RECT 4.930 191.090 6.110 192.270 ;
        RECT 4.930 189.490 6.110 190.670 ;
        RECT 4.930 11.090 6.110 12.270 ;
        RECT 4.930 9.490 6.110 10.670 ;
        RECT 4.930 -2.910 6.110 -1.730 ;
        RECT 4.930 -4.510 6.110 -3.330 ;
        RECT 22.930 3449.090 24.110 3450.270 ;
        RECT 22.930 3447.490 24.110 3448.670 ;
        RECT 22.930 3269.090 24.110 3270.270 ;
        RECT 22.930 3267.490 24.110 3268.670 ;
        RECT 22.930 3089.090 24.110 3090.270 ;
        RECT 22.930 3087.490 24.110 3088.670 ;
        RECT 22.930 2909.090 24.110 2910.270 ;
        RECT 22.930 2907.490 24.110 2908.670 ;
        RECT 22.930 2729.090 24.110 2730.270 ;
        RECT 22.930 2727.490 24.110 2728.670 ;
        RECT 22.930 2549.090 24.110 2550.270 ;
        RECT 22.930 2547.490 24.110 2548.670 ;
        RECT 22.930 2369.090 24.110 2370.270 ;
        RECT 22.930 2367.490 24.110 2368.670 ;
        RECT 22.930 2189.090 24.110 2190.270 ;
        RECT 22.930 2187.490 24.110 2188.670 ;
        RECT 22.930 2009.090 24.110 2010.270 ;
        RECT 22.930 2007.490 24.110 2008.670 ;
        RECT 22.930 1829.090 24.110 1830.270 ;
        RECT 22.930 1827.490 24.110 1828.670 ;
        RECT 22.930 1649.090 24.110 1650.270 ;
        RECT 22.930 1647.490 24.110 1648.670 ;
        RECT 22.930 1469.090 24.110 1470.270 ;
        RECT 22.930 1467.490 24.110 1468.670 ;
        RECT 22.930 1289.090 24.110 1290.270 ;
        RECT 22.930 1287.490 24.110 1288.670 ;
        RECT 22.930 1109.090 24.110 1110.270 ;
        RECT 22.930 1107.490 24.110 1108.670 ;
        RECT 22.930 929.090 24.110 930.270 ;
        RECT 22.930 927.490 24.110 928.670 ;
        RECT 22.930 749.090 24.110 750.270 ;
        RECT 22.930 747.490 24.110 748.670 ;
        RECT 22.930 569.090 24.110 570.270 ;
        RECT 22.930 567.490 24.110 568.670 ;
        RECT 22.930 389.090 24.110 390.270 ;
        RECT 22.930 387.490 24.110 388.670 ;
        RECT 22.930 209.090 24.110 210.270 ;
        RECT 22.930 207.490 24.110 208.670 ;
        RECT 22.930 29.090 24.110 30.270 ;
        RECT 22.930 27.490 24.110 28.670 ;
        RECT -18.470 -12.310 -17.290 -11.130 ;
        RECT -18.470 -13.910 -17.290 -12.730 ;
        RECT 22.930 -12.310 24.110 -11.130 ;
        RECT 22.930 -13.910 24.110 -12.730 ;
        RECT 40.930 3467.090 42.110 3468.270 ;
        RECT 40.930 3465.490 42.110 3466.670 ;
        RECT 40.930 3287.090 42.110 3288.270 ;
        RECT 40.930 3285.490 42.110 3286.670 ;
        RECT 40.930 3107.090 42.110 3108.270 ;
        RECT 40.930 3105.490 42.110 3106.670 ;
        RECT 40.930 2927.090 42.110 2928.270 ;
        RECT 40.930 2925.490 42.110 2926.670 ;
        RECT 40.930 2747.090 42.110 2748.270 ;
        RECT 40.930 2745.490 42.110 2746.670 ;
        RECT 40.930 2567.090 42.110 2568.270 ;
        RECT 40.930 2565.490 42.110 2566.670 ;
        RECT 40.930 2387.090 42.110 2388.270 ;
        RECT 40.930 2385.490 42.110 2386.670 ;
        RECT 40.930 2207.090 42.110 2208.270 ;
        RECT 40.930 2205.490 42.110 2206.670 ;
        RECT 40.930 2027.090 42.110 2028.270 ;
        RECT 40.930 2025.490 42.110 2026.670 ;
        RECT 40.930 1847.090 42.110 1848.270 ;
        RECT 40.930 1845.490 42.110 1846.670 ;
        RECT 40.930 1667.090 42.110 1668.270 ;
        RECT 40.930 1665.490 42.110 1666.670 ;
        RECT 40.930 1487.090 42.110 1488.270 ;
        RECT 40.930 1485.490 42.110 1486.670 ;
        RECT 40.930 1307.090 42.110 1308.270 ;
        RECT 40.930 1305.490 42.110 1306.670 ;
        RECT 40.930 1127.090 42.110 1128.270 ;
        RECT 40.930 1125.490 42.110 1126.670 ;
        RECT 40.930 947.090 42.110 948.270 ;
        RECT 40.930 945.490 42.110 946.670 ;
        RECT 40.930 767.090 42.110 768.270 ;
        RECT 40.930 765.490 42.110 766.670 ;
        RECT 40.930 587.090 42.110 588.270 ;
        RECT 40.930 585.490 42.110 586.670 ;
        RECT 40.930 407.090 42.110 408.270 ;
        RECT 40.930 405.490 42.110 406.670 ;
        RECT 40.930 227.090 42.110 228.270 ;
        RECT 40.930 225.490 42.110 226.670 ;
        RECT 40.930 47.090 42.110 48.270 ;
        RECT 40.930 45.490 42.110 46.670 ;
        RECT -27.870 -21.710 -26.690 -20.530 ;
        RECT -27.870 -23.310 -26.690 -22.130 ;
        RECT 40.930 -21.710 42.110 -20.530 ;
        RECT 40.930 -23.310 42.110 -22.130 ;
        RECT 238.930 3551.210 240.110 3552.390 ;
        RECT 238.930 3549.610 240.110 3550.790 ;
        RECT 220.930 3541.810 222.110 3542.990 ;
        RECT 220.930 3540.210 222.110 3541.390 ;
        RECT 202.930 3532.410 204.110 3533.590 ;
        RECT 202.930 3530.810 204.110 3531.990 ;
        RECT 58.930 3485.090 60.110 3486.270 ;
        RECT 58.930 3483.490 60.110 3484.670 ;
        RECT 58.930 3305.090 60.110 3306.270 ;
        RECT 58.930 3303.490 60.110 3304.670 ;
        RECT 58.930 3125.090 60.110 3126.270 ;
        RECT 58.930 3123.490 60.110 3124.670 ;
        RECT 58.930 2945.090 60.110 2946.270 ;
        RECT 58.930 2943.490 60.110 2944.670 ;
        RECT 58.930 2765.090 60.110 2766.270 ;
        RECT 58.930 2763.490 60.110 2764.670 ;
        RECT 58.930 2585.090 60.110 2586.270 ;
        RECT 58.930 2583.490 60.110 2584.670 ;
        RECT 58.930 2405.090 60.110 2406.270 ;
        RECT 58.930 2403.490 60.110 2404.670 ;
        RECT 58.930 2225.090 60.110 2226.270 ;
        RECT 58.930 2223.490 60.110 2224.670 ;
        RECT 58.930 2045.090 60.110 2046.270 ;
        RECT 58.930 2043.490 60.110 2044.670 ;
        RECT 58.930 1865.090 60.110 1866.270 ;
        RECT 58.930 1863.490 60.110 1864.670 ;
        RECT 58.930 1685.090 60.110 1686.270 ;
        RECT 58.930 1683.490 60.110 1684.670 ;
        RECT 58.930 1505.090 60.110 1506.270 ;
        RECT 58.930 1503.490 60.110 1504.670 ;
        RECT 58.930 1325.090 60.110 1326.270 ;
        RECT 58.930 1323.490 60.110 1324.670 ;
        RECT 58.930 1145.090 60.110 1146.270 ;
        RECT 58.930 1143.490 60.110 1144.670 ;
        RECT 58.930 965.090 60.110 966.270 ;
        RECT 58.930 963.490 60.110 964.670 ;
        RECT 58.930 785.090 60.110 786.270 ;
        RECT 58.930 783.490 60.110 784.670 ;
        RECT 58.930 605.090 60.110 606.270 ;
        RECT 58.930 603.490 60.110 604.670 ;
        RECT 58.930 425.090 60.110 426.270 ;
        RECT 58.930 423.490 60.110 424.670 ;
        RECT 58.930 245.090 60.110 246.270 ;
        RECT 58.930 243.490 60.110 244.670 ;
        RECT 58.930 65.090 60.110 66.270 ;
        RECT 58.930 63.490 60.110 64.670 ;
        RECT -37.270 -31.110 -36.090 -29.930 ;
        RECT -37.270 -32.710 -36.090 -31.530 ;
        RECT 184.930 3523.010 186.110 3524.190 ;
        RECT 184.930 3521.410 186.110 3522.590 ;
        RECT 184.930 3431.090 186.110 3432.270 ;
        RECT 184.930 3429.490 186.110 3430.670 ;
        RECT 184.930 3251.090 186.110 3252.270 ;
        RECT 184.930 3249.490 186.110 3250.670 ;
        RECT 184.930 3071.090 186.110 3072.270 ;
        RECT 184.930 3069.490 186.110 3070.670 ;
        RECT 184.930 2891.090 186.110 2892.270 ;
        RECT 184.930 2889.490 186.110 2890.670 ;
        RECT 184.930 2711.090 186.110 2712.270 ;
        RECT 184.930 2709.490 186.110 2710.670 ;
        RECT 184.930 2531.090 186.110 2532.270 ;
        RECT 184.930 2529.490 186.110 2530.670 ;
        RECT 184.930 2351.090 186.110 2352.270 ;
        RECT 184.930 2349.490 186.110 2350.670 ;
        RECT 184.930 2171.090 186.110 2172.270 ;
        RECT 184.930 2169.490 186.110 2170.670 ;
        RECT 184.930 1991.090 186.110 1992.270 ;
        RECT 184.930 1989.490 186.110 1990.670 ;
        RECT 184.930 1811.090 186.110 1812.270 ;
        RECT 184.930 1809.490 186.110 1810.670 ;
        RECT 184.930 1631.090 186.110 1632.270 ;
        RECT 184.930 1629.490 186.110 1630.670 ;
        RECT 184.930 1451.090 186.110 1452.270 ;
        RECT 184.930 1449.490 186.110 1450.670 ;
        RECT 184.930 1271.090 186.110 1272.270 ;
        RECT 184.930 1269.490 186.110 1270.670 ;
        RECT 184.930 1091.090 186.110 1092.270 ;
        RECT 184.930 1089.490 186.110 1090.670 ;
        RECT 184.930 911.090 186.110 912.270 ;
        RECT 184.930 909.490 186.110 910.670 ;
        RECT 184.930 731.090 186.110 732.270 ;
        RECT 184.930 729.490 186.110 730.670 ;
        RECT 184.930 551.090 186.110 552.270 ;
        RECT 184.930 549.490 186.110 550.670 ;
        RECT 184.930 371.090 186.110 372.270 ;
        RECT 184.930 369.490 186.110 370.670 ;
        RECT 184.930 191.090 186.110 192.270 ;
        RECT 184.930 189.490 186.110 190.670 ;
        RECT 184.930 11.090 186.110 12.270 ;
        RECT 184.930 9.490 186.110 10.670 ;
        RECT 184.930 -2.910 186.110 -1.730 ;
        RECT 184.930 -4.510 186.110 -3.330 ;
        RECT 202.930 3449.090 204.110 3450.270 ;
        RECT 202.930 3447.490 204.110 3448.670 ;
        RECT 202.930 3269.090 204.110 3270.270 ;
        RECT 202.930 3267.490 204.110 3268.670 ;
        RECT 202.930 3089.090 204.110 3090.270 ;
        RECT 202.930 3087.490 204.110 3088.670 ;
        RECT 202.930 2909.090 204.110 2910.270 ;
        RECT 202.930 2907.490 204.110 2908.670 ;
        RECT 202.930 2729.090 204.110 2730.270 ;
        RECT 202.930 2727.490 204.110 2728.670 ;
        RECT 202.930 2549.090 204.110 2550.270 ;
        RECT 202.930 2547.490 204.110 2548.670 ;
        RECT 202.930 2369.090 204.110 2370.270 ;
        RECT 202.930 2367.490 204.110 2368.670 ;
        RECT 202.930 2189.090 204.110 2190.270 ;
        RECT 202.930 2187.490 204.110 2188.670 ;
        RECT 202.930 2009.090 204.110 2010.270 ;
        RECT 202.930 2007.490 204.110 2008.670 ;
        RECT 202.930 1829.090 204.110 1830.270 ;
        RECT 202.930 1827.490 204.110 1828.670 ;
        RECT 202.930 1649.090 204.110 1650.270 ;
        RECT 202.930 1647.490 204.110 1648.670 ;
        RECT 202.930 1469.090 204.110 1470.270 ;
        RECT 202.930 1467.490 204.110 1468.670 ;
        RECT 202.930 1289.090 204.110 1290.270 ;
        RECT 202.930 1287.490 204.110 1288.670 ;
        RECT 202.930 1109.090 204.110 1110.270 ;
        RECT 202.930 1107.490 204.110 1108.670 ;
        RECT 202.930 929.090 204.110 930.270 ;
        RECT 202.930 927.490 204.110 928.670 ;
        RECT 202.930 749.090 204.110 750.270 ;
        RECT 202.930 747.490 204.110 748.670 ;
        RECT 202.930 569.090 204.110 570.270 ;
        RECT 202.930 567.490 204.110 568.670 ;
        RECT 202.930 389.090 204.110 390.270 ;
        RECT 202.930 387.490 204.110 388.670 ;
        RECT 202.930 209.090 204.110 210.270 ;
        RECT 202.930 207.490 204.110 208.670 ;
        RECT 202.930 29.090 204.110 30.270 ;
        RECT 202.930 27.490 204.110 28.670 ;
        RECT 202.930 -12.310 204.110 -11.130 ;
        RECT 202.930 -13.910 204.110 -12.730 ;
        RECT 220.930 3467.090 222.110 3468.270 ;
        RECT 220.930 3465.490 222.110 3466.670 ;
        RECT 220.930 3287.090 222.110 3288.270 ;
        RECT 220.930 3285.490 222.110 3286.670 ;
        RECT 220.930 3107.090 222.110 3108.270 ;
        RECT 220.930 3105.490 222.110 3106.670 ;
        RECT 220.930 2927.090 222.110 2928.270 ;
        RECT 220.930 2925.490 222.110 2926.670 ;
        RECT 220.930 2747.090 222.110 2748.270 ;
        RECT 220.930 2745.490 222.110 2746.670 ;
        RECT 220.930 2567.090 222.110 2568.270 ;
        RECT 220.930 2565.490 222.110 2566.670 ;
        RECT 220.930 2387.090 222.110 2388.270 ;
        RECT 220.930 2385.490 222.110 2386.670 ;
        RECT 220.930 2207.090 222.110 2208.270 ;
        RECT 220.930 2205.490 222.110 2206.670 ;
        RECT 220.930 2027.090 222.110 2028.270 ;
        RECT 220.930 2025.490 222.110 2026.670 ;
        RECT 220.930 1847.090 222.110 1848.270 ;
        RECT 220.930 1845.490 222.110 1846.670 ;
        RECT 220.930 1667.090 222.110 1668.270 ;
        RECT 220.930 1665.490 222.110 1666.670 ;
        RECT 220.930 1487.090 222.110 1488.270 ;
        RECT 220.930 1485.490 222.110 1486.670 ;
        RECT 220.930 1307.090 222.110 1308.270 ;
        RECT 220.930 1305.490 222.110 1306.670 ;
        RECT 220.930 1127.090 222.110 1128.270 ;
        RECT 220.930 1125.490 222.110 1126.670 ;
        RECT 220.930 947.090 222.110 948.270 ;
        RECT 220.930 945.490 222.110 946.670 ;
        RECT 220.930 767.090 222.110 768.270 ;
        RECT 220.930 765.490 222.110 766.670 ;
        RECT 220.930 587.090 222.110 588.270 ;
        RECT 220.930 585.490 222.110 586.670 ;
        RECT 220.930 407.090 222.110 408.270 ;
        RECT 220.930 405.490 222.110 406.670 ;
        RECT 220.930 227.090 222.110 228.270 ;
        RECT 220.930 225.490 222.110 226.670 ;
        RECT 220.930 47.090 222.110 48.270 ;
        RECT 220.930 45.490 222.110 46.670 ;
        RECT 220.930 -21.710 222.110 -20.530 ;
        RECT 220.930 -23.310 222.110 -22.130 ;
        RECT 418.930 3551.210 420.110 3552.390 ;
        RECT 418.930 3549.610 420.110 3550.790 ;
        RECT 400.930 3541.810 402.110 3542.990 ;
        RECT 400.930 3540.210 402.110 3541.390 ;
        RECT 382.930 3532.410 384.110 3533.590 ;
        RECT 382.930 3530.810 384.110 3531.990 ;
        RECT 238.930 3485.090 240.110 3486.270 ;
        RECT 238.930 3483.490 240.110 3484.670 ;
        RECT 238.930 3305.090 240.110 3306.270 ;
        RECT 238.930 3303.490 240.110 3304.670 ;
        RECT 238.930 3125.090 240.110 3126.270 ;
        RECT 238.930 3123.490 240.110 3124.670 ;
        RECT 238.930 2945.090 240.110 2946.270 ;
        RECT 238.930 2943.490 240.110 2944.670 ;
        RECT 364.930 3523.010 366.110 3524.190 ;
        RECT 364.930 3521.410 366.110 3522.590 ;
        RECT 364.930 3431.090 366.110 3432.270 ;
        RECT 364.930 3429.490 366.110 3430.670 ;
        RECT 364.930 3251.090 366.110 3252.270 ;
        RECT 364.930 3249.490 366.110 3250.670 ;
        RECT 364.930 3071.090 366.110 3072.270 ;
        RECT 364.930 3069.490 366.110 3070.670 ;
        RECT 364.930 2891.090 366.110 2892.270 ;
        RECT 364.930 2889.490 366.110 2890.670 ;
        RECT 382.930 3449.090 384.110 3450.270 ;
        RECT 382.930 3447.490 384.110 3448.670 ;
        RECT 382.930 3269.090 384.110 3270.270 ;
        RECT 382.930 3267.490 384.110 3268.670 ;
        RECT 382.930 3089.090 384.110 3090.270 ;
        RECT 382.930 3087.490 384.110 3088.670 ;
        RECT 382.930 2909.090 384.110 2910.270 ;
        RECT 382.930 2907.490 384.110 2908.670 ;
        RECT 400.930 3467.090 402.110 3468.270 ;
        RECT 400.930 3465.490 402.110 3466.670 ;
        RECT 400.930 3287.090 402.110 3288.270 ;
        RECT 400.930 3285.490 402.110 3286.670 ;
        RECT 400.930 3107.090 402.110 3108.270 ;
        RECT 400.930 3105.490 402.110 3106.670 ;
        RECT 400.930 2927.090 402.110 2928.270 ;
        RECT 400.930 2925.490 402.110 2926.670 ;
        RECT 598.930 3551.210 600.110 3552.390 ;
        RECT 598.930 3549.610 600.110 3550.790 ;
        RECT 580.930 3541.810 582.110 3542.990 ;
        RECT 580.930 3540.210 582.110 3541.390 ;
        RECT 562.930 3532.410 564.110 3533.590 ;
        RECT 562.930 3530.810 564.110 3531.990 ;
        RECT 418.930 3485.090 420.110 3486.270 ;
        RECT 418.930 3483.490 420.110 3484.670 ;
        RECT 418.930 3305.090 420.110 3306.270 ;
        RECT 418.930 3303.490 420.110 3304.670 ;
        RECT 418.930 3125.090 420.110 3126.270 ;
        RECT 418.930 3123.490 420.110 3124.670 ;
        RECT 418.930 2945.090 420.110 2946.270 ;
        RECT 418.930 2943.490 420.110 2944.670 ;
        RECT 544.930 3523.010 546.110 3524.190 ;
        RECT 544.930 3521.410 546.110 3522.590 ;
        RECT 544.930 3431.090 546.110 3432.270 ;
        RECT 544.930 3429.490 546.110 3430.670 ;
        RECT 544.930 3251.090 546.110 3252.270 ;
        RECT 544.930 3249.490 546.110 3250.670 ;
        RECT 544.930 3071.090 546.110 3072.270 ;
        RECT 544.930 3069.490 546.110 3070.670 ;
        RECT 544.930 2891.090 546.110 2892.270 ;
        RECT 544.930 2889.490 546.110 2890.670 ;
        RECT 562.930 3449.090 564.110 3450.270 ;
        RECT 562.930 3447.490 564.110 3448.670 ;
        RECT 562.930 3269.090 564.110 3270.270 ;
        RECT 562.930 3267.490 564.110 3268.670 ;
        RECT 562.930 3089.090 564.110 3090.270 ;
        RECT 562.930 3087.490 564.110 3088.670 ;
        RECT 562.930 2909.090 564.110 2910.270 ;
        RECT 562.930 2907.490 564.110 2908.670 ;
        RECT 580.930 3467.090 582.110 3468.270 ;
        RECT 580.930 3465.490 582.110 3466.670 ;
        RECT 580.930 3287.090 582.110 3288.270 ;
        RECT 580.930 3285.490 582.110 3286.670 ;
        RECT 580.930 3107.090 582.110 3108.270 ;
        RECT 580.930 3105.490 582.110 3106.670 ;
        RECT 580.930 2927.090 582.110 2928.270 ;
        RECT 580.930 2925.490 582.110 2926.670 ;
        RECT 778.930 3551.210 780.110 3552.390 ;
        RECT 778.930 3549.610 780.110 3550.790 ;
        RECT 760.930 3541.810 762.110 3542.990 ;
        RECT 760.930 3540.210 762.110 3541.390 ;
        RECT 742.930 3532.410 744.110 3533.590 ;
        RECT 742.930 3530.810 744.110 3531.990 ;
        RECT 598.930 3485.090 600.110 3486.270 ;
        RECT 598.930 3483.490 600.110 3484.670 ;
        RECT 598.930 3305.090 600.110 3306.270 ;
        RECT 598.930 3303.490 600.110 3304.670 ;
        RECT 598.930 3125.090 600.110 3126.270 ;
        RECT 598.930 3123.490 600.110 3124.670 ;
        RECT 598.930 2945.090 600.110 2946.270 ;
        RECT 598.930 2943.490 600.110 2944.670 ;
        RECT 724.930 3523.010 726.110 3524.190 ;
        RECT 724.930 3521.410 726.110 3522.590 ;
        RECT 724.930 3431.090 726.110 3432.270 ;
        RECT 724.930 3429.490 726.110 3430.670 ;
        RECT 724.930 3251.090 726.110 3252.270 ;
        RECT 724.930 3249.490 726.110 3250.670 ;
        RECT 724.930 3071.090 726.110 3072.270 ;
        RECT 724.930 3069.490 726.110 3070.670 ;
        RECT 724.930 2891.090 726.110 2892.270 ;
        RECT 724.930 2889.490 726.110 2890.670 ;
        RECT 238.930 2765.090 240.110 2766.270 ;
        RECT 238.930 2763.490 240.110 2764.670 ;
        RECT 238.930 2585.090 240.110 2586.270 ;
        RECT 238.930 2583.490 240.110 2584.670 ;
        RECT 238.930 2405.090 240.110 2406.270 ;
        RECT 238.930 2403.490 240.110 2404.670 ;
        RECT 682.680 2729.090 683.860 2730.270 ;
        RECT 682.680 2727.490 683.860 2728.670 ;
        RECT 682.680 2711.090 683.860 2712.270 ;
        RECT 682.680 2709.490 683.860 2710.670 ;
        RECT 682.680 2585.090 683.860 2586.270 ;
        RECT 682.680 2583.490 683.860 2584.670 ;
        RECT 682.680 2567.090 683.860 2568.270 ;
        RECT 682.680 2565.490 683.860 2566.670 ;
        RECT 682.680 2549.090 683.860 2550.270 ;
        RECT 682.680 2547.490 683.860 2548.670 ;
        RECT 682.680 2531.090 683.860 2532.270 ;
        RECT 682.680 2529.490 683.860 2530.670 ;
        RECT 682.680 2405.090 683.860 2406.270 ;
        RECT 682.680 2403.490 683.860 2404.670 ;
        RECT 682.680 2387.090 683.860 2388.270 ;
        RECT 682.680 2385.490 683.860 2386.670 ;
        RECT 682.680 2369.090 683.860 2370.270 ;
        RECT 682.680 2367.490 683.860 2368.670 ;
        RECT 682.680 2351.090 683.860 2352.270 ;
        RECT 682.680 2349.490 683.860 2350.670 ;
        RECT 724.930 2711.090 726.110 2712.270 ;
        RECT 724.930 2709.490 726.110 2710.670 ;
        RECT 724.930 2531.090 726.110 2532.270 ;
        RECT 724.930 2529.490 726.110 2530.670 ;
        RECT 724.930 2351.090 726.110 2352.270 ;
        RECT 724.930 2349.490 726.110 2350.670 ;
        RECT 238.930 2225.090 240.110 2226.270 ;
        RECT 238.930 2223.490 240.110 2224.670 ;
        RECT 418.930 2225.090 420.110 2226.270 ;
        RECT 418.930 2223.490 420.110 2224.670 ;
        RECT 598.930 2225.090 600.110 2226.270 ;
        RECT 598.930 2223.490 600.110 2224.670 ;
        RECT 742.930 3449.090 744.110 3450.270 ;
        RECT 742.930 3447.490 744.110 3448.670 ;
        RECT 742.930 3269.090 744.110 3270.270 ;
        RECT 742.930 3267.490 744.110 3268.670 ;
        RECT 742.930 3089.090 744.110 3090.270 ;
        RECT 742.930 3087.490 744.110 3088.670 ;
        RECT 742.930 2909.090 744.110 2910.270 ;
        RECT 742.930 2907.490 744.110 2908.670 ;
        RECT 742.930 2729.090 744.110 2730.270 ;
        RECT 742.930 2727.490 744.110 2728.670 ;
        RECT 742.930 2549.090 744.110 2550.270 ;
        RECT 742.930 2547.490 744.110 2548.670 ;
        RECT 742.930 2369.090 744.110 2370.270 ;
        RECT 742.930 2367.490 744.110 2368.670 ;
        RECT 760.930 3467.090 762.110 3468.270 ;
        RECT 760.930 3465.490 762.110 3466.670 ;
        RECT 760.930 3287.090 762.110 3288.270 ;
        RECT 760.930 3285.490 762.110 3286.670 ;
        RECT 760.930 3107.090 762.110 3108.270 ;
        RECT 760.930 3105.490 762.110 3106.670 ;
        RECT 760.930 2927.090 762.110 2928.270 ;
        RECT 760.930 2925.490 762.110 2926.670 ;
        RECT 760.930 2747.090 762.110 2748.270 ;
        RECT 760.930 2745.490 762.110 2746.670 ;
        RECT 760.930 2567.090 762.110 2568.270 ;
        RECT 760.930 2565.490 762.110 2566.670 ;
        RECT 760.930 2387.090 762.110 2388.270 ;
        RECT 760.930 2385.490 762.110 2386.670 ;
        RECT 958.930 3551.210 960.110 3552.390 ;
        RECT 958.930 3549.610 960.110 3550.790 ;
        RECT 940.930 3541.810 942.110 3542.990 ;
        RECT 940.930 3540.210 942.110 3541.390 ;
        RECT 922.930 3532.410 924.110 3533.590 ;
        RECT 922.930 3530.810 924.110 3531.990 ;
        RECT 778.930 3485.090 780.110 3486.270 ;
        RECT 778.930 3483.490 780.110 3484.670 ;
        RECT 778.930 3305.090 780.110 3306.270 ;
        RECT 778.930 3303.490 780.110 3304.670 ;
        RECT 778.930 3125.090 780.110 3126.270 ;
        RECT 778.930 3123.490 780.110 3124.670 ;
        RECT 778.930 2945.090 780.110 2946.270 ;
        RECT 778.930 2943.490 780.110 2944.670 ;
        RECT 778.930 2765.090 780.110 2766.270 ;
        RECT 778.930 2763.490 780.110 2764.670 ;
        RECT 778.930 2585.090 780.110 2586.270 ;
        RECT 778.930 2583.490 780.110 2584.670 ;
        RECT 778.930 2405.090 780.110 2406.270 ;
        RECT 778.930 2403.490 780.110 2404.670 ;
        RECT 778.930 2225.090 780.110 2226.270 ;
        RECT 778.930 2223.490 780.110 2224.670 ;
        RECT 904.930 3523.010 906.110 3524.190 ;
        RECT 904.930 3521.410 906.110 3522.590 ;
        RECT 904.930 3431.090 906.110 3432.270 ;
        RECT 904.930 3429.490 906.110 3430.670 ;
        RECT 904.930 3251.090 906.110 3252.270 ;
        RECT 904.930 3249.490 906.110 3250.670 ;
        RECT 904.930 3071.090 906.110 3072.270 ;
        RECT 904.930 3069.490 906.110 3070.670 ;
        RECT 904.930 2891.090 906.110 2892.270 ;
        RECT 904.930 2889.490 906.110 2890.670 ;
        RECT 904.930 2711.090 906.110 2712.270 ;
        RECT 904.930 2709.490 906.110 2710.670 ;
        RECT 904.930 2531.090 906.110 2532.270 ;
        RECT 904.930 2529.490 906.110 2530.670 ;
        RECT 904.930 2351.090 906.110 2352.270 ;
        RECT 904.930 2349.490 906.110 2350.670 ;
        RECT 922.930 3449.090 924.110 3450.270 ;
        RECT 922.930 3447.490 924.110 3448.670 ;
        RECT 922.930 3269.090 924.110 3270.270 ;
        RECT 922.930 3267.490 924.110 3268.670 ;
        RECT 922.930 3089.090 924.110 3090.270 ;
        RECT 922.930 3087.490 924.110 3088.670 ;
        RECT 922.930 2909.090 924.110 2910.270 ;
        RECT 922.930 2907.490 924.110 2908.670 ;
        RECT 940.930 3467.090 942.110 3468.270 ;
        RECT 940.930 3465.490 942.110 3466.670 ;
        RECT 940.930 3287.090 942.110 3288.270 ;
        RECT 940.930 3285.490 942.110 3286.670 ;
        RECT 940.930 3107.090 942.110 3108.270 ;
        RECT 940.930 3105.490 942.110 3106.670 ;
        RECT 940.930 2927.090 942.110 2928.270 ;
        RECT 940.930 2925.490 942.110 2926.670 ;
        RECT 1138.930 3551.210 1140.110 3552.390 ;
        RECT 1138.930 3549.610 1140.110 3550.790 ;
        RECT 1120.930 3541.810 1122.110 3542.990 ;
        RECT 1120.930 3540.210 1122.110 3541.390 ;
        RECT 1102.930 3532.410 1104.110 3533.590 ;
        RECT 1102.930 3530.810 1104.110 3531.990 ;
        RECT 958.930 3485.090 960.110 3486.270 ;
        RECT 958.930 3483.490 960.110 3484.670 ;
        RECT 958.930 3305.090 960.110 3306.270 ;
        RECT 958.930 3303.490 960.110 3304.670 ;
        RECT 958.930 3125.090 960.110 3126.270 ;
        RECT 958.930 3123.490 960.110 3124.670 ;
        RECT 958.930 2945.090 960.110 2946.270 ;
        RECT 958.930 2943.490 960.110 2944.670 ;
        RECT 1084.930 3523.010 1086.110 3524.190 ;
        RECT 1084.930 3521.410 1086.110 3522.590 ;
        RECT 1084.930 3431.090 1086.110 3432.270 ;
        RECT 1084.930 3429.490 1086.110 3430.670 ;
        RECT 1084.930 3251.090 1086.110 3252.270 ;
        RECT 1084.930 3249.490 1086.110 3250.670 ;
        RECT 1084.930 3071.090 1086.110 3072.270 ;
        RECT 1084.930 3069.490 1086.110 3070.670 ;
        RECT 1084.930 2891.090 1086.110 2892.270 ;
        RECT 1084.930 2889.490 1086.110 2890.670 ;
        RECT 1102.930 3449.090 1104.110 3450.270 ;
        RECT 1102.930 3447.490 1104.110 3448.670 ;
        RECT 1102.930 3269.090 1104.110 3270.270 ;
        RECT 1102.930 3267.490 1104.110 3268.670 ;
        RECT 1102.930 3089.090 1104.110 3090.270 ;
        RECT 1102.930 3087.490 1104.110 3088.670 ;
        RECT 1102.930 2909.090 1104.110 2910.270 ;
        RECT 1102.930 2907.490 1104.110 2908.670 ;
        RECT 1120.930 3467.090 1122.110 3468.270 ;
        RECT 1120.930 3465.490 1122.110 3466.670 ;
        RECT 1120.930 3287.090 1122.110 3288.270 ;
        RECT 1120.930 3285.490 1122.110 3286.670 ;
        RECT 1120.930 3107.090 1122.110 3108.270 ;
        RECT 1120.930 3105.490 1122.110 3106.670 ;
        RECT 1120.930 2927.090 1122.110 2928.270 ;
        RECT 1120.930 2925.490 1122.110 2926.670 ;
        RECT 1318.930 3551.210 1320.110 3552.390 ;
        RECT 1318.930 3549.610 1320.110 3550.790 ;
        RECT 1300.930 3541.810 1302.110 3542.990 ;
        RECT 1300.930 3540.210 1302.110 3541.390 ;
        RECT 1282.930 3532.410 1284.110 3533.590 ;
        RECT 1282.930 3530.810 1284.110 3531.990 ;
        RECT 1138.930 3485.090 1140.110 3486.270 ;
        RECT 1138.930 3483.490 1140.110 3484.670 ;
        RECT 1138.930 3305.090 1140.110 3306.270 ;
        RECT 1138.930 3303.490 1140.110 3304.670 ;
        RECT 1138.930 3125.090 1140.110 3126.270 ;
        RECT 1138.930 3123.490 1140.110 3124.670 ;
        RECT 1138.930 2945.090 1140.110 2946.270 ;
        RECT 1138.930 2943.490 1140.110 2944.670 ;
        RECT 1264.930 3523.010 1266.110 3524.190 ;
        RECT 1264.930 3521.410 1266.110 3522.590 ;
        RECT 1264.930 3431.090 1266.110 3432.270 ;
        RECT 1264.930 3429.490 1266.110 3430.670 ;
        RECT 1264.930 3251.090 1266.110 3252.270 ;
        RECT 1264.930 3249.490 1266.110 3250.670 ;
        RECT 1264.930 3071.090 1266.110 3072.270 ;
        RECT 1264.930 3069.490 1266.110 3070.670 ;
        RECT 1264.930 2891.090 1266.110 2892.270 ;
        RECT 1264.930 2889.490 1266.110 2890.670 ;
        RECT 1282.930 3449.090 1284.110 3450.270 ;
        RECT 1282.930 3447.490 1284.110 3448.670 ;
        RECT 1282.930 3269.090 1284.110 3270.270 ;
        RECT 1282.930 3267.490 1284.110 3268.670 ;
        RECT 1282.930 3089.090 1284.110 3090.270 ;
        RECT 1282.930 3087.490 1284.110 3088.670 ;
        RECT 1282.930 2909.090 1284.110 2910.270 ;
        RECT 1282.930 2907.490 1284.110 2908.670 ;
        RECT 1300.930 3467.090 1302.110 3468.270 ;
        RECT 1300.930 3465.490 1302.110 3466.670 ;
        RECT 1300.930 3287.090 1302.110 3288.270 ;
        RECT 1300.930 3285.490 1302.110 3286.670 ;
        RECT 1300.930 3107.090 1302.110 3108.270 ;
        RECT 1300.930 3105.490 1302.110 3106.670 ;
        RECT 1300.930 2927.090 1302.110 2928.270 ;
        RECT 1300.930 2925.490 1302.110 2926.670 ;
        RECT 1498.930 3551.210 1500.110 3552.390 ;
        RECT 1498.930 3549.610 1500.110 3550.790 ;
        RECT 1480.930 3541.810 1482.110 3542.990 ;
        RECT 1480.930 3540.210 1482.110 3541.390 ;
        RECT 1462.930 3532.410 1464.110 3533.590 ;
        RECT 1462.930 3530.810 1464.110 3531.990 ;
        RECT 1318.930 3485.090 1320.110 3486.270 ;
        RECT 1318.930 3483.490 1320.110 3484.670 ;
        RECT 1318.930 3305.090 1320.110 3306.270 ;
        RECT 1318.930 3303.490 1320.110 3304.670 ;
        RECT 1318.930 3125.090 1320.110 3126.270 ;
        RECT 1318.930 3123.490 1320.110 3124.670 ;
        RECT 1318.930 2945.090 1320.110 2946.270 ;
        RECT 1318.930 2943.490 1320.110 2944.670 ;
        RECT 1444.930 3523.010 1446.110 3524.190 ;
        RECT 1444.930 3521.410 1446.110 3522.590 ;
        RECT 1444.930 3431.090 1446.110 3432.270 ;
        RECT 1444.930 3429.490 1446.110 3430.670 ;
        RECT 1444.930 3251.090 1446.110 3252.270 ;
        RECT 1444.930 3249.490 1446.110 3250.670 ;
        RECT 1444.930 3071.090 1446.110 3072.270 ;
        RECT 1444.930 3069.490 1446.110 3070.670 ;
        RECT 1444.930 2891.090 1446.110 2892.270 ;
        RECT 1444.930 2889.490 1446.110 2890.670 ;
        RECT 922.930 2729.090 924.110 2730.270 ;
        RECT 922.930 2727.490 924.110 2728.670 ;
        RECT 922.930 2549.090 924.110 2550.270 ;
        RECT 922.930 2547.490 924.110 2548.670 ;
        RECT 922.930 2369.090 924.110 2370.270 ;
        RECT 922.930 2367.490 924.110 2368.670 ;
        RECT 1332.680 2729.090 1333.860 2730.270 ;
        RECT 1332.680 2727.490 1333.860 2728.670 ;
        RECT 1332.680 2711.090 1333.860 2712.270 ;
        RECT 1332.680 2709.490 1333.860 2710.670 ;
        RECT 1332.680 2585.090 1333.860 2586.270 ;
        RECT 1332.680 2583.490 1333.860 2584.670 ;
        RECT 1332.680 2567.090 1333.860 2568.270 ;
        RECT 1332.680 2565.490 1333.860 2566.670 ;
        RECT 1332.680 2549.090 1333.860 2550.270 ;
        RECT 1332.680 2547.490 1333.860 2548.670 ;
        RECT 1332.680 2531.090 1333.860 2532.270 ;
        RECT 1332.680 2529.490 1333.860 2530.670 ;
        RECT 1332.680 2405.090 1333.860 2406.270 ;
        RECT 1332.680 2403.490 1333.860 2404.670 ;
        RECT 1332.680 2387.090 1333.860 2388.270 ;
        RECT 1332.680 2385.490 1333.860 2386.670 ;
        RECT 1332.680 2369.090 1333.860 2370.270 ;
        RECT 1332.680 2367.490 1333.860 2368.670 ;
        RECT 1332.680 2351.090 1333.860 2352.270 ;
        RECT 1332.680 2349.490 1333.860 2350.670 ;
        RECT 1444.930 2711.090 1446.110 2712.270 ;
        RECT 1444.930 2709.490 1446.110 2710.670 ;
        RECT 1444.930 2531.090 1446.110 2532.270 ;
        RECT 1444.930 2529.490 1446.110 2530.670 ;
        RECT 1444.930 2351.090 1446.110 2352.270 ;
        RECT 1444.930 2349.490 1446.110 2350.670 ;
        RECT 958.930 2225.090 960.110 2226.270 ;
        RECT 958.930 2223.490 960.110 2224.670 ;
        RECT 1138.930 2225.090 1140.110 2226.270 ;
        RECT 1138.930 2223.490 1140.110 2224.670 ;
        RECT 1318.930 2225.090 1320.110 2226.270 ;
        RECT 1318.930 2223.490 1320.110 2224.670 ;
        RECT 1462.930 3449.090 1464.110 3450.270 ;
        RECT 1462.930 3447.490 1464.110 3448.670 ;
        RECT 1462.930 3269.090 1464.110 3270.270 ;
        RECT 1462.930 3267.490 1464.110 3268.670 ;
        RECT 1462.930 3089.090 1464.110 3090.270 ;
        RECT 1462.930 3087.490 1464.110 3088.670 ;
        RECT 1462.930 2909.090 1464.110 2910.270 ;
        RECT 1462.930 2907.490 1464.110 2908.670 ;
        RECT 1462.930 2729.090 1464.110 2730.270 ;
        RECT 1462.930 2727.490 1464.110 2728.670 ;
        RECT 1462.930 2549.090 1464.110 2550.270 ;
        RECT 1462.930 2547.490 1464.110 2548.670 ;
        RECT 1462.930 2369.090 1464.110 2370.270 ;
        RECT 1462.930 2367.490 1464.110 2368.670 ;
        RECT 1480.930 3467.090 1482.110 3468.270 ;
        RECT 1480.930 3465.490 1482.110 3466.670 ;
        RECT 1480.930 3287.090 1482.110 3288.270 ;
        RECT 1480.930 3285.490 1482.110 3286.670 ;
        RECT 1480.930 3107.090 1482.110 3108.270 ;
        RECT 1480.930 3105.490 1482.110 3106.670 ;
        RECT 1480.930 2927.090 1482.110 2928.270 ;
        RECT 1480.930 2925.490 1482.110 2926.670 ;
        RECT 1480.930 2747.090 1482.110 2748.270 ;
        RECT 1480.930 2745.490 1482.110 2746.670 ;
        RECT 1480.930 2567.090 1482.110 2568.270 ;
        RECT 1480.930 2565.490 1482.110 2566.670 ;
        RECT 1480.930 2387.090 1482.110 2388.270 ;
        RECT 1480.930 2385.490 1482.110 2386.670 ;
        RECT 1678.930 3551.210 1680.110 3552.390 ;
        RECT 1678.930 3549.610 1680.110 3550.790 ;
        RECT 1660.930 3541.810 1662.110 3542.990 ;
        RECT 1660.930 3540.210 1662.110 3541.390 ;
        RECT 1642.930 3532.410 1644.110 3533.590 ;
        RECT 1642.930 3530.810 1644.110 3531.990 ;
        RECT 1498.930 3485.090 1500.110 3486.270 ;
        RECT 1498.930 3483.490 1500.110 3484.670 ;
        RECT 1498.930 3305.090 1500.110 3306.270 ;
        RECT 1498.930 3303.490 1500.110 3304.670 ;
        RECT 1498.930 3125.090 1500.110 3126.270 ;
        RECT 1498.930 3123.490 1500.110 3124.670 ;
        RECT 1498.930 2945.090 1500.110 2946.270 ;
        RECT 1498.930 2943.490 1500.110 2944.670 ;
        RECT 1624.930 3523.010 1626.110 3524.190 ;
        RECT 1624.930 3521.410 1626.110 3522.590 ;
        RECT 1624.930 3431.090 1626.110 3432.270 ;
        RECT 1624.930 3429.490 1626.110 3430.670 ;
        RECT 1624.930 3251.090 1626.110 3252.270 ;
        RECT 1624.930 3249.490 1626.110 3250.670 ;
        RECT 1624.930 3071.090 1626.110 3072.270 ;
        RECT 1624.930 3069.490 1626.110 3070.670 ;
        RECT 1624.930 2891.090 1626.110 2892.270 ;
        RECT 1624.930 2889.490 1626.110 2890.670 ;
        RECT 1642.930 3449.090 1644.110 3450.270 ;
        RECT 1642.930 3447.490 1644.110 3448.670 ;
        RECT 1642.930 3269.090 1644.110 3270.270 ;
        RECT 1642.930 3267.490 1644.110 3268.670 ;
        RECT 1642.930 3089.090 1644.110 3090.270 ;
        RECT 1642.930 3087.490 1644.110 3088.670 ;
        RECT 1642.930 2909.090 1644.110 2910.270 ;
        RECT 1642.930 2907.490 1644.110 2908.670 ;
        RECT 1660.930 3467.090 1662.110 3468.270 ;
        RECT 1660.930 3465.490 1662.110 3466.670 ;
        RECT 1660.930 3287.090 1662.110 3288.270 ;
        RECT 1660.930 3285.490 1662.110 3286.670 ;
        RECT 1660.930 3107.090 1662.110 3108.270 ;
        RECT 1660.930 3105.490 1662.110 3106.670 ;
        RECT 1660.930 2927.090 1662.110 2928.270 ;
        RECT 1660.930 2925.490 1662.110 2926.670 ;
        RECT 1858.930 3551.210 1860.110 3552.390 ;
        RECT 1858.930 3549.610 1860.110 3550.790 ;
        RECT 1840.930 3541.810 1842.110 3542.990 ;
        RECT 1840.930 3540.210 1842.110 3541.390 ;
        RECT 1822.930 3532.410 1824.110 3533.590 ;
        RECT 1822.930 3530.810 1824.110 3531.990 ;
        RECT 1678.930 3485.090 1680.110 3486.270 ;
        RECT 1678.930 3483.490 1680.110 3484.670 ;
        RECT 1678.930 3305.090 1680.110 3306.270 ;
        RECT 1678.930 3303.490 1680.110 3304.670 ;
        RECT 1678.930 3125.090 1680.110 3126.270 ;
        RECT 1678.930 3123.490 1680.110 3124.670 ;
        RECT 1678.930 2945.090 1680.110 2946.270 ;
        RECT 1678.930 2943.490 1680.110 2944.670 ;
        RECT 1804.930 3523.010 1806.110 3524.190 ;
        RECT 1804.930 3521.410 1806.110 3522.590 ;
        RECT 1804.930 3431.090 1806.110 3432.270 ;
        RECT 1804.930 3429.490 1806.110 3430.670 ;
        RECT 1804.930 3251.090 1806.110 3252.270 ;
        RECT 1804.930 3249.490 1806.110 3250.670 ;
        RECT 1804.930 3071.090 1806.110 3072.270 ;
        RECT 1804.930 3069.490 1806.110 3070.670 ;
        RECT 1804.930 2891.090 1806.110 2892.270 ;
        RECT 1804.930 2889.490 1806.110 2890.670 ;
        RECT 1822.930 3449.090 1824.110 3450.270 ;
        RECT 1822.930 3447.490 1824.110 3448.670 ;
        RECT 1822.930 3269.090 1824.110 3270.270 ;
        RECT 1822.930 3267.490 1824.110 3268.670 ;
        RECT 1822.930 3089.090 1824.110 3090.270 ;
        RECT 1822.930 3087.490 1824.110 3088.670 ;
        RECT 1822.930 2909.090 1824.110 2910.270 ;
        RECT 1822.930 2907.490 1824.110 2908.670 ;
        RECT 1840.930 3467.090 1842.110 3468.270 ;
        RECT 1840.930 3465.490 1842.110 3466.670 ;
        RECT 1840.930 3287.090 1842.110 3288.270 ;
        RECT 1840.930 3285.490 1842.110 3286.670 ;
        RECT 1840.930 3107.090 1842.110 3108.270 ;
        RECT 1840.930 3105.490 1842.110 3106.670 ;
        RECT 1840.930 2927.090 1842.110 2928.270 ;
        RECT 1840.930 2925.490 1842.110 2926.670 ;
        RECT 2038.930 3551.210 2040.110 3552.390 ;
        RECT 2038.930 3549.610 2040.110 3550.790 ;
        RECT 2020.930 3541.810 2022.110 3542.990 ;
        RECT 2020.930 3540.210 2022.110 3541.390 ;
        RECT 2002.930 3532.410 2004.110 3533.590 ;
        RECT 2002.930 3530.810 2004.110 3531.990 ;
        RECT 1858.930 3485.090 1860.110 3486.270 ;
        RECT 1858.930 3483.490 1860.110 3484.670 ;
        RECT 1858.930 3305.090 1860.110 3306.270 ;
        RECT 1858.930 3303.490 1860.110 3304.670 ;
        RECT 1858.930 3125.090 1860.110 3126.270 ;
        RECT 1858.930 3123.490 1860.110 3124.670 ;
        RECT 1858.930 2945.090 1860.110 2946.270 ;
        RECT 1858.930 2943.490 1860.110 2944.670 ;
        RECT 1984.930 3523.010 1986.110 3524.190 ;
        RECT 1984.930 3521.410 1986.110 3522.590 ;
        RECT 1984.930 3431.090 1986.110 3432.270 ;
        RECT 1984.930 3429.490 1986.110 3430.670 ;
        RECT 1984.930 3251.090 1986.110 3252.270 ;
        RECT 1984.930 3249.490 1986.110 3250.670 ;
        RECT 1984.930 3071.090 1986.110 3072.270 ;
        RECT 1984.930 3069.490 1986.110 3070.670 ;
        RECT 1984.930 2891.090 1986.110 2892.270 ;
        RECT 1984.930 2889.490 1986.110 2890.670 ;
        RECT 1498.930 2765.090 1500.110 2766.270 ;
        RECT 1498.930 2763.490 1500.110 2764.670 ;
        RECT 1498.930 2585.090 1500.110 2586.270 ;
        RECT 1498.930 2583.490 1500.110 2584.670 ;
        RECT 1498.930 2405.090 1500.110 2406.270 ;
        RECT 1498.930 2403.490 1500.110 2404.670 ;
        RECT 1932.680 2729.090 1933.860 2730.270 ;
        RECT 1932.680 2727.490 1933.860 2728.670 ;
        RECT 1932.680 2711.090 1933.860 2712.270 ;
        RECT 1932.680 2709.490 1933.860 2710.670 ;
        RECT 1932.680 2585.090 1933.860 2586.270 ;
        RECT 1932.680 2583.490 1933.860 2584.670 ;
        RECT 1932.680 2567.090 1933.860 2568.270 ;
        RECT 1932.680 2565.490 1933.860 2566.670 ;
        RECT 1932.680 2549.090 1933.860 2550.270 ;
        RECT 1932.680 2547.490 1933.860 2548.670 ;
        RECT 1932.680 2531.090 1933.860 2532.270 ;
        RECT 1932.680 2529.490 1933.860 2530.670 ;
        RECT 1932.680 2405.090 1933.860 2406.270 ;
        RECT 1932.680 2403.490 1933.860 2404.670 ;
        RECT 1932.680 2387.090 1933.860 2388.270 ;
        RECT 1932.680 2385.490 1933.860 2386.670 ;
        RECT 1932.680 2369.090 1933.860 2370.270 ;
        RECT 1932.680 2367.490 1933.860 2368.670 ;
        RECT 1932.680 2351.090 1933.860 2352.270 ;
        RECT 1932.680 2349.490 1933.860 2350.670 ;
        RECT 1984.930 2711.090 1986.110 2712.270 ;
        RECT 1984.930 2709.490 1986.110 2710.670 ;
        RECT 1984.930 2531.090 1986.110 2532.270 ;
        RECT 1984.930 2529.490 1986.110 2530.670 ;
        RECT 1984.930 2351.090 1986.110 2352.270 ;
        RECT 1984.930 2349.490 1986.110 2350.670 ;
        RECT 1498.930 2225.090 1500.110 2226.270 ;
        RECT 1498.930 2223.490 1500.110 2224.670 ;
        RECT 238.930 2045.090 240.110 2046.270 ;
        RECT 238.930 2043.490 240.110 2044.670 ;
        RECT 238.930 1865.090 240.110 1866.270 ;
        RECT 238.930 1863.490 240.110 1864.670 ;
        RECT 238.930 1685.090 240.110 1686.270 ;
        RECT 238.930 1683.490 240.110 1684.670 ;
        RECT 238.930 1505.090 240.110 1506.270 ;
        RECT 238.930 1503.490 240.110 1504.670 ;
        RECT 238.930 1325.090 240.110 1326.270 ;
        RECT 238.930 1323.490 240.110 1324.670 ;
        RECT 238.930 1145.090 240.110 1146.270 ;
        RECT 238.930 1143.490 240.110 1144.670 ;
        RECT 321.250 2171.090 322.430 2172.270 ;
        RECT 321.250 2169.490 322.430 2170.670 ;
        RECT 321.250 2045.090 322.430 2046.270 ;
        RECT 321.250 2043.490 322.430 2044.670 ;
        RECT 321.250 2027.090 322.430 2028.270 ;
        RECT 321.250 2025.490 322.430 2026.670 ;
        RECT 321.250 2009.090 322.430 2010.270 ;
        RECT 321.250 2007.490 322.430 2008.670 ;
        RECT 321.250 1991.090 322.430 1992.270 ;
        RECT 321.250 1989.490 322.430 1990.670 ;
        RECT 321.250 1865.090 322.430 1866.270 ;
        RECT 321.250 1863.490 322.430 1864.670 ;
        RECT 321.250 1847.090 322.430 1848.270 ;
        RECT 321.250 1845.490 322.430 1846.670 ;
        RECT 321.250 1829.090 322.430 1830.270 ;
        RECT 321.250 1827.490 322.430 1828.670 ;
        RECT 321.250 1811.090 322.430 1812.270 ;
        RECT 321.250 1809.490 322.430 1810.670 ;
        RECT 321.250 1685.090 322.430 1686.270 ;
        RECT 321.250 1683.490 322.430 1684.670 ;
        RECT 321.250 1667.090 322.430 1668.270 ;
        RECT 321.250 1665.490 322.430 1666.670 ;
        RECT 321.250 1649.090 322.430 1650.270 ;
        RECT 321.250 1647.490 322.430 1648.670 ;
        RECT 321.250 1631.090 322.430 1632.270 ;
        RECT 321.250 1629.490 322.430 1630.670 ;
        RECT 321.250 1505.090 322.430 1506.270 ;
        RECT 321.250 1503.490 322.430 1504.670 ;
        RECT 321.250 1487.090 322.430 1488.270 ;
        RECT 321.250 1485.490 322.430 1486.670 ;
        RECT 321.250 1469.090 322.430 1470.270 ;
        RECT 321.250 1467.490 322.430 1468.670 ;
        RECT 321.250 1451.090 322.430 1452.270 ;
        RECT 321.250 1449.490 322.430 1450.670 ;
        RECT 321.250 1325.090 322.430 1326.270 ;
        RECT 321.250 1323.490 322.430 1324.670 ;
        RECT 321.250 1307.090 322.430 1308.270 ;
        RECT 321.250 1305.490 322.430 1306.670 ;
        RECT 321.250 1289.090 322.430 1290.270 ;
        RECT 321.250 1287.490 322.430 1288.670 ;
        RECT 321.250 1271.090 322.430 1272.270 ;
        RECT 321.250 1269.490 322.430 1270.670 ;
        RECT 321.250 1145.090 322.430 1146.270 ;
        RECT 321.250 1143.490 322.430 1144.670 ;
        RECT 321.250 1127.090 322.430 1128.270 ;
        RECT 321.250 1125.490 322.430 1126.670 ;
        RECT 321.250 1109.090 322.430 1110.270 ;
        RECT 321.250 1107.490 322.430 1108.670 ;
        RECT 321.250 1091.090 322.430 1092.270 ;
        RECT 321.250 1089.490 322.430 1090.670 ;
        RECT 1624.930 2171.090 1626.110 2172.270 ;
        RECT 1624.930 2169.490 1626.110 2170.670 ;
        RECT 1624.930 1991.090 1626.110 1992.270 ;
        RECT 1624.930 1989.490 1626.110 1990.670 ;
        RECT 1624.930 1811.090 1626.110 1812.270 ;
        RECT 1624.930 1809.490 1626.110 1810.670 ;
        RECT 1624.930 1631.090 1626.110 1632.270 ;
        RECT 1624.930 1629.490 1626.110 1630.670 ;
        RECT 1624.930 1451.090 1626.110 1452.270 ;
        RECT 1624.930 1449.490 1626.110 1450.670 ;
        RECT 1624.930 1271.090 1626.110 1272.270 ;
        RECT 1624.930 1269.490 1626.110 1270.670 ;
        RECT 1624.930 1091.090 1626.110 1092.270 ;
        RECT 1624.930 1089.490 1626.110 1090.670 ;
        RECT 238.930 965.090 240.110 966.270 ;
        RECT 238.930 963.490 240.110 964.670 ;
        RECT 238.930 785.090 240.110 786.270 ;
        RECT 238.930 783.490 240.110 784.670 ;
        RECT 238.930 605.090 240.110 606.270 ;
        RECT 238.930 603.490 240.110 604.670 ;
        RECT 238.930 425.090 240.110 426.270 ;
        RECT 238.930 423.490 240.110 424.670 ;
        RECT 238.930 245.090 240.110 246.270 ;
        RECT 238.930 243.490 240.110 244.670 ;
        RECT 238.930 65.090 240.110 66.270 ;
        RECT 238.930 63.490 240.110 64.670 ;
        RECT 58.930 -31.110 60.110 -29.930 ;
        RECT 58.930 -32.710 60.110 -31.530 ;
        RECT 364.930 911.090 366.110 912.270 ;
        RECT 364.930 909.490 366.110 910.670 ;
        RECT 364.930 731.090 366.110 732.270 ;
        RECT 364.930 729.490 366.110 730.670 ;
        RECT 364.930 551.090 366.110 552.270 ;
        RECT 364.930 549.490 366.110 550.670 ;
        RECT 364.930 371.090 366.110 372.270 ;
        RECT 364.930 369.490 366.110 370.670 ;
        RECT 364.930 191.090 366.110 192.270 ;
        RECT 364.930 189.490 366.110 190.670 ;
        RECT 364.930 11.090 366.110 12.270 ;
        RECT 364.930 9.490 366.110 10.670 ;
        RECT 364.930 -2.910 366.110 -1.730 ;
        RECT 364.930 -4.510 366.110 -3.330 ;
        RECT 382.930 929.090 384.110 930.270 ;
        RECT 382.930 927.490 384.110 928.670 ;
        RECT 382.930 749.090 384.110 750.270 ;
        RECT 382.930 747.490 384.110 748.670 ;
        RECT 382.930 569.090 384.110 570.270 ;
        RECT 382.930 567.490 384.110 568.670 ;
        RECT 382.930 389.090 384.110 390.270 ;
        RECT 382.930 387.490 384.110 388.670 ;
        RECT 382.930 209.090 384.110 210.270 ;
        RECT 382.930 207.490 384.110 208.670 ;
        RECT 382.930 29.090 384.110 30.270 ;
        RECT 382.930 27.490 384.110 28.670 ;
        RECT 382.930 -12.310 384.110 -11.130 ;
        RECT 382.930 -13.910 384.110 -12.730 ;
        RECT 400.930 947.090 402.110 948.270 ;
        RECT 400.930 945.490 402.110 946.670 ;
        RECT 400.930 767.090 402.110 768.270 ;
        RECT 400.930 765.490 402.110 766.670 ;
        RECT 400.930 587.090 402.110 588.270 ;
        RECT 400.930 585.490 402.110 586.670 ;
        RECT 400.930 407.090 402.110 408.270 ;
        RECT 400.930 405.490 402.110 406.670 ;
        RECT 400.930 227.090 402.110 228.270 ;
        RECT 400.930 225.490 402.110 226.670 ;
        RECT 400.930 47.090 402.110 48.270 ;
        RECT 400.930 45.490 402.110 46.670 ;
        RECT 400.930 -21.710 402.110 -20.530 ;
        RECT 400.930 -23.310 402.110 -22.130 ;
        RECT 418.930 965.090 420.110 966.270 ;
        RECT 418.930 963.490 420.110 964.670 ;
        RECT 418.930 785.090 420.110 786.270 ;
        RECT 418.930 783.490 420.110 784.670 ;
        RECT 418.930 605.090 420.110 606.270 ;
        RECT 418.930 603.490 420.110 604.670 ;
        RECT 418.930 425.090 420.110 426.270 ;
        RECT 418.930 423.490 420.110 424.670 ;
        RECT 418.930 245.090 420.110 246.270 ;
        RECT 418.930 243.490 420.110 244.670 ;
        RECT 418.930 65.090 420.110 66.270 ;
        RECT 418.930 63.490 420.110 64.670 ;
        RECT 238.930 -31.110 240.110 -29.930 ;
        RECT 238.930 -32.710 240.110 -31.530 ;
        RECT 544.930 911.090 546.110 912.270 ;
        RECT 544.930 909.490 546.110 910.670 ;
        RECT 544.930 731.090 546.110 732.270 ;
        RECT 544.930 729.490 546.110 730.670 ;
        RECT 544.930 551.090 546.110 552.270 ;
        RECT 544.930 549.490 546.110 550.670 ;
        RECT 544.930 371.090 546.110 372.270 ;
        RECT 544.930 369.490 546.110 370.670 ;
        RECT 544.930 191.090 546.110 192.270 ;
        RECT 544.930 189.490 546.110 190.670 ;
        RECT 544.930 11.090 546.110 12.270 ;
        RECT 544.930 9.490 546.110 10.670 ;
        RECT 544.930 -2.910 546.110 -1.730 ;
        RECT 544.930 -4.510 546.110 -3.330 ;
        RECT 562.930 929.090 564.110 930.270 ;
        RECT 562.930 927.490 564.110 928.670 ;
        RECT 562.930 749.090 564.110 750.270 ;
        RECT 562.930 747.490 564.110 748.670 ;
        RECT 562.930 569.090 564.110 570.270 ;
        RECT 562.930 567.490 564.110 568.670 ;
        RECT 562.930 389.090 564.110 390.270 ;
        RECT 562.930 387.490 564.110 388.670 ;
        RECT 562.930 209.090 564.110 210.270 ;
        RECT 562.930 207.490 564.110 208.670 ;
        RECT 562.930 29.090 564.110 30.270 ;
        RECT 562.930 27.490 564.110 28.670 ;
        RECT 562.930 -12.310 564.110 -11.130 ;
        RECT 562.930 -13.910 564.110 -12.730 ;
        RECT 580.930 947.090 582.110 948.270 ;
        RECT 580.930 945.490 582.110 946.670 ;
        RECT 580.930 767.090 582.110 768.270 ;
        RECT 580.930 765.490 582.110 766.670 ;
        RECT 580.930 587.090 582.110 588.270 ;
        RECT 580.930 585.490 582.110 586.670 ;
        RECT 580.930 407.090 582.110 408.270 ;
        RECT 580.930 405.490 582.110 406.670 ;
        RECT 580.930 227.090 582.110 228.270 ;
        RECT 580.930 225.490 582.110 226.670 ;
        RECT 580.930 47.090 582.110 48.270 ;
        RECT 580.930 45.490 582.110 46.670 ;
        RECT 580.930 -21.710 582.110 -20.530 ;
        RECT 580.930 -23.310 582.110 -22.130 ;
        RECT 598.930 965.090 600.110 966.270 ;
        RECT 598.930 963.490 600.110 964.670 ;
        RECT 598.930 785.090 600.110 786.270 ;
        RECT 598.930 783.490 600.110 784.670 ;
        RECT 598.930 605.090 600.110 606.270 ;
        RECT 598.930 603.490 600.110 604.670 ;
        RECT 598.930 425.090 600.110 426.270 ;
        RECT 598.930 423.490 600.110 424.670 ;
        RECT 598.930 245.090 600.110 246.270 ;
        RECT 598.930 243.490 600.110 244.670 ;
        RECT 598.930 65.090 600.110 66.270 ;
        RECT 598.930 63.490 600.110 64.670 ;
        RECT 418.930 -31.110 420.110 -29.930 ;
        RECT 418.930 -32.710 420.110 -31.530 ;
        RECT 724.930 911.090 726.110 912.270 ;
        RECT 724.930 909.490 726.110 910.670 ;
        RECT 724.930 731.090 726.110 732.270 ;
        RECT 724.930 729.490 726.110 730.670 ;
        RECT 724.930 551.090 726.110 552.270 ;
        RECT 724.930 549.490 726.110 550.670 ;
        RECT 724.930 371.090 726.110 372.270 ;
        RECT 724.930 369.490 726.110 370.670 ;
        RECT 724.930 191.090 726.110 192.270 ;
        RECT 724.930 189.490 726.110 190.670 ;
        RECT 724.930 11.090 726.110 12.270 ;
        RECT 724.930 9.490 726.110 10.670 ;
        RECT 724.930 -2.910 726.110 -1.730 ;
        RECT 724.930 -4.510 726.110 -3.330 ;
        RECT 742.930 929.090 744.110 930.270 ;
        RECT 742.930 927.490 744.110 928.670 ;
        RECT 742.930 749.090 744.110 750.270 ;
        RECT 742.930 747.490 744.110 748.670 ;
        RECT 742.930 569.090 744.110 570.270 ;
        RECT 742.930 567.490 744.110 568.670 ;
        RECT 742.930 389.090 744.110 390.270 ;
        RECT 742.930 387.490 744.110 388.670 ;
        RECT 742.930 209.090 744.110 210.270 ;
        RECT 742.930 207.490 744.110 208.670 ;
        RECT 742.930 29.090 744.110 30.270 ;
        RECT 742.930 27.490 744.110 28.670 ;
        RECT 742.930 -12.310 744.110 -11.130 ;
        RECT 742.930 -13.910 744.110 -12.730 ;
        RECT 760.930 947.090 762.110 948.270 ;
        RECT 760.930 945.490 762.110 946.670 ;
        RECT 760.930 767.090 762.110 768.270 ;
        RECT 760.930 765.490 762.110 766.670 ;
        RECT 760.930 587.090 762.110 588.270 ;
        RECT 760.930 585.490 762.110 586.670 ;
        RECT 760.930 407.090 762.110 408.270 ;
        RECT 760.930 405.490 762.110 406.670 ;
        RECT 760.930 227.090 762.110 228.270 ;
        RECT 760.930 225.490 762.110 226.670 ;
        RECT 760.930 47.090 762.110 48.270 ;
        RECT 760.930 45.490 762.110 46.670 ;
        RECT 760.930 -21.710 762.110 -20.530 ;
        RECT 760.930 -23.310 762.110 -22.130 ;
        RECT 778.930 965.090 780.110 966.270 ;
        RECT 778.930 963.490 780.110 964.670 ;
        RECT 778.930 785.090 780.110 786.270 ;
        RECT 778.930 783.490 780.110 784.670 ;
        RECT 778.930 605.090 780.110 606.270 ;
        RECT 778.930 603.490 780.110 604.670 ;
        RECT 778.930 425.090 780.110 426.270 ;
        RECT 778.930 423.490 780.110 424.670 ;
        RECT 778.930 245.090 780.110 246.270 ;
        RECT 778.930 243.490 780.110 244.670 ;
        RECT 778.930 65.090 780.110 66.270 ;
        RECT 778.930 63.490 780.110 64.670 ;
        RECT 598.930 -31.110 600.110 -29.930 ;
        RECT 598.930 -32.710 600.110 -31.530 ;
        RECT 904.930 911.090 906.110 912.270 ;
        RECT 904.930 909.490 906.110 910.670 ;
        RECT 904.930 731.090 906.110 732.270 ;
        RECT 904.930 729.490 906.110 730.670 ;
        RECT 904.930 551.090 906.110 552.270 ;
        RECT 904.930 549.490 906.110 550.670 ;
        RECT 904.930 371.090 906.110 372.270 ;
        RECT 904.930 369.490 906.110 370.670 ;
        RECT 904.930 191.090 906.110 192.270 ;
        RECT 904.930 189.490 906.110 190.670 ;
        RECT 904.930 11.090 906.110 12.270 ;
        RECT 904.930 9.490 906.110 10.670 ;
        RECT 904.930 -2.910 906.110 -1.730 ;
        RECT 904.930 -4.510 906.110 -3.330 ;
        RECT 922.930 929.090 924.110 930.270 ;
        RECT 922.930 927.490 924.110 928.670 ;
        RECT 922.930 749.090 924.110 750.270 ;
        RECT 922.930 747.490 924.110 748.670 ;
        RECT 922.930 569.090 924.110 570.270 ;
        RECT 922.930 567.490 924.110 568.670 ;
        RECT 922.930 389.090 924.110 390.270 ;
        RECT 922.930 387.490 924.110 388.670 ;
        RECT 922.930 209.090 924.110 210.270 ;
        RECT 922.930 207.490 924.110 208.670 ;
        RECT 922.930 29.090 924.110 30.270 ;
        RECT 922.930 27.490 924.110 28.670 ;
        RECT 922.930 -12.310 924.110 -11.130 ;
        RECT 922.930 -13.910 924.110 -12.730 ;
        RECT 940.930 947.090 942.110 948.270 ;
        RECT 940.930 945.490 942.110 946.670 ;
        RECT 940.930 767.090 942.110 768.270 ;
        RECT 940.930 765.490 942.110 766.670 ;
        RECT 940.930 587.090 942.110 588.270 ;
        RECT 940.930 585.490 942.110 586.670 ;
        RECT 940.930 407.090 942.110 408.270 ;
        RECT 940.930 405.490 942.110 406.670 ;
        RECT 940.930 227.090 942.110 228.270 ;
        RECT 940.930 225.490 942.110 226.670 ;
        RECT 940.930 47.090 942.110 48.270 ;
        RECT 940.930 45.490 942.110 46.670 ;
        RECT 940.930 -21.710 942.110 -20.530 ;
        RECT 940.930 -23.310 942.110 -22.130 ;
        RECT 958.930 965.090 960.110 966.270 ;
        RECT 958.930 963.490 960.110 964.670 ;
        RECT 958.930 785.090 960.110 786.270 ;
        RECT 958.930 783.490 960.110 784.670 ;
        RECT 958.930 605.090 960.110 606.270 ;
        RECT 958.930 603.490 960.110 604.670 ;
        RECT 958.930 425.090 960.110 426.270 ;
        RECT 958.930 423.490 960.110 424.670 ;
        RECT 958.930 245.090 960.110 246.270 ;
        RECT 958.930 243.490 960.110 244.670 ;
        RECT 958.930 65.090 960.110 66.270 ;
        RECT 958.930 63.490 960.110 64.670 ;
        RECT 778.930 -31.110 780.110 -29.930 ;
        RECT 778.930 -32.710 780.110 -31.530 ;
        RECT 1084.930 911.090 1086.110 912.270 ;
        RECT 1084.930 909.490 1086.110 910.670 ;
        RECT 1084.930 731.090 1086.110 732.270 ;
        RECT 1084.930 729.490 1086.110 730.670 ;
        RECT 1084.930 551.090 1086.110 552.270 ;
        RECT 1084.930 549.490 1086.110 550.670 ;
        RECT 1084.930 371.090 1086.110 372.270 ;
        RECT 1084.930 369.490 1086.110 370.670 ;
        RECT 1084.930 191.090 1086.110 192.270 ;
        RECT 1084.930 189.490 1086.110 190.670 ;
        RECT 1084.930 11.090 1086.110 12.270 ;
        RECT 1084.930 9.490 1086.110 10.670 ;
        RECT 1084.930 -2.910 1086.110 -1.730 ;
        RECT 1084.930 -4.510 1086.110 -3.330 ;
        RECT 1102.930 929.090 1104.110 930.270 ;
        RECT 1102.930 927.490 1104.110 928.670 ;
        RECT 1102.930 749.090 1104.110 750.270 ;
        RECT 1102.930 747.490 1104.110 748.670 ;
        RECT 1102.930 569.090 1104.110 570.270 ;
        RECT 1102.930 567.490 1104.110 568.670 ;
        RECT 1102.930 389.090 1104.110 390.270 ;
        RECT 1102.930 387.490 1104.110 388.670 ;
        RECT 1102.930 209.090 1104.110 210.270 ;
        RECT 1102.930 207.490 1104.110 208.670 ;
        RECT 1102.930 29.090 1104.110 30.270 ;
        RECT 1102.930 27.490 1104.110 28.670 ;
        RECT 1102.930 -12.310 1104.110 -11.130 ;
        RECT 1102.930 -13.910 1104.110 -12.730 ;
        RECT 1120.930 947.090 1122.110 948.270 ;
        RECT 1120.930 945.490 1122.110 946.670 ;
        RECT 1120.930 767.090 1122.110 768.270 ;
        RECT 1120.930 765.490 1122.110 766.670 ;
        RECT 1120.930 587.090 1122.110 588.270 ;
        RECT 1120.930 585.490 1122.110 586.670 ;
        RECT 1120.930 407.090 1122.110 408.270 ;
        RECT 1120.930 405.490 1122.110 406.670 ;
        RECT 1120.930 227.090 1122.110 228.270 ;
        RECT 1120.930 225.490 1122.110 226.670 ;
        RECT 1120.930 47.090 1122.110 48.270 ;
        RECT 1120.930 45.490 1122.110 46.670 ;
        RECT 1120.930 -21.710 1122.110 -20.530 ;
        RECT 1120.930 -23.310 1122.110 -22.130 ;
        RECT 1138.930 965.090 1140.110 966.270 ;
        RECT 1138.930 963.490 1140.110 964.670 ;
        RECT 1138.930 785.090 1140.110 786.270 ;
        RECT 1138.930 783.490 1140.110 784.670 ;
        RECT 1138.930 605.090 1140.110 606.270 ;
        RECT 1138.930 603.490 1140.110 604.670 ;
        RECT 1138.930 425.090 1140.110 426.270 ;
        RECT 1138.930 423.490 1140.110 424.670 ;
        RECT 1138.930 245.090 1140.110 246.270 ;
        RECT 1138.930 243.490 1140.110 244.670 ;
        RECT 1138.930 65.090 1140.110 66.270 ;
        RECT 1138.930 63.490 1140.110 64.670 ;
        RECT 958.930 -31.110 960.110 -29.930 ;
        RECT 958.930 -32.710 960.110 -31.530 ;
        RECT 1264.930 911.090 1266.110 912.270 ;
        RECT 1264.930 909.490 1266.110 910.670 ;
        RECT 1264.930 731.090 1266.110 732.270 ;
        RECT 1264.930 729.490 1266.110 730.670 ;
        RECT 1264.930 551.090 1266.110 552.270 ;
        RECT 1264.930 549.490 1266.110 550.670 ;
        RECT 1264.930 371.090 1266.110 372.270 ;
        RECT 1264.930 369.490 1266.110 370.670 ;
        RECT 1264.930 191.090 1266.110 192.270 ;
        RECT 1264.930 189.490 1266.110 190.670 ;
        RECT 1264.930 11.090 1266.110 12.270 ;
        RECT 1264.930 9.490 1266.110 10.670 ;
        RECT 1264.930 -2.910 1266.110 -1.730 ;
        RECT 1264.930 -4.510 1266.110 -3.330 ;
        RECT 1282.930 929.090 1284.110 930.270 ;
        RECT 1282.930 927.490 1284.110 928.670 ;
        RECT 1282.930 749.090 1284.110 750.270 ;
        RECT 1282.930 747.490 1284.110 748.670 ;
        RECT 1282.930 569.090 1284.110 570.270 ;
        RECT 1282.930 567.490 1284.110 568.670 ;
        RECT 1282.930 389.090 1284.110 390.270 ;
        RECT 1282.930 387.490 1284.110 388.670 ;
        RECT 1282.930 209.090 1284.110 210.270 ;
        RECT 1282.930 207.490 1284.110 208.670 ;
        RECT 1282.930 29.090 1284.110 30.270 ;
        RECT 1282.930 27.490 1284.110 28.670 ;
        RECT 1282.930 -12.310 1284.110 -11.130 ;
        RECT 1282.930 -13.910 1284.110 -12.730 ;
        RECT 1300.930 947.090 1302.110 948.270 ;
        RECT 1300.930 945.490 1302.110 946.670 ;
        RECT 1300.930 767.090 1302.110 768.270 ;
        RECT 1300.930 765.490 1302.110 766.670 ;
        RECT 1300.930 587.090 1302.110 588.270 ;
        RECT 1300.930 585.490 1302.110 586.670 ;
        RECT 1300.930 407.090 1302.110 408.270 ;
        RECT 1300.930 405.490 1302.110 406.670 ;
        RECT 1300.930 227.090 1302.110 228.270 ;
        RECT 1300.930 225.490 1302.110 226.670 ;
        RECT 1300.930 47.090 1302.110 48.270 ;
        RECT 1300.930 45.490 1302.110 46.670 ;
        RECT 1300.930 -21.710 1302.110 -20.530 ;
        RECT 1300.930 -23.310 1302.110 -22.130 ;
        RECT 1318.930 965.090 1320.110 966.270 ;
        RECT 1318.930 963.490 1320.110 964.670 ;
        RECT 1318.930 785.090 1320.110 786.270 ;
        RECT 1318.930 783.490 1320.110 784.670 ;
        RECT 1318.930 605.090 1320.110 606.270 ;
        RECT 1318.930 603.490 1320.110 604.670 ;
        RECT 1318.930 425.090 1320.110 426.270 ;
        RECT 1318.930 423.490 1320.110 424.670 ;
        RECT 1318.930 245.090 1320.110 246.270 ;
        RECT 1318.930 243.490 1320.110 244.670 ;
        RECT 1318.930 65.090 1320.110 66.270 ;
        RECT 1318.930 63.490 1320.110 64.670 ;
        RECT 1138.930 -31.110 1140.110 -29.930 ;
        RECT 1138.930 -32.710 1140.110 -31.530 ;
        RECT 1444.930 911.090 1446.110 912.270 ;
        RECT 1444.930 909.490 1446.110 910.670 ;
        RECT 1444.930 731.090 1446.110 732.270 ;
        RECT 1444.930 729.490 1446.110 730.670 ;
        RECT 1444.930 551.090 1446.110 552.270 ;
        RECT 1444.930 549.490 1446.110 550.670 ;
        RECT 1444.930 371.090 1446.110 372.270 ;
        RECT 1444.930 369.490 1446.110 370.670 ;
        RECT 1444.930 191.090 1446.110 192.270 ;
        RECT 1444.930 189.490 1446.110 190.670 ;
        RECT 1444.930 11.090 1446.110 12.270 ;
        RECT 1444.930 9.490 1446.110 10.670 ;
        RECT 1444.930 -2.910 1446.110 -1.730 ;
        RECT 1444.930 -4.510 1446.110 -3.330 ;
        RECT 1462.930 929.090 1464.110 930.270 ;
        RECT 1462.930 927.490 1464.110 928.670 ;
        RECT 1462.930 749.090 1464.110 750.270 ;
        RECT 1462.930 747.490 1464.110 748.670 ;
        RECT 1462.930 569.090 1464.110 570.270 ;
        RECT 1462.930 567.490 1464.110 568.670 ;
        RECT 1462.930 389.090 1464.110 390.270 ;
        RECT 1462.930 387.490 1464.110 388.670 ;
        RECT 1462.930 209.090 1464.110 210.270 ;
        RECT 1462.930 207.490 1464.110 208.670 ;
        RECT 1462.930 29.090 1464.110 30.270 ;
        RECT 1462.930 27.490 1464.110 28.670 ;
        RECT 1462.930 -12.310 1464.110 -11.130 ;
        RECT 1462.930 -13.910 1464.110 -12.730 ;
        RECT 1480.930 947.090 1482.110 948.270 ;
        RECT 1480.930 945.490 1482.110 946.670 ;
        RECT 1480.930 767.090 1482.110 768.270 ;
        RECT 1480.930 765.490 1482.110 766.670 ;
        RECT 1480.930 587.090 1482.110 588.270 ;
        RECT 1480.930 585.490 1482.110 586.670 ;
        RECT 1480.930 407.090 1482.110 408.270 ;
        RECT 1480.930 405.490 1482.110 406.670 ;
        RECT 1480.930 227.090 1482.110 228.270 ;
        RECT 1480.930 225.490 1482.110 226.670 ;
        RECT 1480.930 47.090 1482.110 48.270 ;
        RECT 1480.930 45.490 1482.110 46.670 ;
        RECT 1480.930 -21.710 1482.110 -20.530 ;
        RECT 1480.930 -23.310 1482.110 -22.130 ;
        RECT 1498.930 965.090 1500.110 966.270 ;
        RECT 1498.930 963.490 1500.110 964.670 ;
        RECT 1498.930 785.090 1500.110 786.270 ;
        RECT 1498.930 783.490 1500.110 784.670 ;
        RECT 1498.930 605.090 1500.110 606.270 ;
        RECT 1498.930 603.490 1500.110 604.670 ;
        RECT 1498.930 425.090 1500.110 426.270 ;
        RECT 1498.930 423.490 1500.110 424.670 ;
        RECT 1498.930 245.090 1500.110 246.270 ;
        RECT 1498.930 243.490 1500.110 244.670 ;
        RECT 1498.930 65.090 1500.110 66.270 ;
        RECT 1498.930 63.490 1500.110 64.670 ;
        RECT 1318.930 -31.110 1320.110 -29.930 ;
        RECT 1318.930 -32.710 1320.110 -31.530 ;
        RECT 1624.930 911.090 1626.110 912.270 ;
        RECT 1624.930 909.490 1626.110 910.670 ;
        RECT 1624.930 731.090 1626.110 732.270 ;
        RECT 1624.930 729.490 1626.110 730.670 ;
        RECT 1624.930 551.090 1626.110 552.270 ;
        RECT 1624.930 549.490 1626.110 550.670 ;
        RECT 1624.930 371.090 1626.110 372.270 ;
        RECT 1624.930 369.490 1626.110 370.670 ;
        RECT 1624.930 191.090 1626.110 192.270 ;
        RECT 1624.930 189.490 1626.110 190.670 ;
        RECT 1624.930 11.090 1626.110 12.270 ;
        RECT 1624.930 9.490 1626.110 10.670 ;
        RECT 1624.930 -2.910 1626.110 -1.730 ;
        RECT 1624.930 -4.510 1626.110 -3.330 ;
        RECT 1642.930 2189.090 1644.110 2190.270 ;
        RECT 1642.930 2187.490 1644.110 2188.670 ;
        RECT 1642.930 2009.090 1644.110 2010.270 ;
        RECT 1642.930 2007.490 1644.110 2008.670 ;
        RECT 1642.930 1829.090 1644.110 1830.270 ;
        RECT 1642.930 1827.490 1644.110 1828.670 ;
        RECT 1642.930 1649.090 1644.110 1650.270 ;
        RECT 1642.930 1647.490 1644.110 1648.670 ;
        RECT 1642.930 1469.090 1644.110 1470.270 ;
        RECT 1642.930 1467.490 1644.110 1468.670 ;
        RECT 1642.930 1289.090 1644.110 1290.270 ;
        RECT 1642.930 1287.490 1644.110 1288.670 ;
        RECT 1642.930 1109.090 1644.110 1110.270 ;
        RECT 1642.930 1107.490 1644.110 1108.670 ;
        RECT 1642.930 929.090 1644.110 930.270 ;
        RECT 1642.930 927.490 1644.110 928.670 ;
        RECT 1642.930 749.090 1644.110 750.270 ;
        RECT 1642.930 747.490 1644.110 748.670 ;
        RECT 1642.930 569.090 1644.110 570.270 ;
        RECT 1642.930 567.490 1644.110 568.670 ;
        RECT 1642.930 389.090 1644.110 390.270 ;
        RECT 1642.930 387.490 1644.110 388.670 ;
        RECT 1642.930 209.090 1644.110 210.270 ;
        RECT 1642.930 207.490 1644.110 208.670 ;
        RECT 1642.930 29.090 1644.110 30.270 ;
        RECT 1642.930 27.490 1644.110 28.670 ;
        RECT 1642.930 -12.310 1644.110 -11.130 ;
        RECT 1642.930 -13.910 1644.110 -12.730 ;
        RECT 1660.930 2207.090 1662.110 2208.270 ;
        RECT 1660.930 2205.490 1662.110 2206.670 ;
        RECT 1660.930 2027.090 1662.110 2028.270 ;
        RECT 1660.930 2025.490 1662.110 2026.670 ;
        RECT 1660.930 1847.090 1662.110 1848.270 ;
        RECT 1660.930 1845.490 1662.110 1846.670 ;
        RECT 1660.930 1667.090 1662.110 1668.270 ;
        RECT 1660.930 1665.490 1662.110 1666.670 ;
        RECT 1660.930 1487.090 1662.110 1488.270 ;
        RECT 1660.930 1485.490 1662.110 1486.670 ;
        RECT 1660.930 1307.090 1662.110 1308.270 ;
        RECT 1660.930 1305.490 1662.110 1306.670 ;
        RECT 1660.930 1127.090 1662.110 1128.270 ;
        RECT 1660.930 1125.490 1662.110 1126.670 ;
        RECT 1660.930 947.090 1662.110 948.270 ;
        RECT 1660.930 945.490 1662.110 946.670 ;
        RECT 1660.930 767.090 1662.110 768.270 ;
        RECT 1660.930 765.490 1662.110 766.670 ;
        RECT 1660.930 587.090 1662.110 588.270 ;
        RECT 1660.930 585.490 1662.110 586.670 ;
        RECT 1660.930 407.090 1662.110 408.270 ;
        RECT 1660.930 405.490 1662.110 406.670 ;
        RECT 1660.930 227.090 1662.110 228.270 ;
        RECT 1660.930 225.490 1662.110 226.670 ;
        RECT 1660.930 47.090 1662.110 48.270 ;
        RECT 1660.930 45.490 1662.110 46.670 ;
        RECT 1660.930 -21.710 1662.110 -20.530 ;
        RECT 1660.930 -23.310 1662.110 -22.130 ;
        RECT 1678.930 2225.090 1680.110 2226.270 ;
        RECT 1678.930 2223.490 1680.110 2224.670 ;
        RECT 1678.930 2045.090 1680.110 2046.270 ;
        RECT 1678.930 2043.490 1680.110 2044.670 ;
        RECT 1678.930 1865.090 1680.110 1866.270 ;
        RECT 1678.930 1863.490 1680.110 1864.670 ;
        RECT 1678.930 1685.090 1680.110 1686.270 ;
        RECT 1678.930 1683.490 1680.110 1684.670 ;
        RECT 1678.930 1505.090 1680.110 1506.270 ;
        RECT 1678.930 1503.490 1680.110 1504.670 ;
        RECT 1678.930 1325.090 1680.110 1326.270 ;
        RECT 1678.930 1323.490 1680.110 1324.670 ;
        RECT 1678.930 1145.090 1680.110 1146.270 ;
        RECT 1678.930 1143.490 1680.110 1144.670 ;
        RECT 1678.930 965.090 1680.110 966.270 ;
        RECT 1678.930 963.490 1680.110 964.670 ;
        RECT 1678.930 785.090 1680.110 786.270 ;
        RECT 1678.930 783.490 1680.110 784.670 ;
        RECT 1678.930 605.090 1680.110 606.270 ;
        RECT 1678.930 603.490 1680.110 604.670 ;
        RECT 1678.930 425.090 1680.110 426.270 ;
        RECT 1678.930 423.490 1680.110 424.670 ;
        RECT 1678.930 245.090 1680.110 246.270 ;
        RECT 1678.930 243.490 1680.110 244.670 ;
        RECT 1678.930 65.090 1680.110 66.270 ;
        RECT 1678.930 63.490 1680.110 64.670 ;
        RECT 1498.930 -31.110 1500.110 -29.930 ;
        RECT 1498.930 -32.710 1500.110 -31.530 ;
        RECT 1804.930 2171.090 1806.110 2172.270 ;
        RECT 1804.930 2169.490 1806.110 2170.670 ;
        RECT 1804.930 1991.090 1806.110 1992.270 ;
        RECT 1804.930 1989.490 1806.110 1990.670 ;
        RECT 1804.930 1811.090 1806.110 1812.270 ;
        RECT 1804.930 1809.490 1806.110 1810.670 ;
        RECT 1804.930 1631.090 1806.110 1632.270 ;
        RECT 1804.930 1629.490 1806.110 1630.670 ;
        RECT 1804.930 1451.090 1806.110 1452.270 ;
        RECT 1804.930 1449.490 1806.110 1450.670 ;
        RECT 1804.930 1271.090 1806.110 1272.270 ;
        RECT 1804.930 1269.490 1806.110 1270.670 ;
        RECT 1804.930 1091.090 1806.110 1092.270 ;
        RECT 1804.930 1089.490 1806.110 1090.670 ;
        RECT 1804.930 911.090 1806.110 912.270 ;
        RECT 1804.930 909.490 1806.110 910.670 ;
        RECT 1804.930 731.090 1806.110 732.270 ;
        RECT 1804.930 729.490 1806.110 730.670 ;
        RECT 1804.930 551.090 1806.110 552.270 ;
        RECT 1804.930 549.490 1806.110 550.670 ;
        RECT 1804.930 371.090 1806.110 372.270 ;
        RECT 1804.930 369.490 1806.110 370.670 ;
        RECT 1804.930 191.090 1806.110 192.270 ;
        RECT 1804.930 189.490 1806.110 190.670 ;
        RECT 1804.930 11.090 1806.110 12.270 ;
        RECT 1804.930 9.490 1806.110 10.670 ;
        RECT 1804.930 -2.910 1806.110 -1.730 ;
        RECT 1804.930 -4.510 1806.110 -3.330 ;
        RECT 1822.930 2189.090 1824.110 2190.270 ;
        RECT 1822.930 2187.490 1824.110 2188.670 ;
        RECT 1822.930 2009.090 1824.110 2010.270 ;
        RECT 1822.930 2007.490 1824.110 2008.670 ;
        RECT 1822.930 1829.090 1824.110 1830.270 ;
        RECT 1822.930 1827.490 1824.110 1828.670 ;
        RECT 1822.930 1649.090 1824.110 1650.270 ;
        RECT 1822.930 1647.490 1824.110 1648.670 ;
        RECT 1822.930 1469.090 1824.110 1470.270 ;
        RECT 1822.930 1467.490 1824.110 1468.670 ;
        RECT 1822.930 1289.090 1824.110 1290.270 ;
        RECT 1822.930 1287.490 1824.110 1288.670 ;
        RECT 1822.930 1109.090 1824.110 1110.270 ;
        RECT 1822.930 1107.490 1824.110 1108.670 ;
        RECT 1822.930 929.090 1824.110 930.270 ;
        RECT 1822.930 927.490 1824.110 928.670 ;
        RECT 1822.930 749.090 1824.110 750.270 ;
        RECT 1822.930 747.490 1824.110 748.670 ;
        RECT 1822.930 569.090 1824.110 570.270 ;
        RECT 1822.930 567.490 1824.110 568.670 ;
        RECT 1822.930 389.090 1824.110 390.270 ;
        RECT 1822.930 387.490 1824.110 388.670 ;
        RECT 1822.930 209.090 1824.110 210.270 ;
        RECT 1822.930 207.490 1824.110 208.670 ;
        RECT 1822.930 29.090 1824.110 30.270 ;
        RECT 1822.930 27.490 1824.110 28.670 ;
        RECT 1822.930 -12.310 1824.110 -11.130 ;
        RECT 1822.930 -13.910 1824.110 -12.730 ;
        RECT 1840.930 2207.090 1842.110 2208.270 ;
        RECT 1840.930 2205.490 1842.110 2206.670 ;
        RECT 1840.930 2027.090 1842.110 2028.270 ;
        RECT 1840.930 2025.490 1842.110 2026.670 ;
        RECT 1840.930 1847.090 1842.110 1848.270 ;
        RECT 1840.930 1845.490 1842.110 1846.670 ;
        RECT 1840.930 1667.090 1842.110 1668.270 ;
        RECT 1840.930 1665.490 1842.110 1666.670 ;
        RECT 1840.930 1487.090 1842.110 1488.270 ;
        RECT 1840.930 1485.490 1842.110 1486.670 ;
        RECT 1840.930 1307.090 1842.110 1308.270 ;
        RECT 1840.930 1305.490 1842.110 1306.670 ;
        RECT 1840.930 1127.090 1842.110 1128.270 ;
        RECT 1840.930 1125.490 1842.110 1126.670 ;
        RECT 1840.930 947.090 1842.110 948.270 ;
        RECT 1840.930 945.490 1842.110 946.670 ;
        RECT 1840.930 767.090 1842.110 768.270 ;
        RECT 1840.930 765.490 1842.110 766.670 ;
        RECT 1840.930 587.090 1842.110 588.270 ;
        RECT 1840.930 585.490 1842.110 586.670 ;
        RECT 1840.930 407.090 1842.110 408.270 ;
        RECT 1840.930 405.490 1842.110 406.670 ;
        RECT 1840.930 227.090 1842.110 228.270 ;
        RECT 1840.930 225.490 1842.110 226.670 ;
        RECT 1840.930 47.090 1842.110 48.270 ;
        RECT 1840.930 45.490 1842.110 46.670 ;
        RECT 1840.930 -21.710 1842.110 -20.530 ;
        RECT 1840.930 -23.310 1842.110 -22.130 ;
        RECT 1858.930 2225.090 1860.110 2226.270 ;
        RECT 1858.930 2223.490 1860.110 2224.670 ;
        RECT 1858.930 2045.090 1860.110 2046.270 ;
        RECT 1858.930 2043.490 1860.110 2044.670 ;
        RECT 1858.930 1865.090 1860.110 1866.270 ;
        RECT 1858.930 1863.490 1860.110 1864.670 ;
        RECT 1858.930 1685.090 1860.110 1686.270 ;
        RECT 1858.930 1683.490 1860.110 1684.670 ;
        RECT 1858.930 1505.090 1860.110 1506.270 ;
        RECT 1858.930 1503.490 1860.110 1504.670 ;
        RECT 1858.930 1325.090 1860.110 1326.270 ;
        RECT 1858.930 1323.490 1860.110 1324.670 ;
        RECT 1858.930 1145.090 1860.110 1146.270 ;
        RECT 1858.930 1143.490 1860.110 1144.670 ;
        RECT 1858.930 965.090 1860.110 966.270 ;
        RECT 1858.930 963.490 1860.110 964.670 ;
        RECT 1858.930 785.090 1860.110 786.270 ;
        RECT 1858.930 783.490 1860.110 784.670 ;
        RECT 1858.930 605.090 1860.110 606.270 ;
        RECT 1858.930 603.490 1860.110 604.670 ;
        RECT 1858.930 425.090 1860.110 426.270 ;
        RECT 1858.930 423.490 1860.110 424.670 ;
        RECT 1858.930 245.090 1860.110 246.270 ;
        RECT 1858.930 243.490 1860.110 244.670 ;
        RECT 1858.930 65.090 1860.110 66.270 ;
        RECT 1858.930 63.490 1860.110 64.670 ;
        RECT 1678.930 -31.110 1680.110 -29.930 ;
        RECT 1678.930 -32.710 1680.110 -31.530 ;
        RECT 1984.930 2171.090 1986.110 2172.270 ;
        RECT 1984.930 2169.490 1986.110 2170.670 ;
        RECT 1984.930 1991.090 1986.110 1992.270 ;
        RECT 1984.930 1989.490 1986.110 1990.670 ;
        RECT 1984.930 1811.090 1986.110 1812.270 ;
        RECT 1984.930 1809.490 1986.110 1810.670 ;
        RECT 1984.930 1631.090 1986.110 1632.270 ;
        RECT 1984.930 1629.490 1986.110 1630.670 ;
        RECT 1984.930 1451.090 1986.110 1452.270 ;
        RECT 1984.930 1449.490 1986.110 1450.670 ;
        RECT 1984.930 1271.090 1986.110 1272.270 ;
        RECT 1984.930 1269.490 1986.110 1270.670 ;
        RECT 1984.930 1091.090 1986.110 1092.270 ;
        RECT 1984.930 1089.490 1986.110 1090.670 ;
        RECT 1984.930 911.090 1986.110 912.270 ;
        RECT 1984.930 909.490 1986.110 910.670 ;
        RECT 1984.930 731.090 1986.110 732.270 ;
        RECT 1984.930 729.490 1986.110 730.670 ;
        RECT 1984.930 551.090 1986.110 552.270 ;
        RECT 1984.930 549.490 1986.110 550.670 ;
        RECT 1984.930 371.090 1986.110 372.270 ;
        RECT 1984.930 369.490 1986.110 370.670 ;
        RECT 1984.930 191.090 1986.110 192.270 ;
        RECT 1984.930 189.490 1986.110 190.670 ;
        RECT 1984.930 11.090 1986.110 12.270 ;
        RECT 1984.930 9.490 1986.110 10.670 ;
        RECT 1984.930 -2.910 1986.110 -1.730 ;
        RECT 1984.930 -4.510 1986.110 -3.330 ;
        RECT 2002.930 3449.090 2004.110 3450.270 ;
        RECT 2002.930 3447.490 2004.110 3448.670 ;
        RECT 2002.930 3269.090 2004.110 3270.270 ;
        RECT 2002.930 3267.490 2004.110 3268.670 ;
        RECT 2002.930 3089.090 2004.110 3090.270 ;
        RECT 2002.930 3087.490 2004.110 3088.670 ;
        RECT 2002.930 2909.090 2004.110 2910.270 ;
        RECT 2002.930 2907.490 2004.110 2908.670 ;
        RECT 2002.930 2729.090 2004.110 2730.270 ;
        RECT 2002.930 2727.490 2004.110 2728.670 ;
        RECT 2002.930 2549.090 2004.110 2550.270 ;
        RECT 2002.930 2547.490 2004.110 2548.670 ;
        RECT 2002.930 2369.090 2004.110 2370.270 ;
        RECT 2002.930 2367.490 2004.110 2368.670 ;
        RECT 2002.930 2189.090 2004.110 2190.270 ;
        RECT 2002.930 2187.490 2004.110 2188.670 ;
        RECT 2002.930 2009.090 2004.110 2010.270 ;
        RECT 2002.930 2007.490 2004.110 2008.670 ;
        RECT 2002.930 1829.090 2004.110 1830.270 ;
        RECT 2002.930 1827.490 2004.110 1828.670 ;
        RECT 2002.930 1649.090 2004.110 1650.270 ;
        RECT 2002.930 1647.490 2004.110 1648.670 ;
        RECT 2002.930 1469.090 2004.110 1470.270 ;
        RECT 2002.930 1467.490 2004.110 1468.670 ;
        RECT 2002.930 1289.090 2004.110 1290.270 ;
        RECT 2002.930 1287.490 2004.110 1288.670 ;
        RECT 2002.930 1109.090 2004.110 1110.270 ;
        RECT 2002.930 1107.490 2004.110 1108.670 ;
        RECT 2002.930 929.090 2004.110 930.270 ;
        RECT 2002.930 927.490 2004.110 928.670 ;
        RECT 2002.930 749.090 2004.110 750.270 ;
        RECT 2002.930 747.490 2004.110 748.670 ;
        RECT 2002.930 569.090 2004.110 570.270 ;
        RECT 2002.930 567.490 2004.110 568.670 ;
        RECT 2002.930 389.090 2004.110 390.270 ;
        RECT 2002.930 387.490 2004.110 388.670 ;
        RECT 2002.930 209.090 2004.110 210.270 ;
        RECT 2002.930 207.490 2004.110 208.670 ;
        RECT 2002.930 29.090 2004.110 30.270 ;
        RECT 2002.930 27.490 2004.110 28.670 ;
        RECT 2002.930 -12.310 2004.110 -11.130 ;
        RECT 2002.930 -13.910 2004.110 -12.730 ;
        RECT 2020.930 3467.090 2022.110 3468.270 ;
        RECT 2020.930 3465.490 2022.110 3466.670 ;
        RECT 2020.930 3287.090 2022.110 3288.270 ;
        RECT 2020.930 3285.490 2022.110 3286.670 ;
        RECT 2020.930 3107.090 2022.110 3108.270 ;
        RECT 2020.930 3105.490 2022.110 3106.670 ;
        RECT 2020.930 2927.090 2022.110 2928.270 ;
        RECT 2020.930 2925.490 2022.110 2926.670 ;
        RECT 2020.930 2747.090 2022.110 2748.270 ;
        RECT 2020.930 2745.490 2022.110 2746.670 ;
        RECT 2020.930 2567.090 2022.110 2568.270 ;
        RECT 2020.930 2565.490 2022.110 2566.670 ;
        RECT 2020.930 2387.090 2022.110 2388.270 ;
        RECT 2020.930 2385.490 2022.110 2386.670 ;
        RECT 2020.930 2207.090 2022.110 2208.270 ;
        RECT 2020.930 2205.490 2022.110 2206.670 ;
        RECT 2020.930 2027.090 2022.110 2028.270 ;
        RECT 2020.930 2025.490 2022.110 2026.670 ;
        RECT 2020.930 1847.090 2022.110 1848.270 ;
        RECT 2020.930 1845.490 2022.110 1846.670 ;
        RECT 2020.930 1667.090 2022.110 1668.270 ;
        RECT 2020.930 1665.490 2022.110 1666.670 ;
        RECT 2020.930 1487.090 2022.110 1488.270 ;
        RECT 2020.930 1485.490 2022.110 1486.670 ;
        RECT 2020.930 1307.090 2022.110 1308.270 ;
        RECT 2020.930 1305.490 2022.110 1306.670 ;
        RECT 2020.930 1127.090 2022.110 1128.270 ;
        RECT 2020.930 1125.490 2022.110 1126.670 ;
        RECT 2020.930 947.090 2022.110 948.270 ;
        RECT 2020.930 945.490 2022.110 946.670 ;
        RECT 2020.930 767.090 2022.110 768.270 ;
        RECT 2020.930 765.490 2022.110 766.670 ;
        RECT 2020.930 587.090 2022.110 588.270 ;
        RECT 2020.930 585.490 2022.110 586.670 ;
        RECT 2020.930 407.090 2022.110 408.270 ;
        RECT 2020.930 405.490 2022.110 406.670 ;
        RECT 2020.930 227.090 2022.110 228.270 ;
        RECT 2020.930 225.490 2022.110 226.670 ;
        RECT 2020.930 47.090 2022.110 48.270 ;
        RECT 2020.930 45.490 2022.110 46.670 ;
        RECT 2020.930 -21.710 2022.110 -20.530 ;
        RECT 2020.930 -23.310 2022.110 -22.130 ;
        RECT 2218.930 3551.210 2220.110 3552.390 ;
        RECT 2218.930 3549.610 2220.110 3550.790 ;
        RECT 2200.930 3541.810 2202.110 3542.990 ;
        RECT 2200.930 3540.210 2202.110 3541.390 ;
        RECT 2182.930 3532.410 2184.110 3533.590 ;
        RECT 2182.930 3530.810 2184.110 3531.990 ;
        RECT 2038.930 3485.090 2040.110 3486.270 ;
        RECT 2038.930 3483.490 2040.110 3484.670 ;
        RECT 2038.930 3305.090 2040.110 3306.270 ;
        RECT 2038.930 3303.490 2040.110 3304.670 ;
        RECT 2038.930 3125.090 2040.110 3126.270 ;
        RECT 2038.930 3123.490 2040.110 3124.670 ;
        RECT 2038.930 2945.090 2040.110 2946.270 ;
        RECT 2038.930 2943.490 2040.110 2944.670 ;
        RECT 2038.930 2765.090 2040.110 2766.270 ;
        RECT 2038.930 2763.490 2040.110 2764.670 ;
        RECT 2038.930 2585.090 2040.110 2586.270 ;
        RECT 2038.930 2583.490 2040.110 2584.670 ;
        RECT 2038.930 2405.090 2040.110 2406.270 ;
        RECT 2038.930 2403.490 2040.110 2404.670 ;
        RECT 2038.930 2225.090 2040.110 2226.270 ;
        RECT 2038.930 2223.490 2040.110 2224.670 ;
        RECT 2038.930 2045.090 2040.110 2046.270 ;
        RECT 2038.930 2043.490 2040.110 2044.670 ;
        RECT 2038.930 1865.090 2040.110 1866.270 ;
        RECT 2038.930 1863.490 2040.110 1864.670 ;
        RECT 2038.930 1685.090 2040.110 1686.270 ;
        RECT 2038.930 1683.490 2040.110 1684.670 ;
        RECT 2038.930 1505.090 2040.110 1506.270 ;
        RECT 2038.930 1503.490 2040.110 1504.670 ;
        RECT 2038.930 1325.090 2040.110 1326.270 ;
        RECT 2038.930 1323.490 2040.110 1324.670 ;
        RECT 2038.930 1145.090 2040.110 1146.270 ;
        RECT 2038.930 1143.490 2040.110 1144.670 ;
        RECT 2038.930 965.090 2040.110 966.270 ;
        RECT 2038.930 963.490 2040.110 964.670 ;
        RECT 2038.930 785.090 2040.110 786.270 ;
        RECT 2038.930 783.490 2040.110 784.670 ;
        RECT 2038.930 605.090 2040.110 606.270 ;
        RECT 2038.930 603.490 2040.110 604.670 ;
        RECT 2038.930 425.090 2040.110 426.270 ;
        RECT 2038.930 423.490 2040.110 424.670 ;
        RECT 2038.930 245.090 2040.110 246.270 ;
        RECT 2038.930 243.490 2040.110 244.670 ;
        RECT 2038.930 65.090 2040.110 66.270 ;
        RECT 2038.930 63.490 2040.110 64.670 ;
        RECT 1858.930 -31.110 1860.110 -29.930 ;
        RECT 1858.930 -32.710 1860.110 -31.530 ;
        RECT 2164.930 3523.010 2166.110 3524.190 ;
        RECT 2164.930 3521.410 2166.110 3522.590 ;
        RECT 2164.930 3431.090 2166.110 3432.270 ;
        RECT 2164.930 3429.490 2166.110 3430.670 ;
        RECT 2164.930 3251.090 2166.110 3252.270 ;
        RECT 2164.930 3249.490 2166.110 3250.670 ;
        RECT 2164.930 3071.090 2166.110 3072.270 ;
        RECT 2164.930 3069.490 2166.110 3070.670 ;
        RECT 2164.930 2891.090 2166.110 2892.270 ;
        RECT 2164.930 2889.490 2166.110 2890.670 ;
        RECT 2182.930 3449.090 2184.110 3450.270 ;
        RECT 2182.930 3447.490 2184.110 3448.670 ;
        RECT 2182.930 3269.090 2184.110 3270.270 ;
        RECT 2182.930 3267.490 2184.110 3268.670 ;
        RECT 2182.930 3089.090 2184.110 3090.270 ;
        RECT 2182.930 3087.490 2184.110 3088.670 ;
        RECT 2182.930 2909.090 2184.110 2910.270 ;
        RECT 2182.930 2907.490 2184.110 2908.670 ;
        RECT 2200.930 3467.090 2202.110 3468.270 ;
        RECT 2200.930 3465.490 2202.110 3466.670 ;
        RECT 2200.930 3287.090 2202.110 3288.270 ;
        RECT 2200.930 3285.490 2202.110 3286.670 ;
        RECT 2200.930 3107.090 2202.110 3108.270 ;
        RECT 2200.930 3105.490 2202.110 3106.670 ;
        RECT 2200.930 2927.090 2202.110 2928.270 ;
        RECT 2200.930 2925.490 2202.110 2926.670 ;
        RECT 2398.930 3551.210 2400.110 3552.390 ;
        RECT 2398.930 3549.610 2400.110 3550.790 ;
        RECT 2380.930 3541.810 2382.110 3542.990 ;
        RECT 2380.930 3540.210 2382.110 3541.390 ;
        RECT 2362.930 3532.410 2364.110 3533.590 ;
        RECT 2362.930 3530.810 2364.110 3531.990 ;
        RECT 2218.930 3485.090 2220.110 3486.270 ;
        RECT 2218.930 3483.490 2220.110 3484.670 ;
        RECT 2218.930 3305.090 2220.110 3306.270 ;
        RECT 2218.930 3303.490 2220.110 3304.670 ;
        RECT 2218.930 3125.090 2220.110 3126.270 ;
        RECT 2218.930 3123.490 2220.110 3124.670 ;
        RECT 2218.930 2945.090 2220.110 2946.270 ;
        RECT 2218.930 2943.490 2220.110 2944.670 ;
        RECT 2344.930 3523.010 2346.110 3524.190 ;
        RECT 2344.930 3521.410 2346.110 3522.590 ;
        RECT 2344.930 3431.090 2346.110 3432.270 ;
        RECT 2344.930 3429.490 2346.110 3430.670 ;
        RECT 2344.930 3251.090 2346.110 3252.270 ;
        RECT 2344.930 3249.490 2346.110 3250.670 ;
        RECT 2344.930 3071.090 2346.110 3072.270 ;
        RECT 2344.930 3069.490 2346.110 3070.670 ;
        RECT 2344.930 2891.090 2346.110 2892.270 ;
        RECT 2344.930 2889.490 2346.110 2890.670 ;
        RECT 2362.930 3449.090 2364.110 3450.270 ;
        RECT 2362.930 3447.490 2364.110 3448.670 ;
        RECT 2362.930 3269.090 2364.110 3270.270 ;
        RECT 2362.930 3267.490 2364.110 3268.670 ;
        RECT 2362.930 3089.090 2364.110 3090.270 ;
        RECT 2362.930 3087.490 2364.110 3088.670 ;
        RECT 2362.930 2909.090 2364.110 2910.270 ;
        RECT 2362.930 2907.490 2364.110 2908.670 ;
        RECT 2380.930 3467.090 2382.110 3468.270 ;
        RECT 2380.930 3465.490 2382.110 3466.670 ;
        RECT 2380.930 3287.090 2382.110 3288.270 ;
        RECT 2380.930 3285.490 2382.110 3286.670 ;
        RECT 2380.930 3107.090 2382.110 3108.270 ;
        RECT 2380.930 3105.490 2382.110 3106.670 ;
        RECT 2380.930 2927.090 2382.110 2928.270 ;
        RECT 2380.930 2925.490 2382.110 2926.670 ;
        RECT 2578.930 3551.210 2580.110 3552.390 ;
        RECT 2578.930 3549.610 2580.110 3550.790 ;
        RECT 2560.930 3541.810 2562.110 3542.990 ;
        RECT 2560.930 3540.210 2562.110 3541.390 ;
        RECT 2542.930 3532.410 2544.110 3533.590 ;
        RECT 2542.930 3530.810 2544.110 3531.990 ;
        RECT 2398.930 3485.090 2400.110 3486.270 ;
        RECT 2398.930 3483.490 2400.110 3484.670 ;
        RECT 2398.930 3305.090 2400.110 3306.270 ;
        RECT 2398.930 3303.490 2400.110 3304.670 ;
        RECT 2398.930 3125.090 2400.110 3126.270 ;
        RECT 2398.930 3123.490 2400.110 3124.670 ;
        RECT 2398.930 2945.090 2400.110 2946.270 ;
        RECT 2398.930 2943.490 2400.110 2944.670 ;
        RECT 2524.930 3523.010 2526.110 3524.190 ;
        RECT 2524.930 3521.410 2526.110 3522.590 ;
        RECT 2524.930 3431.090 2526.110 3432.270 ;
        RECT 2524.930 3429.490 2526.110 3430.670 ;
        RECT 2524.930 3251.090 2526.110 3252.270 ;
        RECT 2524.930 3249.490 2526.110 3250.670 ;
        RECT 2524.930 3071.090 2526.110 3072.270 ;
        RECT 2524.930 3069.490 2526.110 3070.670 ;
        RECT 2524.930 2891.090 2526.110 2892.270 ;
        RECT 2524.930 2889.490 2526.110 2890.670 ;
        RECT 2542.930 3449.090 2544.110 3450.270 ;
        RECT 2542.930 3447.490 2544.110 3448.670 ;
        RECT 2542.930 3269.090 2544.110 3270.270 ;
        RECT 2542.930 3267.490 2544.110 3268.670 ;
        RECT 2542.930 3089.090 2544.110 3090.270 ;
        RECT 2542.930 3087.490 2544.110 3088.670 ;
        RECT 2542.930 2909.090 2544.110 2910.270 ;
        RECT 2542.930 2907.490 2544.110 2908.670 ;
        RECT 2560.930 3467.090 2562.110 3468.270 ;
        RECT 2560.930 3465.490 2562.110 3466.670 ;
        RECT 2560.930 3287.090 2562.110 3288.270 ;
        RECT 2560.930 3285.490 2562.110 3286.670 ;
        RECT 2560.930 3107.090 2562.110 3108.270 ;
        RECT 2560.930 3105.490 2562.110 3106.670 ;
        RECT 2560.930 2927.090 2562.110 2928.270 ;
        RECT 2560.930 2925.490 2562.110 2926.670 ;
        RECT 2758.930 3551.210 2760.110 3552.390 ;
        RECT 2758.930 3549.610 2760.110 3550.790 ;
        RECT 2740.930 3541.810 2742.110 3542.990 ;
        RECT 2740.930 3540.210 2742.110 3541.390 ;
        RECT 2722.930 3532.410 2724.110 3533.590 ;
        RECT 2722.930 3530.810 2724.110 3531.990 ;
        RECT 2578.930 3485.090 2580.110 3486.270 ;
        RECT 2578.930 3483.490 2580.110 3484.670 ;
        RECT 2578.930 3305.090 2580.110 3306.270 ;
        RECT 2578.930 3303.490 2580.110 3304.670 ;
        RECT 2578.930 3125.090 2580.110 3126.270 ;
        RECT 2578.930 3123.490 2580.110 3124.670 ;
        RECT 2578.930 2945.090 2580.110 2946.270 ;
        RECT 2578.930 2943.490 2580.110 2944.670 ;
        RECT 2704.930 3523.010 2706.110 3524.190 ;
        RECT 2704.930 3521.410 2706.110 3522.590 ;
        RECT 2704.930 3431.090 2706.110 3432.270 ;
        RECT 2704.930 3429.490 2706.110 3430.670 ;
        RECT 2704.930 3251.090 2706.110 3252.270 ;
        RECT 2704.930 3249.490 2706.110 3250.670 ;
        RECT 2704.930 3071.090 2706.110 3072.270 ;
        RECT 2704.930 3069.490 2706.110 3070.670 ;
        RECT 2704.930 2891.090 2706.110 2892.270 ;
        RECT 2704.930 2889.490 2706.110 2890.670 ;
        RECT 2164.930 2711.090 2166.110 2712.270 ;
        RECT 2164.930 2709.490 2166.110 2710.670 ;
        RECT 2164.930 2531.090 2166.110 2532.270 ;
        RECT 2164.930 2529.490 2166.110 2530.670 ;
        RECT 2164.930 2351.090 2166.110 2352.270 ;
        RECT 2164.930 2349.490 2166.110 2350.670 ;
        RECT 2582.680 2729.090 2583.860 2730.270 ;
        RECT 2582.680 2727.490 2583.860 2728.670 ;
        RECT 2582.680 2711.090 2583.860 2712.270 ;
        RECT 2582.680 2709.490 2583.860 2710.670 ;
        RECT 2582.680 2585.090 2583.860 2586.270 ;
        RECT 2582.680 2583.490 2583.860 2584.670 ;
        RECT 2582.680 2567.090 2583.860 2568.270 ;
        RECT 2582.680 2565.490 2583.860 2566.670 ;
        RECT 2582.680 2549.090 2583.860 2550.270 ;
        RECT 2582.680 2547.490 2583.860 2548.670 ;
        RECT 2582.680 2531.090 2583.860 2532.270 ;
        RECT 2582.680 2529.490 2583.860 2530.670 ;
        RECT 2582.680 2405.090 2583.860 2406.270 ;
        RECT 2582.680 2403.490 2583.860 2404.670 ;
        RECT 2582.680 2387.090 2583.860 2388.270 ;
        RECT 2582.680 2385.490 2583.860 2386.670 ;
        RECT 2582.680 2369.090 2583.860 2370.270 ;
        RECT 2582.680 2367.490 2583.860 2368.670 ;
        RECT 2582.680 2351.090 2583.860 2352.270 ;
        RECT 2582.680 2349.490 2583.860 2350.670 ;
        RECT 2704.930 2711.090 2706.110 2712.270 ;
        RECT 2704.930 2709.490 2706.110 2710.670 ;
        RECT 2704.930 2531.090 2706.110 2532.270 ;
        RECT 2704.930 2529.490 2706.110 2530.670 ;
        RECT 2704.930 2351.090 2706.110 2352.270 ;
        RECT 2704.930 2349.490 2706.110 2350.670 ;
        RECT 2164.930 2171.090 2166.110 2172.270 ;
        RECT 2164.930 2169.490 2166.110 2170.670 ;
        RECT 2164.930 1991.090 2166.110 1992.270 ;
        RECT 2164.930 1989.490 2166.110 1990.670 ;
        RECT 2164.930 1811.090 2166.110 1812.270 ;
        RECT 2164.930 1809.490 2166.110 1810.670 ;
        RECT 2164.930 1631.090 2166.110 1632.270 ;
        RECT 2164.930 1629.490 2166.110 1630.670 ;
        RECT 2164.930 1451.090 2166.110 1452.270 ;
        RECT 2164.930 1449.490 2166.110 1450.670 ;
        RECT 2164.930 1271.090 2166.110 1272.270 ;
        RECT 2164.930 1269.490 2166.110 1270.670 ;
        RECT 2164.930 1091.090 2166.110 1092.270 ;
        RECT 2164.930 1089.490 2166.110 1090.670 ;
        RECT 2164.930 911.090 2166.110 912.270 ;
        RECT 2164.930 909.490 2166.110 910.670 ;
        RECT 2164.930 731.090 2166.110 732.270 ;
        RECT 2164.930 729.490 2166.110 730.670 ;
        RECT 2164.930 551.090 2166.110 552.270 ;
        RECT 2164.930 549.490 2166.110 550.670 ;
        RECT 2164.930 371.090 2166.110 372.270 ;
        RECT 2164.930 369.490 2166.110 370.670 ;
        RECT 2164.930 191.090 2166.110 192.270 ;
        RECT 2164.930 189.490 2166.110 190.670 ;
        RECT 2164.930 11.090 2166.110 12.270 ;
        RECT 2164.930 9.490 2166.110 10.670 ;
        RECT 2164.930 -2.910 2166.110 -1.730 ;
        RECT 2164.930 -4.510 2166.110 -3.330 ;
        RECT 2182.930 2189.090 2184.110 2190.270 ;
        RECT 2182.930 2187.490 2184.110 2188.670 ;
        RECT 2182.930 2009.090 2184.110 2010.270 ;
        RECT 2182.930 2007.490 2184.110 2008.670 ;
        RECT 2182.930 1829.090 2184.110 1830.270 ;
        RECT 2182.930 1827.490 2184.110 1828.670 ;
        RECT 2182.930 1649.090 2184.110 1650.270 ;
        RECT 2182.930 1647.490 2184.110 1648.670 ;
        RECT 2182.930 1469.090 2184.110 1470.270 ;
        RECT 2182.930 1467.490 2184.110 1468.670 ;
        RECT 2182.930 1289.090 2184.110 1290.270 ;
        RECT 2182.930 1287.490 2184.110 1288.670 ;
        RECT 2182.930 1109.090 2184.110 1110.270 ;
        RECT 2182.930 1107.490 2184.110 1108.670 ;
        RECT 2182.930 929.090 2184.110 930.270 ;
        RECT 2182.930 927.490 2184.110 928.670 ;
        RECT 2182.930 749.090 2184.110 750.270 ;
        RECT 2182.930 747.490 2184.110 748.670 ;
        RECT 2182.930 569.090 2184.110 570.270 ;
        RECT 2182.930 567.490 2184.110 568.670 ;
        RECT 2182.930 389.090 2184.110 390.270 ;
        RECT 2182.930 387.490 2184.110 388.670 ;
        RECT 2182.930 209.090 2184.110 210.270 ;
        RECT 2182.930 207.490 2184.110 208.670 ;
        RECT 2182.930 29.090 2184.110 30.270 ;
        RECT 2182.930 27.490 2184.110 28.670 ;
        RECT 2182.930 -12.310 2184.110 -11.130 ;
        RECT 2182.930 -13.910 2184.110 -12.730 ;
        RECT 2200.930 2207.090 2202.110 2208.270 ;
        RECT 2200.930 2205.490 2202.110 2206.670 ;
        RECT 2200.930 2027.090 2202.110 2028.270 ;
        RECT 2200.930 2025.490 2202.110 2026.670 ;
        RECT 2200.930 1847.090 2202.110 1848.270 ;
        RECT 2200.930 1845.490 2202.110 1846.670 ;
        RECT 2200.930 1667.090 2202.110 1668.270 ;
        RECT 2200.930 1665.490 2202.110 1666.670 ;
        RECT 2200.930 1487.090 2202.110 1488.270 ;
        RECT 2200.930 1485.490 2202.110 1486.670 ;
        RECT 2200.930 1307.090 2202.110 1308.270 ;
        RECT 2200.930 1305.490 2202.110 1306.670 ;
        RECT 2200.930 1127.090 2202.110 1128.270 ;
        RECT 2200.930 1125.490 2202.110 1126.670 ;
        RECT 2200.930 947.090 2202.110 948.270 ;
        RECT 2200.930 945.490 2202.110 946.670 ;
        RECT 2200.930 767.090 2202.110 768.270 ;
        RECT 2200.930 765.490 2202.110 766.670 ;
        RECT 2200.930 587.090 2202.110 588.270 ;
        RECT 2200.930 585.490 2202.110 586.670 ;
        RECT 2200.930 407.090 2202.110 408.270 ;
        RECT 2200.930 405.490 2202.110 406.670 ;
        RECT 2200.930 227.090 2202.110 228.270 ;
        RECT 2200.930 225.490 2202.110 226.670 ;
        RECT 2200.930 47.090 2202.110 48.270 ;
        RECT 2200.930 45.490 2202.110 46.670 ;
        RECT 2200.930 -21.710 2202.110 -20.530 ;
        RECT 2200.930 -23.310 2202.110 -22.130 ;
        RECT 2218.930 2225.090 2220.110 2226.270 ;
        RECT 2218.930 2223.490 2220.110 2224.670 ;
        RECT 2218.930 2045.090 2220.110 2046.270 ;
        RECT 2218.930 2043.490 2220.110 2044.670 ;
        RECT 2218.930 1865.090 2220.110 1866.270 ;
        RECT 2218.930 1863.490 2220.110 1864.670 ;
        RECT 2218.930 1685.090 2220.110 1686.270 ;
        RECT 2218.930 1683.490 2220.110 1684.670 ;
        RECT 2218.930 1505.090 2220.110 1506.270 ;
        RECT 2218.930 1503.490 2220.110 1504.670 ;
        RECT 2218.930 1325.090 2220.110 1326.270 ;
        RECT 2218.930 1323.490 2220.110 1324.670 ;
        RECT 2218.930 1145.090 2220.110 1146.270 ;
        RECT 2218.930 1143.490 2220.110 1144.670 ;
        RECT 2218.930 965.090 2220.110 966.270 ;
        RECT 2218.930 963.490 2220.110 964.670 ;
        RECT 2218.930 785.090 2220.110 786.270 ;
        RECT 2218.930 783.490 2220.110 784.670 ;
        RECT 2218.930 605.090 2220.110 606.270 ;
        RECT 2218.930 603.490 2220.110 604.670 ;
        RECT 2218.930 425.090 2220.110 426.270 ;
        RECT 2218.930 423.490 2220.110 424.670 ;
        RECT 2218.930 245.090 2220.110 246.270 ;
        RECT 2218.930 243.490 2220.110 244.670 ;
        RECT 2218.930 65.090 2220.110 66.270 ;
        RECT 2218.930 63.490 2220.110 64.670 ;
        RECT 2038.930 -31.110 2040.110 -29.930 ;
        RECT 2038.930 -32.710 2040.110 -31.530 ;
        RECT 2344.930 2171.090 2346.110 2172.270 ;
        RECT 2344.930 2169.490 2346.110 2170.670 ;
        RECT 2344.930 1991.090 2346.110 1992.270 ;
        RECT 2344.930 1989.490 2346.110 1990.670 ;
        RECT 2344.930 1811.090 2346.110 1812.270 ;
        RECT 2344.930 1809.490 2346.110 1810.670 ;
        RECT 2344.930 1631.090 2346.110 1632.270 ;
        RECT 2344.930 1629.490 2346.110 1630.670 ;
        RECT 2344.930 1451.090 2346.110 1452.270 ;
        RECT 2344.930 1449.490 2346.110 1450.670 ;
        RECT 2344.930 1271.090 2346.110 1272.270 ;
        RECT 2344.930 1269.490 2346.110 1270.670 ;
        RECT 2344.930 1091.090 2346.110 1092.270 ;
        RECT 2344.930 1089.490 2346.110 1090.670 ;
        RECT 2344.930 911.090 2346.110 912.270 ;
        RECT 2344.930 909.490 2346.110 910.670 ;
        RECT 2344.930 731.090 2346.110 732.270 ;
        RECT 2344.930 729.490 2346.110 730.670 ;
        RECT 2344.930 551.090 2346.110 552.270 ;
        RECT 2344.930 549.490 2346.110 550.670 ;
        RECT 2344.930 371.090 2346.110 372.270 ;
        RECT 2344.930 369.490 2346.110 370.670 ;
        RECT 2344.930 191.090 2346.110 192.270 ;
        RECT 2344.930 189.490 2346.110 190.670 ;
        RECT 2344.930 11.090 2346.110 12.270 ;
        RECT 2344.930 9.490 2346.110 10.670 ;
        RECT 2344.930 -2.910 2346.110 -1.730 ;
        RECT 2344.930 -4.510 2346.110 -3.330 ;
        RECT 2362.930 2189.090 2364.110 2190.270 ;
        RECT 2362.930 2187.490 2364.110 2188.670 ;
        RECT 2362.930 2009.090 2364.110 2010.270 ;
        RECT 2362.930 2007.490 2364.110 2008.670 ;
        RECT 2362.930 1829.090 2364.110 1830.270 ;
        RECT 2362.930 1827.490 2364.110 1828.670 ;
        RECT 2362.930 1649.090 2364.110 1650.270 ;
        RECT 2362.930 1647.490 2364.110 1648.670 ;
        RECT 2362.930 1469.090 2364.110 1470.270 ;
        RECT 2362.930 1467.490 2364.110 1468.670 ;
        RECT 2362.930 1289.090 2364.110 1290.270 ;
        RECT 2362.930 1287.490 2364.110 1288.670 ;
        RECT 2362.930 1109.090 2364.110 1110.270 ;
        RECT 2362.930 1107.490 2364.110 1108.670 ;
        RECT 2362.930 929.090 2364.110 930.270 ;
        RECT 2362.930 927.490 2364.110 928.670 ;
        RECT 2362.930 749.090 2364.110 750.270 ;
        RECT 2362.930 747.490 2364.110 748.670 ;
        RECT 2362.930 569.090 2364.110 570.270 ;
        RECT 2362.930 567.490 2364.110 568.670 ;
        RECT 2362.930 389.090 2364.110 390.270 ;
        RECT 2362.930 387.490 2364.110 388.670 ;
        RECT 2362.930 209.090 2364.110 210.270 ;
        RECT 2362.930 207.490 2364.110 208.670 ;
        RECT 2362.930 29.090 2364.110 30.270 ;
        RECT 2362.930 27.490 2364.110 28.670 ;
        RECT 2362.930 -12.310 2364.110 -11.130 ;
        RECT 2362.930 -13.910 2364.110 -12.730 ;
        RECT 2380.930 2207.090 2382.110 2208.270 ;
        RECT 2380.930 2205.490 2382.110 2206.670 ;
        RECT 2380.930 2027.090 2382.110 2028.270 ;
        RECT 2380.930 2025.490 2382.110 2026.670 ;
        RECT 2380.930 1847.090 2382.110 1848.270 ;
        RECT 2380.930 1845.490 2382.110 1846.670 ;
        RECT 2380.930 1667.090 2382.110 1668.270 ;
        RECT 2380.930 1665.490 2382.110 1666.670 ;
        RECT 2380.930 1487.090 2382.110 1488.270 ;
        RECT 2380.930 1485.490 2382.110 1486.670 ;
        RECT 2380.930 1307.090 2382.110 1308.270 ;
        RECT 2380.930 1305.490 2382.110 1306.670 ;
        RECT 2380.930 1127.090 2382.110 1128.270 ;
        RECT 2380.930 1125.490 2382.110 1126.670 ;
        RECT 2380.930 947.090 2382.110 948.270 ;
        RECT 2380.930 945.490 2382.110 946.670 ;
        RECT 2380.930 767.090 2382.110 768.270 ;
        RECT 2380.930 765.490 2382.110 766.670 ;
        RECT 2380.930 587.090 2382.110 588.270 ;
        RECT 2380.930 585.490 2382.110 586.670 ;
        RECT 2380.930 407.090 2382.110 408.270 ;
        RECT 2380.930 405.490 2382.110 406.670 ;
        RECT 2380.930 227.090 2382.110 228.270 ;
        RECT 2380.930 225.490 2382.110 226.670 ;
        RECT 2380.930 47.090 2382.110 48.270 ;
        RECT 2380.930 45.490 2382.110 46.670 ;
        RECT 2380.930 -21.710 2382.110 -20.530 ;
        RECT 2380.930 -23.310 2382.110 -22.130 ;
        RECT 2398.930 2225.090 2400.110 2226.270 ;
        RECT 2398.930 2223.490 2400.110 2224.670 ;
        RECT 2398.930 2045.090 2400.110 2046.270 ;
        RECT 2398.930 2043.490 2400.110 2044.670 ;
        RECT 2398.930 1865.090 2400.110 1866.270 ;
        RECT 2398.930 1863.490 2400.110 1864.670 ;
        RECT 2398.930 1685.090 2400.110 1686.270 ;
        RECT 2398.930 1683.490 2400.110 1684.670 ;
        RECT 2398.930 1505.090 2400.110 1506.270 ;
        RECT 2398.930 1503.490 2400.110 1504.670 ;
        RECT 2398.930 1325.090 2400.110 1326.270 ;
        RECT 2398.930 1323.490 2400.110 1324.670 ;
        RECT 2398.930 1145.090 2400.110 1146.270 ;
        RECT 2398.930 1143.490 2400.110 1144.670 ;
        RECT 2398.930 965.090 2400.110 966.270 ;
        RECT 2398.930 963.490 2400.110 964.670 ;
        RECT 2398.930 785.090 2400.110 786.270 ;
        RECT 2398.930 783.490 2400.110 784.670 ;
        RECT 2398.930 605.090 2400.110 606.270 ;
        RECT 2398.930 603.490 2400.110 604.670 ;
        RECT 2398.930 425.090 2400.110 426.270 ;
        RECT 2398.930 423.490 2400.110 424.670 ;
        RECT 2398.930 245.090 2400.110 246.270 ;
        RECT 2398.930 243.490 2400.110 244.670 ;
        RECT 2398.930 65.090 2400.110 66.270 ;
        RECT 2398.930 63.490 2400.110 64.670 ;
        RECT 2218.930 -31.110 2220.110 -29.930 ;
        RECT 2218.930 -32.710 2220.110 -31.530 ;
        RECT 2524.930 2171.090 2526.110 2172.270 ;
        RECT 2524.930 2169.490 2526.110 2170.670 ;
        RECT 2524.930 1991.090 2526.110 1992.270 ;
        RECT 2524.930 1989.490 2526.110 1990.670 ;
        RECT 2524.930 1811.090 2526.110 1812.270 ;
        RECT 2524.930 1809.490 2526.110 1810.670 ;
        RECT 2524.930 1631.090 2526.110 1632.270 ;
        RECT 2524.930 1629.490 2526.110 1630.670 ;
        RECT 2524.930 1451.090 2526.110 1452.270 ;
        RECT 2524.930 1449.490 2526.110 1450.670 ;
        RECT 2524.930 1271.090 2526.110 1272.270 ;
        RECT 2524.930 1269.490 2526.110 1270.670 ;
        RECT 2524.930 1091.090 2526.110 1092.270 ;
        RECT 2524.930 1089.490 2526.110 1090.670 ;
        RECT 2524.930 911.090 2526.110 912.270 ;
        RECT 2524.930 909.490 2526.110 910.670 ;
        RECT 2524.930 731.090 2526.110 732.270 ;
        RECT 2524.930 729.490 2526.110 730.670 ;
        RECT 2524.930 551.090 2526.110 552.270 ;
        RECT 2524.930 549.490 2526.110 550.670 ;
        RECT 2524.930 371.090 2526.110 372.270 ;
        RECT 2524.930 369.490 2526.110 370.670 ;
        RECT 2524.930 191.090 2526.110 192.270 ;
        RECT 2524.930 189.490 2526.110 190.670 ;
        RECT 2524.930 11.090 2526.110 12.270 ;
        RECT 2524.930 9.490 2526.110 10.670 ;
        RECT 2524.930 -2.910 2526.110 -1.730 ;
        RECT 2524.930 -4.510 2526.110 -3.330 ;
        RECT 2542.930 2189.090 2544.110 2190.270 ;
        RECT 2542.930 2187.490 2544.110 2188.670 ;
        RECT 2542.930 2009.090 2544.110 2010.270 ;
        RECT 2542.930 2007.490 2544.110 2008.670 ;
        RECT 2542.930 1829.090 2544.110 1830.270 ;
        RECT 2542.930 1827.490 2544.110 1828.670 ;
        RECT 2542.930 1649.090 2544.110 1650.270 ;
        RECT 2542.930 1647.490 2544.110 1648.670 ;
        RECT 2542.930 1469.090 2544.110 1470.270 ;
        RECT 2542.930 1467.490 2544.110 1468.670 ;
        RECT 2542.930 1289.090 2544.110 1290.270 ;
        RECT 2542.930 1287.490 2544.110 1288.670 ;
        RECT 2542.930 1109.090 2544.110 1110.270 ;
        RECT 2542.930 1107.490 2544.110 1108.670 ;
        RECT 2542.930 929.090 2544.110 930.270 ;
        RECT 2542.930 927.490 2544.110 928.670 ;
        RECT 2542.930 749.090 2544.110 750.270 ;
        RECT 2542.930 747.490 2544.110 748.670 ;
        RECT 2542.930 569.090 2544.110 570.270 ;
        RECT 2542.930 567.490 2544.110 568.670 ;
        RECT 2542.930 389.090 2544.110 390.270 ;
        RECT 2542.930 387.490 2544.110 388.670 ;
        RECT 2542.930 209.090 2544.110 210.270 ;
        RECT 2542.930 207.490 2544.110 208.670 ;
        RECT 2542.930 29.090 2544.110 30.270 ;
        RECT 2542.930 27.490 2544.110 28.670 ;
        RECT 2542.930 -12.310 2544.110 -11.130 ;
        RECT 2542.930 -13.910 2544.110 -12.730 ;
        RECT 2560.930 2207.090 2562.110 2208.270 ;
        RECT 2560.930 2205.490 2562.110 2206.670 ;
        RECT 2560.930 2027.090 2562.110 2028.270 ;
        RECT 2560.930 2025.490 2562.110 2026.670 ;
        RECT 2560.930 1847.090 2562.110 1848.270 ;
        RECT 2560.930 1845.490 2562.110 1846.670 ;
        RECT 2560.930 1667.090 2562.110 1668.270 ;
        RECT 2560.930 1665.490 2562.110 1666.670 ;
        RECT 2560.930 1487.090 2562.110 1488.270 ;
        RECT 2560.930 1485.490 2562.110 1486.670 ;
        RECT 2560.930 1307.090 2562.110 1308.270 ;
        RECT 2560.930 1305.490 2562.110 1306.670 ;
        RECT 2560.930 1127.090 2562.110 1128.270 ;
        RECT 2560.930 1125.490 2562.110 1126.670 ;
        RECT 2560.930 947.090 2562.110 948.270 ;
        RECT 2560.930 945.490 2562.110 946.670 ;
        RECT 2560.930 767.090 2562.110 768.270 ;
        RECT 2560.930 765.490 2562.110 766.670 ;
        RECT 2560.930 587.090 2562.110 588.270 ;
        RECT 2560.930 585.490 2562.110 586.670 ;
        RECT 2560.930 407.090 2562.110 408.270 ;
        RECT 2560.930 405.490 2562.110 406.670 ;
        RECT 2560.930 227.090 2562.110 228.270 ;
        RECT 2560.930 225.490 2562.110 226.670 ;
        RECT 2560.930 47.090 2562.110 48.270 ;
        RECT 2560.930 45.490 2562.110 46.670 ;
        RECT 2560.930 -21.710 2562.110 -20.530 ;
        RECT 2560.930 -23.310 2562.110 -22.130 ;
        RECT 2578.930 2225.090 2580.110 2226.270 ;
        RECT 2578.930 2223.490 2580.110 2224.670 ;
        RECT 2578.930 2045.090 2580.110 2046.270 ;
        RECT 2578.930 2043.490 2580.110 2044.670 ;
        RECT 2578.930 1865.090 2580.110 1866.270 ;
        RECT 2578.930 1863.490 2580.110 1864.670 ;
        RECT 2578.930 1685.090 2580.110 1686.270 ;
        RECT 2578.930 1683.490 2580.110 1684.670 ;
        RECT 2578.930 1505.090 2580.110 1506.270 ;
        RECT 2578.930 1503.490 2580.110 1504.670 ;
        RECT 2578.930 1325.090 2580.110 1326.270 ;
        RECT 2578.930 1323.490 2580.110 1324.670 ;
        RECT 2578.930 1145.090 2580.110 1146.270 ;
        RECT 2578.930 1143.490 2580.110 1144.670 ;
        RECT 2578.930 965.090 2580.110 966.270 ;
        RECT 2578.930 963.490 2580.110 964.670 ;
        RECT 2578.930 785.090 2580.110 786.270 ;
        RECT 2578.930 783.490 2580.110 784.670 ;
        RECT 2578.930 605.090 2580.110 606.270 ;
        RECT 2578.930 603.490 2580.110 604.670 ;
        RECT 2578.930 425.090 2580.110 426.270 ;
        RECT 2578.930 423.490 2580.110 424.670 ;
        RECT 2578.930 245.090 2580.110 246.270 ;
        RECT 2578.930 243.490 2580.110 244.670 ;
        RECT 2578.930 65.090 2580.110 66.270 ;
        RECT 2578.930 63.490 2580.110 64.670 ;
        RECT 2398.930 -31.110 2400.110 -29.930 ;
        RECT 2398.930 -32.710 2400.110 -31.530 ;
        RECT 2704.930 2171.090 2706.110 2172.270 ;
        RECT 2704.930 2169.490 2706.110 2170.670 ;
        RECT 2704.930 1991.090 2706.110 1992.270 ;
        RECT 2704.930 1989.490 2706.110 1990.670 ;
        RECT 2704.930 1811.090 2706.110 1812.270 ;
        RECT 2704.930 1809.490 2706.110 1810.670 ;
        RECT 2704.930 1631.090 2706.110 1632.270 ;
        RECT 2704.930 1629.490 2706.110 1630.670 ;
        RECT 2704.930 1451.090 2706.110 1452.270 ;
        RECT 2704.930 1449.490 2706.110 1450.670 ;
        RECT 2704.930 1271.090 2706.110 1272.270 ;
        RECT 2704.930 1269.490 2706.110 1270.670 ;
        RECT 2704.930 1091.090 2706.110 1092.270 ;
        RECT 2704.930 1089.490 2706.110 1090.670 ;
        RECT 2704.930 911.090 2706.110 912.270 ;
        RECT 2704.930 909.490 2706.110 910.670 ;
        RECT 2704.930 731.090 2706.110 732.270 ;
        RECT 2704.930 729.490 2706.110 730.670 ;
        RECT 2704.930 551.090 2706.110 552.270 ;
        RECT 2704.930 549.490 2706.110 550.670 ;
        RECT 2704.930 371.090 2706.110 372.270 ;
        RECT 2704.930 369.490 2706.110 370.670 ;
        RECT 2704.930 191.090 2706.110 192.270 ;
        RECT 2704.930 189.490 2706.110 190.670 ;
        RECT 2704.930 11.090 2706.110 12.270 ;
        RECT 2704.930 9.490 2706.110 10.670 ;
        RECT 2704.930 -2.910 2706.110 -1.730 ;
        RECT 2704.930 -4.510 2706.110 -3.330 ;
        RECT 2722.930 3449.090 2724.110 3450.270 ;
        RECT 2722.930 3447.490 2724.110 3448.670 ;
        RECT 2722.930 3269.090 2724.110 3270.270 ;
        RECT 2722.930 3267.490 2724.110 3268.670 ;
        RECT 2722.930 3089.090 2724.110 3090.270 ;
        RECT 2722.930 3087.490 2724.110 3088.670 ;
        RECT 2722.930 2909.090 2724.110 2910.270 ;
        RECT 2722.930 2907.490 2724.110 2908.670 ;
        RECT 2722.930 2729.090 2724.110 2730.270 ;
        RECT 2722.930 2727.490 2724.110 2728.670 ;
        RECT 2722.930 2549.090 2724.110 2550.270 ;
        RECT 2722.930 2547.490 2724.110 2548.670 ;
        RECT 2722.930 2369.090 2724.110 2370.270 ;
        RECT 2722.930 2367.490 2724.110 2368.670 ;
        RECT 2722.930 2189.090 2724.110 2190.270 ;
        RECT 2722.930 2187.490 2724.110 2188.670 ;
        RECT 2722.930 2009.090 2724.110 2010.270 ;
        RECT 2722.930 2007.490 2724.110 2008.670 ;
        RECT 2722.930 1829.090 2724.110 1830.270 ;
        RECT 2722.930 1827.490 2724.110 1828.670 ;
        RECT 2722.930 1649.090 2724.110 1650.270 ;
        RECT 2722.930 1647.490 2724.110 1648.670 ;
        RECT 2722.930 1469.090 2724.110 1470.270 ;
        RECT 2722.930 1467.490 2724.110 1468.670 ;
        RECT 2722.930 1289.090 2724.110 1290.270 ;
        RECT 2722.930 1287.490 2724.110 1288.670 ;
        RECT 2722.930 1109.090 2724.110 1110.270 ;
        RECT 2722.930 1107.490 2724.110 1108.670 ;
        RECT 2722.930 929.090 2724.110 930.270 ;
        RECT 2722.930 927.490 2724.110 928.670 ;
        RECT 2722.930 749.090 2724.110 750.270 ;
        RECT 2722.930 747.490 2724.110 748.670 ;
        RECT 2722.930 569.090 2724.110 570.270 ;
        RECT 2722.930 567.490 2724.110 568.670 ;
        RECT 2722.930 389.090 2724.110 390.270 ;
        RECT 2722.930 387.490 2724.110 388.670 ;
        RECT 2722.930 209.090 2724.110 210.270 ;
        RECT 2722.930 207.490 2724.110 208.670 ;
        RECT 2722.930 29.090 2724.110 30.270 ;
        RECT 2722.930 27.490 2724.110 28.670 ;
        RECT 2722.930 -12.310 2724.110 -11.130 ;
        RECT 2722.930 -13.910 2724.110 -12.730 ;
        RECT 2740.930 3467.090 2742.110 3468.270 ;
        RECT 2740.930 3465.490 2742.110 3466.670 ;
        RECT 2740.930 3287.090 2742.110 3288.270 ;
        RECT 2740.930 3285.490 2742.110 3286.670 ;
        RECT 2740.930 3107.090 2742.110 3108.270 ;
        RECT 2740.930 3105.490 2742.110 3106.670 ;
        RECT 2740.930 2927.090 2742.110 2928.270 ;
        RECT 2740.930 2925.490 2742.110 2926.670 ;
        RECT 2740.930 2747.090 2742.110 2748.270 ;
        RECT 2740.930 2745.490 2742.110 2746.670 ;
        RECT 2740.930 2567.090 2742.110 2568.270 ;
        RECT 2740.930 2565.490 2742.110 2566.670 ;
        RECT 2740.930 2387.090 2742.110 2388.270 ;
        RECT 2740.930 2385.490 2742.110 2386.670 ;
        RECT 2740.930 2207.090 2742.110 2208.270 ;
        RECT 2740.930 2205.490 2742.110 2206.670 ;
        RECT 2740.930 2027.090 2742.110 2028.270 ;
        RECT 2740.930 2025.490 2742.110 2026.670 ;
        RECT 2740.930 1847.090 2742.110 1848.270 ;
        RECT 2740.930 1845.490 2742.110 1846.670 ;
        RECT 2740.930 1667.090 2742.110 1668.270 ;
        RECT 2740.930 1665.490 2742.110 1666.670 ;
        RECT 2740.930 1487.090 2742.110 1488.270 ;
        RECT 2740.930 1485.490 2742.110 1486.670 ;
        RECT 2740.930 1307.090 2742.110 1308.270 ;
        RECT 2740.930 1305.490 2742.110 1306.670 ;
        RECT 2740.930 1127.090 2742.110 1128.270 ;
        RECT 2740.930 1125.490 2742.110 1126.670 ;
        RECT 2740.930 947.090 2742.110 948.270 ;
        RECT 2740.930 945.490 2742.110 946.670 ;
        RECT 2740.930 767.090 2742.110 768.270 ;
        RECT 2740.930 765.490 2742.110 766.670 ;
        RECT 2740.930 587.090 2742.110 588.270 ;
        RECT 2740.930 585.490 2742.110 586.670 ;
        RECT 2740.930 407.090 2742.110 408.270 ;
        RECT 2740.930 405.490 2742.110 406.670 ;
        RECT 2740.930 227.090 2742.110 228.270 ;
        RECT 2740.930 225.490 2742.110 226.670 ;
        RECT 2740.930 47.090 2742.110 48.270 ;
        RECT 2740.930 45.490 2742.110 46.670 ;
        RECT 2740.930 -21.710 2742.110 -20.530 ;
        RECT 2740.930 -23.310 2742.110 -22.130 ;
        RECT 2955.710 3551.210 2956.890 3552.390 ;
        RECT 2955.710 3549.610 2956.890 3550.790 ;
        RECT 2946.310 3541.810 2947.490 3542.990 ;
        RECT 2946.310 3540.210 2947.490 3541.390 ;
        RECT 2902.930 3532.410 2904.110 3533.590 ;
        RECT 2902.930 3530.810 2904.110 3531.990 ;
        RECT 2758.930 3485.090 2760.110 3486.270 ;
        RECT 2758.930 3483.490 2760.110 3484.670 ;
        RECT 2758.930 3305.090 2760.110 3306.270 ;
        RECT 2758.930 3303.490 2760.110 3304.670 ;
        RECT 2758.930 3125.090 2760.110 3126.270 ;
        RECT 2758.930 3123.490 2760.110 3124.670 ;
        RECT 2758.930 2945.090 2760.110 2946.270 ;
        RECT 2758.930 2943.490 2760.110 2944.670 ;
        RECT 2758.930 2765.090 2760.110 2766.270 ;
        RECT 2758.930 2763.490 2760.110 2764.670 ;
        RECT 2758.930 2585.090 2760.110 2586.270 ;
        RECT 2758.930 2583.490 2760.110 2584.670 ;
        RECT 2758.930 2405.090 2760.110 2406.270 ;
        RECT 2758.930 2403.490 2760.110 2404.670 ;
        RECT 2758.930 2225.090 2760.110 2226.270 ;
        RECT 2758.930 2223.490 2760.110 2224.670 ;
        RECT 2758.930 2045.090 2760.110 2046.270 ;
        RECT 2758.930 2043.490 2760.110 2044.670 ;
        RECT 2758.930 1865.090 2760.110 1866.270 ;
        RECT 2758.930 1863.490 2760.110 1864.670 ;
        RECT 2758.930 1685.090 2760.110 1686.270 ;
        RECT 2758.930 1683.490 2760.110 1684.670 ;
        RECT 2758.930 1505.090 2760.110 1506.270 ;
        RECT 2758.930 1503.490 2760.110 1504.670 ;
        RECT 2758.930 1325.090 2760.110 1326.270 ;
        RECT 2758.930 1323.490 2760.110 1324.670 ;
        RECT 2758.930 1145.090 2760.110 1146.270 ;
        RECT 2758.930 1143.490 2760.110 1144.670 ;
        RECT 2758.930 965.090 2760.110 966.270 ;
        RECT 2758.930 963.490 2760.110 964.670 ;
        RECT 2758.930 785.090 2760.110 786.270 ;
        RECT 2758.930 783.490 2760.110 784.670 ;
        RECT 2758.930 605.090 2760.110 606.270 ;
        RECT 2758.930 603.490 2760.110 604.670 ;
        RECT 2758.930 425.090 2760.110 426.270 ;
        RECT 2758.930 423.490 2760.110 424.670 ;
        RECT 2758.930 245.090 2760.110 246.270 ;
        RECT 2758.930 243.490 2760.110 244.670 ;
        RECT 2758.930 65.090 2760.110 66.270 ;
        RECT 2758.930 63.490 2760.110 64.670 ;
        RECT 2578.930 -31.110 2580.110 -29.930 ;
        RECT 2578.930 -32.710 2580.110 -31.530 ;
        RECT 2884.930 3523.010 2886.110 3524.190 ;
        RECT 2884.930 3521.410 2886.110 3522.590 ;
        RECT 2884.930 3431.090 2886.110 3432.270 ;
        RECT 2884.930 3429.490 2886.110 3430.670 ;
        RECT 2884.930 3251.090 2886.110 3252.270 ;
        RECT 2884.930 3249.490 2886.110 3250.670 ;
        RECT 2884.930 3071.090 2886.110 3072.270 ;
        RECT 2884.930 3069.490 2886.110 3070.670 ;
        RECT 2884.930 2891.090 2886.110 2892.270 ;
        RECT 2884.930 2889.490 2886.110 2890.670 ;
        RECT 2884.930 2711.090 2886.110 2712.270 ;
        RECT 2884.930 2709.490 2886.110 2710.670 ;
        RECT 2884.930 2531.090 2886.110 2532.270 ;
        RECT 2884.930 2529.490 2886.110 2530.670 ;
        RECT 2884.930 2351.090 2886.110 2352.270 ;
        RECT 2884.930 2349.490 2886.110 2350.670 ;
        RECT 2884.930 2171.090 2886.110 2172.270 ;
        RECT 2884.930 2169.490 2886.110 2170.670 ;
        RECT 2884.930 1991.090 2886.110 1992.270 ;
        RECT 2884.930 1989.490 2886.110 1990.670 ;
        RECT 2884.930 1811.090 2886.110 1812.270 ;
        RECT 2884.930 1809.490 2886.110 1810.670 ;
        RECT 2884.930 1631.090 2886.110 1632.270 ;
        RECT 2884.930 1629.490 2886.110 1630.670 ;
        RECT 2884.930 1451.090 2886.110 1452.270 ;
        RECT 2884.930 1449.490 2886.110 1450.670 ;
        RECT 2884.930 1271.090 2886.110 1272.270 ;
        RECT 2884.930 1269.490 2886.110 1270.670 ;
        RECT 2884.930 1091.090 2886.110 1092.270 ;
        RECT 2884.930 1089.490 2886.110 1090.670 ;
        RECT 2884.930 911.090 2886.110 912.270 ;
        RECT 2884.930 909.490 2886.110 910.670 ;
        RECT 2884.930 731.090 2886.110 732.270 ;
        RECT 2884.930 729.490 2886.110 730.670 ;
        RECT 2884.930 551.090 2886.110 552.270 ;
        RECT 2884.930 549.490 2886.110 550.670 ;
        RECT 2884.930 371.090 2886.110 372.270 ;
        RECT 2884.930 369.490 2886.110 370.670 ;
        RECT 2884.930 191.090 2886.110 192.270 ;
        RECT 2884.930 189.490 2886.110 190.670 ;
        RECT 2884.930 11.090 2886.110 12.270 ;
        RECT 2884.930 9.490 2886.110 10.670 ;
        RECT 2884.930 -2.910 2886.110 -1.730 ;
        RECT 2884.930 -4.510 2886.110 -3.330 ;
        RECT 2936.910 3532.410 2938.090 3533.590 ;
        RECT 2936.910 3530.810 2938.090 3531.990 ;
        RECT 2902.930 3449.090 2904.110 3450.270 ;
        RECT 2902.930 3447.490 2904.110 3448.670 ;
        RECT 2902.930 3269.090 2904.110 3270.270 ;
        RECT 2902.930 3267.490 2904.110 3268.670 ;
        RECT 2902.930 3089.090 2904.110 3090.270 ;
        RECT 2902.930 3087.490 2904.110 3088.670 ;
        RECT 2902.930 2909.090 2904.110 2910.270 ;
        RECT 2902.930 2907.490 2904.110 2908.670 ;
        RECT 2902.930 2729.090 2904.110 2730.270 ;
        RECT 2902.930 2727.490 2904.110 2728.670 ;
        RECT 2902.930 2549.090 2904.110 2550.270 ;
        RECT 2902.930 2547.490 2904.110 2548.670 ;
        RECT 2902.930 2369.090 2904.110 2370.270 ;
        RECT 2902.930 2367.490 2904.110 2368.670 ;
        RECT 2902.930 2189.090 2904.110 2190.270 ;
        RECT 2902.930 2187.490 2904.110 2188.670 ;
        RECT 2902.930 2009.090 2904.110 2010.270 ;
        RECT 2902.930 2007.490 2904.110 2008.670 ;
        RECT 2902.930 1829.090 2904.110 1830.270 ;
        RECT 2902.930 1827.490 2904.110 1828.670 ;
        RECT 2902.930 1649.090 2904.110 1650.270 ;
        RECT 2902.930 1647.490 2904.110 1648.670 ;
        RECT 2902.930 1469.090 2904.110 1470.270 ;
        RECT 2902.930 1467.490 2904.110 1468.670 ;
        RECT 2902.930 1289.090 2904.110 1290.270 ;
        RECT 2902.930 1287.490 2904.110 1288.670 ;
        RECT 2902.930 1109.090 2904.110 1110.270 ;
        RECT 2902.930 1107.490 2904.110 1108.670 ;
        RECT 2902.930 929.090 2904.110 930.270 ;
        RECT 2902.930 927.490 2904.110 928.670 ;
        RECT 2902.930 749.090 2904.110 750.270 ;
        RECT 2902.930 747.490 2904.110 748.670 ;
        RECT 2902.930 569.090 2904.110 570.270 ;
        RECT 2902.930 567.490 2904.110 568.670 ;
        RECT 2902.930 389.090 2904.110 390.270 ;
        RECT 2902.930 387.490 2904.110 388.670 ;
        RECT 2902.930 209.090 2904.110 210.270 ;
        RECT 2902.930 207.490 2904.110 208.670 ;
        RECT 2902.930 29.090 2904.110 30.270 ;
        RECT 2902.930 27.490 2904.110 28.670 ;
        RECT 2927.510 3523.010 2928.690 3524.190 ;
        RECT 2927.510 3521.410 2928.690 3522.590 ;
        RECT 2927.510 3431.090 2928.690 3432.270 ;
        RECT 2927.510 3429.490 2928.690 3430.670 ;
        RECT 2927.510 3251.090 2928.690 3252.270 ;
        RECT 2927.510 3249.490 2928.690 3250.670 ;
        RECT 2927.510 3071.090 2928.690 3072.270 ;
        RECT 2927.510 3069.490 2928.690 3070.670 ;
        RECT 2927.510 2891.090 2928.690 2892.270 ;
        RECT 2927.510 2889.490 2928.690 2890.670 ;
        RECT 2927.510 2711.090 2928.690 2712.270 ;
        RECT 2927.510 2709.490 2928.690 2710.670 ;
        RECT 2927.510 2531.090 2928.690 2532.270 ;
        RECT 2927.510 2529.490 2928.690 2530.670 ;
        RECT 2927.510 2351.090 2928.690 2352.270 ;
        RECT 2927.510 2349.490 2928.690 2350.670 ;
        RECT 2927.510 2171.090 2928.690 2172.270 ;
        RECT 2927.510 2169.490 2928.690 2170.670 ;
        RECT 2927.510 1991.090 2928.690 1992.270 ;
        RECT 2927.510 1989.490 2928.690 1990.670 ;
        RECT 2927.510 1811.090 2928.690 1812.270 ;
        RECT 2927.510 1809.490 2928.690 1810.670 ;
        RECT 2927.510 1631.090 2928.690 1632.270 ;
        RECT 2927.510 1629.490 2928.690 1630.670 ;
        RECT 2927.510 1451.090 2928.690 1452.270 ;
        RECT 2927.510 1449.490 2928.690 1450.670 ;
        RECT 2927.510 1271.090 2928.690 1272.270 ;
        RECT 2927.510 1269.490 2928.690 1270.670 ;
        RECT 2927.510 1091.090 2928.690 1092.270 ;
        RECT 2927.510 1089.490 2928.690 1090.670 ;
        RECT 2927.510 911.090 2928.690 912.270 ;
        RECT 2927.510 909.490 2928.690 910.670 ;
        RECT 2927.510 731.090 2928.690 732.270 ;
        RECT 2927.510 729.490 2928.690 730.670 ;
        RECT 2927.510 551.090 2928.690 552.270 ;
        RECT 2927.510 549.490 2928.690 550.670 ;
        RECT 2927.510 371.090 2928.690 372.270 ;
        RECT 2927.510 369.490 2928.690 370.670 ;
        RECT 2927.510 191.090 2928.690 192.270 ;
        RECT 2927.510 189.490 2928.690 190.670 ;
        RECT 2927.510 11.090 2928.690 12.270 ;
        RECT 2927.510 9.490 2928.690 10.670 ;
        RECT 2927.510 -2.910 2928.690 -1.730 ;
        RECT 2927.510 -4.510 2928.690 -3.330 ;
        RECT 2936.910 3449.090 2938.090 3450.270 ;
        RECT 2936.910 3447.490 2938.090 3448.670 ;
        RECT 2936.910 3269.090 2938.090 3270.270 ;
        RECT 2936.910 3267.490 2938.090 3268.670 ;
        RECT 2936.910 3089.090 2938.090 3090.270 ;
        RECT 2936.910 3087.490 2938.090 3088.670 ;
        RECT 2936.910 2909.090 2938.090 2910.270 ;
        RECT 2936.910 2907.490 2938.090 2908.670 ;
        RECT 2936.910 2729.090 2938.090 2730.270 ;
        RECT 2936.910 2727.490 2938.090 2728.670 ;
        RECT 2936.910 2549.090 2938.090 2550.270 ;
        RECT 2936.910 2547.490 2938.090 2548.670 ;
        RECT 2936.910 2369.090 2938.090 2370.270 ;
        RECT 2936.910 2367.490 2938.090 2368.670 ;
        RECT 2936.910 2189.090 2938.090 2190.270 ;
        RECT 2936.910 2187.490 2938.090 2188.670 ;
        RECT 2936.910 2009.090 2938.090 2010.270 ;
        RECT 2936.910 2007.490 2938.090 2008.670 ;
        RECT 2936.910 1829.090 2938.090 1830.270 ;
        RECT 2936.910 1827.490 2938.090 1828.670 ;
        RECT 2936.910 1649.090 2938.090 1650.270 ;
        RECT 2936.910 1647.490 2938.090 1648.670 ;
        RECT 2936.910 1469.090 2938.090 1470.270 ;
        RECT 2936.910 1467.490 2938.090 1468.670 ;
        RECT 2936.910 1289.090 2938.090 1290.270 ;
        RECT 2936.910 1287.490 2938.090 1288.670 ;
        RECT 2936.910 1109.090 2938.090 1110.270 ;
        RECT 2936.910 1107.490 2938.090 1108.670 ;
        RECT 2936.910 929.090 2938.090 930.270 ;
        RECT 2936.910 927.490 2938.090 928.670 ;
        RECT 2936.910 749.090 2938.090 750.270 ;
        RECT 2936.910 747.490 2938.090 748.670 ;
        RECT 2936.910 569.090 2938.090 570.270 ;
        RECT 2936.910 567.490 2938.090 568.670 ;
        RECT 2936.910 389.090 2938.090 390.270 ;
        RECT 2936.910 387.490 2938.090 388.670 ;
        RECT 2936.910 209.090 2938.090 210.270 ;
        RECT 2936.910 207.490 2938.090 208.670 ;
        RECT 2936.910 29.090 2938.090 30.270 ;
        RECT 2936.910 27.490 2938.090 28.670 ;
        RECT 2902.930 -12.310 2904.110 -11.130 ;
        RECT 2902.930 -13.910 2904.110 -12.730 ;
        RECT 2936.910 -12.310 2938.090 -11.130 ;
        RECT 2936.910 -13.910 2938.090 -12.730 ;
        RECT 2946.310 3467.090 2947.490 3468.270 ;
        RECT 2946.310 3465.490 2947.490 3466.670 ;
        RECT 2946.310 3287.090 2947.490 3288.270 ;
        RECT 2946.310 3285.490 2947.490 3286.670 ;
        RECT 2946.310 3107.090 2947.490 3108.270 ;
        RECT 2946.310 3105.490 2947.490 3106.670 ;
        RECT 2946.310 2927.090 2947.490 2928.270 ;
        RECT 2946.310 2925.490 2947.490 2926.670 ;
        RECT 2946.310 2747.090 2947.490 2748.270 ;
        RECT 2946.310 2745.490 2947.490 2746.670 ;
        RECT 2946.310 2567.090 2947.490 2568.270 ;
        RECT 2946.310 2565.490 2947.490 2566.670 ;
        RECT 2946.310 2387.090 2947.490 2388.270 ;
        RECT 2946.310 2385.490 2947.490 2386.670 ;
        RECT 2946.310 2207.090 2947.490 2208.270 ;
        RECT 2946.310 2205.490 2947.490 2206.670 ;
        RECT 2946.310 2027.090 2947.490 2028.270 ;
        RECT 2946.310 2025.490 2947.490 2026.670 ;
        RECT 2946.310 1847.090 2947.490 1848.270 ;
        RECT 2946.310 1845.490 2947.490 1846.670 ;
        RECT 2946.310 1667.090 2947.490 1668.270 ;
        RECT 2946.310 1665.490 2947.490 1666.670 ;
        RECT 2946.310 1487.090 2947.490 1488.270 ;
        RECT 2946.310 1485.490 2947.490 1486.670 ;
        RECT 2946.310 1307.090 2947.490 1308.270 ;
        RECT 2946.310 1305.490 2947.490 1306.670 ;
        RECT 2946.310 1127.090 2947.490 1128.270 ;
        RECT 2946.310 1125.490 2947.490 1126.670 ;
        RECT 2946.310 947.090 2947.490 948.270 ;
        RECT 2946.310 945.490 2947.490 946.670 ;
        RECT 2946.310 767.090 2947.490 768.270 ;
        RECT 2946.310 765.490 2947.490 766.670 ;
        RECT 2946.310 587.090 2947.490 588.270 ;
        RECT 2946.310 585.490 2947.490 586.670 ;
        RECT 2946.310 407.090 2947.490 408.270 ;
        RECT 2946.310 405.490 2947.490 406.670 ;
        RECT 2946.310 227.090 2947.490 228.270 ;
        RECT 2946.310 225.490 2947.490 226.670 ;
        RECT 2946.310 47.090 2947.490 48.270 ;
        RECT 2946.310 45.490 2947.490 46.670 ;
        RECT 2946.310 -21.710 2947.490 -20.530 ;
        RECT 2946.310 -23.310 2947.490 -22.130 ;
        RECT 2955.710 3485.090 2956.890 3486.270 ;
        RECT 2955.710 3483.490 2956.890 3484.670 ;
        RECT 2955.710 3305.090 2956.890 3306.270 ;
        RECT 2955.710 3303.490 2956.890 3304.670 ;
        RECT 2955.710 3125.090 2956.890 3126.270 ;
        RECT 2955.710 3123.490 2956.890 3124.670 ;
        RECT 2955.710 2945.090 2956.890 2946.270 ;
        RECT 2955.710 2943.490 2956.890 2944.670 ;
        RECT 2955.710 2765.090 2956.890 2766.270 ;
        RECT 2955.710 2763.490 2956.890 2764.670 ;
        RECT 2955.710 2585.090 2956.890 2586.270 ;
        RECT 2955.710 2583.490 2956.890 2584.670 ;
        RECT 2955.710 2405.090 2956.890 2406.270 ;
        RECT 2955.710 2403.490 2956.890 2404.670 ;
        RECT 2955.710 2225.090 2956.890 2226.270 ;
        RECT 2955.710 2223.490 2956.890 2224.670 ;
        RECT 2955.710 2045.090 2956.890 2046.270 ;
        RECT 2955.710 2043.490 2956.890 2044.670 ;
        RECT 2955.710 1865.090 2956.890 1866.270 ;
        RECT 2955.710 1863.490 2956.890 1864.670 ;
        RECT 2955.710 1685.090 2956.890 1686.270 ;
        RECT 2955.710 1683.490 2956.890 1684.670 ;
        RECT 2955.710 1505.090 2956.890 1506.270 ;
        RECT 2955.710 1503.490 2956.890 1504.670 ;
        RECT 2955.710 1325.090 2956.890 1326.270 ;
        RECT 2955.710 1323.490 2956.890 1324.670 ;
        RECT 2955.710 1145.090 2956.890 1146.270 ;
        RECT 2955.710 1143.490 2956.890 1144.670 ;
        RECT 2955.710 965.090 2956.890 966.270 ;
        RECT 2955.710 963.490 2956.890 964.670 ;
        RECT 2955.710 785.090 2956.890 786.270 ;
        RECT 2955.710 783.490 2956.890 784.670 ;
        RECT 2955.710 605.090 2956.890 606.270 ;
        RECT 2955.710 603.490 2956.890 604.670 ;
        RECT 2955.710 425.090 2956.890 426.270 ;
        RECT 2955.710 423.490 2956.890 424.670 ;
        RECT 2955.710 245.090 2956.890 246.270 ;
        RECT 2955.710 243.490 2956.890 244.670 ;
        RECT 2955.710 65.090 2956.890 66.270 ;
        RECT 2955.710 63.490 2956.890 64.670 ;
        RECT 2758.930 -31.110 2760.110 -29.930 ;
        RECT 2758.930 -32.710 2760.110 -31.530 ;
        RECT 2955.710 -31.110 2956.890 -29.930 ;
        RECT 2955.710 -32.710 2956.890 -31.530 ;
      LAYER met5 ;
        RECT -38.180 3552.500 -35.180 3552.510 ;
        RECT 58.020 3552.500 61.020 3552.510 ;
        RECT 238.020 3552.500 241.020 3552.510 ;
        RECT 418.020 3552.500 421.020 3552.510 ;
        RECT 598.020 3552.500 601.020 3552.510 ;
        RECT 778.020 3552.500 781.020 3552.510 ;
        RECT 958.020 3552.500 961.020 3552.510 ;
        RECT 1138.020 3552.500 1141.020 3552.510 ;
        RECT 1318.020 3552.500 1321.020 3552.510 ;
        RECT 1498.020 3552.500 1501.020 3552.510 ;
        RECT 1678.020 3552.500 1681.020 3552.510 ;
        RECT 1858.020 3552.500 1861.020 3552.510 ;
        RECT 2038.020 3552.500 2041.020 3552.510 ;
        RECT 2218.020 3552.500 2221.020 3552.510 ;
        RECT 2398.020 3552.500 2401.020 3552.510 ;
        RECT 2578.020 3552.500 2581.020 3552.510 ;
        RECT 2758.020 3552.500 2761.020 3552.510 ;
        RECT 2954.800 3552.500 2957.800 3552.510 ;
        RECT -38.180 3549.500 2957.800 3552.500 ;
        RECT -38.180 3549.490 -35.180 3549.500 ;
        RECT 58.020 3549.490 61.020 3549.500 ;
        RECT 238.020 3549.490 241.020 3549.500 ;
        RECT 418.020 3549.490 421.020 3549.500 ;
        RECT 598.020 3549.490 601.020 3549.500 ;
        RECT 778.020 3549.490 781.020 3549.500 ;
        RECT 958.020 3549.490 961.020 3549.500 ;
        RECT 1138.020 3549.490 1141.020 3549.500 ;
        RECT 1318.020 3549.490 1321.020 3549.500 ;
        RECT 1498.020 3549.490 1501.020 3549.500 ;
        RECT 1678.020 3549.490 1681.020 3549.500 ;
        RECT 1858.020 3549.490 1861.020 3549.500 ;
        RECT 2038.020 3549.490 2041.020 3549.500 ;
        RECT 2218.020 3549.490 2221.020 3549.500 ;
        RECT 2398.020 3549.490 2401.020 3549.500 ;
        RECT 2578.020 3549.490 2581.020 3549.500 ;
        RECT 2758.020 3549.490 2761.020 3549.500 ;
        RECT 2954.800 3549.490 2957.800 3549.500 ;
        RECT -28.780 3543.100 -25.780 3543.110 ;
        RECT 40.020 3543.100 43.020 3543.110 ;
        RECT 220.020 3543.100 223.020 3543.110 ;
        RECT 400.020 3543.100 403.020 3543.110 ;
        RECT 580.020 3543.100 583.020 3543.110 ;
        RECT 760.020 3543.100 763.020 3543.110 ;
        RECT 940.020 3543.100 943.020 3543.110 ;
        RECT 1120.020 3543.100 1123.020 3543.110 ;
        RECT 1300.020 3543.100 1303.020 3543.110 ;
        RECT 1480.020 3543.100 1483.020 3543.110 ;
        RECT 1660.020 3543.100 1663.020 3543.110 ;
        RECT 1840.020 3543.100 1843.020 3543.110 ;
        RECT 2020.020 3543.100 2023.020 3543.110 ;
        RECT 2200.020 3543.100 2203.020 3543.110 ;
        RECT 2380.020 3543.100 2383.020 3543.110 ;
        RECT 2560.020 3543.100 2563.020 3543.110 ;
        RECT 2740.020 3543.100 2743.020 3543.110 ;
        RECT 2945.400 3543.100 2948.400 3543.110 ;
        RECT -28.780 3540.100 2948.400 3543.100 ;
        RECT -28.780 3540.090 -25.780 3540.100 ;
        RECT 40.020 3540.090 43.020 3540.100 ;
        RECT 220.020 3540.090 223.020 3540.100 ;
        RECT 400.020 3540.090 403.020 3540.100 ;
        RECT 580.020 3540.090 583.020 3540.100 ;
        RECT 760.020 3540.090 763.020 3540.100 ;
        RECT 940.020 3540.090 943.020 3540.100 ;
        RECT 1120.020 3540.090 1123.020 3540.100 ;
        RECT 1300.020 3540.090 1303.020 3540.100 ;
        RECT 1480.020 3540.090 1483.020 3540.100 ;
        RECT 1660.020 3540.090 1663.020 3540.100 ;
        RECT 1840.020 3540.090 1843.020 3540.100 ;
        RECT 2020.020 3540.090 2023.020 3540.100 ;
        RECT 2200.020 3540.090 2203.020 3540.100 ;
        RECT 2380.020 3540.090 2383.020 3540.100 ;
        RECT 2560.020 3540.090 2563.020 3540.100 ;
        RECT 2740.020 3540.090 2743.020 3540.100 ;
        RECT 2945.400 3540.090 2948.400 3540.100 ;
        RECT -19.380 3533.700 -16.380 3533.710 ;
        RECT 22.020 3533.700 25.020 3533.710 ;
        RECT 202.020 3533.700 205.020 3533.710 ;
        RECT 382.020 3533.700 385.020 3533.710 ;
        RECT 562.020 3533.700 565.020 3533.710 ;
        RECT 742.020 3533.700 745.020 3533.710 ;
        RECT 922.020 3533.700 925.020 3533.710 ;
        RECT 1102.020 3533.700 1105.020 3533.710 ;
        RECT 1282.020 3533.700 1285.020 3533.710 ;
        RECT 1462.020 3533.700 1465.020 3533.710 ;
        RECT 1642.020 3533.700 1645.020 3533.710 ;
        RECT 1822.020 3533.700 1825.020 3533.710 ;
        RECT 2002.020 3533.700 2005.020 3533.710 ;
        RECT 2182.020 3533.700 2185.020 3533.710 ;
        RECT 2362.020 3533.700 2365.020 3533.710 ;
        RECT 2542.020 3533.700 2545.020 3533.710 ;
        RECT 2722.020 3533.700 2725.020 3533.710 ;
        RECT 2902.020 3533.700 2905.020 3533.710 ;
        RECT 2936.000 3533.700 2939.000 3533.710 ;
        RECT -19.380 3530.700 2939.000 3533.700 ;
        RECT -19.380 3530.690 -16.380 3530.700 ;
        RECT 22.020 3530.690 25.020 3530.700 ;
        RECT 202.020 3530.690 205.020 3530.700 ;
        RECT 382.020 3530.690 385.020 3530.700 ;
        RECT 562.020 3530.690 565.020 3530.700 ;
        RECT 742.020 3530.690 745.020 3530.700 ;
        RECT 922.020 3530.690 925.020 3530.700 ;
        RECT 1102.020 3530.690 1105.020 3530.700 ;
        RECT 1282.020 3530.690 1285.020 3530.700 ;
        RECT 1462.020 3530.690 1465.020 3530.700 ;
        RECT 1642.020 3530.690 1645.020 3530.700 ;
        RECT 1822.020 3530.690 1825.020 3530.700 ;
        RECT 2002.020 3530.690 2005.020 3530.700 ;
        RECT 2182.020 3530.690 2185.020 3530.700 ;
        RECT 2362.020 3530.690 2365.020 3530.700 ;
        RECT 2542.020 3530.690 2545.020 3530.700 ;
        RECT 2722.020 3530.690 2725.020 3530.700 ;
        RECT 2902.020 3530.690 2905.020 3530.700 ;
        RECT 2936.000 3530.690 2939.000 3530.700 ;
        RECT -9.980 3524.300 -6.980 3524.310 ;
        RECT 4.020 3524.300 7.020 3524.310 ;
        RECT 184.020 3524.300 187.020 3524.310 ;
        RECT 364.020 3524.300 367.020 3524.310 ;
        RECT 544.020 3524.300 547.020 3524.310 ;
        RECT 724.020 3524.300 727.020 3524.310 ;
        RECT 904.020 3524.300 907.020 3524.310 ;
        RECT 1084.020 3524.300 1087.020 3524.310 ;
        RECT 1264.020 3524.300 1267.020 3524.310 ;
        RECT 1444.020 3524.300 1447.020 3524.310 ;
        RECT 1624.020 3524.300 1627.020 3524.310 ;
        RECT 1804.020 3524.300 1807.020 3524.310 ;
        RECT 1984.020 3524.300 1987.020 3524.310 ;
        RECT 2164.020 3524.300 2167.020 3524.310 ;
        RECT 2344.020 3524.300 2347.020 3524.310 ;
        RECT 2524.020 3524.300 2527.020 3524.310 ;
        RECT 2704.020 3524.300 2707.020 3524.310 ;
        RECT 2884.020 3524.300 2887.020 3524.310 ;
        RECT 2926.600 3524.300 2929.600 3524.310 ;
        RECT -9.980 3521.300 2929.600 3524.300 ;
        RECT -9.980 3521.290 -6.980 3521.300 ;
        RECT 4.020 3521.290 7.020 3521.300 ;
        RECT 184.020 3521.290 187.020 3521.300 ;
        RECT 364.020 3521.290 367.020 3521.300 ;
        RECT 544.020 3521.290 547.020 3521.300 ;
        RECT 724.020 3521.290 727.020 3521.300 ;
        RECT 904.020 3521.290 907.020 3521.300 ;
        RECT 1084.020 3521.290 1087.020 3521.300 ;
        RECT 1264.020 3521.290 1267.020 3521.300 ;
        RECT 1444.020 3521.290 1447.020 3521.300 ;
        RECT 1624.020 3521.290 1627.020 3521.300 ;
        RECT 1804.020 3521.290 1807.020 3521.300 ;
        RECT 1984.020 3521.290 1987.020 3521.300 ;
        RECT 2164.020 3521.290 2167.020 3521.300 ;
        RECT 2344.020 3521.290 2347.020 3521.300 ;
        RECT 2524.020 3521.290 2527.020 3521.300 ;
        RECT 2704.020 3521.290 2707.020 3521.300 ;
        RECT 2884.020 3521.290 2887.020 3521.300 ;
        RECT 2926.600 3521.290 2929.600 3521.300 ;
        RECT -38.180 3486.380 -35.180 3486.390 ;
        RECT 58.020 3486.380 61.020 3486.390 ;
        RECT 238.020 3486.380 241.020 3486.390 ;
        RECT 418.020 3486.380 421.020 3486.390 ;
        RECT 598.020 3486.380 601.020 3486.390 ;
        RECT 778.020 3486.380 781.020 3486.390 ;
        RECT 958.020 3486.380 961.020 3486.390 ;
        RECT 1138.020 3486.380 1141.020 3486.390 ;
        RECT 1318.020 3486.380 1321.020 3486.390 ;
        RECT 1498.020 3486.380 1501.020 3486.390 ;
        RECT 1678.020 3486.380 1681.020 3486.390 ;
        RECT 1858.020 3486.380 1861.020 3486.390 ;
        RECT 2038.020 3486.380 2041.020 3486.390 ;
        RECT 2218.020 3486.380 2221.020 3486.390 ;
        RECT 2398.020 3486.380 2401.020 3486.390 ;
        RECT 2578.020 3486.380 2581.020 3486.390 ;
        RECT 2758.020 3486.380 2761.020 3486.390 ;
        RECT 2954.800 3486.380 2957.800 3486.390 ;
        RECT -42.880 3483.380 2962.500 3486.380 ;
        RECT -38.180 3483.370 -35.180 3483.380 ;
        RECT 58.020 3483.370 61.020 3483.380 ;
        RECT 238.020 3483.370 241.020 3483.380 ;
        RECT 418.020 3483.370 421.020 3483.380 ;
        RECT 598.020 3483.370 601.020 3483.380 ;
        RECT 778.020 3483.370 781.020 3483.380 ;
        RECT 958.020 3483.370 961.020 3483.380 ;
        RECT 1138.020 3483.370 1141.020 3483.380 ;
        RECT 1318.020 3483.370 1321.020 3483.380 ;
        RECT 1498.020 3483.370 1501.020 3483.380 ;
        RECT 1678.020 3483.370 1681.020 3483.380 ;
        RECT 1858.020 3483.370 1861.020 3483.380 ;
        RECT 2038.020 3483.370 2041.020 3483.380 ;
        RECT 2218.020 3483.370 2221.020 3483.380 ;
        RECT 2398.020 3483.370 2401.020 3483.380 ;
        RECT 2578.020 3483.370 2581.020 3483.380 ;
        RECT 2758.020 3483.370 2761.020 3483.380 ;
        RECT 2954.800 3483.370 2957.800 3483.380 ;
        RECT -28.780 3468.380 -25.780 3468.390 ;
        RECT 40.020 3468.380 43.020 3468.390 ;
        RECT 220.020 3468.380 223.020 3468.390 ;
        RECT 400.020 3468.380 403.020 3468.390 ;
        RECT 580.020 3468.380 583.020 3468.390 ;
        RECT 760.020 3468.380 763.020 3468.390 ;
        RECT 940.020 3468.380 943.020 3468.390 ;
        RECT 1120.020 3468.380 1123.020 3468.390 ;
        RECT 1300.020 3468.380 1303.020 3468.390 ;
        RECT 1480.020 3468.380 1483.020 3468.390 ;
        RECT 1660.020 3468.380 1663.020 3468.390 ;
        RECT 1840.020 3468.380 1843.020 3468.390 ;
        RECT 2020.020 3468.380 2023.020 3468.390 ;
        RECT 2200.020 3468.380 2203.020 3468.390 ;
        RECT 2380.020 3468.380 2383.020 3468.390 ;
        RECT 2560.020 3468.380 2563.020 3468.390 ;
        RECT 2740.020 3468.380 2743.020 3468.390 ;
        RECT 2945.400 3468.380 2948.400 3468.390 ;
        RECT -33.480 3465.380 2953.100 3468.380 ;
        RECT -28.780 3465.370 -25.780 3465.380 ;
        RECT 40.020 3465.370 43.020 3465.380 ;
        RECT 220.020 3465.370 223.020 3465.380 ;
        RECT 400.020 3465.370 403.020 3465.380 ;
        RECT 580.020 3465.370 583.020 3465.380 ;
        RECT 760.020 3465.370 763.020 3465.380 ;
        RECT 940.020 3465.370 943.020 3465.380 ;
        RECT 1120.020 3465.370 1123.020 3465.380 ;
        RECT 1300.020 3465.370 1303.020 3465.380 ;
        RECT 1480.020 3465.370 1483.020 3465.380 ;
        RECT 1660.020 3465.370 1663.020 3465.380 ;
        RECT 1840.020 3465.370 1843.020 3465.380 ;
        RECT 2020.020 3465.370 2023.020 3465.380 ;
        RECT 2200.020 3465.370 2203.020 3465.380 ;
        RECT 2380.020 3465.370 2383.020 3465.380 ;
        RECT 2560.020 3465.370 2563.020 3465.380 ;
        RECT 2740.020 3465.370 2743.020 3465.380 ;
        RECT 2945.400 3465.370 2948.400 3465.380 ;
        RECT -19.380 3450.380 -16.380 3450.390 ;
        RECT 22.020 3450.380 25.020 3450.390 ;
        RECT 202.020 3450.380 205.020 3450.390 ;
        RECT 382.020 3450.380 385.020 3450.390 ;
        RECT 562.020 3450.380 565.020 3450.390 ;
        RECT 742.020 3450.380 745.020 3450.390 ;
        RECT 922.020 3450.380 925.020 3450.390 ;
        RECT 1102.020 3450.380 1105.020 3450.390 ;
        RECT 1282.020 3450.380 1285.020 3450.390 ;
        RECT 1462.020 3450.380 1465.020 3450.390 ;
        RECT 1642.020 3450.380 1645.020 3450.390 ;
        RECT 1822.020 3450.380 1825.020 3450.390 ;
        RECT 2002.020 3450.380 2005.020 3450.390 ;
        RECT 2182.020 3450.380 2185.020 3450.390 ;
        RECT 2362.020 3450.380 2365.020 3450.390 ;
        RECT 2542.020 3450.380 2545.020 3450.390 ;
        RECT 2722.020 3450.380 2725.020 3450.390 ;
        RECT 2902.020 3450.380 2905.020 3450.390 ;
        RECT 2936.000 3450.380 2939.000 3450.390 ;
        RECT -24.080 3447.380 2943.700 3450.380 ;
        RECT -19.380 3447.370 -16.380 3447.380 ;
        RECT 22.020 3447.370 25.020 3447.380 ;
        RECT 202.020 3447.370 205.020 3447.380 ;
        RECT 382.020 3447.370 385.020 3447.380 ;
        RECT 562.020 3447.370 565.020 3447.380 ;
        RECT 742.020 3447.370 745.020 3447.380 ;
        RECT 922.020 3447.370 925.020 3447.380 ;
        RECT 1102.020 3447.370 1105.020 3447.380 ;
        RECT 1282.020 3447.370 1285.020 3447.380 ;
        RECT 1462.020 3447.370 1465.020 3447.380 ;
        RECT 1642.020 3447.370 1645.020 3447.380 ;
        RECT 1822.020 3447.370 1825.020 3447.380 ;
        RECT 2002.020 3447.370 2005.020 3447.380 ;
        RECT 2182.020 3447.370 2185.020 3447.380 ;
        RECT 2362.020 3447.370 2365.020 3447.380 ;
        RECT 2542.020 3447.370 2545.020 3447.380 ;
        RECT 2722.020 3447.370 2725.020 3447.380 ;
        RECT 2902.020 3447.370 2905.020 3447.380 ;
        RECT 2936.000 3447.370 2939.000 3447.380 ;
        RECT -9.980 3432.380 -6.980 3432.390 ;
        RECT 4.020 3432.380 7.020 3432.390 ;
        RECT 184.020 3432.380 187.020 3432.390 ;
        RECT 364.020 3432.380 367.020 3432.390 ;
        RECT 544.020 3432.380 547.020 3432.390 ;
        RECT 724.020 3432.380 727.020 3432.390 ;
        RECT 904.020 3432.380 907.020 3432.390 ;
        RECT 1084.020 3432.380 1087.020 3432.390 ;
        RECT 1264.020 3432.380 1267.020 3432.390 ;
        RECT 1444.020 3432.380 1447.020 3432.390 ;
        RECT 1624.020 3432.380 1627.020 3432.390 ;
        RECT 1804.020 3432.380 1807.020 3432.390 ;
        RECT 1984.020 3432.380 1987.020 3432.390 ;
        RECT 2164.020 3432.380 2167.020 3432.390 ;
        RECT 2344.020 3432.380 2347.020 3432.390 ;
        RECT 2524.020 3432.380 2527.020 3432.390 ;
        RECT 2704.020 3432.380 2707.020 3432.390 ;
        RECT 2884.020 3432.380 2887.020 3432.390 ;
        RECT 2926.600 3432.380 2929.600 3432.390 ;
        RECT -14.680 3429.380 2934.300 3432.380 ;
        RECT -9.980 3429.370 -6.980 3429.380 ;
        RECT 4.020 3429.370 7.020 3429.380 ;
        RECT 184.020 3429.370 187.020 3429.380 ;
        RECT 364.020 3429.370 367.020 3429.380 ;
        RECT 544.020 3429.370 547.020 3429.380 ;
        RECT 724.020 3429.370 727.020 3429.380 ;
        RECT 904.020 3429.370 907.020 3429.380 ;
        RECT 1084.020 3429.370 1087.020 3429.380 ;
        RECT 1264.020 3429.370 1267.020 3429.380 ;
        RECT 1444.020 3429.370 1447.020 3429.380 ;
        RECT 1624.020 3429.370 1627.020 3429.380 ;
        RECT 1804.020 3429.370 1807.020 3429.380 ;
        RECT 1984.020 3429.370 1987.020 3429.380 ;
        RECT 2164.020 3429.370 2167.020 3429.380 ;
        RECT 2344.020 3429.370 2347.020 3429.380 ;
        RECT 2524.020 3429.370 2527.020 3429.380 ;
        RECT 2704.020 3429.370 2707.020 3429.380 ;
        RECT 2884.020 3429.370 2887.020 3429.380 ;
        RECT 2926.600 3429.370 2929.600 3429.380 ;
        RECT -38.180 3306.380 -35.180 3306.390 ;
        RECT 58.020 3306.380 61.020 3306.390 ;
        RECT 238.020 3306.380 241.020 3306.390 ;
        RECT 418.020 3306.380 421.020 3306.390 ;
        RECT 598.020 3306.380 601.020 3306.390 ;
        RECT 778.020 3306.380 781.020 3306.390 ;
        RECT 958.020 3306.380 961.020 3306.390 ;
        RECT 1138.020 3306.380 1141.020 3306.390 ;
        RECT 1318.020 3306.380 1321.020 3306.390 ;
        RECT 1498.020 3306.380 1501.020 3306.390 ;
        RECT 1678.020 3306.380 1681.020 3306.390 ;
        RECT 1858.020 3306.380 1861.020 3306.390 ;
        RECT 2038.020 3306.380 2041.020 3306.390 ;
        RECT 2218.020 3306.380 2221.020 3306.390 ;
        RECT 2398.020 3306.380 2401.020 3306.390 ;
        RECT 2578.020 3306.380 2581.020 3306.390 ;
        RECT 2758.020 3306.380 2761.020 3306.390 ;
        RECT 2954.800 3306.380 2957.800 3306.390 ;
        RECT -42.880 3303.380 2962.500 3306.380 ;
        RECT -38.180 3303.370 -35.180 3303.380 ;
        RECT 58.020 3303.370 61.020 3303.380 ;
        RECT 238.020 3303.370 241.020 3303.380 ;
        RECT 418.020 3303.370 421.020 3303.380 ;
        RECT 598.020 3303.370 601.020 3303.380 ;
        RECT 778.020 3303.370 781.020 3303.380 ;
        RECT 958.020 3303.370 961.020 3303.380 ;
        RECT 1138.020 3303.370 1141.020 3303.380 ;
        RECT 1318.020 3303.370 1321.020 3303.380 ;
        RECT 1498.020 3303.370 1501.020 3303.380 ;
        RECT 1678.020 3303.370 1681.020 3303.380 ;
        RECT 1858.020 3303.370 1861.020 3303.380 ;
        RECT 2038.020 3303.370 2041.020 3303.380 ;
        RECT 2218.020 3303.370 2221.020 3303.380 ;
        RECT 2398.020 3303.370 2401.020 3303.380 ;
        RECT 2578.020 3303.370 2581.020 3303.380 ;
        RECT 2758.020 3303.370 2761.020 3303.380 ;
        RECT 2954.800 3303.370 2957.800 3303.380 ;
        RECT -28.780 3288.380 -25.780 3288.390 ;
        RECT 40.020 3288.380 43.020 3288.390 ;
        RECT 220.020 3288.380 223.020 3288.390 ;
        RECT 400.020 3288.380 403.020 3288.390 ;
        RECT 580.020 3288.380 583.020 3288.390 ;
        RECT 760.020 3288.380 763.020 3288.390 ;
        RECT 940.020 3288.380 943.020 3288.390 ;
        RECT 1120.020 3288.380 1123.020 3288.390 ;
        RECT 1300.020 3288.380 1303.020 3288.390 ;
        RECT 1480.020 3288.380 1483.020 3288.390 ;
        RECT 1660.020 3288.380 1663.020 3288.390 ;
        RECT 1840.020 3288.380 1843.020 3288.390 ;
        RECT 2020.020 3288.380 2023.020 3288.390 ;
        RECT 2200.020 3288.380 2203.020 3288.390 ;
        RECT 2380.020 3288.380 2383.020 3288.390 ;
        RECT 2560.020 3288.380 2563.020 3288.390 ;
        RECT 2740.020 3288.380 2743.020 3288.390 ;
        RECT 2945.400 3288.380 2948.400 3288.390 ;
        RECT -33.480 3285.380 2953.100 3288.380 ;
        RECT -28.780 3285.370 -25.780 3285.380 ;
        RECT 40.020 3285.370 43.020 3285.380 ;
        RECT 220.020 3285.370 223.020 3285.380 ;
        RECT 400.020 3285.370 403.020 3285.380 ;
        RECT 580.020 3285.370 583.020 3285.380 ;
        RECT 760.020 3285.370 763.020 3285.380 ;
        RECT 940.020 3285.370 943.020 3285.380 ;
        RECT 1120.020 3285.370 1123.020 3285.380 ;
        RECT 1300.020 3285.370 1303.020 3285.380 ;
        RECT 1480.020 3285.370 1483.020 3285.380 ;
        RECT 1660.020 3285.370 1663.020 3285.380 ;
        RECT 1840.020 3285.370 1843.020 3285.380 ;
        RECT 2020.020 3285.370 2023.020 3285.380 ;
        RECT 2200.020 3285.370 2203.020 3285.380 ;
        RECT 2380.020 3285.370 2383.020 3285.380 ;
        RECT 2560.020 3285.370 2563.020 3285.380 ;
        RECT 2740.020 3285.370 2743.020 3285.380 ;
        RECT 2945.400 3285.370 2948.400 3285.380 ;
        RECT -19.380 3270.380 -16.380 3270.390 ;
        RECT 22.020 3270.380 25.020 3270.390 ;
        RECT 202.020 3270.380 205.020 3270.390 ;
        RECT 382.020 3270.380 385.020 3270.390 ;
        RECT 562.020 3270.380 565.020 3270.390 ;
        RECT 742.020 3270.380 745.020 3270.390 ;
        RECT 922.020 3270.380 925.020 3270.390 ;
        RECT 1102.020 3270.380 1105.020 3270.390 ;
        RECT 1282.020 3270.380 1285.020 3270.390 ;
        RECT 1462.020 3270.380 1465.020 3270.390 ;
        RECT 1642.020 3270.380 1645.020 3270.390 ;
        RECT 1822.020 3270.380 1825.020 3270.390 ;
        RECT 2002.020 3270.380 2005.020 3270.390 ;
        RECT 2182.020 3270.380 2185.020 3270.390 ;
        RECT 2362.020 3270.380 2365.020 3270.390 ;
        RECT 2542.020 3270.380 2545.020 3270.390 ;
        RECT 2722.020 3270.380 2725.020 3270.390 ;
        RECT 2902.020 3270.380 2905.020 3270.390 ;
        RECT 2936.000 3270.380 2939.000 3270.390 ;
        RECT -24.080 3267.380 2943.700 3270.380 ;
        RECT -19.380 3267.370 -16.380 3267.380 ;
        RECT 22.020 3267.370 25.020 3267.380 ;
        RECT 202.020 3267.370 205.020 3267.380 ;
        RECT 382.020 3267.370 385.020 3267.380 ;
        RECT 562.020 3267.370 565.020 3267.380 ;
        RECT 742.020 3267.370 745.020 3267.380 ;
        RECT 922.020 3267.370 925.020 3267.380 ;
        RECT 1102.020 3267.370 1105.020 3267.380 ;
        RECT 1282.020 3267.370 1285.020 3267.380 ;
        RECT 1462.020 3267.370 1465.020 3267.380 ;
        RECT 1642.020 3267.370 1645.020 3267.380 ;
        RECT 1822.020 3267.370 1825.020 3267.380 ;
        RECT 2002.020 3267.370 2005.020 3267.380 ;
        RECT 2182.020 3267.370 2185.020 3267.380 ;
        RECT 2362.020 3267.370 2365.020 3267.380 ;
        RECT 2542.020 3267.370 2545.020 3267.380 ;
        RECT 2722.020 3267.370 2725.020 3267.380 ;
        RECT 2902.020 3267.370 2905.020 3267.380 ;
        RECT 2936.000 3267.370 2939.000 3267.380 ;
        RECT -9.980 3252.380 -6.980 3252.390 ;
        RECT 4.020 3252.380 7.020 3252.390 ;
        RECT 184.020 3252.380 187.020 3252.390 ;
        RECT 364.020 3252.380 367.020 3252.390 ;
        RECT 544.020 3252.380 547.020 3252.390 ;
        RECT 724.020 3252.380 727.020 3252.390 ;
        RECT 904.020 3252.380 907.020 3252.390 ;
        RECT 1084.020 3252.380 1087.020 3252.390 ;
        RECT 1264.020 3252.380 1267.020 3252.390 ;
        RECT 1444.020 3252.380 1447.020 3252.390 ;
        RECT 1624.020 3252.380 1627.020 3252.390 ;
        RECT 1804.020 3252.380 1807.020 3252.390 ;
        RECT 1984.020 3252.380 1987.020 3252.390 ;
        RECT 2164.020 3252.380 2167.020 3252.390 ;
        RECT 2344.020 3252.380 2347.020 3252.390 ;
        RECT 2524.020 3252.380 2527.020 3252.390 ;
        RECT 2704.020 3252.380 2707.020 3252.390 ;
        RECT 2884.020 3252.380 2887.020 3252.390 ;
        RECT 2926.600 3252.380 2929.600 3252.390 ;
        RECT -14.680 3249.380 2934.300 3252.380 ;
        RECT -9.980 3249.370 -6.980 3249.380 ;
        RECT 4.020 3249.370 7.020 3249.380 ;
        RECT 184.020 3249.370 187.020 3249.380 ;
        RECT 364.020 3249.370 367.020 3249.380 ;
        RECT 544.020 3249.370 547.020 3249.380 ;
        RECT 724.020 3249.370 727.020 3249.380 ;
        RECT 904.020 3249.370 907.020 3249.380 ;
        RECT 1084.020 3249.370 1087.020 3249.380 ;
        RECT 1264.020 3249.370 1267.020 3249.380 ;
        RECT 1444.020 3249.370 1447.020 3249.380 ;
        RECT 1624.020 3249.370 1627.020 3249.380 ;
        RECT 1804.020 3249.370 1807.020 3249.380 ;
        RECT 1984.020 3249.370 1987.020 3249.380 ;
        RECT 2164.020 3249.370 2167.020 3249.380 ;
        RECT 2344.020 3249.370 2347.020 3249.380 ;
        RECT 2524.020 3249.370 2527.020 3249.380 ;
        RECT 2704.020 3249.370 2707.020 3249.380 ;
        RECT 2884.020 3249.370 2887.020 3249.380 ;
        RECT 2926.600 3249.370 2929.600 3249.380 ;
        RECT -38.180 3126.380 -35.180 3126.390 ;
        RECT 58.020 3126.380 61.020 3126.390 ;
        RECT 238.020 3126.380 241.020 3126.390 ;
        RECT 418.020 3126.380 421.020 3126.390 ;
        RECT 598.020 3126.380 601.020 3126.390 ;
        RECT 778.020 3126.380 781.020 3126.390 ;
        RECT 958.020 3126.380 961.020 3126.390 ;
        RECT 1138.020 3126.380 1141.020 3126.390 ;
        RECT 1318.020 3126.380 1321.020 3126.390 ;
        RECT 1498.020 3126.380 1501.020 3126.390 ;
        RECT 1678.020 3126.380 1681.020 3126.390 ;
        RECT 1858.020 3126.380 1861.020 3126.390 ;
        RECT 2038.020 3126.380 2041.020 3126.390 ;
        RECT 2218.020 3126.380 2221.020 3126.390 ;
        RECT 2398.020 3126.380 2401.020 3126.390 ;
        RECT 2578.020 3126.380 2581.020 3126.390 ;
        RECT 2758.020 3126.380 2761.020 3126.390 ;
        RECT 2954.800 3126.380 2957.800 3126.390 ;
        RECT -42.880 3123.380 2962.500 3126.380 ;
        RECT -38.180 3123.370 -35.180 3123.380 ;
        RECT 58.020 3123.370 61.020 3123.380 ;
        RECT 238.020 3123.370 241.020 3123.380 ;
        RECT 418.020 3123.370 421.020 3123.380 ;
        RECT 598.020 3123.370 601.020 3123.380 ;
        RECT 778.020 3123.370 781.020 3123.380 ;
        RECT 958.020 3123.370 961.020 3123.380 ;
        RECT 1138.020 3123.370 1141.020 3123.380 ;
        RECT 1318.020 3123.370 1321.020 3123.380 ;
        RECT 1498.020 3123.370 1501.020 3123.380 ;
        RECT 1678.020 3123.370 1681.020 3123.380 ;
        RECT 1858.020 3123.370 1861.020 3123.380 ;
        RECT 2038.020 3123.370 2041.020 3123.380 ;
        RECT 2218.020 3123.370 2221.020 3123.380 ;
        RECT 2398.020 3123.370 2401.020 3123.380 ;
        RECT 2578.020 3123.370 2581.020 3123.380 ;
        RECT 2758.020 3123.370 2761.020 3123.380 ;
        RECT 2954.800 3123.370 2957.800 3123.380 ;
        RECT -28.780 3108.380 -25.780 3108.390 ;
        RECT 40.020 3108.380 43.020 3108.390 ;
        RECT 220.020 3108.380 223.020 3108.390 ;
        RECT 400.020 3108.380 403.020 3108.390 ;
        RECT 580.020 3108.380 583.020 3108.390 ;
        RECT 760.020 3108.380 763.020 3108.390 ;
        RECT 940.020 3108.380 943.020 3108.390 ;
        RECT 1120.020 3108.380 1123.020 3108.390 ;
        RECT 1300.020 3108.380 1303.020 3108.390 ;
        RECT 1480.020 3108.380 1483.020 3108.390 ;
        RECT 1660.020 3108.380 1663.020 3108.390 ;
        RECT 1840.020 3108.380 1843.020 3108.390 ;
        RECT 2020.020 3108.380 2023.020 3108.390 ;
        RECT 2200.020 3108.380 2203.020 3108.390 ;
        RECT 2380.020 3108.380 2383.020 3108.390 ;
        RECT 2560.020 3108.380 2563.020 3108.390 ;
        RECT 2740.020 3108.380 2743.020 3108.390 ;
        RECT 2945.400 3108.380 2948.400 3108.390 ;
        RECT -33.480 3105.380 2953.100 3108.380 ;
        RECT -28.780 3105.370 -25.780 3105.380 ;
        RECT 40.020 3105.370 43.020 3105.380 ;
        RECT 220.020 3105.370 223.020 3105.380 ;
        RECT 400.020 3105.370 403.020 3105.380 ;
        RECT 580.020 3105.370 583.020 3105.380 ;
        RECT 760.020 3105.370 763.020 3105.380 ;
        RECT 940.020 3105.370 943.020 3105.380 ;
        RECT 1120.020 3105.370 1123.020 3105.380 ;
        RECT 1300.020 3105.370 1303.020 3105.380 ;
        RECT 1480.020 3105.370 1483.020 3105.380 ;
        RECT 1660.020 3105.370 1663.020 3105.380 ;
        RECT 1840.020 3105.370 1843.020 3105.380 ;
        RECT 2020.020 3105.370 2023.020 3105.380 ;
        RECT 2200.020 3105.370 2203.020 3105.380 ;
        RECT 2380.020 3105.370 2383.020 3105.380 ;
        RECT 2560.020 3105.370 2563.020 3105.380 ;
        RECT 2740.020 3105.370 2743.020 3105.380 ;
        RECT 2945.400 3105.370 2948.400 3105.380 ;
        RECT -19.380 3090.380 -16.380 3090.390 ;
        RECT 22.020 3090.380 25.020 3090.390 ;
        RECT 202.020 3090.380 205.020 3090.390 ;
        RECT 382.020 3090.380 385.020 3090.390 ;
        RECT 562.020 3090.380 565.020 3090.390 ;
        RECT 742.020 3090.380 745.020 3090.390 ;
        RECT 922.020 3090.380 925.020 3090.390 ;
        RECT 1102.020 3090.380 1105.020 3090.390 ;
        RECT 1282.020 3090.380 1285.020 3090.390 ;
        RECT 1462.020 3090.380 1465.020 3090.390 ;
        RECT 1642.020 3090.380 1645.020 3090.390 ;
        RECT 1822.020 3090.380 1825.020 3090.390 ;
        RECT 2002.020 3090.380 2005.020 3090.390 ;
        RECT 2182.020 3090.380 2185.020 3090.390 ;
        RECT 2362.020 3090.380 2365.020 3090.390 ;
        RECT 2542.020 3090.380 2545.020 3090.390 ;
        RECT 2722.020 3090.380 2725.020 3090.390 ;
        RECT 2902.020 3090.380 2905.020 3090.390 ;
        RECT 2936.000 3090.380 2939.000 3090.390 ;
        RECT -24.080 3087.380 2943.700 3090.380 ;
        RECT -19.380 3087.370 -16.380 3087.380 ;
        RECT 22.020 3087.370 25.020 3087.380 ;
        RECT 202.020 3087.370 205.020 3087.380 ;
        RECT 382.020 3087.370 385.020 3087.380 ;
        RECT 562.020 3087.370 565.020 3087.380 ;
        RECT 742.020 3087.370 745.020 3087.380 ;
        RECT 922.020 3087.370 925.020 3087.380 ;
        RECT 1102.020 3087.370 1105.020 3087.380 ;
        RECT 1282.020 3087.370 1285.020 3087.380 ;
        RECT 1462.020 3087.370 1465.020 3087.380 ;
        RECT 1642.020 3087.370 1645.020 3087.380 ;
        RECT 1822.020 3087.370 1825.020 3087.380 ;
        RECT 2002.020 3087.370 2005.020 3087.380 ;
        RECT 2182.020 3087.370 2185.020 3087.380 ;
        RECT 2362.020 3087.370 2365.020 3087.380 ;
        RECT 2542.020 3087.370 2545.020 3087.380 ;
        RECT 2722.020 3087.370 2725.020 3087.380 ;
        RECT 2902.020 3087.370 2905.020 3087.380 ;
        RECT 2936.000 3087.370 2939.000 3087.380 ;
        RECT -9.980 3072.380 -6.980 3072.390 ;
        RECT 4.020 3072.380 7.020 3072.390 ;
        RECT 184.020 3072.380 187.020 3072.390 ;
        RECT 364.020 3072.380 367.020 3072.390 ;
        RECT 544.020 3072.380 547.020 3072.390 ;
        RECT 724.020 3072.380 727.020 3072.390 ;
        RECT 904.020 3072.380 907.020 3072.390 ;
        RECT 1084.020 3072.380 1087.020 3072.390 ;
        RECT 1264.020 3072.380 1267.020 3072.390 ;
        RECT 1444.020 3072.380 1447.020 3072.390 ;
        RECT 1624.020 3072.380 1627.020 3072.390 ;
        RECT 1804.020 3072.380 1807.020 3072.390 ;
        RECT 1984.020 3072.380 1987.020 3072.390 ;
        RECT 2164.020 3072.380 2167.020 3072.390 ;
        RECT 2344.020 3072.380 2347.020 3072.390 ;
        RECT 2524.020 3072.380 2527.020 3072.390 ;
        RECT 2704.020 3072.380 2707.020 3072.390 ;
        RECT 2884.020 3072.380 2887.020 3072.390 ;
        RECT 2926.600 3072.380 2929.600 3072.390 ;
        RECT -14.680 3069.380 2934.300 3072.380 ;
        RECT -9.980 3069.370 -6.980 3069.380 ;
        RECT 4.020 3069.370 7.020 3069.380 ;
        RECT 184.020 3069.370 187.020 3069.380 ;
        RECT 364.020 3069.370 367.020 3069.380 ;
        RECT 544.020 3069.370 547.020 3069.380 ;
        RECT 724.020 3069.370 727.020 3069.380 ;
        RECT 904.020 3069.370 907.020 3069.380 ;
        RECT 1084.020 3069.370 1087.020 3069.380 ;
        RECT 1264.020 3069.370 1267.020 3069.380 ;
        RECT 1444.020 3069.370 1447.020 3069.380 ;
        RECT 1624.020 3069.370 1627.020 3069.380 ;
        RECT 1804.020 3069.370 1807.020 3069.380 ;
        RECT 1984.020 3069.370 1987.020 3069.380 ;
        RECT 2164.020 3069.370 2167.020 3069.380 ;
        RECT 2344.020 3069.370 2347.020 3069.380 ;
        RECT 2524.020 3069.370 2527.020 3069.380 ;
        RECT 2704.020 3069.370 2707.020 3069.380 ;
        RECT 2884.020 3069.370 2887.020 3069.380 ;
        RECT 2926.600 3069.370 2929.600 3069.380 ;
        RECT -38.180 2946.380 -35.180 2946.390 ;
        RECT 58.020 2946.380 61.020 2946.390 ;
        RECT 238.020 2946.380 241.020 2946.390 ;
        RECT 418.020 2946.380 421.020 2946.390 ;
        RECT 598.020 2946.380 601.020 2946.390 ;
        RECT 778.020 2946.380 781.020 2946.390 ;
        RECT 958.020 2946.380 961.020 2946.390 ;
        RECT 1138.020 2946.380 1141.020 2946.390 ;
        RECT 1318.020 2946.380 1321.020 2946.390 ;
        RECT 1498.020 2946.380 1501.020 2946.390 ;
        RECT 1678.020 2946.380 1681.020 2946.390 ;
        RECT 1858.020 2946.380 1861.020 2946.390 ;
        RECT 2038.020 2946.380 2041.020 2946.390 ;
        RECT 2218.020 2946.380 2221.020 2946.390 ;
        RECT 2398.020 2946.380 2401.020 2946.390 ;
        RECT 2578.020 2946.380 2581.020 2946.390 ;
        RECT 2758.020 2946.380 2761.020 2946.390 ;
        RECT 2954.800 2946.380 2957.800 2946.390 ;
        RECT -42.880 2943.380 2962.500 2946.380 ;
        RECT -38.180 2943.370 -35.180 2943.380 ;
        RECT 58.020 2943.370 61.020 2943.380 ;
        RECT 238.020 2943.370 241.020 2943.380 ;
        RECT 418.020 2943.370 421.020 2943.380 ;
        RECT 598.020 2943.370 601.020 2943.380 ;
        RECT 778.020 2943.370 781.020 2943.380 ;
        RECT 958.020 2943.370 961.020 2943.380 ;
        RECT 1138.020 2943.370 1141.020 2943.380 ;
        RECT 1318.020 2943.370 1321.020 2943.380 ;
        RECT 1498.020 2943.370 1501.020 2943.380 ;
        RECT 1678.020 2943.370 1681.020 2943.380 ;
        RECT 1858.020 2943.370 1861.020 2943.380 ;
        RECT 2038.020 2943.370 2041.020 2943.380 ;
        RECT 2218.020 2943.370 2221.020 2943.380 ;
        RECT 2398.020 2943.370 2401.020 2943.380 ;
        RECT 2578.020 2943.370 2581.020 2943.380 ;
        RECT 2758.020 2943.370 2761.020 2943.380 ;
        RECT 2954.800 2943.370 2957.800 2943.380 ;
        RECT -28.780 2928.380 -25.780 2928.390 ;
        RECT 40.020 2928.380 43.020 2928.390 ;
        RECT 220.020 2928.380 223.020 2928.390 ;
        RECT 400.020 2928.380 403.020 2928.390 ;
        RECT 580.020 2928.380 583.020 2928.390 ;
        RECT 760.020 2928.380 763.020 2928.390 ;
        RECT 940.020 2928.380 943.020 2928.390 ;
        RECT 1120.020 2928.380 1123.020 2928.390 ;
        RECT 1300.020 2928.380 1303.020 2928.390 ;
        RECT 1480.020 2928.380 1483.020 2928.390 ;
        RECT 1660.020 2928.380 1663.020 2928.390 ;
        RECT 1840.020 2928.380 1843.020 2928.390 ;
        RECT 2020.020 2928.380 2023.020 2928.390 ;
        RECT 2200.020 2928.380 2203.020 2928.390 ;
        RECT 2380.020 2928.380 2383.020 2928.390 ;
        RECT 2560.020 2928.380 2563.020 2928.390 ;
        RECT 2740.020 2928.380 2743.020 2928.390 ;
        RECT 2945.400 2928.380 2948.400 2928.390 ;
        RECT -33.480 2925.380 2953.100 2928.380 ;
        RECT -28.780 2925.370 -25.780 2925.380 ;
        RECT 40.020 2925.370 43.020 2925.380 ;
        RECT 220.020 2925.370 223.020 2925.380 ;
        RECT 400.020 2925.370 403.020 2925.380 ;
        RECT 580.020 2925.370 583.020 2925.380 ;
        RECT 760.020 2925.370 763.020 2925.380 ;
        RECT 940.020 2925.370 943.020 2925.380 ;
        RECT 1120.020 2925.370 1123.020 2925.380 ;
        RECT 1300.020 2925.370 1303.020 2925.380 ;
        RECT 1480.020 2925.370 1483.020 2925.380 ;
        RECT 1660.020 2925.370 1663.020 2925.380 ;
        RECT 1840.020 2925.370 1843.020 2925.380 ;
        RECT 2020.020 2925.370 2023.020 2925.380 ;
        RECT 2200.020 2925.370 2203.020 2925.380 ;
        RECT 2380.020 2925.370 2383.020 2925.380 ;
        RECT 2560.020 2925.370 2563.020 2925.380 ;
        RECT 2740.020 2925.370 2743.020 2925.380 ;
        RECT 2945.400 2925.370 2948.400 2925.380 ;
        RECT -19.380 2910.380 -16.380 2910.390 ;
        RECT 22.020 2910.380 25.020 2910.390 ;
        RECT 202.020 2910.380 205.020 2910.390 ;
        RECT 382.020 2910.380 385.020 2910.390 ;
        RECT 562.020 2910.380 565.020 2910.390 ;
        RECT 742.020 2910.380 745.020 2910.390 ;
        RECT 922.020 2910.380 925.020 2910.390 ;
        RECT 1102.020 2910.380 1105.020 2910.390 ;
        RECT 1282.020 2910.380 1285.020 2910.390 ;
        RECT 1462.020 2910.380 1465.020 2910.390 ;
        RECT 1642.020 2910.380 1645.020 2910.390 ;
        RECT 1822.020 2910.380 1825.020 2910.390 ;
        RECT 2002.020 2910.380 2005.020 2910.390 ;
        RECT 2182.020 2910.380 2185.020 2910.390 ;
        RECT 2362.020 2910.380 2365.020 2910.390 ;
        RECT 2542.020 2910.380 2545.020 2910.390 ;
        RECT 2722.020 2910.380 2725.020 2910.390 ;
        RECT 2902.020 2910.380 2905.020 2910.390 ;
        RECT 2936.000 2910.380 2939.000 2910.390 ;
        RECT -24.080 2907.380 2943.700 2910.380 ;
        RECT -19.380 2907.370 -16.380 2907.380 ;
        RECT 22.020 2907.370 25.020 2907.380 ;
        RECT 202.020 2907.370 205.020 2907.380 ;
        RECT 382.020 2907.370 385.020 2907.380 ;
        RECT 562.020 2907.370 565.020 2907.380 ;
        RECT 742.020 2907.370 745.020 2907.380 ;
        RECT 922.020 2907.370 925.020 2907.380 ;
        RECT 1102.020 2907.370 1105.020 2907.380 ;
        RECT 1282.020 2907.370 1285.020 2907.380 ;
        RECT 1462.020 2907.370 1465.020 2907.380 ;
        RECT 1642.020 2907.370 1645.020 2907.380 ;
        RECT 1822.020 2907.370 1825.020 2907.380 ;
        RECT 2002.020 2907.370 2005.020 2907.380 ;
        RECT 2182.020 2907.370 2185.020 2907.380 ;
        RECT 2362.020 2907.370 2365.020 2907.380 ;
        RECT 2542.020 2907.370 2545.020 2907.380 ;
        RECT 2722.020 2907.370 2725.020 2907.380 ;
        RECT 2902.020 2907.370 2905.020 2907.380 ;
        RECT 2936.000 2907.370 2939.000 2907.380 ;
        RECT -9.980 2892.380 -6.980 2892.390 ;
        RECT 4.020 2892.380 7.020 2892.390 ;
        RECT 184.020 2892.380 187.020 2892.390 ;
        RECT 364.020 2892.380 367.020 2892.390 ;
        RECT 544.020 2892.380 547.020 2892.390 ;
        RECT 724.020 2892.380 727.020 2892.390 ;
        RECT 904.020 2892.380 907.020 2892.390 ;
        RECT 1084.020 2892.380 1087.020 2892.390 ;
        RECT 1264.020 2892.380 1267.020 2892.390 ;
        RECT 1444.020 2892.380 1447.020 2892.390 ;
        RECT 1624.020 2892.380 1627.020 2892.390 ;
        RECT 1804.020 2892.380 1807.020 2892.390 ;
        RECT 1984.020 2892.380 1987.020 2892.390 ;
        RECT 2164.020 2892.380 2167.020 2892.390 ;
        RECT 2344.020 2892.380 2347.020 2892.390 ;
        RECT 2524.020 2892.380 2527.020 2892.390 ;
        RECT 2704.020 2892.380 2707.020 2892.390 ;
        RECT 2884.020 2892.380 2887.020 2892.390 ;
        RECT 2926.600 2892.380 2929.600 2892.390 ;
        RECT -14.680 2889.380 2934.300 2892.380 ;
        RECT -9.980 2889.370 -6.980 2889.380 ;
        RECT 4.020 2889.370 7.020 2889.380 ;
        RECT 184.020 2889.370 187.020 2889.380 ;
        RECT 364.020 2889.370 367.020 2889.380 ;
        RECT 544.020 2889.370 547.020 2889.380 ;
        RECT 724.020 2889.370 727.020 2889.380 ;
        RECT 904.020 2889.370 907.020 2889.380 ;
        RECT 1084.020 2889.370 1087.020 2889.380 ;
        RECT 1264.020 2889.370 1267.020 2889.380 ;
        RECT 1444.020 2889.370 1447.020 2889.380 ;
        RECT 1624.020 2889.370 1627.020 2889.380 ;
        RECT 1804.020 2889.370 1807.020 2889.380 ;
        RECT 1984.020 2889.370 1987.020 2889.380 ;
        RECT 2164.020 2889.370 2167.020 2889.380 ;
        RECT 2344.020 2889.370 2347.020 2889.380 ;
        RECT 2524.020 2889.370 2527.020 2889.380 ;
        RECT 2704.020 2889.370 2707.020 2889.380 ;
        RECT 2884.020 2889.370 2887.020 2889.380 ;
        RECT 2926.600 2889.370 2929.600 2889.380 ;
        RECT -38.180 2766.380 -35.180 2766.390 ;
        RECT 58.020 2766.380 61.020 2766.390 ;
        RECT 238.020 2766.380 241.020 2766.390 ;
        RECT 778.020 2766.380 781.020 2766.390 ;
        RECT 1498.020 2766.380 1501.020 2766.390 ;
        RECT 2038.020 2766.380 2041.020 2766.390 ;
        RECT 2758.020 2766.380 2761.020 2766.390 ;
        RECT 2954.800 2766.380 2957.800 2766.390 ;
        RECT -42.880 2763.380 2962.500 2766.380 ;
        RECT -38.180 2763.370 -35.180 2763.380 ;
        RECT 58.020 2763.370 61.020 2763.380 ;
        RECT 238.020 2763.370 241.020 2763.380 ;
        RECT 778.020 2763.370 781.020 2763.380 ;
        RECT 1498.020 2763.370 1501.020 2763.380 ;
        RECT 2038.020 2763.370 2041.020 2763.380 ;
        RECT 2758.020 2763.370 2761.020 2763.380 ;
        RECT 2954.800 2763.370 2957.800 2763.380 ;
        RECT -28.780 2748.380 -25.780 2748.390 ;
        RECT 40.020 2748.380 43.020 2748.390 ;
        RECT 220.020 2748.380 223.020 2748.390 ;
        RECT 760.020 2748.380 763.020 2748.390 ;
        RECT 1480.020 2748.380 1483.020 2748.390 ;
        RECT 2020.020 2748.380 2023.020 2748.390 ;
        RECT 2740.020 2748.380 2743.020 2748.390 ;
        RECT 2945.400 2748.380 2948.400 2748.390 ;
        RECT -33.480 2745.380 2953.100 2748.380 ;
        RECT -28.780 2745.370 -25.780 2745.380 ;
        RECT 40.020 2745.370 43.020 2745.380 ;
        RECT 220.020 2745.370 223.020 2745.380 ;
        RECT 760.020 2745.370 763.020 2745.380 ;
        RECT 1480.020 2745.370 1483.020 2745.380 ;
        RECT 2020.020 2745.370 2023.020 2745.380 ;
        RECT 2740.020 2745.370 2743.020 2745.380 ;
        RECT 2945.400 2745.370 2948.400 2745.380 ;
        RECT -19.380 2730.380 -16.380 2730.390 ;
        RECT 22.020 2730.380 25.020 2730.390 ;
        RECT 202.020 2730.380 205.020 2730.390 ;
        RECT 682.470 2730.380 684.070 2730.390 ;
        RECT 742.020 2730.380 745.020 2730.390 ;
        RECT 922.020 2730.380 925.020 2730.390 ;
        RECT 1332.470 2730.380 1334.070 2730.390 ;
        RECT 1462.020 2730.380 1465.020 2730.390 ;
        RECT 1932.470 2730.380 1934.070 2730.390 ;
        RECT 2002.020 2730.380 2005.020 2730.390 ;
        RECT 2582.470 2730.380 2584.070 2730.390 ;
        RECT 2722.020 2730.380 2725.020 2730.390 ;
        RECT 2902.020 2730.380 2905.020 2730.390 ;
        RECT 2936.000 2730.380 2939.000 2730.390 ;
        RECT -24.080 2727.380 2943.700 2730.380 ;
        RECT -19.380 2727.370 -16.380 2727.380 ;
        RECT 22.020 2727.370 25.020 2727.380 ;
        RECT 202.020 2727.370 205.020 2727.380 ;
        RECT 682.470 2727.370 684.070 2727.380 ;
        RECT 742.020 2727.370 745.020 2727.380 ;
        RECT 922.020 2727.370 925.020 2727.380 ;
        RECT 1332.470 2727.370 1334.070 2727.380 ;
        RECT 1462.020 2727.370 1465.020 2727.380 ;
        RECT 1932.470 2727.370 1934.070 2727.380 ;
        RECT 2002.020 2727.370 2005.020 2727.380 ;
        RECT 2582.470 2727.370 2584.070 2727.380 ;
        RECT 2722.020 2727.370 2725.020 2727.380 ;
        RECT 2902.020 2727.370 2905.020 2727.380 ;
        RECT 2936.000 2727.370 2939.000 2727.380 ;
        RECT -9.980 2712.380 -6.980 2712.390 ;
        RECT 4.020 2712.380 7.020 2712.390 ;
        RECT 184.020 2712.380 187.020 2712.390 ;
        RECT 682.470 2712.380 684.070 2712.390 ;
        RECT 724.020 2712.380 727.020 2712.390 ;
        RECT 904.020 2712.380 907.020 2712.390 ;
        RECT 1332.470 2712.380 1334.070 2712.390 ;
        RECT 1444.020 2712.380 1447.020 2712.390 ;
        RECT 1932.470 2712.380 1934.070 2712.390 ;
        RECT 1984.020 2712.380 1987.020 2712.390 ;
        RECT 2164.020 2712.380 2167.020 2712.390 ;
        RECT 2582.470 2712.380 2584.070 2712.390 ;
        RECT 2704.020 2712.380 2707.020 2712.390 ;
        RECT 2884.020 2712.380 2887.020 2712.390 ;
        RECT 2926.600 2712.380 2929.600 2712.390 ;
        RECT -14.680 2709.380 2934.300 2712.380 ;
        RECT -9.980 2709.370 -6.980 2709.380 ;
        RECT 4.020 2709.370 7.020 2709.380 ;
        RECT 184.020 2709.370 187.020 2709.380 ;
        RECT 682.470 2709.370 684.070 2709.380 ;
        RECT 724.020 2709.370 727.020 2709.380 ;
        RECT 904.020 2709.370 907.020 2709.380 ;
        RECT 1332.470 2709.370 1334.070 2709.380 ;
        RECT 1444.020 2709.370 1447.020 2709.380 ;
        RECT 1932.470 2709.370 1934.070 2709.380 ;
        RECT 1984.020 2709.370 1987.020 2709.380 ;
        RECT 2164.020 2709.370 2167.020 2709.380 ;
        RECT 2582.470 2709.370 2584.070 2709.380 ;
        RECT 2704.020 2709.370 2707.020 2709.380 ;
        RECT 2884.020 2709.370 2887.020 2709.380 ;
        RECT 2926.600 2709.370 2929.600 2709.380 ;
        RECT -38.180 2586.380 -35.180 2586.390 ;
        RECT 58.020 2586.380 61.020 2586.390 ;
        RECT 238.020 2586.380 241.020 2586.390 ;
        RECT 682.470 2586.380 684.070 2586.390 ;
        RECT 778.020 2586.380 781.020 2586.390 ;
        RECT 1332.470 2586.380 1334.070 2586.390 ;
        RECT 1498.020 2586.380 1501.020 2586.390 ;
        RECT 1932.470 2586.380 1934.070 2586.390 ;
        RECT 2038.020 2586.380 2041.020 2586.390 ;
        RECT 2582.470 2586.380 2584.070 2586.390 ;
        RECT 2758.020 2586.380 2761.020 2586.390 ;
        RECT 2954.800 2586.380 2957.800 2586.390 ;
        RECT -42.880 2583.380 2962.500 2586.380 ;
        RECT -38.180 2583.370 -35.180 2583.380 ;
        RECT 58.020 2583.370 61.020 2583.380 ;
        RECT 238.020 2583.370 241.020 2583.380 ;
        RECT 682.470 2583.370 684.070 2583.380 ;
        RECT 778.020 2583.370 781.020 2583.380 ;
        RECT 1332.470 2583.370 1334.070 2583.380 ;
        RECT 1498.020 2583.370 1501.020 2583.380 ;
        RECT 1932.470 2583.370 1934.070 2583.380 ;
        RECT 2038.020 2583.370 2041.020 2583.380 ;
        RECT 2582.470 2583.370 2584.070 2583.380 ;
        RECT 2758.020 2583.370 2761.020 2583.380 ;
        RECT 2954.800 2583.370 2957.800 2583.380 ;
        RECT -28.780 2568.380 -25.780 2568.390 ;
        RECT 40.020 2568.380 43.020 2568.390 ;
        RECT 220.020 2568.380 223.020 2568.390 ;
        RECT 682.470 2568.380 684.070 2568.390 ;
        RECT 760.020 2568.380 763.020 2568.390 ;
        RECT 1332.470 2568.380 1334.070 2568.390 ;
        RECT 1480.020 2568.380 1483.020 2568.390 ;
        RECT 1932.470 2568.380 1934.070 2568.390 ;
        RECT 2020.020 2568.380 2023.020 2568.390 ;
        RECT 2582.470 2568.380 2584.070 2568.390 ;
        RECT 2740.020 2568.380 2743.020 2568.390 ;
        RECT 2945.400 2568.380 2948.400 2568.390 ;
        RECT -33.480 2565.380 2953.100 2568.380 ;
        RECT -28.780 2565.370 -25.780 2565.380 ;
        RECT 40.020 2565.370 43.020 2565.380 ;
        RECT 220.020 2565.370 223.020 2565.380 ;
        RECT 682.470 2565.370 684.070 2565.380 ;
        RECT 760.020 2565.370 763.020 2565.380 ;
        RECT 1332.470 2565.370 1334.070 2565.380 ;
        RECT 1480.020 2565.370 1483.020 2565.380 ;
        RECT 1932.470 2565.370 1934.070 2565.380 ;
        RECT 2020.020 2565.370 2023.020 2565.380 ;
        RECT 2582.470 2565.370 2584.070 2565.380 ;
        RECT 2740.020 2565.370 2743.020 2565.380 ;
        RECT 2945.400 2565.370 2948.400 2565.380 ;
        RECT -19.380 2550.380 -16.380 2550.390 ;
        RECT 22.020 2550.380 25.020 2550.390 ;
        RECT 202.020 2550.380 205.020 2550.390 ;
        RECT 682.470 2550.380 684.070 2550.390 ;
        RECT 742.020 2550.380 745.020 2550.390 ;
        RECT 922.020 2550.380 925.020 2550.390 ;
        RECT 1332.470 2550.380 1334.070 2550.390 ;
        RECT 1462.020 2550.380 1465.020 2550.390 ;
        RECT 1932.470 2550.380 1934.070 2550.390 ;
        RECT 2002.020 2550.380 2005.020 2550.390 ;
        RECT 2582.470 2550.380 2584.070 2550.390 ;
        RECT 2722.020 2550.380 2725.020 2550.390 ;
        RECT 2902.020 2550.380 2905.020 2550.390 ;
        RECT 2936.000 2550.380 2939.000 2550.390 ;
        RECT -24.080 2547.380 2943.700 2550.380 ;
        RECT -19.380 2547.370 -16.380 2547.380 ;
        RECT 22.020 2547.370 25.020 2547.380 ;
        RECT 202.020 2547.370 205.020 2547.380 ;
        RECT 682.470 2547.370 684.070 2547.380 ;
        RECT 742.020 2547.370 745.020 2547.380 ;
        RECT 922.020 2547.370 925.020 2547.380 ;
        RECT 1332.470 2547.370 1334.070 2547.380 ;
        RECT 1462.020 2547.370 1465.020 2547.380 ;
        RECT 1932.470 2547.370 1934.070 2547.380 ;
        RECT 2002.020 2547.370 2005.020 2547.380 ;
        RECT 2582.470 2547.370 2584.070 2547.380 ;
        RECT 2722.020 2547.370 2725.020 2547.380 ;
        RECT 2902.020 2547.370 2905.020 2547.380 ;
        RECT 2936.000 2547.370 2939.000 2547.380 ;
        RECT -9.980 2532.380 -6.980 2532.390 ;
        RECT 4.020 2532.380 7.020 2532.390 ;
        RECT 184.020 2532.380 187.020 2532.390 ;
        RECT 682.470 2532.380 684.070 2532.390 ;
        RECT 724.020 2532.380 727.020 2532.390 ;
        RECT 904.020 2532.380 907.020 2532.390 ;
        RECT 1332.470 2532.380 1334.070 2532.390 ;
        RECT 1444.020 2532.380 1447.020 2532.390 ;
        RECT 1932.470 2532.380 1934.070 2532.390 ;
        RECT 1984.020 2532.380 1987.020 2532.390 ;
        RECT 2164.020 2532.380 2167.020 2532.390 ;
        RECT 2582.470 2532.380 2584.070 2532.390 ;
        RECT 2704.020 2532.380 2707.020 2532.390 ;
        RECT 2884.020 2532.380 2887.020 2532.390 ;
        RECT 2926.600 2532.380 2929.600 2532.390 ;
        RECT -14.680 2529.380 2934.300 2532.380 ;
        RECT -9.980 2529.370 -6.980 2529.380 ;
        RECT 4.020 2529.370 7.020 2529.380 ;
        RECT 184.020 2529.370 187.020 2529.380 ;
        RECT 682.470 2529.370 684.070 2529.380 ;
        RECT 724.020 2529.370 727.020 2529.380 ;
        RECT 904.020 2529.370 907.020 2529.380 ;
        RECT 1332.470 2529.370 1334.070 2529.380 ;
        RECT 1444.020 2529.370 1447.020 2529.380 ;
        RECT 1932.470 2529.370 1934.070 2529.380 ;
        RECT 1984.020 2529.370 1987.020 2529.380 ;
        RECT 2164.020 2529.370 2167.020 2529.380 ;
        RECT 2582.470 2529.370 2584.070 2529.380 ;
        RECT 2704.020 2529.370 2707.020 2529.380 ;
        RECT 2884.020 2529.370 2887.020 2529.380 ;
        RECT 2926.600 2529.370 2929.600 2529.380 ;
        RECT -38.180 2406.380 -35.180 2406.390 ;
        RECT 58.020 2406.380 61.020 2406.390 ;
        RECT 238.020 2406.380 241.020 2406.390 ;
        RECT 682.470 2406.380 684.070 2406.390 ;
        RECT 778.020 2406.380 781.020 2406.390 ;
        RECT 1332.470 2406.380 1334.070 2406.390 ;
        RECT 1498.020 2406.380 1501.020 2406.390 ;
        RECT 1932.470 2406.380 1934.070 2406.390 ;
        RECT 2038.020 2406.380 2041.020 2406.390 ;
        RECT 2582.470 2406.380 2584.070 2406.390 ;
        RECT 2758.020 2406.380 2761.020 2406.390 ;
        RECT 2954.800 2406.380 2957.800 2406.390 ;
        RECT -42.880 2403.380 2962.500 2406.380 ;
        RECT -38.180 2403.370 -35.180 2403.380 ;
        RECT 58.020 2403.370 61.020 2403.380 ;
        RECT 238.020 2403.370 241.020 2403.380 ;
        RECT 682.470 2403.370 684.070 2403.380 ;
        RECT 778.020 2403.370 781.020 2403.380 ;
        RECT 1332.470 2403.370 1334.070 2403.380 ;
        RECT 1498.020 2403.370 1501.020 2403.380 ;
        RECT 1932.470 2403.370 1934.070 2403.380 ;
        RECT 2038.020 2403.370 2041.020 2403.380 ;
        RECT 2582.470 2403.370 2584.070 2403.380 ;
        RECT 2758.020 2403.370 2761.020 2403.380 ;
        RECT 2954.800 2403.370 2957.800 2403.380 ;
        RECT -28.780 2388.380 -25.780 2388.390 ;
        RECT 40.020 2388.380 43.020 2388.390 ;
        RECT 220.020 2388.380 223.020 2388.390 ;
        RECT 682.470 2388.380 684.070 2388.390 ;
        RECT 760.020 2388.380 763.020 2388.390 ;
        RECT 1332.470 2388.380 1334.070 2388.390 ;
        RECT 1480.020 2388.380 1483.020 2388.390 ;
        RECT 1932.470 2388.380 1934.070 2388.390 ;
        RECT 2020.020 2388.380 2023.020 2388.390 ;
        RECT 2582.470 2388.380 2584.070 2388.390 ;
        RECT 2740.020 2388.380 2743.020 2388.390 ;
        RECT 2945.400 2388.380 2948.400 2388.390 ;
        RECT -33.480 2385.380 2953.100 2388.380 ;
        RECT -28.780 2385.370 -25.780 2385.380 ;
        RECT 40.020 2385.370 43.020 2385.380 ;
        RECT 220.020 2385.370 223.020 2385.380 ;
        RECT 682.470 2385.370 684.070 2385.380 ;
        RECT 760.020 2385.370 763.020 2385.380 ;
        RECT 1332.470 2385.370 1334.070 2385.380 ;
        RECT 1480.020 2385.370 1483.020 2385.380 ;
        RECT 1932.470 2385.370 1934.070 2385.380 ;
        RECT 2020.020 2385.370 2023.020 2385.380 ;
        RECT 2582.470 2385.370 2584.070 2385.380 ;
        RECT 2740.020 2385.370 2743.020 2385.380 ;
        RECT 2945.400 2385.370 2948.400 2385.380 ;
        RECT -19.380 2370.380 -16.380 2370.390 ;
        RECT 22.020 2370.380 25.020 2370.390 ;
        RECT 202.020 2370.380 205.020 2370.390 ;
        RECT 682.470 2370.380 684.070 2370.390 ;
        RECT 742.020 2370.380 745.020 2370.390 ;
        RECT 922.020 2370.380 925.020 2370.390 ;
        RECT 1332.470 2370.380 1334.070 2370.390 ;
        RECT 1462.020 2370.380 1465.020 2370.390 ;
        RECT 1932.470 2370.380 1934.070 2370.390 ;
        RECT 2002.020 2370.380 2005.020 2370.390 ;
        RECT 2582.470 2370.380 2584.070 2370.390 ;
        RECT 2722.020 2370.380 2725.020 2370.390 ;
        RECT 2902.020 2370.380 2905.020 2370.390 ;
        RECT 2936.000 2370.380 2939.000 2370.390 ;
        RECT -24.080 2367.380 2943.700 2370.380 ;
        RECT -19.380 2367.370 -16.380 2367.380 ;
        RECT 22.020 2367.370 25.020 2367.380 ;
        RECT 202.020 2367.370 205.020 2367.380 ;
        RECT 682.470 2367.370 684.070 2367.380 ;
        RECT 742.020 2367.370 745.020 2367.380 ;
        RECT 922.020 2367.370 925.020 2367.380 ;
        RECT 1332.470 2367.370 1334.070 2367.380 ;
        RECT 1462.020 2367.370 1465.020 2367.380 ;
        RECT 1932.470 2367.370 1934.070 2367.380 ;
        RECT 2002.020 2367.370 2005.020 2367.380 ;
        RECT 2582.470 2367.370 2584.070 2367.380 ;
        RECT 2722.020 2367.370 2725.020 2367.380 ;
        RECT 2902.020 2367.370 2905.020 2367.380 ;
        RECT 2936.000 2367.370 2939.000 2367.380 ;
        RECT -9.980 2352.380 -6.980 2352.390 ;
        RECT 4.020 2352.380 7.020 2352.390 ;
        RECT 184.020 2352.380 187.020 2352.390 ;
        RECT 682.470 2352.380 684.070 2352.390 ;
        RECT 724.020 2352.380 727.020 2352.390 ;
        RECT 904.020 2352.380 907.020 2352.390 ;
        RECT 1332.470 2352.380 1334.070 2352.390 ;
        RECT 1444.020 2352.380 1447.020 2352.390 ;
        RECT 1932.470 2352.380 1934.070 2352.390 ;
        RECT 1984.020 2352.380 1987.020 2352.390 ;
        RECT 2164.020 2352.380 2167.020 2352.390 ;
        RECT 2582.470 2352.380 2584.070 2352.390 ;
        RECT 2704.020 2352.380 2707.020 2352.390 ;
        RECT 2884.020 2352.380 2887.020 2352.390 ;
        RECT 2926.600 2352.380 2929.600 2352.390 ;
        RECT -14.680 2349.380 2934.300 2352.380 ;
        RECT -9.980 2349.370 -6.980 2349.380 ;
        RECT 4.020 2349.370 7.020 2349.380 ;
        RECT 184.020 2349.370 187.020 2349.380 ;
        RECT 682.470 2349.370 684.070 2349.380 ;
        RECT 724.020 2349.370 727.020 2349.380 ;
        RECT 904.020 2349.370 907.020 2349.380 ;
        RECT 1332.470 2349.370 1334.070 2349.380 ;
        RECT 1444.020 2349.370 1447.020 2349.380 ;
        RECT 1932.470 2349.370 1934.070 2349.380 ;
        RECT 1984.020 2349.370 1987.020 2349.380 ;
        RECT 2164.020 2349.370 2167.020 2349.380 ;
        RECT 2582.470 2349.370 2584.070 2349.380 ;
        RECT 2704.020 2349.370 2707.020 2349.380 ;
        RECT 2884.020 2349.370 2887.020 2349.380 ;
        RECT 2926.600 2349.370 2929.600 2349.380 ;
        RECT -38.180 2226.380 -35.180 2226.390 ;
        RECT 58.020 2226.380 61.020 2226.390 ;
        RECT 238.020 2226.380 241.020 2226.390 ;
        RECT 418.020 2226.380 421.020 2226.390 ;
        RECT 598.020 2226.380 601.020 2226.390 ;
        RECT 778.020 2226.380 781.020 2226.390 ;
        RECT 958.020 2226.380 961.020 2226.390 ;
        RECT 1138.020 2226.380 1141.020 2226.390 ;
        RECT 1318.020 2226.380 1321.020 2226.390 ;
        RECT 1498.020 2226.380 1501.020 2226.390 ;
        RECT 1678.020 2226.380 1681.020 2226.390 ;
        RECT 1858.020 2226.380 1861.020 2226.390 ;
        RECT 2038.020 2226.380 2041.020 2226.390 ;
        RECT 2218.020 2226.380 2221.020 2226.390 ;
        RECT 2398.020 2226.380 2401.020 2226.390 ;
        RECT 2578.020 2226.380 2581.020 2226.390 ;
        RECT 2758.020 2226.380 2761.020 2226.390 ;
        RECT 2954.800 2226.380 2957.800 2226.390 ;
        RECT -42.880 2223.380 2962.500 2226.380 ;
        RECT -38.180 2223.370 -35.180 2223.380 ;
        RECT 58.020 2223.370 61.020 2223.380 ;
        RECT 238.020 2223.370 241.020 2223.380 ;
        RECT 418.020 2223.370 421.020 2223.380 ;
        RECT 598.020 2223.370 601.020 2223.380 ;
        RECT 778.020 2223.370 781.020 2223.380 ;
        RECT 958.020 2223.370 961.020 2223.380 ;
        RECT 1138.020 2223.370 1141.020 2223.380 ;
        RECT 1318.020 2223.370 1321.020 2223.380 ;
        RECT 1498.020 2223.370 1501.020 2223.380 ;
        RECT 1678.020 2223.370 1681.020 2223.380 ;
        RECT 1858.020 2223.370 1861.020 2223.380 ;
        RECT 2038.020 2223.370 2041.020 2223.380 ;
        RECT 2218.020 2223.370 2221.020 2223.380 ;
        RECT 2398.020 2223.370 2401.020 2223.380 ;
        RECT 2578.020 2223.370 2581.020 2223.380 ;
        RECT 2758.020 2223.370 2761.020 2223.380 ;
        RECT 2954.800 2223.370 2957.800 2223.380 ;
        RECT -28.780 2208.380 -25.780 2208.390 ;
        RECT 40.020 2208.380 43.020 2208.390 ;
        RECT 220.020 2208.380 223.020 2208.390 ;
        RECT 1660.020 2208.380 1663.020 2208.390 ;
        RECT 1840.020 2208.380 1843.020 2208.390 ;
        RECT 2020.020 2208.380 2023.020 2208.390 ;
        RECT 2200.020 2208.380 2203.020 2208.390 ;
        RECT 2380.020 2208.380 2383.020 2208.390 ;
        RECT 2560.020 2208.380 2563.020 2208.390 ;
        RECT 2740.020 2208.380 2743.020 2208.390 ;
        RECT 2945.400 2208.380 2948.400 2208.390 ;
        RECT -33.480 2205.380 2953.100 2208.380 ;
        RECT -28.780 2205.370 -25.780 2205.380 ;
        RECT 40.020 2205.370 43.020 2205.380 ;
        RECT 220.020 2205.370 223.020 2205.380 ;
        RECT 1660.020 2205.370 1663.020 2205.380 ;
        RECT 1840.020 2205.370 1843.020 2205.380 ;
        RECT 2020.020 2205.370 2023.020 2205.380 ;
        RECT 2200.020 2205.370 2203.020 2205.380 ;
        RECT 2380.020 2205.370 2383.020 2205.380 ;
        RECT 2560.020 2205.370 2563.020 2205.380 ;
        RECT 2740.020 2205.370 2743.020 2205.380 ;
        RECT 2945.400 2205.370 2948.400 2205.380 ;
        RECT -19.380 2190.380 -16.380 2190.390 ;
        RECT 22.020 2190.380 25.020 2190.390 ;
        RECT 202.020 2190.380 205.020 2190.390 ;
        RECT 1642.020 2190.380 1645.020 2190.390 ;
        RECT 1822.020 2190.380 1825.020 2190.390 ;
        RECT 2002.020 2190.380 2005.020 2190.390 ;
        RECT 2182.020 2190.380 2185.020 2190.390 ;
        RECT 2362.020 2190.380 2365.020 2190.390 ;
        RECT 2542.020 2190.380 2545.020 2190.390 ;
        RECT 2722.020 2190.380 2725.020 2190.390 ;
        RECT 2902.020 2190.380 2905.020 2190.390 ;
        RECT 2936.000 2190.380 2939.000 2190.390 ;
        RECT -24.080 2187.380 2943.700 2190.380 ;
        RECT -19.380 2187.370 -16.380 2187.380 ;
        RECT 22.020 2187.370 25.020 2187.380 ;
        RECT 202.020 2187.370 205.020 2187.380 ;
        RECT 1642.020 2187.370 1645.020 2187.380 ;
        RECT 1822.020 2187.370 1825.020 2187.380 ;
        RECT 2002.020 2187.370 2005.020 2187.380 ;
        RECT 2182.020 2187.370 2185.020 2187.380 ;
        RECT 2362.020 2187.370 2365.020 2187.380 ;
        RECT 2542.020 2187.370 2545.020 2187.380 ;
        RECT 2722.020 2187.370 2725.020 2187.380 ;
        RECT 2902.020 2187.370 2905.020 2187.380 ;
        RECT 2936.000 2187.370 2939.000 2187.380 ;
        RECT -9.980 2172.380 -6.980 2172.390 ;
        RECT 4.020 2172.380 7.020 2172.390 ;
        RECT 184.020 2172.380 187.020 2172.390 ;
        RECT 321.040 2172.380 322.640 2172.390 ;
        RECT 1624.020 2172.380 1627.020 2172.390 ;
        RECT 1804.020 2172.380 1807.020 2172.390 ;
        RECT 1984.020 2172.380 1987.020 2172.390 ;
        RECT 2164.020 2172.380 2167.020 2172.390 ;
        RECT 2344.020 2172.380 2347.020 2172.390 ;
        RECT 2524.020 2172.380 2527.020 2172.390 ;
        RECT 2704.020 2172.380 2707.020 2172.390 ;
        RECT 2884.020 2172.380 2887.020 2172.390 ;
        RECT 2926.600 2172.380 2929.600 2172.390 ;
        RECT -14.680 2169.380 2934.300 2172.380 ;
        RECT -9.980 2169.370 -6.980 2169.380 ;
        RECT 4.020 2169.370 7.020 2169.380 ;
        RECT 184.020 2169.370 187.020 2169.380 ;
        RECT 321.040 2169.370 322.640 2169.380 ;
        RECT 1624.020 2169.370 1627.020 2169.380 ;
        RECT 1804.020 2169.370 1807.020 2169.380 ;
        RECT 1984.020 2169.370 1987.020 2169.380 ;
        RECT 2164.020 2169.370 2167.020 2169.380 ;
        RECT 2344.020 2169.370 2347.020 2169.380 ;
        RECT 2524.020 2169.370 2527.020 2169.380 ;
        RECT 2704.020 2169.370 2707.020 2169.380 ;
        RECT 2884.020 2169.370 2887.020 2169.380 ;
        RECT 2926.600 2169.370 2929.600 2169.380 ;
        RECT -38.180 2046.380 -35.180 2046.390 ;
        RECT 58.020 2046.380 61.020 2046.390 ;
        RECT 238.020 2046.380 241.020 2046.390 ;
        RECT 321.040 2046.380 322.640 2046.390 ;
        RECT 1678.020 2046.380 1681.020 2046.390 ;
        RECT 1858.020 2046.380 1861.020 2046.390 ;
        RECT 2038.020 2046.380 2041.020 2046.390 ;
        RECT 2218.020 2046.380 2221.020 2046.390 ;
        RECT 2398.020 2046.380 2401.020 2046.390 ;
        RECT 2578.020 2046.380 2581.020 2046.390 ;
        RECT 2758.020 2046.380 2761.020 2046.390 ;
        RECT 2954.800 2046.380 2957.800 2046.390 ;
        RECT -42.880 2043.380 2962.500 2046.380 ;
        RECT -38.180 2043.370 -35.180 2043.380 ;
        RECT 58.020 2043.370 61.020 2043.380 ;
        RECT 238.020 2043.370 241.020 2043.380 ;
        RECT 321.040 2043.370 322.640 2043.380 ;
        RECT 1678.020 2043.370 1681.020 2043.380 ;
        RECT 1858.020 2043.370 1861.020 2043.380 ;
        RECT 2038.020 2043.370 2041.020 2043.380 ;
        RECT 2218.020 2043.370 2221.020 2043.380 ;
        RECT 2398.020 2043.370 2401.020 2043.380 ;
        RECT 2578.020 2043.370 2581.020 2043.380 ;
        RECT 2758.020 2043.370 2761.020 2043.380 ;
        RECT 2954.800 2043.370 2957.800 2043.380 ;
        RECT -28.780 2028.380 -25.780 2028.390 ;
        RECT 40.020 2028.380 43.020 2028.390 ;
        RECT 220.020 2028.380 223.020 2028.390 ;
        RECT 321.040 2028.380 322.640 2028.390 ;
        RECT 1660.020 2028.380 1663.020 2028.390 ;
        RECT 1840.020 2028.380 1843.020 2028.390 ;
        RECT 2020.020 2028.380 2023.020 2028.390 ;
        RECT 2200.020 2028.380 2203.020 2028.390 ;
        RECT 2380.020 2028.380 2383.020 2028.390 ;
        RECT 2560.020 2028.380 2563.020 2028.390 ;
        RECT 2740.020 2028.380 2743.020 2028.390 ;
        RECT 2945.400 2028.380 2948.400 2028.390 ;
        RECT -33.480 2025.380 2953.100 2028.380 ;
        RECT -28.780 2025.370 -25.780 2025.380 ;
        RECT 40.020 2025.370 43.020 2025.380 ;
        RECT 220.020 2025.370 223.020 2025.380 ;
        RECT 321.040 2025.370 322.640 2025.380 ;
        RECT 1660.020 2025.370 1663.020 2025.380 ;
        RECT 1840.020 2025.370 1843.020 2025.380 ;
        RECT 2020.020 2025.370 2023.020 2025.380 ;
        RECT 2200.020 2025.370 2203.020 2025.380 ;
        RECT 2380.020 2025.370 2383.020 2025.380 ;
        RECT 2560.020 2025.370 2563.020 2025.380 ;
        RECT 2740.020 2025.370 2743.020 2025.380 ;
        RECT 2945.400 2025.370 2948.400 2025.380 ;
        RECT -19.380 2010.380 -16.380 2010.390 ;
        RECT 22.020 2010.380 25.020 2010.390 ;
        RECT 202.020 2010.380 205.020 2010.390 ;
        RECT 321.040 2010.380 322.640 2010.390 ;
        RECT 1642.020 2010.380 1645.020 2010.390 ;
        RECT 1822.020 2010.380 1825.020 2010.390 ;
        RECT 2002.020 2010.380 2005.020 2010.390 ;
        RECT 2182.020 2010.380 2185.020 2010.390 ;
        RECT 2362.020 2010.380 2365.020 2010.390 ;
        RECT 2542.020 2010.380 2545.020 2010.390 ;
        RECT 2722.020 2010.380 2725.020 2010.390 ;
        RECT 2902.020 2010.380 2905.020 2010.390 ;
        RECT 2936.000 2010.380 2939.000 2010.390 ;
        RECT -24.080 2007.380 2943.700 2010.380 ;
        RECT -19.380 2007.370 -16.380 2007.380 ;
        RECT 22.020 2007.370 25.020 2007.380 ;
        RECT 202.020 2007.370 205.020 2007.380 ;
        RECT 321.040 2007.370 322.640 2007.380 ;
        RECT 1642.020 2007.370 1645.020 2007.380 ;
        RECT 1822.020 2007.370 1825.020 2007.380 ;
        RECT 2002.020 2007.370 2005.020 2007.380 ;
        RECT 2182.020 2007.370 2185.020 2007.380 ;
        RECT 2362.020 2007.370 2365.020 2007.380 ;
        RECT 2542.020 2007.370 2545.020 2007.380 ;
        RECT 2722.020 2007.370 2725.020 2007.380 ;
        RECT 2902.020 2007.370 2905.020 2007.380 ;
        RECT 2936.000 2007.370 2939.000 2007.380 ;
        RECT -9.980 1992.380 -6.980 1992.390 ;
        RECT 4.020 1992.380 7.020 1992.390 ;
        RECT 184.020 1992.380 187.020 1992.390 ;
        RECT 321.040 1992.380 322.640 1992.390 ;
        RECT 1624.020 1992.380 1627.020 1992.390 ;
        RECT 1804.020 1992.380 1807.020 1992.390 ;
        RECT 1984.020 1992.380 1987.020 1992.390 ;
        RECT 2164.020 1992.380 2167.020 1992.390 ;
        RECT 2344.020 1992.380 2347.020 1992.390 ;
        RECT 2524.020 1992.380 2527.020 1992.390 ;
        RECT 2704.020 1992.380 2707.020 1992.390 ;
        RECT 2884.020 1992.380 2887.020 1992.390 ;
        RECT 2926.600 1992.380 2929.600 1992.390 ;
        RECT -14.680 1989.380 2934.300 1992.380 ;
        RECT -9.980 1989.370 -6.980 1989.380 ;
        RECT 4.020 1989.370 7.020 1989.380 ;
        RECT 184.020 1989.370 187.020 1989.380 ;
        RECT 321.040 1989.370 322.640 1989.380 ;
        RECT 1624.020 1989.370 1627.020 1989.380 ;
        RECT 1804.020 1989.370 1807.020 1989.380 ;
        RECT 1984.020 1989.370 1987.020 1989.380 ;
        RECT 2164.020 1989.370 2167.020 1989.380 ;
        RECT 2344.020 1989.370 2347.020 1989.380 ;
        RECT 2524.020 1989.370 2527.020 1989.380 ;
        RECT 2704.020 1989.370 2707.020 1989.380 ;
        RECT 2884.020 1989.370 2887.020 1989.380 ;
        RECT 2926.600 1989.370 2929.600 1989.380 ;
        RECT -38.180 1866.380 -35.180 1866.390 ;
        RECT 58.020 1866.380 61.020 1866.390 ;
        RECT 238.020 1866.380 241.020 1866.390 ;
        RECT 321.040 1866.380 322.640 1866.390 ;
        RECT 1678.020 1866.380 1681.020 1866.390 ;
        RECT 1858.020 1866.380 1861.020 1866.390 ;
        RECT 2038.020 1866.380 2041.020 1866.390 ;
        RECT 2218.020 1866.380 2221.020 1866.390 ;
        RECT 2398.020 1866.380 2401.020 1866.390 ;
        RECT 2578.020 1866.380 2581.020 1866.390 ;
        RECT 2758.020 1866.380 2761.020 1866.390 ;
        RECT 2954.800 1866.380 2957.800 1866.390 ;
        RECT -42.880 1863.380 2962.500 1866.380 ;
        RECT -38.180 1863.370 -35.180 1863.380 ;
        RECT 58.020 1863.370 61.020 1863.380 ;
        RECT 238.020 1863.370 241.020 1863.380 ;
        RECT 321.040 1863.370 322.640 1863.380 ;
        RECT 1678.020 1863.370 1681.020 1863.380 ;
        RECT 1858.020 1863.370 1861.020 1863.380 ;
        RECT 2038.020 1863.370 2041.020 1863.380 ;
        RECT 2218.020 1863.370 2221.020 1863.380 ;
        RECT 2398.020 1863.370 2401.020 1863.380 ;
        RECT 2578.020 1863.370 2581.020 1863.380 ;
        RECT 2758.020 1863.370 2761.020 1863.380 ;
        RECT 2954.800 1863.370 2957.800 1863.380 ;
        RECT -28.780 1848.380 -25.780 1848.390 ;
        RECT 40.020 1848.380 43.020 1848.390 ;
        RECT 220.020 1848.380 223.020 1848.390 ;
        RECT 321.040 1848.380 322.640 1848.390 ;
        RECT 1660.020 1848.380 1663.020 1848.390 ;
        RECT 1840.020 1848.380 1843.020 1848.390 ;
        RECT 2020.020 1848.380 2023.020 1848.390 ;
        RECT 2200.020 1848.380 2203.020 1848.390 ;
        RECT 2380.020 1848.380 2383.020 1848.390 ;
        RECT 2560.020 1848.380 2563.020 1848.390 ;
        RECT 2740.020 1848.380 2743.020 1848.390 ;
        RECT 2945.400 1848.380 2948.400 1848.390 ;
        RECT -33.480 1845.380 2953.100 1848.380 ;
        RECT -28.780 1845.370 -25.780 1845.380 ;
        RECT 40.020 1845.370 43.020 1845.380 ;
        RECT 220.020 1845.370 223.020 1845.380 ;
        RECT 321.040 1845.370 322.640 1845.380 ;
        RECT 1660.020 1845.370 1663.020 1845.380 ;
        RECT 1840.020 1845.370 1843.020 1845.380 ;
        RECT 2020.020 1845.370 2023.020 1845.380 ;
        RECT 2200.020 1845.370 2203.020 1845.380 ;
        RECT 2380.020 1845.370 2383.020 1845.380 ;
        RECT 2560.020 1845.370 2563.020 1845.380 ;
        RECT 2740.020 1845.370 2743.020 1845.380 ;
        RECT 2945.400 1845.370 2948.400 1845.380 ;
        RECT -19.380 1830.380 -16.380 1830.390 ;
        RECT 22.020 1830.380 25.020 1830.390 ;
        RECT 202.020 1830.380 205.020 1830.390 ;
        RECT 321.040 1830.380 322.640 1830.390 ;
        RECT 1642.020 1830.380 1645.020 1830.390 ;
        RECT 1822.020 1830.380 1825.020 1830.390 ;
        RECT 2002.020 1830.380 2005.020 1830.390 ;
        RECT 2182.020 1830.380 2185.020 1830.390 ;
        RECT 2362.020 1830.380 2365.020 1830.390 ;
        RECT 2542.020 1830.380 2545.020 1830.390 ;
        RECT 2722.020 1830.380 2725.020 1830.390 ;
        RECT 2902.020 1830.380 2905.020 1830.390 ;
        RECT 2936.000 1830.380 2939.000 1830.390 ;
        RECT -24.080 1827.380 2943.700 1830.380 ;
        RECT -19.380 1827.370 -16.380 1827.380 ;
        RECT 22.020 1827.370 25.020 1827.380 ;
        RECT 202.020 1827.370 205.020 1827.380 ;
        RECT 321.040 1827.370 322.640 1827.380 ;
        RECT 1642.020 1827.370 1645.020 1827.380 ;
        RECT 1822.020 1827.370 1825.020 1827.380 ;
        RECT 2002.020 1827.370 2005.020 1827.380 ;
        RECT 2182.020 1827.370 2185.020 1827.380 ;
        RECT 2362.020 1827.370 2365.020 1827.380 ;
        RECT 2542.020 1827.370 2545.020 1827.380 ;
        RECT 2722.020 1827.370 2725.020 1827.380 ;
        RECT 2902.020 1827.370 2905.020 1827.380 ;
        RECT 2936.000 1827.370 2939.000 1827.380 ;
        RECT -9.980 1812.380 -6.980 1812.390 ;
        RECT 4.020 1812.380 7.020 1812.390 ;
        RECT 184.020 1812.380 187.020 1812.390 ;
        RECT 321.040 1812.380 322.640 1812.390 ;
        RECT 1624.020 1812.380 1627.020 1812.390 ;
        RECT 1804.020 1812.380 1807.020 1812.390 ;
        RECT 1984.020 1812.380 1987.020 1812.390 ;
        RECT 2164.020 1812.380 2167.020 1812.390 ;
        RECT 2344.020 1812.380 2347.020 1812.390 ;
        RECT 2524.020 1812.380 2527.020 1812.390 ;
        RECT 2704.020 1812.380 2707.020 1812.390 ;
        RECT 2884.020 1812.380 2887.020 1812.390 ;
        RECT 2926.600 1812.380 2929.600 1812.390 ;
        RECT -14.680 1809.380 2934.300 1812.380 ;
        RECT -9.980 1809.370 -6.980 1809.380 ;
        RECT 4.020 1809.370 7.020 1809.380 ;
        RECT 184.020 1809.370 187.020 1809.380 ;
        RECT 321.040 1809.370 322.640 1809.380 ;
        RECT 1624.020 1809.370 1627.020 1809.380 ;
        RECT 1804.020 1809.370 1807.020 1809.380 ;
        RECT 1984.020 1809.370 1987.020 1809.380 ;
        RECT 2164.020 1809.370 2167.020 1809.380 ;
        RECT 2344.020 1809.370 2347.020 1809.380 ;
        RECT 2524.020 1809.370 2527.020 1809.380 ;
        RECT 2704.020 1809.370 2707.020 1809.380 ;
        RECT 2884.020 1809.370 2887.020 1809.380 ;
        RECT 2926.600 1809.370 2929.600 1809.380 ;
        RECT -38.180 1686.380 -35.180 1686.390 ;
        RECT 58.020 1686.380 61.020 1686.390 ;
        RECT 238.020 1686.380 241.020 1686.390 ;
        RECT 321.040 1686.380 322.640 1686.390 ;
        RECT 1678.020 1686.380 1681.020 1686.390 ;
        RECT 1858.020 1686.380 1861.020 1686.390 ;
        RECT 2038.020 1686.380 2041.020 1686.390 ;
        RECT 2218.020 1686.380 2221.020 1686.390 ;
        RECT 2398.020 1686.380 2401.020 1686.390 ;
        RECT 2578.020 1686.380 2581.020 1686.390 ;
        RECT 2758.020 1686.380 2761.020 1686.390 ;
        RECT 2954.800 1686.380 2957.800 1686.390 ;
        RECT -42.880 1683.380 2962.500 1686.380 ;
        RECT -38.180 1683.370 -35.180 1683.380 ;
        RECT 58.020 1683.370 61.020 1683.380 ;
        RECT 238.020 1683.370 241.020 1683.380 ;
        RECT 321.040 1683.370 322.640 1683.380 ;
        RECT 1678.020 1683.370 1681.020 1683.380 ;
        RECT 1858.020 1683.370 1861.020 1683.380 ;
        RECT 2038.020 1683.370 2041.020 1683.380 ;
        RECT 2218.020 1683.370 2221.020 1683.380 ;
        RECT 2398.020 1683.370 2401.020 1683.380 ;
        RECT 2578.020 1683.370 2581.020 1683.380 ;
        RECT 2758.020 1683.370 2761.020 1683.380 ;
        RECT 2954.800 1683.370 2957.800 1683.380 ;
        RECT -28.780 1668.380 -25.780 1668.390 ;
        RECT 40.020 1668.380 43.020 1668.390 ;
        RECT 220.020 1668.380 223.020 1668.390 ;
        RECT 321.040 1668.380 322.640 1668.390 ;
        RECT 1660.020 1668.380 1663.020 1668.390 ;
        RECT 1840.020 1668.380 1843.020 1668.390 ;
        RECT 2020.020 1668.380 2023.020 1668.390 ;
        RECT 2200.020 1668.380 2203.020 1668.390 ;
        RECT 2380.020 1668.380 2383.020 1668.390 ;
        RECT 2560.020 1668.380 2563.020 1668.390 ;
        RECT 2740.020 1668.380 2743.020 1668.390 ;
        RECT 2945.400 1668.380 2948.400 1668.390 ;
        RECT -33.480 1665.380 2953.100 1668.380 ;
        RECT -28.780 1665.370 -25.780 1665.380 ;
        RECT 40.020 1665.370 43.020 1665.380 ;
        RECT 220.020 1665.370 223.020 1665.380 ;
        RECT 321.040 1665.370 322.640 1665.380 ;
        RECT 1660.020 1665.370 1663.020 1665.380 ;
        RECT 1840.020 1665.370 1843.020 1665.380 ;
        RECT 2020.020 1665.370 2023.020 1665.380 ;
        RECT 2200.020 1665.370 2203.020 1665.380 ;
        RECT 2380.020 1665.370 2383.020 1665.380 ;
        RECT 2560.020 1665.370 2563.020 1665.380 ;
        RECT 2740.020 1665.370 2743.020 1665.380 ;
        RECT 2945.400 1665.370 2948.400 1665.380 ;
        RECT -19.380 1650.380 -16.380 1650.390 ;
        RECT 22.020 1650.380 25.020 1650.390 ;
        RECT 202.020 1650.380 205.020 1650.390 ;
        RECT 321.040 1650.380 322.640 1650.390 ;
        RECT 1642.020 1650.380 1645.020 1650.390 ;
        RECT 1822.020 1650.380 1825.020 1650.390 ;
        RECT 2002.020 1650.380 2005.020 1650.390 ;
        RECT 2182.020 1650.380 2185.020 1650.390 ;
        RECT 2362.020 1650.380 2365.020 1650.390 ;
        RECT 2542.020 1650.380 2545.020 1650.390 ;
        RECT 2722.020 1650.380 2725.020 1650.390 ;
        RECT 2902.020 1650.380 2905.020 1650.390 ;
        RECT 2936.000 1650.380 2939.000 1650.390 ;
        RECT -24.080 1647.380 2943.700 1650.380 ;
        RECT -19.380 1647.370 -16.380 1647.380 ;
        RECT 22.020 1647.370 25.020 1647.380 ;
        RECT 202.020 1647.370 205.020 1647.380 ;
        RECT 321.040 1647.370 322.640 1647.380 ;
        RECT 1642.020 1647.370 1645.020 1647.380 ;
        RECT 1822.020 1647.370 1825.020 1647.380 ;
        RECT 2002.020 1647.370 2005.020 1647.380 ;
        RECT 2182.020 1647.370 2185.020 1647.380 ;
        RECT 2362.020 1647.370 2365.020 1647.380 ;
        RECT 2542.020 1647.370 2545.020 1647.380 ;
        RECT 2722.020 1647.370 2725.020 1647.380 ;
        RECT 2902.020 1647.370 2905.020 1647.380 ;
        RECT 2936.000 1647.370 2939.000 1647.380 ;
        RECT -9.980 1632.380 -6.980 1632.390 ;
        RECT 4.020 1632.380 7.020 1632.390 ;
        RECT 184.020 1632.380 187.020 1632.390 ;
        RECT 321.040 1632.380 322.640 1632.390 ;
        RECT 1624.020 1632.380 1627.020 1632.390 ;
        RECT 1804.020 1632.380 1807.020 1632.390 ;
        RECT 1984.020 1632.380 1987.020 1632.390 ;
        RECT 2164.020 1632.380 2167.020 1632.390 ;
        RECT 2344.020 1632.380 2347.020 1632.390 ;
        RECT 2524.020 1632.380 2527.020 1632.390 ;
        RECT 2704.020 1632.380 2707.020 1632.390 ;
        RECT 2884.020 1632.380 2887.020 1632.390 ;
        RECT 2926.600 1632.380 2929.600 1632.390 ;
        RECT -14.680 1629.380 2934.300 1632.380 ;
        RECT -9.980 1629.370 -6.980 1629.380 ;
        RECT 4.020 1629.370 7.020 1629.380 ;
        RECT 184.020 1629.370 187.020 1629.380 ;
        RECT 321.040 1629.370 322.640 1629.380 ;
        RECT 1624.020 1629.370 1627.020 1629.380 ;
        RECT 1804.020 1629.370 1807.020 1629.380 ;
        RECT 1984.020 1629.370 1987.020 1629.380 ;
        RECT 2164.020 1629.370 2167.020 1629.380 ;
        RECT 2344.020 1629.370 2347.020 1629.380 ;
        RECT 2524.020 1629.370 2527.020 1629.380 ;
        RECT 2704.020 1629.370 2707.020 1629.380 ;
        RECT 2884.020 1629.370 2887.020 1629.380 ;
        RECT 2926.600 1629.370 2929.600 1629.380 ;
        RECT -38.180 1506.380 -35.180 1506.390 ;
        RECT 58.020 1506.380 61.020 1506.390 ;
        RECT 238.020 1506.380 241.020 1506.390 ;
        RECT 321.040 1506.380 322.640 1506.390 ;
        RECT 1678.020 1506.380 1681.020 1506.390 ;
        RECT 1858.020 1506.380 1861.020 1506.390 ;
        RECT 2038.020 1506.380 2041.020 1506.390 ;
        RECT 2218.020 1506.380 2221.020 1506.390 ;
        RECT 2398.020 1506.380 2401.020 1506.390 ;
        RECT 2578.020 1506.380 2581.020 1506.390 ;
        RECT 2758.020 1506.380 2761.020 1506.390 ;
        RECT 2954.800 1506.380 2957.800 1506.390 ;
        RECT -42.880 1503.380 2962.500 1506.380 ;
        RECT -38.180 1503.370 -35.180 1503.380 ;
        RECT 58.020 1503.370 61.020 1503.380 ;
        RECT 238.020 1503.370 241.020 1503.380 ;
        RECT 321.040 1503.370 322.640 1503.380 ;
        RECT 1678.020 1503.370 1681.020 1503.380 ;
        RECT 1858.020 1503.370 1861.020 1503.380 ;
        RECT 2038.020 1503.370 2041.020 1503.380 ;
        RECT 2218.020 1503.370 2221.020 1503.380 ;
        RECT 2398.020 1503.370 2401.020 1503.380 ;
        RECT 2578.020 1503.370 2581.020 1503.380 ;
        RECT 2758.020 1503.370 2761.020 1503.380 ;
        RECT 2954.800 1503.370 2957.800 1503.380 ;
        RECT -28.780 1488.380 -25.780 1488.390 ;
        RECT 40.020 1488.380 43.020 1488.390 ;
        RECT 220.020 1488.380 223.020 1488.390 ;
        RECT 321.040 1488.380 322.640 1488.390 ;
        RECT 1660.020 1488.380 1663.020 1488.390 ;
        RECT 1840.020 1488.380 1843.020 1488.390 ;
        RECT 2020.020 1488.380 2023.020 1488.390 ;
        RECT 2200.020 1488.380 2203.020 1488.390 ;
        RECT 2380.020 1488.380 2383.020 1488.390 ;
        RECT 2560.020 1488.380 2563.020 1488.390 ;
        RECT 2740.020 1488.380 2743.020 1488.390 ;
        RECT 2945.400 1488.380 2948.400 1488.390 ;
        RECT -33.480 1485.380 2953.100 1488.380 ;
        RECT -28.780 1485.370 -25.780 1485.380 ;
        RECT 40.020 1485.370 43.020 1485.380 ;
        RECT 220.020 1485.370 223.020 1485.380 ;
        RECT 321.040 1485.370 322.640 1485.380 ;
        RECT 1660.020 1485.370 1663.020 1485.380 ;
        RECT 1840.020 1485.370 1843.020 1485.380 ;
        RECT 2020.020 1485.370 2023.020 1485.380 ;
        RECT 2200.020 1485.370 2203.020 1485.380 ;
        RECT 2380.020 1485.370 2383.020 1485.380 ;
        RECT 2560.020 1485.370 2563.020 1485.380 ;
        RECT 2740.020 1485.370 2743.020 1485.380 ;
        RECT 2945.400 1485.370 2948.400 1485.380 ;
        RECT -19.380 1470.380 -16.380 1470.390 ;
        RECT 22.020 1470.380 25.020 1470.390 ;
        RECT 202.020 1470.380 205.020 1470.390 ;
        RECT 321.040 1470.380 322.640 1470.390 ;
        RECT 1642.020 1470.380 1645.020 1470.390 ;
        RECT 1822.020 1470.380 1825.020 1470.390 ;
        RECT 2002.020 1470.380 2005.020 1470.390 ;
        RECT 2182.020 1470.380 2185.020 1470.390 ;
        RECT 2362.020 1470.380 2365.020 1470.390 ;
        RECT 2542.020 1470.380 2545.020 1470.390 ;
        RECT 2722.020 1470.380 2725.020 1470.390 ;
        RECT 2902.020 1470.380 2905.020 1470.390 ;
        RECT 2936.000 1470.380 2939.000 1470.390 ;
        RECT -24.080 1467.380 2943.700 1470.380 ;
        RECT -19.380 1467.370 -16.380 1467.380 ;
        RECT 22.020 1467.370 25.020 1467.380 ;
        RECT 202.020 1467.370 205.020 1467.380 ;
        RECT 321.040 1467.370 322.640 1467.380 ;
        RECT 1642.020 1467.370 1645.020 1467.380 ;
        RECT 1822.020 1467.370 1825.020 1467.380 ;
        RECT 2002.020 1467.370 2005.020 1467.380 ;
        RECT 2182.020 1467.370 2185.020 1467.380 ;
        RECT 2362.020 1467.370 2365.020 1467.380 ;
        RECT 2542.020 1467.370 2545.020 1467.380 ;
        RECT 2722.020 1467.370 2725.020 1467.380 ;
        RECT 2902.020 1467.370 2905.020 1467.380 ;
        RECT 2936.000 1467.370 2939.000 1467.380 ;
        RECT -9.980 1452.380 -6.980 1452.390 ;
        RECT 4.020 1452.380 7.020 1452.390 ;
        RECT 184.020 1452.380 187.020 1452.390 ;
        RECT 321.040 1452.380 322.640 1452.390 ;
        RECT 1624.020 1452.380 1627.020 1452.390 ;
        RECT 1804.020 1452.380 1807.020 1452.390 ;
        RECT 1984.020 1452.380 1987.020 1452.390 ;
        RECT 2164.020 1452.380 2167.020 1452.390 ;
        RECT 2344.020 1452.380 2347.020 1452.390 ;
        RECT 2524.020 1452.380 2527.020 1452.390 ;
        RECT 2704.020 1452.380 2707.020 1452.390 ;
        RECT 2884.020 1452.380 2887.020 1452.390 ;
        RECT 2926.600 1452.380 2929.600 1452.390 ;
        RECT -14.680 1449.380 2934.300 1452.380 ;
        RECT -9.980 1449.370 -6.980 1449.380 ;
        RECT 4.020 1449.370 7.020 1449.380 ;
        RECT 184.020 1449.370 187.020 1449.380 ;
        RECT 321.040 1449.370 322.640 1449.380 ;
        RECT 1624.020 1449.370 1627.020 1449.380 ;
        RECT 1804.020 1449.370 1807.020 1449.380 ;
        RECT 1984.020 1449.370 1987.020 1449.380 ;
        RECT 2164.020 1449.370 2167.020 1449.380 ;
        RECT 2344.020 1449.370 2347.020 1449.380 ;
        RECT 2524.020 1449.370 2527.020 1449.380 ;
        RECT 2704.020 1449.370 2707.020 1449.380 ;
        RECT 2884.020 1449.370 2887.020 1449.380 ;
        RECT 2926.600 1449.370 2929.600 1449.380 ;
        RECT -38.180 1326.380 -35.180 1326.390 ;
        RECT 58.020 1326.380 61.020 1326.390 ;
        RECT 238.020 1326.380 241.020 1326.390 ;
        RECT 321.040 1326.380 322.640 1326.390 ;
        RECT 1678.020 1326.380 1681.020 1326.390 ;
        RECT 1858.020 1326.380 1861.020 1326.390 ;
        RECT 2038.020 1326.380 2041.020 1326.390 ;
        RECT 2218.020 1326.380 2221.020 1326.390 ;
        RECT 2398.020 1326.380 2401.020 1326.390 ;
        RECT 2578.020 1326.380 2581.020 1326.390 ;
        RECT 2758.020 1326.380 2761.020 1326.390 ;
        RECT 2954.800 1326.380 2957.800 1326.390 ;
        RECT -42.880 1323.380 2962.500 1326.380 ;
        RECT -38.180 1323.370 -35.180 1323.380 ;
        RECT 58.020 1323.370 61.020 1323.380 ;
        RECT 238.020 1323.370 241.020 1323.380 ;
        RECT 321.040 1323.370 322.640 1323.380 ;
        RECT 1678.020 1323.370 1681.020 1323.380 ;
        RECT 1858.020 1323.370 1861.020 1323.380 ;
        RECT 2038.020 1323.370 2041.020 1323.380 ;
        RECT 2218.020 1323.370 2221.020 1323.380 ;
        RECT 2398.020 1323.370 2401.020 1323.380 ;
        RECT 2578.020 1323.370 2581.020 1323.380 ;
        RECT 2758.020 1323.370 2761.020 1323.380 ;
        RECT 2954.800 1323.370 2957.800 1323.380 ;
        RECT -28.780 1308.380 -25.780 1308.390 ;
        RECT 40.020 1308.380 43.020 1308.390 ;
        RECT 220.020 1308.380 223.020 1308.390 ;
        RECT 321.040 1308.380 322.640 1308.390 ;
        RECT 1660.020 1308.380 1663.020 1308.390 ;
        RECT 1840.020 1308.380 1843.020 1308.390 ;
        RECT 2020.020 1308.380 2023.020 1308.390 ;
        RECT 2200.020 1308.380 2203.020 1308.390 ;
        RECT 2380.020 1308.380 2383.020 1308.390 ;
        RECT 2560.020 1308.380 2563.020 1308.390 ;
        RECT 2740.020 1308.380 2743.020 1308.390 ;
        RECT 2945.400 1308.380 2948.400 1308.390 ;
        RECT -33.480 1305.380 2953.100 1308.380 ;
        RECT -28.780 1305.370 -25.780 1305.380 ;
        RECT 40.020 1305.370 43.020 1305.380 ;
        RECT 220.020 1305.370 223.020 1305.380 ;
        RECT 321.040 1305.370 322.640 1305.380 ;
        RECT 1660.020 1305.370 1663.020 1305.380 ;
        RECT 1840.020 1305.370 1843.020 1305.380 ;
        RECT 2020.020 1305.370 2023.020 1305.380 ;
        RECT 2200.020 1305.370 2203.020 1305.380 ;
        RECT 2380.020 1305.370 2383.020 1305.380 ;
        RECT 2560.020 1305.370 2563.020 1305.380 ;
        RECT 2740.020 1305.370 2743.020 1305.380 ;
        RECT 2945.400 1305.370 2948.400 1305.380 ;
        RECT -19.380 1290.380 -16.380 1290.390 ;
        RECT 22.020 1290.380 25.020 1290.390 ;
        RECT 202.020 1290.380 205.020 1290.390 ;
        RECT 321.040 1290.380 322.640 1290.390 ;
        RECT 1642.020 1290.380 1645.020 1290.390 ;
        RECT 1822.020 1290.380 1825.020 1290.390 ;
        RECT 2002.020 1290.380 2005.020 1290.390 ;
        RECT 2182.020 1290.380 2185.020 1290.390 ;
        RECT 2362.020 1290.380 2365.020 1290.390 ;
        RECT 2542.020 1290.380 2545.020 1290.390 ;
        RECT 2722.020 1290.380 2725.020 1290.390 ;
        RECT 2902.020 1290.380 2905.020 1290.390 ;
        RECT 2936.000 1290.380 2939.000 1290.390 ;
        RECT -24.080 1287.380 2943.700 1290.380 ;
        RECT -19.380 1287.370 -16.380 1287.380 ;
        RECT 22.020 1287.370 25.020 1287.380 ;
        RECT 202.020 1287.370 205.020 1287.380 ;
        RECT 321.040 1287.370 322.640 1287.380 ;
        RECT 1642.020 1287.370 1645.020 1287.380 ;
        RECT 1822.020 1287.370 1825.020 1287.380 ;
        RECT 2002.020 1287.370 2005.020 1287.380 ;
        RECT 2182.020 1287.370 2185.020 1287.380 ;
        RECT 2362.020 1287.370 2365.020 1287.380 ;
        RECT 2542.020 1287.370 2545.020 1287.380 ;
        RECT 2722.020 1287.370 2725.020 1287.380 ;
        RECT 2902.020 1287.370 2905.020 1287.380 ;
        RECT 2936.000 1287.370 2939.000 1287.380 ;
        RECT -9.980 1272.380 -6.980 1272.390 ;
        RECT 4.020 1272.380 7.020 1272.390 ;
        RECT 184.020 1272.380 187.020 1272.390 ;
        RECT 321.040 1272.380 322.640 1272.390 ;
        RECT 1624.020 1272.380 1627.020 1272.390 ;
        RECT 1804.020 1272.380 1807.020 1272.390 ;
        RECT 1984.020 1272.380 1987.020 1272.390 ;
        RECT 2164.020 1272.380 2167.020 1272.390 ;
        RECT 2344.020 1272.380 2347.020 1272.390 ;
        RECT 2524.020 1272.380 2527.020 1272.390 ;
        RECT 2704.020 1272.380 2707.020 1272.390 ;
        RECT 2884.020 1272.380 2887.020 1272.390 ;
        RECT 2926.600 1272.380 2929.600 1272.390 ;
        RECT -14.680 1269.380 2934.300 1272.380 ;
        RECT -9.980 1269.370 -6.980 1269.380 ;
        RECT 4.020 1269.370 7.020 1269.380 ;
        RECT 184.020 1269.370 187.020 1269.380 ;
        RECT 321.040 1269.370 322.640 1269.380 ;
        RECT 1624.020 1269.370 1627.020 1269.380 ;
        RECT 1804.020 1269.370 1807.020 1269.380 ;
        RECT 1984.020 1269.370 1987.020 1269.380 ;
        RECT 2164.020 1269.370 2167.020 1269.380 ;
        RECT 2344.020 1269.370 2347.020 1269.380 ;
        RECT 2524.020 1269.370 2527.020 1269.380 ;
        RECT 2704.020 1269.370 2707.020 1269.380 ;
        RECT 2884.020 1269.370 2887.020 1269.380 ;
        RECT 2926.600 1269.370 2929.600 1269.380 ;
        RECT -38.180 1146.380 -35.180 1146.390 ;
        RECT 58.020 1146.380 61.020 1146.390 ;
        RECT 238.020 1146.380 241.020 1146.390 ;
        RECT 321.040 1146.380 322.640 1146.390 ;
        RECT 1678.020 1146.380 1681.020 1146.390 ;
        RECT 1858.020 1146.380 1861.020 1146.390 ;
        RECT 2038.020 1146.380 2041.020 1146.390 ;
        RECT 2218.020 1146.380 2221.020 1146.390 ;
        RECT 2398.020 1146.380 2401.020 1146.390 ;
        RECT 2578.020 1146.380 2581.020 1146.390 ;
        RECT 2758.020 1146.380 2761.020 1146.390 ;
        RECT 2954.800 1146.380 2957.800 1146.390 ;
        RECT -42.880 1143.380 2962.500 1146.380 ;
        RECT -38.180 1143.370 -35.180 1143.380 ;
        RECT 58.020 1143.370 61.020 1143.380 ;
        RECT 238.020 1143.370 241.020 1143.380 ;
        RECT 321.040 1143.370 322.640 1143.380 ;
        RECT 1678.020 1143.370 1681.020 1143.380 ;
        RECT 1858.020 1143.370 1861.020 1143.380 ;
        RECT 2038.020 1143.370 2041.020 1143.380 ;
        RECT 2218.020 1143.370 2221.020 1143.380 ;
        RECT 2398.020 1143.370 2401.020 1143.380 ;
        RECT 2578.020 1143.370 2581.020 1143.380 ;
        RECT 2758.020 1143.370 2761.020 1143.380 ;
        RECT 2954.800 1143.370 2957.800 1143.380 ;
        RECT -28.780 1128.380 -25.780 1128.390 ;
        RECT 40.020 1128.380 43.020 1128.390 ;
        RECT 220.020 1128.380 223.020 1128.390 ;
        RECT 321.040 1128.380 322.640 1128.390 ;
        RECT 1660.020 1128.380 1663.020 1128.390 ;
        RECT 1840.020 1128.380 1843.020 1128.390 ;
        RECT 2020.020 1128.380 2023.020 1128.390 ;
        RECT 2200.020 1128.380 2203.020 1128.390 ;
        RECT 2380.020 1128.380 2383.020 1128.390 ;
        RECT 2560.020 1128.380 2563.020 1128.390 ;
        RECT 2740.020 1128.380 2743.020 1128.390 ;
        RECT 2945.400 1128.380 2948.400 1128.390 ;
        RECT -33.480 1125.380 2953.100 1128.380 ;
        RECT -28.780 1125.370 -25.780 1125.380 ;
        RECT 40.020 1125.370 43.020 1125.380 ;
        RECT 220.020 1125.370 223.020 1125.380 ;
        RECT 321.040 1125.370 322.640 1125.380 ;
        RECT 1660.020 1125.370 1663.020 1125.380 ;
        RECT 1840.020 1125.370 1843.020 1125.380 ;
        RECT 2020.020 1125.370 2023.020 1125.380 ;
        RECT 2200.020 1125.370 2203.020 1125.380 ;
        RECT 2380.020 1125.370 2383.020 1125.380 ;
        RECT 2560.020 1125.370 2563.020 1125.380 ;
        RECT 2740.020 1125.370 2743.020 1125.380 ;
        RECT 2945.400 1125.370 2948.400 1125.380 ;
        RECT -19.380 1110.380 -16.380 1110.390 ;
        RECT 22.020 1110.380 25.020 1110.390 ;
        RECT 202.020 1110.380 205.020 1110.390 ;
        RECT 321.040 1110.380 322.640 1110.390 ;
        RECT 1642.020 1110.380 1645.020 1110.390 ;
        RECT 1822.020 1110.380 1825.020 1110.390 ;
        RECT 2002.020 1110.380 2005.020 1110.390 ;
        RECT 2182.020 1110.380 2185.020 1110.390 ;
        RECT 2362.020 1110.380 2365.020 1110.390 ;
        RECT 2542.020 1110.380 2545.020 1110.390 ;
        RECT 2722.020 1110.380 2725.020 1110.390 ;
        RECT 2902.020 1110.380 2905.020 1110.390 ;
        RECT 2936.000 1110.380 2939.000 1110.390 ;
        RECT -24.080 1107.380 2943.700 1110.380 ;
        RECT -19.380 1107.370 -16.380 1107.380 ;
        RECT 22.020 1107.370 25.020 1107.380 ;
        RECT 202.020 1107.370 205.020 1107.380 ;
        RECT 321.040 1107.370 322.640 1107.380 ;
        RECT 1642.020 1107.370 1645.020 1107.380 ;
        RECT 1822.020 1107.370 1825.020 1107.380 ;
        RECT 2002.020 1107.370 2005.020 1107.380 ;
        RECT 2182.020 1107.370 2185.020 1107.380 ;
        RECT 2362.020 1107.370 2365.020 1107.380 ;
        RECT 2542.020 1107.370 2545.020 1107.380 ;
        RECT 2722.020 1107.370 2725.020 1107.380 ;
        RECT 2902.020 1107.370 2905.020 1107.380 ;
        RECT 2936.000 1107.370 2939.000 1107.380 ;
        RECT -9.980 1092.380 -6.980 1092.390 ;
        RECT 4.020 1092.380 7.020 1092.390 ;
        RECT 184.020 1092.380 187.020 1092.390 ;
        RECT 321.040 1092.380 322.640 1092.390 ;
        RECT 1624.020 1092.380 1627.020 1092.390 ;
        RECT 1804.020 1092.380 1807.020 1092.390 ;
        RECT 1984.020 1092.380 1987.020 1092.390 ;
        RECT 2164.020 1092.380 2167.020 1092.390 ;
        RECT 2344.020 1092.380 2347.020 1092.390 ;
        RECT 2524.020 1092.380 2527.020 1092.390 ;
        RECT 2704.020 1092.380 2707.020 1092.390 ;
        RECT 2884.020 1092.380 2887.020 1092.390 ;
        RECT 2926.600 1092.380 2929.600 1092.390 ;
        RECT -14.680 1089.380 2934.300 1092.380 ;
        RECT -9.980 1089.370 -6.980 1089.380 ;
        RECT 4.020 1089.370 7.020 1089.380 ;
        RECT 184.020 1089.370 187.020 1089.380 ;
        RECT 321.040 1089.370 322.640 1089.380 ;
        RECT 1624.020 1089.370 1627.020 1089.380 ;
        RECT 1804.020 1089.370 1807.020 1089.380 ;
        RECT 1984.020 1089.370 1987.020 1089.380 ;
        RECT 2164.020 1089.370 2167.020 1089.380 ;
        RECT 2344.020 1089.370 2347.020 1089.380 ;
        RECT 2524.020 1089.370 2527.020 1089.380 ;
        RECT 2704.020 1089.370 2707.020 1089.380 ;
        RECT 2884.020 1089.370 2887.020 1089.380 ;
        RECT 2926.600 1089.370 2929.600 1089.380 ;
        RECT -38.180 966.380 -35.180 966.390 ;
        RECT 58.020 966.380 61.020 966.390 ;
        RECT 238.020 966.380 241.020 966.390 ;
        RECT 418.020 966.380 421.020 966.390 ;
        RECT 598.020 966.380 601.020 966.390 ;
        RECT 778.020 966.380 781.020 966.390 ;
        RECT 958.020 966.380 961.020 966.390 ;
        RECT 1138.020 966.380 1141.020 966.390 ;
        RECT 1318.020 966.380 1321.020 966.390 ;
        RECT 1498.020 966.380 1501.020 966.390 ;
        RECT 1678.020 966.380 1681.020 966.390 ;
        RECT 1858.020 966.380 1861.020 966.390 ;
        RECT 2038.020 966.380 2041.020 966.390 ;
        RECT 2218.020 966.380 2221.020 966.390 ;
        RECT 2398.020 966.380 2401.020 966.390 ;
        RECT 2578.020 966.380 2581.020 966.390 ;
        RECT 2758.020 966.380 2761.020 966.390 ;
        RECT 2954.800 966.380 2957.800 966.390 ;
        RECT -42.880 963.380 2962.500 966.380 ;
        RECT -38.180 963.370 -35.180 963.380 ;
        RECT 58.020 963.370 61.020 963.380 ;
        RECT 238.020 963.370 241.020 963.380 ;
        RECT 418.020 963.370 421.020 963.380 ;
        RECT 598.020 963.370 601.020 963.380 ;
        RECT 778.020 963.370 781.020 963.380 ;
        RECT 958.020 963.370 961.020 963.380 ;
        RECT 1138.020 963.370 1141.020 963.380 ;
        RECT 1318.020 963.370 1321.020 963.380 ;
        RECT 1498.020 963.370 1501.020 963.380 ;
        RECT 1678.020 963.370 1681.020 963.380 ;
        RECT 1858.020 963.370 1861.020 963.380 ;
        RECT 2038.020 963.370 2041.020 963.380 ;
        RECT 2218.020 963.370 2221.020 963.380 ;
        RECT 2398.020 963.370 2401.020 963.380 ;
        RECT 2578.020 963.370 2581.020 963.380 ;
        RECT 2758.020 963.370 2761.020 963.380 ;
        RECT 2954.800 963.370 2957.800 963.380 ;
        RECT -28.780 948.380 -25.780 948.390 ;
        RECT 40.020 948.380 43.020 948.390 ;
        RECT 220.020 948.380 223.020 948.390 ;
        RECT 400.020 948.380 403.020 948.390 ;
        RECT 580.020 948.380 583.020 948.390 ;
        RECT 760.020 948.380 763.020 948.390 ;
        RECT 940.020 948.380 943.020 948.390 ;
        RECT 1120.020 948.380 1123.020 948.390 ;
        RECT 1300.020 948.380 1303.020 948.390 ;
        RECT 1480.020 948.380 1483.020 948.390 ;
        RECT 1660.020 948.380 1663.020 948.390 ;
        RECT 1840.020 948.380 1843.020 948.390 ;
        RECT 2020.020 948.380 2023.020 948.390 ;
        RECT 2200.020 948.380 2203.020 948.390 ;
        RECT 2380.020 948.380 2383.020 948.390 ;
        RECT 2560.020 948.380 2563.020 948.390 ;
        RECT 2740.020 948.380 2743.020 948.390 ;
        RECT 2945.400 948.380 2948.400 948.390 ;
        RECT -33.480 945.380 2953.100 948.380 ;
        RECT -28.780 945.370 -25.780 945.380 ;
        RECT 40.020 945.370 43.020 945.380 ;
        RECT 220.020 945.370 223.020 945.380 ;
        RECT 400.020 945.370 403.020 945.380 ;
        RECT 580.020 945.370 583.020 945.380 ;
        RECT 760.020 945.370 763.020 945.380 ;
        RECT 940.020 945.370 943.020 945.380 ;
        RECT 1120.020 945.370 1123.020 945.380 ;
        RECT 1300.020 945.370 1303.020 945.380 ;
        RECT 1480.020 945.370 1483.020 945.380 ;
        RECT 1660.020 945.370 1663.020 945.380 ;
        RECT 1840.020 945.370 1843.020 945.380 ;
        RECT 2020.020 945.370 2023.020 945.380 ;
        RECT 2200.020 945.370 2203.020 945.380 ;
        RECT 2380.020 945.370 2383.020 945.380 ;
        RECT 2560.020 945.370 2563.020 945.380 ;
        RECT 2740.020 945.370 2743.020 945.380 ;
        RECT 2945.400 945.370 2948.400 945.380 ;
        RECT -19.380 930.380 -16.380 930.390 ;
        RECT 22.020 930.380 25.020 930.390 ;
        RECT 202.020 930.380 205.020 930.390 ;
        RECT 382.020 930.380 385.020 930.390 ;
        RECT 562.020 930.380 565.020 930.390 ;
        RECT 742.020 930.380 745.020 930.390 ;
        RECT 922.020 930.380 925.020 930.390 ;
        RECT 1102.020 930.380 1105.020 930.390 ;
        RECT 1282.020 930.380 1285.020 930.390 ;
        RECT 1462.020 930.380 1465.020 930.390 ;
        RECT 1642.020 930.380 1645.020 930.390 ;
        RECT 1822.020 930.380 1825.020 930.390 ;
        RECT 2002.020 930.380 2005.020 930.390 ;
        RECT 2182.020 930.380 2185.020 930.390 ;
        RECT 2362.020 930.380 2365.020 930.390 ;
        RECT 2542.020 930.380 2545.020 930.390 ;
        RECT 2722.020 930.380 2725.020 930.390 ;
        RECT 2902.020 930.380 2905.020 930.390 ;
        RECT 2936.000 930.380 2939.000 930.390 ;
        RECT -24.080 927.380 2943.700 930.380 ;
        RECT -19.380 927.370 -16.380 927.380 ;
        RECT 22.020 927.370 25.020 927.380 ;
        RECT 202.020 927.370 205.020 927.380 ;
        RECT 382.020 927.370 385.020 927.380 ;
        RECT 562.020 927.370 565.020 927.380 ;
        RECT 742.020 927.370 745.020 927.380 ;
        RECT 922.020 927.370 925.020 927.380 ;
        RECT 1102.020 927.370 1105.020 927.380 ;
        RECT 1282.020 927.370 1285.020 927.380 ;
        RECT 1462.020 927.370 1465.020 927.380 ;
        RECT 1642.020 927.370 1645.020 927.380 ;
        RECT 1822.020 927.370 1825.020 927.380 ;
        RECT 2002.020 927.370 2005.020 927.380 ;
        RECT 2182.020 927.370 2185.020 927.380 ;
        RECT 2362.020 927.370 2365.020 927.380 ;
        RECT 2542.020 927.370 2545.020 927.380 ;
        RECT 2722.020 927.370 2725.020 927.380 ;
        RECT 2902.020 927.370 2905.020 927.380 ;
        RECT 2936.000 927.370 2939.000 927.380 ;
        RECT -9.980 912.380 -6.980 912.390 ;
        RECT 4.020 912.380 7.020 912.390 ;
        RECT 184.020 912.380 187.020 912.390 ;
        RECT 364.020 912.380 367.020 912.390 ;
        RECT 544.020 912.380 547.020 912.390 ;
        RECT 724.020 912.380 727.020 912.390 ;
        RECT 904.020 912.380 907.020 912.390 ;
        RECT 1084.020 912.380 1087.020 912.390 ;
        RECT 1264.020 912.380 1267.020 912.390 ;
        RECT 1444.020 912.380 1447.020 912.390 ;
        RECT 1624.020 912.380 1627.020 912.390 ;
        RECT 1804.020 912.380 1807.020 912.390 ;
        RECT 1984.020 912.380 1987.020 912.390 ;
        RECT 2164.020 912.380 2167.020 912.390 ;
        RECT 2344.020 912.380 2347.020 912.390 ;
        RECT 2524.020 912.380 2527.020 912.390 ;
        RECT 2704.020 912.380 2707.020 912.390 ;
        RECT 2884.020 912.380 2887.020 912.390 ;
        RECT 2926.600 912.380 2929.600 912.390 ;
        RECT -14.680 909.380 2934.300 912.380 ;
        RECT -9.980 909.370 -6.980 909.380 ;
        RECT 4.020 909.370 7.020 909.380 ;
        RECT 184.020 909.370 187.020 909.380 ;
        RECT 364.020 909.370 367.020 909.380 ;
        RECT 544.020 909.370 547.020 909.380 ;
        RECT 724.020 909.370 727.020 909.380 ;
        RECT 904.020 909.370 907.020 909.380 ;
        RECT 1084.020 909.370 1087.020 909.380 ;
        RECT 1264.020 909.370 1267.020 909.380 ;
        RECT 1444.020 909.370 1447.020 909.380 ;
        RECT 1624.020 909.370 1627.020 909.380 ;
        RECT 1804.020 909.370 1807.020 909.380 ;
        RECT 1984.020 909.370 1987.020 909.380 ;
        RECT 2164.020 909.370 2167.020 909.380 ;
        RECT 2344.020 909.370 2347.020 909.380 ;
        RECT 2524.020 909.370 2527.020 909.380 ;
        RECT 2704.020 909.370 2707.020 909.380 ;
        RECT 2884.020 909.370 2887.020 909.380 ;
        RECT 2926.600 909.370 2929.600 909.380 ;
        RECT -38.180 786.380 -35.180 786.390 ;
        RECT 58.020 786.380 61.020 786.390 ;
        RECT 238.020 786.380 241.020 786.390 ;
        RECT 418.020 786.380 421.020 786.390 ;
        RECT 598.020 786.380 601.020 786.390 ;
        RECT 778.020 786.380 781.020 786.390 ;
        RECT 958.020 786.380 961.020 786.390 ;
        RECT 1138.020 786.380 1141.020 786.390 ;
        RECT 1318.020 786.380 1321.020 786.390 ;
        RECT 1498.020 786.380 1501.020 786.390 ;
        RECT 1678.020 786.380 1681.020 786.390 ;
        RECT 1858.020 786.380 1861.020 786.390 ;
        RECT 2038.020 786.380 2041.020 786.390 ;
        RECT 2218.020 786.380 2221.020 786.390 ;
        RECT 2398.020 786.380 2401.020 786.390 ;
        RECT 2578.020 786.380 2581.020 786.390 ;
        RECT 2758.020 786.380 2761.020 786.390 ;
        RECT 2954.800 786.380 2957.800 786.390 ;
        RECT -42.880 783.380 2962.500 786.380 ;
        RECT -38.180 783.370 -35.180 783.380 ;
        RECT 58.020 783.370 61.020 783.380 ;
        RECT 238.020 783.370 241.020 783.380 ;
        RECT 418.020 783.370 421.020 783.380 ;
        RECT 598.020 783.370 601.020 783.380 ;
        RECT 778.020 783.370 781.020 783.380 ;
        RECT 958.020 783.370 961.020 783.380 ;
        RECT 1138.020 783.370 1141.020 783.380 ;
        RECT 1318.020 783.370 1321.020 783.380 ;
        RECT 1498.020 783.370 1501.020 783.380 ;
        RECT 1678.020 783.370 1681.020 783.380 ;
        RECT 1858.020 783.370 1861.020 783.380 ;
        RECT 2038.020 783.370 2041.020 783.380 ;
        RECT 2218.020 783.370 2221.020 783.380 ;
        RECT 2398.020 783.370 2401.020 783.380 ;
        RECT 2578.020 783.370 2581.020 783.380 ;
        RECT 2758.020 783.370 2761.020 783.380 ;
        RECT 2954.800 783.370 2957.800 783.380 ;
        RECT -28.780 768.380 -25.780 768.390 ;
        RECT 40.020 768.380 43.020 768.390 ;
        RECT 220.020 768.380 223.020 768.390 ;
        RECT 400.020 768.380 403.020 768.390 ;
        RECT 580.020 768.380 583.020 768.390 ;
        RECT 760.020 768.380 763.020 768.390 ;
        RECT 940.020 768.380 943.020 768.390 ;
        RECT 1120.020 768.380 1123.020 768.390 ;
        RECT 1300.020 768.380 1303.020 768.390 ;
        RECT 1480.020 768.380 1483.020 768.390 ;
        RECT 1660.020 768.380 1663.020 768.390 ;
        RECT 1840.020 768.380 1843.020 768.390 ;
        RECT 2020.020 768.380 2023.020 768.390 ;
        RECT 2200.020 768.380 2203.020 768.390 ;
        RECT 2380.020 768.380 2383.020 768.390 ;
        RECT 2560.020 768.380 2563.020 768.390 ;
        RECT 2740.020 768.380 2743.020 768.390 ;
        RECT 2945.400 768.380 2948.400 768.390 ;
        RECT -33.480 765.380 2953.100 768.380 ;
        RECT -28.780 765.370 -25.780 765.380 ;
        RECT 40.020 765.370 43.020 765.380 ;
        RECT 220.020 765.370 223.020 765.380 ;
        RECT 400.020 765.370 403.020 765.380 ;
        RECT 580.020 765.370 583.020 765.380 ;
        RECT 760.020 765.370 763.020 765.380 ;
        RECT 940.020 765.370 943.020 765.380 ;
        RECT 1120.020 765.370 1123.020 765.380 ;
        RECT 1300.020 765.370 1303.020 765.380 ;
        RECT 1480.020 765.370 1483.020 765.380 ;
        RECT 1660.020 765.370 1663.020 765.380 ;
        RECT 1840.020 765.370 1843.020 765.380 ;
        RECT 2020.020 765.370 2023.020 765.380 ;
        RECT 2200.020 765.370 2203.020 765.380 ;
        RECT 2380.020 765.370 2383.020 765.380 ;
        RECT 2560.020 765.370 2563.020 765.380 ;
        RECT 2740.020 765.370 2743.020 765.380 ;
        RECT 2945.400 765.370 2948.400 765.380 ;
        RECT -19.380 750.380 -16.380 750.390 ;
        RECT 22.020 750.380 25.020 750.390 ;
        RECT 202.020 750.380 205.020 750.390 ;
        RECT 382.020 750.380 385.020 750.390 ;
        RECT 562.020 750.380 565.020 750.390 ;
        RECT 742.020 750.380 745.020 750.390 ;
        RECT 922.020 750.380 925.020 750.390 ;
        RECT 1102.020 750.380 1105.020 750.390 ;
        RECT 1282.020 750.380 1285.020 750.390 ;
        RECT 1462.020 750.380 1465.020 750.390 ;
        RECT 1642.020 750.380 1645.020 750.390 ;
        RECT 1822.020 750.380 1825.020 750.390 ;
        RECT 2002.020 750.380 2005.020 750.390 ;
        RECT 2182.020 750.380 2185.020 750.390 ;
        RECT 2362.020 750.380 2365.020 750.390 ;
        RECT 2542.020 750.380 2545.020 750.390 ;
        RECT 2722.020 750.380 2725.020 750.390 ;
        RECT 2902.020 750.380 2905.020 750.390 ;
        RECT 2936.000 750.380 2939.000 750.390 ;
        RECT -24.080 747.380 2943.700 750.380 ;
        RECT -19.380 747.370 -16.380 747.380 ;
        RECT 22.020 747.370 25.020 747.380 ;
        RECT 202.020 747.370 205.020 747.380 ;
        RECT 382.020 747.370 385.020 747.380 ;
        RECT 562.020 747.370 565.020 747.380 ;
        RECT 742.020 747.370 745.020 747.380 ;
        RECT 922.020 747.370 925.020 747.380 ;
        RECT 1102.020 747.370 1105.020 747.380 ;
        RECT 1282.020 747.370 1285.020 747.380 ;
        RECT 1462.020 747.370 1465.020 747.380 ;
        RECT 1642.020 747.370 1645.020 747.380 ;
        RECT 1822.020 747.370 1825.020 747.380 ;
        RECT 2002.020 747.370 2005.020 747.380 ;
        RECT 2182.020 747.370 2185.020 747.380 ;
        RECT 2362.020 747.370 2365.020 747.380 ;
        RECT 2542.020 747.370 2545.020 747.380 ;
        RECT 2722.020 747.370 2725.020 747.380 ;
        RECT 2902.020 747.370 2905.020 747.380 ;
        RECT 2936.000 747.370 2939.000 747.380 ;
        RECT -9.980 732.380 -6.980 732.390 ;
        RECT 4.020 732.380 7.020 732.390 ;
        RECT 184.020 732.380 187.020 732.390 ;
        RECT 364.020 732.380 367.020 732.390 ;
        RECT 544.020 732.380 547.020 732.390 ;
        RECT 724.020 732.380 727.020 732.390 ;
        RECT 904.020 732.380 907.020 732.390 ;
        RECT 1084.020 732.380 1087.020 732.390 ;
        RECT 1264.020 732.380 1267.020 732.390 ;
        RECT 1444.020 732.380 1447.020 732.390 ;
        RECT 1624.020 732.380 1627.020 732.390 ;
        RECT 1804.020 732.380 1807.020 732.390 ;
        RECT 1984.020 732.380 1987.020 732.390 ;
        RECT 2164.020 732.380 2167.020 732.390 ;
        RECT 2344.020 732.380 2347.020 732.390 ;
        RECT 2524.020 732.380 2527.020 732.390 ;
        RECT 2704.020 732.380 2707.020 732.390 ;
        RECT 2884.020 732.380 2887.020 732.390 ;
        RECT 2926.600 732.380 2929.600 732.390 ;
        RECT -14.680 729.380 2934.300 732.380 ;
        RECT -9.980 729.370 -6.980 729.380 ;
        RECT 4.020 729.370 7.020 729.380 ;
        RECT 184.020 729.370 187.020 729.380 ;
        RECT 364.020 729.370 367.020 729.380 ;
        RECT 544.020 729.370 547.020 729.380 ;
        RECT 724.020 729.370 727.020 729.380 ;
        RECT 904.020 729.370 907.020 729.380 ;
        RECT 1084.020 729.370 1087.020 729.380 ;
        RECT 1264.020 729.370 1267.020 729.380 ;
        RECT 1444.020 729.370 1447.020 729.380 ;
        RECT 1624.020 729.370 1627.020 729.380 ;
        RECT 1804.020 729.370 1807.020 729.380 ;
        RECT 1984.020 729.370 1987.020 729.380 ;
        RECT 2164.020 729.370 2167.020 729.380 ;
        RECT 2344.020 729.370 2347.020 729.380 ;
        RECT 2524.020 729.370 2527.020 729.380 ;
        RECT 2704.020 729.370 2707.020 729.380 ;
        RECT 2884.020 729.370 2887.020 729.380 ;
        RECT 2926.600 729.370 2929.600 729.380 ;
        RECT -38.180 606.380 -35.180 606.390 ;
        RECT 58.020 606.380 61.020 606.390 ;
        RECT 238.020 606.380 241.020 606.390 ;
        RECT 418.020 606.380 421.020 606.390 ;
        RECT 598.020 606.380 601.020 606.390 ;
        RECT 778.020 606.380 781.020 606.390 ;
        RECT 958.020 606.380 961.020 606.390 ;
        RECT 1138.020 606.380 1141.020 606.390 ;
        RECT 1318.020 606.380 1321.020 606.390 ;
        RECT 1498.020 606.380 1501.020 606.390 ;
        RECT 1678.020 606.380 1681.020 606.390 ;
        RECT 1858.020 606.380 1861.020 606.390 ;
        RECT 2038.020 606.380 2041.020 606.390 ;
        RECT 2218.020 606.380 2221.020 606.390 ;
        RECT 2398.020 606.380 2401.020 606.390 ;
        RECT 2578.020 606.380 2581.020 606.390 ;
        RECT 2758.020 606.380 2761.020 606.390 ;
        RECT 2954.800 606.380 2957.800 606.390 ;
        RECT -42.880 603.380 2962.500 606.380 ;
        RECT -38.180 603.370 -35.180 603.380 ;
        RECT 58.020 603.370 61.020 603.380 ;
        RECT 238.020 603.370 241.020 603.380 ;
        RECT 418.020 603.370 421.020 603.380 ;
        RECT 598.020 603.370 601.020 603.380 ;
        RECT 778.020 603.370 781.020 603.380 ;
        RECT 958.020 603.370 961.020 603.380 ;
        RECT 1138.020 603.370 1141.020 603.380 ;
        RECT 1318.020 603.370 1321.020 603.380 ;
        RECT 1498.020 603.370 1501.020 603.380 ;
        RECT 1678.020 603.370 1681.020 603.380 ;
        RECT 1858.020 603.370 1861.020 603.380 ;
        RECT 2038.020 603.370 2041.020 603.380 ;
        RECT 2218.020 603.370 2221.020 603.380 ;
        RECT 2398.020 603.370 2401.020 603.380 ;
        RECT 2578.020 603.370 2581.020 603.380 ;
        RECT 2758.020 603.370 2761.020 603.380 ;
        RECT 2954.800 603.370 2957.800 603.380 ;
        RECT -28.780 588.380 -25.780 588.390 ;
        RECT 40.020 588.380 43.020 588.390 ;
        RECT 220.020 588.380 223.020 588.390 ;
        RECT 400.020 588.380 403.020 588.390 ;
        RECT 580.020 588.380 583.020 588.390 ;
        RECT 760.020 588.380 763.020 588.390 ;
        RECT 940.020 588.380 943.020 588.390 ;
        RECT 1120.020 588.380 1123.020 588.390 ;
        RECT 1300.020 588.380 1303.020 588.390 ;
        RECT 1480.020 588.380 1483.020 588.390 ;
        RECT 1660.020 588.380 1663.020 588.390 ;
        RECT 1840.020 588.380 1843.020 588.390 ;
        RECT 2020.020 588.380 2023.020 588.390 ;
        RECT 2200.020 588.380 2203.020 588.390 ;
        RECT 2380.020 588.380 2383.020 588.390 ;
        RECT 2560.020 588.380 2563.020 588.390 ;
        RECT 2740.020 588.380 2743.020 588.390 ;
        RECT 2945.400 588.380 2948.400 588.390 ;
        RECT -33.480 585.380 2953.100 588.380 ;
        RECT -28.780 585.370 -25.780 585.380 ;
        RECT 40.020 585.370 43.020 585.380 ;
        RECT 220.020 585.370 223.020 585.380 ;
        RECT 400.020 585.370 403.020 585.380 ;
        RECT 580.020 585.370 583.020 585.380 ;
        RECT 760.020 585.370 763.020 585.380 ;
        RECT 940.020 585.370 943.020 585.380 ;
        RECT 1120.020 585.370 1123.020 585.380 ;
        RECT 1300.020 585.370 1303.020 585.380 ;
        RECT 1480.020 585.370 1483.020 585.380 ;
        RECT 1660.020 585.370 1663.020 585.380 ;
        RECT 1840.020 585.370 1843.020 585.380 ;
        RECT 2020.020 585.370 2023.020 585.380 ;
        RECT 2200.020 585.370 2203.020 585.380 ;
        RECT 2380.020 585.370 2383.020 585.380 ;
        RECT 2560.020 585.370 2563.020 585.380 ;
        RECT 2740.020 585.370 2743.020 585.380 ;
        RECT 2945.400 585.370 2948.400 585.380 ;
        RECT -19.380 570.380 -16.380 570.390 ;
        RECT 22.020 570.380 25.020 570.390 ;
        RECT 202.020 570.380 205.020 570.390 ;
        RECT 382.020 570.380 385.020 570.390 ;
        RECT 562.020 570.380 565.020 570.390 ;
        RECT 742.020 570.380 745.020 570.390 ;
        RECT 922.020 570.380 925.020 570.390 ;
        RECT 1102.020 570.380 1105.020 570.390 ;
        RECT 1282.020 570.380 1285.020 570.390 ;
        RECT 1462.020 570.380 1465.020 570.390 ;
        RECT 1642.020 570.380 1645.020 570.390 ;
        RECT 1822.020 570.380 1825.020 570.390 ;
        RECT 2002.020 570.380 2005.020 570.390 ;
        RECT 2182.020 570.380 2185.020 570.390 ;
        RECT 2362.020 570.380 2365.020 570.390 ;
        RECT 2542.020 570.380 2545.020 570.390 ;
        RECT 2722.020 570.380 2725.020 570.390 ;
        RECT 2902.020 570.380 2905.020 570.390 ;
        RECT 2936.000 570.380 2939.000 570.390 ;
        RECT -24.080 567.380 2943.700 570.380 ;
        RECT -19.380 567.370 -16.380 567.380 ;
        RECT 22.020 567.370 25.020 567.380 ;
        RECT 202.020 567.370 205.020 567.380 ;
        RECT 382.020 567.370 385.020 567.380 ;
        RECT 562.020 567.370 565.020 567.380 ;
        RECT 742.020 567.370 745.020 567.380 ;
        RECT 922.020 567.370 925.020 567.380 ;
        RECT 1102.020 567.370 1105.020 567.380 ;
        RECT 1282.020 567.370 1285.020 567.380 ;
        RECT 1462.020 567.370 1465.020 567.380 ;
        RECT 1642.020 567.370 1645.020 567.380 ;
        RECT 1822.020 567.370 1825.020 567.380 ;
        RECT 2002.020 567.370 2005.020 567.380 ;
        RECT 2182.020 567.370 2185.020 567.380 ;
        RECT 2362.020 567.370 2365.020 567.380 ;
        RECT 2542.020 567.370 2545.020 567.380 ;
        RECT 2722.020 567.370 2725.020 567.380 ;
        RECT 2902.020 567.370 2905.020 567.380 ;
        RECT 2936.000 567.370 2939.000 567.380 ;
        RECT -9.980 552.380 -6.980 552.390 ;
        RECT 4.020 552.380 7.020 552.390 ;
        RECT 184.020 552.380 187.020 552.390 ;
        RECT 364.020 552.380 367.020 552.390 ;
        RECT 544.020 552.380 547.020 552.390 ;
        RECT 724.020 552.380 727.020 552.390 ;
        RECT 904.020 552.380 907.020 552.390 ;
        RECT 1084.020 552.380 1087.020 552.390 ;
        RECT 1264.020 552.380 1267.020 552.390 ;
        RECT 1444.020 552.380 1447.020 552.390 ;
        RECT 1624.020 552.380 1627.020 552.390 ;
        RECT 1804.020 552.380 1807.020 552.390 ;
        RECT 1984.020 552.380 1987.020 552.390 ;
        RECT 2164.020 552.380 2167.020 552.390 ;
        RECT 2344.020 552.380 2347.020 552.390 ;
        RECT 2524.020 552.380 2527.020 552.390 ;
        RECT 2704.020 552.380 2707.020 552.390 ;
        RECT 2884.020 552.380 2887.020 552.390 ;
        RECT 2926.600 552.380 2929.600 552.390 ;
        RECT -14.680 549.380 2934.300 552.380 ;
        RECT -9.980 549.370 -6.980 549.380 ;
        RECT 4.020 549.370 7.020 549.380 ;
        RECT 184.020 549.370 187.020 549.380 ;
        RECT 364.020 549.370 367.020 549.380 ;
        RECT 544.020 549.370 547.020 549.380 ;
        RECT 724.020 549.370 727.020 549.380 ;
        RECT 904.020 549.370 907.020 549.380 ;
        RECT 1084.020 549.370 1087.020 549.380 ;
        RECT 1264.020 549.370 1267.020 549.380 ;
        RECT 1444.020 549.370 1447.020 549.380 ;
        RECT 1624.020 549.370 1627.020 549.380 ;
        RECT 1804.020 549.370 1807.020 549.380 ;
        RECT 1984.020 549.370 1987.020 549.380 ;
        RECT 2164.020 549.370 2167.020 549.380 ;
        RECT 2344.020 549.370 2347.020 549.380 ;
        RECT 2524.020 549.370 2527.020 549.380 ;
        RECT 2704.020 549.370 2707.020 549.380 ;
        RECT 2884.020 549.370 2887.020 549.380 ;
        RECT 2926.600 549.370 2929.600 549.380 ;
        RECT -38.180 426.380 -35.180 426.390 ;
        RECT 58.020 426.380 61.020 426.390 ;
        RECT 238.020 426.380 241.020 426.390 ;
        RECT 418.020 426.380 421.020 426.390 ;
        RECT 598.020 426.380 601.020 426.390 ;
        RECT 778.020 426.380 781.020 426.390 ;
        RECT 958.020 426.380 961.020 426.390 ;
        RECT 1138.020 426.380 1141.020 426.390 ;
        RECT 1318.020 426.380 1321.020 426.390 ;
        RECT 1498.020 426.380 1501.020 426.390 ;
        RECT 1678.020 426.380 1681.020 426.390 ;
        RECT 1858.020 426.380 1861.020 426.390 ;
        RECT 2038.020 426.380 2041.020 426.390 ;
        RECT 2218.020 426.380 2221.020 426.390 ;
        RECT 2398.020 426.380 2401.020 426.390 ;
        RECT 2578.020 426.380 2581.020 426.390 ;
        RECT 2758.020 426.380 2761.020 426.390 ;
        RECT 2954.800 426.380 2957.800 426.390 ;
        RECT -42.880 423.380 2962.500 426.380 ;
        RECT -38.180 423.370 -35.180 423.380 ;
        RECT 58.020 423.370 61.020 423.380 ;
        RECT 238.020 423.370 241.020 423.380 ;
        RECT 418.020 423.370 421.020 423.380 ;
        RECT 598.020 423.370 601.020 423.380 ;
        RECT 778.020 423.370 781.020 423.380 ;
        RECT 958.020 423.370 961.020 423.380 ;
        RECT 1138.020 423.370 1141.020 423.380 ;
        RECT 1318.020 423.370 1321.020 423.380 ;
        RECT 1498.020 423.370 1501.020 423.380 ;
        RECT 1678.020 423.370 1681.020 423.380 ;
        RECT 1858.020 423.370 1861.020 423.380 ;
        RECT 2038.020 423.370 2041.020 423.380 ;
        RECT 2218.020 423.370 2221.020 423.380 ;
        RECT 2398.020 423.370 2401.020 423.380 ;
        RECT 2578.020 423.370 2581.020 423.380 ;
        RECT 2758.020 423.370 2761.020 423.380 ;
        RECT 2954.800 423.370 2957.800 423.380 ;
        RECT -28.780 408.380 -25.780 408.390 ;
        RECT 40.020 408.380 43.020 408.390 ;
        RECT 220.020 408.380 223.020 408.390 ;
        RECT 400.020 408.380 403.020 408.390 ;
        RECT 580.020 408.380 583.020 408.390 ;
        RECT 760.020 408.380 763.020 408.390 ;
        RECT 940.020 408.380 943.020 408.390 ;
        RECT 1120.020 408.380 1123.020 408.390 ;
        RECT 1300.020 408.380 1303.020 408.390 ;
        RECT 1480.020 408.380 1483.020 408.390 ;
        RECT 1660.020 408.380 1663.020 408.390 ;
        RECT 1840.020 408.380 1843.020 408.390 ;
        RECT 2020.020 408.380 2023.020 408.390 ;
        RECT 2200.020 408.380 2203.020 408.390 ;
        RECT 2380.020 408.380 2383.020 408.390 ;
        RECT 2560.020 408.380 2563.020 408.390 ;
        RECT 2740.020 408.380 2743.020 408.390 ;
        RECT 2945.400 408.380 2948.400 408.390 ;
        RECT -33.480 405.380 2953.100 408.380 ;
        RECT -28.780 405.370 -25.780 405.380 ;
        RECT 40.020 405.370 43.020 405.380 ;
        RECT 220.020 405.370 223.020 405.380 ;
        RECT 400.020 405.370 403.020 405.380 ;
        RECT 580.020 405.370 583.020 405.380 ;
        RECT 760.020 405.370 763.020 405.380 ;
        RECT 940.020 405.370 943.020 405.380 ;
        RECT 1120.020 405.370 1123.020 405.380 ;
        RECT 1300.020 405.370 1303.020 405.380 ;
        RECT 1480.020 405.370 1483.020 405.380 ;
        RECT 1660.020 405.370 1663.020 405.380 ;
        RECT 1840.020 405.370 1843.020 405.380 ;
        RECT 2020.020 405.370 2023.020 405.380 ;
        RECT 2200.020 405.370 2203.020 405.380 ;
        RECT 2380.020 405.370 2383.020 405.380 ;
        RECT 2560.020 405.370 2563.020 405.380 ;
        RECT 2740.020 405.370 2743.020 405.380 ;
        RECT 2945.400 405.370 2948.400 405.380 ;
        RECT -19.380 390.380 -16.380 390.390 ;
        RECT 22.020 390.380 25.020 390.390 ;
        RECT 202.020 390.380 205.020 390.390 ;
        RECT 382.020 390.380 385.020 390.390 ;
        RECT 562.020 390.380 565.020 390.390 ;
        RECT 742.020 390.380 745.020 390.390 ;
        RECT 922.020 390.380 925.020 390.390 ;
        RECT 1102.020 390.380 1105.020 390.390 ;
        RECT 1282.020 390.380 1285.020 390.390 ;
        RECT 1462.020 390.380 1465.020 390.390 ;
        RECT 1642.020 390.380 1645.020 390.390 ;
        RECT 1822.020 390.380 1825.020 390.390 ;
        RECT 2002.020 390.380 2005.020 390.390 ;
        RECT 2182.020 390.380 2185.020 390.390 ;
        RECT 2362.020 390.380 2365.020 390.390 ;
        RECT 2542.020 390.380 2545.020 390.390 ;
        RECT 2722.020 390.380 2725.020 390.390 ;
        RECT 2902.020 390.380 2905.020 390.390 ;
        RECT 2936.000 390.380 2939.000 390.390 ;
        RECT -24.080 387.380 2943.700 390.380 ;
        RECT -19.380 387.370 -16.380 387.380 ;
        RECT 22.020 387.370 25.020 387.380 ;
        RECT 202.020 387.370 205.020 387.380 ;
        RECT 382.020 387.370 385.020 387.380 ;
        RECT 562.020 387.370 565.020 387.380 ;
        RECT 742.020 387.370 745.020 387.380 ;
        RECT 922.020 387.370 925.020 387.380 ;
        RECT 1102.020 387.370 1105.020 387.380 ;
        RECT 1282.020 387.370 1285.020 387.380 ;
        RECT 1462.020 387.370 1465.020 387.380 ;
        RECT 1642.020 387.370 1645.020 387.380 ;
        RECT 1822.020 387.370 1825.020 387.380 ;
        RECT 2002.020 387.370 2005.020 387.380 ;
        RECT 2182.020 387.370 2185.020 387.380 ;
        RECT 2362.020 387.370 2365.020 387.380 ;
        RECT 2542.020 387.370 2545.020 387.380 ;
        RECT 2722.020 387.370 2725.020 387.380 ;
        RECT 2902.020 387.370 2905.020 387.380 ;
        RECT 2936.000 387.370 2939.000 387.380 ;
        RECT -9.980 372.380 -6.980 372.390 ;
        RECT 4.020 372.380 7.020 372.390 ;
        RECT 184.020 372.380 187.020 372.390 ;
        RECT 364.020 372.380 367.020 372.390 ;
        RECT 544.020 372.380 547.020 372.390 ;
        RECT 724.020 372.380 727.020 372.390 ;
        RECT 904.020 372.380 907.020 372.390 ;
        RECT 1084.020 372.380 1087.020 372.390 ;
        RECT 1264.020 372.380 1267.020 372.390 ;
        RECT 1444.020 372.380 1447.020 372.390 ;
        RECT 1624.020 372.380 1627.020 372.390 ;
        RECT 1804.020 372.380 1807.020 372.390 ;
        RECT 1984.020 372.380 1987.020 372.390 ;
        RECT 2164.020 372.380 2167.020 372.390 ;
        RECT 2344.020 372.380 2347.020 372.390 ;
        RECT 2524.020 372.380 2527.020 372.390 ;
        RECT 2704.020 372.380 2707.020 372.390 ;
        RECT 2884.020 372.380 2887.020 372.390 ;
        RECT 2926.600 372.380 2929.600 372.390 ;
        RECT -14.680 369.380 2934.300 372.380 ;
        RECT -9.980 369.370 -6.980 369.380 ;
        RECT 4.020 369.370 7.020 369.380 ;
        RECT 184.020 369.370 187.020 369.380 ;
        RECT 364.020 369.370 367.020 369.380 ;
        RECT 544.020 369.370 547.020 369.380 ;
        RECT 724.020 369.370 727.020 369.380 ;
        RECT 904.020 369.370 907.020 369.380 ;
        RECT 1084.020 369.370 1087.020 369.380 ;
        RECT 1264.020 369.370 1267.020 369.380 ;
        RECT 1444.020 369.370 1447.020 369.380 ;
        RECT 1624.020 369.370 1627.020 369.380 ;
        RECT 1804.020 369.370 1807.020 369.380 ;
        RECT 1984.020 369.370 1987.020 369.380 ;
        RECT 2164.020 369.370 2167.020 369.380 ;
        RECT 2344.020 369.370 2347.020 369.380 ;
        RECT 2524.020 369.370 2527.020 369.380 ;
        RECT 2704.020 369.370 2707.020 369.380 ;
        RECT 2884.020 369.370 2887.020 369.380 ;
        RECT 2926.600 369.370 2929.600 369.380 ;
        RECT -38.180 246.380 -35.180 246.390 ;
        RECT 58.020 246.380 61.020 246.390 ;
        RECT 238.020 246.380 241.020 246.390 ;
        RECT 418.020 246.380 421.020 246.390 ;
        RECT 598.020 246.380 601.020 246.390 ;
        RECT 778.020 246.380 781.020 246.390 ;
        RECT 958.020 246.380 961.020 246.390 ;
        RECT 1138.020 246.380 1141.020 246.390 ;
        RECT 1318.020 246.380 1321.020 246.390 ;
        RECT 1498.020 246.380 1501.020 246.390 ;
        RECT 1678.020 246.380 1681.020 246.390 ;
        RECT 1858.020 246.380 1861.020 246.390 ;
        RECT 2038.020 246.380 2041.020 246.390 ;
        RECT 2218.020 246.380 2221.020 246.390 ;
        RECT 2398.020 246.380 2401.020 246.390 ;
        RECT 2578.020 246.380 2581.020 246.390 ;
        RECT 2758.020 246.380 2761.020 246.390 ;
        RECT 2954.800 246.380 2957.800 246.390 ;
        RECT -42.880 243.380 2962.500 246.380 ;
        RECT -38.180 243.370 -35.180 243.380 ;
        RECT 58.020 243.370 61.020 243.380 ;
        RECT 238.020 243.370 241.020 243.380 ;
        RECT 418.020 243.370 421.020 243.380 ;
        RECT 598.020 243.370 601.020 243.380 ;
        RECT 778.020 243.370 781.020 243.380 ;
        RECT 958.020 243.370 961.020 243.380 ;
        RECT 1138.020 243.370 1141.020 243.380 ;
        RECT 1318.020 243.370 1321.020 243.380 ;
        RECT 1498.020 243.370 1501.020 243.380 ;
        RECT 1678.020 243.370 1681.020 243.380 ;
        RECT 1858.020 243.370 1861.020 243.380 ;
        RECT 2038.020 243.370 2041.020 243.380 ;
        RECT 2218.020 243.370 2221.020 243.380 ;
        RECT 2398.020 243.370 2401.020 243.380 ;
        RECT 2578.020 243.370 2581.020 243.380 ;
        RECT 2758.020 243.370 2761.020 243.380 ;
        RECT 2954.800 243.370 2957.800 243.380 ;
        RECT -28.780 228.380 -25.780 228.390 ;
        RECT 40.020 228.380 43.020 228.390 ;
        RECT 220.020 228.380 223.020 228.390 ;
        RECT 400.020 228.380 403.020 228.390 ;
        RECT 580.020 228.380 583.020 228.390 ;
        RECT 760.020 228.380 763.020 228.390 ;
        RECT 940.020 228.380 943.020 228.390 ;
        RECT 1120.020 228.380 1123.020 228.390 ;
        RECT 1300.020 228.380 1303.020 228.390 ;
        RECT 1480.020 228.380 1483.020 228.390 ;
        RECT 1660.020 228.380 1663.020 228.390 ;
        RECT 1840.020 228.380 1843.020 228.390 ;
        RECT 2020.020 228.380 2023.020 228.390 ;
        RECT 2200.020 228.380 2203.020 228.390 ;
        RECT 2380.020 228.380 2383.020 228.390 ;
        RECT 2560.020 228.380 2563.020 228.390 ;
        RECT 2740.020 228.380 2743.020 228.390 ;
        RECT 2945.400 228.380 2948.400 228.390 ;
        RECT -33.480 225.380 2953.100 228.380 ;
        RECT -28.780 225.370 -25.780 225.380 ;
        RECT 40.020 225.370 43.020 225.380 ;
        RECT 220.020 225.370 223.020 225.380 ;
        RECT 400.020 225.370 403.020 225.380 ;
        RECT 580.020 225.370 583.020 225.380 ;
        RECT 760.020 225.370 763.020 225.380 ;
        RECT 940.020 225.370 943.020 225.380 ;
        RECT 1120.020 225.370 1123.020 225.380 ;
        RECT 1300.020 225.370 1303.020 225.380 ;
        RECT 1480.020 225.370 1483.020 225.380 ;
        RECT 1660.020 225.370 1663.020 225.380 ;
        RECT 1840.020 225.370 1843.020 225.380 ;
        RECT 2020.020 225.370 2023.020 225.380 ;
        RECT 2200.020 225.370 2203.020 225.380 ;
        RECT 2380.020 225.370 2383.020 225.380 ;
        RECT 2560.020 225.370 2563.020 225.380 ;
        RECT 2740.020 225.370 2743.020 225.380 ;
        RECT 2945.400 225.370 2948.400 225.380 ;
        RECT -19.380 210.380 -16.380 210.390 ;
        RECT 22.020 210.380 25.020 210.390 ;
        RECT 202.020 210.380 205.020 210.390 ;
        RECT 382.020 210.380 385.020 210.390 ;
        RECT 562.020 210.380 565.020 210.390 ;
        RECT 742.020 210.380 745.020 210.390 ;
        RECT 922.020 210.380 925.020 210.390 ;
        RECT 1102.020 210.380 1105.020 210.390 ;
        RECT 1282.020 210.380 1285.020 210.390 ;
        RECT 1462.020 210.380 1465.020 210.390 ;
        RECT 1642.020 210.380 1645.020 210.390 ;
        RECT 1822.020 210.380 1825.020 210.390 ;
        RECT 2002.020 210.380 2005.020 210.390 ;
        RECT 2182.020 210.380 2185.020 210.390 ;
        RECT 2362.020 210.380 2365.020 210.390 ;
        RECT 2542.020 210.380 2545.020 210.390 ;
        RECT 2722.020 210.380 2725.020 210.390 ;
        RECT 2902.020 210.380 2905.020 210.390 ;
        RECT 2936.000 210.380 2939.000 210.390 ;
        RECT -24.080 207.380 2943.700 210.380 ;
        RECT -19.380 207.370 -16.380 207.380 ;
        RECT 22.020 207.370 25.020 207.380 ;
        RECT 202.020 207.370 205.020 207.380 ;
        RECT 382.020 207.370 385.020 207.380 ;
        RECT 562.020 207.370 565.020 207.380 ;
        RECT 742.020 207.370 745.020 207.380 ;
        RECT 922.020 207.370 925.020 207.380 ;
        RECT 1102.020 207.370 1105.020 207.380 ;
        RECT 1282.020 207.370 1285.020 207.380 ;
        RECT 1462.020 207.370 1465.020 207.380 ;
        RECT 1642.020 207.370 1645.020 207.380 ;
        RECT 1822.020 207.370 1825.020 207.380 ;
        RECT 2002.020 207.370 2005.020 207.380 ;
        RECT 2182.020 207.370 2185.020 207.380 ;
        RECT 2362.020 207.370 2365.020 207.380 ;
        RECT 2542.020 207.370 2545.020 207.380 ;
        RECT 2722.020 207.370 2725.020 207.380 ;
        RECT 2902.020 207.370 2905.020 207.380 ;
        RECT 2936.000 207.370 2939.000 207.380 ;
        RECT -9.980 192.380 -6.980 192.390 ;
        RECT 4.020 192.380 7.020 192.390 ;
        RECT 184.020 192.380 187.020 192.390 ;
        RECT 364.020 192.380 367.020 192.390 ;
        RECT 544.020 192.380 547.020 192.390 ;
        RECT 724.020 192.380 727.020 192.390 ;
        RECT 904.020 192.380 907.020 192.390 ;
        RECT 1084.020 192.380 1087.020 192.390 ;
        RECT 1264.020 192.380 1267.020 192.390 ;
        RECT 1444.020 192.380 1447.020 192.390 ;
        RECT 1624.020 192.380 1627.020 192.390 ;
        RECT 1804.020 192.380 1807.020 192.390 ;
        RECT 1984.020 192.380 1987.020 192.390 ;
        RECT 2164.020 192.380 2167.020 192.390 ;
        RECT 2344.020 192.380 2347.020 192.390 ;
        RECT 2524.020 192.380 2527.020 192.390 ;
        RECT 2704.020 192.380 2707.020 192.390 ;
        RECT 2884.020 192.380 2887.020 192.390 ;
        RECT 2926.600 192.380 2929.600 192.390 ;
        RECT -14.680 189.380 2934.300 192.380 ;
        RECT -9.980 189.370 -6.980 189.380 ;
        RECT 4.020 189.370 7.020 189.380 ;
        RECT 184.020 189.370 187.020 189.380 ;
        RECT 364.020 189.370 367.020 189.380 ;
        RECT 544.020 189.370 547.020 189.380 ;
        RECT 724.020 189.370 727.020 189.380 ;
        RECT 904.020 189.370 907.020 189.380 ;
        RECT 1084.020 189.370 1087.020 189.380 ;
        RECT 1264.020 189.370 1267.020 189.380 ;
        RECT 1444.020 189.370 1447.020 189.380 ;
        RECT 1624.020 189.370 1627.020 189.380 ;
        RECT 1804.020 189.370 1807.020 189.380 ;
        RECT 1984.020 189.370 1987.020 189.380 ;
        RECT 2164.020 189.370 2167.020 189.380 ;
        RECT 2344.020 189.370 2347.020 189.380 ;
        RECT 2524.020 189.370 2527.020 189.380 ;
        RECT 2704.020 189.370 2707.020 189.380 ;
        RECT 2884.020 189.370 2887.020 189.380 ;
        RECT 2926.600 189.370 2929.600 189.380 ;
        RECT -38.180 66.380 -35.180 66.390 ;
        RECT 58.020 66.380 61.020 66.390 ;
        RECT 238.020 66.380 241.020 66.390 ;
        RECT 418.020 66.380 421.020 66.390 ;
        RECT 598.020 66.380 601.020 66.390 ;
        RECT 778.020 66.380 781.020 66.390 ;
        RECT 958.020 66.380 961.020 66.390 ;
        RECT 1138.020 66.380 1141.020 66.390 ;
        RECT 1318.020 66.380 1321.020 66.390 ;
        RECT 1498.020 66.380 1501.020 66.390 ;
        RECT 1678.020 66.380 1681.020 66.390 ;
        RECT 1858.020 66.380 1861.020 66.390 ;
        RECT 2038.020 66.380 2041.020 66.390 ;
        RECT 2218.020 66.380 2221.020 66.390 ;
        RECT 2398.020 66.380 2401.020 66.390 ;
        RECT 2578.020 66.380 2581.020 66.390 ;
        RECT 2758.020 66.380 2761.020 66.390 ;
        RECT 2954.800 66.380 2957.800 66.390 ;
        RECT -42.880 63.380 2962.500 66.380 ;
        RECT -38.180 63.370 -35.180 63.380 ;
        RECT 58.020 63.370 61.020 63.380 ;
        RECT 238.020 63.370 241.020 63.380 ;
        RECT 418.020 63.370 421.020 63.380 ;
        RECT 598.020 63.370 601.020 63.380 ;
        RECT 778.020 63.370 781.020 63.380 ;
        RECT 958.020 63.370 961.020 63.380 ;
        RECT 1138.020 63.370 1141.020 63.380 ;
        RECT 1318.020 63.370 1321.020 63.380 ;
        RECT 1498.020 63.370 1501.020 63.380 ;
        RECT 1678.020 63.370 1681.020 63.380 ;
        RECT 1858.020 63.370 1861.020 63.380 ;
        RECT 2038.020 63.370 2041.020 63.380 ;
        RECT 2218.020 63.370 2221.020 63.380 ;
        RECT 2398.020 63.370 2401.020 63.380 ;
        RECT 2578.020 63.370 2581.020 63.380 ;
        RECT 2758.020 63.370 2761.020 63.380 ;
        RECT 2954.800 63.370 2957.800 63.380 ;
        RECT -28.780 48.380 -25.780 48.390 ;
        RECT 40.020 48.380 43.020 48.390 ;
        RECT 220.020 48.380 223.020 48.390 ;
        RECT 400.020 48.380 403.020 48.390 ;
        RECT 580.020 48.380 583.020 48.390 ;
        RECT 760.020 48.380 763.020 48.390 ;
        RECT 940.020 48.380 943.020 48.390 ;
        RECT 1120.020 48.380 1123.020 48.390 ;
        RECT 1300.020 48.380 1303.020 48.390 ;
        RECT 1480.020 48.380 1483.020 48.390 ;
        RECT 1660.020 48.380 1663.020 48.390 ;
        RECT 1840.020 48.380 1843.020 48.390 ;
        RECT 2020.020 48.380 2023.020 48.390 ;
        RECT 2200.020 48.380 2203.020 48.390 ;
        RECT 2380.020 48.380 2383.020 48.390 ;
        RECT 2560.020 48.380 2563.020 48.390 ;
        RECT 2740.020 48.380 2743.020 48.390 ;
        RECT 2945.400 48.380 2948.400 48.390 ;
        RECT -33.480 45.380 2953.100 48.380 ;
        RECT -28.780 45.370 -25.780 45.380 ;
        RECT 40.020 45.370 43.020 45.380 ;
        RECT 220.020 45.370 223.020 45.380 ;
        RECT 400.020 45.370 403.020 45.380 ;
        RECT 580.020 45.370 583.020 45.380 ;
        RECT 760.020 45.370 763.020 45.380 ;
        RECT 940.020 45.370 943.020 45.380 ;
        RECT 1120.020 45.370 1123.020 45.380 ;
        RECT 1300.020 45.370 1303.020 45.380 ;
        RECT 1480.020 45.370 1483.020 45.380 ;
        RECT 1660.020 45.370 1663.020 45.380 ;
        RECT 1840.020 45.370 1843.020 45.380 ;
        RECT 2020.020 45.370 2023.020 45.380 ;
        RECT 2200.020 45.370 2203.020 45.380 ;
        RECT 2380.020 45.370 2383.020 45.380 ;
        RECT 2560.020 45.370 2563.020 45.380 ;
        RECT 2740.020 45.370 2743.020 45.380 ;
        RECT 2945.400 45.370 2948.400 45.380 ;
        RECT -19.380 30.380 -16.380 30.390 ;
        RECT 22.020 30.380 25.020 30.390 ;
        RECT 202.020 30.380 205.020 30.390 ;
        RECT 382.020 30.380 385.020 30.390 ;
        RECT 562.020 30.380 565.020 30.390 ;
        RECT 742.020 30.380 745.020 30.390 ;
        RECT 922.020 30.380 925.020 30.390 ;
        RECT 1102.020 30.380 1105.020 30.390 ;
        RECT 1282.020 30.380 1285.020 30.390 ;
        RECT 1462.020 30.380 1465.020 30.390 ;
        RECT 1642.020 30.380 1645.020 30.390 ;
        RECT 1822.020 30.380 1825.020 30.390 ;
        RECT 2002.020 30.380 2005.020 30.390 ;
        RECT 2182.020 30.380 2185.020 30.390 ;
        RECT 2362.020 30.380 2365.020 30.390 ;
        RECT 2542.020 30.380 2545.020 30.390 ;
        RECT 2722.020 30.380 2725.020 30.390 ;
        RECT 2902.020 30.380 2905.020 30.390 ;
        RECT 2936.000 30.380 2939.000 30.390 ;
        RECT -24.080 27.380 2943.700 30.380 ;
        RECT -19.380 27.370 -16.380 27.380 ;
        RECT 22.020 27.370 25.020 27.380 ;
        RECT 202.020 27.370 205.020 27.380 ;
        RECT 382.020 27.370 385.020 27.380 ;
        RECT 562.020 27.370 565.020 27.380 ;
        RECT 742.020 27.370 745.020 27.380 ;
        RECT 922.020 27.370 925.020 27.380 ;
        RECT 1102.020 27.370 1105.020 27.380 ;
        RECT 1282.020 27.370 1285.020 27.380 ;
        RECT 1462.020 27.370 1465.020 27.380 ;
        RECT 1642.020 27.370 1645.020 27.380 ;
        RECT 1822.020 27.370 1825.020 27.380 ;
        RECT 2002.020 27.370 2005.020 27.380 ;
        RECT 2182.020 27.370 2185.020 27.380 ;
        RECT 2362.020 27.370 2365.020 27.380 ;
        RECT 2542.020 27.370 2545.020 27.380 ;
        RECT 2722.020 27.370 2725.020 27.380 ;
        RECT 2902.020 27.370 2905.020 27.380 ;
        RECT 2936.000 27.370 2939.000 27.380 ;
        RECT -9.980 12.380 -6.980 12.390 ;
        RECT 4.020 12.380 7.020 12.390 ;
        RECT 184.020 12.380 187.020 12.390 ;
        RECT 364.020 12.380 367.020 12.390 ;
        RECT 544.020 12.380 547.020 12.390 ;
        RECT 724.020 12.380 727.020 12.390 ;
        RECT 904.020 12.380 907.020 12.390 ;
        RECT 1084.020 12.380 1087.020 12.390 ;
        RECT 1264.020 12.380 1267.020 12.390 ;
        RECT 1444.020 12.380 1447.020 12.390 ;
        RECT 1624.020 12.380 1627.020 12.390 ;
        RECT 1804.020 12.380 1807.020 12.390 ;
        RECT 1984.020 12.380 1987.020 12.390 ;
        RECT 2164.020 12.380 2167.020 12.390 ;
        RECT 2344.020 12.380 2347.020 12.390 ;
        RECT 2524.020 12.380 2527.020 12.390 ;
        RECT 2704.020 12.380 2707.020 12.390 ;
        RECT 2884.020 12.380 2887.020 12.390 ;
        RECT 2926.600 12.380 2929.600 12.390 ;
        RECT -14.680 9.380 2934.300 12.380 ;
        RECT -9.980 9.370 -6.980 9.380 ;
        RECT 4.020 9.370 7.020 9.380 ;
        RECT 184.020 9.370 187.020 9.380 ;
        RECT 364.020 9.370 367.020 9.380 ;
        RECT 544.020 9.370 547.020 9.380 ;
        RECT 724.020 9.370 727.020 9.380 ;
        RECT 904.020 9.370 907.020 9.380 ;
        RECT 1084.020 9.370 1087.020 9.380 ;
        RECT 1264.020 9.370 1267.020 9.380 ;
        RECT 1444.020 9.370 1447.020 9.380 ;
        RECT 1624.020 9.370 1627.020 9.380 ;
        RECT 1804.020 9.370 1807.020 9.380 ;
        RECT 1984.020 9.370 1987.020 9.380 ;
        RECT 2164.020 9.370 2167.020 9.380 ;
        RECT 2344.020 9.370 2347.020 9.380 ;
        RECT 2524.020 9.370 2527.020 9.380 ;
        RECT 2704.020 9.370 2707.020 9.380 ;
        RECT 2884.020 9.370 2887.020 9.380 ;
        RECT 2926.600 9.370 2929.600 9.380 ;
        RECT -9.980 -1.620 -6.980 -1.610 ;
        RECT 4.020 -1.620 7.020 -1.610 ;
        RECT 184.020 -1.620 187.020 -1.610 ;
        RECT 364.020 -1.620 367.020 -1.610 ;
        RECT 544.020 -1.620 547.020 -1.610 ;
        RECT 724.020 -1.620 727.020 -1.610 ;
        RECT 904.020 -1.620 907.020 -1.610 ;
        RECT 1084.020 -1.620 1087.020 -1.610 ;
        RECT 1264.020 -1.620 1267.020 -1.610 ;
        RECT 1444.020 -1.620 1447.020 -1.610 ;
        RECT 1624.020 -1.620 1627.020 -1.610 ;
        RECT 1804.020 -1.620 1807.020 -1.610 ;
        RECT 1984.020 -1.620 1987.020 -1.610 ;
        RECT 2164.020 -1.620 2167.020 -1.610 ;
        RECT 2344.020 -1.620 2347.020 -1.610 ;
        RECT 2524.020 -1.620 2527.020 -1.610 ;
        RECT 2704.020 -1.620 2707.020 -1.610 ;
        RECT 2884.020 -1.620 2887.020 -1.610 ;
        RECT 2926.600 -1.620 2929.600 -1.610 ;
        RECT -9.980 -4.620 2929.600 -1.620 ;
        RECT -9.980 -4.630 -6.980 -4.620 ;
        RECT 4.020 -4.630 7.020 -4.620 ;
        RECT 184.020 -4.630 187.020 -4.620 ;
        RECT 364.020 -4.630 367.020 -4.620 ;
        RECT 544.020 -4.630 547.020 -4.620 ;
        RECT 724.020 -4.630 727.020 -4.620 ;
        RECT 904.020 -4.630 907.020 -4.620 ;
        RECT 1084.020 -4.630 1087.020 -4.620 ;
        RECT 1264.020 -4.630 1267.020 -4.620 ;
        RECT 1444.020 -4.630 1447.020 -4.620 ;
        RECT 1624.020 -4.630 1627.020 -4.620 ;
        RECT 1804.020 -4.630 1807.020 -4.620 ;
        RECT 1984.020 -4.630 1987.020 -4.620 ;
        RECT 2164.020 -4.630 2167.020 -4.620 ;
        RECT 2344.020 -4.630 2347.020 -4.620 ;
        RECT 2524.020 -4.630 2527.020 -4.620 ;
        RECT 2704.020 -4.630 2707.020 -4.620 ;
        RECT 2884.020 -4.630 2887.020 -4.620 ;
        RECT 2926.600 -4.630 2929.600 -4.620 ;
        RECT -19.380 -11.020 -16.380 -11.010 ;
        RECT 22.020 -11.020 25.020 -11.010 ;
        RECT 202.020 -11.020 205.020 -11.010 ;
        RECT 382.020 -11.020 385.020 -11.010 ;
        RECT 562.020 -11.020 565.020 -11.010 ;
        RECT 742.020 -11.020 745.020 -11.010 ;
        RECT 922.020 -11.020 925.020 -11.010 ;
        RECT 1102.020 -11.020 1105.020 -11.010 ;
        RECT 1282.020 -11.020 1285.020 -11.010 ;
        RECT 1462.020 -11.020 1465.020 -11.010 ;
        RECT 1642.020 -11.020 1645.020 -11.010 ;
        RECT 1822.020 -11.020 1825.020 -11.010 ;
        RECT 2002.020 -11.020 2005.020 -11.010 ;
        RECT 2182.020 -11.020 2185.020 -11.010 ;
        RECT 2362.020 -11.020 2365.020 -11.010 ;
        RECT 2542.020 -11.020 2545.020 -11.010 ;
        RECT 2722.020 -11.020 2725.020 -11.010 ;
        RECT 2902.020 -11.020 2905.020 -11.010 ;
        RECT 2936.000 -11.020 2939.000 -11.010 ;
        RECT -19.380 -14.020 2939.000 -11.020 ;
        RECT -19.380 -14.030 -16.380 -14.020 ;
        RECT 22.020 -14.030 25.020 -14.020 ;
        RECT 202.020 -14.030 205.020 -14.020 ;
        RECT 382.020 -14.030 385.020 -14.020 ;
        RECT 562.020 -14.030 565.020 -14.020 ;
        RECT 742.020 -14.030 745.020 -14.020 ;
        RECT 922.020 -14.030 925.020 -14.020 ;
        RECT 1102.020 -14.030 1105.020 -14.020 ;
        RECT 1282.020 -14.030 1285.020 -14.020 ;
        RECT 1462.020 -14.030 1465.020 -14.020 ;
        RECT 1642.020 -14.030 1645.020 -14.020 ;
        RECT 1822.020 -14.030 1825.020 -14.020 ;
        RECT 2002.020 -14.030 2005.020 -14.020 ;
        RECT 2182.020 -14.030 2185.020 -14.020 ;
        RECT 2362.020 -14.030 2365.020 -14.020 ;
        RECT 2542.020 -14.030 2545.020 -14.020 ;
        RECT 2722.020 -14.030 2725.020 -14.020 ;
        RECT 2902.020 -14.030 2905.020 -14.020 ;
        RECT 2936.000 -14.030 2939.000 -14.020 ;
        RECT -28.780 -20.420 -25.780 -20.410 ;
        RECT 40.020 -20.420 43.020 -20.410 ;
        RECT 220.020 -20.420 223.020 -20.410 ;
        RECT 400.020 -20.420 403.020 -20.410 ;
        RECT 580.020 -20.420 583.020 -20.410 ;
        RECT 760.020 -20.420 763.020 -20.410 ;
        RECT 940.020 -20.420 943.020 -20.410 ;
        RECT 1120.020 -20.420 1123.020 -20.410 ;
        RECT 1300.020 -20.420 1303.020 -20.410 ;
        RECT 1480.020 -20.420 1483.020 -20.410 ;
        RECT 1660.020 -20.420 1663.020 -20.410 ;
        RECT 1840.020 -20.420 1843.020 -20.410 ;
        RECT 2020.020 -20.420 2023.020 -20.410 ;
        RECT 2200.020 -20.420 2203.020 -20.410 ;
        RECT 2380.020 -20.420 2383.020 -20.410 ;
        RECT 2560.020 -20.420 2563.020 -20.410 ;
        RECT 2740.020 -20.420 2743.020 -20.410 ;
        RECT 2945.400 -20.420 2948.400 -20.410 ;
        RECT -28.780 -23.420 2948.400 -20.420 ;
        RECT -28.780 -23.430 -25.780 -23.420 ;
        RECT 40.020 -23.430 43.020 -23.420 ;
        RECT 220.020 -23.430 223.020 -23.420 ;
        RECT 400.020 -23.430 403.020 -23.420 ;
        RECT 580.020 -23.430 583.020 -23.420 ;
        RECT 760.020 -23.430 763.020 -23.420 ;
        RECT 940.020 -23.430 943.020 -23.420 ;
        RECT 1120.020 -23.430 1123.020 -23.420 ;
        RECT 1300.020 -23.430 1303.020 -23.420 ;
        RECT 1480.020 -23.430 1483.020 -23.420 ;
        RECT 1660.020 -23.430 1663.020 -23.420 ;
        RECT 1840.020 -23.430 1843.020 -23.420 ;
        RECT 2020.020 -23.430 2023.020 -23.420 ;
        RECT 2200.020 -23.430 2203.020 -23.420 ;
        RECT 2380.020 -23.430 2383.020 -23.420 ;
        RECT 2560.020 -23.430 2563.020 -23.420 ;
        RECT 2740.020 -23.430 2743.020 -23.420 ;
        RECT 2945.400 -23.430 2948.400 -23.420 ;
        RECT -38.180 -29.820 -35.180 -29.810 ;
        RECT 58.020 -29.820 61.020 -29.810 ;
        RECT 238.020 -29.820 241.020 -29.810 ;
        RECT 418.020 -29.820 421.020 -29.810 ;
        RECT 598.020 -29.820 601.020 -29.810 ;
        RECT 778.020 -29.820 781.020 -29.810 ;
        RECT 958.020 -29.820 961.020 -29.810 ;
        RECT 1138.020 -29.820 1141.020 -29.810 ;
        RECT 1318.020 -29.820 1321.020 -29.810 ;
        RECT 1498.020 -29.820 1501.020 -29.810 ;
        RECT 1678.020 -29.820 1681.020 -29.810 ;
        RECT 1858.020 -29.820 1861.020 -29.810 ;
        RECT 2038.020 -29.820 2041.020 -29.810 ;
        RECT 2218.020 -29.820 2221.020 -29.810 ;
        RECT 2398.020 -29.820 2401.020 -29.810 ;
        RECT 2578.020 -29.820 2581.020 -29.810 ;
        RECT 2758.020 -29.820 2761.020 -29.810 ;
        RECT 2954.800 -29.820 2957.800 -29.810 ;
        RECT -38.180 -32.820 2957.800 -29.820 ;
        RECT -38.180 -32.830 -35.180 -32.820 ;
        RECT 58.020 -32.830 61.020 -32.820 ;
        RECT 238.020 -32.830 241.020 -32.820 ;
        RECT 418.020 -32.830 421.020 -32.820 ;
        RECT 598.020 -32.830 601.020 -32.820 ;
        RECT 778.020 -32.830 781.020 -32.820 ;
        RECT 958.020 -32.830 961.020 -32.820 ;
        RECT 1138.020 -32.830 1141.020 -32.820 ;
        RECT 1318.020 -32.830 1321.020 -32.820 ;
        RECT 1498.020 -32.830 1501.020 -32.820 ;
        RECT 1678.020 -32.830 1681.020 -32.820 ;
        RECT 1858.020 -32.830 1861.020 -32.820 ;
        RECT 2038.020 -32.830 2041.020 -32.820 ;
        RECT 2218.020 -32.830 2221.020 -32.820 ;
        RECT 2398.020 -32.830 2401.020 -32.820 ;
        RECT 2578.020 -32.830 2581.020 -32.820 ;
        RECT 2758.020 -32.830 2761.020 -32.820 ;
        RECT 2954.800 -32.830 2957.800 -32.820 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 681.040 2751.235 686.300 2752.140 ;
        RECT 1331.040 2751.235 1336.300 2752.140 ;
        RECT 1931.040 2751.235 1936.300 2752.140 ;
        RECT 2581.040 2751.235 2586.300 2752.140 ;
        RECT 681.480 2750.400 686.300 2751.235 ;
        RECT 1331.480 2750.400 1336.300 2751.235 ;
        RECT 1931.480 2750.400 1936.300 2751.235 ;
        RECT 2581.480 2750.400 2586.300 2751.235 ;
      LAYER via3 ;
        RECT 684.720 2750.440 686.240 2752.050 ;
        RECT 1334.720 2750.440 1336.240 2752.050 ;
        RECT 1934.720 2750.440 1936.240 2752.050 ;
        RECT 2584.720 2750.440 2586.240 2752.050 ;
      LAYER met4 ;
        RECT -42.880 -37.520 -39.880 3557.200 ;
        RECT -33.480 -28.120 -30.480 3547.800 ;
        RECT -24.080 -18.720 -21.080 3538.400 ;
        RECT -14.680 -9.320 -11.680 3529.000 ;
        RECT 94.020 -9.320 97.020 3529.000 ;
        RECT 112.020 -18.720 115.020 3538.400 ;
        RECT 130.020 -28.120 133.020 3547.800 ;
        RECT 148.020 -37.520 151.020 3557.200 ;
        RECT 274.020 -9.320 277.020 3529.000 ;
        RECT 292.020 2771.235 295.020 3538.400 ;
        RECT 310.020 2771.235 313.020 3547.800 ;
        RECT 328.020 2771.235 331.020 3557.200 ;
        RECT 454.020 2771.235 457.020 3529.000 ;
        RECT 472.020 2771.235 475.020 3538.400 ;
        RECT 490.020 2771.235 493.020 3547.800 ;
        RECT 508.020 2771.235 511.020 3557.200 ;
        RECT 634.020 2771.235 637.020 3529.000 ;
        RECT 652.020 2771.235 655.020 3538.400 ;
        RECT 670.020 2771.235 673.020 3547.800 ;
        RECT 688.020 2771.235 691.020 3557.200 ;
        RECT 684.690 2304.060 686.310 2752.140 ;
        RECT 292.020 2215.000 295.020 2285.000 ;
        RECT 454.020 2215.000 457.020 2285.000 ;
        RECT 472.020 2215.000 475.020 2285.000 ;
        RECT 634.020 2215.000 637.020 2285.000 ;
        RECT 652.020 2215.000 655.020 2285.000 ;
        RECT 814.020 2215.000 817.020 3529.000 ;
        RECT 832.020 2215.000 835.020 3538.400 ;
        RECT 850.020 2215.000 853.020 3547.800 ;
        RECT 868.020 2215.000 871.020 3557.200 ;
        RECT 994.020 2771.235 997.020 3529.000 ;
        RECT 1012.020 2771.235 1015.020 3538.400 ;
        RECT 1030.020 2771.235 1033.020 3547.800 ;
        RECT 1048.020 2771.235 1051.020 3557.200 ;
        RECT 1174.020 2771.235 1177.020 3529.000 ;
        RECT 1192.020 2771.235 1195.020 3538.400 ;
        RECT 1210.020 2771.235 1213.020 3547.800 ;
        RECT 1228.020 2771.235 1231.020 3557.200 ;
        RECT 1334.690 2304.060 1336.310 2752.140 ;
        RECT 994.020 2215.000 997.020 2285.000 ;
        RECT 1012.020 2215.000 1015.020 2285.000 ;
        RECT 1174.020 2215.000 1177.020 2285.000 ;
        RECT 1192.020 2215.000 1195.020 2285.000 ;
        RECT 1354.020 2215.000 1357.020 3529.000 ;
        RECT 1372.020 2215.000 1375.020 3538.400 ;
        RECT 1390.020 2215.000 1393.020 3547.800 ;
        RECT 1408.020 2215.000 1411.020 3557.200 ;
        RECT 1534.020 2771.235 1537.020 3529.000 ;
        RECT 1552.020 2771.235 1555.020 3538.400 ;
        RECT 1570.020 2771.235 1573.020 3547.800 ;
        RECT 1588.020 2771.235 1591.020 3557.200 ;
        RECT 1714.020 2771.235 1717.020 3529.000 ;
        RECT 1732.020 2771.235 1735.020 3538.400 ;
        RECT 1750.020 2771.235 1753.020 3547.800 ;
        RECT 1768.020 2771.235 1771.020 3557.200 ;
        RECT 1894.020 2771.235 1897.020 3529.000 ;
        RECT 1912.020 2771.235 1915.020 3538.400 ;
        RECT 1930.020 2771.235 1933.020 3547.800 ;
        RECT 1948.020 2771.235 1951.020 3557.200 ;
        RECT 1934.690 2304.060 1936.310 2752.140 ;
        RECT 397.840 1010.640 399.440 2188.880 ;
        RECT 292.020 -18.720 295.020 985.000 ;
        RECT 310.020 -28.120 313.020 985.000 ;
        RECT 328.020 -37.520 331.020 985.000 ;
        RECT 454.020 -9.320 457.020 985.000 ;
        RECT 472.020 -18.720 475.020 985.000 ;
        RECT 490.020 -28.120 493.020 985.000 ;
        RECT 508.020 -37.520 511.020 985.000 ;
        RECT 634.020 -9.320 637.020 985.000 ;
        RECT 652.020 -18.720 655.020 985.000 ;
        RECT 670.020 -28.120 673.020 985.000 ;
        RECT 688.020 -37.520 691.020 985.000 ;
        RECT 814.020 -9.320 817.020 985.000 ;
        RECT 832.020 -18.720 835.020 985.000 ;
        RECT 850.020 -28.120 853.020 985.000 ;
        RECT 868.020 -37.520 871.020 985.000 ;
        RECT 994.020 -9.320 997.020 985.000 ;
        RECT 1012.020 -18.720 1015.020 985.000 ;
        RECT 1030.020 -28.120 1033.020 985.000 ;
        RECT 1048.020 -37.520 1051.020 985.000 ;
        RECT 1174.020 -9.320 1177.020 985.000 ;
        RECT 1192.020 -18.720 1195.020 985.000 ;
        RECT 1210.020 -28.120 1213.020 985.000 ;
        RECT 1228.020 -37.520 1231.020 985.000 ;
        RECT 1354.020 -9.320 1357.020 985.000 ;
        RECT 1372.020 -18.720 1375.020 985.000 ;
        RECT 1390.020 -28.120 1393.020 985.000 ;
        RECT 1408.020 -37.520 1411.020 985.000 ;
        RECT 1534.020 -9.320 1537.020 2285.000 ;
        RECT 1552.020 -18.720 1555.020 2285.000 ;
        RECT 1570.020 -28.120 1573.020 2285.000 ;
        RECT 1588.020 -37.520 1591.020 2285.000 ;
        RECT 1714.020 -9.320 1717.020 2285.000 ;
        RECT 1732.020 -18.720 1735.020 2285.000 ;
        RECT 1750.020 -28.120 1753.020 2285.000 ;
        RECT 1768.020 -37.520 1771.020 2285.000 ;
        RECT 1894.020 -9.320 1897.020 2285.000 ;
        RECT 1912.020 -18.720 1915.020 2285.000 ;
        RECT 1930.020 -28.120 1933.020 2285.000 ;
        RECT 1948.020 -37.520 1951.020 2285.000 ;
        RECT 2074.020 -9.320 2077.020 3529.000 ;
        RECT 2092.020 -18.720 2095.020 3538.400 ;
        RECT 2110.020 -28.120 2113.020 3547.800 ;
        RECT 2128.020 -37.520 2131.020 3557.200 ;
        RECT 2254.020 2771.235 2257.020 3529.000 ;
        RECT 2272.020 2771.235 2275.020 3538.400 ;
        RECT 2290.020 2771.235 2293.020 3547.800 ;
        RECT 2308.020 2771.235 2311.020 3557.200 ;
        RECT 2434.020 2771.235 2437.020 3529.000 ;
        RECT 2452.020 2771.235 2455.020 3538.400 ;
        RECT 2470.020 2771.235 2473.020 3547.800 ;
        RECT 2488.020 2771.235 2491.020 3557.200 ;
        RECT 2584.690 2304.060 2586.310 2752.140 ;
        RECT 2254.020 -9.320 2257.020 2285.000 ;
        RECT 2272.020 -18.720 2275.020 2285.000 ;
        RECT 2290.020 -28.120 2293.020 2285.000 ;
        RECT 2308.020 -37.520 2311.020 2285.000 ;
        RECT 2434.020 -9.320 2437.020 2285.000 ;
        RECT 2452.020 -18.720 2455.020 2285.000 ;
        RECT 2470.020 -28.120 2473.020 2285.000 ;
        RECT 2488.020 -37.520 2491.020 2285.000 ;
        RECT 2614.020 -9.320 2617.020 3529.000 ;
        RECT 2632.020 -18.720 2635.020 3538.400 ;
        RECT 2650.020 -28.120 2653.020 3547.800 ;
        RECT 2668.020 -37.520 2671.020 3557.200 ;
        RECT 2794.020 -9.320 2797.020 3529.000 ;
        RECT 2812.020 -18.720 2815.020 3538.400 ;
        RECT 2830.020 -28.120 2833.020 3547.800 ;
        RECT 2848.020 -37.520 2851.020 3557.200 ;
        RECT 2931.300 -9.320 2934.300 3529.000 ;
        RECT 2940.700 -18.720 2943.700 3538.400 ;
        RECT 2950.100 -28.120 2953.100 3547.800 ;
        RECT 2959.500 -37.520 2962.500 3557.200 ;
      LAYER via4 ;
        RECT -41.970 3555.910 -40.790 3557.090 ;
        RECT -41.970 3554.310 -40.790 3555.490 ;
        RECT 148.930 3555.910 150.110 3557.090 ;
        RECT 148.930 3554.310 150.110 3555.490 ;
        RECT -41.970 3395.090 -40.790 3396.270 ;
        RECT -41.970 3393.490 -40.790 3394.670 ;
        RECT -41.970 3215.090 -40.790 3216.270 ;
        RECT -41.970 3213.490 -40.790 3214.670 ;
        RECT -41.970 3035.090 -40.790 3036.270 ;
        RECT -41.970 3033.490 -40.790 3034.670 ;
        RECT -41.970 2855.090 -40.790 2856.270 ;
        RECT -41.970 2853.490 -40.790 2854.670 ;
        RECT -41.970 2675.090 -40.790 2676.270 ;
        RECT -41.970 2673.490 -40.790 2674.670 ;
        RECT -41.970 2495.090 -40.790 2496.270 ;
        RECT -41.970 2493.490 -40.790 2494.670 ;
        RECT -41.970 2315.090 -40.790 2316.270 ;
        RECT -41.970 2313.490 -40.790 2314.670 ;
        RECT -41.970 2135.090 -40.790 2136.270 ;
        RECT -41.970 2133.490 -40.790 2134.670 ;
        RECT -41.970 1955.090 -40.790 1956.270 ;
        RECT -41.970 1953.490 -40.790 1954.670 ;
        RECT -41.970 1775.090 -40.790 1776.270 ;
        RECT -41.970 1773.490 -40.790 1774.670 ;
        RECT -41.970 1595.090 -40.790 1596.270 ;
        RECT -41.970 1593.490 -40.790 1594.670 ;
        RECT -41.970 1415.090 -40.790 1416.270 ;
        RECT -41.970 1413.490 -40.790 1414.670 ;
        RECT -41.970 1235.090 -40.790 1236.270 ;
        RECT -41.970 1233.490 -40.790 1234.670 ;
        RECT -41.970 1055.090 -40.790 1056.270 ;
        RECT -41.970 1053.490 -40.790 1054.670 ;
        RECT -41.970 875.090 -40.790 876.270 ;
        RECT -41.970 873.490 -40.790 874.670 ;
        RECT -41.970 695.090 -40.790 696.270 ;
        RECT -41.970 693.490 -40.790 694.670 ;
        RECT -41.970 515.090 -40.790 516.270 ;
        RECT -41.970 513.490 -40.790 514.670 ;
        RECT -41.970 335.090 -40.790 336.270 ;
        RECT -41.970 333.490 -40.790 334.670 ;
        RECT -41.970 155.090 -40.790 156.270 ;
        RECT -41.970 153.490 -40.790 154.670 ;
        RECT -32.570 3546.510 -31.390 3547.690 ;
        RECT -32.570 3544.910 -31.390 3546.090 ;
        RECT 130.930 3546.510 132.110 3547.690 ;
        RECT 130.930 3544.910 132.110 3546.090 ;
        RECT -32.570 3377.090 -31.390 3378.270 ;
        RECT -32.570 3375.490 -31.390 3376.670 ;
        RECT -32.570 3197.090 -31.390 3198.270 ;
        RECT -32.570 3195.490 -31.390 3196.670 ;
        RECT -32.570 3017.090 -31.390 3018.270 ;
        RECT -32.570 3015.490 -31.390 3016.670 ;
        RECT -32.570 2837.090 -31.390 2838.270 ;
        RECT -32.570 2835.490 -31.390 2836.670 ;
        RECT -32.570 2657.090 -31.390 2658.270 ;
        RECT -32.570 2655.490 -31.390 2656.670 ;
        RECT -32.570 2477.090 -31.390 2478.270 ;
        RECT -32.570 2475.490 -31.390 2476.670 ;
        RECT -32.570 2297.090 -31.390 2298.270 ;
        RECT -32.570 2295.490 -31.390 2296.670 ;
        RECT -32.570 2117.090 -31.390 2118.270 ;
        RECT -32.570 2115.490 -31.390 2116.670 ;
        RECT -32.570 1937.090 -31.390 1938.270 ;
        RECT -32.570 1935.490 -31.390 1936.670 ;
        RECT -32.570 1757.090 -31.390 1758.270 ;
        RECT -32.570 1755.490 -31.390 1756.670 ;
        RECT -32.570 1577.090 -31.390 1578.270 ;
        RECT -32.570 1575.490 -31.390 1576.670 ;
        RECT -32.570 1397.090 -31.390 1398.270 ;
        RECT -32.570 1395.490 -31.390 1396.670 ;
        RECT -32.570 1217.090 -31.390 1218.270 ;
        RECT -32.570 1215.490 -31.390 1216.670 ;
        RECT -32.570 1037.090 -31.390 1038.270 ;
        RECT -32.570 1035.490 -31.390 1036.670 ;
        RECT -32.570 857.090 -31.390 858.270 ;
        RECT -32.570 855.490 -31.390 856.670 ;
        RECT -32.570 677.090 -31.390 678.270 ;
        RECT -32.570 675.490 -31.390 676.670 ;
        RECT -32.570 497.090 -31.390 498.270 ;
        RECT -32.570 495.490 -31.390 496.670 ;
        RECT -32.570 317.090 -31.390 318.270 ;
        RECT -32.570 315.490 -31.390 316.670 ;
        RECT -32.570 137.090 -31.390 138.270 ;
        RECT -32.570 135.490 -31.390 136.670 ;
        RECT -23.170 3537.110 -21.990 3538.290 ;
        RECT -23.170 3535.510 -21.990 3536.690 ;
        RECT 112.930 3537.110 114.110 3538.290 ;
        RECT 112.930 3535.510 114.110 3536.690 ;
        RECT -23.170 3359.090 -21.990 3360.270 ;
        RECT -23.170 3357.490 -21.990 3358.670 ;
        RECT -23.170 3179.090 -21.990 3180.270 ;
        RECT -23.170 3177.490 -21.990 3178.670 ;
        RECT -23.170 2999.090 -21.990 3000.270 ;
        RECT -23.170 2997.490 -21.990 2998.670 ;
        RECT -23.170 2819.090 -21.990 2820.270 ;
        RECT -23.170 2817.490 -21.990 2818.670 ;
        RECT -23.170 2639.090 -21.990 2640.270 ;
        RECT -23.170 2637.490 -21.990 2638.670 ;
        RECT -23.170 2459.090 -21.990 2460.270 ;
        RECT -23.170 2457.490 -21.990 2458.670 ;
        RECT -23.170 2279.090 -21.990 2280.270 ;
        RECT -23.170 2277.490 -21.990 2278.670 ;
        RECT -23.170 2099.090 -21.990 2100.270 ;
        RECT -23.170 2097.490 -21.990 2098.670 ;
        RECT -23.170 1919.090 -21.990 1920.270 ;
        RECT -23.170 1917.490 -21.990 1918.670 ;
        RECT -23.170 1739.090 -21.990 1740.270 ;
        RECT -23.170 1737.490 -21.990 1738.670 ;
        RECT -23.170 1559.090 -21.990 1560.270 ;
        RECT -23.170 1557.490 -21.990 1558.670 ;
        RECT -23.170 1379.090 -21.990 1380.270 ;
        RECT -23.170 1377.490 -21.990 1378.670 ;
        RECT -23.170 1199.090 -21.990 1200.270 ;
        RECT -23.170 1197.490 -21.990 1198.670 ;
        RECT -23.170 1019.090 -21.990 1020.270 ;
        RECT -23.170 1017.490 -21.990 1018.670 ;
        RECT -23.170 839.090 -21.990 840.270 ;
        RECT -23.170 837.490 -21.990 838.670 ;
        RECT -23.170 659.090 -21.990 660.270 ;
        RECT -23.170 657.490 -21.990 658.670 ;
        RECT -23.170 479.090 -21.990 480.270 ;
        RECT -23.170 477.490 -21.990 478.670 ;
        RECT -23.170 299.090 -21.990 300.270 ;
        RECT -23.170 297.490 -21.990 298.670 ;
        RECT -23.170 119.090 -21.990 120.270 ;
        RECT -23.170 117.490 -21.990 118.670 ;
        RECT -13.770 3527.710 -12.590 3528.890 ;
        RECT -13.770 3526.110 -12.590 3527.290 ;
        RECT -13.770 3341.090 -12.590 3342.270 ;
        RECT -13.770 3339.490 -12.590 3340.670 ;
        RECT -13.770 3161.090 -12.590 3162.270 ;
        RECT -13.770 3159.490 -12.590 3160.670 ;
        RECT -13.770 2981.090 -12.590 2982.270 ;
        RECT -13.770 2979.490 -12.590 2980.670 ;
        RECT -13.770 2801.090 -12.590 2802.270 ;
        RECT -13.770 2799.490 -12.590 2800.670 ;
        RECT -13.770 2621.090 -12.590 2622.270 ;
        RECT -13.770 2619.490 -12.590 2620.670 ;
        RECT -13.770 2441.090 -12.590 2442.270 ;
        RECT -13.770 2439.490 -12.590 2440.670 ;
        RECT -13.770 2261.090 -12.590 2262.270 ;
        RECT -13.770 2259.490 -12.590 2260.670 ;
        RECT -13.770 2081.090 -12.590 2082.270 ;
        RECT -13.770 2079.490 -12.590 2080.670 ;
        RECT -13.770 1901.090 -12.590 1902.270 ;
        RECT -13.770 1899.490 -12.590 1900.670 ;
        RECT -13.770 1721.090 -12.590 1722.270 ;
        RECT -13.770 1719.490 -12.590 1720.670 ;
        RECT -13.770 1541.090 -12.590 1542.270 ;
        RECT -13.770 1539.490 -12.590 1540.670 ;
        RECT -13.770 1361.090 -12.590 1362.270 ;
        RECT -13.770 1359.490 -12.590 1360.670 ;
        RECT -13.770 1181.090 -12.590 1182.270 ;
        RECT -13.770 1179.490 -12.590 1180.670 ;
        RECT -13.770 1001.090 -12.590 1002.270 ;
        RECT -13.770 999.490 -12.590 1000.670 ;
        RECT -13.770 821.090 -12.590 822.270 ;
        RECT -13.770 819.490 -12.590 820.670 ;
        RECT -13.770 641.090 -12.590 642.270 ;
        RECT -13.770 639.490 -12.590 640.670 ;
        RECT -13.770 461.090 -12.590 462.270 ;
        RECT -13.770 459.490 -12.590 460.670 ;
        RECT -13.770 281.090 -12.590 282.270 ;
        RECT -13.770 279.490 -12.590 280.670 ;
        RECT -13.770 101.090 -12.590 102.270 ;
        RECT -13.770 99.490 -12.590 100.670 ;
        RECT -13.770 -7.610 -12.590 -6.430 ;
        RECT -13.770 -9.210 -12.590 -8.030 ;
        RECT 94.930 3527.710 96.110 3528.890 ;
        RECT 94.930 3526.110 96.110 3527.290 ;
        RECT 94.930 3341.090 96.110 3342.270 ;
        RECT 94.930 3339.490 96.110 3340.670 ;
        RECT 94.930 3161.090 96.110 3162.270 ;
        RECT 94.930 3159.490 96.110 3160.670 ;
        RECT 94.930 2981.090 96.110 2982.270 ;
        RECT 94.930 2979.490 96.110 2980.670 ;
        RECT 94.930 2801.090 96.110 2802.270 ;
        RECT 94.930 2799.490 96.110 2800.670 ;
        RECT 94.930 2621.090 96.110 2622.270 ;
        RECT 94.930 2619.490 96.110 2620.670 ;
        RECT 94.930 2441.090 96.110 2442.270 ;
        RECT 94.930 2439.490 96.110 2440.670 ;
        RECT 94.930 2261.090 96.110 2262.270 ;
        RECT 94.930 2259.490 96.110 2260.670 ;
        RECT 94.930 2081.090 96.110 2082.270 ;
        RECT 94.930 2079.490 96.110 2080.670 ;
        RECT 94.930 1901.090 96.110 1902.270 ;
        RECT 94.930 1899.490 96.110 1900.670 ;
        RECT 94.930 1721.090 96.110 1722.270 ;
        RECT 94.930 1719.490 96.110 1720.670 ;
        RECT 94.930 1541.090 96.110 1542.270 ;
        RECT 94.930 1539.490 96.110 1540.670 ;
        RECT 94.930 1361.090 96.110 1362.270 ;
        RECT 94.930 1359.490 96.110 1360.670 ;
        RECT 94.930 1181.090 96.110 1182.270 ;
        RECT 94.930 1179.490 96.110 1180.670 ;
        RECT 94.930 1001.090 96.110 1002.270 ;
        RECT 94.930 999.490 96.110 1000.670 ;
        RECT 94.930 821.090 96.110 822.270 ;
        RECT 94.930 819.490 96.110 820.670 ;
        RECT 94.930 641.090 96.110 642.270 ;
        RECT 94.930 639.490 96.110 640.670 ;
        RECT 94.930 461.090 96.110 462.270 ;
        RECT 94.930 459.490 96.110 460.670 ;
        RECT 94.930 281.090 96.110 282.270 ;
        RECT 94.930 279.490 96.110 280.670 ;
        RECT 94.930 101.090 96.110 102.270 ;
        RECT 94.930 99.490 96.110 100.670 ;
        RECT 94.930 -7.610 96.110 -6.430 ;
        RECT 94.930 -9.210 96.110 -8.030 ;
        RECT 112.930 3359.090 114.110 3360.270 ;
        RECT 112.930 3357.490 114.110 3358.670 ;
        RECT 112.930 3179.090 114.110 3180.270 ;
        RECT 112.930 3177.490 114.110 3178.670 ;
        RECT 112.930 2999.090 114.110 3000.270 ;
        RECT 112.930 2997.490 114.110 2998.670 ;
        RECT 112.930 2819.090 114.110 2820.270 ;
        RECT 112.930 2817.490 114.110 2818.670 ;
        RECT 112.930 2639.090 114.110 2640.270 ;
        RECT 112.930 2637.490 114.110 2638.670 ;
        RECT 112.930 2459.090 114.110 2460.270 ;
        RECT 112.930 2457.490 114.110 2458.670 ;
        RECT 112.930 2279.090 114.110 2280.270 ;
        RECT 112.930 2277.490 114.110 2278.670 ;
        RECT 112.930 2099.090 114.110 2100.270 ;
        RECT 112.930 2097.490 114.110 2098.670 ;
        RECT 112.930 1919.090 114.110 1920.270 ;
        RECT 112.930 1917.490 114.110 1918.670 ;
        RECT 112.930 1739.090 114.110 1740.270 ;
        RECT 112.930 1737.490 114.110 1738.670 ;
        RECT 112.930 1559.090 114.110 1560.270 ;
        RECT 112.930 1557.490 114.110 1558.670 ;
        RECT 112.930 1379.090 114.110 1380.270 ;
        RECT 112.930 1377.490 114.110 1378.670 ;
        RECT 112.930 1199.090 114.110 1200.270 ;
        RECT 112.930 1197.490 114.110 1198.670 ;
        RECT 112.930 1019.090 114.110 1020.270 ;
        RECT 112.930 1017.490 114.110 1018.670 ;
        RECT 112.930 839.090 114.110 840.270 ;
        RECT 112.930 837.490 114.110 838.670 ;
        RECT 112.930 659.090 114.110 660.270 ;
        RECT 112.930 657.490 114.110 658.670 ;
        RECT 112.930 479.090 114.110 480.270 ;
        RECT 112.930 477.490 114.110 478.670 ;
        RECT 112.930 299.090 114.110 300.270 ;
        RECT 112.930 297.490 114.110 298.670 ;
        RECT 112.930 119.090 114.110 120.270 ;
        RECT 112.930 117.490 114.110 118.670 ;
        RECT -23.170 -17.010 -21.990 -15.830 ;
        RECT -23.170 -18.610 -21.990 -17.430 ;
        RECT 112.930 -17.010 114.110 -15.830 ;
        RECT 112.930 -18.610 114.110 -17.430 ;
        RECT 130.930 3377.090 132.110 3378.270 ;
        RECT 130.930 3375.490 132.110 3376.670 ;
        RECT 130.930 3197.090 132.110 3198.270 ;
        RECT 130.930 3195.490 132.110 3196.670 ;
        RECT 130.930 3017.090 132.110 3018.270 ;
        RECT 130.930 3015.490 132.110 3016.670 ;
        RECT 130.930 2837.090 132.110 2838.270 ;
        RECT 130.930 2835.490 132.110 2836.670 ;
        RECT 130.930 2657.090 132.110 2658.270 ;
        RECT 130.930 2655.490 132.110 2656.670 ;
        RECT 130.930 2477.090 132.110 2478.270 ;
        RECT 130.930 2475.490 132.110 2476.670 ;
        RECT 130.930 2297.090 132.110 2298.270 ;
        RECT 130.930 2295.490 132.110 2296.670 ;
        RECT 130.930 2117.090 132.110 2118.270 ;
        RECT 130.930 2115.490 132.110 2116.670 ;
        RECT 130.930 1937.090 132.110 1938.270 ;
        RECT 130.930 1935.490 132.110 1936.670 ;
        RECT 130.930 1757.090 132.110 1758.270 ;
        RECT 130.930 1755.490 132.110 1756.670 ;
        RECT 130.930 1577.090 132.110 1578.270 ;
        RECT 130.930 1575.490 132.110 1576.670 ;
        RECT 130.930 1397.090 132.110 1398.270 ;
        RECT 130.930 1395.490 132.110 1396.670 ;
        RECT 130.930 1217.090 132.110 1218.270 ;
        RECT 130.930 1215.490 132.110 1216.670 ;
        RECT 130.930 1037.090 132.110 1038.270 ;
        RECT 130.930 1035.490 132.110 1036.670 ;
        RECT 130.930 857.090 132.110 858.270 ;
        RECT 130.930 855.490 132.110 856.670 ;
        RECT 130.930 677.090 132.110 678.270 ;
        RECT 130.930 675.490 132.110 676.670 ;
        RECT 130.930 497.090 132.110 498.270 ;
        RECT 130.930 495.490 132.110 496.670 ;
        RECT 130.930 317.090 132.110 318.270 ;
        RECT 130.930 315.490 132.110 316.670 ;
        RECT 130.930 137.090 132.110 138.270 ;
        RECT 130.930 135.490 132.110 136.670 ;
        RECT -32.570 -26.410 -31.390 -25.230 ;
        RECT -32.570 -28.010 -31.390 -26.830 ;
        RECT 130.930 -26.410 132.110 -25.230 ;
        RECT 130.930 -28.010 132.110 -26.830 ;
        RECT 328.930 3555.910 330.110 3557.090 ;
        RECT 328.930 3554.310 330.110 3555.490 ;
        RECT 310.930 3546.510 312.110 3547.690 ;
        RECT 310.930 3544.910 312.110 3546.090 ;
        RECT 292.930 3537.110 294.110 3538.290 ;
        RECT 292.930 3535.510 294.110 3536.690 ;
        RECT 148.930 3395.090 150.110 3396.270 ;
        RECT 148.930 3393.490 150.110 3394.670 ;
        RECT 148.930 3215.090 150.110 3216.270 ;
        RECT 148.930 3213.490 150.110 3214.670 ;
        RECT 148.930 3035.090 150.110 3036.270 ;
        RECT 148.930 3033.490 150.110 3034.670 ;
        RECT 148.930 2855.090 150.110 2856.270 ;
        RECT 148.930 2853.490 150.110 2854.670 ;
        RECT 148.930 2675.090 150.110 2676.270 ;
        RECT 148.930 2673.490 150.110 2674.670 ;
        RECT 148.930 2495.090 150.110 2496.270 ;
        RECT 148.930 2493.490 150.110 2494.670 ;
        RECT 148.930 2315.090 150.110 2316.270 ;
        RECT 148.930 2313.490 150.110 2314.670 ;
        RECT 148.930 2135.090 150.110 2136.270 ;
        RECT 148.930 2133.490 150.110 2134.670 ;
        RECT 148.930 1955.090 150.110 1956.270 ;
        RECT 148.930 1953.490 150.110 1954.670 ;
        RECT 148.930 1775.090 150.110 1776.270 ;
        RECT 148.930 1773.490 150.110 1774.670 ;
        RECT 148.930 1595.090 150.110 1596.270 ;
        RECT 148.930 1593.490 150.110 1594.670 ;
        RECT 148.930 1415.090 150.110 1416.270 ;
        RECT 148.930 1413.490 150.110 1414.670 ;
        RECT 148.930 1235.090 150.110 1236.270 ;
        RECT 148.930 1233.490 150.110 1234.670 ;
        RECT 148.930 1055.090 150.110 1056.270 ;
        RECT 148.930 1053.490 150.110 1054.670 ;
        RECT 148.930 875.090 150.110 876.270 ;
        RECT 148.930 873.490 150.110 874.670 ;
        RECT 148.930 695.090 150.110 696.270 ;
        RECT 148.930 693.490 150.110 694.670 ;
        RECT 148.930 515.090 150.110 516.270 ;
        RECT 148.930 513.490 150.110 514.670 ;
        RECT 148.930 335.090 150.110 336.270 ;
        RECT 148.930 333.490 150.110 334.670 ;
        RECT 148.930 155.090 150.110 156.270 ;
        RECT 148.930 153.490 150.110 154.670 ;
        RECT -41.970 -35.810 -40.790 -34.630 ;
        RECT -41.970 -37.410 -40.790 -36.230 ;
        RECT 274.930 3527.710 276.110 3528.890 ;
        RECT 274.930 3526.110 276.110 3527.290 ;
        RECT 274.930 3341.090 276.110 3342.270 ;
        RECT 274.930 3339.490 276.110 3340.670 ;
        RECT 274.930 3161.090 276.110 3162.270 ;
        RECT 274.930 3159.490 276.110 3160.670 ;
        RECT 274.930 2981.090 276.110 2982.270 ;
        RECT 274.930 2979.490 276.110 2980.670 ;
        RECT 274.930 2801.090 276.110 2802.270 ;
        RECT 274.930 2799.490 276.110 2800.670 ;
        RECT 292.930 3359.090 294.110 3360.270 ;
        RECT 292.930 3357.490 294.110 3358.670 ;
        RECT 292.930 3179.090 294.110 3180.270 ;
        RECT 292.930 3177.490 294.110 3178.670 ;
        RECT 292.930 2999.090 294.110 3000.270 ;
        RECT 292.930 2997.490 294.110 2998.670 ;
        RECT 292.930 2819.090 294.110 2820.270 ;
        RECT 292.930 2817.490 294.110 2818.670 ;
        RECT 310.930 3377.090 312.110 3378.270 ;
        RECT 310.930 3375.490 312.110 3376.670 ;
        RECT 310.930 3197.090 312.110 3198.270 ;
        RECT 310.930 3195.490 312.110 3196.670 ;
        RECT 310.930 3017.090 312.110 3018.270 ;
        RECT 310.930 3015.490 312.110 3016.670 ;
        RECT 310.930 2837.090 312.110 2838.270 ;
        RECT 310.930 2835.490 312.110 2836.670 ;
        RECT 508.930 3555.910 510.110 3557.090 ;
        RECT 508.930 3554.310 510.110 3555.490 ;
        RECT 490.930 3546.510 492.110 3547.690 ;
        RECT 490.930 3544.910 492.110 3546.090 ;
        RECT 472.930 3537.110 474.110 3538.290 ;
        RECT 472.930 3535.510 474.110 3536.690 ;
        RECT 328.930 3395.090 330.110 3396.270 ;
        RECT 328.930 3393.490 330.110 3394.670 ;
        RECT 328.930 3215.090 330.110 3216.270 ;
        RECT 328.930 3213.490 330.110 3214.670 ;
        RECT 328.930 3035.090 330.110 3036.270 ;
        RECT 328.930 3033.490 330.110 3034.670 ;
        RECT 328.930 2855.090 330.110 2856.270 ;
        RECT 328.930 2853.490 330.110 2854.670 ;
        RECT 454.930 3527.710 456.110 3528.890 ;
        RECT 454.930 3526.110 456.110 3527.290 ;
        RECT 454.930 3341.090 456.110 3342.270 ;
        RECT 454.930 3339.490 456.110 3340.670 ;
        RECT 454.930 3161.090 456.110 3162.270 ;
        RECT 454.930 3159.490 456.110 3160.670 ;
        RECT 454.930 2981.090 456.110 2982.270 ;
        RECT 454.930 2979.490 456.110 2980.670 ;
        RECT 454.930 2801.090 456.110 2802.270 ;
        RECT 454.930 2799.490 456.110 2800.670 ;
        RECT 472.930 3359.090 474.110 3360.270 ;
        RECT 472.930 3357.490 474.110 3358.670 ;
        RECT 472.930 3179.090 474.110 3180.270 ;
        RECT 472.930 3177.490 474.110 3178.670 ;
        RECT 472.930 2999.090 474.110 3000.270 ;
        RECT 472.930 2997.490 474.110 2998.670 ;
        RECT 472.930 2819.090 474.110 2820.270 ;
        RECT 472.930 2817.490 474.110 2818.670 ;
        RECT 490.930 3377.090 492.110 3378.270 ;
        RECT 490.930 3375.490 492.110 3376.670 ;
        RECT 490.930 3197.090 492.110 3198.270 ;
        RECT 490.930 3195.490 492.110 3196.670 ;
        RECT 490.930 3017.090 492.110 3018.270 ;
        RECT 490.930 3015.490 492.110 3016.670 ;
        RECT 490.930 2837.090 492.110 2838.270 ;
        RECT 490.930 2835.490 492.110 2836.670 ;
        RECT 688.930 3555.910 690.110 3557.090 ;
        RECT 688.930 3554.310 690.110 3555.490 ;
        RECT 670.930 3546.510 672.110 3547.690 ;
        RECT 670.930 3544.910 672.110 3546.090 ;
        RECT 652.930 3537.110 654.110 3538.290 ;
        RECT 652.930 3535.510 654.110 3536.690 ;
        RECT 508.930 3395.090 510.110 3396.270 ;
        RECT 508.930 3393.490 510.110 3394.670 ;
        RECT 508.930 3215.090 510.110 3216.270 ;
        RECT 508.930 3213.490 510.110 3214.670 ;
        RECT 508.930 3035.090 510.110 3036.270 ;
        RECT 508.930 3033.490 510.110 3034.670 ;
        RECT 508.930 2855.090 510.110 2856.270 ;
        RECT 508.930 2853.490 510.110 2854.670 ;
        RECT 634.930 3527.710 636.110 3528.890 ;
        RECT 634.930 3526.110 636.110 3527.290 ;
        RECT 634.930 3341.090 636.110 3342.270 ;
        RECT 634.930 3339.490 636.110 3340.670 ;
        RECT 634.930 3161.090 636.110 3162.270 ;
        RECT 634.930 3159.490 636.110 3160.670 ;
        RECT 634.930 2981.090 636.110 2982.270 ;
        RECT 634.930 2979.490 636.110 2980.670 ;
        RECT 634.930 2801.090 636.110 2802.270 ;
        RECT 634.930 2799.490 636.110 2800.670 ;
        RECT 652.930 3359.090 654.110 3360.270 ;
        RECT 652.930 3357.490 654.110 3358.670 ;
        RECT 652.930 3179.090 654.110 3180.270 ;
        RECT 652.930 3177.490 654.110 3178.670 ;
        RECT 652.930 2999.090 654.110 3000.270 ;
        RECT 652.930 2997.490 654.110 2998.670 ;
        RECT 652.930 2819.090 654.110 2820.270 ;
        RECT 652.930 2817.490 654.110 2818.670 ;
        RECT 670.930 3377.090 672.110 3378.270 ;
        RECT 670.930 3375.490 672.110 3376.670 ;
        RECT 670.930 3197.090 672.110 3198.270 ;
        RECT 670.930 3195.490 672.110 3196.670 ;
        RECT 670.930 3017.090 672.110 3018.270 ;
        RECT 670.930 3015.490 672.110 3016.670 ;
        RECT 670.930 2837.090 672.110 2838.270 ;
        RECT 670.930 2835.490 672.110 2836.670 ;
        RECT 868.930 3555.910 870.110 3557.090 ;
        RECT 868.930 3554.310 870.110 3555.490 ;
        RECT 850.930 3546.510 852.110 3547.690 ;
        RECT 850.930 3544.910 852.110 3546.090 ;
        RECT 832.930 3537.110 834.110 3538.290 ;
        RECT 832.930 3535.510 834.110 3536.690 ;
        RECT 688.930 3395.090 690.110 3396.270 ;
        RECT 688.930 3393.490 690.110 3394.670 ;
        RECT 688.930 3215.090 690.110 3216.270 ;
        RECT 688.930 3213.490 690.110 3214.670 ;
        RECT 688.930 3035.090 690.110 3036.270 ;
        RECT 688.930 3033.490 690.110 3034.670 ;
        RECT 688.930 2855.090 690.110 2856.270 ;
        RECT 688.930 2853.490 690.110 2854.670 ;
        RECT 814.930 3527.710 816.110 3528.890 ;
        RECT 814.930 3526.110 816.110 3527.290 ;
        RECT 814.930 3341.090 816.110 3342.270 ;
        RECT 814.930 3339.490 816.110 3340.670 ;
        RECT 814.930 3161.090 816.110 3162.270 ;
        RECT 814.930 3159.490 816.110 3160.670 ;
        RECT 814.930 2981.090 816.110 2982.270 ;
        RECT 814.930 2979.490 816.110 2980.670 ;
        RECT 814.930 2801.090 816.110 2802.270 ;
        RECT 814.930 2799.490 816.110 2800.670 ;
        RECT 274.930 2621.090 276.110 2622.270 ;
        RECT 274.930 2619.490 276.110 2620.670 ;
        RECT 274.930 2441.090 276.110 2442.270 ;
        RECT 274.930 2439.490 276.110 2440.670 ;
        RECT 684.910 2675.090 686.090 2676.270 ;
        RECT 684.910 2673.490 686.090 2674.670 ;
        RECT 684.910 2657.090 686.090 2658.270 ;
        RECT 684.910 2655.490 686.090 2656.670 ;
        RECT 684.910 2639.090 686.090 2640.270 ;
        RECT 684.910 2637.490 686.090 2638.670 ;
        RECT 684.910 2621.090 686.090 2622.270 ;
        RECT 684.910 2619.490 686.090 2620.670 ;
        RECT 684.910 2495.090 686.090 2496.270 ;
        RECT 684.910 2493.490 686.090 2494.670 ;
        RECT 684.910 2477.090 686.090 2478.270 ;
        RECT 684.910 2475.490 686.090 2476.670 ;
        RECT 684.910 2459.090 686.090 2460.270 ;
        RECT 684.910 2457.490 686.090 2458.670 ;
        RECT 684.910 2441.090 686.090 2442.270 ;
        RECT 684.910 2439.490 686.090 2440.670 ;
        RECT 684.910 2315.090 686.090 2316.270 ;
        RECT 684.910 2313.490 686.090 2314.670 ;
        RECT 814.930 2621.090 816.110 2622.270 ;
        RECT 814.930 2619.490 816.110 2620.670 ;
        RECT 814.930 2441.090 816.110 2442.270 ;
        RECT 814.930 2439.490 816.110 2440.670 ;
        RECT 274.930 2261.090 276.110 2262.270 ;
        RECT 274.930 2259.490 276.110 2260.670 ;
        RECT 292.930 2279.090 294.110 2280.270 ;
        RECT 292.930 2277.490 294.110 2278.670 ;
        RECT 454.930 2261.090 456.110 2262.270 ;
        RECT 454.930 2259.490 456.110 2260.670 ;
        RECT 472.930 2279.090 474.110 2280.270 ;
        RECT 472.930 2277.490 474.110 2278.670 ;
        RECT 634.930 2261.090 636.110 2262.270 ;
        RECT 634.930 2259.490 636.110 2260.670 ;
        RECT 652.930 2279.090 654.110 2280.270 ;
        RECT 652.930 2277.490 654.110 2278.670 ;
        RECT 814.930 2261.090 816.110 2262.270 ;
        RECT 814.930 2259.490 816.110 2260.670 ;
        RECT 832.930 3359.090 834.110 3360.270 ;
        RECT 832.930 3357.490 834.110 3358.670 ;
        RECT 832.930 3179.090 834.110 3180.270 ;
        RECT 832.930 3177.490 834.110 3178.670 ;
        RECT 832.930 2999.090 834.110 3000.270 ;
        RECT 832.930 2997.490 834.110 2998.670 ;
        RECT 832.930 2819.090 834.110 2820.270 ;
        RECT 832.930 2817.490 834.110 2818.670 ;
        RECT 832.930 2639.090 834.110 2640.270 ;
        RECT 832.930 2637.490 834.110 2638.670 ;
        RECT 832.930 2459.090 834.110 2460.270 ;
        RECT 832.930 2457.490 834.110 2458.670 ;
        RECT 832.930 2279.090 834.110 2280.270 ;
        RECT 832.930 2277.490 834.110 2278.670 ;
        RECT 850.930 3377.090 852.110 3378.270 ;
        RECT 850.930 3375.490 852.110 3376.670 ;
        RECT 850.930 3197.090 852.110 3198.270 ;
        RECT 850.930 3195.490 852.110 3196.670 ;
        RECT 850.930 3017.090 852.110 3018.270 ;
        RECT 850.930 3015.490 852.110 3016.670 ;
        RECT 850.930 2837.090 852.110 2838.270 ;
        RECT 850.930 2835.490 852.110 2836.670 ;
        RECT 850.930 2657.090 852.110 2658.270 ;
        RECT 850.930 2655.490 852.110 2656.670 ;
        RECT 850.930 2477.090 852.110 2478.270 ;
        RECT 850.930 2475.490 852.110 2476.670 ;
        RECT 850.930 2297.090 852.110 2298.270 ;
        RECT 850.930 2295.490 852.110 2296.670 ;
        RECT 1048.930 3555.910 1050.110 3557.090 ;
        RECT 1048.930 3554.310 1050.110 3555.490 ;
        RECT 1030.930 3546.510 1032.110 3547.690 ;
        RECT 1030.930 3544.910 1032.110 3546.090 ;
        RECT 1012.930 3537.110 1014.110 3538.290 ;
        RECT 1012.930 3535.510 1014.110 3536.690 ;
        RECT 868.930 3395.090 870.110 3396.270 ;
        RECT 868.930 3393.490 870.110 3394.670 ;
        RECT 868.930 3215.090 870.110 3216.270 ;
        RECT 868.930 3213.490 870.110 3214.670 ;
        RECT 868.930 3035.090 870.110 3036.270 ;
        RECT 868.930 3033.490 870.110 3034.670 ;
        RECT 868.930 2855.090 870.110 2856.270 ;
        RECT 868.930 2853.490 870.110 2854.670 ;
        RECT 994.930 3527.710 996.110 3528.890 ;
        RECT 994.930 3526.110 996.110 3527.290 ;
        RECT 994.930 3341.090 996.110 3342.270 ;
        RECT 994.930 3339.490 996.110 3340.670 ;
        RECT 994.930 3161.090 996.110 3162.270 ;
        RECT 994.930 3159.490 996.110 3160.670 ;
        RECT 994.930 2981.090 996.110 2982.270 ;
        RECT 994.930 2979.490 996.110 2980.670 ;
        RECT 994.930 2801.090 996.110 2802.270 ;
        RECT 994.930 2799.490 996.110 2800.670 ;
        RECT 1012.930 3359.090 1014.110 3360.270 ;
        RECT 1012.930 3357.490 1014.110 3358.670 ;
        RECT 1012.930 3179.090 1014.110 3180.270 ;
        RECT 1012.930 3177.490 1014.110 3178.670 ;
        RECT 1012.930 2999.090 1014.110 3000.270 ;
        RECT 1012.930 2997.490 1014.110 2998.670 ;
        RECT 1012.930 2819.090 1014.110 2820.270 ;
        RECT 1012.930 2817.490 1014.110 2818.670 ;
        RECT 1030.930 3377.090 1032.110 3378.270 ;
        RECT 1030.930 3375.490 1032.110 3376.670 ;
        RECT 1030.930 3197.090 1032.110 3198.270 ;
        RECT 1030.930 3195.490 1032.110 3196.670 ;
        RECT 1030.930 3017.090 1032.110 3018.270 ;
        RECT 1030.930 3015.490 1032.110 3016.670 ;
        RECT 1030.930 2837.090 1032.110 2838.270 ;
        RECT 1030.930 2835.490 1032.110 2836.670 ;
        RECT 1228.930 3555.910 1230.110 3557.090 ;
        RECT 1228.930 3554.310 1230.110 3555.490 ;
        RECT 1210.930 3546.510 1212.110 3547.690 ;
        RECT 1210.930 3544.910 1212.110 3546.090 ;
        RECT 1192.930 3537.110 1194.110 3538.290 ;
        RECT 1192.930 3535.510 1194.110 3536.690 ;
        RECT 1048.930 3395.090 1050.110 3396.270 ;
        RECT 1048.930 3393.490 1050.110 3394.670 ;
        RECT 1048.930 3215.090 1050.110 3216.270 ;
        RECT 1048.930 3213.490 1050.110 3214.670 ;
        RECT 1048.930 3035.090 1050.110 3036.270 ;
        RECT 1048.930 3033.490 1050.110 3034.670 ;
        RECT 1048.930 2855.090 1050.110 2856.270 ;
        RECT 1048.930 2853.490 1050.110 2854.670 ;
        RECT 1174.930 3527.710 1176.110 3528.890 ;
        RECT 1174.930 3526.110 1176.110 3527.290 ;
        RECT 1174.930 3341.090 1176.110 3342.270 ;
        RECT 1174.930 3339.490 1176.110 3340.670 ;
        RECT 1174.930 3161.090 1176.110 3162.270 ;
        RECT 1174.930 3159.490 1176.110 3160.670 ;
        RECT 1174.930 2981.090 1176.110 2982.270 ;
        RECT 1174.930 2979.490 1176.110 2980.670 ;
        RECT 1174.930 2801.090 1176.110 2802.270 ;
        RECT 1174.930 2799.490 1176.110 2800.670 ;
        RECT 1192.930 3359.090 1194.110 3360.270 ;
        RECT 1192.930 3357.490 1194.110 3358.670 ;
        RECT 1192.930 3179.090 1194.110 3180.270 ;
        RECT 1192.930 3177.490 1194.110 3178.670 ;
        RECT 1192.930 2999.090 1194.110 3000.270 ;
        RECT 1192.930 2997.490 1194.110 2998.670 ;
        RECT 1192.930 2819.090 1194.110 2820.270 ;
        RECT 1192.930 2817.490 1194.110 2818.670 ;
        RECT 1210.930 3377.090 1212.110 3378.270 ;
        RECT 1210.930 3375.490 1212.110 3376.670 ;
        RECT 1210.930 3197.090 1212.110 3198.270 ;
        RECT 1210.930 3195.490 1212.110 3196.670 ;
        RECT 1210.930 3017.090 1212.110 3018.270 ;
        RECT 1210.930 3015.490 1212.110 3016.670 ;
        RECT 1210.930 2837.090 1212.110 2838.270 ;
        RECT 1210.930 2835.490 1212.110 2836.670 ;
        RECT 1408.930 3555.910 1410.110 3557.090 ;
        RECT 1408.930 3554.310 1410.110 3555.490 ;
        RECT 1390.930 3546.510 1392.110 3547.690 ;
        RECT 1390.930 3544.910 1392.110 3546.090 ;
        RECT 1372.930 3537.110 1374.110 3538.290 ;
        RECT 1372.930 3535.510 1374.110 3536.690 ;
        RECT 1228.930 3395.090 1230.110 3396.270 ;
        RECT 1228.930 3393.490 1230.110 3394.670 ;
        RECT 1228.930 3215.090 1230.110 3216.270 ;
        RECT 1228.930 3213.490 1230.110 3214.670 ;
        RECT 1228.930 3035.090 1230.110 3036.270 ;
        RECT 1228.930 3033.490 1230.110 3034.670 ;
        RECT 1228.930 2855.090 1230.110 2856.270 ;
        RECT 1228.930 2853.490 1230.110 2854.670 ;
        RECT 1354.930 3527.710 1356.110 3528.890 ;
        RECT 1354.930 3526.110 1356.110 3527.290 ;
        RECT 1354.930 3341.090 1356.110 3342.270 ;
        RECT 1354.930 3339.490 1356.110 3340.670 ;
        RECT 1354.930 3161.090 1356.110 3162.270 ;
        RECT 1354.930 3159.490 1356.110 3160.670 ;
        RECT 1354.930 2981.090 1356.110 2982.270 ;
        RECT 1354.930 2979.490 1356.110 2980.670 ;
        RECT 1354.930 2801.090 1356.110 2802.270 ;
        RECT 1354.930 2799.490 1356.110 2800.670 ;
        RECT 868.930 2675.090 870.110 2676.270 ;
        RECT 868.930 2673.490 870.110 2674.670 ;
        RECT 868.930 2495.090 870.110 2496.270 ;
        RECT 868.930 2493.490 870.110 2494.670 ;
        RECT 868.930 2315.090 870.110 2316.270 ;
        RECT 868.930 2313.490 870.110 2314.670 ;
        RECT 1334.910 2675.090 1336.090 2676.270 ;
        RECT 1334.910 2673.490 1336.090 2674.670 ;
        RECT 1334.910 2657.090 1336.090 2658.270 ;
        RECT 1334.910 2655.490 1336.090 2656.670 ;
        RECT 1334.910 2639.090 1336.090 2640.270 ;
        RECT 1334.910 2637.490 1336.090 2638.670 ;
        RECT 1334.910 2621.090 1336.090 2622.270 ;
        RECT 1334.910 2619.490 1336.090 2620.670 ;
        RECT 1334.910 2495.090 1336.090 2496.270 ;
        RECT 1334.910 2493.490 1336.090 2494.670 ;
        RECT 1334.910 2477.090 1336.090 2478.270 ;
        RECT 1334.910 2475.490 1336.090 2476.670 ;
        RECT 1334.910 2459.090 1336.090 2460.270 ;
        RECT 1334.910 2457.490 1336.090 2458.670 ;
        RECT 1334.910 2441.090 1336.090 2442.270 ;
        RECT 1334.910 2439.490 1336.090 2440.670 ;
        RECT 1334.910 2315.090 1336.090 2316.270 ;
        RECT 1334.910 2313.490 1336.090 2314.670 ;
        RECT 1354.930 2621.090 1356.110 2622.270 ;
        RECT 1354.930 2619.490 1356.110 2620.670 ;
        RECT 1354.930 2441.090 1356.110 2442.270 ;
        RECT 1354.930 2439.490 1356.110 2440.670 ;
        RECT 994.930 2261.090 996.110 2262.270 ;
        RECT 994.930 2259.490 996.110 2260.670 ;
        RECT 1012.930 2279.090 1014.110 2280.270 ;
        RECT 1012.930 2277.490 1014.110 2278.670 ;
        RECT 1174.930 2261.090 1176.110 2262.270 ;
        RECT 1174.930 2259.490 1176.110 2260.670 ;
        RECT 1192.930 2279.090 1194.110 2280.270 ;
        RECT 1192.930 2277.490 1194.110 2278.670 ;
        RECT 1354.930 2261.090 1356.110 2262.270 ;
        RECT 1354.930 2259.490 1356.110 2260.670 ;
        RECT 1372.930 3359.090 1374.110 3360.270 ;
        RECT 1372.930 3357.490 1374.110 3358.670 ;
        RECT 1372.930 3179.090 1374.110 3180.270 ;
        RECT 1372.930 3177.490 1374.110 3178.670 ;
        RECT 1372.930 2999.090 1374.110 3000.270 ;
        RECT 1372.930 2997.490 1374.110 2998.670 ;
        RECT 1372.930 2819.090 1374.110 2820.270 ;
        RECT 1372.930 2817.490 1374.110 2818.670 ;
        RECT 1372.930 2639.090 1374.110 2640.270 ;
        RECT 1372.930 2637.490 1374.110 2638.670 ;
        RECT 1372.930 2459.090 1374.110 2460.270 ;
        RECT 1372.930 2457.490 1374.110 2458.670 ;
        RECT 1372.930 2279.090 1374.110 2280.270 ;
        RECT 1372.930 2277.490 1374.110 2278.670 ;
        RECT 1390.930 3377.090 1392.110 3378.270 ;
        RECT 1390.930 3375.490 1392.110 3376.670 ;
        RECT 1390.930 3197.090 1392.110 3198.270 ;
        RECT 1390.930 3195.490 1392.110 3196.670 ;
        RECT 1390.930 3017.090 1392.110 3018.270 ;
        RECT 1390.930 3015.490 1392.110 3016.670 ;
        RECT 1390.930 2837.090 1392.110 2838.270 ;
        RECT 1390.930 2835.490 1392.110 2836.670 ;
        RECT 1390.930 2657.090 1392.110 2658.270 ;
        RECT 1390.930 2655.490 1392.110 2656.670 ;
        RECT 1390.930 2477.090 1392.110 2478.270 ;
        RECT 1390.930 2475.490 1392.110 2476.670 ;
        RECT 1390.930 2297.090 1392.110 2298.270 ;
        RECT 1390.930 2295.490 1392.110 2296.670 ;
        RECT 1588.930 3555.910 1590.110 3557.090 ;
        RECT 1588.930 3554.310 1590.110 3555.490 ;
        RECT 1570.930 3546.510 1572.110 3547.690 ;
        RECT 1570.930 3544.910 1572.110 3546.090 ;
        RECT 1552.930 3537.110 1554.110 3538.290 ;
        RECT 1552.930 3535.510 1554.110 3536.690 ;
        RECT 1408.930 3395.090 1410.110 3396.270 ;
        RECT 1408.930 3393.490 1410.110 3394.670 ;
        RECT 1408.930 3215.090 1410.110 3216.270 ;
        RECT 1408.930 3213.490 1410.110 3214.670 ;
        RECT 1408.930 3035.090 1410.110 3036.270 ;
        RECT 1408.930 3033.490 1410.110 3034.670 ;
        RECT 1408.930 2855.090 1410.110 2856.270 ;
        RECT 1408.930 2853.490 1410.110 2854.670 ;
        RECT 1534.930 3527.710 1536.110 3528.890 ;
        RECT 1534.930 3526.110 1536.110 3527.290 ;
        RECT 1534.930 3341.090 1536.110 3342.270 ;
        RECT 1534.930 3339.490 1536.110 3340.670 ;
        RECT 1534.930 3161.090 1536.110 3162.270 ;
        RECT 1534.930 3159.490 1536.110 3160.670 ;
        RECT 1534.930 2981.090 1536.110 2982.270 ;
        RECT 1534.930 2979.490 1536.110 2980.670 ;
        RECT 1534.930 2801.090 1536.110 2802.270 ;
        RECT 1534.930 2799.490 1536.110 2800.670 ;
        RECT 1552.930 3359.090 1554.110 3360.270 ;
        RECT 1552.930 3357.490 1554.110 3358.670 ;
        RECT 1552.930 3179.090 1554.110 3180.270 ;
        RECT 1552.930 3177.490 1554.110 3178.670 ;
        RECT 1552.930 2999.090 1554.110 3000.270 ;
        RECT 1552.930 2997.490 1554.110 2998.670 ;
        RECT 1552.930 2819.090 1554.110 2820.270 ;
        RECT 1552.930 2817.490 1554.110 2818.670 ;
        RECT 1570.930 3377.090 1572.110 3378.270 ;
        RECT 1570.930 3375.490 1572.110 3376.670 ;
        RECT 1570.930 3197.090 1572.110 3198.270 ;
        RECT 1570.930 3195.490 1572.110 3196.670 ;
        RECT 1570.930 3017.090 1572.110 3018.270 ;
        RECT 1570.930 3015.490 1572.110 3016.670 ;
        RECT 1570.930 2837.090 1572.110 2838.270 ;
        RECT 1570.930 2835.490 1572.110 2836.670 ;
        RECT 1768.930 3555.910 1770.110 3557.090 ;
        RECT 1768.930 3554.310 1770.110 3555.490 ;
        RECT 1750.930 3546.510 1752.110 3547.690 ;
        RECT 1750.930 3544.910 1752.110 3546.090 ;
        RECT 1732.930 3537.110 1734.110 3538.290 ;
        RECT 1732.930 3535.510 1734.110 3536.690 ;
        RECT 1588.930 3395.090 1590.110 3396.270 ;
        RECT 1588.930 3393.490 1590.110 3394.670 ;
        RECT 1588.930 3215.090 1590.110 3216.270 ;
        RECT 1588.930 3213.490 1590.110 3214.670 ;
        RECT 1588.930 3035.090 1590.110 3036.270 ;
        RECT 1588.930 3033.490 1590.110 3034.670 ;
        RECT 1588.930 2855.090 1590.110 2856.270 ;
        RECT 1588.930 2853.490 1590.110 2854.670 ;
        RECT 1714.930 3527.710 1716.110 3528.890 ;
        RECT 1714.930 3526.110 1716.110 3527.290 ;
        RECT 1714.930 3341.090 1716.110 3342.270 ;
        RECT 1714.930 3339.490 1716.110 3340.670 ;
        RECT 1714.930 3161.090 1716.110 3162.270 ;
        RECT 1714.930 3159.490 1716.110 3160.670 ;
        RECT 1714.930 2981.090 1716.110 2982.270 ;
        RECT 1714.930 2979.490 1716.110 2980.670 ;
        RECT 1714.930 2801.090 1716.110 2802.270 ;
        RECT 1714.930 2799.490 1716.110 2800.670 ;
        RECT 1732.930 3359.090 1734.110 3360.270 ;
        RECT 1732.930 3357.490 1734.110 3358.670 ;
        RECT 1732.930 3179.090 1734.110 3180.270 ;
        RECT 1732.930 3177.490 1734.110 3178.670 ;
        RECT 1732.930 2999.090 1734.110 3000.270 ;
        RECT 1732.930 2997.490 1734.110 2998.670 ;
        RECT 1732.930 2819.090 1734.110 2820.270 ;
        RECT 1732.930 2817.490 1734.110 2818.670 ;
        RECT 1750.930 3377.090 1752.110 3378.270 ;
        RECT 1750.930 3375.490 1752.110 3376.670 ;
        RECT 1750.930 3197.090 1752.110 3198.270 ;
        RECT 1750.930 3195.490 1752.110 3196.670 ;
        RECT 1750.930 3017.090 1752.110 3018.270 ;
        RECT 1750.930 3015.490 1752.110 3016.670 ;
        RECT 1750.930 2837.090 1752.110 2838.270 ;
        RECT 1750.930 2835.490 1752.110 2836.670 ;
        RECT 1948.930 3555.910 1950.110 3557.090 ;
        RECT 1948.930 3554.310 1950.110 3555.490 ;
        RECT 1930.930 3546.510 1932.110 3547.690 ;
        RECT 1930.930 3544.910 1932.110 3546.090 ;
        RECT 1912.930 3537.110 1914.110 3538.290 ;
        RECT 1912.930 3535.510 1914.110 3536.690 ;
        RECT 1768.930 3395.090 1770.110 3396.270 ;
        RECT 1768.930 3393.490 1770.110 3394.670 ;
        RECT 1768.930 3215.090 1770.110 3216.270 ;
        RECT 1768.930 3213.490 1770.110 3214.670 ;
        RECT 1768.930 3035.090 1770.110 3036.270 ;
        RECT 1768.930 3033.490 1770.110 3034.670 ;
        RECT 1768.930 2855.090 1770.110 2856.270 ;
        RECT 1768.930 2853.490 1770.110 2854.670 ;
        RECT 1894.930 3527.710 1896.110 3528.890 ;
        RECT 1894.930 3526.110 1896.110 3527.290 ;
        RECT 1894.930 3341.090 1896.110 3342.270 ;
        RECT 1894.930 3339.490 1896.110 3340.670 ;
        RECT 1894.930 3161.090 1896.110 3162.270 ;
        RECT 1894.930 3159.490 1896.110 3160.670 ;
        RECT 1894.930 2981.090 1896.110 2982.270 ;
        RECT 1894.930 2979.490 1896.110 2980.670 ;
        RECT 1894.930 2801.090 1896.110 2802.270 ;
        RECT 1894.930 2799.490 1896.110 2800.670 ;
        RECT 1912.930 3359.090 1914.110 3360.270 ;
        RECT 1912.930 3357.490 1914.110 3358.670 ;
        RECT 1912.930 3179.090 1914.110 3180.270 ;
        RECT 1912.930 3177.490 1914.110 3178.670 ;
        RECT 1912.930 2999.090 1914.110 3000.270 ;
        RECT 1912.930 2997.490 1914.110 2998.670 ;
        RECT 1912.930 2819.090 1914.110 2820.270 ;
        RECT 1912.930 2817.490 1914.110 2818.670 ;
        RECT 1930.930 3377.090 1932.110 3378.270 ;
        RECT 1930.930 3375.490 1932.110 3376.670 ;
        RECT 1930.930 3197.090 1932.110 3198.270 ;
        RECT 1930.930 3195.490 1932.110 3196.670 ;
        RECT 1930.930 3017.090 1932.110 3018.270 ;
        RECT 1930.930 3015.490 1932.110 3016.670 ;
        RECT 1930.930 2837.090 1932.110 2838.270 ;
        RECT 1930.930 2835.490 1932.110 2836.670 ;
        RECT 2128.930 3555.910 2130.110 3557.090 ;
        RECT 2128.930 3554.310 2130.110 3555.490 ;
        RECT 2110.930 3546.510 2112.110 3547.690 ;
        RECT 2110.930 3544.910 2112.110 3546.090 ;
        RECT 2092.930 3537.110 2094.110 3538.290 ;
        RECT 2092.930 3535.510 2094.110 3536.690 ;
        RECT 1948.930 3395.090 1950.110 3396.270 ;
        RECT 1948.930 3393.490 1950.110 3394.670 ;
        RECT 1948.930 3215.090 1950.110 3216.270 ;
        RECT 1948.930 3213.490 1950.110 3214.670 ;
        RECT 1948.930 3035.090 1950.110 3036.270 ;
        RECT 1948.930 3033.490 1950.110 3034.670 ;
        RECT 1948.930 2855.090 1950.110 2856.270 ;
        RECT 1948.930 2853.490 1950.110 2854.670 ;
        RECT 2074.930 3527.710 2076.110 3528.890 ;
        RECT 2074.930 3526.110 2076.110 3527.290 ;
        RECT 2074.930 3341.090 2076.110 3342.270 ;
        RECT 2074.930 3339.490 2076.110 3340.670 ;
        RECT 2074.930 3161.090 2076.110 3162.270 ;
        RECT 2074.930 3159.490 2076.110 3160.670 ;
        RECT 2074.930 2981.090 2076.110 2982.270 ;
        RECT 2074.930 2979.490 2076.110 2980.670 ;
        RECT 2074.930 2801.090 2076.110 2802.270 ;
        RECT 2074.930 2799.490 2076.110 2800.670 ;
        RECT 1408.930 2675.090 1410.110 2676.270 ;
        RECT 1408.930 2673.490 1410.110 2674.670 ;
        RECT 1408.930 2495.090 1410.110 2496.270 ;
        RECT 1408.930 2493.490 1410.110 2494.670 ;
        RECT 1408.930 2315.090 1410.110 2316.270 ;
        RECT 1408.930 2313.490 1410.110 2314.670 ;
        RECT 1934.910 2675.090 1936.090 2676.270 ;
        RECT 1934.910 2673.490 1936.090 2674.670 ;
        RECT 1934.910 2657.090 1936.090 2658.270 ;
        RECT 1934.910 2655.490 1936.090 2656.670 ;
        RECT 1934.910 2639.090 1936.090 2640.270 ;
        RECT 1934.910 2637.490 1936.090 2638.670 ;
        RECT 1934.910 2621.090 1936.090 2622.270 ;
        RECT 1934.910 2619.490 1936.090 2620.670 ;
        RECT 1934.910 2495.090 1936.090 2496.270 ;
        RECT 1934.910 2493.490 1936.090 2494.670 ;
        RECT 1934.910 2477.090 1936.090 2478.270 ;
        RECT 1934.910 2475.490 1936.090 2476.670 ;
        RECT 1934.910 2459.090 1936.090 2460.270 ;
        RECT 1934.910 2457.490 1936.090 2458.670 ;
        RECT 1934.910 2441.090 1936.090 2442.270 ;
        RECT 1934.910 2439.490 1936.090 2440.670 ;
        RECT 1934.910 2315.090 1936.090 2316.270 ;
        RECT 1934.910 2313.490 1936.090 2314.670 ;
        RECT 2074.930 2621.090 2076.110 2622.270 ;
        RECT 2074.930 2619.490 2076.110 2620.670 ;
        RECT 2074.930 2441.090 2076.110 2442.270 ;
        RECT 2074.930 2439.490 2076.110 2440.670 ;
        RECT 1534.930 2261.090 1536.110 2262.270 ;
        RECT 1534.930 2259.490 1536.110 2260.670 ;
        RECT 274.930 2081.090 276.110 2082.270 ;
        RECT 274.930 2079.490 276.110 2080.670 ;
        RECT 274.930 1901.090 276.110 1902.270 ;
        RECT 274.930 1899.490 276.110 1900.670 ;
        RECT 274.930 1721.090 276.110 1722.270 ;
        RECT 274.930 1719.490 276.110 1720.670 ;
        RECT 274.930 1541.090 276.110 1542.270 ;
        RECT 274.930 1539.490 276.110 1540.670 ;
        RECT 274.930 1361.090 276.110 1362.270 ;
        RECT 274.930 1359.490 276.110 1360.670 ;
        RECT 274.930 1181.090 276.110 1182.270 ;
        RECT 274.930 1179.490 276.110 1180.670 ;
        RECT 398.050 2135.090 399.230 2136.270 ;
        RECT 398.050 2133.490 399.230 2134.670 ;
        RECT 398.050 2117.090 399.230 2118.270 ;
        RECT 398.050 2115.490 399.230 2116.670 ;
        RECT 398.050 2099.090 399.230 2100.270 ;
        RECT 398.050 2097.490 399.230 2098.670 ;
        RECT 398.050 2081.090 399.230 2082.270 ;
        RECT 398.050 2079.490 399.230 2080.670 ;
        RECT 398.050 1955.090 399.230 1956.270 ;
        RECT 398.050 1953.490 399.230 1954.670 ;
        RECT 398.050 1937.090 399.230 1938.270 ;
        RECT 398.050 1935.490 399.230 1936.670 ;
        RECT 398.050 1919.090 399.230 1920.270 ;
        RECT 398.050 1917.490 399.230 1918.670 ;
        RECT 398.050 1901.090 399.230 1902.270 ;
        RECT 398.050 1899.490 399.230 1900.670 ;
        RECT 398.050 1775.090 399.230 1776.270 ;
        RECT 398.050 1773.490 399.230 1774.670 ;
        RECT 398.050 1757.090 399.230 1758.270 ;
        RECT 398.050 1755.490 399.230 1756.670 ;
        RECT 398.050 1739.090 399.230 1740.270 ;
        RECT 398.050 1737.490 399.230 1738.670 ;
        RECT 398.050 1721.090 399.230 1722.270 ;
        RECT 398.050 1719.490 399.230 1720.670 ;
        RECT 398.050 1595.090 399.230 1596.270 ;
        RECT 398.050 1593.490 399.230 1594.670 ;
        RECT 398.050 1577.090 399.230 1578.270 ;
        RECT 398.050 1575.490 399.230 1576.670 ;
        RECT 398.050 1559.090 399.230 1560.270 ;
        RECT 398.050 1557.490 399.230 1558.670 ;
        RECT 398.050 1541.090 399.230 1542.270 ;
        RECT 398.050 1539.490 399.230 1540.670 ;
        RECT 398.050 1415.090 399.230 1416.270 ;
        RECT 398.050 1413.490 399.230 1414.670 ;
        RECT 398.050 1397.090 399.230 1398.270 ;
        RECT 398.050 1395.490 399.230 1396.670 ;
        RECT 398.050 1379.090 399.230 1380.270 ;
        RECT 398.050 1377.490 399.230 1378.670 ;
        RECT 398.050 1361.090 399.230 1362.270 ;
        RECT 398.050 1359.490 399.230 1360.670 ;
        RECT 398.050 1235.090 399.230 1236.270 ;
        RECT 398.050 1233.490 399.230 1234.670 ;
        RECT 398.050 1217.090 399.230 1218.270 ;
        RECT 398.050 1215.490 399.230 1216.670 ;
        RECT 398.050 1199.090 399.230 1200.270 ;
        RECT 398.050 1197.490 399.230 1198.670 ;
        RECT 398.050 1181.090 399.230 1182.270 ;
        RECT 398.050 1179.490 399.230 1180.670 ;
        RECT 398.050 1055.090 399.230 1056.270 ;
        RECT 398.050 1053.490 399.230 1054.670 ;
        RECT 398.050 1037.090 399.230 1038.270 ;
        RECT 398.050 1035.490 399.230 1036.670 ;
        RECT 398.050 1019.090 399.230 1020.270 ;
        RECT 398.050 1017.490 399.230 1018.670 ;
        RECT 1534.930 2081.090 1536.110 2082.270 ;
        RECT 1534.930 2079.490 1536.110 2080.670 ;
        RECT 1534.930 1901.090 1536.110 1902.270 ;
        RECT 1534.930 1899.490 1536.110 1900.670 ;
        RECT 1534.930 1721.090 1536.110 1722.270 ;
        RECT 1534.930 1719.490 1536.110 1720.670 ;
        RECT 1534.930 1541.090 1536.110 1542.270 ;
        RECT 1534.930 1539.490 1536.110 1540.670 ;
        RECT 1534.930 1361.090 1536.110 1362.270 ;
        RECT 1534.930 1359.490 1536.110 1360.670 ;
        RECT 1534.930 1181.090 1536.110 1182.270 ;
        RECT 1534.930 1179.490 1536.110 1180.670 ;
        RECT 274.930 1001.090 276.110 1002.270 ;
        RECT 274.930 999.490 276.110 1000.670 ;
        RECT 1534.930 1001.090 1536.110 1002.270 ;
        RECT 1534.930 999.490 1536.110 1000.670 ;
        RECT 274.930 821.090 276.110 822.270 ;
        RECT 274.930 819.490 276.110 820.670 ;
        RECT 274.930 641.090 276.110 642.270 ;
        RECT 274.930 639.490 276.110 640.670 ;
        RECT 274.930 461.090 276.110 462.270 ;
        RECT 274.930 459.490 276.110 460.670 ;
        RECT 274.930 281.090 276.110 282.270 ;
        RECT 274.930 279.490 276.110 280.670 ;
        RECT 274.930 101.090 276.110 102.270 ;
        RECT 274.930 99.490 276.110 100.670 ;
        RECT 274.930 -7.610 276.110 -6.430 ;
        RECT 274.930 -9.210 276.110 -8.030 ;
        RECT 292.930 839.090 294.110 840.270 ;
        RECT 292.930 837.490 294.110 838.670 ;
        RECT 292.930 659.090 294.110 660.270 ;
        RECT 292.930 657.490 294.110 658.670 ;
        RECT 292.930 479.090 294.110 480.270 ;
        RECT 292.930 477.490 294.110 478.670 ;
        RECT 292.930 299.090 294.110 300.270 ;
        RECT 292.930 297.490 294.110 298.670 ;
        RECT 292.930 119.090 294.110 120.270 ;
        RECT 292.930 117.490 294.110 118.670 ;
        RECT 292.930 -17.010 294.110 -15.830 ;
        RECT 292.930 -18.610 294.110 -17.430 ;
        RECT 310.930 857.090 312.110 858.270 ;
        RECT 310.930 855.490 312.110 856.670 ;
        RECT 310.930 677.090 312.110 678.270 ;
        RECT 310.930 675.490 312.110 676.670 ;
        RECT 310.930 497.090 312.110 498.270 ;
        RECT 310.930 495.490 312.110 496.670 ;
        RECT 310.930 317.090 312.110 318.270 ;
        RECT 310.930 315.490 312.110 316.670 ;
        RECT 310.930 137.090 312.110 138.270 ;
        RECT 310.930 135.490 312.110 136.670 ;
        RECT 310.930 -26.410 312.110 -25.230 ;
        RECT 310.930 -28.010 312.110 -26.830 ;
        RECT 328.930 875.090 330.110 876.270 ;
        RECT 328.930 873.490 330.110 874.670 ;
        RECT 328.930 695.090 330.110 696.270 ;
        RECT 328.930 693.490 330.110 694.670 ;
        RECT 328.930 515.090 330.110 516.270 ;
        RECT 328.930 513.490 330.110 514.670 ;
        RECT 328.930 335.090 330.110 336.270 ;
        RECT 328.930 333.490 330.110 334.670 ;
        RECT 328.930 155.090 330.110 156.270 ;
        RECT 328.930 153.490 330.110 154.670 ;
        RECT 148.930 -35.810 150.110 -34.630 ;
        RECT 148.930 -37.410 150.110 -36.230 ;
        RECT 454.930 821.090 456.110 822.270 ;
        RECT 454.930 819.490 456.110 820.670 ;
        RECT 454.930 641.090 456.110 642.270 ;
        RECT 454.930 639.490 456.110 640.670 ;
        RECT 454.930 461.090 456.110 462.270 ;
        RECT 454.930 459.490 456.110 460.670 ;
        RECT 454.930 281.090 456.110 282.270 ;
        RECT 454.930 279.490 456.110 280.670 ;
        RECT 454.930 101.090 456.110 102.270 ;
        RECT 454.930 99.490 456.110 100.670 ;
        RECT 454.930 -7.610 456.110 -6.430 ;
        RECT 454.930 -9.210 456.110 -8.030 ;
        RECT 472.930 839.090 474.110 840.270 ;
        RECT 472.930 837.490 474.110 838.670 ;
        RECT 472.930 659.090 474.110 660.270 ;
        RECT 472.930 657.490 474.110 658.670 ;
        RECT 472.930 479.090 474.110 480.270 ;
        RECT 472.930 477.490 474.110 478.670 ;
        RECT 472.930 299.090 474.110 300.270 ;
        RECT 472.930 297.490 474.110 298.670 ;
        RECT 472.930 119.090 474.110 120.270 ;
        RECT 472.930 117.490 474.110 118.670 ;
        RECT 472.930 -17.010 474.110 -15.830 ;
        RECT 472.930 -18.610 474.110 -17.430 ;
        RECT 490.930 857.090 492.110 858.270 ;
        RECT 490.930 855.490 492.110 856.670 ;
        RECT 490.930 677.090 492.110 678.270 ;
        RECT 490.930 675.490 492.110 676.670 ;
        RECT 490.930 497.090 492.110 498.270 ;
        RECT 490.930 495.490 492.110 496.670 ;
        RECT 490.930 317.090 492.110 318.270 ;
        RECT 490.930 315.490 492.110 316.670 ;
        RECT 490.930 137.090 492.110 138.270 ;
        RECT 490.930 135.490 492.110 136.670 ;
        RECT 490.930 -26.410 492.110 -25.230 ;
        RECT 490.930 -28.010 492.110 -26.830 ;
        RECT 508.930 875.090 510.110 876.270 ;
        RECT 508.930 873.490 510.110 874.670 ;
        RECT 508.930 695.090 510.110 696.270 ;
        RECT 508.930 693.490 510.110 694.670 ;
        RECT 508.930 515.090 510.110 516.270 ;
        RECT 508.930 513.490 510.110 514.670 ;
        RECT 508.930 335.090 510.110 336.270 ;
        RECT 508.930 333.490 510.110 334.670 ;
        RECT 508.930 155.090 510.110 156.270 ;
        RECT 508.930 153.490 510.110 154.670 ;
        RECT 328.930 -35.810 330.110 -34.630 ;
        RECT 328.930 -37.410 330.110 -36.230 ;
        RECT 634.930 821.090 636.110 822.270 ;
        RECT 634.930 819.490 636.110 820.670 ;
        RECT 634.930 641.090 636.110 642.270 ;
        RECT 634.930 639.490 636.110 640.670 ;
        RECT 634.930 461.090 636.110 462.270 ;
        RECT 634.930 459.490 636.110 460.670 ;
        RECT 634.930 281.090 636.110 282.270 ;
        RECT 634.930 279.490 636.110 280.670 ;
        RECT 634.930 101.090 636.110 102.270 ;
        RECT 634.930 99.490 636.110 100.670 ;
        RECT 634.930 -7.610 636.110 -6.430 ;
        RECT 634.930 -9.210 636.110 -8.030 ;
        RECT 652.930 839.090 654.110 840.270 ;
        RECT 652.930 837.490 654.110 838.670 ;
        RECT 652.930 659.090 654.110 660.270 ;
        RECT 652.930 657.490 654.110 658.670 ;
        RECT 652.930 479.090 654.110 480.270 ;
        RECT 652.930 477.490 654.110 478.670 ;
        RECT 652.930 299.090 654.110 300.270 ;
        RECT 652.930 297.490 654.110 298.670 ;
        RECT 652.930 119.090 654.110 120.270 ;
        RECT 652.930 117.490 654.110 118.670 ;
        RECT 652.930 -17.010 654.110 -15.830 ;
        RECT 652.930 -18.610 654.110 -17.430 ;
        RECT 670.930 857.090 672.110 858.270 ;
        RECT 670.930 855.490 672.110 856.670 ;
        RECT 670.930 677.090 672.110 678.270 ;
        RECT 670.930 675.490 672.110 676.670 ;
        RECT 670.930 497.090 672.110 498.270 ;
        RECT 670.930 495.490 672.110 496.670 ;
        RECT 670.930 317.090 672.110 318.270 ;
        RECT 670.930 315.490 672.110 316.670 ;
        RECT 670.930 137.090 672.110 138.270 ;
        RECT 670.930 135.490 672.110 136.670 ;
        RECT 670.930 -26.410 672.110 -25.230 ;
        RECT 670.930 -28.010 672.110 -26.830 ;
        RECT 688.930 875.090 690.110 876.270 ;
        RECT 688.930 873.490 690.110 874.670 ;
        RECT 688.930 695.090 690.110 696.270 ;
        RECT 688.930 693.490 690.110 694.670 ;
        RECT 688.930 515.090 690.110 516.270 ;
        RECT 688.930 513.490 690.110 514.670 ;
        RECT 688.930 335.090 690.110 336.270 ;
        RECT 688.930 333.490 690.110 334.670 ;
        RECT 688.930 155.090 690.110 156.270 ;
        RECT 688.930 153.490 690.110 154.670 ;
        RECT 508.930 -35.810 510.110 -34.630 ;
        RECT 508.930 -37.410 510.110 -36.230 ;
        RECT 814.930 821.090 816.110 822.270 ;
        RECT 814.930 819.490 816.110 820.670 ;
        RECT 814.930 641.090 816.110 642.270 ;
        RECT 814.930 639.490 816.110 640.670 ;
        RECT 814.930 461.090 816.110 462.270 ;
        RECT 814.930 459.490 816.110 460.670 ;
        RECT 814.930 281.090 816.110 282.270 ;
        RECT 814.930 279.490 816.110 280.670 ;
        RECT 814.930 101.090 816.110 102.270 ;
        RECT 814.930 99.490 816.110 100.670 ;
        RECT 814.930 -7.610 816.110 -6.430 ;
        RECT 814.930 -9.210 816.110 -8.030 ;
        RECT 832.930 839.090 834.110 840.270 ;
        RECT 832.930 837.490 834.110 838.670 ;
        RECT 832.930 659.090 834.110 660.270 ;
        RECT 832.930 657.490 834.110 658.670 ;
        RECT 832.930 479.090 834.110 480.270 ;
        RECT 832.930 477.490 834.110 478.670 ;
        RECT 832.930 299.090 834.110 300.270 ;
        RECT 832.930 297.490 834.110 298.670 ;
        RECT 832.930 119.090 834.110 120.270 ;
        RECT 832.930 117.490 834.110 118.670 ;
        RECT 832.930 -17.010 834.110 -15.830 ;
        RECT 832.930 -18.610 834.110 -17.430 ;
        RECT 850.930 857.090 852.110 858.270 ;
        RECT 850.930 855.490 852.110 856.670 ;
        RECT 850.930 677.090 852.110 678.270 ;
        RECT 850.930 675.490 852.110 676.670 ;
        RECT 850.930 497.090 852.110 498.270 ;
        RECT 850.930 495.490 852.110 496.670 ;
        RECT 850.930 317.090 852.110 318.270 ;
        RECT 850.930 315.490 852.110 316.670 ;
        RECT 850.930 137.090 852.110 138.270 ;
        RECT 850.930 135.490 852.110 136.670 ;
        RECT 850.930 -26.410 852.110 -25.230 ;
        RECT 850.930 -28.010 852.110 -26.830 ;
        RECT 868.930 875.090 870.110 876.270 ;
        RECT 868.930 873.490 870.110 874.670 ;
        RECT 868.930 695.090 870.110 696.270 ;
        RECT 868.930 693.490 870.110 694.670 ;
        RECT 868.930 515.090 870.110 516.270 ;
        RECT 868.930 513.490 870.110 514.670 ;
        RECT 868.930 335.090 870.110 336.270 ;
        RECT 868.930 333.490 870.110 334.670 ;
        RECT 868.930 155.090 870.110 156.270 ;
        RECT 868.930 153.490 870.110 154.670 ;
        RECT 688.930 -35.810 690.110 -34.630 ;
        RECT 688.930 -37.410 690.110 -36.230 ;
        RECT 994.930 821.090 996.110 822.270 ;
        RECT 994.930 819.490 996.110 820.670 ;
        RECT 994.930 641.090 996.110 642.270 ;
        RECT 994.930 639.490 996.110 640.670 ;
        RECT 994.930 461.090 996.110 462.270 ;
        RECT 994.930 459.490 996.110 460.670 ;
        RECT 994.930 281.090 996.110 282.270 ;
        RECT 994.930 279.490 996.110 280.670 ;
        RECT 994.930 101.090 996.110 102.270 ;
        RECT 994.930 99.490 996.110 100.670 ;
        RECT 994.930 -7.610 996.110 -6.430 ;
        RECT 994.930 -9.210 996.110 -8.030 ;
        RECT 1012.930 839.090 1014.110 840.270 ;
        RECT 1012.930 837.490 1014.110 838.670 ;
        RECT 1012.930 659.090 1014.110 660.270 ;
        RECT 1012.930 657.490 1014.110 658.670 ;
        RECT 1012.930 479.090 1014.110 480.270 ;
        RECT 1012.930 477.490 1014.110 478.670 ;
        RECT 1012.930 299.090 1014.110 300.270 ;
        RECT 1012.930 297.490 1014.110 298.670 ;
        RECT 1012.930 119.090 1014.110 120.270 ;
        RECT 1012.930 117.490 1014.110 118.670 ;
        RECT 1012.930 -17.010 1014.110 -15.830 ;
        RECT 1012.930 -18.610 1014.110 -17.430 ;
        RECT 1030.930 857.090 1032.110 858.270 ;
        RECT 1030.930 855.490 1032.110 856.670 ;
        RECT 1030.930 677.090 1032.110 678.270 ;
        RECT 1030.930 675.490 1032.110 676.670 ;
        RECT 1030.930 497.090 1032.110 498.270 ;
        RECT 1030.930 495.490 1032.110 496.670 ;
        RECT 1030.930 317.090 1032.110 318.270 ;
        RECT 1030.930 315.490 1032.110 316.670 ;
        RECT 1030.930 137.090 1032.110 138.270 ;
        RECT 1030.930 135.490 1032.110 136.670 ;
        RECT 1030.930 -26.410 1032.110 -25.230 ;
        RECT 1030.930 -28.010 1032.110 -26.830 ;
        RECT 1048.930 875.090 1050.110 876.270 ;
        RECT 1048.930 873.490 1050.110 874.670 ;
        RECT 1048.930 695.090 1050.110 696.270 ;
        RECT 1048.930 693.490 1050.110 694.670 ;
        RECT 1048.930 515.090 1050.110 516.270 ;
        RECT 1048.930 513.490 1050.110 514.670 ;
        RECT 1048.930 335.090 1050.110 336.270 ;
        RECT 1048.930 333.490 1050.110 334.670 ;
        RECT 1048.930 155.090 1050.110 156.270 ;
        RECT 1048.930 153.490 1050.110 154.670 ;
        RECT 868.930 -35.810 870.110 -34.630 ;
        RECT 868.930 -37.410 870.110 -36.230 ;
        RECT 1174.930 821.090 1176.110 822.270 ;
        RECT 1174.930 819.490 1176.110 820.670 ;
        RECT 1174.930 641.090 1176.110 642.270 ;
        RECT 1174.930 639.490 1176.110 640.670 ;
        RECT 1174.930 461.090 1176.110 462.270 ;
        RECT 1174.930 459.490 1176.110 460.670 ;
        RECT 1174.930 281.090 1176.110 282.270 ;
        RECT 1174.930 279.490 1176.110 280.670 ;
        RECT 1174.930 101.090 1176.110 102.270 ;
        RECT 1174.930 99.490 1176.110 100.670 ;
        RECT 1174.930 -7.610 1176.110 -6.430 ;
        RECT 1174.930 -9.210 1176.110 -8.030 ;
        RECT 1192.930 839.090 1194.110 840.270 ;
        RECT 1192.930 837.490 1194.110 838.670 ;
        RECT 1192.930 659.090 1194.110 660.270 ;
        RECT 1192.930 657.490 1194.110 658.670 ;
        RECT 1192.930 479.090 1194.110 480.270 ;
        RECT 1192.930 477.490 1194.110 478.670 ;
        RECT 1192.930 299.090 1194.110 300.270 ;
        RECT 1192.930 297.490 1194.110 298.670 ;
        RECT 1192.930 119.090 1194.110 120.270 ;
        RECT 1192.930 117.490 1194.110 118.670 ;
        RECT 1192.930 -17.010 1194.110 -15.830 ;
        RECT 1192.930 -18.610 1194.110 -17.430 ;
        RECT 1210.930 857.090 1212.110 858.270 ;
        RECT 1210.930 855.490 1212.110 856.670 ;
        RECT 1210.930 677.090 1212.110 678.270 ;
        RECT 1210.930 675.490 1212.110 676.670 ;
        RECT 1210.930 497.090 1212.110 498.270 ;
        RECT 1210.930 495.490 1212.110 496.670 ;
        RECT 1210.930 317.090 1212.110 318.270 ;
        RECT 1210.930 315.490 1212.110 316.670 ;
        RECT 1210.930 137.090 1212.110 138.270 ;
        RECT 1210.930 135.490 1212.110 136.670 ;
        RECT 1210.930 -26.410 1212.110 -25.230 ;
        RECT 1210.930 -28.010 1212.110 -26.830 ;
        RECT 1228.930 875.090 1230.110 876.270 ;
        RECT 1228.930 873.490 1230.110 874.670 ;
        RECT 1228.930 695.090 1230.110 696.270 ;
        RECT 1228.930 693.490 1230.110 694.670 ;
        RECT 1228.930 515.090 1230.110 516.270 ;
        RECT 1228.930 513.490 1230.110 514.670 ;
        RECT 1228.930 335.090 1230.110 336.270 ;
        RECT 1228.930 333.490 1230.110 334.670 ;
        RECT 1228.930 155.090 1230.110 156.270 ;
        RECT 1228.930 153.490 1230.110 154.670 ;
        RECT 1048.930 -35.810 1050.110 -34.630 ;
        RECT 1048.930 -37.410 1050.110 -36.230 ;
        RECT 1354.930 821.090 1356.110 822.270 ;
        RECT 1354.930 819.490 1356.110 820.670 ;
        RECT 1354.930 641.090 1356.110 642.270 ;
        RECT 1354.930 639.490 1356.110 640.670 ;
        RECT 1354.930 461.090 1356.110 462.270 ;
        RECT 1354.930 459.490 1356.110 460.670 ;
        RECT 1354.930 281.090 1356.110 282.270 ;
        RECT 1354.930 279.490 1356.110 280.670 ;
        RECT 1354.930 101.090 1356.110 102.270 ;
        RECT 1354.930 99.490 1356.110 100.670 ;
        RECT 1354.930 -7.610 1356.110 -6.430 ;
        RECT 1354.930 -9.210 1356.110 -8.030 ;
        RECT 1372.930 839.090 1374.110 840.270 ;
        RECT 1372.930 837.490 1374.110 838.670 ;
        RECT 1372.930 659.090 1374.110 660.270 ;
        RECT 1372.930 657.490 1374.110 658.670 ;
        RECT 1372.930 479.090 1374.110 480.270 ;
        RECT 1372.930 477.490 1374.110 478.670 ;
        RECT 1372.930 299.090 1374.110 300.270 ;
        RECT 1372.930 297.490 1374.110 298.670 ;
        RECT 1372.930 119.090 1374.110 120.270 ;
        RECT 1372.930 117.490 1374.110 118.670 ;
        RECT 1372.930 -17.010 1374.110 -15.830 ;
        RECT 1372.930 -18.610 1374.110 -17.430 ;
        RECT 1390.930 857.090 1392.110 858.270 ;
        RECT 1390.930 855.490 1392.110 856.670 ;
        RECT 1390.930 677.090 1392.110 678.270 ;
        RECT 1390.930 675.490 1392.110 676.670 ;
        RECT 1390.930 497.090 1392.110 498.270 ;
        RECT 1390.930 495.490 1392.110 496.670 ;
        RECT 1390.930 317.090 1392.110 318.270 ;
        RECT 1390.930 315.490 1392.110 316.670 ;
        RECT 1390.930 137.090 1392.110 138.270 ;
        RECT 1390.930 135.490 1392.110 136.670 ;
        RECT 1390.930 -26.410 1392.110 -25.230 ;
        RECT 1390.930 -28.010 1392.110 -26.830 ;
        RECT 1408.930 875.090 1410.110 876.270 ;
        RECT 1408.930 873.490 1410.110 874.670 ;
        RECT 1408.930 695.090 1410.110 696.270 ;
        RECT 1408.930 693.490 1410.110 694.670 ;
        RECT 1408.930 515.090 1410.110 516.270 ;
        RECT 1408.930 513.490 1410.110 514.670 ;
        RECT 1408.930 335.090 1410.110 336.270 ;
        RECT 1408.930 333.490 1410.110 334.670 ;
        RECT 1408.930 155.090 1410.110 156.270 ;
        RECT 1408.930 153.490 1410.110 154.670 ;
        RECT 1228.930 -35.810 1230.110 -34.630 ;
        RECT 1228.930 -37.410 1230.110 -36.230 ;
        RECT 1534.930 821.090 1536.110 822.270 ;
        RECT 1534.930 819.490 1536.110 820.670 ;
        RECT 1534.930 641.090 1536.110 642.270 ;
        RECT 1534.930 639.490 1536.110 640.670 ;
        RECT 1534.930 461.090 1536.110 462.270 ;
        RECT 1534.930 459.490 1536.110 460.670 ;
        RECT 1534.930 281.090 1536.110 282.270 ;
        RECT 1534.930 279.490 1536.110 280.670 ;
        RECT 1534.930 101.090 1536.110 102.270 ;
        RECT 1534.930 99.490 1536.110 100.670 ;
        RECT 1534.930 -7.610 1536.110 -6.430 ;
        RECT 1534.930 -9.210 1536.110 -8.030 ;
        RECT 1552.930 2279.090 1554.110 2280.270 ;
        RECT 1552.930 2277.490 1554.110 2278.670 ;
        RECT 1552.930 2099.090 1554.110 2100.270 ;
        RECT 1552.930 2097.490 1554.110 2098.670 ;
        RECT 1552.930 1919.090 1554.110 1920.270 ;
        RECT 1552.930 1917.490 1554.110 1918.670 ;
        RECT 1552.930 1739.090 1554.110 1740.270 ;
        RECT 1552.930 1737.490 1554.110 1738.670 ;
        RECT 1552.930 1559.090 1554.110 1560.270 ;
        RECT 1552.930 1557.490 1554.110 1558.670 ;
        RECT 1552.930 1379.090 1554.110 1380.270 ;
        RECT 1552.930 1377.490 1554.110 1378.670 ;
        RECT 1552.930 1199.090 1554.110 1200.270 ;
        RECT 1552.930 1197.490 1554.110 1198.670 ;
        RECT 1552.930 1019.090 1554.110 1020.270 ;
        RECT 1552.930 1017.490 1554.110 1018.670 ;
        RECT 1552.930 839.090 1554.110 840.270 ;
        RECT 1552.930 837.490 1554.110 838.670 ;
        RECT 1552.930 659.090 1554.110 660.270 ;
        RECT 1552.930 657.490 1554.110 658.670 ;
        RECT 1552.930 479.090 1554.110 480.270 ;
        RECT 1552.930 477.490 1554.110 478.670 ;
        RECT 1552.930 299.090 1554.110 300.270 ;
        RECT 1552.930 297.490 1554.110 298.670 ;
        RECT 1552.930 119.090 1554.110 120.270 ;
        RECT 1552.930 117.490 1554.110 118.670 ;
        RECT 1552.930 -17.010 1554.110 -15.830 ;
        RECT 1552.930 -18.610 1554.110 -17.430 ;
        RECT 1570.930 2117.090 1572.110 2118.270 ;
        RECT 1570.930 2115.490 1572.110 2116.670 ;
        RECT 1570.930 1937.090 1572.110 1938.270 ;
        RECT 1570.930 1935.490 1572.110 1936.670 ;
        RECT 1570.930 1757.090 1572.110 1758.270 ;
        RECT 1570.930 1755.490 1572.110 1756.670 ;
        RECT 1570.930 1577.090 1572.110 1578.270 ;
        RECT 1570.930 1575.490 1572.110 1576.670 ;
        RECT 1570.930 1397.090 1572.110 1398.270 ;
        RECT 1570.930 1395.490 1572.110 1396.670 ;
        RECT 1570.930 1217.090 1572.110 1218.270 ;
        RECT 1570.930 1215.490 1572.110 1216.670 ;
        RECT 1570.930 1037.090 1572.110 1038.270 ;
        RECT 1570.930 1035.490 1572.110 1036.670 ;
        RECT 1570.930 857.090 1572.110 858.270 ;
        RECT 1570.930 855.490 1572.110 856.670 ;
        RECT 1570.930 677.090 1572.110 678.270 ;
        RECT 1570.930 675.490 1572.110 676.670 ;
        RECT 1570.930 497.090 1572.110 498.270 ;
        RECT 1570.930 495.490 1572.110 496.670 ;
        RECT 1570.930 317.090 1572.110 318.270 ;
        RECT 1570.930 315.490 1572.110 316.670 ;
        RECT 1570.930 137.090 1572.110 138.270 ;
        RECT 1570.930 135.490 1572.110 136.670 ;
        RECT 1570.930 -26.410 1572.110 -25.230 ;
        RECT 1570.930 -28.010 1572.110 -26.830 ;
        RECT 1588.930 2135.090 1590.110 2136.270 ;
        RECT 1588.930 2133.490 1590.110 2134.670 ;
        RECT 1588.930 1955.090 1590.110 1956.270 ;
        RECT 1588.930 1953.490 1590.110 1954.670 ;
        RECT 1588.930 1775.090 1590.110 1776.270 ;
        RECT 1588.930 1773.490 1590.110 1774.670 ;
        RECT 1588.930 1595.090 1590.110 1596.270 ;
        RECT 1588.930 1593.490 1590.110 1594.670 ;
        RECT 1588.930 1415.090 1590.110 1416.270 ;
        RECT 1588.930 1413.490 1590.110 1414.670 ;
        RECT 1588.930 1235.090 1590.110 1236.270 ;
        RECT 1588.930 1233.490 1590.110 1234.670 ;
        RECT 1588.930 1055.090 1590.110 1056.270 ;
        RECT 1588.930 1053.490 1590.110 1054.670 ;
        RECT 1588.930 875.090 1590.110 876.270 ;
        RECT 1588.930 873.490 1590.110 874.670 ;
        RECT 1588.930 695.090 1590.110 696.270 ;
        RECT 1588.930 693.490 1590.110 694.670 ;
        RECT 1588.930 515.090 1590.110 516.270 ;
        RECT 1588.930 513.490 1590.110 514.670 ;
        RECT 1588.930 335.090 1590.110 336.270 ;
        RECT 1588.930 333.490 1590.110 334.670 ;
        RECT 1588.930 155.090 1590.110 156.270 ;
        RECT 1588.930 153.490 1590.110 154.670 ;
        RECT 1408.930 -35.810 1410.110 -34.630 ;
        RECT 1408.930 -37.410 1410.110 -36.230 ;
        RECT 1714.930 2261.090 1716.110 2262.270 ;
        RECT 1714.930 2259.490 1716.110 2260.670 ;
        RECT 1714.930 2081.090 1716.110 2082.270 ;
        RECT 1714.930 2079.490 1716.110 2080.670 ;
        RECT 1714.930 1901.090 1716.110 1902.270 ;
        RECT 1714.930 1899.490 1716.110 1900.670 ;
        RECT 1714.930 1721.090 1716.110 1722.270 ;
        RECT 1714.930 1719.490 1716.110 1720.670 ;
        RECT 1714.930 1541.090 1716.110 1542.270 ;
        RECT 1714.930 1539.490 1716.110 1540.670 ;
        RECT 1714.930 1361.090 1716.110 1362.270 ;
        RECT 1714.930 1359.490 1716.110 1360.670 ;
        RECT 1714.930 1181.090 1716.110 1182.270 ;
        RECT 1714.930 1179.490 1716.110 1180.670 ;
        RECT 1714.930 1001.090 1716.110 1002.270 ;
        RECT 1714.930 999.490 1716.110 1000.670 ;
        RECT 1714.930 821.090 1716.110 822.270 ;
        RECT 1714.930 819.490 1716.110 820.670 ;
        RECT 1714.930 641.090 1716.110 642.270 ;
        RECT 1714.930 639.490 1716.110 640.670 ;
        RECT 1714.930 461.090 1716.110 462.270 ;
        RECT 1714.930 459.490 1716.110 460.670 ;
        RECT 1714.930 281.090 1716.110 282.270 ;
        RECT 1714.930 279.490 1716.110 280.670 ;
        RECT 1714.930 101.090 1716.110 102.270 ;
        RECT 1714.930 99.490 1716.110 100.670 ;
        RECT 1714.930 -7.610 1716.110 -6.430 ;
        RECT 1714.930 -9.210 1716.110 -8.030 ;
        RECT 1732.930 2279.090 1734.110 2280.270 ;
        RECT 1732.930 2277.490 1734.110 2278.670 ;
        RECT 1732.930 2099.090 1734.110 2100.270 ;
        RECT 1732.930 2097.490 1734.110 2098.670 ;
        RECT 1732.930 1919.090 1734.110 1920.270 ;
        RECT 1732.930 1917.490 1734.110 1918.670 ;
        RECT 1732.930 1739.090 1734.110 1740.270 ;
        RECT 1732.930 1737.490 1734.110 1738.670 ;
        RECT 1732.930 1559.090 1734.110 1560.270 ;
        RECT 1732.930 1557.490 1734.110 1558.670 ;
        RECT 1732.930 1379.090 1734.110 1380.270 ;
        RECT 1732.930 1377.490 1734.110 1378.670 ;
        RECT 1732.930 1199.090 1734.110 1200.270 ;
        RECT 1732.930 1197.490 1734.110 1198.670 ;
        RECT 1732.930 1019.090 1734.110 1020.270 ;
        RECT 1732.930 1017.490 1734.110 1018.670 ;
        RECT 1732.930 839.090 1734.110 840.270 ;
        RECT 1732.930 837.490 1734.110 838.670 ;
        RECT 1732.930 659.090 1734.110 660.270 ;
        RECT 1732.930 657.490 1734.110 658.670 ;
        RECT 1732.930 479.090 1734.110 480.270 ;
        RECT 1732.930 477.490 1734.110 478.670 ;
        RECT 1732.930 299.090 1734.110 300.270 ;
        RECT 1732.930 297.490 1734.110 298.670 ;
        RECT 1732.930 119.090 1734.110 120.270 ;
        RECT 1732.930 117.490 1734.110 118.670 ;
        RECT 1732.930 -17.010 1734.110 -15.830 ;
        RECT 1732.930 -18.610 1734.110 -17.430 ;
        RECT 1750.930 2117.090 1752.110 2118.270 ;
        RECT 1750.930 2115.490 1752.110 2116.670 ;
        RECT 1750.930 1937.090 1752.110 1938.270 ;
        RECT 1750.930 1935.490 1752.110 1936.670 ;
        RECT 1750.930 1757.090 1752.110 1758.270 ;
        RECT 1750.930 1755.490 1752.110 1756.670 ;
        RECT 1750.930 1577.090 1752.110 1578.270 ;
        RECT 1750.930 1575.490 1752.110 1576.670 ;
        RECT 1750.930 1397.090 1752.110 1398.270 ;
        RECT 1750.930 1395.490 1752.110 1396.670 ;
        RECT 1750.930 1217.090 1752.110 1218.270 ;
        RECT 1750.930 1215.490 1752.110 1216.670 ;
        RECT 1750.930 1037.090 1752.110 1038.270 ;
        RECT 1750.930 1035.490 1752.110 1036.670 ;
        RECT 1750.930 857.090 1752.110 858.270 ;
        RECT 1750.930 855.490 1752.110 856.670 ;
        RECT 1750.930 677.090 1752.110 678.270 ;
        RECT 1750.930 675.490 1752.110 676.670 ;
        RECT 1750.930 497.090 1752.110 498.270 ;
        RECT 1750.930 495.490 1752.110 496.670 ;
        RECT 1750.930 317.090 1752.110 318.270 ;
        RECT 1750.930 315.490 1752.110 316.670 ;
        RECT 1750.930 137.090 1752.110 138.270 ;
        RECT 1750.930 135.490 1752.110 136.670 ;
        RECT 1750.930 -26.410 1752.110 -25.230 ;
        RECT 1750.930 -28.010 1752.110 -26.830 ;
        RECT 1768.930 2135.090 1770.110 2136.270 ;
        RECT 1768.930 2133.490 1770.110 2134.670 ;
        RECT 1768.930 1955.090 1770.110 1956.270 ;
        RECT 1768.930 1953.490 1770.110 1954.670 ;
        RECT 1768.930 1775.090 1770.110 1776.270 ;
        RECT 1768.930 1773.490 1770.110 1774.670 ;
        RECT 1768.930 1595.090 1770.110 1596.270 ;
        RECT 1768.930 1593.490 1770.110 1594.670 ;
        RECT 1768.930 1415.090 1770.110 1416.270 ;
        RECT 1768.930 1413.490 1770.110 1414.670 ;
        RECT 1768.930 1235.090 1770.110 1236.270 ;
        RECT 1768.930 1233.490 1770.110 1234.670 ;
        RECT 1768.930 1055.090 1770.110 1056.270 ;
        RECT 1768.930 1053.490 1770.110 1054.670 ;
        RECT 1768.930 875.090 1770.110 876.270 ;
        RECT 1768.930 873.490 1770.110 874.670 ;
        RECT 1768.930 695.090 1770.110 696.270 ;
        RECT 1768.930 693.490 1770.110 694.670 ;
        RECT 1768.930 515.090 1770.110 516.270 ;
        RECT 1768.930 513.490 1770.110 514.670 ;
        RECT 1768.930 335.090 1770.110 336.270 ;
        RECT 1768.930 333.490 1770.110 334.670 ;
        RECT 1768.930 155.090 1770.110 156.270 ;
        RECT 1768.930 153.490 1770.110 154.670 ;
        RECT 1588.930 -35.810 1590.110 -34.630 ;
        RECT 1588.930 -37.410 1590.110 -36.230 ;
        RECT 1894.930 2261.090 1896.110 2262.270 ;
        RECT 1894.930 2259.490 1896.110 2260.670 ;
        RECT 1894.930 2081.090 1896.110 2082.270 ;
        RECT 1894.930 2079.490 1896.110 2080.670 ;
        RECT 1894.930 1901.090 1896.110 1902.270 ;
        RECT 1894.930 1899.490 1896.110 1900.670 ;
        RECT 1894.930 1721.090 1896.110 1722.270 ;
        RECT 1894.930 1719.490 1896.110 1720.670 ;
        RECT 1894.930 1541.090 1896.110 1542.270 ;
        RECT 1894.930 1539.490 1896.110 1540.670 ;
        RECT 1894.930 1361.090 1896.110 1362.270 ;
        RECT 1894.930 1359.490 1896.110 1360.670 ;
        RECT 1894.930 1181.090 1896.110 1182.270 ;
        RECT 1894.930 1179.490 1896.110 1180.670 ;
        RECT 1894.930 1001.090 1896.110 1002.270 ;
        RECT 1894.930 999.490 1896.110 1000.670 ;
        RECT 1894.930 821.090 1896.110 822.270 ;
        RECT 1894.930 819.490 1896.110 820.670 ;
        RECT 1894.930 641.090 1896.110 642.270 ;
        RECT 1894.930 639.490 1896.110 640.670 ;
        RECT 1894.930 461.090 1896.110 462.270 ;
        RECT 1894.930 459.490 1896.110 460.670 ;
        RECT 1894.930 281.090 1896.110 282.270 ;
        RECT 1894.930 279.490 1896.110 280.670 ;
        RECT 1894.930 101.090 1896.110 102.270 ;
        RECT 1894.930 99.490 1896.110 100.670 ;
        RECT 1894.930 -7.610 1896.110 -6.430 ;
        RECT 1894.930 -9.210 1896.110 -8.030 ;
        RECT 1912.930 2279.090 1914.110 2280.270 ;
        RECT 1912.930 2277.490 1914.110 2278.670 ;
        RECT 1912.930 2099.090 1914.110 2100.270 ;
        RECT 1912.930 2097.490 1914.110 2098.670 ;
        RECT 1912.930 1919.090 1914.110 1920.270 ;
        RECT 1912.930 1917.490 1914.110 1918.670 ;
        RECT 1912.930 1739.090 1914.110 1740.270 ;
        RECT 1912.930 1737.490 1914.110 1738.670 ;
        RECT 1912.930 1559.090 1914.110 1560.270 ;
        RECT 1912.930 1557.490 1914.110 1558.670 ;
        RECT 1912.930 1379.090 1914.110 1380.270 ;
        RECT 1912.930 1377.490 1914.110 1378.670 ;
        RECT 1912.930 1199.090 1914.110 1200.270 ;
        RECT 1912.930 1197.490 1914.110 1198.670 ;
        RECT 1912.930 1019.090 1914.110 1020.270 ;
        RECT 1912.930 1017.490 1914.110 1018.670 ;
        RECT 1912.930 839.090 1914.110 840.270 ;
        RECT 1912.930 837.490 1914.110 838.670 ;
        RECT 1912.930 659.090 1914.110 660.270 ;
        RECT 1912.930 657.490 1914.110 658.670 ;
        RECT 1912.930 479.090 1914.110 480.270 ;
        RECT 1912.930 477.490 1914.110 478.670 ;
        RECT 1912.930 299.090 1914.110 300.270 ;
        RECT 1912.930 297.490 1914.110 298.670 ;
        RECT 1912.930 119.090 1914.110 120.270 ;
        RECT 1912.930 117.490 1914.110 118.670 ;
        RECT 1912.930 -17.010 1914.110 -15.830 ;
        RECT 1912.930 -18.610 1914.110 -17.430 ;
        RECT 1930.930 2117.090 1932.110 2118.270 ;
        RECT 1930.930 2115.490 1932.110 2116.670 ;
        RECT 1930.930 1937.090 1932.110 1938.270 ;
        RECT 1930.930 1935.490 1932.110 1936.670 ;
        RECT 1930.930 1757.090 1932.110 1758.270 ;
        RECT 1930.930 1755.490 1932.110 1756.670 ;
        RECT 1930.930 1577.090 1932.110 1578.270 ;
        RECT 1930.930 1575.490 1932.110 1576.670 ;
        RECT 1930.930 1397.090 1932.110 1398.270 ;
        RECT 1930.930 1395.490 1932.110 1396.670 ;
        RECT 1930.930 1217.090 1932.110 1218.270 ;
        RECT 1930.930 1215.490 1932.110 1216.670 ;
        RECT 1930.930 1037.090 1932.110 1038.270 ;
        RECT 1930.930 1035.490 1932.110 1036.670 ;
        RECT 1930.930 857.090 1932.110 858.270 ;
        RECT 1930.930 855.490 1932.110 856.670 ;
        RECT 1930.930 677.090 1932.110 678.270 ;
        RECT 1930.930 675.490 1932.110 676.670 ;
        RECT 1930.930 497.090 1932.110 498.270 ;
        RECT 1930.930 495.490 1932.110 496.670 ;
        RECT 1930.930 317.090 1932.110 318.270 ;
        RECT 1930.930 315.490 1932.110 316.670 ;
        RECT 1930.930 137.090 1932.110 138.270 ;
        RECT 1930.930 135.490 1932.110 136.670 ;
        RECT 1930.930 -26.410 1932.110 -25.230 ;
        RECT 1930.930 -28.010 1932.110 -26.830 ;
        RECT 1948.930 2135.090 1950.110 2136.270 ;
        RECT 1948.930 2133.490 1950.110 2134.670 ;
        RECT 1948.930 1955.090 1950.110 1956.270 ;
        RECT 1948.930 1953.490 1950.110 1954.670 ;
        RECT 1948.930 1775.090 1950.110 1776.270 ;
        RECT 1948.930 1773.490 1950.110 1774.670 ;
        RECT 1948.930 1595.090 1950.110 1596.270 ;
        RECT 1948.930 1593.490 1950.110 1594.670 ;
        RECT 1948.930 1415.090 1950.110 1416.270 ;
        RECT 1948.930 1413.490 1950.110 1414.670 ;
        RECT 1948.930 1235.090 1950.110 1236.270 ;
        RECT 1948.930 1233.490 1950.110 1234.670 ;
        RECT 1948.930 1055.090 1950.110 1056.270 ;
        RECT 1948.930 1053.490 1950.110 1054.670 ;
        RECT 1948.930 875.090 1950.110 876.270 ;
        RECT 1948.930 873.490 1950.110 874.670 ;
        RECT 1948.930 695.090 1950.110 696.270 ;
        RECT 1948.930 693.490 1950.110 694.670 ;
        RECT 1948.930 515.090 1950.110 516.270 ;
        RECT 1948.930 513.490 1950.110 514.670 ;
        RECT 1948.930 335.090 1950.110 336.270 ;
        RECT 1948.930 333.490 1950.110 334.670 ;
        RECT 1948.930 155.090 1950.110 156.270 ;
        RECT 1948.930 153.490 1950.110 154.670 ;
        RECT 1768.930 -35.810 1770.110 -34.630 ;
        RECT 1768.930 -37.410 1770.110 -36.230 ;
        RECT 2074.930 2261.090 2076.110 2262.270 ;
        RECT 2074.930 2259.490 2076.110 2260.670 ;
        RECT 2074.930 2081.090 2076.110 2082.270 ;
        RECT 2074.930 2079.490 2076.110 2080.670 ;
        RECT 2074.930 1901.090 2076.110 1902.270 ;
        RECT 2074.930 1899.490 2076.110 1900.670 ;
        RECT 2074.930 1721.090 2076.110 1722.270 ;
        RECT 2074.930 1719.490 2076.110 1720.670 ;
        RECT 2074.930 1541.090 2076.110 1542.270 ;
        RECT 2074.930 1539.490 2076.110 1540.670 ;
        RECT 2074.930 1361.090 2076.110 1362.270 ;
        RECT 2074.930 1359.490 2076.110 1360.670 ;
        RECT 2074.930 1181.090 2076.110 1182.270 ;
        RECT 2074.930 1179.490 2076.110 1180.670 ;
        RECT 2074.930 1001.090 2076.110 1002.270 ;
        RECT 2074.930 999.490 2076.110 1000.670 ;
        RECT 2074.930 821.090 2076.110 822.270 ;
        RECT 2074.930 819.490 2076.110 820.670 ;
        RECT 2074.930 641.090 2076.110 642.270 ;
        RECT 2074.930 639.490 2076.110 640.670 ;
        RECT 2074.930 461.090 2076.110 462.270 ;
        RECT 2074.930 459.490 2076.110 460.670 ;
        RECT 2074.930 281.090 2076.110 282.270 ;
        RECT 2074.930 279.490 2076.110 280.670 ;
        RECT 2074.930 101.090 2076.110 102.270 ;
        RECT 2074.930 99.490 2076.110 100.670 ;
        RECT 2074.930 -7.610 2076.110 -6.430 ;
        RECT 2074.930 -9.210 2076.110 -8.030 ;
        RECT 2092.930 3359.090 2094.110 3360.270 ;
        RECT 2092.930 3357.490 2094.110 3358.670 ;
        RECT 2092.930 3179.090 2094.110 3180.270 ;
        RECT 2092.930 3177.490 2094.110 3178.670 ;
        RECT 2092.930 2999.090 2094.110 3000.270 ;
        RECT 2092.930 2997.490 2094.110 2998.670 ;
        RECT 2092.930 2819.090 2094.110 2820.270 ;
        RECT 2092.930 2817.490 2094.110 2818.670 ;
        RECT 2092.930 2639.090 2094.110 2640.270 ;
        RECT 2092.930 2637.490 2094.110 2638.670 ;
        RECT 2092.930 2459.090 2094.110 2460.270 ;
        RECT 2092.930 2457.490 2094.110 2458.670 ;
        RECT 2092.930 2279.090 2094.110 2280.270 ;
        RECT 2092.930 2277.490 2094.110 2278.670 ;
        RECT 2092.930 2099.090 2094.110 2100.270 ;
        RECT 2092.930 2097.490 2094.110 2098.670 ;
        RECT 2092.930 1919.090 2094.110 1920.270 ;
        RECT 2092.930 1917.490 2094.110 1918.670 ;
        RECT 2092.930 1739.090 2094.110 1740.270 ;
        RECT 2092.930 1737.490 2094.110 1738.670 ;
        RECT 2092.930 1559.090 2094.110 1560.270 ;
        RECT 2092.930 1557.490 2094.110 1558.670 ;
        RECT 2092.930 1379.090 2094.110 1380.270 ;
        RECT 2092.930 1377.490 2094.110 1378.670 ;
        RECT 2092.930 1199.090 2094.110 1200.270 ;
        RECT 2092.930 1197.490 2094.110 1198.670 ;
        RECT 2092.930 1019.090 2094.110 1020.270 ;
        RECT 2092.930 1017.490 2094.110 1018.670 ;
        RECT 2092.930 839.090 2094.110 840.270 ;
        RECT 2092.930 837.490 2094.110 838.670 ;
        RECT 2092.930 659.090 2094.110 660.270 ;
        RECT 2092.930 657.490 2094.110 658.670 ;
        RECT 2092.930 479.090 2094.110 480.270 ;
        RECT 2092.930 477.490 2094.110 478.670 ;
        RECT 2092.930 299.090 2094.110 300.270 ;
        RECT 2092.930 297.490 2094.110 298.670 ;
        RECT 2092.930 119.090 2094.110 120.270 ;
        RECT 2092.930 117.490 2094.110 118.670 ;
        RECT 2092.930 -17.010 2094.110 -15.830 ;
        RECT 2092.930 -18.610 2094.110 -17.430 ;
        RECT 2110.930 3377.090 2112.110 3378.270 ;
        RECT 2110.930 3375.490 2112.110 3376.670 ;
        RECT 2110.930 3197.090 2112.110 3198.270 ;
        RECT 2110.930 3195.490 2112.110 3196.670 ;
        RECT 2110.930 3017.090 2112.110 3018.270 ;
        RECT 2110.930 3015.490 2112.110 3016.670 ;
        RECT 2110.930 2837.090 2112.110 2838.270 ;
        RECT 2110.930 2835.490 2112.110 2836.670 ;
        RECT 2110.930 2657.090 2112.110 2658.270 ;
        RECT 2110.930 2655.490 2112.110 2656.670 ;
        RECT 2110.930 2477.090 2112.110 2478.270 ;
        RECT 2110.930 2475.490 2112.110 2476.670 ;
        RECT 2110.930 2297.090 2112.110 2298.270 ;
        RECT 2110.930 2295.490 2112.110 2296.670 ;
        RECT 2110.930 2117.090 2112.110 2118.270 ;
        RECT 2110.930 2115.490 2112.110 2116.670 ;
        RECT 2110.930 1937.090 2112.110 1938.270 ;
        RECT 2110.930 1935.490 2112.110 1936.670 ;
        RECT 2110.930 1757.090 2112.110 1758.270 ;
        RECT 2110.930 1755.490 2112.110 1756.670 ;
        RECT 2110.930 1577.090 2112.110 1578.270 ;
        RECT 2110.930 1575.490 2112.110 1576.670 ;
        RECT 2110.930 1397.090 2112.110 1398.270 ;
        RECT 2110.930 1395.490 2112.110 1396.670 ;
        RECT 2110.930 1217.090 2112.110 1218.270 ;
        RECT 2110.930 1215.490 2112.110 1216.670 ;
        RECT 2110.930 1037.090 2112.110 1038.270 ;
        RECT 2110.930 1035.490 2112.110 1036.670 ;
        RECT 2110.930 857.090 2112.110 858.270 ;
        RECT 2110.930 855.490 2112.110 856.670 ;
        RECT 2110.930 677.090 2112.110 678.270 ;
        RECT 2110.930 675.490 2112.110 676.670 ;
        RECT 2110.930 497.090 2112.110 498.270 ;
        RECT 2110.930 495.490 2112.110 496.670 ;
        RECT 2110.930 317.090 2112.110 318.270 ;
        RECT 2110.930 315.490 2112.110 316.670 ;
        RECT 2110.930 137.090 2112.110 138.270 ;
        RECT 2110.930 135.490 2112.110 136.670 ;
        RECT 2110.930 -26.410 2112.110 -25.230 ;
        RECT 2110.930 -28.010 2112.110 -26.830 ;
        RECT 2308.930 3555.910 2310.110 3557.090 ;
        RECT 2308.930 3554.310 2310.110 3555.490 ;
        RECT 2290.930 3546.510 2292.110 3547.690 ;
        RECT 2290.930 3544.910 2292.110 3546.090 ;
        RECT 2272.930 3537.110 2274.110 3538.290 ;
        RECT 2272.930 3535.510 2274.110 3536.690 ;
        RECT 2128.930 3395.090 2130.110 3396.270 ;
        RECT 2128.930 3393.490 2130.110 3394.670 ;
        RECT 2128.930 3215.090 2130.110 3216.270 ;
        RECT 2128.930 3213.490 2130.110 3214.670 ;
        RECT 2128.930 3035.090 2130.110 3036.270 ;
        RECT 2128.930 3033.490 2130.110 3034.670 ;
        RECT 2128.930 2855.090 2130.110 2856.270 ;
        RECT 2128.930 2853.490 2130.110 2854.670 ;
        RECT 2254.930 3527.710 2256.110 3528.890 ;
        RECT 2254.930 3526.110 2256.110 3527.290 ;
        RECT 2254.930 3341.090 2256.110 3342.270 ;
        RECT 2254.930 3339.490 2256.110 3340.670 ;
        RECT 2254.930 3161.090 2256.110 3162.270 ;
        RECT 2254.930 3159.490 2256.110 3160.670 ;
        RECT 2254.930 2981.090 2256.110 2982.270 ;
        RECT 2254.930 2979.490 2256.110 2980.670 ;
        RECT 2254.930 2801.090 2256.110 2802.270 ;
        RECT 2254.930 2799.490 2256.110 2800.670 ;
        RECT 2272.930 3359.090 2274.110 3360.270 ;
        RECT 2272.930 3357.490 2274.110 3358.670 ;
        RECT 2272.930 3179.090 2274.110 3180.270 ;
        RECT 2272.930 3177.490 2274.110 3178.670 ;
        RECT 2272.930 2999.090 2274.110 3000.270 ;
        RECT 2272.930 2997.490 2274.110 2998.670 ;
        RECT 2272.930 2819.090 2274.110 2820.270 ;
        RECT 2272.930 2817.490 2274.110 2818.670 ;
        RECT 2290.930 3377.090 2292.110 3378.270 ;
        RECT 2290.930 3375.490 2292.110 3376.670 ;
        RECT 2290.930 3197.090 2292.110 3198.270 ;
        RECT 2290.930 3195.490 2292.110 3196.670 ;
        RECT 2290.930 3017.090 2292.110 3018.270 ;
        RECT 2290.930 3015.490 2292.110 3016.670 ;
        RECT 2290.930 2837.090 2292.110 2838.270 ;
        RECT 2290.930 2835.490 2292.110 2836.670 ;
        RECT 2488.930 3555.910 2490.110 3557.090 ;
        RECT 2488.930 3554.310 2490.110 3555.490 ;
        RECT 2470.930 3546.510 2472.110 3547.690 ;
        RECT 2470.930 3544.910 2472.110 3546.090 ;
        RECT 2452.930 3537.110 2454.110 3538.290 ;
        RECT 2452.930 3535.510 2454.110 3536.690 ;
        RECT 2308.930 3395.090 2310.110 3396.270 ;
        RECT 2308.930 3393.490 2310.110 3394.670 ;
        RECT 2308.930 3215.090 2310.110 3216.270 ;
        RECT 2308.930 3213.490 2310.110 3214.670 ;
        RECT 2308.930 3035.090 2310.110 3036.270 ;
        RECT 2308.930 3033.490 2310.110 3034.670 ;
        RECT 2308.930 2855.090 2310.110 2856.270 ;
        RECT 2308.930 2853.490 2310.110 2854.670 ;
        RECT 2434.930 3527.710 2436.110 3528.890 ;
        RECT 2434.930 3526.110 2436.110 3527.290 ;
        RECT 2434.930 3341.090 2436.110 3342.270 ;
        RECT 2434.930 3339.490 2436.110 3340.670 ;
        RECT 2434.930 3161.090 2436.110 3162.270 ;
        RECT 2434.930 3159.490 2436.110 3160.670 ;
        RECT 2434.930 2981.090 2436.110 2982.270 ;
        RECT 2434.930 2979.490 2436.110 2980.670 ;
        RECT 2434.930 2801.090 2436.110 2802.270 ;
        RECT 2434.930 2799.490 2436.110 2800.670 ;
        RECT 2452.930 3359.090 2454.110 3360.270 ;
        RECT 2452.930 3357.490 2454.110 3358.670 ;
        RECT 2452.930 3179.090 2454.110 3180.270 ;
        RECT 2452.930 3177.490 2454.110 3178.670 ;
        RECT 2452.930 2999.090 2454.110 3000.270 ;
        RECT 2452.930 2997.490 2454.110 2998.670 ;
        RECT 2452.930 2819.090 2454.110 2820.270 ;
        RECT 2452.930 2817.490 2454.110 2818.670 ;
        RECT 2470.930 3377.090 2472.110 3378.270 ;
        RECT 2470.930 3375.490 2472.110 3376.670 ;
        RECT 2470.930 3197.090 2472.110 3198.270 ;
        RECT 2470.930 3195.490 2472.110 3196.670 ;
        RECT 2470.930 3017.090 2472.110 3018.270 ;
        RECT 2470.930 3015.490 2472.110 3016.670 ;
        RECT 2470.930 2837.090 2472.110 2838.270 ;
        RECT 2470.930 2835.490 2472.110 2836.670 ;
        RECT 2668.930 3555.910 2670.110 3557.090 ;
        RECT 2668.930 3554.310 2670.110 3555.490 ;
        RECT 2650.930 3546.510 2652.110 3547.690 ;
        RECT 2650.930 3544.910 2652.110 3546.090 ;
        RECT 2632.930 3537.110 2634.110 3538.290 ;
        RECT 2632.930 3535.510 2634.110 3536.690 ;
        RECT 2488.930 3395.090 2490.110 3396.270 ;
        RECT 2488.930 3393.490 2490.110 3394.670 ;
        RECT 2488.930 3215.090 2490.110 3216.270 ;
        RECT 2488.930 3213.490 2490.110 3214.670 ;
        RECT 2488.930 3035.090 2490.110 3036.270 ;
        RECT 2488.930 3033.490 2490.110 3034.670 ;
        RECT 2488.930 2855.090 2490.110 2856.270 ;
        RECT 2488.930 2853.490 2490.110 2854.670 ;
        RECT 2614.930 3527.710 2616.110 3528.890 ;
        RECT 2614.930 3526.110 2616.110 3527.290 ;
        RECT 2614.930 3341.090 2616.110 3342.270 ;
        RECT 2614.930 3339.490 2616.110 3340.670 ;
        RECT 2614.930 3161.090 2616.110 3162.270 ;
        RECT 2614.930 3159.490 2616.110 3160.670 ;
        RECT 2614.930 2981.090 2616.110 2982.270 ;
        RECT 2614.930 2979.490 2616.110 2980.670 ;
        RECT 2614.930 2801.090 2616.110 2802.270 ;
        RECT 2614.930 2799.490 2616.110 2800.670 ;
        RECT 2128.930 2675.090 2130.110 2676.270 ;
        RECT 2128.930 2673.490 2130.110 2674.670 ;
        RECT 2128.930 2495.090 2130.110 2496.270 ;
        RECT 2128.930 2493.490 2130.110 2494.670 ;
        RECT 2128.930 2315.090 2130.110 2316.270 ;
        RECT 2128.930 2313.490 2130.110 2314.670 ;
        RECT 2584.910 2675.090 2586.090 2676.270 ;
        RECT 2584.910 2673.490 2586.090 2674.670 ;
        RECT 2584.910 2657.090 2586.090 2658.270 ;
        RECT 2584.910 2655.490 2586.090 2656.670 ;
        RECT 2584.910 2639.090 2586.090 2640.270 ;
        RECT 2584.910 2637.490 2586.090 2638.670 ;
        RECT 2584.910 2621.090 2586.090 2622.270 ;
        RECT 2584.910 2619.490 2586.090 2620.670 ;
        RECT 2584.910 2495.090 2586.090 2496.270 ;
        RECT 2584.910 2493.490 2586.090 2494.670 ;
        RECT 2584.910 2477.090 2586.090 2478.270 ;
        RECT 2584.910 2475.490 2586.090 2476.670 ;
        RECT 2584.910 2459.090 2586.090 2460.270 ;
        RECT 2584.910 2457.490 2586.090 2458.670 ;
        RECT 2584.910 2441.090 2586.090 2442.270 ;
        RECT 2584.910 2439.490 2586.090 2440.670 ;
        RECT 2584.910 2315.090 2586.090 2316.270 ;
        RECT 2584.910 2313.490 2586.090 2314.670 ;
        RECT 2614.930 2621.090 2616.110 2622.270 ;
        RECT 2614.930 2619.490 2616.110 2620.670 ;
        RECT 2614.930 2441.090 2616.110 2442.270 ;
        RECT 2614.930 2439.490 2616.110 2440.670 ;
        RECT 2128.930 2135.090 2130.110 2136.270 ;
        RECT 2128.930 2133.490 2130.110 2134.670 ;
        RECT 2128.930 1955.090 2130.110 1956.270 ;
        RECT 2128.930 1953.490 2130.110 1954.670 ;
        RECT 2128.930 1775.090 2130.110 1776.270 ;
        RECT 2128.930 1773.490 2130.110 1774.670 ;
        RECT 2128.930 1595.090 2130.110 1596.270 ;
        RECT 2128.930 1593.490 2130.110 1594.670 ;
        RECT 2128.930 1415.090 2130.110 1416.270 ;
        RECT 2128.930 1413.490 2130.110 1414.670 ;
        RECT 2128.930 1235.090 2130.110 1236.270 ;
        RECT 2128.930 1233.490 2130.110 1234.670 ;
        RECT 2128.930 1055.090 2130.110 1056.270 ;
        RECT 2128.930 1053.490 2130.110 1054.670 ;
        RECT 2128.930 875.090 2130.110 876.270 ;
        RECT 2128.930 873.490 2130.110 874.670 ;
        RECT 2128.930 695.090 2130.110 696.270 ;
        RECT 2128.930 693.490 2130.110 694.670 ;
        RECT 2128.930 515.090 2130.110 516.270 ;
        RECT 2128.930 513.490 2130.110 514.670 ;
        RECT 2128.930 335.090 2130.110 336.270 ;
        RECT 2128.930 333.490 2130.110 334.670 ;
        RECT 2128.930 155.090 2130.110 156.270 ;
        RECT 2128.930 153.490 2130.110 154.670 ;
        RECT 1948.930 -35.810 1950.110 -34.630 ;
        RECT 1948.930 -37.410 1950.110 -36.230 ;
        RECT 2254.930 2261.090 2256.110 2262.270 ;
        RECT 2254.930 2259.490 2256.110 2260.670 ;
        RECT 2254.930 2081.090 2256.110 2082.270 ;
        RECT 2254.930 2079.490 2256.110 2080.670 ;
        RECT 2254.930 1901.090 2256.110 1902.270 ;
        RECT 2254.930 1899.490 2256.110 1900.670 ;
        RECT 2254.930 1721.090 2256.110 1722.270 ;
        RECT 2254.930 1719.490 2256.110 1720.670 ;
        RECT 2254.930 1541.090 2256.110 1542.270 ;
        RECT 2254.930 1539.490 2256.110 1540.670 ;
        RECT 2254.930 1361.090 2256.110 1362.270 ;
        RECT 2254.930 1359.490 2256.110 1360.670 ;
        RECT 2254.930 1181.090 2256.110 1182.270 ;
        RECT 2254.930 1179.490 2256.110 1180.670 ;
        RECT 2254.930 1001.090 2256.110 1002.270 ;
        RECT 2254.930 999.490 2256.110 1000.670 ;
        RECT 2254.930 821.090 2256.110 822.270 ;
        RECT 2254.930 819.490 2256.110 820.670 ;
        RECT 2254.930 641.090 2256.110 642.270 ;
        RECT 2254.930 639.490 2256.110 640.670 ;
        RECT 2254.930 461.090 2256.110 462.270 ;
        RECT 2254.930 459.490 2256.110 460.670 ;
        RECT 2254.930 281.090 2256.110 282.270 ;
        RECT 2254.930 279.490 2256.110 280.670 ;
        RECT 2254.930 101.090 2256.110 102.270 ;
        RECT 2254.930 99.490 2256.110 100.670 ;
        RECT 2254.930 -7.610 2256.110 -6.430 ;
        RECT 2254.930 -9.210 2256.110 -8.030 ;
        RECT 2272.930 2279.090 2274.110 2280.270 ;
        RECT 2272.930 2277.490 2274.110 2278.670 ;
        RECT 2272.930 2099.090 2274.110 2100.270 ;
        RECT 2272.930 2097.490 2274.110 2098.670 ;
        RECT 2272.930 1919.090 2274.110 1920.270 ;
        RECT 2272.930 1917.490 2274.110 1918.670 ;
        RECT 2272.930 1739.090 2274.110 1740.270 ;
        RECT 2272.930 1737.490 2274.110 1738.670 ;
        RECT 2272.930 1559.090 2274.110 1560.270 ;
        RECT 2272.930 1557.490 2274.110 1558.670 ;
        RECT 2272.930 1379.090 2274.110 1380.270 ;
        RECT 2272.930 1377.490 2274.110 1378.670 ;
        RECT 2272.930 1199.090 2274.110 1200.270 ;
        RECT 2272.930 1197.490 2274.110 1198.670 ;
        RECT 2272.930 1019.090 2274.110 1020.270 ;
        RECT 2272.930 1017.490 2274.110 1018.670 ;
        RECT 2272.930 839.090 2274.110 840.270 ;
        RECT 2272.930 837.490 2274.110 838.670 ;
        RECT 2272.930 659.090 2274.110 660.270 ;
        RECT 2272.930 657.490 2274.110 658.670 ;
        RECT 2272.930 479.090 2274.110 480.270 ;
        RECT 2272.930 477.490 2274.110 478.670 ;
        RECT 2272.930 299.090 2274.110 300.270 ;
        RECT 2272.930 297.490 2274.110 298.670 ;
        RECT 2272.930 119.090 2274.110 120.270 ;
        RECT 2272.930 117.490 2274.110 118.670 ;
        RECT 2272.930 -17.010 2274.110 -15.830 ;
        RECT 2272.930 -18.610 2274.110 -17.430 ;
        RECT 2290.930 2117.090 2292.110 2118.270 ;
        RECT 2290.930 2115.490 2292.110 2116.670 ;
        RECT 2290.930 1937.090 2292.110 1938.270 ;
        RECT 2290.930 1935.490 2292.110 1936.670 ;
        RECT 2290.930 1757.090 2292.110 1758.270 ;
        RECT 2290.930 1755.490 2292.110 1756.670 ;
        RECT 2290.930 1577.090 2292.110 1578.270 ;
        RECT 2290.930 1575.490 2292.110 1576.670 ;
        RECT 2290.930 1397.090 2292.110 1398.270 ;
        RECT 2290.930 1395.490 2292.110 1396.670 ;
        RECT 2290.930 1217.090 2292.110 1218.270 ;
        RECT 2290.930 1215.490 2292.110 1216.670 ;
        RECT 2290.930 1037.090 2292.110 1038.270 ;
        RECT 2290.930 1035.490 2292.110 1036.670 ;
        RECT 2290.930 857.090 2292.110 858.270 ;
        RECT 2290.930 855.490 2292.110 856.670 ;
        RECT 2290.930 677.090 2292.110 678.270 ;
        RECT 2290.930 675.490 2292.110 676.670 ;
        RECT 2290.930 497.090 2292.110 498.270 ;
        RECT 2290.930 495.490 2292.110 496.670 ;
        RECT 2290.930 317.090 2292.110 318.270 ;
        RECT 2290.930 315.490 2292.110 316.670 ;
        RECT 2290.930 137.090 2292.110 138.270 ;
        RECT 2290.930 135.490 2292.110 136.670 ;
        RECT 2290.930 -26.410 2292.110 -25.230 ;
        RECT 2290.930 -28.010 2292.110 -26.830 ;
        RECT 2308.930 2135.090 2310.110 2136.270 ;
        RECT 2308.930 2133.490 2310.110 2134.670 ;
        RECT 2308.930 1955.090 2310.110 1956.270 ;
        RECT 2308.930 1953.490 2310.110 1954.670 ;
        RECT 2308.930 1775.090 2310.110 1776.270 ;
        RECT 2308.930 1773.490 2310.110 1774.670 ;
        RECT 2308.930 1595.090 2310.110 1596.270 ;
        RECT 2308.930 1593.490 2310.110 1594.670 ;
        RECT 2308.930 1415.090 2310.110 1416.270 ;
        RECT 2308.930 1413.490 2310.110 1414.670 ;
        RECT 2308.930 1235.090 2310.110 1236.270 ;
        RECT 2308.930 1233.490 2310.110 1234.670 ;
        RECT 2308.930 1055.090 2310.110 1056.270 ;
        RECT 2308.930 1053.490 2310.110 1054.670 ;
        RECT 2308.930 875.090 2310.110 876.270 ;
        RECT 2308.930 873.490 2310.110 874.670 ;
        RECT 2308.930 695.090 2310.110 696.270 ;
        RECT 2308.930 693.490 2310.110 694.670 ;
        RECT 2308.930 515.090 2310.110 516.270 ;
        RECT 2308.930 513.490 2310.110 514.670 ;
        RECT 2308.930 335.090 2310.110 336.270 ;
        RECT 2308.930 333.490 2310.110 334.670 ;
        RECT 2308.930 155.090 2310.110 156.270 ;
        RECT 2308.930 153.490 2310.110 154.670 ;
        RECT 2128.930 -35.810 2130.110 -34.630 ;
        RECT 2128.930 -37.410 2130.110 -36.230 ;
        RECT 2434.930 2261.090 2436.110 2262.270 ;
        RECT 2434.930 2259.490 2436.110 2260.670 ;
        RECT 2434.930 2081.090 2436.110 2082.270 ;
        RECT 2434.930 2079.490 2436.110 2080.670 ;
        RECT 2434.930 1901.090 2436.110 1902.270 ;
        RECT 2434.930 1899.490 2436.110 1900.670 ;
        RECT 2434.930 1721.090 2436.110 1722.270 ;
        RECT 2434.930 1719.490 2436.110 1720.670 ;
        RECT 2434.930 1541.090 2436.110 1542.270 ;
        RECT 2434.930 1539.490 2436.110 1540.670 ;
        RECT 2434.930 1361.090 2436.110 1362.270 ;
        RECT 2434.930 1359.490 2436.110 1360.670 ;
        RECT 2434.930 1181.090 2436.110 1182.270 ;
        RECT 2434.930 1179.490 2436.110 1180.670 ;
        RECT 2434.930 1001.090 2436.110 1002.270 ;
        RECT 2434.930 999.490 2436.110 1000.670 ;
        RECT 2434.930 821.090 2436.110 822.270 ;
        RECT 2434.930 819.490 2436.110 820.670 ;
        RECT 2434.930 641.090 2436.110 642.270 ;
        RECT 2434.930 639.490 2436.110 640.670 ;
        RECT 2434.930 461.090 2436.110 462.270 ;
        RECT 2434.930 459.490 2436.110 460.670 ;
        RECT 2434.930 281.090 2436.110 282.270 ;
        RECT 2434.930 279.490 2436.110 280.670 ;
        RECT 2434.930 101.090 2436.110 102.270 ;
        RECT 2434.930 99.490 2436.110 100.670 ;
        RECT 2434.930 -7.610 2436.110 -6.430 ;
        RECT 2434.930 -9.210 2436.110 -8.030 ;
        RECT 2452.930 2279.090 2454.110 2280.270 ;
        RECT 2452.930 2277.490 2454.110 2278.670 ;
        RECT 2452.930 2099.090 2454.110 2100.270 ;
        RECT 2452.930 2097.490 2454.110 2098.670 ;
        RECT 2452.930 1919.090 2454.110 1920.270 ;
        RECT 2452.930 1917.490 2454.110 1918.670 ;
        RECT 2452.930 1739.090 2454.110 1740.270 ;
        RECT 2452.930 1737.490 2454.110 1738.670 ;
        RECT 2452.930 1559.090 2454.110 1560.270 ;
        RECT 2452.930 1557.490 2454.110 1558.670 ;
        RECT 2452.930 1379.090 2454.110 1380.270 ;
        RECT 2452.930 1377.490 2454.110 1378.670 ;
        RECT 2452.930 1199.090 2454.110 1200.270 ;
        RECT 2452.930 1197.490 2454.110 1198.670 ;
        RECT 2452.930 1019.090 2454.110 1020.270 ;
        RECT 2452.930 1017.490 2454.110 1018.670 ;
        RECT 2452.930 839.090 2454.110 840.270 ;
        RECT 2452.930 837.490 2454.110 838.670 ;
        RECT 2452.930 659.090 2454.110 660.270 ;
        RECT 2452.930 657.490 2454.110 658.670 ;
        RECT 2452.930 479.090 2454.110 480.270 ;
        RECT 2452.930 477.490 2454.110 478.670 ;
        RECT 2452.930 299.090 2454.110 300.270 ;
        RECT 2452.930 297.490 2454.110 298.670 ;
        RECT 2452.930 119.090 2454.110 120.270 ;
        RECT 2452.930 117.490 2454.110 118.670 ;
        RECT 2452.930 -17.010 2454.110 -15.830 ;
        RECT 2452.930 -18.610 2454.110 -17.430 ;
        RECT 2470.930 2117.090 2472.110 2118.270 ;
        RECT 2470.930 2115.490 2472.110 2116.670 ;
        RECT 2470.930 1937.090 2472.110 1938.270 ;
        RECT 2470.930 1935.490 2472.110 1936.670 ;
        RECT 2470.930 1757.090 2472.110 1758.270 ;
        RECT 2470.930 1755.490 2472.110 1756.670 ;
        RECT 2470.930 1577.090 2472.110 1578.270 ;
        RECT 2470.930 1575.490 2472.110 1576.670 ;
        RECT 2470.930 1397.090 2472.110 1398.270 ;
        RECT 2470.930 1395.490 2472.110 1396.670 ;
        RECT 2470.930 1217.090 2472.110 1218.270 ;
        RECT 2470.930 1215.490 2472.110 1216.670 ;
        RECT 2470.930 1037.090 2472.110 1038.270 ;
        RECT 2470.930 1035.490 2472.110 1036.670 ;
        RECT 2470.930 857.090 2472.110 858.270 ;
        RECT 2470.930 855.490 2472.110 856.670 ;
        RECT 2470.930 677.090 2472.110 678.270 ;
        RECT 2470.930 675.490 2472.110 676.670 ;
        RECT 2470.930 497.090 2472.110 498.270 ;
        RECT 2470.930 495.490 2472.110 496.670 ;
        RECT 2470.930 317.090 2472.110 318.270 ;
        RECT 2470.930 315.490 2472.110 316.670 ;
        RECT 2470.930 137.090 2472.110 138.270 ;
        RECT 2470.930 135.490 2472.110 136.670 ;
        RECT 2470.930 -26.410 2472.110 -25.230 ;
        RECT 2470.930 -28.010 2472.110 -26.830 ;
        RECT 2488.930 2135.090 2490.110 2136.270 ;
        RECT 2488.930 2133.490 2490.110 2134.670 ;
        RECT 2488.930 1955.090 2490.110 1956.270 ;
        RECT 2488.930 1953.490 2490.110 1954.670 ;
        RECT 2488.930 1775.090 2490.110 1776.270 ;
        RECT 2488.930 1773.490 2490.110 1774.670 ;
        RECT 2488.930 1595.090 2490.110 1596.270 ;
        RECT 2488.930 1593.490 2490.110 1594.670 ;
        RECT 2488.930 1415.090 2490.110 1416.270 ;
        RECT 2488.930 1413.490 2490.110 1414.670 ;
        RECT 2488.930 1235.090 2490.110 1236.270 ;
        RECT 2488.930 1233.490 2490.110 1234.670 ;
        RECT 2488.930 1055.090 2490.110 1056.270 ;
        RECT 2488.930 1053.490 2490.110 1054.670 ;
        RECT 2488.930 875.090 2490.110 876.270 ;
        RECT 2488.930 873.490 2490.110 874.670 ;
        RECT 2488.930 695.090 2490.110 696.270 ;
        RECT 2488.930 693.490 2490.110 694.670 ;
        RECT 2488.930 515.090 2490.110 516.270 ;
        RECT 2488.930 513.490 2490.110 514.670 ;
        RECT 2488.930 335.090 2490.110 336.270 ;
        RECT 2488.930 333.490 2490.110 334.670 ;
        RECT 2488.930 155.090 2490.110 156.270 ;
        RECT 2488.930 153.490 2490.110 154.670 ;
        RECT 2308.930 -35.810 2310.110 -34.630 ;
        RECT 2308.930 -37.410 2310.110 -36.230 ;
        RECT 2614.930 2261.090 2616.110 2262.270 ;
        RECT 2614.930 2259.490 2616.110 2260.670 ;
        RECT 2614.930 2081.090 2616.110 2082.270 ;
        RECT 2614.930 2079.490 2616.110 2080.670 ;
        RECT 2614.930 1901.090 2616.110 1902.270 ;
        RECT 2614.930 1899.490 2616.110 1900.670 ;
        RECT 2614.930 1721.090 2616.110 1722.270 ;
        RECT 2614.930 1719.490 2616.110 1720.670 ;
        RECT 2614.930 1541.090 2616.110 1542.270 ;
        RECT 2614.930 1539.490 2616.110 1540.670 ;
        RECT 2614.930 1361.090 2616.110 1362.270 ;
        RECT 2614.930 1359.490 2616.110 1360.670 ;
        RECT 2614.930 1181.090 2616.110 1182.270 ;
        RECT 2614.930 1179.490 2616.110 1180.670 ;
        RECT 2614.930 1001.090 2616.110 1002.270 ;
        RECT 2614.930 999.490 2616.110 1000.670 ;
        RECT 2614.930 821.090 2616.110 822.270 ;
        RECT 2614.930 819.490 2616.110 820.670 ;
        RECT 2614.930 641.090 2616.110 642.270 ;
        RECT 2614.930 639.490 2616.110 640.670 ;
        RECT 2614.930 461.090 2616.110 462.270 ;
        RECT 2614.930 459.490 2616.110 460.670 ;
        RECT 2614.930 281.090 2616.110 282.270 ;
        RECT 2614.930 279.490 2616.110 280.670 ;
        RECT 2614.930 101.090 2616.110 102.270 ;
        RECT 2614.930 99.490 2616.110 100.670 ;
        RECT 2614.930 -7.610 2616.110 -6.430 ;
        RECT 2614.930 -9.210 2616.110 -8.030 ;
        RECT 2632.930 3359.090 2634.110 3360.270 ;
        RECT 2632.930 3357.490 2634.110 3358.670 ;
        RECT 2632.930 3179.090 2634.110 3180.270 ;
        RECT 2632.930 3177.490 2634.110 3178.670 ;
        RECT 2632.930 2999.090 2634.110 3000.270 ;
        RECT 2632.930 2997.490 2634.110 2998.670 ;
        RECT 2632.930 2819.090 2634.110 2820.270 ;
        RECT 2632.930 2817.490 2634.110 2818.670 ;
        RECT 2632.930 2639.090 2634.110 2640.270 ;
        RECT 2632.930 2637.490 2634.110 2638.670 ;
        RECT 2632.930 2459.090 2634.110 2460.270 ;
        RECT 2632.930 2457.490 2634.110 2458.670 ;
        RECT 2632.930 2279.090 2634.110 2280.270 ;
        RECT 2632.930 2277.490 2634.110 2278.670 ;
        RECT 2632.930 2099.090 2634.110 2100.270 ;
        RECT 2632.930 2097.490 2634.110 2098.670 ;
        RECT 2632.930 1919.090 2634.110 1920.270 ;
        RECT 2632.930 1917.490 2634.110 1918.670 ;
        RECT 2632.930 1739.090 2634.110 1740.270 ;
        RECT 2632.930 1737.490 2634.110 1738.670 ;
        RECT 2632.930 1559.090 2634.110 1560.270 ;
        RECT 2632.930 1557.490 2634.110 1558.670 ;
        RECT 2632.930 1379.090 2634.110 1380.270 ;
        RECT 2632.930 1377.490 2634.110 1378.670 ;
        RECT 2632.930 1199.090 2634.110 1200.270 ;
        RECT 2632.930 1197.490 2634.110 1198.670 ;
        RECT 2632.930 1019.090 2634.110 1020.270 ;
        RECT 2632.930 1017.490 2634.110 1018.670 ;
        RECT 2632.930 839.090 2634.110 840.270 ;
        RECT 2632.930 837.490 2634.110 838.670 ;
        RECT 2632.930 659.090 2634.110 660.270 ;
        RECT 2632.930 657.490 2634.110 658.670 ;
        RECT 2632.930 479.090 2634.110 480.270 ;
        RECT 2632.930 477.490 2634.110 478.670 ;
        RECT 2632.930 299.090 2634.110 300.270 ;
        RECT 2632.930 297.490 2634.110 298.670 ;
        RECT 2632.930 119.090 2634.110 120.270 ;
        RECT 2632.930 117.490 2634.110 118.670 ;
        RECT 2632.930 -17.010 2634.110 -15.830 ;
        RECT 2632.930 -18.610 2634.110 -17.430 ;
        RECT 2650.930 3377.090 2652.110 3378.270 ;
        RECT 2650.930 3375.490 2652.110 3376.670 ;
        RECT 2650.930 3197.090 2652.110 3198.270 ;
        RECT 2650.930 3195.490 2652.110 3196.670 ;
        RECT 2650.930 3017.090 2652.110 3018.270 ;
        RECT 2650.930 3015.490 2652.110 3016.670 ;
        RECT 2650.930 2837.090 2652.110 2838.270 ;
        RECT 2650.930 2835.490 2652.110 2836.670 ;
        RECT 2650.930 2657.090 2652.110 2658.270 ;
        RECT 2650.930 2655.490 2652.110 2656.670 ;
        RECT 2650.930 2477.090 2652.110 2478.270 ;
        RECT 2650.930 2475.490 2652.110 2476.670 ;
        RECT 2650.930 2297.090 2652.110 2298.270 ;
        RECT 2650.930 2295.490 2652.110 2296.670 ;
        RECT 2650.930 2117.090 2652.110 2118.270 ;
        RECT 2650.930 2115.490 2652.110 2116.670 ;
        RECT 2650.930 1937.090 2652.110 1938.270 ;
        RECT 2650.930 1935.490 2652.110 1936.670 ;
        RECT 2650.930 1757.090 2652.110 1758.270 ;
        RECT 2650.930 1755.490 2652.110 1756.670 ;
        RECT 2650.930 1577.090 2652.110 1578.270 ;
        RECT 2650.930 1575.490 2652.110 1576.670 ;
        RECT 2650.930 1397.090 2652.110 1398.270 ;
        RECT 2650.930 1395.490 2652.110 1396.670 ;
        RECT 2650.930 1217.090 2652.110 1218.270 ;
        RECT 2650.930 1215.490 2652.110 1216.670 ;
        RECT 2650.930 1037.090 2652.110 1038.270 ;
        RECT 2650.930 1035.490 2652.110 1036.670 ;
        RECT 2650.930 857.090 2652.110 858.270 ;
        RECT 2650.930 855.490 2652.110 856.670 ;
        RECT 2650.930 677.090 2652.110 678.270 ;
        RECT 2650.930 675.490 2652.110 676.670 ;
        RECT 2650.930 497.090 2652.110 498.270 ;
        RECT 2650.930 495.490 2652.110 496.670 ;
        RECT 2650.930 317.090 2652.110 318.270 ;
        RECT 2650.930 315.490 2652.110 316.670 ;
        RECT 2650.930 137.090 2652.110 138.270 ;
        RECT 2650.930 135.490 2652.110 136.670 ;
        RECT 2650.930 -26.410 2652.110 -25.230 ;
        RECT 2650.930 -28.010 2652.110 -26.830 ;
        RECT 2848.930 3555.910 2850.110 3557.090 ;
        RECT 2848.930 3554.310 2850.110 3555.490 ;
        RECT 2830.930 3546.510 2832.110 3547.690 ;
        RECT 2830.930 3544.910 2832.110 3546.090 ;
        RECT 2812.930 3537.110 2814.110 3538.290 ;
        RECT 2812.930 3535.510 2814.110 3536.690 ;
        RECT 2668.930 3395.090 2670.110 3396.270 ;
        RECT 2668.930 3393.490 2670.110 3394.670 ;
        RECT 2668.930 3215.090 2670.110 3216.270 ;
        RECT 2668.930 3213.490 2670.110 3214.670 ;
        RECT 2668.930 3035.090 2670.110 3036.270 ;
        RECT 2668.930 3033.490 2670.110 3034.670 ;
        RECT 2668.930 2855.090 2670.110 2856.270 ;
        RECT 2668.930 2853.490 2670.110 2854.670 ;
        RECT 2668.930 2675.090 2670.110 2676.270 ;
        RECT 2668.930 2673.490 2670.110 2674.670 ;
        RECT 2668.930 2495.090 2670.110 2496.270 ;
        RECT 2668.930 2493.490 2670.110 2494.670 ;
        RECT 2668.930 2315.090 2670.110 2316.270 ;
        RECT 2668.930 2313.490 2670.110 2314.670 ;
        RECT 2668.930 2135.090 2670.110 2136.270 ;
        RECT 2668.930 2133.490 2670.110 2134.670 ;
        RECT 2668.930 1955.090 2670.110 1956.270 ;
        RECT 2668.930 1953.490 2670.110 1954.670 ;
        RECT 2668.930 1775.090 2670.110 1776.270 ;
        RECT 2668.930 1773.490 2670.110 1774.670 ;
        RECT 2668.930 1595.090 2670.110 1596.270 ;
        RECT 2668.930 1593.490 2670.110 1594.670 ;
        RECT 2668.930 1415.090 2670.110 1416.270 ;
        RECT 2668.930 1413.490 2670.110 1414.670 ;
        RECT 2668.930 1235.090 2670.110 1236.270 ;
        RECT 2668.930 1233.490 2670.110 1234.670 ;
        RECT 2668.930 1055.090 2670.110 1056.270 ;
        RECT 2668.930 1053.490 2670.110 1054.670 ;
        RECT 2668.930 875.090 2670.110 876.270 ;
        RECT 2668.930 873.490 2670.110 874.670 ;
        RECT 2668.930 695.090 2670.110 696.270 ;
        RECT 2668.930 693.490 2670.110 694.670 ;
        RECT 2668.930 515.090 2670.110 516.270 ;
        RECT 2668.930 513.490 2670.110 514.670 ;
        RECT 2668.930 335.090 2670.110 336.270 ;
        RECT 2668.930 333.490 2670.110 334.670 ;
        RECT 2668.930 155.090 2670.110 156.270 ;
        RECT 2668.930 153.490 2670.110 154.670 ;
        RECT 2488.930 -35.810 2490.110 -34.630 ;
        RECT 2488.930 -37.410 2490.110 -36.230 ;
        RECT 2794.930 3527.710 2796.110 3528.890 ;
        RECT 2794.930 3526.110 2796.110 3527.290 ;
        RECT 2794.930 3341.090 2796.110 3342.270 ;
        RECT 2794.930 3339.490 2796.110 3340.670 ;
        RECT 2794.930 3161.090 2796.110 3162.270 ;
        RECT 2794.930 3159.490 2796.110 3160.670 ;
        RECT 2794.930 2981.090 2796.110 2982.270 ;
        RECT 2794.930 2979.490 2796.110 2980.670 ;
        RECT 2794.930 2801.090 2796.110 2802.270 ;
        RECT 2794.930 2799.490 2796.110 2800.670 ;
        RECT 2794.930 2621.090 2796.110 2622.270 ;
        RECT 2794.930 2619.490 2796.110 2620.670 ;
        RECT 2794.930 2441.090 2796.110 2442.270 ;
        RECT 2794.930 2439.490 2796.110 2440.670 ;
        RECT 2794.930 2261.090 2796.110 2262.270 ;
        RECT 2794.930 2259.490 2796.110 2260.670 ;
        RECT 2794.930 2081.090 2796.110 2082.270 ;
        RECT 2794.930 2079.490 2796.110 2080.670 ;
        RECT 2794.930 1901.090 2796.110 1902.270 ;
        RECT 2794.930 1899.490 2796.110 1900.670 ;
        RECT 2794.930 1721.090 2796.110 1722.270 ;
        RECT 2794.930 1719.490 2796.110 1720.670 ;
        RECT 2794.930 1541.090 2796.110 1542.270 ;
        RECT 2794.930 1539.490 2796.110 1540.670 ;
        RECT 2794.930 1361.090 2796.110 1362.270 ;
        RECT 2794.930 1359.490 2796.110 1360.670 ;
        RECT 2794.930 1181.090 2796.110 1182.270 ;
        RECT 2794.930 1179.490 2796.110 1180.670 ;
        RECT 2794.930 1001.090 2796.110 1002.270 ;
        RECT 2794.930 999.490 2796.110 1000.670 ;
        RECT 2794.930 821.090 2796.110 822.270 ;
        RECT 2794.930 819.490 2796.110 820.670 ;
        RECT 2794.930 641.090 2796.110 642.270 ;
        RECT 2794.930 639.490 2796.110 640.670 ;
        RECT 2794.930 461.090 2796.110 462.270 ;
        RECT 2794.930 459.490 2796.110 460.670 ;
        RECT 2794.930 281.090 2796.110 282.270 ;
        RECT 2794.930 279.490 2796.110 280.670 ;
        RECT 2794.930 101.090 2796.110 102.270 ;
        RECT 2794.930 99.490 2796.110 100.670 ;
        RECT 2794.930 -7.610 2796.110 -6.430 ;
        RECT 2794.930 -9.210 2796.110 -8.030 ;
        RECT 2812.930 3359.090 2814.110 3360.270 ;
        RECT 2812.930 3357.490 2814.110 3358.670 ;
        RECT 2812.930 3179.090 2814.110 3180.270 ;
        RECT 2812.930 3177.490 2814.110 3178.670 ;
        RECT 2812.930 2999.090 2814.110 3000.270 ;
        RECT 2812.930 2997.490 2814.110 2998.670 ;
        RECT 2812.930 2819.090 2814.110 2820.270 ;
        RECT 2812.930 2817.490 2814.110 2818.670 ;
        RECT 2812.930 2639.090 2814.110 2640.270 ;
        RECT 2812.930 2637.490 2814.110 2638.670 ;
        RECT 2812.930 2459.090 2814.110 2460.270 ;
        RECT 2812.930 2457.490 2814.110 2458.670 ;
        RECT 2812.930 2279.090 2814.110 2280.270 ;
        RECT 2812.930 2277.490 2814.110 2278.670 ;
        RECT 2812.930 2099.090 2814.110 2100.270 ;
        RECT 2812.930 2097.490 2814.110 2098.670 ;
        RECT 2812.930 1919.090 2814.110 1920.270 ;
        RECT 2812.930 1917.490 2814.110 1918.670 ;
        RECT 2812.930 1739.090 2814.110 1740.270 ;
        RECT 2812.930 1737.490 2814.110 1738.670 ;
        RECT 2812.930 1559.090 2814.110 1560.270 ;
        RECT 2812.930 1557.490 2814.110 1558.670 ;
        RECT 2812.930 1379.090 2814.110 1380.270 ;
        RECT 2812.930 1377.490 2814.110 1378.670 ;
        RECT 2812.930 1199.090 2814.110 1200.270 ;
        RECT 2812.930 1197.490 2814.110 1198.670 ;
        RECT 2812.930 1019.090 2814.110 1020.270 ;
        RECT 2812.930 1017.490 2814.110 1018.670 ;
        RECT 2812.930 839.090 2814.110 840.270 ;
        RECT 2812.930 837.490 2814.110 838.670 ;
        RECT 2812.930 659.090 2814.110 660.270 ;
        RECT 2812.930 657.490 2814.110 658.670 ;
        RECT 2812.930 479.090 2814.110 480.270 ;
        RECT 2812.930 477.490 2814.110 478.670 ;
        RECT 2812.930 299.090 2814.110 300.270 ;
        RECT 2812.930 297.490 2814.110 298.670 ;
        RECT 2812.930 119.090 2814.110 120.270 ;
        RECT 2812.930 117.490 2814.110 118.670 ;
        RECT 2812.930 -17.010 2814.110 -15.830 ;
        RECT 2812.930 -18.610 2814.110 -17.430 ;
        RECT 2830.930 3377.090 2832.110 3378.270 ;
        RECT 2830.930 3375.490 2832.110 3376.670 ;
        RECT 2830.930 3197.090 2832.110 3198.270 ;
        RECT 2830.930 3195.490 2832.110 3196.670 ;
        RECT 2830.930 3017.090 2832.110 3018.270 ;
        RECT 2830.930 3015.490 2832.110 3016.670 ;
        RECT 2830.930 2837.090 2832.110 2838.270 ;
        RECT 2830.930 2835.490 2832.110 2836.670 ;
        RECT 2830.930 2657.090 2832.110 2658.270 ;
        RECT 2830.930 2655.490 2832.110 2656.670 ;
        RECT 2830.930 2477.090 2832.110 2478.270 ;
        RECT 2830.930 2475.490 2832.110 2476.670 ;
        RECT 2830.930 2297.090 2832.110 2298.270 ;
        RECT 2830.930 2295.490 2832.110 2296.670 ;
        RECT 2830.930 2117.090 2832.110 2118.270 ;
        RECT 2830.930 2115.490 2832.110 2116.670 ;
        RECT 2830.930 1937.090 2832.110 1938.270 ;
        RECT 2830.930 1935.490 2832.110 1936.670 ;
        RECT 2830.930 1757.090 2832.110 1758.270 ;
        RECT 2830.930 1755.490 2832.110 1756.670 ;
        RECT 2830.930 1577.090 2832.110 1578.270 ;
        RECT 2830.930 1575.490 2832.110 1576.670 ;
        RECT 2830.930 1397.090 2832.110 1398.270 ;
        RECT 2830.930 1395.490 2832.110 1396.670 ;
        RECT 2830.930 1217.090 2832.110 1218.270 ;
        RECT 2830.930 1215.490 2832.110 1216.670 ;
        RECT 2830.930 1037.090 2832.110 1038.270 ;
        RECT 2830.930 1035.490 2832.110 1036.670 ;
        RECT 2830.930 857.090 2832.110 858.270 ;
        RECT 2830.930 855.490 2832.110 856.670 ;
        RECT 2830.930 677.090 2832.110 678.270 ;
        RECT 2830.930 675.490 2832.110 676.670 ;
        RECT 2830.930 497.090 2832.110 498.270 ;
        RECT 2830.930 495.490 2832.110 496.670 ;
        RECT 2830.930 317.090 2832.110 318.270 ;
        RECT 2830.930 315.490 2832.110 316.670 ;
        RECT 2830.930 137.090 2832.110 138.270 ;
        RECT 2830.930 135.490 2832.110 136.670 ;
        RECT 2830.930 -26.410 2832.110 -25.230 ;
        RECT 2830.930 -28.010 2832.110 -26.830 ;
        RECT 2960.410 3555.910 2961.590 3557.090 ;
        RECT 2960.410 3554.310 2961.590 3555.490 ;
        RECT 2951.010 3546.510 2952.190 3547.690 ;
        RECT 2951.010 3544.910 2952.190 3546.090 ;
        RECT 2941.610 3537.110 2942.790 3538.290 ;
        RECT 2941.610 3535.510 2942.790 3536.690 ;
        RECT 2848.930 3395.090 2850.110 3396.270 ;
        RECT 2848.930 3393.490 2850.110 3394.670 ;
        RECT 2848.930 3215.090 2850.110 3216.270 ;
        RECT 2848.930 3213.490 2850.110 3214.670 ;
        RECT 2848.930 3035.090 2850.110 3036.270 ;
        RECT 2848.930 3033.490 2850.110 3034.670 ;
        RECT 2848.930 2855.090 2850.110 2856.270 ;
        RECT 2848.930 2853.490 2850.110 2854.670 ;
        RECT 2848.930 2675.090 2850.110 2676.270 ;
        RECT 2848.930 2673.490 2850.110 2674.670 ;
        RECT 2848.930 2495.090 2850.110 2496.270 ;
        RECT 2848.930 2493.490 2850.110 2494.670 ;
        RECT 2848.930 2315.090 2850.110 2316.270 ;
        RECT 2848.930 2313.490 2850.110 2314.670 ;
        RECT 2848.930 2135.090 2850.110 2136.270 ;
        RECT 2848.930 2133.490 2850.110 2134.670 ;
        RECT 2848.930 1955.090 2850.110 1956.270 ;
        RECT 2848.930 1953.490 2850.110 1954.670 ;
        RECT 2848.930 1775.090 2850.110 1776.270 ;
        RECT 2848.930 1773.490 2850.110 1774.670 ;
        RECT 2848.930 1595.090 2850.110 1596.270 ;
        RECT 2848.930 1593.490 2850.110 1594.670 ;
        RECT 2848.930 1415.090 2850.110 1416.270 ;
        RECT 2848.930 1413.490 2850.110 1414.670 ;
        RECT 2848.930 1235.090 2850.110 1236.270 ;
        RECT 2848.930 1233.490 2850.110 1234.670 ;
        RECT 2848.930 1055.090 2850.110 1056.270 ;
        RECT 2848.930 1053.490 2850.110 1054.670 ;
        RECT 2848.930 875.090 2850.110 876.270 ;
        RECT 2848.930 873.490 2850.110 874.670 ;
        RECT 2848.930 695.090 2850.110 696.270 ;
        RECT 2848.930 693.490 2850.110 694.670 ;
        RECT 2848.930 515.090 2850.110 516.270 ;
        RECT 2848.930 513.490 2850.110 514.670 ;
        RECT 2848.930 335.090 2850.110 336.270 ;
        RECT 2848.930 333.490 2850.110 334.670 ;
        RECT 2848.930 155.090 2850.110 156.270 ;
        RECT 2848.930 153.490 2850.110 154.670 ;
        RECT 2668.930 -35.810 2670.110 -34.630 ;
        RECT 2668.930 -37.410 2670.110 -36.230 ;
        RECT 2932.210 3527.710 2933.390 3528.890 ;
        RECT 2932.210 3526.110 2933.390 3527.290 ;
        RECT 2932.210 3341.090 2933.390 3342.270 ;
        RECT 2932.210 3339.490 2933.390 3340.670 ;
        RECT 2932.210 3161.090 2933.390 3162.270 ;
        RECT 2932.210 3159.490 2933.390 3160.670 ;
        RECT 2932.210 2981.090 2933.390 2982.270 ;
        RECT 2932.210 2979.490 2933.390 2980.670 ;
        RECT 2932.210 2801.090 2933.390 2802.270 ;
        RECT 2932.210 2799.490 2933.390 2800.670 ;
        RECT 2932.210 2621.090 2933.390 2622.270 ;
        RECT 2932.210 2619.490 2933.390 2620.670 ;
        RECT 2932.210 2441.090 2933.390 2442.270 ;
        RECT 2932.210 2439.490 2933.390 2440.670 ;
        RECT 2932.210 2261.090 2933.390 2262.270 ;
        RECT 2932.210 2259.490 2933.390 2260.670 ;
        RECT 2932.210 2081.090 2933.390 2082.270 ;
        RECT 2932.210 2079.490 2933.390 2080.670 ;
        RECT 2932.210 1901.090 2933.390 1902.270 ;
        RECT 2932.210 1899.490 2933.390 1900.670 ;
        RECT 2932.210 1721.090 2933.390 1722.270 ;
        RECT 2932.210 1719.490 2933.390 1720.670 ;
        RECT 2932.210 1541.090 2933.390 1542.270 ;
        RECT 2932.210 1539.490 2933.390 1540.670 ;
        RECT 2932.210 1361.090 2933.390 1362.270 ;
        RECT 2932.210 1359.490 2933.390 1360.670 ;
        RECT 2932.210 1181.090 2933.390 1182.270 ;
        RECT 2932.210 1179.490 2933.390 1180.670 ;
        RECT 2932.210 1001.090 2933.390 1002.270 ;
        RECT 2932.210 999.490 2933.390 1000.670 ;
        RECT 2932.210 821.090 2933.390 822.270 ;
        RECT 2932.210 819.490 2933.390 820.670 ;
        RECT 2932.210 641.090 2933.390 642.270 ;
        RECT 2932.210 639.490 2933.390 640.670 ;
        RECT 2932.210 461.090 2933.390 462.270 ;
        RECT 2932.210 459.490 2933.390 460.670 ;
        RECT 2932.210 281.090 2933.390 282.270 ;
        RECT 2932.210 279.490 2933.390 280.670 ;
        RECT 2932.210 101.090 2933.390 102.270 ;
        RECT 2932.210 99.490 2933.390 100.670 ;
        RECT 2932.210 -7.610 2933.390 -6.430 ;
        RECT 2932.210 -9.210 2933.390 -8.030 ;
        RECT 2941.610 3359.090 2942.790 3360.270 ;
        RECT 2941.610 3357.490 2942.790 3358.670 ;
        RECT 2941.610 3179.090 2942.790 3180.270 ;
        RECT 2941.610 3177.490 2942.790 3178.670 ;
        RECT 2941.610 2999.090 2942.790 3000.270 ;
        RECT 2941.610 2997.490 2942.790 2998.670 ;
        RECT 2941.610 2819.090 2942.790 2820.270 ;
        RECT 2941.610 2817.490 2942.790 2818.670 ;
        RECT 2941.610 2639.090 2942.790 2640.270 ;
        RECT 2941.610 2637.490 2942.790 2638.670 ;
        RECT 2941.610 2459.090 2942.790 2460.270 ;
        RECT 2941.610 2457.490 2942.790 2458.670 ;
        RECT 2941.610 2279.090 2942.790 2280.270 ;
        RECT 2941.610 2277.490 2942.790 2278.670 ;
        RECT 2941.610 2099.090 2942.790 2100.270 ;
        RECT 2941.610 2097.490 2942.790 2098.670 ;
        RECT 2941.610 1919.090 2942.790 1920.270 ;
        RECT 2941.610 1917.490 2942.790 1918.670 ;
        RECT 2941.610 1739.090 2942.790 1740.270 ;
        RECT 2941.610 1737.490 2942.790 1738.670 ;
        RECT 2941.610 1559.090 2942.790 1560.270 ;
        RECT 2941.610 1557.490 2942.790 1558.670 ;
        RECT 2941.610 1379.090 2942.790 1380.270 ;
        RECT 2941.610 1377.490 2942.790 1378.670 ;
        RECT 2941.610 1199.090 2942.790 1200.270 ;
        RECT 2941.610 1197.490 2942.790 1198.670 ;
        RECT 2941.610 1019.090 2942.790 1020.270 ;
        RECT 2941.610 1017.490 2942.790 1018.670 ;
        RECT 2941.610 839.090 2942.790 840.270 ;
        RECT 2941.610 837.490 2942.790 838.670 ;
        RECT 2941.610 659.090 2942.790 660.270 ;
        RECT 2941.610 657.490 2942.790 658.670 ;
        RECT 2941.610 479.090 2942.790 480.270 ;
        RECT 2941.610 477.490 2942.790 478.670 ;
        RECT 2941.610 299.090 2942.790 300.270 ;
        RECT 2941.610 297.490 2942.790 298.670 ;
        RECT 2941.610 119.090 2942.790 120.270 ;
        RECT 2941.610 117.490 2942.790 118.670 ;
        RECT 2941.610 -17.010 2942.790 -15.830 ;
        RECT 2941.610 -18.610 2942.790 -17.430 ;
        RECT 2951.010 3377.090 2952.190 3378.270 ;
        RECT 2951.010 3375.490 2952.190 3376.670 ;
        RECT 2951.010 3197.090 2952.190 3198.270 ;
        RECT 2951.010 3195.490 2952.190 3196.670 ;
        RECT 2951.010 3017.090 2952.190 3018.270 ;
        RECT 2951.010 3015.490 2952.190 3016.670 ;
        RECT 2951.010 2837.090 2952.190 2838.270 ;
        RECT 2951.010 2835.490 2952.190 2836.670 ;
        RECT 2951.010 2657.090 2952.190 2658.270 ;
        RECT 2951.010 2655.490 2952.190 2656.670 ;
        RECT 2951.010 2477.090 2952.190 2478.270 ;
        RECT 2951.010 2475.490 2952.190 2476.670 ;
        RECT 2951.010 2297.090 2952.190 2298.270 ;
        RECT 2951.010 2295.490 2952.190 2296.670 ;
        RECT 2951.010 2117.090 2952.190 2118.270 ;
        RECT 2951.010 2115.490 2952.190 2116.670 ;
        RECT 2951.010 1937.090 2952.190 1938.270 ;
        RECT 2951.010 1935.490 2952.190 1936.670 ;
        RECT 2951.010 1757.090 2952.190 1758.270 ;
        RECT 2951.010 1755.490 2952.190 1756.670 ;
        RECT 2951.010 1577.090 2952.190 1578.270 ;
        RECT 2951.010 1575.490 2952.190 1576.670 ;
        RECT 2951.010 1397.090 2952.190 1398.270 ;
        RECT 2951.010 1395.490 2952.190 1396.670 ;
        RECT 2951.010 1217.090 2952.190 1218.270 ;
        RECT 2951.010 1215.490 2952.190 1216.670 ;
        RECT 2951.010 1037.090 2952.190 1038.270 ;
        RECT 2951.010 1035.490 2952.190 1036.670 ;
        RECT 2951.010 857.090 2952.190 858.270 ;
        RECT 2951.010 855.490 2952.190 856.670 ;
        RECT 2951.010 677.090 2952.190 678.270 ;
        RECT 2951.010 675.490 2952.190 676.670 ;
        RECT 2951.010 497.090 2952.190 498.270 ;
        RECT 2951.010 495.490 2952.190 496.670 ;
        RECT 2951.010 317.090 2952.190 318.270 ;
        RECT 2951.010 315.490 2952.190 316.670 ;
        RECT 2951.010 137.090 2952.190 138.270 ;
        RECT 2951.010 135.490 2952.190 136.670 ;
        RECT 2951.010 -26.410 2952.190 -25.230 ;
        RECT 2951.010 -28.010 2952.190 -26.830 ;
        RECT 2960.410 3395.090 2961.590 3396.270 ;
        RECT 2960.410 3393.490 2961.590 3394.670 ;
        RECT 2960.410 3215.090 2961.590 3216.270 ;
        RECT 2960.410 3213.490 2961.590 3214.670 ;
        RECT 2960.410 3035.090 2961.590 3036.270 ;
        RECT 2960.410 3033.490 2961.590 3034.670 ;
        RECT 2960.410 2855.090 2961.590 2856.270 ;
        RECT 2960.410 2853.490 2961.590 2854.670 ;
        RECT 2960.410 2675.090 2961.590 2676.270 ;
        RECT 2960.410 2673.490 2961.590 2674.670 ;
        RECT 2960.410 2495.090 2961.590 2496.270 ;
        RECT 2960.410 2493.490 2961.590 2494.670 ;
        RECT 2960.410 2315.090 2961.590 2316.270 ;
        RECT 2960.410 2313.490 2961.590 2314.670 ;
        RECT 2960.410 2135.090 2961.590 2136.270 ;
        RECT 2960.410 2133.490 2961.590 2134.670 ;
        RECT 2960.410 1955.090 2961.590 1956.270 ;
        RECT 2960.410 1953.490 2961.590 1954.670 ;
        RECT 2960.410 1775.090 2961.590 1776.270 ;
        RECT 2960.410 1773.490 2961.590 1774.670 ;
        RECT 2960.410 1595.090 2961.590 1596.270 ;
        RECT 2960.410 1593.490 2961.590 1594.670 ;
        RECT 2960.410 1415.090 2961.590 1416.270 ;
        RECT 2960.410 1413.490 2961.590 1414.670 ;
        RECT 2960.410 1235.090 2961.590 1236.270 ;
        RECT 2960.410 1233.490 2961.590 1234.670 ;
        RECT 2960.410 1055.090 2961.590 1056.270 ;
        RECT 2960.410 1053.490 2961.590 1054.670 ;
        RECT 2960.410 875.090 2961.590 876.270 ;
        RECT 2960.410 873.490 2961.590 874.670 ;
        RECT 2960.410 695.090 2961.590 696.270 ;
        RECT 2960.410 693.490 2961.590 694.670 ;
        RECT 2960.410 515.090 2961.590 516.270 ;
        RECT 2960.410 513.490 2961.590 514.670 ;
        RECT 2960.410 335.090 2961.590 336.270 ;
        RECT 2960.410 333.490 2961.590 334.670 ;
        RECT 2960.410 155.090 2961.590 156.270 ;
        RECT 2960.410 153.490 2961.590 154.670 ;
        RECT 2848.930 -35.810 2850.110 -34.630 ;
        RECT 2848.930 -37.410 2850.110 -36.230 ;
        RECT 2960.410 -35.810 2961.590 -34.630 ;
        RECT 2960.410 -37.410 2961.590 -36.230 ;
      LAYER met5 ;
        RECT -42.880 3557.200 -39.880 3557.210 ;
        RECT 148.020 3557.200 151.020 3557.210 ;
        RECT 328.020 3557.200 331.020 3557.210 ;
        RECT 508.020 3557.200 511.020 3557.210 ;
        RECT 688.020 3557.200 691.020 3557.210 ;
        RECT 868.020 3557.200 871.020 3557.210 ;
        RECT 1048.020 3557.200 1051.020 3557.210 ;
        RECT 1228.020 3557.200 1231.020 3557.210 ;
        RECT 1408.020 3557.200 1411.020 3557.210 ;
        RECT 1588.020 3557.200 1591.020 3557.210 ;
        RECT 1768.020 3557.200 1771.020 3557.210 ;
        RECT 1948.020 3557.200 1951.020 3557.210 ;
        RECT 2128.020 3557.200 2131.020 3557.210 ;
        RECT 2308.020 3557.200 2311.020 3557.210 ;
        RECT 2488.020 3557.200 2491.020 3557.210 ;
        RECT 2668.020 3557.200 2671.020 3557.210 ;
        RECT 2848.020 3557.200 2851.020 3557.210 ;
        RECT 2959.500 3557.200 2962.500 3557.210 ;
        RECT -42.880 3554.200 2962.500 3557.200 ;
        RECT -42.880 3554.190 -39.880 3554.200 ;
        RECT 148.020 3554.190 151.020 3554.200 ;
        RECT 328.020 3554.190 331.020 3554.200 ;
        RECT 508.020 3554.190 511.020 3554.200 ;
        RECT 688.020 3554.190 691.020 3554.200 ;
        RECT 868.020 3554.190 871.020 3554.200 ;
        RECT 1048.020 3554.190 1051.020 3554.200 ;
        RECT 1228.020 3554.190 1231.020 3554.200 ;
        RECT 1408.020 3554.190 1411.020 3554.200 ;
        RECT 1588.020 3554.190 1591.020 3554.200 ;
        RECT 1768.020 3554.190 1771.020 3554.200 ;
        RECT 1948.020 3554.190 1951.020 3554.200 ;
        RECT 2128.020 3554.190 2131.020 3554.200 ;
        RECT 2308.020 3554.190 2311.020 3554.200 ;
        RECT 2488.020 3554.190 2491.020 3554.200 ;
        RECT 2668.020 3554.190 2671.020 3554.200 ;
        RECT 2848.020 3554.190 2851.020 3554.200 ;
        RECT 2959.500 3554.190 2962.500 3554.200 ;
        RECT -33.480 3547.800 -30.480 3547.810 ;
        RECT 130.020 3547.800 133.020 3547.810 ;
        RECT 310.020 3547.800 313.020 3547.810 ;
        RECT 490.020 3547.800 493.020 3547.810 ;
        RECT 670.020 3547.800 673.020 3547.810 ;
        RECT 850.020 3547.800 853.020 3547.810 ;
        RECT 1030.020 3547.800 1033.020 3547.810 ;
        RECT 1210.020 3547.800 1213.020 3547.810 ;
        RECT 1390.020 3547.800 1393.020 3547.810 ;
        RECT 1570.020 3547.800 1573.020 3547.810 ;
        RECT 1750.020 3547.800 1753.020 3547.810 ;
        RECT 1930.020 3547.800 1933.020 3547.810 ;
        RECT 2110.020 3547.800 2113.020 3547.810 ;
        RECT 2290.020 3547.800 2293.020 3547.810 ;
        RECT 2470.020 3547.800 2473.020 3547.810 ;
        RECT 2650.020 3547.800 2653.020 3547.810 ;
        RECT 2830.020 3547.800 2833.020 3547.810 ;
        RECT 2950.100 3547.800 2953.100 3547.810 ;
        RECT -33.480 3544.800 2953.100 3547.800 ;
        RECT -33.480 3544.790 -30.480 3544.800 ;
        RECT 130.020 3544.790 133.020 3544.800 ;
        RECT 310.020 3544.790 313.020 3544.800 ;
        RECT 490.020 3544.790 493.020 3544.800 ;
        RECT 670.020 3544.790 673.020 3544.800 ;
        RECT 850.020 3544.790 853.020 3544.800 ;
        RECT 1030.020 3544.790 1033.020 3544.800 ;
        RECT 1210.020 3544.790 1213.020 3544.800 ;
        RECT 1390.020 3544.790 1393.020 3544.800 ;
        RECT 1570.020 3544.790 1573.020 3544.800 ;
        RECT 1750.020 3544.790 1753.020 3544.800 ;
        RECT 1930.020 3544.790 1933.020 3544.800 ;
        RECT 2110.020 3544.790 2113.020 3544.800 ;
        RECT 2290.020 3544.790 2293.020 3544.800 ;
        RECT 2470.020 3544.790 2473.020 3544.800 ;
        RECT 2650.020 3544.790 2653.020 3544.800 ;
        RECT 2830.020 3544.790 2833.020 3544.800 ;
        RECT 2950.100 3544.790 2953.100 3544.800 ;
        RECT -24.080 3538.400 -21.080 3538.410 ;
        RECT 112.020 3538.400 115.020 3538.410 ;
        RECT 292.020 3538.400 295.020 3538.410 ;
        RECT 472.020 3538.400 475.020 3538.410 ;
        RECT 652.020 3538.400 655.020 3538.410 ;
        RECT 832.020 3538.400 835.020 3538.410 ;
        RECT 1012.020 3538.400 1015.020 3538.410 ;
        RECT 1192.020 3538.400 1195.020 3538.410 ;
        RECT 1372.020 3538.400 1375.020 3538.410 ;
        RECT 1552.020 3538.400 1555.020 3538.410 ;
        RECT 1732.020 3538.400 1735.020 3538.410 ;
        RECT 1912.020 3538.400 1915.020 3538.410 ;
        RECT 2092.020 3538.400 2095.020 3538.410 ;
        RECT 2272.020 3538.400 2275.020 3538.410 ;
        RECT 2452.020 3538.400 2455.020 3538.410 ;
        RECT 2632.020 3538.400 2635.020 3538.410 ;
        RECT 2812.020 3538.400 2815.020 3538.410 ;
        RECT 2940.700 3538.400 2943.700 3538.410 ;
        RECT -24.080 3535.400 2943.700 3538.400 ;
        RECT -24.080 3535.390 -21.080 3535.400 ;
        RECT 112.020 3535.390 115.020 3535.400 ;
        RECT 292.020 3535.390 295.020 3535.400 ;
        RECT 472.020 3535.390 475.020 3535.400 ;
        RECT 652.020 3535.390 655.020 3535.400 ;
        RECT 832.020 3535.390 835.020 3535.400 ;
        RECT 1012.020 3535.390 1015.020 3535.400 ;
        RECT 1192.020 3535.390 1195.020 3535.400 ;
        RECT 1372.020 3535.390 1375.020 3535.400 ;
        RECT 1552.020 3535.390 1555.020 3535.400 ;
        RECT 1732.020 3535.390 1735.020 3535.400 ;
        RECT 1912.020 3535.390 1915.020 3535.400 ;
        RECT 2092.020 3535.390 2095.020 3535.400 ;
        RECT 2272.020 3535.390 2275.020 3535.400 ;
        RECT 2452.020 3535.390 2455.020 3535.400 ;
        RECT 2632.020 3535.390 2635.020 3535.400 ;
        RECT 2812.020 3535.390 2815.020 3535.400 ;
        RECT 2940.700 3535.390 2943.700 3535.400 ;
        RECT -14.680 3529.000 -11.680 3529.010 ;
        RECT 94.020 3529.000 97.020 3529.010 ;
        RECT 274.020 3529.000 277.020 3529.010 ;
        RECT 454.020 3529.000 457.020 3529.010 ;
        RECT 634.020 3529.000 637.020 3529.010 ;
        RECT 814.020 3529.000 817.020 3529.010 ;
        RECT 994.020 3529.000 997.020 3529.010 ;
        RECT 1174.020 3529.000 1177.020 3529.010 ;
        RECT 1354.020 3529.000 1357.020 3529.010 ;
        RECT 1534.020 3529.000 1537.020 3529.010 ;
        RECT 1714.020 3529.000 1717.020 3529.010 ;
        RECT 1894.020 3529.000 1897.020 3529.010 ;
        RECT 2074.020 3529.000 2077.020 3529.010 ;
        RECT 2254.020 3529.000 2257.020 3529.010 ;
        RECT 2434.020 3529.000 2437.020 3529.010 ;
        RECT 2614.020 3529.000 2617.020 3529.010 ;
        RECT 2794.020 3529.000 2797.020 3529.010 ;
        RECT 2931.300 3529.000 2934.300 3529.010 ;
        RECT -14.680 3526.000 2934.300 3529.000 ;
        RECT -14.680 3525.990 -11.680 3526.000 ;
        RECT 94.020 3525.990 97.020 3526.000 ;
        RECT 274.020 3525.990 277.020 3526.000 ;
        RECT 454.020 3525.990 457.020 3526.000 ;
        RECT 634.020 3525.990 637.020 3526.000 ;
        RECT 814.020 3525.990 817.020 3526.000 ;
        RECT 994.020 3525.990 997.020 3526.000 ;
        RECT 1174.020 3525.990 1177.020 3526.000 ;
        RECT 1354.020 3525.990 1357.020 3526.000 ;
        RECT 1534.020 3525.990 1537.020 3526.000 ;
        RECT 1714.020 3525.990 1717.020 3526.000 ;
        RECT 1894.020 3525.990 1897.020 3526.000 ;
        RECT 2074.020 3525.990 2077.020 3526.000 ;
        RECT 2254.020 3525.990 2257.020 3526.000 ;
        RECT 2434.020 3525.990 2437.020 3526.000 ;
        RECT 2614.020 3525.990 2617.020 3526.000 ;
        RECT 2794.020 3525.990 2797.020 3526.000 ;
        RECT 2931.300 3525.990 2934.300 3526.000 ;
        RECT -42.880 3396.380 -39.880 3396.390 ;
        RECT 148.020 3396.380 151.020 3396.390 ;
        RECT 328.020 3396.380 331.020 3396.390 ;
        RECT 508.020 3396.380 511.020 3396.390 ;
        RECT 688.020 3396.380 691.020 3396.390 ;
        RECT 868.020 3396.380 871.020 3396.390 ;
        RECT 1048.020 3396.380 1051.020 3396.390 ;
        RECT 1228.020 3396.380 1231.020 3396.390 ;
        RECT 1408.020 3396.380 1411.020 3396.390 ;
        RECT 1588.020 3396.380 1591.020 3396.390 ;
        RECT 1768.020 3396.380 1771.020 3396.390 ;
        RECT 1948.020 3396.380 1951.020 3396.390 ;
        RECT 2128.020 3396.380 2131.020 3396.390 ;
        RECT 2308.020 3396.380 2311.020 3396.390 ;
        RECT 2488.020 3396.380 2491.020 3396.390 ;
        RECT 2668.020 3396.380 2671.020 3396.390 ;
        RECT 2848.020 3396.380 2851.020 3396.390 ;
        RECT 2959.500 3396.380 2962.500 3396.390 ;
        RECT -42.880 3393.380 2962.500 3396.380 ;
        RECT -42.880 3393.370 -39.880 3393.380 ;
        RECT 148.020 3393.370 151.020 3393.380 ;
        RECT 328.020 3393.370 331.020 3393.380 ;
        RECT 508.020 3393.370 511.020 3393.380 ;
        RECT 688.020 3393.370 691.020 3393.380 ;
        RECT 868.020 3393.370 871.020 3393.380 ;
        RECT 1048.020 3393.370 1051.020 3393.380 ;
        RECT 1228.020 3393.370 1231.020 3393.380 ;
        RECT 1408.020 3393.370 1411.020 3393.380 ;
        RECT 1588.020 3393.370 1591.020 3393.380 ;
        RECT 1768.020 3393.370 1771.020 3393.380 ;
        RECT 1948.020 3393.370 1951.020 3393.380 ;
        RECT 2128.020 3393.370 2131.020 3393.380 ;
        RECT 2308.020 3393.370 2311.020 3393.380 ;
        RECT 2488.020 3393.370 2491.020 3393.380 ;
        RECT 2668.020 3393.370 2671.020 3393.380 ;
        RECT 2848.020 3393.370 2851.020 3393.380 ;
        RECT 2959.500 3393.370 2962.500 3393.380 ;
        RECT -33.480 3378.380 -30.480 3378.390 ;
        RECT 130.020 3378.380 133.020 3378.390 ;
        RECT 310.020 3378.380 313.020 3378.390 ;
        RECT 490.020 3378.380 493.020 3378.390 ;
        RECT 670.020 3378.380 673.020 3378.390 ;
        RECT 850.020 3378.380 853.020 3378.390 ;
        RECT 1030.020 3378.380 1033.020 3378.390 ;
        RECT 1210.020 3378.380 1213.020 3378.390 ;
        RECT 1390.020 3378.380 1393.020 3378.390 ;
        RECT 1570.020 3378.380 1573.020 3378.390 ;
        RECT 1750.020 3378.380 1753.020 3378.390 ;
        RECT 1930.020 3378.380 1933.020 3378.390 ;
        RECT 2110.020 3378.380 2113.020 3378.390 ;
        RECT 2290.020 3378.380 2293.020 3378.390 ;
        RECT 2470.020 3378.380 2473.020 3378.390 ;
        RECT 2650.020 3378.380 2653.020 3378.390 ;
        RECT 2830.020 3378.380 2833.020 3378.390 ;
        RECT 2950.100 3378.380 2953.100 3378.390 ;
        RECT -33.480 3375.380 2953.100 3378.380 ;
        RECT -33.480 3375.370 -30.480 3375.380 ;
        RECT 130.020 3375.370 133.020 3375.380 ;
        RECT 310.020 3375.370 313.020 3375.380 ;
        RECT 490.020 3375.370 493.020 3375.380 ;
        RECT 670.020 3375.370 673.020 3375.380 ;
        RECT 850.020 3375.370 853.020 3375.380 ;
        RECT 1030.020 3375.370 1033.020 3375.380 ;
        RECT 1210.020 3375.370 1213.020 3375.380 ;
        RECT 1390.020 3375.370 1393.020 3375.380 ;
        RECT 1570.020 3375.370 1573.020 3375.380 ;
        RECT 1750.020 3375.370 1753.020 3375.380 ;
        RECT 1930.020 3375.370 1933.020 3375.380 ;
        RECT 2110.020 3375.370 2113.020 3375.380 ;
        RECT 2290.020 3375.370 2293.020 3375.380 ;
        RECT 2470.020 3375.370 2473.020 3375.380 ;
        RECT 2650.020 3375.370 2653.020 3375.380 ;
        RECT 2830.020 3375.370 2833.020 3375.380 ;
        RECT 2950.100 3375.370 2953.100 3375.380 ;
        RECT -24.080 3360.380 -21.080 3360.390 ;
        RECT 112.020 3360.380 115.020 3360.390 ;
        RECT 292.020 3360.380 295.020 3360.390 ;
        RECT 472.020 3360.380 475.020 3360.390 ;
        RECT 652.020 3360.380 655.020 3360.390 ;
        RECT 832.020 3360.380 835.020 3360.390 ;
        RECT 1012.020 3360.380 1015.020 3360.390 ;
        RECT 1192.020 3360.380 1195.020 3360.390 ;
        RECT 1372.020 3360.380 1375.020 3360.390 ;
        RECT 1552.020 3360.380 1555.020 3360.390 ;
        RECT 1732.020 3360.380 1735.020 3360.390 ;
        RECT 1912.020 3360.380 1915.020 3360.390 ;
        RECT 2092.020 3360.380 2095.020 3360.390 ;
        RECT 2272.020 3360.380 2275.020 3360.390 ;
        RECT 2452.020 3360.380 2455.020 3360.390 ;
        RECT 2632.020 3360.380 2635.020 3360.390 ;
        RECT 2812.020 3360.380 2815.020 3360.390 ;
        RECT 2940.700 3360.380 2943.700 3360.390 ;
        RECT -24.080 3357.380 2943.700 3360.380 ;
        RECT -24.080 3357.370 -21.080 3357.380 ;
        RECT 112.020 3357.370 115.020 3357.380 ;
        RECT 292.020 3357.370 295.020 3357.380 ;
        RECT 472.020 3357.370 475.020 3357.380 ;
        RECT 652.020 3357.370 655.020 3357.380 ;
        RECT 832.020 3357.370 835.020 3357.380 ;
        RECT 1012.020 3357.370 1015.020 3357.380 ;
        RECT 1192.020 3357.370 1195.020 3357.380 ;
        RECT 1372.020 3357.370 1375.020 3357.380 ;
        RECT 1552.020 3357.370 1555.020 3357.380 ;
        RECT 1732.020 3357.370 1735.020 3357.380 ;
        RECT 1912.020 3357.370 1915.020 3357.380 ;
        RECT 2092.020 3357.370 2095.020 3357.380 ;
        RECT 2272.020 3357.370 2275.020 3357.380 ;
        RECT 2452.020 3357.370 2455.020 3357.380 ;
        RECT 2632.020 3357.370 2635.020 3357.380 ;
        RECT 2812.020 3357.370 2815.020 3357.380 ;
        RECT 2940.700 3357.370 2943.700 3357.380 ;
        RECT -14.680 3342.380 -11.680 3342.390 ;
        RECT 94.020 3342.380 97.020 3342.390 ;
        RECT 274.020 3342.380 277.020 3342.390 ;
        RECT 454.020 3342.380 457.020 3342.390 ;
        RECT 634.020 3342.380 637.020 3342.390 ;
        RECT 814.020 3342.380 817.020 3342.390 ;
        RECT 994.020 3342.380 997.020 3342.390 ;
        RECT 1174.020 3342.380 1177.020 3342.390 ;
        RECT 1354.020 3342.380 1357.020 3342.390 ;
        RECT 1534.020 3342.380 1537.020 3342.390 ;
        RECT 1714.020 3342.380 1717.020 3342.390 ;
        RECT 1894.020 3342.380 1897.020 3342.390 ;
        RECT 2074.020 3342.380 2077.020 3342.390 ;
        RECT 2254.020 3342.380 2257.020 3342.390 ;
        RECT 2434.020 3342.380 2437.020 3342.390 ;
        RECT 2614.020 3342.380 2617.020 3342.390 ;
        RECT 2794.020 3342.380 2797.020 3342.390 ;
        RECT 2931.300 3342.380 2934.300 3342.390 ;
        RECT -14.680 3339.380 2934.300 3342.380 ;
        RECT -14.680 3339.370 -11.680 3339.380 ;
        RECT 94.020 3339.370 97.020 3339.380 ;
        RECT 274.020 3339.370 277.020 3339.380 ;
        RECT 454.020 3339.370 457.020 3339.380 ;
        RECT 634.020 3339.370 637.020 3339.380 ;
        RECT 814.020 3339.370 817.020 3339.380 ;
        RECT 994.020 3339.370 997.020 3339.380 ;
        RECT 1174.020 3339.370 1177.020 3339.380 ;
        RECT 1354.020 3339.370 1357.020 3339.380 ;
        RECT 1534.020 3339.370 1537.020 3339.380 ;
        RECT 1714.020 3339.370 1717.020 3339.380 ;
        RECT 1894.020 3339.370 1897.020 3339.380 ;
        RECT 2074.020 3339.370 2077.020 3339.380 ;
        RECT 2254.020 3339.370 2257.020 3339.380 ;
        RECT 2434.020 3339.370 2437.020 3339.380 ;
        RECT 2614.020 3339.370 2617.020 3339.380 ;
        RECT 2794.020 3339.370 2797.020 3339.380 ;
        RECT 2931.300 3339.370 2934.300 3339.380 ;
        RECT -42.880 3216.380 -39.880 3216.390 ;
        RECT 148.020 3216.380 151.020 3216.390 ;
        RECT 328.020 3216.380 331.020 3216.390 ;
        RECT 508.020 3216.380 511.020 3216.390 ;
        RECT 688.020 3216.380 691.020 3216.390 ;
        RECT 868.020 3216.380 871.020 3216.390 ;
        RECT 1048.020 3216.380 1051.020 3216.390 ;
        RECT 1228.020 3216.380 1231.020 3216.390 ;
        RECT 1408.020 3216.380 1411.020 3216.390 ;
        RECT 1588.020 3216.380 1591.020 3216.390 ;
        RECT 1768.020 3216.380 1771.020 3216.390 ;
        RECT 1948.020 3216.380 1951.020 3216.390 ;
        RECT 2128.020 3216.380 2131.020 3216.390 ;
        RECT 2308.020 3216.380 2311.020 3216.390 ;
        RECT 2488.020 3216.380 2491.020 3216.390 ;
        RECT 2668.020 3216.380 2671.020 3216.390 ;
        RECT 2848.020 3216.380 2851.020 3216.390 ;
        RECT 2959.500 3216.380 2962.500 3216.390 ;
        RECT -42.880 3213.380 2962.500 3216.380 ;
        RECT -42.880 3213.370 -39.880 3213.380 ;
        RECT 148.020 3213.370 151.020 3213.380 ;
        RECT 328.020 3213.370 331.020 3213.380 ;
        RECT 508.020 3213.370 511.020 3213.380 ;
        RECT 688.020 3213.370 691.020 3213.380 ;
        RECT 868.020 3213.370 871.020 3213.380 ;
        RECT 1048.020 3213.370 1051.020 3213.380 ;
        RECT 1228.020 3213.370 1231.020 3213.380 ;
        RECT 1408.020 3213.370 1411.020 3213.380 ;
        RECT 1588.020 3213.370 1591.020 3213.380 ;
        RECT 1768.020 3213.370 1771.020 3213.380 ;
        RECT 1948.020 3213.370 1951.020 3213.380 ;
        RECT 2128.020 3213.370 2131.020 3213.380 ;
        RECT 2308.020 3213.370 2311.020 3213.380 ;
        RECT 2488.020 3213.370 2491.020 3213.380 ;
        RECT 2668.020 3213.370 2671.020 3213.380 ;
        RECT 2848.020 3213.370 2851.020 3213.380 ;
        RECT 2959.500 3213.370 2962.500 3213.380 ;
        RECT -33.480 3198.380 -30.480 3198.390 ;
        RECT 130.020 3198.380 133.020 3198.390 ;
        RECT 310.020 3198.380 313.020 3198.390 ;
        RECT 490.020 3198.380 493.020 3198.390 ;
        RECT 670.020 3198.380 673.020 3198.390 ;
        RECT 850.020 3198.380 853.020 3198.390 ;
        RECT 1030.020 3198.380 1033.020 3198.390 ;
        RECT 1210.020 3198.380 1213.020 3198.390 ;
        RECT 1390.020 3198.380 1393.020 3198.390 ;
        RECT 1570.020 3198.380 1573.020 3198.390 ;
        RECT 1750.020 3198.380 1753.020 3198.390 ;
        RECT 1930.020 3198.380 1933.020 3198.390 ;
        RECT 2110.020 3198.380 2113.020 3198.390 ;
        RECT 2290.020 3198.380 2293.020 3198.390 ;
        RECT 2470.020 3198.380 2473.020 3198.390 ;
        RECT 2650.020 3198.380 2653.020 3198.390 ;
        RECT 2830.020 3198.380 2833.020 3198.390 ;
        RECT 2950.100 3198.380 2953.100 3198.390 ;
        RECT -33.480 3195.380 2953.100 3198.380 ;
        RECT -33.480 3195.370 -30.480 3195.380 ;
        RECT 130.020 3195.370 133.020 3195.380 ;
        RECT 310.020 3195.370 313.020 3195.380 ;
        RECT 490.020 3195.370 493.020 3195.380 ;
        RECT 670.020 3195.370 673.020 3195.380 ;
        RECT 850.020 3195.370 853.020 3195.380 ;
        RECT 1030.020 3195.370 1033.020 3195.380 ;
        RECT 1210.020 3195.370 1213.020 3195.380 ;
        RECT 1390.020 3195.370 1393.020 3195.380 ;
        RECT 1570.020 3195.370 1573.020 3195.380 ;
        RECT 1750.020 3195.370 1753.020 3195.380 ;
        RECT 1930.020 3195.370 1933.020 3195.380 ;
        RECT 2110.020 3195.370 2113.020 3195.380 ;
        RECT 2290.020 3195.370 2293.020 3195.380 ;
        RECT 2470.020 3195.370 2473.020 3195.380 ;
        RECT 2650.020 3195.370 2653.020 3195.380 ;
        RECT 2830.020 3195.370 2833.020 3195.380 ;
        RECT 2950.100 3195.370 2953.100 3195.380 ;
        RECT -24.080 3180.380 -21.080 3180.390 ;
        RECT 112.020 3180.380 115.020 3180.390 ;
        RECT 292.020 3180.380 295.020 3180.390 ;
        RECT 472.020 3180.380 475.020 3180.390 ;
        RECT 652.020 3180.380 655.020 3180.390 ;
        RECT 832.020 3180.380 835.020 3180.390 ;
        RECT 1012.020 3180.380 1015.020 3180.390 ;
        RECT 1192.020 3180.380 1195.020 3180.390 ;
        RECT 1372.020 3180.380 1375.020 3180.390 ;
        RECT 1552.020 3180.380 1555.020 3180.390 ;
        RECT 1732.020 3180.380 1735.020 3180.390 ;
        RECT 1912.020 3180.380 1915.020 3180.390 ;
        RECT 2092.020 3180.380 2095.020 3180.390 ;
        RECT 2272.020 3180.380 2275.020 3180.390 ;
        RECT 2452.020 3180.380 2455.020 3180.390 ;
        RECT 2632.020 3180.380 2635.020 3180.390 ;
        RECT 2812.020 3180.380 2815.020 3180.390 ;
        RECT 2940.700 3180.380 2943.700 3180.390 ;
        RECT -24.080 3177.380 2943.700 3180.380 ;
        RECT -24.080 3177.370 -21.080 3177.380 ;
        RECT 112.020 3177.370 115.020 3177.380 ;
        RECT 292.020 3177.370 295.020 3177.380 ;
        RECT 472.020 3177.370 475.020 3177.380 ;
        RECT 652.020 3177.370 655.020 3177.380 ;
        RECT 832.020 3177.370 835.020 3177.380 ;
        RECT 1012.020 3177.370 1015.020 3177.380 ;
        RECT 1192.020 3177.370 1195.020 3177.380 ;
        RECT 1372.020 3177.370 1375.020 3177.380 ;
        RECT 1552.020 3177.370 1555.020 3177.380 ;
        RECT 1732.020 3177.370 1735.020 3177.380 ;
        RECT 1912.020 3177.370 1915.020 3177.380 ;
        RECT 2092.020 3177.370 2095.020 3177.380 ;
        RECT 2272.020 3177.370 2275.020 3177.380 ;
        RECT 2452.020 3177.370 2455.020 3177.380 ;
        RECT 2632.020 3177.370 2635.020 3177.380 ;
        RECT 2812.020 3177.370 2815.020 3177.380 ;
        RECT 2940.700 3177.370 2943.700 3177.380 ;
        RECT -14.680 3162.380 -11.680 3162.390 ;
        RECT 94.020 3162.380 97.020 3162.390 ;
        RECT 274.020 3162.380 277.020 3162.390 ;
        RECT 454.020 3162.380 457.020 3162.390 ;
        RECT 634.020 3162.380 637.020 3162.390 ;
        RECT 814.020 3162.380 817.020 3162.390 ;
        RECT 994.020 3162.380 997.020 3162.390 ;
        RECT 1174.020 3162.380 1177.020 3162.390 ;
        RECT 1354.020 3162.380 1357.020 3162.390 ;
        RECT 1534.020 3162.380 1537.020 3162.390 ;
        RECT 1714.020 3162.380 1717.020 3162.390 ;
        RECT 1894.020 3162.380 1897.020 3162.390 ;
        RECT 2074.020 3162.380 2077.020 3162.390 ;
        RECT 2254.020 3162.380 2257.020 3162.390 ;
        RECT 2434.020 3162.380 2437.020 3162.390 ;
        RECT 2614.020 3162.380 2617.020 3162.390 ;
        RECT 2794.020 3162.380 2797.020 3162.390 ;
        RECT 2931.300 3162.380 2934.300 3162.390 ;
        RECT -14.680 3159.380 2934.300 3162.380 ;
        RECT -14.680 3159.370 -11.680 3159.380 ;
        RECT 94.020 3159.370 97.020 3159.380 ;
        RECT 274.020 3159.370 277.020 3159.380 ;
        RECT 454.020 3159.370 457.020 3159.380 ;
        RECT 634.020 3159.370 637.020 3159.380 ;
        RECT 814.020 3159.370 817.020 3159.380 ;
        RECT 994.020 3159.370 997.020 3159.380 ;
        RECT 1174.020 3159.370 1177.020 3159.380 ;
        RECT 1354.020 3159.370 1357.020 3159.380 ;
        RECT 1534.020 3159.370 1537.020 3159.380 ;
        RECT 1714.020 3159.370 1717.020 3159.380 ;
        RECT 1894.020 3159.370 1897.020 3159.380 ;
        RECT 2074.020 3159.370 2077.020 3159.380 ;
        RECT 2254.020 3159.370 2257.020 3159.380 ;
        RECT 2434.020 3159.370 2437.020 3159.380 ;
        RECT 2614.020 3159.370 2617.020 3159.380 ;
        RECT 2794.020 3159.370 2797.020 3159.380 ;
        RECT 2931.300 3159.370 2934.300 3159.380 ;
        RECT -42.880 3036.380 -39.880 3036.390 ;
        RECT 148.020 3036.380 151.020 3036.390 ;
        RECT 328.020 3036.380 331.020 3036.390 ;
        RECT 508.020 3036.380 511.020 3036.390 ;
        RECT 688.020 3036.380 691.020 3036.390 ;
        RECT 868.020 3036.380 871.020 3036.390 ;
        RECT 1048.020 3036.380 1051.020 3036.390 ;
        RECT 1228.020 3036.380 1231.020 3036.390 ;
        RECT 1408.020 3036.380 1411.020 3036.390 ;
        RECT 1588.020 3036.380 1591.020 3036.390 ;
        RECT 1768.020 3036.380 1771.020 3036.390 ;
        RECT 1948.020 3036.380 1951.020 3036.390 ;
        RECT 2128.020 3036.380 2131.020 3036.390 ;
        RECT 2308.020 3036.380 2311.020 3036.390 ;
        RECT 2488.020 3036.380 2491.020 3036.390 ;
        RECT 2668.020 3036.380 2671.020 3036.390 ;
        RECT 2848.020 3036.380 2851.020 3036.390 ;
        RECT 2959.500 3036.380 2962.500 3036.390 ;
        RECT -42.880 3033.380 2962.500 3036.380 ;
        RECT -42.880 3033.370 -39.880 3033.380 ;
        RECT 148.020 3033.370 151.020 3033.380 ;
        RECT 328.020 3033.370 331.020 3033.380 ;
        RECT 508.020 3033.370 511.020 3033.380 ;
        RECT 688.020 3033.370 691.020 3033.380 ;
        RECT 868.020 3033.370 871.020 3033.380 ;
        RECT 1048.020 3033.370 1051.020 3033.380 ;
        RECT 1228.020 3033.370 1231.020 3033.380 ;
        RECT 1408.020 3033.370 1411.020 3033.380 ;
        RECT 1588.020 3033.370 1591.020 3033.380 ;
        RECT 1768.020 3033.370 1771.020 3033.380 ;
        RECT 1948.020 3033.370 1951.020 3033.380 ;
        RECT 2128.020 3033.370 2131.020 3033.380 ;
        RECT 2308.020 3033.370 2311.020 3033.380 ;
        RECT 2488.020 3033.370 2491.020 3033.380 ;
        RECT 2668.020 3033.370 2671.020 3033.380 ;
        RECT 2848.020 3033.370 2851.020 3033.380 ;
        RECT 2959.500 3033.370 2962.500 3033.380 ;
        RECT -33.480 3018.380 -30.480 3018.390 ;
        RECT 130.020 3018.380 133.020 3018.390 ;
        RECT 310.020 3018.380 313.020 3018.390 ;
        RECT 490.020 3018.380 493.020 3018.390 ;
        RECT 670.020 3018.380 673.020 3018.390 ;
        RECT 850.020 3018.380 853.020 3018.390 ;
        RECT 1030.020 3018.380 1033.020 3018.390 ;
        RECT 1210.020 3018.380 1213.020 3018.390 ;
        RECT 1390.020 3018.380 1393.020 3018.390 ;
        RECT 1570.020 3018.380 1573.020 3018.390 ;
        RECT 1750.020 3018.380 1753.020 3018.390 ;
        RECT 1930.020 3018.380 1933.020 3018.390 ;
        RECT 2110.020 3018.380 2113.020 3018.390 ;
        RECT 2290.020 3018.380 2293.020 3018.390 ;
        RECT 2470.020 3018.380 2473.020 3018.390 ;
        RECT 2650.020 3018.380 2653.020 3018.390 ;
        RECT 2830.020 3018.380 2833.020 3018.390 ;
        RECT 2950.100 3018.380 2953.100 3018.390 ;
        RECT -33.480 3015.380 2953.100 3018.380 ;
        RECT -33.480 3015.370 -30.480 3015.380 ;
        RECT 130.020 3015.370 133.020 3015.380 ;
        RECT 310.020 3015.370 313.020 3015.380 ;
        RECT 490.020 3015.370 493.020 3015.380 ;
        RECT 670.020 3015.370 673.020 3015.380 ;
        RECT 850.020 3015.370 853.020 3015.380 ;
        RECT 1030.020 3015.370 1033.020 3015.380 ;
        RECT 1210.020 3015.370 1213.020 3015.380 ;
        RECT 1390.020 3015.370 1393.020 3015.380 ;
        RECT 1570.020 3015.370 1573.020 3015.380 ;
        RECT 1750.020 3015.370 1753.020 3015.380 ;
        RECT 1930.020 3015.370 1933.020 3015.380 ;
        RECT 2110.020 3015.370 2113.020 3015.380 ;
        RECT 2290.020 3015.370 2293.020 3015.380 ;
        RECT 2470.020 3015.370 2473.020 3015.380 ;
        RECT 2650.020 3015.370 2653.020 3015.380 ;
        RECT 2830.020 3015.370 2833.020 3015.380 ;
        RECT 2950.100 3015.370 2953.100 3015.380 ;
        RECT -24.080 3000.380 -21.080 3000.390 ;
        RECT 112.020 3000.380 115.020 3000.390 ;
        RECT 292.020 3000.380 295.020 3000.390 ;
        RECT 472.020 3000.380 475.020 3000.390 ;
        RECT 652.020 3000.380 655.020 3000.390 ;
        RECT 832.020 3000.380 835.020 3000.390 ;
        RECT 1012.020 3000.380 1015.020 3000.390 ;
        RECT 1192.020 3000.380 1195.020 3000.390 ;
        RECT 1372.020 3000.380 1375.020 3000.390 ;
        RECT 1552.020 3000.380 1555.020 3000.390 ;
        RECT 1732.020 3000.380 1735.020 3000.390 ;
        RECT 1912.020 3000.380 1915.020 3000.390 ;
        RECT 2092.020 3000.380 2095.020 3000.390 ;
        RECT 2272.020 3000.380 2275.020 3000.390 ;
        RECT 2452.020 3000.380 2455.020 3000.390 ;
        RECT 2632.020 3000.380 2635.020 3000.390 ;
        RECT 2812.020 3000.380 2815.020 3000.390 ;
        RECT 2940.700 3000.380 2943.700 3000.390 ;
        RECT -24.080 2997.380 2943.700 3000.380 ;
        RECT -24.080 2997.370 -21.080 2997.380 ;
        RECT 112.020 2997.370 115.020 2997.380 ;
        RECT 292.020 2997.370 295.020 2997.380 ;
        RECT 472.020 2997.370 475.020 2997.380 ;
        RECT 652.020 2997.370 655.020 2997.380 ;
        RECT 832.020 2997.370 835.020 2997.380 ;
        RECT 1012.020 2997.370 1015.020 2997.380 ;
        RECT 1192.020 2997.370 1195.020 2997.380 ;
        RECT 1372.020 2997.370 1375.020 2997.380 ;
        RECT 1552.020 2997.370 1555.020 2997.380 ;
        RECT 1732.020 2997.370 1735.020 2997.380 ;
        RECT 1912.020 2997.370 1915.020 2997.380 ;
        RECT 2092.020 2997.370 2095.020 2997.380 ;
        RECT 2272.020 2997.370 2275.020 2997.380 ;
        RECT 2452.020 2997.370 2455.020 2997.380 ;
        RECT 2632.020 2997.370 2635.020 2997.380 ;
        RECT 2812.020 2997.370 2815.020 2997.380 ;
        RECT 2940.700 2997.370 2943.700 2997.380 ;
        RECT -14.680 2982.380 -11.680 2982.390 ;
        RECT 94.020 2982.380 97.020 2982.390 ;
        RECT 274.020 2982.380 277.020 2982.390 ;
        RECT 454.020 2982.380 457.020 2982.390 ;
        RECT 634.020 2982.380 637.020 2982.390 ;
        RECT 814.020 2982.380 817.020 2982.390 ;
        RECT 994.020 2982.380 997.020 2982.390 ;
        RECT 1174.020 2982.380 1177.020 2982.390 ;
        RECT 1354.020 2982.380 1357.020 2982.390 ;
        RECT 1534.020 2982.380 1537.020 2982.390 ;
        RECT 1714.020 2982.380 1717.020 2982.390 ;
        RECT 1894.020 2982.380 1897.020 2982.390 ;
        RECT 2074.020 2982.380 2077.020 2982.390 ;
        RECT 2254.020 2982.380 2257.020 2982.390 ;
        RECT 2434.020 2982.380 2437.020 2982.390 ;
        RECT 2614.020 2982.380 2617.020 2982.390 ;
        RECT 2794.020 2982.380 2797.020 2982.390 ;
        RECT 2931.300 2982.380 2934.300 2982.390 ;
        RECT -14.680 2979.380 2934.300 2982.380 ;
        RECT -14.680 2979.370 -11.680 2979.380 ;
        RECT 94.020 2979.370 97.020 2979.380 ;
        RECT 274.020 2979.370 277.020 2979.380 ;
        RECT 454.020 2979.370 457.020 2979.380 ;
        RECT 634.020 2979.370 637.020 2979.380 ;
        RECT 814.020 2979.370 817.020 2979.380 ;
        RECT 994.020 2979.370 997.020 2979.380 ;
        RECT 1174.020 2979.370 1177.020 2979.380 ;
        RECT 1354.020 2979.370 1357.020 2979.380 ;
        RECT 1534.020 2979.370 1537.020 2979.380 ;
        RECT 1714.020 2979.370 1717.020 2979.380 ;
        RECT 1894.020 2979.370 1897.020 2979.380 ;
        RECT 2074.020 2979.370 2077.020 2979.380 ;
        RECT 2254.020 2979.370 2257.020 2979.380 ;
        RECT 2434.020 2979.370 2437.020 2979.380 ;
        RECT 2614.020 2979.370 2617.020 2979.380 ;
        RECT 2794.020 2979.370 2797.020 2979.380 ;
        RECT 2931.300 2979.370 2934.300 2979.380 ;
        RECT -42.880 2856.380 -39.880 2856.390 ;
        RECT 148.020 2856.380 151.020 2856.390 ;
        RECT 328.020 2856.380 331.020 2856.390 ;
        RECT 508.020 2856.380 511.020 2856.390 ;
        RECT 688.020 2856.380 691.020 2856.390 ;
        RECT 868.020 2856.380 871.020 2856.390 ;
        RECT 1048.020 2856.380 1051.020 2856.390 ;
        RECT 1228.020 2856.380 1231.020 2856.390 ;
        RECT 1408.020 2856.380 1411.020 2856.390 ;
        RECT 1588.020 2856.380 1591.020 2856.390 ;
        RECT 1768.020 2856.380 1771.020 2856.390 ;
        RECT 1948.020 2856.380 1951.020 2856.390 ;
        RECT 2128.020 2856.380 2131.020 2856.390 ;
        RECT 2308.020 2856.380 2311.020 2856.390 ;
        RECT 2488.020 2856.380 2491.020 2856.390 ;
        RECT 2668.020 2856.380 2671.020 2856.390 ;
        RECT 2848.020 2856.380 2851.020 2856.390 ;
        RECT 2959.500 2856.380 2962.500 2856.390 ;
        RECT -42.880 2853.380 2962.500 2856.380 ;
        RECT -42.880 2853.370 -39.880 2853.380 ;
        RECT 148.020 2853.370 151.020 2853.380 ;
        RECT 328.020 2853.370 331.020 2853.380 ;
        RECT 508.020 2853.370 511.020 2853.380 ;
        RECT 688.020 2853.370 691.020 2853.380 ;
        RECT 868.020 2853.370 871.020 2853.380 ;
        RECT 1048.020 2853.370 1051.020 2853.380 ;
        RECT 1228.020 2853.370 1231.020 2853.380 ;
        RECT 1408.020 2853.370 1411.020 2853.380 ;
        RECT 1588.020 2853.370 1591.020 2853.380 ;
        RECT 1768.020 2853.370 1771.020 2853.380 ;
        RECT 1948.020 2853.370 1951.020 2853.380 ;
        RECT 2128.020 2853.370 2131.020 2853.380 ;
        RECT 2308.020 2853.370 2311.020 2853.380 ;
        RECT 2488.020 2853.370 2491.020 2853.380 ;
        RECT 2668.020 2853.370 2671.020 2853.380 ;
        RECT 2848.020 2853.370 2851.020 2853.380 ;
        RECT 2959.500 2853.370 2962.500 2853.380 ;
        RECT -33.480 2838.380 -30.480 2838.390 ;
        RECT 130.020 2838.380 133.020 2838.390 ;
        RECT 310.020 2838.380 313.020 2838.390 ;
        RECT 490.020 2838.380 493.020 2838.390 ;
        RECT 670.020 2838.380 673.020 2838.390 ;
        RECT 850.020 2838.380 853.020 2838.390 ;
        RECT 1030.020 2838.380 1033.020 2838.390 ;
        RECT 1210.020 2838.380 1213.020 2838.390 ;
        RECT 1390.020 2838.380 1393.020 2838.390 ;
        RECT 1570.020 2838.380 1573.020 2838.390 ;
        RECT 1750.020 2838.380 1753.020 2838.390 ;
        RECT 1930.020 2838.380 1933.020 2838.390 ;
        RECT 2110.020 2838.380 2113.020 2838.390 ;
        RECT 2290.020 2838.380 2293.020 2838.390 ;
        RECT 2470.020 2838.380 2473.020 2838.390 ;
        RECT 2650.020 2838.380 2653.020 2838.390 ;
        RECT 2830.020 2838.380 2833.020 2838.390 ;
        RECT 2950.100 2838.380 2953.100 2838.390 ;
        RECT -33.480 2835.380 2953.100 2838.380 ;
        RECT -33.480 2835.370 -30.480 2835.380 ;
        RECT 130.020 2835.370 133.020 2835.380 ;
        RECT 310.020 2835.370 313.020 2835.380 ;
        RECT 490.020 2835.370 493.020 2835.380 ;
        RECT 670.020 2835.370 673.020 2835.380 ;
        RECT 850.020 2835.370 853.020 2835.380 ;
        RECT 1030.020 2835.370 1033.020 2835.380 ;
        RECT 1210.020 2835.370 1213.020 2835.380 ;
        RECT 1390.020 2835.370 1393.020 2835.380 ;
        RECT 1570.020 2835.370 1573.020 2835.380 ;
        RECT 1750.020 2835.370 1753.020 2835.380 ;
        RECT 1930.020 2835.370 1933.020 2835.380 ;
        RECT 2110.020 2835.370 2113.020 2835.380 ;
        RECT 2290.020 2835.370 2293.020 2835.380 ;
        RECT 2470.020 2835.370 2473.020 2835.380 ;
        RECT 2650.020 2835.370 2653.020 2835.380 ;
        RECT 2830.020 2835.370 2833.020 2835.380 ;
        RECT 2950.100 2835.370 2953.100 2835.380 ;
        RECT -24.080 2820.380 -21.080 2820.390 ;
        RECT 112.020 2820.380 115.020 2820.390 ;
        RECT 292.020 2820.380 295.020 2820.390 ;
        RECT 472.020 2820.380 475.020 2820.390 ;
        RECT 652.020 2820.380 655.020 2820.390 ;
        RECT 832.020 2820.380 835.020 2820.390 ;
        RECT 1012.020 2820.380 1015.020 2820.390 ;
        RECT 1192.020 2820.380 1195.020 2820.390 ;
        RECT 1372.020 2820.380 1375.020 2820.390 ;
        RECT 1552.020 2820.380 1555.020 2820.390 ;
        RECT 1732.020 2820.380 1735.020 2820.390 ;
        RECT 1912.020 2820.380 1915.020 2820.390 ;
        RECT 2092.020 2820.380 2095.020 2820.390 ;
        RECT 2272.020 2820.380 2275.020 2820.390 ;
        RECT 2452.020 2820.380 2455.020 2820.390 ;
        RECT 2632.020 2820.380 2635.020 2820.390 ;
        RECT 2812.020 2820.380 2815.020 2820.390 ;
        RECT 2940.700 2820.380 2943.700 2820.390 ;
        RECT -24.080 2817.380 2943.700 2820.380 ;
        RECT -24.080 2817.370 -21.080 2817.380 ;
        RECT 112.020 2817.370 115.020 2817.380 ;
        RECT 292.020 2817.370 295.020 2817.380 ;
        RECT 472.020 2817.370 475.020 2817.380 ;
        RECT 652.020 2817.370 655.020 2817.380 ;
        RECT 832.020 2817.370 835.020 2817.380 ;
        RECT 1012.020 2817.370 1015.020 2817.380 ;
        RECT 1192.020 2817.370 1195.020 2817.380 ;
        RECT 1372.020 2817.370 1375.020 2817.380 ;
        RECT 1552.020 2817.370 1555.020 2817.380 ;
        RECT 1732.020 2817.370 1735.020 2817.380 ;
        RECT 1912.020 2817.370 1915.020 2817.380 ;
        RECT 2092.020 2817.370 2095.020 2817.380 ;
        RECT 2272.020 2817.370 2275.020 2817.380 ;
        RECT 2452.020 2817.370 2455.020 2817.380 ;
        RECT 2632.020 2817.370 2635.020 2817.380 ;
        RECT 2812.020 2817.370 2815.020 2817.380 ;
        RECT 2940.700 2817.370 2943.700 2817.380 ;
        RECT -14.680 2802.380 -11.680 2802.390 ;
        RECT 94.020 2802.380 97.020 2802.390 ;
        RECT 274.020 2802.380 277.020 2802.390 ;
        RECT 454.020 2802.380 457.020 2802.390 ;
        RECT 634.020 2802.380 637.020 2802.390 ;
        RECT 814.020 2802.380 817.020 2802.390 ;
        RECT 994.020 2802.380 997.020 2802.390 ;
        RECT 1174.020 2802.380 1177.020 2802.390 ;
        RECT 1354.020 2802.380 1357.020 2802.390 ;
        RECT 1534.020 2802.380 1537.020 2802.390 ;
        RECT 1714.020 2802.380 1717.020 2802.390 ;
        RECT 1894.020 2802.380 1897.020 2802.390 ;
        RECT 2074.020 2802.380 2077.020 2802.390 ;
        RECT 2254.020 2802.380 2257.020 2802.390 ;
        RECT 2434.020 2802.380 2437.020 2802.390 ;
        RECT 2614.020 2802.380 2617.020 2802.390 ;
        RECT 2794.020 2802.380 2797.020 2802.390 ;
        RECT 2931.300 2802.380 2934.300 2802.390 ;
        RECT -14.680 2799.380 2934.300 2802.380 ;
        RECT -14.680 2799.370 -11.680 2799.380 ;
        RECT 94.020 2799.370 97.020 2799.380 ;
        RECT 274.020 2799.370 277.020 2799.380 ;
        RECT 454.020 2799.370 457.020 2799.380 ;
        RECT 634.020 2799.370 637.020 2799.380 ;
        RECT 814.020 2799.370 817.020 2799.380 ;
        RECT 994.020 2799.370 997.020 2799.380 ;
        RECT 1174.020 2799.370 1177.020 2799.380 ;
        RECT 1354.020 2799.370 1357.020 2799.380 ;
        RECT 1534.020 2799.370 1537.020 2799.380 ;
        RECT 1714.020 2799.370 1717.020 2799.380 ;
        RECT 1894.020 2799.370 1897.020 2799.380 ;
        RECT 2074.020 2799.370 2077.020 2799.380 ;
        RECT 2254.020 2799.370 2257.020 2799.380 ;
        RECT 2434.020 2799.370 2437.020 2799.380 ;
        RECT 2614.020 2799.370 2617.020 2799.380 ;
        RECT 2794.020 2799.370 2797.020 2799.380 ;
        RECT 2931.300 2799.370 2934.300 2799.380 ;
        RECT -42.880 2676.380 -39.880 2676.390 ;
        RECT 148.020 2676.380 151.020 2676.390 ;
        RECT 684.690 2676.380 686.310 2676.390 ;
        RECT 868.020 2676.380 871.020 2676.390 ;
        RECT 1334.690 2676.380 1336.310 2676.390 ;
        RECT 1408.020 2676.380 1411.020 2676.390 ;
        RECT 1934.690 2676.380 1936.310 2676.390 ;
        RECT 2128.020 2676.380 2131.020 2676.390 ;
        RECT 2584.690 2676.380 2586.310 2676.390 ;
        RECT 2668.020 2676.380 2671.020 2676.390 ;
        RECT 2848.020 2676.380 2851.020 2676.390 ;
        RECT 2959.500 2676.380 2962.500 2676.390 ;
        RECT -42.880 2673.380 2962.500 2676.380 ;
        RECT -42.880 2673.370 -39.880 2673.380 ;
        RECT 148.020 2673.370 151.020 2673.380 ;
        RECT 684.690 2673.370 686.310 2673.380 ;
        RECT 868.020 2673.370 871.020 2673.380 ;
        RECT 1334.690 2673.370 1336.310 2673.380 ;
        RECT 1408.020 2673.370 1411.020 2673.380 ;
        RECT 1934.690 2673.370 1936.310 2673.380 ;
        RECT 2128.020 2673.370 2131.020 2673.380 ;
        RECT 2584.690 2673.370 2586.310 2673.380 ;
        RECT 2668.020 2673.370 2671.020 2673.380 ;
        RECT 2848.020 2673.370 2851.020 2673.380 ;
        RECT 2959.500 2673.370 2962.500 2673.380 ;
        RECT -33.480 2658.380 -30.480 2658.390 ;
        RECT 130.020 2658.380 133.020 2658.390 ;
        RECT 684.690 2658.380 686.310 2658.390 ;
        RECT 850.020 2658.380 853.020 2658.390 ;
        RECT 1334.690 2658.380 1336.310 2658.390 ;
        RECT 1390.020 2658.380 1393.020 2658.390 ;
        RECT 1934.690 2658.380 1936.310 2658.390 ;
        RECT 2110.020 2658.380 2113.020 2658.390 ;
        RECT 2584.690 2658.380 2586.310 2658.390 ;
        RECT 2650.020 2658.380 2653.020 2658.390 ;
        RECT 2830.020 2658.380 2833.020 2658.390 ;
        RECT 2950.100 2658.380 2953.100 2658.390 ;
        RECT -33.480 2655.380 2953.100 2658.380 ;
        RECT -33.480 2655.370 -30.480 2655.380 ;
        RECT 130.020 2655.370 133.020 2655.380 ;
        RECT 684.690 2655.370 686.310 2655.380 ;
        RECT 850.020 2655.370 853.020 2655.380 ;
        RECT 1334.690 2655.370 1336.310 2655.380 ;
        RECT 1390.020 2655.370 1393.020 2655.380 ;
        RECT 1934.690 2655.370 1936.310 2655.380 ;
        RECT 2110.020 2655.370 2113.020 2655.380 ;
        RECT 2584.690 2655.370 2586.310 2655.380 ;
        RECT 2650.020 2655.370 2653.020 2655.380 ;
        RECT 2830.020 2655.370 2833.020 2655.380 ;
        RECT 2950.100 2655.370 2953.100 2655.380 ;
        RECT -24.080 2640.380 -21.080 2640.390 ;
        RECT 112.020 2640.380 115.020 2640.390 ;
        RECT 684.690 2640.380 686.310 2640.390 ;
        RECT 832.020 2640.380 835.020 2640.390 ;
        RECT 1334.690 2640.380 1336.310 2640.390 ;
        RECT 1372.020 2640.380 1375.020 2640.390 ;
        RECT 1934.690 2640.380 1936.310 2640.390 ;
        RECT 2092.020 2640.380 2095.020 2640.390 ;
        RECT 2584.690 2640.380 2586.310 2640.390 ;
        RECT 2632.020 2640.380 2635.020 2640.390 ;
        RECT 2812.020 2640.380 2815.020 2640.390 ;
        RECT 2940.700 2640.380 2943.700 2640.390 ;
        RECT -24.080 2637.380 2943.700 2640.380 ;
        RECT -24.080 2637.370 -21.080 2637.380 ;
        RECT 112.020 2637.370 115.020 2637.380 ;
        RECT 684.690 2637.370 686.310 2637.380 ;
        RECT 832.020 2637.370 835.020 2637.380 ;
        RECT 1334.690 2637.370 1336.310 2637.380 ;
        RECT 1372.020 2637.370 1375.020 2637.380 ;
        RECT 1934.690 2637.370 1936.310 2637.380 ;
        RECT 2092.020 2637.370 2095.020 2637.380 ;
        RECT 2584.690 2637.370 2586.310 2637.380 ;
        RECT 2632.020 2637.370 2635.020 2637.380 ;
        RECT 2812.020 2637.370 2815.020 2637.380 ;
        RECT 2940.700 2637.370 2943.700 2637.380 ;
        RECT -14.680 2622.380 -11.680 2622.390 ;
        RECT 94.020 2622.380 97.020 2622.390 ;
        RECT 274.020 2622.380 277.020 2622.390 ;
        RECT 684.690 2622.380 686.310 2622.390 ;
        RECT 814.020 2622.380 817.020 2622.390 ;
        RECT 1334.690 2622.380 1336.310 2622.390 ;
        RECT 1354.020 2622.380 1357.020 2622.390 ;
        RECT 1934.690 2622.380 1936.310 2622.390 ;
        RECT 2074.020 2622.380 2077.020 2622.390 ;
        RECT 2584.690 2622.380 2586.310 2622.390 ;
        RECT 2614.020 2622.380 2617.020 2622.390 ;
        RECT 2794.020 2622.380 2797.020 2622.390 ;
        RECT 2931.300 2622.380 2934.300 2622.390 ;
        RECT -14.680 2619.380 2934.300 2622.380 ;
        RECT -14.680 2619.370 -11.680 2619.380 ;
        RECT 94.020 2619.370 97.020 2619.380 ;
        RECT 274.020 2619.370 277.020 2619.380 ;
        RECT 684.690 2619.370 686.310 2619.380 ;
        RECT 814.020 2619.370 817.020 2619.380 ;
        RECT 1334.690 2619.370 1336.310 2619.380 ;
        RECT 1354.020 2619.370 1357.020 2619.380 ;
        RECT 1934.690 2619.370 1936.310 2619.380 ;
        RECT 2074.020 2619.370 2077.020 2619.380 ;
        RECT 2584.690 2619.370 2586.310 2619.380 ;
        RECT 2614.020 2619.370 2617.020 2619.380 ;
        RECT 2794.020 2619.370 2797.020 2619.380 ;
        RECT 2931.300 2619.370 2934.300 2619.380 ;
        RECT -42.880 2496.380 -39.880 2496.390 ;
        RECT 148.020 2496.380 151.020 2496.390 ;
        RECT 684.690 2496.380 686.310 2496.390 ;
        RECT 868.020 2496.380 871.020 2496.390 ;
        RECT 1334.690 2496.380 1336.310 2496.390 ;
        RECT 1408.020 2496.380 1411.020 2496.390 ;
        RECT 1934.690 2496.380 1936.310 2496.390 ;
        RECT 2128.020 2496.380 2131.020 2496.390 ;
        RECT 2584.690 2496.380 2586.310 2496.390 ;
        RECT 2668.020 2496.380 2671.020 2496.390 ;
        RECT 2848.020 2496.380 2851.020 2496.390 ;
        RECT 2959.500 2496.380 2962.500 2496.390 ;
        RECT -42.880 2493.380 2962.500 2496.380 ;
        RECT -42.880 2493.370 -39.880 2493.380 ;
        RECT 148.020 2493.370 151.020 2493.380 ;
        RECT 684.690 2493.370 686.310 2493.380 ;
        RECT 868.020 2493.370 871.020 2493.380 ;
        RECT 1334.690 2493.370 1336.310 2493.380 ;
        RECT 1408.020 2493.370 1411.020 2493.380 ;
        RECT 1934.690 2493.370 1936.310 2493.380 ;
        RECT 2128.020 2493.370 2131.020 2493.380 ;
        RECT 2584.690 2493.370 2586.310 2493.380 ;
        RECT 2668.020 2493.370 2671.020 2493.380 ;
        RECT 2848.020 2493.370 2851.020 2493.380 ;
        RECT 2959.500 2493.370 2962.500 2493.380 ;
        RECT -33.480 2478.380 -30.480 2478.390 ;
        RECT 130.020 2478.380 133.020 2478.390 ;
        RECT 684.690 2478.380 686.310 2478.390 ;
        RECT 850.020 2478.380 853.020 2478.390 ;
        RECT 1334.690 2478.380 1336.310 2478.390 ;
        RECT 1390.020 2478.380 1393.020 2478.390 ;
        RECT 1934.690 2478.380 1936.310 2478.390 ;
        RECT 2110.020 2478.380 2113.020 2478.390 ;
        RECT 2584.690 2478.380 2586.310 2478.390 ;
        RECT 2650.020 2478.380 2653.020 2478.390 ;
        RECT 2830.020 2478.380 2833.020 2478.390 ;
        RECT 2950.100 2478.380 2953.100 2478.390 ;
        RECT -33.480 2475.380 2953.100 2478.380 ;
        RECT -33.480 2475.370 -30.480 2475.380 ;
        RECT 130.020 2475.370 133.020 2475.380 ;
        RECT 684.690 2475.370 686.310 2475.380 ;
        RECT 850.020 2475.370 853.020 2475.380 ;
        RECT 1334.690 2475.370 1336.310 2475.380 ;
        RECT 1390.020 2475.370 1393.020 2475.380 ;
        RECT 1934.690 2475.370 1936.310 2475.380 ;
        RECT 2110.020 2475.370 2113.020 2475.380 ;
        RECT 2584.690 2475.370 2586.310 2475.380 ;
        RECT 2650.020 2475.370 2653.020 2475.380 ;
        RECT 2830.020 2475.370 2833.020 2475.380 ;
        RECT 2950.100 2475.370 2953.100 2475.380 ;
        RECT -24.080 2460.380 -21.080 2460.390 ;
        RECT 112.020 2460.380 115.020 2460.390 ;
        RECT 684.690 2460.380 686.310 2460.390 ;
        RECT 832.020 2460.380 835.020 2460.390 ;
        RECT 1334.690 2460.380 1336.310 2460.390 ;
        RECT 1372.020 2460.380 1375.020 2460.390 ;
        RECT 1934.690 2460.380 1936.310 2460.390 ;
        RECT 2092.020 2460.380 2095.020 2460.390 ;
        RECT 2584.690 2460.380 2586.310 2460.390 ;
        RECT 2632.020 2460.380 2635.020 2460.390 ;
        RECT 2812.020 2460.380 2815.020 2460.390 ;
        RECT 2940.700 2460.380 2943.700 2460.390 ;
        RECT -24.080 2457.380 2943.700 2460.380 ;
        RECT -24.080 2457.370 -21.080 2457.380 ;
        RECT 112.020 2457.370 115.020 2457.380 ;
        RECT 684.690 2457.370 686.310 2457.380 ;
        RECT 832.020 2457.370 835.020 2457.380 ;
        RECT 1334.690 2457.370 1336.310 2457.380 ;
        RECT 1372.020 2457.370 1375.020 2457.380 ;
        RECT 1934.690 2457.370 1936.310 2457.380 ;
        RECT 2092.020 2457.370 2095.020 2457.380 ;
        RECT 2584.690 2457.370 2586.310 2457.380 ;
        RECT 2632.020 2457.370 2635.020 2457.380 ;
        RECT 2812.020 2457.370 2815.020 2457.380 ;
        RECT 2940.700 2457.370 2943.700 2457.380 ;
        RECT -14.680 2442.380 -11.680 2442.390 ;
        RECT 94.020 2442.380 97.020 2442.390 ;
        RECT 274.020 2442.380 277.020 2442.390 ;
        RECT 684.690 2442.380 686.310 2442.390 ;
        RECT 814.020 2442.380 817.020 2442.390 ;
        RECT 1334.690 2442.380 1336.310 2442.390 ;
        RECT 1354.020 2442.380 1357.020 2442.390 ;
        RECT 1934.690 2442.380 1936.310 2442.390 ;
        RECT 2074.020 2442.380 2077.020 2442.390 ;
        RECT 2584.690 2442.380 2586.310 2442.390 ;
        RECT 2614.020 2442.380 2617.020 2442.390 ;
        RECT 2794.020 2442.380 2797.020 2442.390 ;
        RECT 2931.300 2442.380 2934.300 2442.390 ;
        RECT -14.680 2439.380 2934.300 2442.380 ;
        RECT -14.680 2439.370 -11.680 2439.380 ;
        RECT 94.020 2439.370 97.020 2439.380 ;
        RECT 274.020 2439.370 277.020 2439.380 ;
        RECT 684.690 2439.370 686.310 2439.380 ;
        RECT 814.020 2439.370 817.020 2439.380 ;
        RECT 1334.690 2439.370 1336.310 2439.380 ;
        RECT 1354.020 2439.370 1357.020 2439.380 ;
        RECT 1934.690 2439.370 1936.310 2439.380 ;
        RECT 2074.020 2439.370 2077.020 2439.380 ;
        RECT 2584.690 2439.370 2586.310 2439.380 ;
        RECT 2614.020 2439.370 2617.020 2439.380 ;
        RECT 2794.020 2439.370 2797.020 2439.380 ;
        RECT 2931.300 2439.370 2934.300 2439.380 ;
        RECT -42.880 2316.380 -39.880 2316.390 ;
        RECT 148.020 2316.380 151.020 2316.390 ;
        RECT 684.690 2316.380 686.310 2316.390 ;
        RECT 868.020 2316.380 871.020 2316.390 ;
        RECT 1334.690 2316.380 1336.310 2316.390 ;
        RECT 1408.020 2316.380 1411.020 2316.390 ;
        RECT 1934.690 2316.380 1936.310 2316.390 ;
        RECT 2128.020 2316.380 2131.020 2316.390 ;
        RECT 2584.690 2316.380 2586.310 2316.390 ;
        RECT 2668.020 2316.380 2671.020 2316.390 ;
        RECT 2848.020 2316.380 2851.020 2316.390 ;
        RECT 2959.500 2316.380 2962.500 2316.390 ;
        RECT -42.880 2313.380 2962.500 2316.380 ;
        RECT -42.880 2313.370 -39.880 2313.380 ;
        RECT 148.020 2313.370 151.020 2313.380 ;
        RECT 684.690 2313.370 686.310 2313.380 ;
        RECT 868.020 2313.370 871.020 2313.380 ;
        RECT 1334.690 2313.370 1336.310 2313.380 ;
        RECT 1408.020 2313.370 1411.020 2313.380 ;
        RECT 1934.690 2313.370 1936.310 2313.380 ;
        RECT 2128.020 2313.370 2131.020 2313.380 ;
        RECT 2584.690 2313.370 2586.310 2313.380 ;
        RECT 2668.020 2313.370 2671.020 2313.380 ;
        RECT 2848.020 2313.370 2851.020 2313.380 ;
        RECT 2959.500 2313.370 2962.500 2313.380 ;
        RECT -33.480 2298.380 -30.480 2298.390 ;
        RECT 130.020 2298.380 133.020 2298.390 ;
        RECT 850.020 2298.380 853.020 2298.390 ;
        RECT 1390.020 2298.380 1393.020 2298.390 ;
        RECT 2110.020 2298.380 2113.020 2298.390 ;
        RECT 2650.020 2298.380 2653.020 2298.390 ;
        RECT 2830.020 2298.380 2833.020 2298.390 ;
        RECT 2950.100 2298.380 2953.100 2298.390 ;
        RECT -33.480 2295.380 2953.100 2298.380 ;
        RECT -33.480 2295.370 -30.480 2295.380 ;
        RECT 130.020 2295.370 133.020 2295.380 ;
        RECT 850.020 2295.370 853.020 2295.380 ;
        RECT 1390.020 2295.370 1393.020 2295.380 ;
        RECT 2110.020 2295.370 2113.020 2295.380 ;
        RECT 2650.020 2295.370 2653.020 2295.380 ;
        RECT 2830.020 2295.370 2833.020 2295.380 ;
        RECT 2950.100 2295.370 2953.100 2295.380 ;
        RECT -24.080 2280.380 -21.080 2280.390 ;
        RECT 112.020 2280.380 115.020 2280.390 ;
        RECT 292.020 2280.380 295.020 2280.390 ;
        RECT 472.020 2280.380 475.020 2280.390 ;
        RECT 652.020 2280.380 655.020 2280.390 ;
        RECT 832.020 2280.380 835.020 2280.390 ;
        RECT 1012.020 2280.380 1015.020 2280.390 ;
        RECT 1192.020 2280.380 1195.020 2280.390 ;
        RECT 1372.020 2280.380 1375.020 2280.390 ;
        RECT 1552.020 2280.380 1555.020 2280.390 ;
        RECT 1732.020 2280.380 1735.020 2280.390 ;
        RECT 1912.020 2280.380 1915.020 2280.390 ;
        RECT 2092.020 2280.380 2095.020 2280.390 ;
        RECT 2272.020 2280.380 2275.020 2280.390 ;
        RECT 2452.020 2280.380 2455.020 2280.390 ;
        RECT 2632.020 2280.380 2635.020 2280.390 ;
        RECT 2812.020 2280.380 2815.020 2280.390 ;
        RECT 2940.700 2280.380 2943.700 2280.390 ;
        RECT -24.080 2277.380 2943.700 2280.380 ;
        RECT -24.080 2277.370 -21.080 2277.380 ;
        RECT 112.020 2277.370 115.020 2277.380 ;
        RECT 292.020 2277.370 295.020 2277.380 ;
        RECT 472.020 2277.370 475.020 2277.380 ;
        RECT 652.020 2277.370 655.020 2277.380 ;
        RECT 832.020 2277.370 835.020 2277.380 ;
        RECT 1012.020 2277.370 1015.020 2277.380 ;
        RECT 1192.020 2277.370 1195.020 2277.380 ;
        RECT 1372.020 2277.370 1375.020 2277.380 ;
        RECT 1552.020 2277.370 1555.020 2277.380 ;
        RECT 1732.020 2277.370 1735.020 2277.380 ;
        RECT 1912.020 2277.370 1915.020 2277.380 ;
        RECT 2092.020 2277.370 2095.020 2277.380 ;
        RECT 2272.020 2277.370 2275.020 2277.380 ;
        RECT 2452.020 2277.370 2455.020 2277.380 ;
        RECT 2632.020 2277.370 2635.020 2277.380 ;
        RECT 2812.020 2277.370 2815.020 2277.380 ;
        RECT 2940.700 2277.370 2943.700 2277.380 ;
        RECT -14.680 2262.380 -11.680 2262.390 ;
        RECT 94.020 2262.380 97.020 2262.390 ;
        RECT 274.020 2262.380 277.020 2262.390 ;
        RECT 454.020 2262.380 457.020 2262.390 ;
        RECT 634.020 2262.380 637.020 2262.390 ;
        RECT 814.020 2262.380 817.020 2262.390 ;
        RECT 994.020 2262.380 997.020 2262.390 ;
        RECT 1174.020 2262.380 1177.020 2262.390 ;
        RECT 1354.020 2262.380 1357.020 2262.390 ;
        RECT 1534.020 2262.380 1537.020 2262.390 ;
        RECT 1714.020 2262.380 1717.020 2262.390 ;
        RECT 1894.020 2262.380 1897.020 2262.390 ;
        RECT 2074.020 2262.380 2077.020 2262.390 ;
        RECT 2254.020 2262.380 2257.020 2262.390 ;
        RECT 2434.020 2262.380 2437.020 2262.390 ;
        RECT 2614.020 2262.380 2617.020 2262.390 ;
        RECT 2794.020 2262.380 2797.020 2262.390 ;
        RECT 2931.300 2262.380 2934.300 2262.390 ;
        RECT -14.680 2259.380 2934.300 2262.380 ;
        RECT -14.680 2259.370 -11.680 2259.380 ;
        RECT 94.020 2259.370 97.020 2259.380 ;
        RECT 274.020 2259.370 277.020 2259.380 ;
        RECT 454.020 2259.370 457.020 2259.380 ;
        RECT 634.020 2259.370 637.020 2259.380 ;
        RECT 814.020 2259.370 817.020 2259.380 ;
        RECT 994.020 2259.370 997.020 2259.380 ;
        RECT 1174.020 2259.370 1177.020 2259.380 ;
        RECT 1354.020 2259.370 1357.020 2259.380 ;
        RECT 1534.020 2259.370 1537.020 2259.380 ;
        RECT 1714.020 2259.370 1717.020 2259.380 ;
        RECT 1894.020 2259.370 1897.020 2259.380 ;
        RECT 2074.020 2259.370 2077.020 2259.380 ;
        RECT 2254.020 2259.370 2257.020 2259.380 ;
        RECT 2434.020 2259.370 2437.020 2259.380 ;
        RECT 2614.020 2259.370 2617.020 2259.380 ;
        RECT 2794.020 2259.370 2797.020 2259.380 ;
        RECT 2931.300 2259.370 2934.300 2259.380 ;
        RECT -42.880 2136.380 -39.880 2136.390 ;
        RECT 148.020 2136.380 151.020 2136.390 ;
        RECT 397.840 2136.380 399.440 2136.390 ;
        RECT 1588.020 2136.380 1591.020 2136.390 ;
        RECT 1768.020 2136.380 1771.020 2136.390 ;
        RECT 1948.020 2136.380 1951.020 2136.390 ;
        RECT 2128.020 2136.380 2131.020 2136.390 ;
        RECT 2308.020 2136.380 2311.020 2136.390 ;
        RECT 2488.020 2136.380 2491.020 2136.390 ;
        RECT 2668.020 2136.380 2671.020 2136.390 ;
        RECT 2848.020 2136.380 2851.020 2136.390 ;
        RECT 2959.500 2136.380 2962.500 2136.390 ;
        RECT -42.880 2133.380 2962.500 2136.380 ;
        RECT -42.880 2133.370 -39.880 2133.380 ;
        RECT 148.020 2133.370 151.020 2133.380 ;
        RECT 397.840 2133.370 399.440 2133.380 ;
        RECT 1588.020 2133.370 1591.020 2133.380 ;
        RECT 1768.020 2133.370 1771.020 2133.380 ;
        RECT 1948.020 2133.370 1951.020 2133.380 ;
        RECT 2128.020 2133.370 2131.020 2133.380 ;
        RECT 2308.020 2133.370 2311.020 2133.380 ;
        RECT 2488.020 2133.370 2491.020 2133.380 ;
        RECT 2668.020 2133.370 2671.020 2133.380 ;
        RECT 2848.020 2133.370 2851.020 2133.380 ;
        RECT 2959.500 2133.370 2962.500 2133.380 ;
        RECT -33.480 2118.380 -30.480 2118.390 ;
        RECT 130.020 2118.380 133.020 2118.390 ;
        RECT 397.840 2118.380 399.440 2118.390 ;
        RECT 1570.020 2118.380 1573.020 2118.390 ;
        RECT 1750.020 2118.380 1753.020 2118.390 ;
        RECT 1930.020 2118.380 1933.020 2118.390 ;
        RECT 2110.020 2118.380 2113.020 2118.390 ;
        RECT 2290.020 2118.380 2293.020 2118.390 ;
        RECT 2470.020 2118.380 2473.020 2118.390 ;
        RECT 2650.020 2118.380 2653.020 2118.390 ;
        RECT 2830.020 2118.380 2833.020 2118.390 ;
        RECT 2950.100 2118.380 2953.100 2118.390 ;
        RECT -33.480 2115.380 2953.100 2118.380 ;
        RECT -33.480 2115.370 -30.480 2115.380 ;
        RECT 130.020 2115.370 133.020 2115.380 ;
        RECT 397.840 2115.370 399.440 2115.380 ;
        RECT 1570.020 2115.370 1573.020 2115.380 ;
        RECT 1750.020 2115.370 1753.020 2115.380 ;
        RECT 1930.020 2115.370 1933.020 2115.380 ;
        RECT 2110.020 2115.370 2113.020 2115.380 ;
        RECT 2290.020 2115.370 2293.020 2115.380 ;
        RECT 2470.020 2115.370 2473.020 2115.380 ;
        RECT 2650.020 2115.370 2653.020 2115.380 ;
        RECT 2830.020 2115.370 2833.020 2115.380 ;
        RECT 2950.100 2115.370 2953.100 2115.380 ;
        RECT -24.080 2100.380 -21.080 2100.390 ;
        RECT 112.020 2100.380 115.020 2100.390 ;
        RECT 397.840 2100.380 399.440 2100.390 ;
        RECT 1552.020 2100.380 1555.020 2100.390 ;
        RECT 1732.020 2100.380 1735.020 2100.390 ;
        RECT 1912.020 2100.380 1915.020 2100.390 ;
        RECT 2092.020 2100.380 2095.020 2100.390 ;
        RECT 2272.020 2100.380 2275.020 2100.390 ;
        RECT 2452.020 2100.380 2455.020 2100.390 ;
        RECT 2632.020 2100.380 2635.020 2100.390 ;
        RECT 2812.020 2100.380 2815.020 2100.390 ;
        RECT 2940.700 2100.380 2943.700 2100.390 ;
        RECT -24.080 2097.380 2943.700 2100.380 ;
        RECT -24.080 2097.370 -21.080 2097.380 ;
        RECT 112.020 2097.370 115.020 2097.380 ;
        RECT 397.840 2097.370 399.440 2097.380 ;
        RECT 1552.020 2097.370 1555.020 2097.380 ;
        RECT 1732.020 2097.370 1735.020 2097.380 ;
        RECT 1912.020 2097.370 1915.020 2097.380 ;
        RECT 2092.020 2097.370 2095.020 2097.380 ;
        RECT 2272.020 2097.370 2275.020 2097.380 ;
        RECT 2452.020 2097.370 2455.020 2097.380 ;
        RECT 2632.020 2097.370 2635.020 2097.380 ;
        RECT 2812.020 2097.370 2815.020 2097.380 ;
        RECT 2940.700 2097.370 2943.700 2097.380 ;
        RECT -14.680 2082.380 -11.680 2082.390 ;
        RECT 94.020 2082.380 97.020 2082.390 ;
        RECT 274.020 2082.380 277.020 2082.390 ;
        RECT 397.840 2082.380 399.440 2082.390 ;
        RECT 1534.020 2082.380 1537.020 2082.390 ;
        RECT 1714.020 2082.380 1717.020 2082.390 ;
        RECT 1894.020 2082.380 1897.020 2082.390 ;
        RECT 2074.020 2082.380 2077.020 2082.390 ;
        RECT 2254.020 2082.380 2257.020 2082.390 ;
        RECT 2434.020 2082.380 2437.020 2082.390 ;
        RECT 2614.020 2082.380 2617.020 2082.390 ;
        RECT 2794.020 2082.380 2797.020 2082.390 ;
        RECT 2931.300 2082.380 2934.300 2082.390 ;
        RECT -14.680 2079.380 2934.300 2082.380 ;
        RECT -14.680 2079.370 -11.680 2079.380 ;
        RECT 94.020 2079.370 97.020 2079.380 ;
        RECT 274.020 2079.370 277.020 2079.380 ;
        RECT 397.840 2079.370 399.440 2079.380 ;
        RECT 1534.020 2079.370 1537.020 2079.380 ;
        RECT 1714.020 2079.370 1717.020 2079.380 ;
        RECT 1894.020 2079.370 1897.020 2079.380 ;
        RECT 2074.020 2079.370 2077.020 2079.380 ;
        RECT 2254.020 2079.370 2257.020 2079.380 ;
        RECT 2434.020 2079.370 2437.020 2079.380 ;
        RECT 2614.020 2079.370 2617.020 2079.380 ;
        RECT 2794.020 2079.370 2797.020 2079.380 ;
        RECT 2931.300 2079.370 2934.300 2079.380 ;
        RECT -42.880 1956.380 -39.880 1956.390 ;
        RECT 148.020 1956.380 151.020 1956.390 ;
        RECT 397.840 1956.380 399.440 1956.390 ;
        RECT 1588.020 1956.380 1591.020 1956.390 ;
        RECT 1768.020 1956.380 1771.020 1956.390 ;
        RECT 1948.020 1956.380 1951.020 1956.390 ;
        RECT 2128.020 1956.380 2131.020 1956.390 ;
        RECT 2308.020 1956.380 2311.020 1956.390 ;
        RECT 2488.020 1956.380 2491.020 1956.390 ;
        RECT 2668.020 1956.380 2671.020 1956.390 ;
        RECT 2848.020 1956.380 2851.020 1956.390 ;
        RECT 2959.500 1956.380 2962.500 1956.390 ;
        RECT -42.880 1953.380 2962.500 1956.380 ;
        RECT -42.880 1953.370 -39.880 1953.380 ;
        RECT 148.020 1953.370 151.020 1953.380 ;
        RECT 397.840 1953.370 399.440 1953.380 ;
        RECT 1588.020 1953.370 1591.020 1953.380 ;
        RECT 1768.020 1953.370 1771.020 1953.380 ;
        RECT 1948.020 1953.370 1951.020 1953.380 ;
        RECT 2128.020 1953.370 2131.020 1953.380 ;
        RECT 2308.020 1953.370 2311.020 1953.380 ;
        RECT 2488.020 1953.370 2491.020 1953.380 ;
        RECT 2668.020 1953.370 2671.020 1953.380 ;
        RECT 2848.020 1953.370 2851.020 1953.380 ;
        RECT 2959.500 1953.370 2962.500 1953.380 ;
        RECT -33.480 1938.380 -30.480 1938.390 ;
        RECT 130.020 1938.380 133.020 1938.390 ;
        RECT 397.840 1938.380 399.440 1938.390 ;
        RECT 1570.020 1938.380 1573.020 1938.390 ;
        RECT 1750.020 1938.380 1753.020 1938.390 ;
        RECT 1930.020 1938.380 1933.020 1938.390 ;
        RECT 2110.020 1938.380 2113.020 1938.390 ;
        RECT 2290.020 1938.380 2293.020 1938.390 ;
        RECT 2470.020 1938.380 2473.020 1938.390 ;
        RECT 2650.020 1938.380 2653.020 1938.390 ;
        RECT 2830.020 1938.380 2833.020 1938.390 ;
        RECT 2950.100 1938.380 2953.100 1938.390 ;
        RECT -33.480 1935.380 2953.100 1938.380 ;
        RECT -33.480 1935.370 -30.480 1935.380 ;
        RECT 130.020 1935.370 133.020 1935.380 ;
        RECT 397.840 1935.370 399.440 1935.380 ;
        RECT 1570.020 1935.370 1573.020 1935.380 ;
        RECT 1750.020 1935.370 1753.020 1935.380 ;
        RECT 1930.020 1935.370 1933.020 1935.380 ;
        RECT 2110.020 1935.370 2113.020 1935.380 ;
        RECT 2290.020 1935.370 2293.020 1935.380 ;
        RECT 2470.020 1935.370 2473.020 1935.380 ;
        RECT 2650.020 1935.370 2653.020 1935.380 ;
        RECT 2830.020 1935.370 2833.020 1935.380 ;
        RECT 2950.100 1935.370 2953.100 1935.380 ;
        RECT -24.080 1920.380 -21.080 1920.390 ;
        RECT 112.020 1920.380 115.020 1920.390 ;
        RECT 397.840 1920.380 399.440 1920.390 ;
        RECT 1552.020 1920.380 1555.020 1920.390 ;
        RECT 1732.020 1920.380 1735.020 1920.390 ;
        RECT 1912.020 1920.380 1915.020 1920.390 ;
        RECT 2092.020 1920.380 2095.020 1920.390 ;
        RECT 2272.020 1920.380 2275.020 1920.390 ;
        RECT 2452.020 1920.380 2455.020 1920.390 ;
        RECT 2632.020 1920.380 2635.020 1920.390 ;
        RECT 2812.020 1920.380 2815.020 1920.390 ;
        RECT 2940.700 1920.380 2943.700 1920.390 ;
        RECT -24.080 1917.380 2943.700 1920.380 ;
        RECT -24.080 1917.370 -21.080 1917.380 ;
        RECT 112.020 1917.370 115.020 1917.380 ;
        RECT 397.840 1917.370 399.440 1917.380 ;
        RECT 1552.020 1917.370 1555.020 1917.380 ;
        RECT 1732.020 1917.370 1735.020 1917.380 ;
        RECT 1912.020 1917.370 1915.020 1917.380 ;
        RECT 2092.020 1917.370 2095.020 1917.380 ;
        RECT 2272.020 1917.370 2275.020 1917.380 ;
        RECT 2452.020 1917.370 2455.020 1917.380 ;
        RECT 2632.020 1917.370 2635.020 1917.380 ;
        RECT 2812.020 1917.370 2815.020 1917.380 ;
        RECT 2940.700 1917.370 2943.700 1917.380 ;
        RECT -14.680 1902.380 -11.680 1902.390 ;
        RECT 94.020 1902.380 97.020 1902.390 ;
        RECT 274.020 1902.380 277.020 1902.390 ;
        RECT 397.840 1902.380 399.440 1902.390 ;
        RECT 1534.020 1902.380 1537.020 1902.390 ;
        RECT 1714.020 1902.380 1717.020 1902.390 ;
        RECT 1894.020 1902.380 1897.020 1902.390 ;
        RECT 2074.020 1902.380 2077.020 1902.390 ;
        RECT 2254.020 1902.380 2257.020 1902.390 ;
        RECT 2434.020 1902.380 2437.020 1902.390 ;
        RECT 2614.020 1902.380 2617.020 1902.390 ;
        RECT 2794.020 1902.380 2797.020 1902.390 ;
        RECT 2931.300 1902.380 2934.300 1902.390 ;
        RECT -14.680 1899.380 2934.300 1902.380 ;
        RECT -14.680 1899.370 -11.680 1899.380 ;
        RECT 94.020 1899.370 97.020 1899.380 ;
        RECT 274.020 1899.370 277.020 1899.380 ;
        RECT 397.840 1899.370 399.440 1899.380 ;
        RECT 1534.020 1899.370 1537.020 1899.380 ;
        RECT 1714.020 1899.370 1717.020 1899.380 ;
        RECT 1894.020 1899.370 1897.020 1899.380 ;
        RECT 2074.020 1899.370 2077.020 1899.380 ;
        RECT 2254.020 1899.370 2257.020 1899.380 ;
        RECT 2434.020 1899.370 2437.020 1899.380 ;
        RECT 2614.020 1899.370 2617.020 1899.380 ;
        RECT 2794.020 1899.370 2797.020 1899.380 ;
        RECT 2931.300 1899.370 2934.300 1899.380 ;
        RECT -42.880 1776.380 -39.880 1776.390 ;
        RECT 148.020 1776.380 151.020 1776.390 ;
        RECT 397.840 1776.380 399.440 1776.390 ;
        RECT 1588.020 1776.380 1591.020 1776.390 ;
        RECT 1768.020 1776.380 1771.020 1776.390 ;
        RECT 1948.020 1776.380 1951.020 1776.390 ;
        RECT 2128.020 1776.380 2131.020 1776.390 ;
        RECT 2308.020 1776.380 2311.020 1776.390 ;
        RECT 2488.020 1776.380 2491.020 1776.390 ;
        RECT 2668.020 1776.380 2671.020 1776.390 ;
        RECT 2848.020 1776.380 2851.020 1776.390 ;
        RECT 2959.500 1776.380 2962.500 1776.390 ;
        RECT -42.880 1773.380 2962.500 1776.380 ;
        RECT -42.880 1773.370 -39.880 1773.380 ;
        RECT 148.020 1773.370 151.020 1773.380 ;
        RECT 397.840 1773.370 399.440 1773.380 ;
        RECT 1588.020 1773.370 1591.020 1773.380 ;
        RECT 1768.020 1773.370 1771.020 1773.380 ;
        RECT 1948.020 1773.370 1951.020 1773.380 ;
        RECT 2128.020 1773.370 2131.020 1773.380 ;
        RECT 2308.020 1773.370 2311.020 1773.380 ;
        RECT 2488.020 1773.370 2491.020 1773.380 ;
        RECT 2668.020 1773.370 2671.020 1773.380 ;
        RECT 2848.020 1773.370 2851.020 1773.380 ;
        RECT 2959.500 1773.370 2962.500 1773.380 ;
        RECT -33.480 1758.380 -30.480 1758.390 ;
        RECT 130.020 1758.380 133.020 1758.390 ;
        RECT 397.840 1758.380 399.440 1758.390 ;
        RECT 1570.020 1758.380 1573.020 1758.390 ;
        RECT 1750.020 1758.380 1753.020 1758.390 ;
        RECT 1930.020 1758.380 1933.020 1758.390 ;
        RECT 2110.020 1758.380 2113.020 1758.390 ;
        RECT 2290.020 1758.380 2293.020 1758.390 ;
        RECT 2470.020 1758.380 2473.020 1758.390 ;
        RECT 2650.020 1758.380 2653.020 1758.390 ;
        RECT 2830.020 1758.380 2833.020 1758.390 ;
        RECT 2950.100 1758.380 2953.100 1758.390 ;
        RECT -33.480 1755.380 2953.100 1758.380 ;
        RECT -33.480 1755.370 -30.480 1755.380 ;
        RECT 130.020 1755.370 133.020 1755.380 ;
        RECT 397.840 1755.370 399.440 1755.380 ;
        RECT 1570.020 1755.370 1573.020 1755.380 ;
        RECT 1750.020 1755.370 1753.020 1755.380 ;
        RECT 1930.020 1755.370 1933.020 1755.380 ;
        RECT 2110.020 1755.370 2113.020 1755.380 ;
        RECT 2290.020 1755.370 2293.020 1755.380 ;
        RECT 2470.020 1755.370 2473.020 1755.380 ;
        RECT 2650.020 1755.370 2653.020 1755.380 ;
        RECT 2830.020 1755.370 2833.020 1755.380 ;
        RECT 2950.100 1755.370 2953.100 1755.380 ;
        RECT -24.080 1740.380 -21.080 1740.390 ;
        RECT 112.020 1740.380 115.020 1740.390 ;
        RECT 397.840 1740.380 399.440 1740.390 ;
        RECT 1552.020 1740.380 1555.020 1740.390 ;
        RECT 1732.020 1740.380 1735.020 1740.390 ;
        RECT 1912.020 1740.380 1915.020 1740.390 ;
        RECT 2092.020 1740.380 2095.020 1740.390 ;
        RECT 2272.020 1740.380 2275.020 1740.390 ;
        RECT 2452.020 1740.380 2455.020 1740.390 ;
        RECT 2632.020 1740.380 2635.020 1740.390 ;
        RECT 2812.020 1740.380 2815.020 1740.390 ;
        RECT 2940.700 1740.380 2943.700 1740.390 ;
        RECT -24.080 1737.380 2943.700 1740.380 ;
        RECT -24.080 1737.370 -21.080 1737.380 ;
        RECT 112.020 1737.370 115.020 1737.380 ;
        RECT 397.840 1737.370 399.440 1737.380 ;
        RECT 1552.020 1737.370 1555.020 1737.380 ;
        RECT 1732.020 1737.370 1735.020 1737.380 ;
        RECT 1912.020 1737.370 1915.020 1737.380 ;
        RECT 2092.020 1737.370 2095.020 1737.380 ;
        RECT 2272.020 1737.370 2275.020 1737.380 ;
        RECT 2452.020 1737.370 2455.020 1737.380 ;
        RECT 2632.020 1737.370 2635.020 1737.380 ;
        RECT 2812.020 1737.370 2815.020 1737.380 ;
        RECT 2940.700 1737.370 2943.700 1737.380 ;
        RECT -14.680 1722.380 -11.680 1722.390 ;
        RECT 94.020 1722.380 97.020 1722.390 ;
        RECT 274.020 1722.380 277.020 1722.390 ;
        RECT 397.840 1722.380 399.440 1722.390 ;
        RECT 1534.020 1722.380 1537.020 1722.390 ;
        RECT 1714.020 1722.380 1717.020 1722.390 ;
        RECT 1894.020 1722.380 1897.020 1722.390 ;
        RECT 2074.020 1722.380 2077.020 1722.390 ;
        RECT 2254.020 1722.380 2257.020 1722.390 ;
        RECT 2434.020 1722.380 2437.020 1722.390 ;
        RECT 2614.020 1722.380 2617.020 1722.390 ;
        RECT 2794.020 1722.380 2797.020 1722.390 ;
        RECT 2931.300 1722.380 2934.300 1722.390 ;
        RECT -14.680 1719.380 2934.300 1722.380 ;
        RECT -14.680 1719.370 -11.680 1719.380 ;
        RECT 94.020 1719.370 97.020 1719.380 ;
        RECT 274.020 1719.370 277.020 1719.380 ;
        RECT 397.840 1719.370 399.440 1719.380 ;
        RECT 1534.020 1719.370 1537.020 1719.380 ;
        RECT 1714.020 1719.370 1717.020 1719.380 ;
        RECT 1894.020 1719.370 1897.020 1719.380 ;
        RECT 2074.020 1719.370 2077.020 1719.380 ;
        RECT 2254.020 1719.370 2257.020 1719.380 ;
        RECT 2434.020 1719.370 2437.020 1719.380 ;
        RECT 2614.020 1719.370 2617.020 1719.380 ;
        RECT 2794.020 1719.370 2797.020 1719.380 ;
        RECT 2931.300 1719.370 2934.300 1719.380 ;
        RECT -42.880 1596.380 -39.880 1596.390 ;
        RECT 148.020 1596.380 151.020 1596.390 ;
        RECT 397.840 1596.380 399.440 1596.390 ;
        RECT 1588.020 1596.380 1591.020 1596.390 ;
        RECT 1768.020 1596.380 1771.020 1596.390 ;
        RECT 1948.020 1596.380 1951.020 1596.390 ;
        RECT 2128.020 1596.380 2131.020 1596.390 ;
        RECT 2308.020 1596.380 2311.020 1596.390 ;
        RECT 2488.020 1596.380 2491.020 1596.390 ;
        RECT 2668.020 1596.380 2671.020 1596.390 ;
        RECT 2848.020 1596.380 2851.020 1596.390 ;
        RECT 2959.500 1596.380 2962.500 1596.390 ;
        RECT -42.880 1593.380 2962.500 1596.380 ;
        RECT -42.880 1593.370 -39.880 1593.380 ;
        RECT 148.020 1593.370 151.020 1593.380 ;
        RECT 397.840 1593.370 399.440 1593.380 ;
        RECT 1588.020 1593.370 1591.020 1593.380 ;
        RECT 1768.020 1593.370 1771.020 1593.380 ;
        RECT 1948.020 1593.370 1951.020 1593.380 ;
        RECT 2128.020 1593.370 2131.020 1593.380 ;
        RECT 2308.020 1593.370 2311.020 1593.380 ;
        RECT 2488.020 1593.370 2491.020 1593.380 ;
        RECT 2668.020 1593.370 2671.020 1593.380 ;
        RECT 2848.020 1593.370 2851.020 1593.380 ;
        RECT 2959.500 1593.370 2962.500 1593.380 ;
        RECT -33.480 1578.380 -30.480 1578.390 ;
        RECT 130.020 1578.380 133.020 1578.390 ;
        RECT 397.840 1578.380 399.440 1578.390 ;
        RECT 1570.020 1578.380 1573.020 1578.390 ;
        RECT 1750.020 1578.380 1753.020 1578.390 ;
        RECT 1930.020 1578.380 1933.020 1578.390 ;
        RECT 2110.020 1578.380 2113.020 1578.390 ;
        RECT 2290.020 1578.380 2293.020 1578.390 ;
        RECT 2470.020 1578.380 2473.020 1578.390 ;
        RECT 2650.020 1578.380 2653.020 1578.390 ;
        RECT 2830.020 1578.380 2833.020 1578.390 ;
        RECT 2950.100 1578.380 2953.100 1578.390 ;
        RECT -33.480 1575.380 2953.100 1578.380 ;
        RECT -33.480 1575.370 -30.480 1575.380 ;
        RECT 130.020 1575.370 133.020 1575.380 ;
        RECT 397.840 1575.370 399.440 1575.380 ;
        RECT 1570.020 1575.370 1573.020 1575.380 ;
        RECT 1750.020 1575.370 1753.020 1575.380 ;
        RECT 1930.020 1575.370 1933.020 1575.380 ;
        RECT 2110.020 1575.370 2113.020 1575.380 ;
        RECT 2290.020 1575.370 2293.020 1575.380 ;
        RECT 2470.020 1575.370 2473.020 1575.380 ;
        RECT 2650.020 1575.370 2653.020 1575.380 ;
        RECT 2830.020 1575.370 2833.020 1575.380 ;
        RECT 2950.100 1575.370 2953.100 1575.380 ;
        RECT -24.080 1560.380 -21.080 1560.390 ;
        RECT 112.020 1560.380 115.020 1560.390 ;
        RECT 397.840 1560.380 399.440 1560.390 ;
        RECT 1552.020 1560.380 1555.020 1560.390 ;
        RECT 1732.020 1560.380 1735.020 1560.390 ;
        RECT 1912.020 1560.380 1915.020 1560.390 ;
        RECT 2092.020 1560.380 2095.020 1560.390 ;
        RECT 2272.020 1560.380 2275.020 1560.390 ;
        RECT 2452.020 1560.380 2455.020 1560.390 ;
        RECT 2632.020 1560.380 2635.020 1560.390 ;
        RECT 2812.020 1560.380 2815.020 1560.390 ;
        RECT 2940.700 1560.380 2943.700 1560.390 ;
        RECT -24.080 1557.380 2943.700 1560.380 ;
        RECT -24.080 1557.370 -21.080 1557.380 ;
        RECT 112.020 1557.370 115.020 1557.380 ;
        RECT 397.840 1557.370 399.440 1557.380 ;
        RECT 1552.020 1557.370 1555.020 1557.380 ;
        RECT 1732.020 1557.370 1735.020 1557.380 ;
        RECT 1912.020 1557.370 1915.020 1557.380 ;
        RECT 2092.020 1557.370 2095.020 1557.380 ;
        RECT 2272.020 1557.370 2275.020 1557.380 ;
        RECT 2452.020 1557.370 2455.020 1557.380 ;
        RECT 2632.020 1557.370 2635.020 1557.380 ;
        RECT 2812.020 1557.370 2815.020 1557.380 ;
        RECT 2940.700 1557.370 2943.700 1557.380 ;
        RECT -14.680 1542.380 -11.680 1542.390 ;
        RECT 94.020 1542.380 97.020 1542.390 ;
        RECT 274.020 1542.380 277.020 1542.390 ;
        RECT 397.840 1542.380 399.440 1542.390 ;
        RECT 1534.020 1542.380 1537.020 1542.390 ;
        RECT 1714.020 1542.380 1717.020 1542.390 ;
        RECT 1894.020 1542.380 1897.020 1542.390 ;
        RECT 2074.020 1542.380 2077.020 1542.390 ;
        RECT 2254.020 1542.380 2257.020 1542.390 ;
        RECT 2434.020 1542.380 2437.020 1542.390 ;
        RECT 2614.020 1542.380 2617.020 1542.390 ;
        RECT 2794.020 1542.380 2797.020 1542.390 ;
        RECT 2931.300 1542.380 2934.300 1542.390 ;
        RECT -14.680 1539.380 2934.300 1542.380 ;
        RECT -14.680 1539.370 -11.680 1539.380 ;
        RECT 94.020 1539.370 97.020 1539.380 ;
        RECT 274.020 1539.370 277.020 1539.380 ;
        RECT 397.840 1539.370 399.440 1539.380 ;
        RECT 1534.020 1539.370 1537.020 1539.380 ;
        RECT 1714.020 1539.370 1717.020 1539.380 ;
        RECT 1894.020 1539.370 1897.020 1539.380 ;
        RECT 2074.020 1539.370 2077.020 1539.380 ;
        RECT 2254.020 1539.370 2257.020 1539.380 ;
        RECT 2434.020 1539.370 2437.020 1539.380 ;
        RECT 2614.020 1539.370 2617.020 1539.380 ;
        RECT 2794.020 1539.370 2797.020 1539.380 ;
        RECT 2931.300 1539.370 2934.300 1539.380 ;
        RECT -42.880 1416.380 -39.880 1416.390 ;
        RECT 148.020 1416.380 151.020 1416.390 ;
        RECT 397.840 1416.380 399.440 1416.390 ;
        RECT 1588.020 1416.380 1591.020 1416.390 ;
        RECT 1768.020 1416.380 1771.020 1416.390 ;
        RECT 1948.020 1416.380 1951.020 1416.390 ;
        RECT 2128.020 1416.380 2131.020 1416.390 ;
        RECT 2308.020 1416.380 2311.020 1416.390 ;
        RECT 2488.020 1416.380 2491.020 1416.390 ;
        RECT 2668.020 1416.380 2671.020 1416.390 ;
        RECT 2848.020 1416.380 2851.020 1416.390 ;
        RECT 2959.500 1416.380 2962.500 1416.390 ;
        RECT -42.880 1413.380 2962.500 1416.380 ;
        RECT -42.880 1413.370 -39.880 1413.380 ;
        RECT 148.020 1413.370 151.020 1413.380 ;
        RECT 397.840 1413.370 399.440 1413.380 ;
        RECT 1588.020 1413.370 1591.020 1413.380 ;
        RECT 1768.020 1413.370 1771.020 1413.380 ;
        RECT 1948.020 1413.370 1951.020 1413.380 ;
        RECT 2128.020 1413.370 2131.020 1413.380 ;
        RECT 2308.020 1413.370 2311.020 1413.380 ;
        RECT 2488.020 1413.370 2491.020 1413.380 ;
        RECT 2668.020 1413.370 2671.020 1413.380 ;
        RECT 2848.020 1413.370 2851.020 1413.380 ;
        RECT 2959.500 1413.370 2962.500 1413.380 ;
        RECT -33.480 1398.380 -30.480 1398.390 ;
        RECT 130.020 1398.380 133.020 1398.390 ;
        RECT 397.840 1398.380 399.440 1398.390 ;
        RECT 1570.020 1398.380 1573.020 1398.390 ;
        RECT 1750.020 1398.380 1753.020 1398.390 ;
        RECT 1930.020 1398.380 1933.020 1398.390 ;
        RECT 2110.020 1398.380 2113.020 1398.390 ;
        RECT 2290.020 1398.380 2293.020 1398.390 ;
        RECT 2470.020 1398.380 2473.020 1398.390 ;
        RECT 2650.020 1398.380 2653.020 1398.390 ;
        RECT 2830.020 1398.380 2833.020 1398.390 ;
        RECT 2950.100 1398.380 2953.100 1398.390 ;
        RECT -33.480 1395.380 2953.100 1398.380 ;
        RECT -33.480 1395.370 -30.480 1395.380 ;
        RECT 130.020 1395.370 133.020 1395.380 ;
        RECT 397.840 1395.370 399.440 1395.380 ;
        RECT 1570.020 1395.370 1573.020 1395.380 ;
        RECT 1750.020 1395.370 1753.020 1395.380 ;
        RECT 1930.020 1395.370 1933.020 1395.380 ;
        RECT 2110.020 1395.370 2113.020 1395.380 ;
        RECT 2290.020 1395.370 2293.020 1395.380 ;
        RECT 2470.020 1395.370 2473.020 1395.380 ;
        RECT 2650.020 1395.370 2653.020 1395.380 ;
        RECT 2830.020 1395.370 2833.020 1395.380 ;
        RECT 2950.100 1395.370 2953.100 1395.380 ;
        RECT -24.080 1380.380 -21.080 1380.390 ;
        RECT 112.020 1380.380 115.020 1380.390 ;
        RECT 397.840 1380.380 399.440 1380.390 ;
        RECT 1552.020 1380.380 1555.020 1380.390 ;
        RECT 1732.020 1380.380 1735.020 1380.390 ;
        RECT 1912.020 1380.380 1915.020 1380.390 ;
        RECT 2092.020 1380.380 2095.020 1380.390 ;
        RECT 2272.020 1380.380 2275.020 1380.390 ;
        RECT 2452.020 1380.380 2455.020 1380.390 ;
        RECT 2632.020 1380.380 2635.020 1380.390 ;
        RECT 2812.020 1380.380 2815.020 1380.390 ;
        RECT 2940.700 1380.380 2943.700 1380.390 ;
        RECT -24.080 1377.380 2943.700 1380.380 ;
        RECT -24.080 1377.370 -21.080 1377.380 ;
        RECT 112.020 1377.370 115.020 1377.380 ;
        RECT 397.840 1377.370 399.440 1377.380 ;
        RECT 1552.020 1377.370 1555.020 1377.380 ;
        RECT 1732.020 1377.370 1735.020 1377.380 ;
        RECT 1912.020 1377.370 1915.020 1377.380 ;
        RECT 2092.020 1377.370 2095.020 1377.380 ;
        RECT 2272.020 1377.370 2275.020 1377.380 ;
        RECT 2452.020 1377.370 2455.020 1377.380 ;
        RECT 2632.020 1377.370 2635.020 1377.380 ;
        RECT 2812.020 1377.370 2815.020 1377.380 ;
        RECT 2940.700 1377.370 2943.700 1377.380 ;
        RECT -14.680 1362.380 -11.680 1362.390 ;
        RECT 94.020 1362.380 97.020 1362.390 ;
        RECT 274.020 1362.380 277.020 1362.390 ;
        RECT 397.840 1362.380 399.440 1362.390 ;
        RECT 1534.020 1362.380 1537.020 1362.390 ;
        RECT 1714.020 1362.380 1717.020 1362.390 ;
        RECT 1894.020 1362.380 1897.020 1362.390 ;
        RECT 2074.020 1362.380 2077.020 1362.390 ;
        RECT 2254.020 1362.380 2257.020 1362.390 ;
        RECT 2434.020 1362.380 2437.020 1362.390 ;
        RECT 2614.020 1362.380 2617.020 1362.390 ;
        RECT 2794.020 1362.380 2797.020 1362.390 ;
        RECT 2931.300 1362.380 2934.300 1362.390 ;
        RECT -14.680 1359.380 2934.300 1362.380 ;
        RECT -14.680 1359.370 -11.680 1359.380 ;
        RECT 94.020 1359.370 97.020 1359.380 ;
        RECT 274.020 1359.370 277.020 1359.380 ;
        RECT 397.840 1359.370 399.440 1359.380 ;
        RECT 1534.020 1359.370 1537.020 1359.380 ;
        RECT 1714.020 1359.370 1717.020 1359.380 ;
        RECT 1894.020 1359.370 1897.020 1359.380 ;
        RECT 2074.020 1359.370 2077.020 1359.380 ;
        RECT 2254.020 1359.370 2257.020 1359.380 ;
        RECT 2434.020 1359.370 2437.020 1359.380 ;
        RECT 2614.020 1359.370 2617.020 1359.380 ;
        RECT 2794.020 1359.370 2797.020 1359.380 ;
        RECT 2931.300 1359.370 2934.300 1359.380 ;
        RECT -42.880 1236.380 -39.880 1236.390 ;
        RECT 148.020 1236.380 151.020 1236.390 ;
        RECT 397.840 1236.380 399.440 1236.390 ;
        RECT 1588.020 1236.380 1591.020 1236.390 ;
        RECT 1768.020 1236.380 1771.020 1236.390 ;
        RECT 1948.020 1236.380 1951.020 1236.390 ;
        RECT 2128.020 1236.380 2131.020 1236.390 ;
        RECT 2308.020 1236.380 2311.020 1236.390 ;
        RECT 2488.020 1236.380 2491.020 1236.390 ;
        RECT 2668.020 1236.380 2671.020 1236.390 ;
        RECT 2848.020 1236.380 2851.020 1236.390 ;
        RECT 2959.500 1236.380 2962.500 1236.390 ;
        RECT -42.880 1233.380 2962.500 1236.380 ;
        RECT -42.880 1233.370 -39.880 1233.380 ;
        RECT 148.020 1233.370 151.020 1233.380 ;
        RECT 397.840 1233.370 399.440 1233.380 ;
        RECT 1588.020 1233.370 1591.020 1233.380 ;
        RECT 1768.020 1233.370 1771.020 1233.380 ;
        RECT 1948.020 1233.370 1951.020 1233.380 ;
        RECT 2128.020 1233.370 2131.020 1233.380 ;
        RECT 2308.020 1233.370 2311.020 1233.380 ;
        RECT 2488.020 1233.370 2491.020 1233.380 ;
        RECT 2668.020 1233.370 2671.020 1233.380 ;
        RECT 2848.020 1233.370 2851.020 1233.380 ;
        RECT 2959.500 1233.370 2962.500 1233.380 ;
        RECT -33.480 1218.380 -30.480 1218.390 ;
        RECT 130.020 1218.380 133.020 1218.390 ;
        RECT 397.840 1218.380 399.440 1218.390 ;
        RECT 1570.020 1218.380 1573.020 1218.390 ;
        RECT 1750.020 1218.380 1753.020 1218.390 ;
        RECT 1930.020 1218.380 1933.020 1218.390 ;
        RECT 2110.020 1218.380 2113.020 1218.390 ;
        RECT 2290.020 1218.380 2293.020 1218.390 ;
        RECT 2470.020 1218.380 2473.020 1218.390 ;
        RECT 2650.020 1218.380 2653.020 1218.390 ;
        RECT 2830.020 1218.380 2833.020 1218.390 ;
        RECT 2950.100 1218.380 2953.100 1218.390 ;
        RECT -33.480 1215.380 2953.100 1218.380 ;
        RECT -33.480 1215.370 -30.480 1215.380 ;
        RECT 130.020 1215.370 133.020 1215.380 ;
        RECT 397.840 1215.370 399.440 1215.380 ;
        RECT 1570.020 1215.370 1573.020 1215.380 ;
        RECT 1750.020 1215.370 1753.020 1215.380 ;
        RECT 1930.020 1215.370 1933.020 1215.380 ;
        RECT 2110.020 1215.370 2113.020 1215.380 ;
        RECT 2290.020 1215.370 2293.020 1215.380 ;
        RECT 2470.020 1215.370 2473.020 1215.380 ;
        RECT 2650.020 1215.370 2653.020 1215.380 ;
        RECT 2830.020 1215.370 2833.020 1215.380 ;
        RECT 2950.100 1215.370 2953.100 1215.380 ;
        RECT -24.080 1200.380 -21.080 1200.390 ;
        RECT 112.020 1200.380 115.020 1200.390 ;
        RECT 397.840 1200.380 399.440 1200.390 ;
        RECT 1552.020 1200.380 1555.020 1200.390 ;
        RECT 1732.020 1200.380 1735.020 1200.390 ;
        RECT 1912.020 1200.380 1915.020 1200.390 ;
        RECT 2092.020 1200.380 2095.020 1200.390 ;
        RECT 2272.020 1200.380 2275.020 1200.390 ;
        RECT 2452.020 1200.380 2455.020 1200.390 ;
        RECT 2632.020 1200.380 2635.020 1200.390 ;
        RECT 2812.020 1200.380 2815.020 1200.390 ;
        RECT 2940.700 1200.380 2943.700 1200.390 ;
        RECT -24.080 1197.380 2943.700 1200.380 ;
        RECT -24.080 1197.370 -21.080 1197.380 ;
        RECT 112.020 1197.370 115.020 1197.380 ;
        RECT 397.840 1197.370 399.440 1197.380 ;
        RECT 1552.020 1197.370 1555.020 1197.380 ;
        RECT 1732.020 1197.370 1735.020 1197.380 ;
        RECT 1912.020 1197.370 1915.020 1197.380 ;
        RECT 2092.020 1197.370 2095.020 1197.380 ;
        RECT 2272.020 1197.370 2275.020 1197.380 ;
        RECT 2452.020 1197.370 2455.020 1197.380 ;
        RECT 2632.020 1197.370 2635.020 1197.380 ;
        RECT 2812.020 1197.370 2815.020 1197.380 ;
        RECT 2940.700 1197.370 2943.700 1197.380 ;
        RECT -14.680 1182.380 -11.680 1182.390 ;
        RECT 94.020 1182.380 97.020 1182.390 ;
        RECT 274.020 1182.380 277.020 1182.390 ;
        RECT 397.840 1182.380 399.440 1182.390 ;
        RECT 1534.020 1182.380 1537.020 1182.390 ;
        RECT 1714.020 1182.380 1717.020 1182.390 ;
        RECT 1894.020 1182.380 1897.020 1182.390 ;
        RECT 2074.020 1182.380 2077.020 1182.390 ;
        RECT 2254.020 1182.380 2257.020 1182.390 ;
        RECT 2434.020 1182.380 2437.020 1182.390 ;
        RECT 2614.020 1182.380 2617.020 1182.390 ;
        RECT 2794.020 1182.380 2797.020 1182.390 ;
        RECT 2931.300 1182.380 2934.300 1182.390 ;
        RECT -14.680 1179.380 2934.300 1182.380 ;
        RECT -14.680 1179.370 -11.680 1179.380 ;
        RECT 94.020 1179.370 97.020 1179.380 ;
        RECT 274.020 1179.370 277.020 1179.380 ;
        RECT 397.840 1179.370 399.440 1179.380 ;
        RECT 1534.020 1179.370 1537.020 1179.380 ;
        RECT 1714.020 1179.370 1717.020 1179.380 ;
        RECT 1894.020 1179.370 1897.020 1179.380 ;
        RECT 2074.020 1179.370 2077.020 1179.380 ;
        RECT 2254.020 1179.370 2257.020 1179.380 ;
        RECT 2434.020 1179.370 2437.020 1179.380 ;
        RECT 2614.020 1179.370 2617.020 1179.380 ;
        RECT 2794.020 1179.370 2797.020 1179.380 ;
        RECT 2931.300 1179.370 2934.300 1179.380 ;
        RECT -42.880 1056.380 -39.880 1056.390 ;
        RECT 148.020 1056.380 151.020 1056.390 ;
        RECT 397.840 1056.380 399.440 1056.390 ;
        RECT 1588.020 1056.380 1591.020 1056.390 ;
        RECT 1768.020 1056.380 1771.020 1056.390 ;
        RECT 1948.020 1056.380 1951.020 1056.390 ;
        RECT 2128.020 1056.380 2131.020 1056.390 ;
        RECT 2308.020 1056.380 2311.020 1056.390 ;
        RECT 2488.020 1056.380 2491.020 1056.390 ;
        RECT 2668.020 1056.380 2671.020 1056.390 ;
        RECT 2848.020 1056.380 2851.020 1056.390 ;
        RECT 2959.500 1056.380 2962.500 1056.390 ;
        RECT -42.880 1053.380 2962.500 1056.380 ;
        RECT -42.880 1053.370 -39.880 1053.380 ;
        RECT 148.020 1053.370 151.020 1053.380 ;
        RECT 397.840 1053.370 399.440 1053.380 ;
        RECT 1588.020 1053.370 1591.020 1053.380 ;
        RECT 1768.020 1053.370 1771.020 1053.380 ;
        RECT 1948.020 1053.370 1951.020 1053.380 ;
        RECT 2128.020 1053.370 2131.020 1053.380 ;
        RECT 2308.020 1053.370 2311.020 1053.380 ;
        RECT 2488.020 1053.370 2491.020 1053.380 ;
        RECT 2668.020 1053.370 2671.020 1053.380 ;
        RECT 2848.020 1053.370 2851.020 1053.380 ;
        RECT 2959.500 1053.370 2962.500 1053.380 ;
        RECT -33.480 1038.380 -30.480 1038.390 ;
        RECT 130.020 1038.380 133.020 1038.390 ;
        RECT 397.840 1038.380 399.440 1038.390 ;
        RECT 1570.020 1038.380 1573.020 1038.390 ;
        RECT 1750.020 1038.380 1753.020 1038.390 ;
        RECT 1930.020 1038.380 1933.020 1038.390 ;
        RECT 2110.020 1038.380 2113.020 1038.390 ;
        RECT 2290.020 1038.380 2293.020 1038.390 ;
        RECT 2470.020 1038.380 2473.020 1038.390 ;
        RECT 2650.020 1038.380 2653.020 1038.390 ;
        RECT 2830.020 1038.380 2833.020 1038.390 ;
        RECT 2950.100 1038.380 2953.100 1038.390 ;
        RECT -33.480 1035.380 2953.100 1038.380 ;
        RECT -33.480 1035.370 -30.480 1035.380 ;
        RECT 130.020 1035.370 133.020 1035.380 ;
        RECT 397.840 1035.370 399.440 1035.380 ;
        RECT 1570.020 1035.370 1573.020 1035.380 ;
        RECT 1750.020 1035.370 1753.020 1035.380 ;
        RECT 1930.020 1035.370 1933.020 1035.380 ;
        RECT 2110.020 1035.370 2113.020 1035.380 ;
        RECT 2290.020 1035.370 2293.020 1035.380 ;
        RECT 2470.020 1035.370 2473.020 1035.380 ;
        RECT 2650.020 1035.370 2653.020 1035.380 ;
        RECT 2830.020 1035.370 2833.020 1035.380 ;
        RECT 2950.100 1035.370 2953.100 1035.380 ;
        RECT -24.080 1020.380 -21.080 1020.390 ;
        RECT 112.020 1020.380 115.020 1020.390 ;
        RECT 397.840 1020.380 399.440 1020.390 ;
        RECT 1552.020 1020.380 1555.020 1020.390 ;
        RECT 1732.020 1020.380 1735.020 1020.390 ;
        RECT 1912.020 1020.380 1915.020 1020.390 ;
        RECT 2092.020 1020.380 2095.020 1020.390 ;
        RECT 2272.020 1020.380 2275.020 1020.390 ;
        RECT 2452.020 1020.380 2455.020 1020.390 ;
        RECT 2632.020 1020.380 2635.020 1020.390 ;
        RECT 2812.020 1020.380 2815.020 1020.390 ;
        RECT 2940.700 1020.380 2943.700 1020.390 ;
        RECT -24.080 1017.380 2943.700 1020.380 ;
        RECT -24.080 1017.370 -21.080 1017.380 ;
        RECT 112.020 1017.370 115.020 1017.380 ;
        RECT 397.840 1017.370 399.440 1017.380 ;
        RECT 1552.020 1017.370 1555.020 1017.380 ;
        RECT 1732.020 1017.370 1735.020 1017.380 ;
        RECT 1912.020 1017.370 1915.020 1017.380 ;
        RECT 2092.020 1017.370 2095.020 1017.380 ;
        RECT 2272.020 1017.370 2275.020 1017.380 ;
        RECT 2452.020 1017.370 2455.020 1017.380 ;
        RECT 2632.020 1017.370 2635.020 1017.380 ;
        RECT 2812.020 1017.370 2815.020 1017.380 ;
        RECT 2940.700 1017.370 2943.700 1017.380 ;
        RECT -14.680 1002.380 -11.680 1002.390 ;
        RECT 94.020 1002.380 97.020 1002.390 ;
        RECT 274.020 1002.380 277.020 1002.390 ;
        RECT 1534.020 1002.380 1537.020 1002.390 ;
        RECT 1714.020 1002.380 1717.020 1002.390 ;
        RECT 1894.020 1002.380 1897.020 1002.390 ;
        RECT 2074.020 1002.380 2077.020 1002.390 ;
        RECT 2254.020 1002.380 2257.020 1002.390 ;
        RECT 2434.020 1002.380 2437.020 1002.390 ;
        RECT 2614.020 1002.380 2617.020 1002.390 ;
        RECT 2794.020 1002.380 2797.020 1002.390 ;
        RECT 2931.300 1002.380 2934.300 1002.390 ;
        RECT -14.680 999.380 2934.300 1002.380 ;
        RECT -14.680 999.370 -11.680 999.380 ;
        RECT 94.020 999.370 97.020 999.380 ;
        RECT 274.020 999.370 277.020 999.380 ;
        RECT 1534.020 999.370 1537.020 999.380 ;
        RECT 1714.020 999.370 1717.020 999.380 ;
        RECT 1894.020 999.370 1897.020 999.380 ;
        RECT 2074.020 999.370 2077.020 999.380 ;
        RECT 2254.020 999.370 2257.020 999.380 ;
        RECT 2434.020 999.370 2437.020 999.380 ;
        RECT 2614.020 999.370 2617.020 999.380 ;
        RECT 2794.020 999.370 2797.020 999.380 ;
        RECT 2931.300 999.370 2934.300 999.380 ;
        RECT -42.880 876.380 -39.880 876.390 ;
        RECT 148.020 876.380 151.020 876.390 ;
        RECT 328.020 876.380 331.020 876.390 ;
        RECT 508.020 876.380 511.020 876.390 ;
        RECT 688.020 876.380 691.020 876.390 ;
        RECT 868.020 876.380 871.020 876.390 ;
        RECT 1048.020 876.380 1051.020 876.390 ;
        RECT 1228.020 876.380 1231.020 876.390 ;
        RECT 1408.020 876.380 1411.020 876.390 ;
        RECT 1588.020 876.380 1591.020 876.390 ;
        RECT 1768.020 876.380 1771.020 876.390 ;
        RECT 1948.020 876.380 1951.020 876.390 ;
        RECT 2128.020 876.380 2131.020 876.390 ;
        RECT 2308.020 876.380 2311.020 876.390 ;
        RECT 2488.020 876.380 2491.020 876.390 ;
        RECT 2668.020 876.380 2671.020 876.390 ;
        RECT 2848.020 876.380 2851.020 876.390 ;
        RECT 2959.500 876.380 2962.500 876.390 ;
        RECT -42.880 873.380 2962.500 876.380 ;
        RECT -42.880 873.370 -39.880 873.380 ;
        RECT 148.020 873.370 151.020 873.380 ;
        RECT 328.020 873.370 331.020 873.380 ;
        RECT 508.020 873.370 511.020 873.380 ;
        RECT 688.020 873.370 691.020 873.380 ;
        RECT 868.020 873.370 871.020 873.380 ;
        RECT 1048.020 873.370 1051.020 873.380 ;
        RECT 1228.020 873.370 1231.020 873.380 ;
        RECT 1408.020 873.370 1411.020 873.380 ;
        RECT 1588.020 873.370 1591.020 873.380 ;
        RECT 1768.020 873.370 1771.020 873.380 ;
        RECT 1948.020 873.370 1951.020 873.380 ;
        RECT 2128.020 873.370 2131.020 873.380 ;
        RECT 2308.020 873.370 2311.020 873.380 ;
        RECT 2488.020 873.370 2491.020 873.380 ;
        RECT 2668.020 873.370 2671.020 873.380 ;
        RECT 2848.020 873.370 2851.020 873.380 ;
        RECT 2959.500 873.370 2962.500 873.380 ;
        RECT -33.480 858.380 -30.480 858.390 ;
        RECT 130.020 858.380 133.020 858.390 ;
        RECT 310.020 858.380 313.020 858.390 ;
        RECT 490.020 858.380 493.020 858.390 ;
        RECT 670.020 858.380 673.020 858.390 ;
        RECT 850.020 858.380 853.020 858.390 ;
        RECT 1030.020 858.380 1033.020 858.390 ;
        RECT 1210.020 858.380 1213.020 858.390 ;
        RECT 1390.020 858.380 1393.020 858.390 ;
        RECT 1570.020 858.380 1573.020 858.390 ;
        RECT 1750.020 858.380 1753.020 858.390 ;
        RECT 1930.020 858.380 1933.020 858.390 ;
        RECT 2110.020 858.380 2113.020 858.390 ;
        RECT 2290.020 858.380 2293.020 858.390 ;
        RECT 2470.020 858.380 2473.020 858.390 ;
        RECT 2650.020 858.380 2653.020 858.390 ;
        RECT 2830.020 858.380 2833.020 858.390 ;
        RECT 2950.100 858.380 2953.100 858.390 ;
        RECT -33.480 855.380 2953.100 858.380 ;
        RECT -33.480 855.370 -30.480 855.380 ;
        RECT 130.020 855.370 133.020 855.380 ;
        RECT 310.020 855.370 313.020 855.380 ;
        RECT 490.020 855.370 493.020 855.380 ;
        RECT 670.020 855.370 673.020 855.380 ;
        RECT 850.020 855.370 853.020 855.380 ;
        RECT 1030.020 855.370 1033.020 855.380 ;
        RECT 1210.020 855.370 1213.020 855.380 ;
        RECT 1390.020 855.370 1393.020 855.380 ;
        RECT 1570.020 855.370 1573.020 855.380 ;
        RECT 1750.020 855.370 1753.020 855.380 ;
        RECT 1930.020 855.370 1933.020 855.380 ;
        RECT 2110.020 855.370 2113.020 855.380 ;
        RECT 2290.020 855.370 2293.020 855.380 ;
        RECT 2470.020 855.370 2473.020 855.380 ;
        RECT 2650.020 855.370 2653.020 855.380 ;
        RECT 2830.020 855.370 2833.020 855.380 ;
        RECT 2950.100 855.370 2953.100 855.380 ;
        RECT -24.080 840.380 -21.080 840.390 ;
        RECT 112.020 840.380 115.020 840.390 ;
        RECT 292.020 840.380 295.020 840.390 ;
        RECT 472.020 840.380 475.020 840.390 ;
        RECT 652.020 840.380 655.020 840.390 ;
        RECT 832.020 840.380 835.020 840.390 ;
        RECT 1012.020 840.380 1015.020 840.390 ;
        RECT 1192.020 840.380 1195.020 840.390 ;
        RECT 1372.020 840.380 1375.020 840.390 ;
        RECT 1552.020 840.380 1555.020 840.390 ;
        RECT 1732.020 840.380 1735.020 840.390 ;
        RECT 1912.020 840.380 1915.020 840.390 ;
        RECT 2092.020 840.380 2095.020 840.390 ;
        RECT 2272.020 840.380 2275.020 840.390 ;
        RECT 2452.020 840.380 2455.020 840.390 ;
        RECT 2632.020 840.380 2635.020 840.390 ;
        RECT 2812.020 840.380 2815.020 840.390 ;
        RECT 2940.700 840.380 2943.700 840.390 ;
        RECT -24.080 837.380 2943.700 840.380 ;
        RECT -24.080 837.370 -21.080 837.380 ;
        RECT 112.020 837.370 115.020 837.380 ;
        RECT 292.020 837.370 295.020 837.380 ;
        RECT 472.020 837.370 475.020 837.380 ;
        RECT 652.020 837.370 655.020 837.380 ;
        RECT 832.020 837.370 835.020 837.380 ;
        RECT 1012.020 837.370 1015.020 837.380 ;
        RECT 1192.020 837.370 1195.020 837.380 ;
        RECT 1372.020 837.370 1375.020 837.380 ;
        RECT 1552.020 837.370 1555.020 837.380 ;
        RECT 1732.020 837.370 1735.020 837.380 ;
        RECT 1912.020 837.370 1915.020 837.380 ;
        RECT 2092.020 837.370 2095.020 837.380 ;
        RECT 2272.020 837.370 2275.020 837.380 ;
        RECT 2452.020 837.370 2455.020 837.380 ;
        RECT 2632.020 837.370 2635.020 837.380 ;
        RECT 2812.020 837.370 2815.020 837.380 ;
        RECT 2940.700 837.370 2943.700 837.380 ;
        RECT -14.680 822.380 -11.680 822.390 ;
        RECT 94.020 822.380 97.020 822.390 ;
        RECT 274.020 822.380 277.020 822.390 ;
        RECT 454.020 822.380 457.020 822.390 ;
        RECT 634.020 822.380 637.020 822.390 ;
        RECT 814.020 822.380 817.020 822.390 ;
        RECT 994.020 822.380 997.020 822.390 ;
        RECT 1174.020 822.380 1177.020 822.390 ;
        RECT 1354.020 822.380 1357.020 822.390 ;
        RECT 1534.020 822.380 1537.020 822.390 ;
        RECT 1714.020 822.380 1717.020 822.390 ;
        RECT 1894.020 822.380 1897.020 822.390 ;
        RECT 2074.020 822.380 2077.020 822.390 ;
        RECT 2254.020 822.380 2257.020 822.390 ;
        RECT 2434.020 822.380 2437.020 822.390 ;
        RECT 2614.020 822.380 2617.020 822.390 ;
        RECT 2794.020 822.380 2797.020 822.390 ;
        RECT 2931.300 822.380 2934.300 822.390 ;
        RECT -14.680 819.380 2934.300 822.380 ;
        RECT -14.680 819.370 -11.680 819.380 ;
        RECT 94.020 819.370 97.020 819.380 ;
        RECT 274.020 819.370 277.020 819.380 ;
        RECT 454.020 819.370 457.020 819.380 ;
        RECT 634.020 819.370 637.020 819.380 ;
        RECT 814.020 819.370 817.020 819.380 ;
        RECT 994.020 819.370 997.020 819.380 ;
        RECT 1174.020 819.370 1177.020 819.380 ;
        RECT 1354.020 819.370 1357.020 819.380 ;
        RECT 1534.020 819.370 1537.020 819.380 ;
        RECT 1714.020 819.370 1717.020 819.380 ;
        RECT 1894.020 819.370 1897.020 819.380 ;
        RECT 2074.020 819.370 2077.020 819.380 ;
        RECT 2254.020 819.370 2257.020 819.380 ;
        RECT 2434.020 819.370 2437.020 819.380 ;
        RECT 2614.020 819.370 2617.020 819.380 ;
        RECT 2794.020 819.370 2797.020 819.380 ;
        RECT 2931.300 819.370 2934.300 819.380 ;
        RECT -42.880 696.380 -39.880 696.390 ;
        RECT 148.020 696.380 151.020 696.390 ;
        RECT 328.020 696.380 331.020 696.390 ;
        RECT 508.020 696.380 511.020 696.390 ;
        RECT 688.020 696.380 691.020 696.390 ;
        RECT 868.020 696.380 871.020 696.390 ;
        RECT 1048.020 696.380 1051.020 696.390 ;
        RECT 1228.020 696.380 1231.020 696.390 ;
        RECT 1408.020 696.380 1411.020 696.390 ;
        RECT 1588.020 696.380 1591.020 696.390 ;
        RECT 1768.020 696.380 1771.020 696.390 ;
        RECT 1948.020 696.380 1951.020 696.390 ;
        RECT 2128.020 696.380 2131.020 696.390 ;
        RECT 2308.020 696.380 2311.020 696.390 ;
        RECT 2488.020 696.380 2491.020 696.390 ;
        RECT 2668.020 696.380 2671.020 696.390 ;
        RECT 2848.020 696.380 2851.020 696.390 ;
        RECT 2959.500 696.380 2962.500 696.390 ;
        RECT -42.880 693.380 2962.500 696.380 ;
        RECT -42.880 693.370 -39.880 693.380 ;
        RECT 148.020 693.370 151.020 693.380 ;
        RECT 328.020 693.370 331.020 693.380 ;
        RECT 508.020 693.370 511.020 693.380 ;
        RECT 688.020 693.370 691.020 693.380 ;
        RECT 868.020 693.370 871.020 693.380 ;
        RECT 1048.020 693.370 1051.020 693.380 ;
        RECT 1228.020 693.370 1231.020 693.380 ;
        RECT 1408.020 693.370 1411.020 693.380 ;
        RECT 1588.020 693.370 1591.020 693.380 ;
        RECT 1768.020 693.370 1771.020 693.380 ;
        RECT 1948.020 693.370 1951.020 693.380 ;
        RECT 2128.020 693.370 2131.020 693.380 ;
        RECT 2308.020 693.370 2311.020 693.380 ;
        RECT 2488.020 693.370 2491.020 693.380 ;
        RECT 2668.020 693.370 2671.020 693.380 ;
        RECT 2848.020 693.370 2851.020 693.380 ;
        RECT 2959.500 693.370 2962.500 693.380 ;
        RECT -33.480 678.380 -30.480 678.390 ;
        RECT 130.020 678.380 133.020 678.390 ;
        RECT 310.020 678.380 313.020 678.390 ;
        RECT 490.020 678.380 493.020 678.390 ;
        RECT 670.020 678.380 673.020 678.390 ;
        RECT 850.020 678.380 853.020 678.390 ;
        RECT 1030.020 678.380 1033.020 678.390 ;
        RECT 1210.020 678.380 1213.020 678.390 ;
        RECT 1390.020 678.380 1393.020 678.390 ;
        RECT 1570.020 678.380 1573.020 678.390 ;
        RECT 1750.020 678.380 1753.020 678.390 ;
        RECT 1930.020 678.380 1933.020 678.390 ;
        RECT 2110.020 678.380 2113.020 678.390 ;
        RECT 2290.020 678.380 2293.020 678.390 ;
        RECT 2470.020 678.380 2473.020 678.390 ;
        RECT 2650.020 678.380 2653.020 678.390 ;
        RECT 2830.020 678.380 2833.020 678.390 ;
        RECT 2950.100 678.380 2953.100 678.390 ;
        RECT -33.480 675.380 2953.100 678.380 ;
        RECT -33.480 675.370 -30.480 675.380 ;
        RECT 130.020 675.370 133.020 675.380 ;
        RECT 310.020 675.370 313.020 675.380 ;
        RECT 490.020 675.370 493.020 675.380 ;
        RECT 670.020 675.370 673.020 675.380 ;
        RECT 850.020 675.370 853.020 675.380 ;
        RECT 1030.020 675.370 1033.020 675.380 ;
        RECT 1210.020 675.370 1213.020 675.380 ;
        RECT 1390.020 675.370 1393.020 675.380 ;
        RECT 1570.020 675.370 1573.020 675.380 ;
        RECT 1750.020 675.370 1753.020 675.380 ;
        RECT 1930.020 675.370 1933.020 675.380 ;
        RECT 2110.020 675.370 2113.020 675.380 ;
        RECT 2290.020 675.370 2293.020 675.380 ;
        RECT 2470.020 675.370 2473.020 675.380 ;
        RECT 2650.020 675.370 2653.020 675.380 ;
        RECT 2830.020 675.370 2833.020 675.380 ;
        RECT 2950.100 675.370 2953.100 675.380 ;
        RECT -24.080 660.380 -21.080 660.390 ;
        RECT 112.020 660.380 115.020 660.390 ;
        RECT 292.020 660.380 295.020 660.390 ;
        RECT 472.020 660.380 475.020 660.390 ;
        RECT 652.020 660.380 655.020 660.390 ;
        RECT 832.020 660.380 835.020 660.390 ;
        RECT 1012.020 660.380 1015.020 660.390 ;
        RECT 1192.020 660.380 1195.020 660.390 ;
        RECT 1372.020 660.380 1375.020 660.390 ;
        RECT 1552.020 660.380 1555.020 660.390 ;
        RECT 1732.020 660.380 1735.020 660.390 ;
        RECT 1912.020 660.380 1915.020 660.390 ;
        RECT 2092.020 660.380 2095.020 660.390 ;
        RECT 2272.020 660.380 2275.020 660.390 ;
        RECT 2452.020 660.380 2455.020 660.390 ;
        RECT 2632.020 660.380 2635.020 660.390 ;
        RECT 2812.020 660.380 2815.020 660.390 ;
        RECT 2940.700 660.380 2943.700 660.390 ;
        RECT -24.080 657.380 2943.700 660.380 ;
        RECT -24.080 657.370 -21.080 657.380 ;
        RECT 112.020 657.370 115.020 657.380 ;
        RECT 292.020 657.370 295.020 657.380 ;
        RECT 472.020 657.370 475.020 657.380 ;
        RECT 652.020 657.370 655.020 657.380 ;
        RECT 832.020 657.370 835.020 657.380 ;
        RECT 1012.020 657.370 1015.020 657.380 ;
        RECT 1192.020 657.370 1195.020 657.380 ;
        RECT 1372.020 657.370 1375.020 657.380 ;
        RECT 1552.020 657.370 1555.020 657.380 ;
        RECT 1732.020 657.370 1735.020 657.380 ;
        RECT 1912.020 657.370 1915.020 657.380 ;
        RECT 2092.020 657.370 2095.020 657.380 ;
        RECT 2272.020 657.370 2275.020 657.380 ;
        RECT 2452.020 657.370 2455.020 657.380 ;
        RECT 2632.020 657.370 2635.020 657.380 ;
        RECT 2812.020 657.370 2815.020 657.380 ;
        RECT 2940.700 657.370 2943.700 657.380 ;
        RECT -14.680 642.380 -11.680 642.390 ;
        RECT 94.020 642.380 97.020 642.390 ;
        RECT 274.020 642.380 277.020 642.390 ;
        RECT 454.020 642.380 457.020 642.390 ;
        RECT 634.020 642.380 637.020 642.390 ;
        RECT 814.020 642.380 817.020 642.390 ;
        RECT 994.020 642.380 997.020 642.390 ;
        RECT 1174.020 642.380 1177.020 642.390 ;
        RECT 1354.020 642.380 1357.020 642.390 ;
        RECT 1534.020 642.380 1537.020 642.390 ;
        RECT 1714.020 642.380 1717.020 642.390 ;
        RECT 1894.020 642.380 1897.020 642.390 ;
        RECT 2074.020 642.380 2077.020 642.390 ;
        RECT 2254.020 642.380 2257.020 642.390 ;
        RECT 2434.020 642.380 2437.020 642.390 ;
        RECT 2614.020 642.380 2617.020 642.390 ;
        RECT 2794.020 642.380 2797.020 642.390 ;
        RECT 2931.300 642.380 2934.300 642.390 ;
        RECT -14.680 639.380 2934.300 642.380 ;
        RECT -14.680 639.370 -11.680 639.380 ;
        RECT 94.020 639.370 97.020 639.380 ;
        RECT 274.020 639.370 277.020 639.380 ;
        RECT 454.020 639.370 457.020 639.380 ;
        RECT 634.020 639.370 637.020 639.380 ;
        RECT 814.020 639.370 817.020 639.380 ;
        RECT 994.020 639.370 997.020 639.380 ;
        RECT 1174.020 639.370 1177.020 639.380 ;
        RECT 1354.020 639.370 1357.020 639.380 ;
        RECT 1534.020 639.370 1537.020 639.380 ;
        RECT 1714.020 639.370 1717.020 639.380 ;
        RECT 1894.020 639.370 1897.020 639.380 ;
        RECT 2074.020 639.370 2077.020 639.380 ;
        RECT 2254.020 639.370 2257.020 639.380 ;
        RECT 2434.020 639.370 2437.020 639.380 ;
        RECT 2614.020 639.370 2617.020 639.380 ;
        RECT 2794.020 639.370 2797.020 639.380 ;
        RECT 2931.300 639.370 2934.300 639.380 ;
        RECT -42.880 516.380 -39.880 516.390 ;
        RECT 148.020 516.380 151.020 516.390 ;
        RECT 328.020 516.380 331.020 516.390 ;
        RECT 508.020 516.380 511.020 516.390 ;
        RECT 688.020 516.380 691.020 516.390 ;
        RECT 868.020 516.380 871.020 516.390 ;
        RECT 1048.020 516.380 1051.020 516.390 ;
        RECT 1228.020 516.380 1231.020 516.390 ;
        RECT 1408.020 516.380 1411.020 516.390 ;
        RECT 1588.020 516.380 1591.020 516.390 ;
        RECT 1768.020 516.380 1771.020 516.390 ;
        RECT 1948.020 516.380 1951.020 516.390 ;
        RECT 2128.020 516.380 2131.020 516.390 ;
        RECT 2308.020 516.380 2311.020 516.390 ;
        RECT 2488.020 516.380 2491.020 516.390 ;
        RECT 2668.020 516.380 2671.020 516.390 ;
        RECT 2848.020 516.380 2851.020 516.390 ;
        RECT 2959.500 516.380 2962.500 516.390 ;
        RECT -42.880 513.380 2962.500 516.380 ;
        RECT -42.880 513.370 -39.880 513.380 ;
        RECT 148.020 513.370 151.020 513.380 ;
        RECT 328.020 513.370 331.020 513.380 ;
        RECT 508.020 513.370 511.020 513.380 ;
        RECT 688.020 513.370 691.020 513.380 ;
        RECT 868.020 513.370 871.020 513.380 ;
        RECT 1048.020 513.370 1051.020 513.380 ;
        RECT 1228.020 513.370 1231.020 513.380 ;
        RECT 1408.020 513.370 1411.020 513.380 ;
        RECT 1588.020 513.370 1591.020 513.380 ;
        RECT 1768.020 513.370 1771.020 513.380 ;
        RECT 1948.020 513.370 1951.020 513.380 ;
        RECT 2128.020 513.370 2131.020 513.380 ;
        RECT 2308.020 513.370 2311.020 513.380 ;
        RECT 2488.020 513.370 2491.020 513.380 ;
        RECT 2668.020 513.370 2671.020 513.380 ;
        RECT 2848.020 513.370 2851.020 513.380 ;
        RECT 2959.500 513.370 2962.500 513.380 ;
        RECT -33.480 498.380 -30.480 498.390 ;
        RECT 130.020 498.380 133.020 498.390 ;
        RECT 310.020 498.380 313.020 498.390 ;
        RECT 490.020 498.380 493.020 498.390 ;
        RECT 670.020 498.380 673.020 498.390 ;
        RECT 850.020 498.380 853.020 498.390 ;
        RECT 1030.020 498.380 1033.020 498.390 ;
        RECT 1210.020 498.380 1213.020 498.390 ;
        RECT 1390.020 498.380 1393.020 498.390 ;
        RECT 1570.020 498.380 1573.020 498.390 ;
        RECT 1750.020 498.380 1753.020 498.390 ;
        RECT 1930.020 498.380 1933.020 498.390 ;
        RECT 2110.020 498.380 2113.020 498.390 ;
        RECT 2290.020 498.380 2293.020 498.390 ;
        RECT 2470.020 498.380 2473.020 498.390 ;
        RECT 2650.020 498.380 2653.020 498.390 ;
        RECT 2830.020 498.380 2833.020 498.390 ;
        RECT 2950.100 498.380 2953.100 498.390 ;
        RECT -33.480 495.380 2953.100 498.380 ;
        RECT -33.480 495.370 -30.480 495.380 ;
        RECT 130.020 495.370 133.020 495.380 ;
        RECT 310.020 495.370 313.020 495.380 ;
        RECT 490.020 495.370 493.020 495.380 ;
        RECT 670.020 495.370 673.020 495.380 ;
        RECT 850.020 495.370 853.020 495.380 ;
        RECT 1030.020 495.370 1033.020 495.380 ;
        RECT 1210.020 495.370 1213.020 495.380 ;
        RECT 1390.020 495.370 1393.020 495.380 ;
        RECT 1570.020 495.370 1573.020 495.380 ;
        RECT 1750.020 495.370 1753.020 495.380 ;
        RECT 1930.020 495.370 1933.020 495.380 ;
        RECT 2110.020 495.370 2113.020 495.380 ;
        RECT 2290.020 495.370 2293.020 495.380 ;
        RECT 2470.020 495.370 2473.020 495.380 ;
        RECT 2650.020 495.370 2653.020 495.380 ;
        RECT 2830.020 495.370 2833.020 495.380 ;
        RECT 2950.100 495.370 2953.100 495.380 ;
        RECT -24.080 480.380 -21.080 480.390 ;
        RECT 112.020 480.380 115.020 480.390 ;
        RECT 292.020 480.380 295.020 480.390 ;
        RECT 472.020 480.380 475.020 480.390 ;
        RECT 652.020 480.380 655.020 480.390 ;
        RECT 832.020 480.380 835.020 480.390 ;
        RECT 1012.020 480.380 1015.020 480.390 ;
        RECT 1192.020 480.380 1195.020 480.390 ;
        RECT 1372.020 480.380 1375.020 480.390 ;
        RECT 1552.020 480.380 1555.020 480.390 ;
        RECT 1732.020 480.380 1735.020 480.390 ;
        RECT 1912.020 480.380 1915.020 480.390 ;
        RECT 2092.020 480.380 2095.020 480.390 ;
        RECT 2272.020 480.380 2275.020 480.390 ;
        RECT 2452.020 480.380 2455.020 480.390 ;
        RECT 2632.020 480.380 2635.020 480.390 ;
        RECT 2812.020 480.380 2815.020 480.390 ;
        RECT 2940.700 480.380 2943.700 480.390 ;
        RECT -24.080 477.380 2943.700 480.380 ;
        RECT -24.080 477.370 -21.080 477.380 ;
        RECT 112.020 477.370 115.020 477.380 ;
        RECT 292.020 477.370 295.020 477.380 ;
        RECT 472.020 477.370 475.020 477.380 ;
        RECT 652.020 477.370 655.020 477.380 ;
        RECT 832.020 477.370 835.020 477.380 ;
        RECT 1012.020 477.370 1015.020 477.380 ;
        RECT 1192.020 477.370 1195.020 477.380 ;
        RECT 1372.020 477.370 1375.020 477.380 ;
        RECT 1552.020 477.370 1555.020 477.380 ;
        RECT 1732.020 477.370 1735.020 477.380 ;
        RECT 1912.020 477.370 1915.020 477.380 ;
        RECT 2092.020 477.370 2095.020 477.380 ;
        RECT 2272.020 477.370 2275.020 477.380 ;
        RECT 2452.020 477.370 2455.020 477.380 ;
        RECT 2632.020 477.370 2635.020 477.380 ;
        RECT 2812.020 477.370 2815.020 477.380 ;
        RECT 2940.700 477.370 2943.700 477.380 ;
        RECT -14.680 462.380 -11.680 462.390 ;
        RECT 94.020 462.380 97.020 462.390 ;
        RECT 274.020 462.380 277.020 462.390 ;
        RECT 454.020 462.380 457.020 462.390 ;
        RECT 634.020 462.380 637.020 462.390 ;
        RECT 814.020 462.380 817.020 462.390 ;
        RECT 994.020 462.380 997.020 462.390 ;
        RECT 1174.020 462.380 1177.020 462.390 ;
        RECT 1354.020 462.380 1357.020 462.390 ;
        RECT 1534.020 462.380 1537.020 462.390 ;
        RECT 1714.020 462.380 1717.020 462.390 ;
        RECT 1894.020 462.380 1897.020 462.390 ;
        RECT 2074.020 462.380 2077.020 462.390 ;
        RECT 2254.020 462.380 2257.020 462.390 ;
        RECT 2434.020 462.380 2437.020 462.390 ;
        RECT 2614.020 462.380 2617.020 462.390 ;
        RECT 2794.020 462.380 2797.020 462.390 ;
        RECT 2931.300 462.380 2934.300 462.390 ;
        RECT -14.680 459.380 2934.300 462.380 ;
        RECT -14.680 459.370 -11.680 459.380 ;
        RECT 94.020 459.370 97.020 459.380 ;
        RECT 274.020 459.370 277.020 459.380 ;
        RECT 454.020 459.370 457.020 459.380 ;
        RECT 634.020 459.370 637.020 459.380 ;
        RECT 814.020 459.370 817.020 459.380 ;
        RECT 994.020 459.370 997.020 459.380 ;
        RECT 1174.020 459.370 1177.020 459.380 ;
        RECT 1354.020 459.370 1357.020 459.380 ;
        RECT 1534.020 459.370 1537.020 459.380 ;
        RECT 1714.020 459.370 1717.020 459.380 ;
        RECT 1894.020 459.370 1897.020 459.380 ;
        RECT 2074.020 459.370 2077.020 459.380 ;
        RECT 2254.020 459.370 2257.020 459.380 ;
        RECT 2434.020 459.370 2437.020 459.380 ;
        RECT 2614.020 459.370 2617.020 459.380 ;
        RECT 2794.020 459.370 2797.020 459.380 ;
        RECT 2931.300 459.370 2934.300 459.380 ;
        RECT -42.880 336.380 -39.880 336.390 ;
        RECT 148.020 336.380 151.020 336.390 ;
        RECT 328.020 336.380 331.020 336.390 ;
        RECT 508.020 336.380 511.020 336.390 ;
        RECT 688.020 336.380 691.020 336.390 ;
        RECT 868.020 336.380 871.020 336.390 ;
        RECT 1048.020 336.380 1051.020 336.390 ;
        RECT 1228.020 336.380 1231.020 336.390 ;
        RECT 1408.020 336.380 1411.020 336.390 ;
        RECT 1588.020 336.380 1591.020 336.390 ;
        RECT 1768.020 336.380 1771.020 336.390 ;
        RECT 1948.020 336.380 1951.020 336.390 ;
        RECT 2128.020 336.380 2131.020 336.390 ;
        RECT 2308.020 336.380 2311.020 336.390 ;
        RECT 2488.020 336.380 2491.020 336.390 ;
        RECT 2668.020 336.380 2671.020 336.390 ;
        RECT 2848.020 336.380 2851.020 336.390 ;
        RECT 2959.500 336.380 2962.500 336.390 ;
        RECT -42.880 333.380 2962.500 336.380 ;
        RECT -42.880 333.370 -39.880 333.380 ;
        RECT 148.020 333.370 151.020 333.380 ;
        RECT 328.020 333.370 331.020 333.380 ;
        RECT 508.020 333.370 511.020 333.380 ;
        RECT 688.020 333.370 691.020 333.380 ;
        RECT 868.020 333.370 871.020 333.380 ;
        RECT 1048.020 333.370 1051.020 333.380 ;
        RECT 1228.020 333.370 1231.020 333.380 ;
        RECT 1408.020 333.370 1411.020 333.380 ;
        RECT 1588.020 333.370 1591.020 333.380 ;
        RECT 1768.020 333.370 1771.020 333.380 ;
        RECT 1948.020 333.370 1951.020 333.380 ;
        RECT 2128.020 333.370 2131.020 333.380 ;
        RECT 2308.020 333.370 2311.020 333.380 ;
        RECT 2488.020 333.370 2491.020 333.380 ;
        RECT 2668.020 333.370 2671.020 333.380 ;
        RECT 2848.020 333.370 2851.020 333.380 ;
        RECT 2959.500 333.370 2962.500 333.380 ;
        RECT -33.480 318.380 -30.480 318.390 ;
        RECT 130.020 318.380 133.020 318.390 ;
        RECT 310.020 318.380 313.020 318.390 ;
        RECT 490.020 318.380 493.020 318.390 ;
        RECT 670.020 318.380 673.020 318.390 ;
        RECT 850.020 318.380 853.020 318.390 ;
        RECT 1030.020 318.380 1033.020 318.390 ;
        RECT 1210.020 318.380 1213.020 318.390 ;
        RECT 1390.020 318.380 1393.020 318.390 ;
        RECT 1570.020 318.380 1573.020 318.390 ;
        RECT 1750.020 318.380 1753.020 318.390 ;
        RECT 1930.020 318.380 1933.020 318.390 ;
        RECT 2110.020 318.380 2113.020 318.390 ;
        RECT 2290.020 318.380 2293.020 318.390 ;
        RECT 2470.020 318.380 2473.020 318.390 ;
        RECT 2650.020 318.380 2653.020 318.390 ;
        RECT 2830.020 318.380 2833.020 318.390 ;
        RECT 2950.100 318.380 2953.100 318.390 ;
        RECT -33.480 315.380 2953.100 318.380 ;
        RECT -33.480 315.370 -30.480 315.380 ;
        RECT 130.020 315.370 133.020 315.380 ;
        RECT 310.020 315.370 313.020 315.380 ;
        RECT 490.020 315.370 493.020 315.380 ;
        RECT 670.020 315.370 673.020 315.380 ;
        RECT 850.020 315.370 853.020 315.380 ;
        RECT 1030.020 315.370 1033.020 315.380 ;
        RECT 1210.020 315.370 1213.020 315.380 ;
        RECT 1390.020 315.370 1393.020 315.380 ;
        RECT 1570.020 315.370 1573.020 315.380 ;
        RECT 1750.020 315.370 1753.020 315.380 ;
        RECT 1930.020 315.370 1933.020 315.380 ;
        RECT 2110.020 315.370 2113.020 315.380 ;
        RECT 2290.020 315.370 2293.020 315.380 ;
        RECT 2470.020 315.370 2473.020 315.380 ;
        RECT 2650.020 315.370 2653.020 315.380 ;
        RECT 2830.020 315.370 2833.020 315.380 ;
        RECT 2950.100 315.370 2953.100 315.380 ;
        RECT -24.080 300.380 -21.080 300.390 ;
        RECT 112.020 300.380 115.020 300.390 ;
        RECT 292.020 300.380 295.020 300.390 ;
        RECT 472.020 300.380 475.020 300.390 ;
        RECT 652.020 300.380 655.020 300.390 ;
        RECT 832.020 300.380 835.020 300.390 ;
        RECT 1012.020 300.380 1015.020 300.390 ;
        RECT 1192.020 300.380 1195.020 300.390 ;
        RECT 1372.020 300.380 1375.020 300.390 ;
        RECT 1552.020 300.380 1555.020 300.390 ;
        RECT 1732.020 300.380 1735.020 300.390 ;
        RECT 1912.020 300.380 1915.020 300.390 ;
        RECT 2092.020 300.380 2095.020 300.390 ;
        RECT 2272.020 300.380 2275.020 300.390 ;
        RECT 2452.020 300.380 2455.020 300.390 ;
        RECT 2632.020 300.380 2635.020 300.390 ;
        RECT 2812.020 300.380 2815.020 300.390 ;
        RECT 2940.700 300.380 2943.700 300.390 ;
        RECT -24.080 297.380 2943.700 300.380 ;
        RECT -24.080 297.370 -21.080 297.380 ;
        RECT 112.020 297.370 115.020 297.380 ;
        RECT 292.020 297.370 295.020 297.380 ;
        RECT 472.020 297.370 475.020 297.380 ;
        RECT 652.020 297.370 655.020 297.380 ;
        RECT 832.020 297.370 835.020 297.380 ;
        RECT 1012.020 297.370 1015.020 297.380 ;
        RECT 1192.020 297.370 1195.020 297.380 ;
        RECT 1372.020 297.370 1375.020 297.380 ;
        RECT 1552.020 297.370 1555.020 297.380 ;
        RECT 1732.020 297.370 1735.020 297.380 ;
        RECT 1912.020 297.370 1915.020 297.380 ;
        RECT 2092.020 297.370 2095.020 297.380 ;
        RECT 2272.020 297.370 2275.020 297.380 ;
        RECT 2452.020 297.370 2455.020 297.380 ;
        RECT 2632.020 297.370 2635.020 297.380 ;
        RECT 2812.020 297.370 2815.020 297.380 ;
        RECT 2940.700 297.370 2943.700 297.380 ;
        RECT -14.680 282.380 -11.680 282.390 ;
        RECT 94.020 282.380 97.020 282.390 ;
        RECT 274.020 282.380 277.020 282.390 ;
        RECT 454.020 282.380 457.020 282.390 ;
        RECT 634.020 282.380 637.020 282.390 ;
        RECT 814.020 282.380 817.020 282.390 ;
        RECT 994.020 282.380 997.020 282.390 ;
        RECT 1174.020 282.380 1177.020 282.390 ;
        RECT 1354.020 282.380 1357.020 282.390 ;
        RECT 1534.020 282.380 1537.020 282.390 ;
        RECT 1714.020 282.380 1717.020 282.390 ;
        RECT 1894.020 282.380 1897.020 282.390 ;
        RECT 2074.020 282.380 2077.020 282.390 ;
        RECT 2254.020 282.380 2257.020 282.390 ;
        RECT 2434.020 282.380 2437.020 282.390 ;
        RECT 2614.020 282.380 2617.020 282.390 ;
        RECT 2794.020 282.380 2797.020 282.390 ;
        RECT 2931.300 282.380 2934.300 282.390 ;
        RECT -14.680 279.380 2934.300 282.380 ;
        RECT -14.680 279.370 -11.680 279.380 ;
        RECT 94.020 279.370 97.020 279.380 ;
        RECT 274.020 279.370 277.020 279.380 ;
        RECT 454.020 279.370 457.020 279.380 ;
        RECT 634.020 279.370 637.020 279.380 ;
        RECT 814.020 279.370 817.020 279.380 ;
        RECT 994.020 279.370 997.020 279.380 ;
        RECT 1174.020 279.370 1177.020 279.380 ;
        RECT 1354.020 279.370 1357.020 279.380 ;
        RECT 1534.020 279.370 1537.020 279.380 ;
        RECT 1714.020 279.370 1717.020 279.380 ;
        RECT 1894.020 279.370 1897.020 279.380 ;
        RECT 2074.020 279.370 2077.020 279.380 ;
        RECT 2254.020 279.370 2257.020 279.380 ;
        RECT 2434.020 279.370 2437.020 279.380 ;
        RECT 2614.020 279.370 2617.020 279.380 ;
        RECT 2794.020 279.370 2797.020 279.380 ;
        RECT 2931.300 279.370 2934.300 279.380 ;
        RECT -42.880 156.380 -39.880 156.390 ;
        RECT 148.020 156.380 151.020 156.390 ;
        RECT 328.020 156.380 331.020 156.390 ;
        RECT 508.020 156.380 511.020 156.390 ;
        RECT 688.020 156.380 691.020 156.390 ;
        RECT 868.020 156.380 871.020 156.390 ;
        RECT 1048.020 156.380 1051.020 156.390 ;
        RECT 1228.020 156.380 1231.020 156.390 ;
        RECT 1408.020 156.380 1411.020 156.390 ;
        RECT 1588.020 156.380 1591.020 156.390 ;
        RECT 1768.020 156.380 1771.020 156.390 ;
        RECT 1948.020 156.380 1951.020 156.390 ;
        RECT 2128.020 156.380 2131.020 156.390 ;
        RECT 2308.020 156.380 2311.020 156.390 ;
        RECT 2488.020 156.380 2491.020 156.390 ;
        RECT 2668.020 156.380 2671.020 156.390 ;
        RECT 2848.020 156.380 2851.020 156.390 ;
        RECT 2959.500 156.380 2962.500 156.390 ;
        RECT -42.880 153.380 2962.500 156.380 ;
        RECT -42.880 153.370 -39.880 153.380 ;
        RECT 148.020 153.370 151.020 153.380 ;
        RECT 328.020 153.370 331.020 153.380 ;
        RECT 508.020 153.370 511.020 153.380 ;
        RECT 688.020 153.370 691.020 153.380 ;
        RECT 868.020 153.370 871.020 153.380 ;
        RECT 1048.020 153.370 1051.020 153.380 ;
        RECT 1228.020 153.370 1231.020 153.380 ;
        RECT 1408.020 153.370 1411.020 153.380 ;
        RECT 1588.020 153.370 1591.020 153.380 ;
        RECT 1768.020 153.370 1771.020 153.380 ;
        RECT 1948.020 153.370 1951.020 153.380 ;
        RECT 2128.020 153.370 2131.020 153.380 ;
        RECT 2308.020 153.370 2311.020 153.380 ;
        RECT 2488.020 153.370 2491.020 153.380 ;
        RECT 2668.020 153.370 2671.020 153.380 ;
        RECT 2848.020 153.370 2851.020 153.380 ;
        RECT 2959.500 153.370 2962.500 153.380 ;
        RECT -33.480 138.380 -30.480 138.390 ;
        RECT 130.020 138.380 133.020 138.390 ;
        RECT 310.020 138.380 313.020 138.390 ;
        RECT 490.020 138.380 493.020 138.390 ;
        RECT 670.020 138.380 673.020 138.390 ;
        RECT 850.020 138.380 853.020 138.390 ;
        RECT 1030.020 138.380 1033.020 138.390 ;
        RECT 1210.020 138.380 1213.020 138.390 ;
        RECT 1390.020 138.380 1393.020 138.390 ;
        RECT 1570.020 138.380 1573.020 138.390 ;
        RECT 1750.020 138.380 1753.020 138.390 ;
        RECT 1930.020 138.380 1933.020 138.390 ;
        RECT 2110.020 138.380 2113.020 138.390 ;
        RECT 2290.020 138.380 2293.020 138.390 ;
        RECT 2470.020 138.380 2473.020 138.390 ;
        RECT 2650.020 138.380 2653.020 138.390 ;
        RECT 2830.020 138.380 2833.020 138.390 ;
        RECT 2950.100 138.380 2953.100 138.390 ;
        RECT -33.480 135.380 2953.100 138.380 ;
        RECT -33.480 135.370 -30.480 135.380 ;
        RECT 130.020 135.370 133.020 135.380 ;
        RECT 310.020 135.370 313.020 135.380 ;
        RECT 490.020 135.370 493.020 135.380 ;
        RECT 670.020 135.370 673.020 135.380 ;
        RECT 850.020 135.370 853.020 135.380 ;
        RECT 1030.020 135.370 1033.020 135.380 ;
        RECT 1210.020 135.370 1213.020 135.380 ;
        RECT 1390.020 135.370 1393.020 135.380 ;
        RECT 1570.020 135.370 1573.020 135.380 ;
        RECT 1750.020 135.370 1753.020 135.380 ;
        RECT 1930.020 135.370 1933.020 135.380 ;
        RECT 2110.020 135.370 2113.020 135.380 ;
        RECT 2290.020 135.370 2293.020 135.380 ;
        RECT 2470.020 135.370 2473.020 135.380 ;
        RECT 2650.020 135.370 2653.020 135.380 ;
        RECT 2830.020 135.370 2833.020 135.380 ;
        RECT 2950.100 135.370 2953.100 135.380 ;
        RECT -24.080 120.380 -21.080 120.390 ;
        RECT 112.020 120.380 115.020 120.390 ;
        RECT 292.020 120.380 295.020 120.390 ;
        RECT 472.020 120.380 475.020 120.390 ;
        RECT 652.020 120.380 655.020 120.390 ;
        RECT 832.020 120.380 835.020 120.390 ;
        RECT 1012.020 120.380 1015.020 120.390 ;
        RECT 1192.020 120.380 1195.020 120.390 ;
        RECT 1372.020 120.380 1375.020 120.390 ;
        RECT 1552.020 120.380 1555.020 120.390 ;
        RECT 1732.020 120.380 1735.020 120.390 ;
        RECT 1912.020 120.380 1915.020 120.390 ;
        RECT 2092.020 120.380 2095.020 120.390 ;
        RECT 2272.020 120.380 2275.020 120.390 ;
        RECT 2452.020 120.380 2455.020 120.390 ;
        RECT 2632.020 120.380 2635.020 120.390 ;
        RECT 2812.020 120.380 2815.020 120.390 ;
        RECT 2940.700 120.380 2943.700 120.390 ;
        RECT -24.080 117.380 2943.700 120.380 ;
        RECT -24.080 117.370 -21.080 117.380 ;
        RECT 112.020 117.370 115.020 117.380 ;
        RECT 292.020 117.370 295.020 117.380 ;
        RECT 472.020 117.370 475.020 117.380 ;
        RECT 652.020 117.370 655.020 117.380 ;
        RECT 832.020 117.370 835.020 117.380 ;
        RECT 1012.020 117.370 1015.020 117.380 ;
        RECT 1192.020 117.370 1195.020 117.380 ;
        RECT 1372.020 117.370 1375.020 117.380 ;
        RECT 1552.020 117.370 1555.020 117.380 ;
        RECT 1732.020 117.370 1735.020 117.380 ;
        RECT 1912.020 117.370 1915.020 117.380 ;
        RECT 2092.020 117.370 2095.020 117.380 ;
        RECT 2272.020 117.370 2275.020 117.380 ;
        RECT 2452.020 117.370 2455.020 117.380 ;
        RECT 2632.020 117.370 2635.020 117.380 ;
        RECT 2812.020 117.370 2815.020 117.380 ;
        RECT 2940.700 117.370 2943.700 117.380 ;
        RECT -14.680 102.380 -11.680 102.390 ;
        RECT 94.020 102.380 97.020 102.390 ;
        RECT 274.020 102.380 277.020 102.390 ;
        RECT 454.020 102.380 457.020 102.390 ;
        RECT 634.020 102.380 637.020 102.390 ;
        RECT 814.020 102.380 817.020 102.390 ;
        RECT 994.020 102.380 997.020 102.390 ;
        RECT 1174.020 102.380 1177.020 102.390 ;
        RECT 1354.020 102.380 1357.020 102.390 ;
        RECT 1534.020 102.380 1537.020 102.390 ;
        RECT 1714.020 102.380 1717.020 102.390 ;
        RECT 1894.020 102.380 1897.020 102.390 ;
        RECT 2074.020 102.380 2077.020 102.390 ;
        RECT 2254.020 102.380 2257.020 102.390 ;
        RECT 2434.020 102.380 2437.020 102.390 ;
        RECT 2614.020 102.380 2617.020 102.390 ;
        RECT 2794.020 102.380 2797.020 102.390 ;
        RECT 2931.300 102.380 2934.300 102.390 ;
        RECT -14.680 99.380 2934.300 102.380 ;
        RECT -14.680 99.370 -11.680 99.380 ;
        RECT 94.020 99.370 97.020 99.380 ;
        RECT 274.020 99.370 277.020 99.380 ;
        RECT 454.020 99.370 457.020 99.380 ;
        RECT 634.020 99.370 637.020 99.380 ;
        RECT 814.020 99.370 817.020 99.380 ;
        RECT 994.020 99.370 997.020 99.380 ;
        RECT 1174.020 99.370 1177.020 99.380 ;
        RECT 1354.020 99.370 1357.020 99.380 ;
        RECT 1534.020 99.370 1537.020 99.380 ;
        RECT 1714.020 99.370 1717.020 99.380 ;
        RECT 1894.020 99.370 1897.020 99.380 ;
        RECT 2074.020 99.370 2077.020 99.380 ;
        RECT 2254.020 99.370 2257.020 99.380 ;
        RECT 2434.020 99.370 2437.020 99.380 ;
        RECT 2614.020 99.370 2617.020 99.380 ;
        RECT 2794.020 99.370 2797.020 99.380 ;
        RECT 2931.300 99.370 2934.300 99.380 ;
        RECT -14.680 -6.320 -11.680 -6.310 ;
        RECT 94.020 -6.320 97.020 -6.310 ;
        RECT 274.020 -6.320 277.020 -6.310 ;
        RECT 454.020 -6.320 457.020 -6.310 ;
        RECT 634.020 -6.320 637.020 -6.310 ;
        RECT 814.020 -6.320 817.020 -6.310 ;
        RECT 994.020 -6.320 997.020 -6.310 ;
        RECT 1174.020 -6.320 1177.020 -6.310 ;
        RECT 1354.020 -6.320 1357.020 -6.310 ;
        RECT 1534.020 -6.320 1537.020 -6.310 ;
        RECT 1714.020 -6.320 1717.020 -6.310 ;
        RECT 1894.020 -6.320 1897.020 -6.310 ;
        RECT 2074.020 -6.320 2077.020 -6.310 ;
        RECT 2254.020 -6.320 2257.020 -6.310 ;
        RECT 2434.020 -6.320 2437.020 -6.310 ;
        RECT 2614.020 -6.320 2617.020 -6.310 ;
        RECT 2794.020 -6.320 2797.020 -6.310 ;
        RECT 2931.300 -6.320 2934.300 -6.310 ;
        RECT -14.680 -9.320 2934.300 -6.320 ;
        RECT -14.680 -9.330 -11.680 -9.320 ;
        RECT 94.020 -9.330 97.020 -9.320 ;
        RECT 274.020 -9.330 277.020 -9.320 ;
        RECT 454.020 -9.330 457.020 -9.320 ;
        RECT 634.020 -9.330 637.020 -9.320 ;
        RECT 814.020 -9.330 817.020 -9.320 ;
        RECT 994.020 -9.330 997.020 -9.320 ;
        RECT 1174.020 -9.330 1177.020 -9.320 ;
        RECT 1354.020 -9.330 1357.020 -9.320 ;
        RECT 1534.020 -9.330 1537.020 -9.320 ;
        RECT 1714.020 -9.330 1717.020 -9.320 ;
        RECT 1894.020 -9.330 1897.020 -9.320 ;
        RECT 2074.020 -9.330 2077.020 -9.320 ;
        RECT 2254.020 -9.330 2257.020 -9.320 ;
        RECT 2434.020 -9.330 2437.020 -9.320 ;
        RECT 2614.020 -9.330 2617.020 -9.320 ;
        RECT 2794.020 -9.330 2797.020 -9.320 ;
        RECT 2931.300 -9.330 2934.300 -9.320 ;
        RECT -24.080 -15.720 -21.080 -15.710 ;
        RECT 112.020 -15.720 115.020 -15.710 ;
        RECT 292.020 -15.720 295.020 -15.710 ;
        RECT 472.020 -15.720 475.020 -15.710 ;
        RECT 652.020 -15.720 655.020 -15.710 ;
        RECT 832.020 -15.720 835.020 -15.710 ;
        RECT 1012.020 -15.720 1015.020 -15.710 ;
        RECT 1192.020 -15.720 1195.020 -15.710 ;
        RECT 1372.020 -15.720 1375.020 -15.710 ;
        RECT 1552.020 -15.720 1555.020 -15.710 ;
        RECT 1732.020 -15.720 1735.020 -15.710 ;
        RECT 1912.020 -15.720 1915.020 -15.710 ;
        RECT 2092.020 -15.720 2095.020 -15.710 ;
        RECT 2272.020 -15.720 2275.020 -15.710 ;
        RECT 2452.020 -15.720 2455.020 -15.710 ;
        RECT 2632.020 -15.720 2635.020 -15.710 ;
        RECT 2812.020 -15.720 2815.020 -15.710 ;
        RECT 2940.700 -15.720 2943.700 -15.710 ;
        RECT -24.080 -18.720 2943.700 -15.720 ;
        RECT -24.080 -18.730 -21.080 -18.720 ;
        RECT 112.020 -18.730 115.020 -18.720 ;
        RECT 292.020 -18.730 295.020 -18.720 ;
        RECT 472.020 -18.730 475.020 -18.720 ;
        RECT 652.020 -18.730 655.020 -18.720 ;
        RECT 832.020 -18.730 835.020 -18.720 ;
        RECT 1012.020 -18.730 1015.020 -18.720 ;
        RECT 1192.020 -18.730 1195.020 -18.720 ;
        RECT 1372.020 -18.730 1375.020 -18.720 ;
        RECT 1552.020 -18.730 1555.020 -18.720 ;
        RECT 1732.020 -18.730 1735.020 -18.720 ;
        RECT 1912.020 -18.730 1915.020 -18.720 ;
        RECT 2092.020 -18.730 2095.020 -18.720 ;
        RECT 2272.020 -18.730 2275.020 -18.720 ;
        RECT 2452.020 -18.730 2455.020 -18.720 ;
        RECT 2632.020 -18.730 2635.020 -18.720 ;
        RECT 2812.020 -18.730 2815.020 -18.720 ;
        RECT 2940.700 -18.730 2943.700 -18.720 ;
        RECT -33.480 -25.120 -30.480 -25.110 ;
        RECT 130.020 -25.120 133.020 -25.110 ;
        RECT 310.020 -25.120 313.020 -25.110 ;
        RECT 490.020 -25.120 493.020 -25.110 ;
        RECT 670.020 -25.120 673.020 -25.110 ;
        RECT 850.020 -25.120 853.020 -25.110 ;
        RECT 1030.020 -25.120 1033.020 -25.110 ;
        RECT 1210.020 -25.120 1213.020 -25.110 ;
        RECT 1390.020 -25.120 1393.020 -25.110 ;
        RECT 1570.020 -25.120 1573.020 -25.110 ;
        RECT 1750.020 -25.120 1753.020 -25.110 ;
        RECT 1930.020 -25.120 1933.020 -25.110 ;
        RECT 2110.020 -25.120 2113.020 -25.110 ;
        RECT 2290.020 -25.120 2293.020 -25.110 ;
        RECT 2470.020 -25.120 2473.020 -25.110 ;
        RECT 2650.020 -25.120 2653.020 -25.110 ;
        RECT 2830.020 -25.120 2833.020 -25.110 ;
        RECT 2950.100 -25.120 2953.100 -25.110 ;
        RECT -33.480 -28.120 2953.100 -25.120 ;
        RECT -33.480 -28.130 -30.480 -28.120 ;
        RECT 130.020 -28.130 133.020 -28.120 ;
        RECT 310.020 -28.130 313.020 -28.120 ;
        RECT 490.020 -28.130 493.020 -28.120 ;
        RECT 670.020 -28.130 673.020 -28.120 ;
        RECT 850.020 -28.130 853.020 -28.120 ;
        RECT 1030.020 -28.130 1033.020 -28.120 ;
        RECT 1210.020 -28.130 1213.020 -28.120 ;
        RECT 1390.020 -28.130 1393.020 -28.120 ;
        RECT 1570.020 -28.130 1573.020 -28.120 ;
        RECT 1750.020 -28.130 1753.020 -28.120 ;
        RECT 1930.020 -28.130 1933.020 -28.120 ;
        RECT 2110.020 -28.130 2113.020 -28.120 ;
        RECT 2290.020 -28.130 2293.020 -28.120 ;
        RECT 2470.020 -28.130 2473.020 -28.120 ;
        RECT 2650.020 -28.130 2653.020 -28.120 ;
        RECT 2830.020 -28.130 2833.020 -28.120 ;
        RECT 2950.100 -28.130 2953.100 -28.120 ;
        RECT -42.880 -34.520 -39.880 -34.510 ;
        RECT 148.020 -34.520 151.020 -34.510 ;
        RECT 328.020 -34.520 331.020 -34.510 ;
        RECT 508.020 -34.520 511.020 -34.510 ;
        RECT 688.020 -34.520 691.020 -34.510 ;
        RECT 868.020 -34.520 871.020 -34.510 ;
        RECT 1048.020 -34.520 1051.020 -34.510 ;
        RECT 1228.020 -34.520 1231.020 -34.510 ;
        RECT 1408.020 -34.520 1411.020 -34.510 ;
        RECT 1588.020 -34.520 1591.020 -34.510 ;
        RECT 1768.020 -34.520 1771.020 -34.510 ;
        RECT 1948.020 -34.520 1951.020 -34.510 ;
        RECT 2128.020 -34.520 2131.020 -34.510 ;
        RECT 2308.020 -34.520 2311.020 -34.510 ;
        RECT 2488.020 -34.520 2491.020 -34.510 ;
        RECT 2668.020 -34.520 2671.020 -34.510 ;
        RECT 2848.020 -34.520 2851.020 -34.510 ;
        RECT 2959.500 -34.520 2962.500 -34.510 ;
        RECT -42.880 -37.520 2962.500 -34.520 ;
        RECT -42.880 -37.530 -39.880 -37.520 ;
        RECT 148.020 -37.530 151.020 -37.520 ;
        RECT 328.020 -37.530 331.020 -37.520 ;
        RECT 508.020 -37.530 511.020 -37.520 ;
        RECT 688.020 -37.530 691.020 -37.520 ;
        RECT 868.020 -37.530 871.020 -37.520 ;
        RECT 1048.020 -37.530 1051.020 -37.520 ;
        RECT 1228.020 -37.530 1231.020 -37.520 ;
        RECT 1408.020 -37.530 1411.020 -37.520 ;
        RECT 1588.020 -37.530 1591.020 -37.520 ;
        RECT 1768.020 -37.530 1771.020 -37.520 ;
        RECT 1948.020 -37.530 1951.020 -37.520 ;
        RECT 2128.020 -37.530 2131.020 -37.520 ;
        RECT 2308.020 -37.530 2311.020 -37.520 ;
        RECT 2488.020 -37.530 2491.020 -37.520 ;
        RECT 2668.020 -37.530 2671.020 -37.520 ;
        RECT 2848.020 -37.530 2851.020 -37.520 ;
        RECT 2959.500 -37.530 2962.500 -37.520 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 305.000 2305.000 681.480 2751.235 ;
        RECT 955.000 2305.000 1331.480 2751.235 ;
        RECT 1555.000 2305.000 1931.480 2751.235 ;
        RECT 2205.000 2305.000 2581.480 2751.235 ;
        RECT 305.520 1010.795 1494.160 2188.725 ;
      LAYER met1 ;
        RECT 1318.890 2770.220 1319.210 2770.280 ;
        RECT 1892.510 2770.220 1892.830 2770.280 ;
        RECT 1318.890 2770.080 1892.830 2770.220 ;
        RECT 1318.890 2770.020 1319.210 2770.080 ;
        RECT 1892.510 2770.020 1892.830 2770.080 ;
        RECT 2539.270 2770.220 2539.590 2770.280 ;
        RECT 2566.870 2770.220 2567.190 2770.280 ;
        RECT 2539.270 2770.080 2567.190 2770.220 ;
        RECT 2539.270 2770.020 2539.590 2770.080 ;
        RECT 2566.870 2770.020 2567.190 2770.080 ;
        RECT 668.450 2767.160 668.770 2767.220 ;
        RECT 697.890 2767.160 698.210 2767.220 ;
        RECT 1295.890 2767.160 1296.210 2767.220 ;
        RECT 1318.890 2767.160 1319.210 2767.220 ;
        RECT 668.450 2767.020 1319.210 2767.160 ;
        RECT 668.450 2766.960 668.770 2767.020 ;
        RECT 697.890 2766.960 698.210 2767.020 ;
        RECT 1295.890 2766.960 1296.210 2767.020 ;
        RECT 1318.890 2766.960 1319.210 2767.020 ;
        RECT 1892.510 2767.160 1892.830 2767.220 ;
        RECT 1914.590 2767.160 1914.910 2767.220 ;
        RECT 1946.790 2767.160 1947.110 2767.220 ;
        RECT 2539.270 2767.160 2539.590 2767.220 ;
        RECT 1892.510 2767.020 2539.590 2767.160 ;
        RECT 1892.510 2766.960 1892.830 2767.020 ;
        RECT 1914.590 2766.960 1914.910 2767.020 ;
        RECT 1946.790 2766.960 1947.110 2767.020 ;
        RECT 2539.270 2766.960 2539.590 2767.020 ;
        RECT 696.970 2751.520 697.290 2751.580 ;
        RECT 1332.230 2751.520 1332.550 2751.580 ;
        RECT 696.970 2751.380 1332.550 2751.520 ;
        RECT 696.970 2751.320 697.290 2751.380 ;
        RECT 1332.230 2751.320 1332.550 2751.380 ;
        RECT 1511.170 2751.520 1511.490 2751.580 ;
        RECT 1945.870 2751.520 1946.190 2751.580 ;
        RECT 2582.050 2751.520 2582.370 2751.580 ;
        RECT 1511.170 2751.380 2582.370 2751.520 ;
        RECT 1511.170 2751.320 1511.490 2751.380 ;
        RECT 1945.870 2751.320 1946.190 2751.380 ;
        RECT 2582.050 2751.320 2582.370 2751.380 ;
      LAYER met1 ;
        RECT 305.000 2305.000 681.480 2751.235 ;
      LAYER met1 ;
        RECT 751.710 2732.480 752.030 2732.540 ;
        RECT 938.470 2732.480 938.790 2732.540 ;
        RECT 751.710 2732.340 938.790 2732.480 ;
        RECT 751.710 2732.280 752.030 2732.340 ;
        RECT 938.470 2732.280 938.790 2732.340 ;
        RECT 737.910 2725.680 738.230 2725.740 ;
        RECT 938.470 2725.680 938.790 2725.740 ;
        RECT 737.910 2725.540 938.790 2725.680 ;
        RECT 737.910 2725.480 738.230 2725.540 ;
        RECT 938.470 2725.480 938.790 2725.540 ;
        RECT 724.110 2718.880 724.430 2718.940 ;
        RECT 938.470 2718.880 938.790 2718.940 ;
        RECT 724.110 2718.740 938.790 2718.880 ;
        RECT 724.110 2718.680 724.430 2718.740 ;
        RECT 938.470 2718.680 938.790 2718.740 ;
        RECT 717.210 2712.080 717.530 2712.140 ;
        RECT 938.470 2712.080 938.790 2712.140 ;
        RECT 717.210 2711.940 938.790 2712.080 ;
        RECT 717.210 2711.880 717.530 2711.940 ;
        RECT 938.470 2711.880 938.790 2711.940 ;
        RECT 703.410 2698.480 703.730 2698.540 ;
        RECT 938.930 2698.480 939.250 2698.540 ;
        RECT 703.410 2698.340 939.250 2698.480 ;
        RECT 703.410 2698.280 703.730 2698.340 ;
        RECT 938.930 2698.280 939.250 2698.340 ;
        RECT 696.510 2698.140 696.830 2698.200 ;
        RECT 938.470 2698.140 938.790 2698.200 ;
        RECT 696.510 2698.000 938.790 2698.140 ;
        RECT 696.510 2697.940 696.830 2698.000 ;
        RECT 938.470 2697.940 938.790 2698.000 ;
      LAYER met1 ;
        RECT 955.000 2305.000 1331.480 2751.235 ;
      LAYER met1 ;
        RECT 1352.010 2746.420 1352.330 2746.480 ;
        RECT 1511.170 2746.420 1511.490 2746.480 ;
        RECT 1352.010 2746.280 1511.490 2746.420 ;
        RECT 1352.010 2746.220 1352.330 2746.280 ;
        RECT 1511.170 2746.220 1511.490 2746.280 ;
        RECT 1522.210 2725.680 1522.530 2725.740 ;
        RECT 1538.310 2725.680 1538.630 2725.740 ;
        RECT 1522.210 2725.540 1538.630 2725.680 ;
        RECT 1522.210 2725.480 1522.530 2725.540 ;
        RECT 1538.310 2725.480 1538.630 2725.540 ;
        RECT 1521.750 2712.080 1522.070 2712.140 ;
        RECT 1536.010 2712.080 1536.330 2712.140 ;
        RECT 1521.750 2711.940 1536.330 2712.080 ;
        RECT 1521.750 2711.880 1522.070 2711.940 ;
        RECT 1536.010 2711.880 1536.330 2711.940 ;
        RECT 1521.290 2698.140 1521.610 2698.200 ;
        RECT 1538.310 2698.140 1538.630 2698.200 ;
        RECT 1521.290 2698.000 1538.630 2698.140 ;
        RECT 1521.290 2697.940 1521.610 2698.000 ;
        RECT 1538.310 2697.940 1538.630 2698.000 ;
        RECT 1345.570 2422.060 1345.890 2422.120 ;
        RECT 1514.390 2422.060 1514.710 2422.120 ;
        RECT 1345.570 2421.920 1514.710 2422.060 ;
        RECT 1345.570 2421.860 1345.890 2421.920 ;
        RECT 1514.390 2421.860 1514.710 2421.920 ;
        RECT 1514.850 2387.720 1515.170 2387.780 ;
        RECT 1535.550 2387.720 1535.870 2387.780 ;
        RECT 1514.850 2387.580 1535.870 2387.720 ;
        RECT 1514.850 2387.520 1515.170 2387.580 ;
        RECT 1535.550 2387.520 1535.870 2387.580 ;
      LAYER met1 ;
        RECT 1555.000 2305.000 1931.480 2751.235 ;
      LAYER met1 ;
        RECT 1997.390 2732.480 1997.710 2732.540 ;
        RECT 2187.370 2732.480 2187.690 2732.540 ;
        RECT 1997.390 2732.340 2187.690 2732.480 ;
        RECT 1997.390 2732.280 1997.710 2732.340 ;
        RECT 2187.370 2732.280 2187.690 2732.340 ;
        RECT 1990.490 2725.680 1990.810 2725.740 ;
        RECT 2187.370 2725.680 2187.690 2725.740 ;
        RECT 1990.490 2725.540 2187.690 2725.680 ;
        RECT 1990.490 2725.480 1990.810 2725.540 ;
        RECT 2187.370 2725.480 2187.690 2725.540 ;
        RECT 1976.690 2718.880 1977.010 2718.940 ;
        RECT 2187.370 2718.880 2187.690 2718.940 ;
        RECT 1976.690 2718.740 2187.690 2718.880 ;
        RECT 1976.690 2718.680 1977.010 2718.740 ;
        RECT 2187.370 2718.680 2187.690 2718.740 ;
        RECT 1969.790 2712.080 1970.110 2712.140 ;
        RECT 2187.370 2712.080 2187.690 2712.140 ;
        RECT 1969.790 2711.940 2187.690 2712.080 ;
        RECT 1969.790 2711.880 1970.110 2711.940 ;
        RECT 2187.370 2711.880 2187.690 2711.940 ;
        RECT 1962.890 2698.480 1963.210 2698.540 ;
        RECT 2187.830 2698.480 2188.150 2698.540 ;
        RECT 1962.890 2698.340 2188.150 2698.480 ;
        RECT 1962.890 2698.280 1963.210 2698.340 ;
        RECT 2187.830 2698.280 2188.150 2698.340 ;
        RECT 1955.990 2698.140 1956.310 2698.200 ;
        RECT 2187.370 2698.140 2187.690 2698.200 ;
        RECT 1955.990 2698.000 2187.690 2698.140 ;
        RECT 1955.990 2697.940 1956.310 2698.000 ;
        RECT 2187.370 2697.940 2187.690 2698.000 ;
        RECT 1942.190 2684.200 1942.510 2684.260 ;
        RECT 2187.370 2684.200 2187.690 2684.260 ;
        RECT 1942.190 2684.060 2187.690 2684.200 ;
        RECT 1942.190 2684.000 1942.510 2684.060 ;
        RECT 2187.370 2684.000 2187.690 2684.060 ;
        RECT 2011.190 2401.320 2011.510 2401.380 ;
        RECT 2187.370 2401.320 2187.690 2401.380 ;
        RECT 2011.190 2401.180 2187.690 2401.320 ;
        RECT 2011.190 2401.120 2011.510 2401.180 ;
        RECT 2187.370 2401.120 2187.690 2401.180 ;
      LAYER met1 ;
        RECT 2205.000 2305.000 2581.480 2751.235 ;
      LAYER met1 ;
        RECT 944.450 2301.020 944.770 2301.080 ;
        RECT 1514.850 2301.020 1515.170 2301.080 ;
        RECT 944.450 2300.880 1515.170 2301.020 ;
        RECT 944.450 2300.820 944.770 2300.880 ;
        RECT 1514.850 2300.820 1515.170 2300.880 ;
        RECT 299.070 2297.620 299.390 2297.680 ;
        RECT 944.450 2297.620 944.770 2297.680 ;
        RECT 299.070 2297.480 944.770 2297.620 ;
        RECT 299.070 2297.420 299.390 2297.480 ;
        RECT 944.450 2297.420 944.770 2297.480 ;
        RECT 1514.850 2297.620 1515.170 2297.680 ;
        RECT 2190.590 2297.620 2190.910 2297.680 ;
        RECT 1514.850 2297.480 2190.910 2297.620 ;
        RECT 1514.850 2297.420 1515.170 2297.480 ;
        RECT 2190.590 2297.420 2190.910 2297.480 ;
        RECT 1514.390 2297.280 1514.710 2297.340 ;
        RECT 1945.870 2297.280 1946.190 2297.340 ;
        RECT 1514.390 2297.140 1946.190 2297.280 ;
        RECT 1514.390 2297.080 1514.710 2297.140 ;
        RECT 1945.870 2297.080 1946.190 2297.140 ;
        RECT 386.470 2290.820 386.790 2290.880 ;
        RECT 431.550 2290.820 431.870 2290.880 ;
        RECT 434.310 2290.820 434.630 2290.880 ;
        RECT 386.470 2290.680 434.630 2290.820 ;
        RECT 386.470 2290.620 386.790 2290.680 ;
        RECT 431.550 2290.620 431.870 2290.680 ;
        RECT 434.310 2290.620 434.630 2290.680 ;
        RECT 496.870 2290.820 497.190 2290.880 ;
        RECT 526.770 2290.820 527.090 2290.880 ;
        RECT 496.870 2290.680 527.090 2290.820 ;
        RECT 496.870 2290.620 497.190 2290.680 ;
        RECT 526.770 2290.620 527.090 2290.680 ;
        RECT 613.710 2290.820 614.030 2290.880 ;
        RECT 635.330 2290.820 635.650 2290.880 ;
        RECT 613.710 2290.680 635.650 2290.820 ;
        RECT 613.710 2290.620 614.030 2290.680 ;
        RECT 635.330 2290.620 635.650 2290.680 ;
        RECT 710.310 2290.820 710.630 2290.880 ;
        RECT 734.690 2290.820 735.010 2290.880 ;
        RECT 710.310 2290.680 735.010 2290.820 ;
        RECT 710.310 2290.620 710.630 2290.680 ;
        RECT 734.690 2290.620 735.010 2290.680 ;
        RECT 806.910 2290.820 807.230 2290.880 ;
        RECT 952.270 2290.820 952.590 2290.880 ;
        RECT 806.910 2290.680 952.590 2290.820 ;
        RECT 806.910 2290.620 807.230 2290.680 ;
        RECT 952.270 2290.620 952.590 2290.680 ;
        RECT 1000.110 2290.820 1000.430 2290.880 ;
        RECT 1048.870 2290.820 1049.190 2290.880 ;
        RECT 1000.110 2290.680 1049.190 2290.820 ;
        RECT 1000.110 2290.620 1000.430 2290.680 ;
        RECT 1048.870 2290.620 1049.190 2290.680 ;
        RECT 1076.470 2290.820 1076.790 2290.880 ;
        RECT 1086.130 2290.820 1086.450 2290.880 ;
        RECT 1076.470 2290.680 1086.450 2290.820 ;
        RECT 1076.470 2290.620 1076.790 2290.680 ;
        RECT 1086.130 2290.620 1086.450 2290.680 ;
        RECT 1096.710 2290.820 1097.030 2290.880 ;
        RECT 1131.670 2290.820 1131.990 2290.880 ;
        RECT 1096.710 2290.680 1131.990 2290.820 ;
        RECT 1096.710 2290.620 1097.030 2290.680 ;
        RECT 1131.670 2290.620 1131.990 2290.680 ;
        RECT 1676.770 2290.820 1677.090 2290.880 ;
        RECT 1723.690 2290.820 1724.010 2290.880 ;
        RECT 1766.470 2290.820 1766.790 2290.880 ;
        RECT 1676.770 2290.680 1766.790 2290.820 ;
        RECT 1676.770 2290.620 1677.090 2290.680 ;
        RECT 1723.690 2290.620 1724.010 2290.680 ;
        RECT 1766.470 2290.620 1766.790 2290.680 ;
        RECT 1770.150 2290.820 1770.470 2290.880 ;
        RECT 2421.970 2290.820 2422.290 2290.880 ;
        RECT 1770.150 2290.680 2422.290 2290.820 ;
        RECT 1770.150 2290.620 1770.470 2290.680 ;
        RECT 2421.970 2290.620 2422.290 2290.680 ;
        RECT 399.810 2290.480 400.130 2290.540 ;
        RECT 445.350 2290.480 445.670 2290.540 ;
        RECT 399.810 2290.340 445.670 2290.480 ;
        RECT 399.810 2290.280 400.130 2290.340 ;
        RECT 445.350 2290.280 445.670 2290.340 ;
        RECT 455.470 2290.480 455.790 2290.540 ;
        RECT 502.850 2290.480 503.170 2290.540 ;
        RECT 455.470 2290.340 503.170 2290.480 ;
        RECT 455.470 2290.280 455.790 2290.340 ;
        RECT 502.850 2290.280 503.170 2290.340 ;
        RECT 538.270 2290.480 538.590 2290.540 ;
        RECT 1117.870 2290.480 1118.190 2290.540 ;
        RECT 538.270 2290.340 1118.190 2290.480 ;
        RECT 538.270 2290.280 538.590 2290.340 ;
        RECT 1117.870 2290.280 1118.190 2290.340 ;
        RECT 1118.330 2290.480 1118.650 2290.540 ;
        RECT 1159.270 2290.480 1159.590 2290.540 ;
        RECT 1118.330 2290.340 1159.590 2290.480 ;
        RECT 1118.330 2290.280 1118.650 2290.340 ;
        RECT 1159.270 2290.280 1159.590 2290.340 ;
        RECT 1645.490 2290.480 1645.810 2290.540 ;
        RECT 1690.110 2290.480 1690.430 2290.540 ;
        RECT 1645.490 2290.340 1690.430 2290.480 ;
        RECT 1645.490 2290.280 1645.810 2290.340 ;
        RECT 1690.110 2290.280 1690.430 2290.340 ;
        RECT 1721.850 2290.480 1722.170 2290.540 ;
        RECT 1759.570 2290.480 1759.890 2290.540 ;
        RECT 1721.850 2290.340 1759.890 2290.480 ;
        RECT 1721.850 2290.280 1722.170 2290.340 ;
        RECT 1759.570 2290.280 1759.890 2290.340 ;
        RECT 1763.710 2290.480 1764.030 2290.540 ;
        RECT 2415.070 2290.480 2415.390 2290.540 ;
        RECT 1763.710 2290.340 2415.390 2290.480 ;
        RECT 1763.710 2290.280 1764.030 2290.340 ;
        RECT 2415.070 2290.280 2415.390 2290.340 ;
        RECT 379.110 2290.140 379.430 2290.200 ;
        RECT 420.970 2290.140 421.290 2290.200 ;
        RECT 467.890 2290.140 468.210 2290.200 ;
        RECT 513.890 2290.140 514.210 2290.200 ;
        RECT 379.110 2290.000 514.210 2290.140 ;
        RECT 379.110 2289.940 379.430 2290.000 ;
        RECT 420.970 2289.940 421.290 2290.000 ;
        RECT 467.890 2289.940 468.210 2290.000 ;
        RECT 513.890 2289.940 514.210 2290.000 ;
        RECT 531.370 2290.140 531.690 2290.200 ;
        RECT 1104.070 2290.140 1104.390 2290.200 ;
        RECT 531.370 2290.000 1104.390 2290.140 ;
        RECT 531.370 2289.940 531.690 2290.000 ;
        RECT 1104.070 2289.940 1104.390 2290.000 ;
        RECT 1121.550 2290.140 1121.870 2290.200 ;
        RECT 1166.170 2290.140 1166.490 2290.200 ;
        RECT 1121.550 2290.000 1166.490 2290.140 ;
        RECT 1121.550 2289.940 1121.870 2290.000 ;
        RECT 1166.170 2289.940 1166.490 2290.000 ;
        RECT 1717.710 2290.140 1718.030 2290.200 ;
        RECT 1759.110 2290.140 1759.430 2290.200 ;
        RECT 1717.710 2290.000 1759.430 2290.140 ;
        RECT 1717.710 2289.940 1718.030 2290.000 ;
        RECT 1759.110 2289.940 1759.430 2290.000 ;
        RECT 1769.690 2290.140 1770.010 2290.200 ;
        RECT 2415.990 2290.140 2416.310 2290.200 ;
        RECT 1769.690 2290.000 2416.310 2290.140 ;
        RECT 1769.690 2289.940 1770.010 2290.000 ;
        RECT 2415.990 2289.940 2416.310 2290.000 ;
        RECT 434.310 2289.800 434.630 2289.860 ;
        RECT 478.930 2289.800 479.250 2289.860 ;
        RECT 496.870 2289.800 497.190 2289.860 ;
        RECT 434.310 2289.660 497.190 2289.800 ;
        RECT 434.310 2289.600 434.630 2289.660 ;
        RECT 478.930 2289.600 479.250 2289.660 ;
        RECT 496.870 2289.600 497.190 2289.660 ;
        RECT 543.790 2289.800 544.110 2289.860 ;
        RECT 613.710 2289.800 614.030 2289.860 ;
        RECT 543.790 2289.660 614.030 2289.800 ;
        RECT 543.790 2289.600 544.110 2289.660 ;
        RECT 613.710 2289.600 614.030 2289.660 ;
        RECT 635.330 2289.800 635.650 2289.860 ;
        RECT 710.310 2289.800 710.630 2289.860 ;
        RECT 635.330 2289.660 710.630 2289.800 ;
        RECT 635.330 2289.600 635.650 2289.660 ;
        RECT 710.310 2289.600 710.630 2289.660 ;
        RECT 734.690 2289.800 735.010 2289.860 ;
        RECT 806.910 2289.800 807.230 2289.860 ;
        RECT 734.690 2289.660 807.230 2289.800 ;
        RECT 734.690 2289.600 735.010 2289.660 ;
        RECT 806.910 2289.600 807.230 2289.660 ;
        RECT 952.270 2289.800 952.590 2289.860 ;
        RECT 1000.110 2289.800 1000.430 2289.860 ;
        RECT 952.270 2289.660 1000.430 2289.800 ;
        RECT 952.270 2289.600 952.590 2289.660 ;
        RECT 1000.110 2289.600 1000.430 2289.660 ;
        RECT 1124.770 2289.800 1125.090 2289.860 ;
        RECT 1129.370 2289.800 1129.690 2289.860 ;
        RECT 1173.070 2289.800 1173.390 2289.860 ;
        RECT 1124.770 2289.660 1173.390 2289.800 ;
        RECT 1124.770 2289.600 1125.090 2289.660 ;
        RECT 1129.370 2289.600 1129.690 2289.660 ;
        RECT 1173.070 2289.600 1173.390 2289.660 ;
        RECT 1682.750 2289.800 1683.070 2289.860 ;
        RECT 1729.670 2289.800 1729.990 2289.860 ;
        RECT 1768.310 2289.800 1768.630 2289.860 ;
        RECT 1682.750 2289.660 1768.630 2289.800 ;
        RECT 1682.750 2289.600 1683.070 2289.660 ;
        RECT 1729.670 2289.600 1729.990 2289.660 ;
        RECT 1768.310 2289.600 1768.630 2289.660 ;
        RECT 2358.950 2289.800 2359.270 2289.860 ;
        RECT 2402.190 2289.800 2402.510 2289.860 ;
        RECT 2358.950 2289.660 2402.510 2289.800 ;
        RECT 2358.950 2289.600 2359.270 2289.660 ;
        RECT 2402.190 2289.600 2402.510 2289.660 ;
        RECT 406.710 2289.460 407.030 2289.520 ;
        RECT 450.870 2289.460 451.190 2289.520 ;
        RECT 497.330 2289.460 497.650 2289.520 ;
        RECT 543.880 2289.460 544.020 2289.600 ;
        RECT 406.710 2289.320 544.020 2289.460 ;
        RECT 1041.050 2289.460 1041.370 2289.520 ;
        RECT 1083.370 2289.460 1083.690 2289.520 ;
        RECT 1085.670 2289.460 1085.990 2289.520 ;
        RECT 1041.050 2289.320 1085.990 2289.460 ;
        RECT 406.710 2289.260 407.030 2289.320 ;
        RECT 450.870 2289.260 451.190 2289.320 ;
        RECT 497.330 2289.260 497.650 2289.320 ;
        RECT 1041.050 2289.260 1041.370 2289.320 ;
        RECT 1083.370 2289.260 1083.690 2289.320 ;
        RECT 1085.670 2289.260 1085.990 2289.320 ;
        RECT 1086.130 2289.460 1086.450 2289.520 ;
        RECT 1121.550 2289.460 1121.870 2289.520 ;
        RECT 1086.130 2289.320 1121.870 2289.460 ;
        RECT 1086.130 2289.260 1086.450 2289.320 ;
        RECT 1121.550 2289.260 1121.870 2289.320 ;
        RECT 1656.530 2289.460 1656.850 2289.520 ;
        RECT 1659.290 2289.460 1659.610 2289.520 ;
        RECT 1706.210 2289.460 1706.530 2289.520 ;
        RECT 1752.670 2289.460 1752.990 2289.520 ;
        RECT 1656.530 2289.320 1752.990 2289.460 ;
        RECT 1656.530 2289.260 1656.850 2289.320 ;
        RECT 1659.290 2289.260 1659.610 2289.320 ;
        RECT 1706.210 2289.260 1706.530 2289.320 ;
        RECT 1752.670 2289.260 1752.990 2289.320 ;
        RECT 1753.130 2289.460 1753.450 2289.520 ;
        RECT 1780.270 2289.460 1780.590 2289.520 ;
        RECT 1753.130 2289.320 1780.590 2289.460 ;
        RECT 1753.130 2289.260 1753.450 2289.320 ;
        RECT 1780.270 2289.260 1780.590 2289.320 ;
        RECT 2300.990 2289.460 2301.310 2289.520 ;
        RECT 2343.770 2289.460 2344.090 2289.520 ;
        RECT 2391.610 2289.460 2391.930 2289.520 ;
        RECT 2435.770 2289.460 2436.090 2289.520 ;
        RECT 2300.990 2289.320 2436.090 2289.460 ;
        RECT 2300.990 2289.260 2301.310 2289.320 ;
        RECT 2343.770 2289.260 2344.090 2289.320 ;
        RECT 2391.610 2289.260 2391.930 2289.320 ;
        RECT 2435.770 2289.260 2436.090 2289.320 ;
        RECT 392.910 2289.120 393.230 2289.180 ;
        RECT 439.370 2289.120 439.690 2289.180 ;
        RECT 485.830 2289.120 486.150 2289.180 ;
        RECT 489.510 2289.120 489.830 2289.180 ;
        RECT 392.910 2288.980 489.830 2289.120 ;
        RECT 392.910 2288.920 393.230 2288.980 ;
        RECT 439.370 2288.920 439.690 2288.980 ;
        RECT 485.830 2288.920 486.150 2288.980 ;
        RECT 489.510 2288.920 489.830 2288.980 ;
        RECT 1065.430 2289.120 1065.750 2289.180 ;
        RECT 1112.810 2289.120 1113.130 2289.180 ;
        RECT 1159.270 2289.120 1159.590 2289.180 ;
        RECT 1065.430 2288.980 1159.590 2289.120 ;
        RECT 1065.430 2288.920 1065.750 2288.980 ;
        RECT 1112.810 2288.920 1113.130 2288.980 ;
        RECT 1159.270 2288.920 1159.590 2288.980 ;
        RECT 1695.170 2289.120 1695.490 2289.180 ;
        RECT 1704.370 2289.120 1704.690 2289.180 ;
        RECT 1695.170 2288.980 1704.690 2289.120 ;
        RECT 1695.170 2288.920 1695.490 2288.980 ;
        RECT 1704.370 2288.920 1704.690 2288.980 ;
        RECT 2324.910 2289.120 2325.230 2289.180 ;
        RECT 2357.570 2289.120 2357.890 2289.180 ;
        RECT 2377.350 2289.120 2377.670 2289.180 ;
        RECT 2421.970 2289.120 2422.290 2289.180 ;
        RECT 2324.910 2288.980 2357.340 2289.120 ;
        RECT 2324.910 2288.920 2325.230 2288.980 ;
        RECT 445.350 2288.780 445.670 2288.840 ;
        RECT 492.730 2288.780 493.050 2288.840 ;
        RECT 538.270 2288.780 538.590 2288.840 ;
        RECT 445.350 2288.640 538.590 2288.780 ;
        RECT 445.350 2288.580 445.670 2288.640 ;
        RECT 492.730 2288.580 493.050 2288.640 ;
        RECT 538.270 2288.580 538.590 2288.640 ;
        RECT 1070.030 2288.780 1070.350 2288.840 ;
        RECT 1118.330 2288.780 1118.650 2288.840 ;
        RECT 1070.030 2288.640 1118.650 2288.780 ;
        RECT 1070.030 2288.580 1070.350 2288.640 ;
        RECT 1118.330 2288.580 1118.650 2288.640 ;
        RECT 1132.130 2288.780 1132.450 2288.840 ;
        RECT 1135.810 2288.780 1136.130 2288.840 ;
        RECT 1179.970 2288.780 1180.290 2288.840 ;
        RECT 1132.130 2288.640 1180.290 2288.780 ;
        RECT 1132.130 2288.580 1132.450 2288.640 ;
        RECT 1135.810 2288.580 1136.130 2288.640 ;
        RECT 1179.970 2288.580 1180.290 2288.640 ;
        RECT 1662.970 2288.780 1663.290 2288.840 ;
        RECT 1665.730 2288.780 1666.050 2288.840 ;
        RECT 1712.650 2288.780 1712.970 2288.840 ;
        RECT 1717.710 2288.780 1718.030 2288.840 ;
        RECT 1662.970 2288.640 1718.030 2288.780 ;
        RECT 1662.970 2288.580 1663.290 2288.640 ;
        RECT 1665.730 2288.580 1666.050 2288.640 ;
        RECT 1712.650 2288.580 1712.970 2288.640 ;
        RECT 1717.710 2288.580 1718.030 2288.640 ;
        RECT 1746.230 2288.780 1746.550 2288.840 ;
        RECT 1748.530 2288.780 1748.850 2288.840 ;
        RECT 2267.410 2288.780 2267.730 2288.840 ;
        RECT 2315.250 2288.780 2315.570 2288.840 ;
        RECT 2356.650 2288.780 2356.970 2288.840 ;
        RECT 1746.230 2288.640 1748.300 2288.780 ;
        RECT 1746.230 2288.580 1746.550 2288.640 ;
        RECT 365.310 2288.440 365.630 2288.500 ;
        RECT 409.470 2288.440 409.790 2288.500 ;
        RECT 455.470 2288.440 455.790 2288.500 ;
        RECT 365.310 2288.300 455.790 2288.440 ;
        RECT 365.310 2288.240 365.630 2288.300 ;
        RECT 409.470 2288.240 409.790 2288.300 ;
        RECT 455.470 2288.240 455.790 2288.300 ;
        RECT 489.510 2288.440 489.830 2288.500 ;
        RECT 531.370 2288.440 531.690 2288.500 ;
        RECT 489.510 2288.300 531.690 2288.440 ;
        RECT 489.510 2288.240 489.830 2288.300 ;
        RECT 531.370 2288.240 531.690 2288.300 ;
        RECT 882.810 2288.440 883.130 2288.500 ;
        RECT 1007.470 2288.440 1007.790 2288.500 ;
        RECT 882.810 2288.300 1007.790 2288.440 ;
        RECT 882.810 2288.240 883.130 2288.300 ;
        RECT 1007.470 2288.240 1007.790 2288.300 ;
        RECT 1038.750 2288.440 1039.070 2288.500 ;
        RECT 1048.410 2288.440 1048.730 2288.500 ;
        RECT 1094.410 2288.440 1094.730 2288.500 ;
        RECT 1141.790 2288.440 1142.110 2288.500 ;
        RECT 1186.870 2288.440 1187.190 2288.500 ;
        RECT 1038.750 2288.300 1187.190 2288.440 ;
        RECT 1038.750 2288.240 1039.070 2288.300 ;
        RECT 1048.410 2288.240 1048.730 2288.300 ;
        RECT 1094.410 2288.240 1094.730 2288.300 ;
        RECT 1141.790 2288.240 1142.110 2288.300 ;
        RECT 1186.870 2288.240 1187.190 2288.300 ;
        RECT 1690.110 2288.440 1690.430 2288.500 ;
        RECT 1734.270 2288.440 1734.590 2288.500 ;
        RECT 1748.160 2288.440 1748.300 2288.640 ;
        RECT 1748.530 2288.640 1768.080 2288.780 ;
        RECT 1748.530 2288.580 1748.850 2288.640 ;
        RECT 1767.940 2288.440 1768.080 2288.640 ;
        RECT 2267.410 2288.640 2356.970 2288.780 ;
        RECT 2357.200 2288.780 2357.340 2288.980 ;
        RECT 2357.570 2288.980 2422.290 2289.120 ;
        RECT 2357.570 2288.920 2357.890 2288.980 ;
        RECT 2377.350 2288.920 2377.670 2288.980 ;
        RECT 2421.970 2288.920 2422.290 2288.980 ;
        RECT 2367.230 2288.780 2367.550 2288.840 ;
        RECT 2401.270 2288.780 2401.590 2288.840 ;
        RECT 2357.200 2288.640 2401.590 2288.780 ;
        RECT 2267.410 2288.580 2267.730 2288.640 ;
        RECT 2315.250 2288.580 2315.570 2288.640 ;
        RECT 2356.650 2288.580 2356.970 2288.640 ;
        RECT 2367.230 2288.580 2367.550 2288.640 ;
        RECT 2401.270 2288.580 2401.590 2288.640 ;
        RECT 1787.170 2288.440 1787.490 2288.500 ;
        RECT 1690.110 2288.300 1746.920 2288.440 ;
        RECT 1748.160 2288.300 1767.620 2288.440 ;
        RECT 1767.940 2288.300 1787.490 2288.440 ;
        RECT 1690.110 2288.240 1690.430 2288.300 ;
        RECT 1734.270 2288.240 1734.590 2288.300 ;
        RECT 370.830 2288.100 371.150 2288.160 ;
        RECT 414.070 2288.100 414.390 2288.160 ;
        RECT 462.370 2288.100 462.690 2288.160 ;
        RECT 509.290 2288.100 509.610 2288.160 ;
        RECT 370.830 2287.960 509.610 2288.100 ;
        RECT 370.830 2287.900 371.150 2287.960 ;
        RECT 414.070 2287.900 414.390 2287.960 ;
        RECT 462.370 2287.900 462.690 2287.960 ;
        RECT 509.290 2287.900 509.610 2287.960 ;
        RECT 875.910 2288.100 876.230 2288.160 ;
        RECT 1001.030 2288.100 1001.350 2288.160 ;
        RECT 875.910 2287.960 1001.350 2288.100 ;
        RECT 875.910 2287.900 876.230 2287.960 ;
        RECT 1001.030 2287.900 1001.350 2287.960 ;
        RECT 1045.650 2288.100 1045.970 2288.160 ;
        RECT 1052.550 2288.100 1052.870 2288.160 ;
        RECT 1100.850 2288.100 1101.170 2288.160 ;
        RECT 1147.770 2288.100 1148.090 2288.160 ;
        RECT 1193.770 2288.100 1194.090 2288.160 ;
        RECT 1045.650 2287.960 1194.090 2288.100 ;
        RECT 1045.650 2287.900 1045.970 2287.960 ;
        RECT 1052.550 2287.900 1052.870 2287.960 ;
        RECT 1100.850 2287.900 1101.170 2287.960 ;
        RECT 1147.770 2287.900 1148.090 2287.960 ;
        RECT 1193.770 2287.900 1194.090 2287.960 ;
        RECT 1699.310 2288.100 1699.630 2288.160 ;
        RECT 1746.230 2288.100 1746.550 2288.160 ;
        RECT 1699.310 2287.960 1746.550 2288.100 ;
        RECT 1746.780 2288.100 1746.920 2288.300 ;
        RECT 1753.130 2288.100 1753.450 2288.160 ;
        RECT 1746.780 2287.960 1753.450 2288.100 ;
        RECT 1767.480 2288.100 1767.620 2288.300 ;
        RECT 1787.170 2288.240 1787.490 2288.300 ;
        RECT 1797.290 2288.440 1797.610 2288.500 ;
        RECT 2290.870 2288.440 2291.190 2288.500 ;
        RECT 1797.290 2288.300 2291.190 2288.440 ;
        RECT 1797.290 2288.240 1797.610 2288.300 ;
        RECT 2290.870 2288.240 2291.190 2288.300 ;
        RECT 2301.910 2288.440 2302.230 2288.500 ;
        RECT 2349.750 2288.440 2350.070 2288.500 ;
        RECT 2397.130 2288.440 2397.450 2288.500 ;
        RECT 2442.670 2288.440 2442.990 2288.500 ;
        RECT 2301.910 2288.300 2442.990 2288.440 ;
        RECT 2301.910 2288.240 2302.230 2288.300 ;
        RECT 2349.750 2288.240 2350.070 2288.300 ;
        RECT 2397.130 2288.240 2397.450 2288.300 ;
        RECT 2442.670 2288.240 2442.990 2288.300 ;
        RECT 1794.070 2288.100 1794.390 2288.160 ;
        RECT 1767.480 2287.960 1794.390 2288.100 ;
        RECT 1699.310 2287.900 1699.630 2287.960 ;
        RECT 1746.230 2287.900 1746.550 2287.960 ;
        RECT 1753.130 2287.900 1753.450 2287.960 ;
        RECT 1794.070 2287.900 1794.390 2287.960 ;
        RECT 2266.490 2288.100 2266.810 2288.160 ;
        RECT 2308.810 2288.100 2309.130 2288.160 ;
        RECT 2358.950 2288.100 2359.270 2288.160 ;
        RECT 2361.250 2288.100 2361.570 2288.160 ;
        RECT 2408.170 2288.100 2408.490 2288.160 ;
        RECT 2266.490 2287.960 2359.270 2288.100 ;
        RECT 2266.490 2287.900 2266.810 2287.960 ;
        RECT 2308.810 2287.900 2309.130 2287.960 ;
        RECT 2358.950 2287.900 2359.270 2287.960 ;
        RECT 2359.500 2287.960 2408.490 2288.100 ;
        RECT 386.010 2287.760 386.330 2287.820 ;
        RECT 427.410 2287.760 427.730 2287.820 ;
        RECT 473.870 2287.760 474.190 2287.820 ;
        RECT 521.250 2287.760 521.570 2287.820 ;
        RECT 386.010 2287.620 521.570 2287.760 ;
        RECT 386.010 2287.560 386.330 2287.620 ;
        RECT 427.410 2287.560 427.730 2287.620 ;
        RECT 473.870 2287.560 474.190 2287.620 ;
        RECT 521.250 2287.560 521.570 2287.620 ;
        RECT 862.110 2287.760 862.430 2287.820 ;
        RECT 993.670 2287.760 993.990 2287.820 ;
        RECT 862.110 2287.620 993.990 2287.760 ;
        RECT 862.110 2287.560 862.430 2287.620 ;
        RECT 993.670 2287.560 993.990 2287.620 ;
        RECT 1062.210 2287.760 1062.530 2287.820 ;
        RECT 1106.830 2287.760 1107.150 2287.820 ;
        RECT 1152.370 2287.760 1152.690 2287.820 ;
        RECT 1062.210 2287.620 1152.690 2287.760 ;
        RECT 1062.210 2287.560 1062.530 2287.620 ;
        RECT 1106.830 2287.560 1107.150 2287.620 ;
        RECT 1152.370 2287.560 1152.690 2287.620 ;
        RECT 1670.330 2287.760 1670.650 2287.820 ;
        RECT 1721.850 2287.760 1722.170 2287.820 ;
        RECT 1670.330 2287.620 1722.170 2287.760 ;
        RECT 1670.330 2287.560 1670.650 2287.620 ;
        RECT 1721.850 2287.560 1722.170 2287.620 ;
        RECT 1768.310 2287.760 1768.630 2287.820 ;
        RECT 1775.210 2287.760 1775.530 2287.820 ;
        RECT 1768.310 2287.620 1775.530 2287.760 ;
        RECT 1768.310 2287.560 1768.630 2287.620 ;
        RECT 1775.210 2287.560 1775.530 2287.620 ;
        RECT 1790.390 2287.760 1790.710 2287.820 ;
        RECT 2283.970 2287.760 2284.290 2287.820 ;
        RECT 1790.390 2287.620 2284.290 2287.760 ;
        RECT 1790.390 2287.560 1790.710 2287.620 ;
        RECT 2283.970 2287.560 2284.290 2287.620 ;
        RECT 2325.830 2287.760 2326.150 2287.820 ;
        RECT 2356.190 2287.760 2356.510 2287.820 ;
        RECT 2325.830 2287.620 2356.510 2287.760 ;
        RECT 2325.830 2287.560 2326.150 2287.620 ;
        RECT 2356.190 2287.560 2356.510 2287.620 ;
        RECT 2356.650 2287.760 2356.970 2287.820 ;
        RECT 2359.500 2287.760 2359.640 2287.960 ;
        RECT 2361.250 2287.900 2361.570 2287.960 ;
        RECT 2408.170 2287.900 2408.490 2287.960 ;
        RECT 2356.650 2287.620 2359.640 2287.760 ;
        RECT 2381.490 2287.760 2381.810 2287.820 ;
        RECT 2384.710 2287.760 2385.030 2287.820 ;
        RECT 2428.870 2287.760 2429.190 2287.820 ;
        RECT 2381.490 2287.620 2429.190 2287.760 ;
        RECT 2356.650 2287.560 2356.970 2287.620 ;
        RECT 2381.490 2287.560 2381.810 2287.620 ;
        RECT 2384.710 2287.560 2385.030 2287.620 ;
        RECT 2428.870 2287.560 2429.190 2287.620 ;
        RECT 2218.190 2287.420 2218.510 2287.480 ;
        RECT 2297.770 2287.420 2298.090 2287.480 ;
        RECT 2218.190 2287.280 2298.090 2287.420 ;
        RECT 2218.190 2287.220 2218.510 2287.280 ;
        RECT 2297.770 2287.220 2298.090 2287.280 ;
        RECT 2328.590 2287.420 2328.910 2287.480 ;
        RECT 2435.770 2287.420 2436.090 2287.480 ;
        RECT 2328.590 2287.280 2436.090 2287.420 ;
        RECT 2328.590 2287.220 2328.910 2287.280 ;
        RECT 2435.770 2287.220 2436.090 2287.280 ;
        RECT 855.210 2287.080 855.530 2287.140 ;
        RECT 986.770 2287.080 987.090 2287.140 ;
        RECT 855.210 2286.940 987.090 2287.080 ;
        RECT 855.210 2286.880 855.530 2286.940 ;
        RECT 986.770 2286.880 987.090 2286.940 ;
        RECT 1045.190 2287.080 1045.510 2287.140 ;
        RECT 1085.670 2287.080 1085.990 2287.140 ;
        RECT 1124.770 2287.080 1125.090 2287.140 ;
        RECT 1045.190 2286.940 1078.540 2287.080 ;
        RECT 1045.190 2286.880 1045.510 2286.940 ;
        RECT 668.910 2286.740 669.230 2286.800 ;
        RECT 979.870 2286.740 980.190 2286.800 ;
        RECT 668.910 2286.600 980.190 2286.740 ;
        RECT 668.910 2286.540 669.230 2286.600 ;
        RECT 979.870 2286.540 980.190 2286.600 ;
        RECT 1010.690 2286.740 1011.010 2286.800 ;
        RECT 1062.210 2286.740 1062.530 2286.800 ;
        RECT 1010.690 2286.600 1062.530 2286.740 ;
        RECT 1078.400 2286.740 1078.540 2286.940 ;
        RECT 1085.670 2286.940 1125.090 2287.080 ;
        RECT 1085.670 2286.880 1085.990 2286.940 ;
        RECT 1124.770 2286.880 1125.090 2286.940 ;
        RECT 1548.890 2287.080 1549.210 2287.140 ;
        RECT 1656.070 2287.080 1656.390 2287.140 ;
        RECT 1548.890 2286.940 1656.390 2287.080 ;
        RECT 1548.890 2286.880 1549.210 2286.940 ;
        RECT 1656.070 2286.880 1656.390 2286.940 ;
        RECT 1704.370 2287.080 1704.690 2287.140 ;
        RECT 1741.170 2287.080 1741.490 2287.140 ;
        RECT 1748.530 2287.080 1748.850 2287.140 ;
        RECT 1704.370 2286.940 1748.850 2287.080 ;
        RECT 1704.370 2286.880 1704.690 2286.940 ;
        RECT 1741.170 2286.880 1741.490 2286.940 ;
        RECT 1748.530 2286.880 1748.850 2286.940 ;
        RECT 1776.590 2287.080 1776.910 2287.140 ;
        RECT 2270.170 2287.080 2270.490 2287.140 ;
        RECT 1776.590 2286.940 2270.490 2287.080 ;
        RECT 1776.590 2286.880 1776.910 2286.940 ;
        RECT 2270.170 2286.880 2270.490 2286.940 ;
        RECT 2273.390 2287.080 2273.710 2287.140 ;
        RECT 2324.910 2287.080 2325.230 2287.140 ;
        RECT 2273.390 2286.940 2325.230 2287.080 ;
        RECT 2273.390 2286.880 2273.710 2286.940 ;
        RECT 2324.910 2286.880 2325.230 2286.940 ;
        RECT 2335.490 2287.080 2335.810 2287.140 ;
        RECT 2442.670 2287.080 2442.990 2287.140 ;
        RECT 2335.490 2286.940 2442.990 2287.080 ;
        RECT 2335.490 2286.880 2335.810 2286.940 ;
        RECT 2442.670 2286.880 2442.990 2286.940 ;
        RECT 1087.970 2286.740 1088.290 2286.800 ;
        RECT 1132.130 2286.740 1132.450 2286.800 ;
        RECT 1078.400 2286.600 1132.450 2286.740 ;
        RECT 1010.690 2286.540 1011.010 2286.600 ;
        RECT 1062.210 2286.540 1062.530 2286.600 ;
        RECT 1087.970 2286.540 1088.290 2286.600 ;
        RECT 1132.130 2286.540 1132.450 2286.600 ;
        RECT 1610.990 2286.740 1611.310 2286.800 ;
        RECT 1656.530 2286.740 1656.850 2286.800 ;
        RECT 1610.990 2286.600 1656.850 2286.740 ;
        RECT 1610.990 2286.540 1611.310 2286.600 ;
        RECT 1656.530 2286.540 1656.850 2286.600 ;
        RECT 1714.490 2286.740 1714.810 2286.800 ;
        RECT 2263.270 2286.740 2263.590 2286.800 ;
        RECT 1714.490 2286.600 2263.590 2286.740 ;
        RECT 1714.490 2286.540 1714.810 2286.600 ;
        RECT 2263.270 2286.540 2263.590 2286.600 ;
        RECT 2321.690 2286.740 2322.010 2286.800 ;
        RECT 2428.870 2286.740 2429.190 2286.800 ;
        RECT 2321.690 2286.600 2429.190 2286.740 ;
        RECT 2321.690 2286.540 2322.010 2286.600 ;
        RECT 2428.870 2286.540 2429.190 2286.600 ;
        RECT 502.850 2286.400 503.170 2286.460 ;
        RECT 1048.870 2286.400 1049.190 2286.460 ;
        RECT 502.850 2286.260 1049.190 2286.400 ;
        RECT 502.850 2286.200 503.170 2286.260 ;
        RECT 1048.870 2286.200 1049.190 2286.260 ;
        RECT 1049.330 2286.400 1049.650 2286.460 ;
        RECT 1096.710 2286.400 1097.030 2286.460 ;
        RECT 1049.330 2286.260 1097.030 2286.400 ;
        RECT 1049.330 2286.200 1049.650 2286.260 ;
        RECT 1096.710 2286.200 1097.030 2286.260 ;
        RECT 1562.690 2286.400 1563.010 2286.460 ;
        RECT 1649.170 2286.400 1649.490 2286.460 ;
        RECT 1562.690 2286.260 1649.490 2286.400 ;
        RECT 1562.690 2286.200 1563.010 2286.260 ;
        RECT 1649.170 2286.200 1649.490 2286.260 ;
        RECT 1748.990 2286.400 1749.310 2286.460 ;
        RECT 2387.470 2286.400 2387.790 2286.460 ;
        RECT 1748.990 2286.260 2387.790 2286.400 ;
        RECT 1748.990 2286.200 1749.310 2286.260 ;
        RECT 2387.470 2286.200 2387.790 2286.260 ;
        RECT 2401.270 2286.400 2401.590 2286.460 ;
        RECT 2415.530 2286.400 2415.850 2286.460 ;
        RECT 2401.270 2286.260 2415.850 2286.400 ;
        RECT 2401.270 2286.200 2401.590 2286.260 ;
        RECT 2415.530 2286.200 2415.850 2286.260 ;
        RECT 509.290 2286.060 509.610 2286.120 ;
        RECT 1062.670 2286.060 1062.990 2286.120 ;
        RECT 509.290 2285.920 1062.990 2286.060 ;
        RECT 509.290 2285.860 509.610 2285.920 ;
        RECT 1062.670 2285.860 1062.990 2285.920 ;
        RECT 1639.510 2286.060 1639.830 2286.120 ;
        RECT 1682.750 2286.060 1683.070 2286.120 ;
        RECT 1639.510 2285.920 1683.070 2286.060 ;
        RECT 1639.510 2285.860 1639.830 2285.920 ;
        RECT 1682.750 2285.860 1683.070 2285.920 ;
        RECT 1755.890 2286.060 1756.210 2286.120 ;
        RECT 2394.370 2286.060 2394.690 2286.120 ;
        RECT 1755.890 2285.920 2394.690 2286.060 ;
        RECT 1755.890 2285.860 1756.210 2285.920 ;
        RECT 2394.370 2285.860 2394.690 2285.920 ;
        RECT 317.010 2285.720 317.330 2285.780 ;
        RECT 365.770 2285.720 366.090 2285.780 ;
        RECT 317.010 2285.580 366.090 2285.720 ;
        RECT 317.010 2285.520 317.330 2285.580 ;
        RECT 365.770 2285.520 366.090 2285.580 ;
        RECT 513.890 2285.720 514.210 2285.780 ;
        RECT 1069.570 2285.720 1069.890 2285.780 ;
        RECT 513.890 2285.580 1069.890 2285.720 ;
        RECT 513.890 2285.520 514.210 2285.580 ;
        RECT 1069.570 2285.520 1069.890 2285.580 ;
        RECT 1076.010 2285.720 1076.330 2285.780 ;
        RECT 1231.490 2285.720 1231.810 2285.780 ;
        RECT 1076.010 2285.580 1231.810 2285.720 ;
        RECT 1076.010 2285.520 1076.330 2285.580 ;
        RECT 1231.490 2285.520 1231.810 2285.580 ;
        RECT 1576.490 2285.720 1576.810 2285.780 ;
        RECT 1642.270 2285.720 1642.590 2285.780 ;
        RECT 1576.490 2285.580 1642.590 2285.720 ;
        RECT 1576.490 2285.520 1576.810 2285.580 ;
        RECT 1642.270 2285.520 1642.590 2285.580 ;
        RECT 1646.410 2285.720 1646.730 2285.780 ;
        RECT 1695.170 2285.720 1695.490 2285.780 ;
        RECT 1646.410 2285.580 1695.490 2285.720 ;
        RECT 1646.410 2285.520 1646.730 2285.580 ;
        RECT 1695.170 2285.520 1695.490 2285.580 ;
        RECT 1762.790 2285.720 1763.110 2285.780 ;
        RECT 2402.650 2285.720 2402.970 2285.780 ;
        RECT 1762.790 2285.580 2402.970 2285.720 ;
        RECT 1762.790 2285.520 1763.110 2285.580 ;
        RECT 2402.650 2285.520 2402.970 2285.580 ;
        RECT 351.510 2285.380 351.830 2285.440 ;
        RECT 386.470 2285.380 386.790 2285.440 ;
        RECT 351.510 2285.240 386.790 2285.380 ;
        RECT 351.510 2285.180 351.830 2285.240 ;
        RECT 386.470 2285.180 386.790 2285.240 ;
        RECT 521.250 2285.380 521.570 2285.440 ;
        RECT 1083.370 2285.380 1083.690 2285.440 ;
        RECT 521.250 2285.240 1083.690 2285.380 ;
        RECT 521.250 2285.180 521.570 2285.240 ;
        RECT 1083.370 2285.180 1083.690 2285.240 ;
        RECT 1617.890 2285.380 1618.210 2285.440 ;
        RECT 1662.970 2285.380 1663.290 2285.440 ;
        RECT 1617.890 2285.240 1663.290 2285.380 ;
        RECT 1617.890 2285.180 1618.210 2285.240 ;
        RECT 1662.970 2285.180 1663.290 2285.240 ;
        RECT 1763.250 2285.380 1763.570 2285.440 ;
        RECT 2408.170 2285.380 2408.490 2285.440 ;
        RECT 1763.250 2285.240 2408.490 2285.380 ;
        RECT 1763.250 2285.180 1763.570 2285.240 ;
        RECT 2408.170 2285.180 2408.490 2285.240 ;
        RECT 344.610 2285.040 344.930 2285.100 ;
        RECT 379.570 2285.040 379.890 2285.100 ;
        RECT 344.610 2284.900 379.890 2285.040 ;
        RECT 344.610 2284.840 344.930 2284.900 ;
        RECT 379.570 2284.840 379.890 2284.900 ;
        RECT 526.770 2285.040 527.090 2285.100 ;
        RECT 1097.170 2285.040 1097.490 2285.100 ;
        RECT 526.770 2284.900 1097.490 2285.040 ;
        RECT 526.770 2284.840 527.090 2284.900 ;
        RECT 1097.170 2284.840 1097.490 2284.900 ;
        RECT 1541.990 2285.040 1542.310 2285.100 ;
        RECT 1587.070 2285.040 1587.390 2285.100 ;
        RECT 1541.990 2284.900 1587.390 2285.040 ;
        RECT 1541.990 2284.840 1542.310 2284.900 ;
        RECT 1587.070 2284.840 1587.390 2284.900 ;
        RECT 1735.190 2285.040 1735.510 2285.100 ;
        RECT 2380.570 2285.040 2380.890 2285.100 ;
        RECT 1735.190 2284.900 2380.890 2285.040 ;
        RECT 1735.190 2284.840 1735.510 2284.900 ;
        RECT 2380.570 2284.840 2380.890 2284.900 ;
        RECT 330.810 2284.700 331.130 2284.760 ;
        RECT 373.590 2284.700 373.910 2284.760 ;
        RECT 330.810 2284.560 373.910 2284.700 ;
        RECT 330.810 2284.500 331.130 2284.560 ;
        RECT 373.590 2284.500 373.910 2284.560 ;
        RECT 1034.150 2284.700 1034.470 2284.760 ;
        RECT 1076.470 2284.700 1076.790 2284.760 ;
        RECT 1034.150 2284.560 1076.790 2284.700 ;
        RECT 1034.150 2284.500 1034.470 2284.560 ;
        RECT 1076.470 2284.500 1076.790 2284.560 ;
        RECT 1624.790 2284.700 1625.110 2284.760 ;
        RECT 1670.330 2284.700 1670.650 2284.760 ;
        RECT 1624.790 2284.560 1670.650 2284.700 ;
        RECT 1624.790 2284.500 1625.110 2284.560 ;
        RECT 1670.330 2284.500 1670.650 2284.560 ;
        RECT 2296.850 2284.700 2297.170 2284.760 ;
        RECT 2340.090 2284.700 2340.410 2284.760 ;
        RECT 2381.490 2284.700 2381.810 2284.760 ;
        RECT 2296.850 2284.560 2381.810 2284.700 ;
        RECT 2296.850 2284.500 2297.170 2284.560 ;
        RECT 2340.090 2284.500 2340.410 2284.560 ;
        RECT 2381.490 2284.500 2381.810 2284.560 ;
        RECT 365.310 2284.360 365.630 2284.420 ;
        RECT 393.830 2284.360 394.150 2284.420 ;
        RECT 365.310 2284.220 394.150 2284.360 ;
        RECT 365.310 2284.160 365.630 2284.220 ;
        RECT 393.830 2284.160 394.150 2284.220 ;
        RECT 1027.250 2284.360 1027.570 2284.420 ;
        RECT 1070.030 2284.360 1070.350 2284.420 ;
        RECT 1027.250 2284.220 1070.350 2284.360 ;
        RECT 1027.250 2284.160 1027.570 2284.220 ;
        RECT 1070.030 2284.160 1070.350 2284.220 ;
        RECT 1082.910 2284.360 1083.230 2284.420 ;
        RECT 1224.590 2284.360 1224.910 2284.420 ;
        RECT 1082.910 2284.220 1224.910 2284.360 ;
        RECT 1082.910 2284.160 1083.230 2284.220 ;
        RECT 1224.590 2284.160 1224.910 2284.220 ;
        RECT 1631.690 2284.360 1632.010 2284.420 ;
        RECT 1677.230 2284.360 1677.550 2284.420 ;
        RECT 1631.690 2284.220 1677.550 2284.360 ;
        RECT 1631.690 2284.160 1632.010 2284.220 ;
        RECT 1677.230 2284.160 1677.550 2284.220 ;
        RECT 1783.490 2284.360 1783.810 2284.420 ;
        RECT 2277.070 2284.360 2277.390 2284.420 ;
        RECT 1783.490 2284.220 2277.390 2284.360 ;
        RECT 1783.490 2284.160 1783.810 2284.220 ;
        RECT 2277.070 2284.160 2277.390 2284.220 ;
        RECT 2283.510 2284.360 2283.830 2284.420 ;
        RECT 2325.830 2284.360 2326.150 2284.420 ;
        RECT 2333.190 2284.360 2333.510 2284.420 ;
        RECT 2355.730 2284.360 2356.050 2284.420 ;
        RECT 2283.510 2284.220 2326.150 2284.360 ;
        RECT 2283.510 2284.160 2283.830 2284.220 ;
        RECT 2325.830 2284.160 2326.150 2284.220 ;
        RECT 2330.060 2284.220 2356.050 2284.360 ;
        RECT 310.110 2284.020 310.430 2284.080 ;
        RECT 358.870 2284.020 359.190 2284.080 ;
        RECT 310.110 2283.880 359.190 2284.020 ;
        RECT 310.110 2283.820 310.430 2283.880 ;
        RECT 358.870 2283.820 359.190 2283.880 ;
        RECT 382.790 2284.020 383.110 2284.080 ;
        RECT 393.370 2284.020 393.690 2284.080 ;
        RECT 382.790 2283.880 393.690 2284.020 ;
        RECT 382.790 2283.820 383.110 2283.880 ;
        RECT 393.370 2283.820 393.690 2283.880 ;
        RECT 1017.590 2284.020 1017.910 2284.080 ;
        RECT 1065.430 2284.020 1065.750 2284.080 ;
        RECT 1017.590 2283.880 1065.750 2284.020 ;
        RECT 1017.590 2283.820 1017.910 2283.880 ;
        RECT 1065.430 2283.820 1065.750 2283.880 ;
        RECT 1089.810 2284.020 1090.130 2284.080 ;
        RECT 1210.790 2284.020 1211.110 2284.080 ;
        RECT 1089.810 2283.880 1211.110 2284.020 ;
        RECT 1089.810 2283.820 1090.130 2283.880 ;
        RECT 1210.790 2283.820 1211.110 2283.880 ;
        RECT 1583.390 2284.020 1583.710 2284.080 ;
        RECT 1621.570 2284.020 1621.890 2284.080 ;
        RECT 1583.390 2283.880 1621.890 2284.020 ;
        RECT 1583.390 2283.820 1583.710 2283.880 ;
        RECT 1621.570 2283.820 1621.890 2283.880 ;
        RECT 1652.390 2284.020 1652.710 2284.080 ;
        RECT 1699.310 2284.020 1699.630 2284.080 ;
        RECT 1652.390 2283.880 1699.630 2284.020 ;
        RECT 1652.390 2283.820 1652.710 2283.880 ;
        RECT 1699.310 2283.820 1699.630 2283.880 ;
        RECT 2290.410 2284.020 2290.730 2284.080 ;
        RECT 2330.060 2284.020 2330.200 2284.220 ;
        RECT 2333.190 2284.160 2333.510 2284.220 ;
        RECT 2355.730 2284.160 2356.050 2284.220 ;
        RECT 2356.190 2284.360 2356.510 2284.420 ;
        RECT 2374.130 2284.360 2374.450 2284.420 ;
        RECT 2415.070 2284.360 2415.390 2284.420 ;
        RECT 2356.190 2284.220 2415.390 2284.360 ;
        RECT 2356.190 2284.160 2356.510 2284.220 ;
        RECT 2374.130 2284.160 2374.450 2284.220 ;
        RECT 2415.070 2284.160 2415.390 2284.220 ;
        RECT 2290.410 2283.880 2330.200 2284.020 ;
        RECT 2290.410 2283.820 2290.730 2283.880 ;
        RECT 1638.130 2222.140 1638.450 2222.200 ;
        RECT 1638.590 2222.140 1638.910 2222.200 ;
        RECT 1638.130 2222.000 1638.910 2222.140 ;
        RECT 1638.130 2221.940 1638.450 2222.000 ;
        RECT 1638.590 2221.940 1638.910 2222.000 ;
        RECT 1211.710 2216.360 1212.030 2216.420 ;
        RECT 1225.510 2216.360 1225.830 2216.420 ;
        RECT 1211.710 2216.220 1225.830 2216.360 ;
        RECT 1211.710 2216.160 1212.030 2216.220 ;
        RECT 1225.510 2216.160 1225.830 2216.220 ;
        RECT 305.510 2214.660 305.830 2214.720 ;
        RECT 310.110 2214.660 310.430 2214.720 ;
        RECT 305.510 2214.520 310.430 2214.660 ;
        RECT 305.510 2214.460 305.830 2214.520 ;
        RECT 310.110 2214.460 310.430 2214.520 ;
        RECT 339.090 2214.660 339.410 2214.720 ;
        RECT 344.610 2214.660 344.930 2214.720 ;
        RECT 339.090 2214.520 344.930 2214.660 ;
        RECT 339.090 2214.460 339.410 2214.520 ;
        RECT 344.610 2214.460 344.930 2214.520 ;
        RECT 373.130 2214.660 373.450 2214.720 ;
        RECT 382.790 2214.660 383.110 2214.720 ;
        RECT 373.130 2214.520 383.110 2214.660 ;
        RECT 373.130 2214.460 373.450 2214.520 ;
        RECT 382.790 2214.460 383.110 2214.520 ;
        RECT 384.630 2214.660 384.950 2214.720 ;
        RECT 400.270 2214.660 400.590 2214.720 ;
        RECT 384.630 2214.520 400.590 2214.660 ;
        RECT 384.630 2214.460 384.950 2214.520 ;
        RECT 400.270 2214.460 400.590 2214.520 ;
        RECT 407.170 2214.660 407.490 2214.720 ;
        RECT 414.070 2214.660 414.390 2214.720 ;
        RECT 407.170 2214.520 414.390 2214.660 ;
        RECT 407.170 2214.460 407.490 2214.520 ;
        RECT 414.070 2214.460 414.390 2214.520 ;
        RECT 434.310 2214.660 434.630 2214.720 ;
        RECT 439.830 2214.660 440.150 2214.720 ;
        RECT 434.310 2214.520 440.150 2214.660 ;
        RECT 434.310 2214.460 434.630 2214.520 ;
        RECT 439.830 2214.460 440.150 2214.520 ;
        RECT 441.210 2214.660 441.530 2214.720 ;
        RECT 452.250 2214.660 452.570 2214.720 ;
        RECT 441.210 2214.520 452.570 2214.660 ;
        RECT 441.210 2214.460 441.530 2214.520 ;
        RECT 452.250 2214.460 452.570 2214.520 ;
        RECT 461.910 2214.660 462.230 2214.720 ;
        RECT 486.290 2214.660 486.610 2214.720 ;
        RECT 461.910 2214.520 486.610 2214.660 ;
        RECT 461.910 2214.460 462.230 2214.520 ;
        RECT 486.290 2214.460 486.610 2214.520 ;
        RECT 489.510 2214.660 489.830 2214.720 ;
        RECT 542.870 2214.660 543.190 2214.720 ;
        RECT 489.510 2214.520 543.190 2214.660 ;
        RECT 489.510 2214.460 489.830 2214.520 ;
        RECT 542.870 2214.460 543.190 2214.520 ;
        RECT 551.610 2214.660 551.930 2214.720 ;
        RECT 656.490 2214.660 656.810 2214.720 ;
        RECT 551.610 2214.520 656.810 2214.660 ;
        RECT 551.610 2214.460 551.930 2214.520 ;
        RECT 656.490 2214.460 656.810 2214.520 ;
        RECT 690.070 2214.660 690.390 2214.720 ;
        RECT 696.510 2214.660 696.830 2214.720 ;
        RECT 690.070 2214.520 696.830 2214.660 ;
        RECT 690.070 2214.460 690.390 2214.520 ;
        RECT 696.510 2214.460 696.830 2214.520 ;
        RECT 696.970 2214.660 697.290 2214.720 ;
        RECT 941.690 2214.660 942.010 2214.720 ;
        RECT 696.970 2214.520 942.010 2214.660 ;
        RECT 696.970 2214.460 697.290 2214.520 ;
        RECT 941.690 2214.460 942.010 2214.520 ;
        RECT 1030.010 2214.660 1030.330 2214.720 ;
        RECT 1038.750 2214.660 1039.070 2214.720 ;
        RECT 1030.010 2214.520 1039.070 2214.660 ;
        RECT 1030.010 2214.460 1030.330 2214.520 ;
        RECT 1038.750 2214.460 1039.070 2214.520 ;
        RECT 1041.050 2214.660 1041.370 2214.720 ;
        RECT 1045.650 2214.660 1045.970 2214.720 ;
        RECT 1041.050 2214.520 1045.970 2214.660 ;
        RECT 1041.050 2214.460 1041.370 2214.520 ;
        RECT 1045.650 2214.460 1045.970 2214.520 ;
        RECT 1124.310 2214.660 1124.630 2214.720 ;
        RECT 1346.950 2214.660 1347.270 2214.720 ;
        RECT 1124.310 2214.520 1347.270 2214.660 ;
        RECT 1124.310 2214.460 1124.630 2214.520 ;
        RECT 1346.950 2214.460 1347.270 2214.520 ;
        RECT 337.710 2214.320 338.030 2214.380 ;
        RECT 712.610 2214.320 712.930 2214.380 ;
        RECT 337.710 2214.180 712.930 2214.320 ;
        RECT 337.710 2214.120 338.030 2214.180 ;
        RECT 712.610 2214.120 712.930 2214.180 ;
        RECT 713.070 2214.320 713.390 2214.380 ;
        RECT 717.210 2214.320 717.530 2214.380 ;
        RECT 713.070 2214.180 717.530 2214.320 ;
        RECT 713.070 2214.120 713.390 2214.180 ;
        RECT 717.210 2214.120 717.530 2214.180 ;
        RECT 746.650 2214.320 746.970 2214.380 ;
        RECT 751.710 2214.320 752.030 2214.380 ;
        RECT 746.650 2214.180 752.030 2214.320 ;
        RECT 746.650 2214.120 746.970 2214.180 ;
        RECT 751.710 2214.120 752.030 2214.180 ;
        RECT 1131.210 2214.320 1131.530 2214.380 ;
        RECT 1358.450 2214.320 1358.770 2214.380 ;
        RECT 1131.210 2214.180 1358.770 2214.320 ;
        RECT 1131.210 2214.120 1131.530 2214.180 ;
        RECT 1358.450 2214.120 1358.770 2214.180 ;
        RECT 285.270 2213.980 285.590 2214.040 ;
        RECT 769.650 2213.980 769.970 2214.040 ;
        RECT 285.270 2213.840 769.970 2213.980 ;
        RECT 285.270 2213.780 285.590 2213.840 ;
        RECT 769.650 2213.780 769.970 2213.840 ;
        RECT 1007.470 2213.980 1007.790 2214.040 ;
        RECT 1038.290 2213.980 1038.610 2214.040 ;
        RECT 1007.470 2213.840 1038.610 2213.980 ;
        RECT 1007.470 2213.780 1007.790 2213.840 ;
        RECT 1038.290 2213.780 1038.610 2213.840 ;
        RECT 1130.750 2213.980 1131.070 2214.040 ;
        RECT 1369.490 2213.980 1369.810 2214.040 ;
        RECT 1130.750 2213.840 1369.810 2213.980 ;
        RECT 1130.750 2213.780 1131.070 2213.840 ;
        RECT 1369.490 2213.780 1369.810 2213.840 ;
        RECT 285.730 2213.640 286.050 2213.700 ;
        RECT 780.690 2213.640 781.010 2213.700 ;
        RECT 285.730 2213.500 781.010 2213.640 ;
        RECT 285.730 2213.440 286.050 2213.500 ;
        RECT 780.690 2213.440 781.010 2213.500 ;
        RECT 1138.110 2213.640 1138.430 2213.700 ;
        RECT 1380.990 2213.640 1381.310 2213.700 ;
        RECT 1138.110 2213.500 1381.310 2213.640 ;
        RECT 1138.110 2213.440 1138.430 2213.500 ;
        RECT 1380.990 2213.440 1381.310 2213.500 ;
        RECT 283.890 2213.300 284.210 2213.360 ;
        RECT 792.190 2213.300 792.510 2213.360 ;
        RECT 283.890 2213.160 792.510 2213.300 ;
        RECT 283.890 2213.100 284.210 2213.160 ;
        RECT 792.190 2213.100 792.510 2213.160 ;
        RECT 995.970 2213.300 996.290 2213.360 ;
        RECT 1031.390 2213.300 1031.710 2213.360 ;
        RECT 995.970 2213.160 1031.710 2213.300 ;
        RECT 995.970 2213.100 996.290 2213.160 ;
        RECT 1031.390 2213.100 1031.710 2213.160 ;
        RECT 1145.010 2213.300 1145.330 2213.360 ;
        RECT 1392.030 2213.300 1392.350 2213.360 ;
        RECT 1145.010 2213.160 1392.350 2213.300 ;
        RECT 1145.010 2213.100 1145.330 2213.160 ;
        RECT 1392.030 2213.100 1392.350 2213.160 ;
        RECT 286.650 2212.960 286.970 2213.020 ;
        RECT 803.230 2212.960 803.550 2213.020 ;
        RECT 286.650 2212.820 803.550 2212.960 ;
        RECT 286.650 2212.760 286.970 2212.820 ;
        RECT 803.230 2212.760 803.550 2212.820 ;
        RECT 939.390 2212.960 939.710 2213.020 ;
        RECT 944.910 2212.960 945.230 2213.020 ;
        RECT 939.390 2212.820 945.230 2212.960 ;
        RECT 939.390 2212.760 939.710 2212.820 ;
        RECT 944.910 2212.760 945.230 2212.820 ;
        RECT 1013.910 2212.960 1014.230 2213.020 ;
        RECT 1143.170 2212.960 1143.490 2213.020 ;
        RECT 1013.910 2212.820 1143.490 2212.960 ;
        RECT 1013.910 2212.760 1014.230 2212.820 ;
        RECT 1143.170 2212.760 1143.490 2212.820 ;
        RECT 1151.910 2212.960 1152.230 2213.020 ;
        RECT 1403.530 2212.960 1403.850 2213.020 ;
        RECT 1151.910 2212.820 1403.850 2212.960 ;
        RECT 1151.910 2212.760 1152.230 2212.820 ;
        RECT 1403.530 2212.760 1403.850 2212.820 ;
        RECT 344.150 2212.620 344.470 2212.680 ;
        RECT 893.850 2212.620 894.170 2212.680 ;
        RECT 344.150 2212.480 894.170 2212.620 ;
        RECT 344.150 2212.420 344.470 2212.480 ;
        RECT 893.850 2212.420 894.170 2212.480 ;
        RECT 1020.810 2212.620 1021.130 2212.680 ;
        RECT 1154.210 2212.620 1154.530 2212.680 ;
        RECT 1020.810 2212.480 1154.530 2212.620 ;
        RECT 1020.810 2212.420 1021.130 2212.480 ;
        RECT 1154.210 2212.420 1154.530 2212.480 ;
        RECT 1158.810 2212.620 1159.130 2212.680 ;
        RECT 1415.030 2212.620 1415.350 2212.680 ;
        RECT 1158.810 2212.480 1415.350 2212.620 ;
        RECT 1158.810 2212.420 1159.130 2212.480 ;
        RECT 1415.030 2212.420 1415.350 2212.480 ;
        RECT 350.590 2212.280 350.910 2212.340 ;
        RECT 905.350 2212.280 905.670 2212.340 ;
        RECT 350.590 2212.140 905.670 2212.280 ;
        RECT 350.590 2212.080 350.910 2212.140 ;
        RECT 905.350 2212.080 905.670 2212.140 ;
        RECT 1027.710 2212.280 1028.030 2212.340 ;
        RECT 1163.870 2212.280 1164.190 2212.340 ;
        RECT 1027.710 2212.140 1164.190 2212.280 ;
        RECT 1027.710 2212.080 1028.030 2212.140 ;
        RECT 1163.870 2212.080 1164.190 2212.140 ;
        RECT 1165.250 2212.280 1165.570 2212.340 ;
        RECT 1426.070 2212.280 1426.390 2212.340 ;
        RECT 1165.250 2212.140 1426.390 2212.280 ;
        RECT 1165.250 2212.080 1165.570 2212.140 ;
        RECT 1426.070 2212.080 1426.390 2212.140 ;
        RECT 351.050 2211.940 351.370 2212.000 ;
        RECT 916.850 2211.940 917.170 2212.000 ;
        RECT 351.050 2211.800 917.170 2211.940 ;
        RECT 351.050 2211.740 351.370 2211.800 ;
        RECT 916.850 2211.740 917.170 2211.800 ;
        RECT 973.430 2211.940 973.750 2212.000 ;
        RECT 1017.590 2211.940 1017.910 2212.000 ;
        RECT 973.430 2211.800 1017.910 2211.940 ;
        RECT 973.430 2211.740 973.750 2211.800 ;
        RECT 1017.590 2211.740 1017.910 2211.800 ;
        RECT 1034.610 2211.940 1034.930 2212.000 ;
        RECT 1177.210 2211.940 1177.530 2212.000 ;
        RECT 1034.610 2211.800 1177.530 2211.940 ;
        RECT 1034.610 2211.740 1034.930 2211.800 ;
        RECT 1177.210 2211.740 1177.530 2211.800 ;
        RECT 1179.510 2211.940 1179.830 2212.000 ;
        RECT 1460.110 2211.940 1460.430 2212.000 ;
        RECT 1179.510 2211.800 1460.430 2211.940 ;
        RECT 1179.510 2211.740 1179.830 2211.800 ;
        RECT 1460.110 2211.740 1460.430 2211.800 ;
        RECT 358.410 2211.600 358.730 2211.660 ;
        RECT 927.890 2211.600 928.210 2211.660 ;
        RECT 358.410 2211.460 928.210 2211.600 ;
        RECT 358.410 2211.400 358.730 2211.460 ;
        RECT 927.890 2211.400 928.210 2211.460 ;
        RECT 984.470 2211.600 984.790 2211.660 ;
        RECT 1024.490 2211.600 1024.810 2211.660 ;
        RECT 984.470 2211.460 1024.810 2211.600 ;
        RECT 984.470 2211.400 984.790 2211.460 ;
        RECT 1024.490 2211.400 1024.810 2211.460 ;
        RECT 1041.510 2211.600 1041.830 2211.660 ;
        RECT 1188.250 2211.600 1188.570 2211.660 ;
        RECT 1041.510 2211.460 1188.570 2211.600 ;
        RECT 1041.510 2211.400 1041.830 2211.460 ;
        RECT 1188.250 2211.400 1188.570 2211.460 ;
        RECT 1193.310 2211.600 1193.630 2211.660 ;
        RECT 1482.650 2211.600 1482.970 2211.660 ;
        RECT 1193.310 2211.460 1482.970 2211.600 ;
        RECT 1193.310 2211.400 1193.630 2211.460 ;
        RECT 1482.650 2211.400 1482.970 2211.460 ;
        RECT 284.810 2211.260 285.130 2211.320 ;
        RECT 950.430 2211.260 950.750 2211.320 ;
        RECT 284.810 2211.120 950.750 2211.260 ;
        RECT 284.810 2211.060 285.130 2211.120 ;
        RECT 950.430 2211.060 950.750 2211.120 ;
        RECT 961.930 2211.260 962.250 2211.320 ;
        RECT 1010.690 2211.260 1011.010 2211.320 ;
        RECT 961.930 2211.120 1011.010 2211.260 ;
        RECT 961.930 2211.060 962.250 2211.120 ;
        RECT 1010.690 2211.060 1011.010 2211.120 ;
        RECT 1048.410 2211.260 1048.730 2211.320 ;
        RECT 1199.750 2211.260 1200.070 2211.320 ;
        RECT 1048.410 2211.120 1200.070 2211.260 ;
        RECT 1048.410 2211.060 1048.730 2211.120 ;
        RECT 1199.750 2211.060 1200.070 2211.120 ;
        RECT 1210.330 2211.260 1210.650 2211.320 ;
        RECT 1231.030 2211.260 1231.350 2211.320 ;
        RECT 1210.330 2211.120 1231.350 2211.260 ;
        RECT 1210.330 2211.060 1210.650 2211.120 ;
        RECT 1231.030 2211.060 1231.350 2211.120 ;
        RECT 1231.490 2211.260 1231.810 2211.320 ;
        RECT 1256.330 2211.260 1256.650 2211.320 ;
        RECT 1231.490 2211.120 1256.650 2211.260 ;
        RECT 1231.490 2211.060 1231.810 2211.120 ;
        RECT 1256.330 2211.060 1256.650 2211.120 ;
        RECT 1256.790 2211.260 1257.110 2211.320 ;
        RECT 1494.150 2211.260 1494.470 2211.320 ;
        RECT 1256.790 2211.120 1494.470 2211.260 ;
        RECT 1256.790 2211.060 1257.110 2211.120 ;
        RECT 1494.150 2211.060 1494.470 2211.120 ;
        RECT 395.670 2210.920 395.990 2210.980 ;
        RECT 406.710 2210.920 407.030 2210.980 ;
        RECT 395.670 2210.780 407.030 2210.920 ;
        RECT 395.670 2210.720 395.990 2210.780 ;
        RECT 406.710 2210.720 407.030 2210.780 ;
        RECT 448.110 2210.920 448.430 2210.980 ;
        RECT 463.750 2210.920 464.070 2210.980 ;
        RECT 448.110 2210.780 464.070 2210.920 ;
        RECT 448.110 2210.720 448.430 2210.780 ;
        RECT 463.750 2210.720 464.070 2210.780 ;
        RECT 482.610 2210.920 482.930 2210.980 ;
        RECT 531.830 2210.920 532.150 2210.980 ;
        RECT 482.610 2210.780 532.150 2210.920 ;
        RECT 482.610 2210.720 482.930 2210.780 ;
        RECT 531.830 2210.720 532.150 2210.780 ;
        RECT 544.710 2210.920 545.030 2210.980 ;
        RECT 644.990 2210.920 645.310 2210.980 ;
        RECT 544.710 2210.780 645.310 2210.920 ;
        RECT 544.710 2210.720 545.030 2210.780 ;
        RECT 644.990 2210.720 645.310 2210.780 ;
        RECT 679.030 2210.920 679.350 2210.980 ;
        RECT 696.970 2210.920 697.290 2210.980 ;
        RECT 679.030 2210.780 697.290 2210.920 ;
        RECT 679.030 2210.720 679.350 2210.780 ;
        RECT 696.970 2210.720 697.290 2210.780 ;
        RECT 712.610 2210.920 712.930 2210.980 ;
        RECT 758.150 2210.920 758.470 2210.980 ;
        RECT 712.610 2210.780 758.470 2210.920 ;
        RECT 712.610 2210.720 712.930 2210.780 ;
        RECT 758.150 2210.720 758.470 2210.780 ;
        RECT 871.310 2210.920 871.630 2210.980 ;
        RECT 875.910 2210.920 876.230 2210.980 ;
        RECT 871.310 2210.780 876.230 2210.920 ;
        RECT 871.310 2210.720 871.630 2210.780 ;
        RECT 875.910 2210.720 876.230 2210.780 ;
        RECT 1117.410 2210.920 1117.730 2210.980 ;
        RECT 1335.450 2210.920 1335.770 2210.980 ;
        RECT 1117.410 2210.780 1335.770 2210.920 ;
        RECT 1117.410 2210.720 1117.730 2210.780 ;
        RECT 1335.450 2210.720 1335.770 2210.780 ;
        RECT 475.710 2210.580 476.030 2210.640 ;
        RECT 520.330 2210.580 520.650 2210.640 ;
        RECT 475.710 2210.440 520.650 2210.580 ;
        RECT 475.710 2210.380 476.030 2210.440 ;
        RECT 520.330 2210.380 520.650 2210.440 ;
        RECT 530.910 2210.580 531.230 2210.640 ;
        RECT 622.450 2210.580 622.770 2210.640 ;
        RECT 530.910 2210.440 622.770 2210.580 ;
        RECT 530.910 2210.380 531.230 2210.440 ;
        RECT 622.450 2210.380 622.770 2210.440 ;
        RECT 1103.610 2210.580 1103.930 2210.640 ;
        RECT 1312.910 2210.580 1313.230 2210.640 ;
        RECT 1103.610 2210.440 1313.230 2210.580 ;
        RECT 1103.610 2210.380 1103.930 2210.440 ;
        RECT 1312.910 2210.380 1313.230 2210.440 ;
        RECT 468.350 2210.240 468.670 2210.300 ;
        RECT 509.290 2210.240 509.610 2210.300 ;
        RECT 468.350 2210.100 509.610 2210.240 ;
        RECT 468.350 2210.040 468.670 2210.100 ;
        RECT 509.290 2210.040 509.610 2210.100 ;
        RECT 537.810 2210.240 538.130 2210.300 ;
        RECT 633.490 2210.240 633.810 2210.300 ;
        RECT 537.810 2210.100 633.810 2210.240 ;
        RECT 537.810 2210.040 538.130 2210.100 ;
        RECT 633.490 2210.040 633.810 2210.100 ;
        RECT 1110.510 2210.240 1110.830 2210.300 ;
        RECT 1324.410 2210.240 1324.730 2210.300 ;
        RECT 1110.510 2210.100 1324.730 2210.240 ;
        RECT 1110.510 2210.040 1110.830 2210.100 ;
        RECT 1324.410 2210.040 1324.730 2210.100 ;
        RECT 468.810 2209.900 469.130 2209.960 ;
        RECT 497.790 2209.900 498.110 2209.960 ;
        RECT 468.810 2209.760 498.110 2209.900 ;
        RECT 468.810 2209.700 469.130 2209.760 ;
        RECT 497.790 2209.700 498.110 2209.760 ;
        RECT 524.010 2209.900 524.330 2209.960 ;
        RECT 610.950 2209.900 611.270 2209.960 ;
        RECT 524.010 2209.760 611.270 2209.900 ;
        RECT 524.010 2209.700 524.330 2209.760 ;
        RECT 610.950 2209.700 611.270 2209.760 ;
        RECT 848.770 2209.900 849.090 2209.960 ;
        RECT 855.210 2209.900 855.530 2209.960 ;
        RECT 848.770 2209.760 855.530 2209.900 ;
        RECT 848.770 2209.700 849.090 2209.760 ;
        RECT 855.210 2209.700 855.530 2209.760 ;
        RECT 1089.350 2209.900 1089.670 2209.960 ;
        RECT 1290.370 2209.900 1290.690 2209.960 ;
        RECT 1089.350 2209.760 1290.690 2209.900 ;
        RECT 1089.350 2209.700 1089.670 2209.760 ;
        RECT 1290.370 2209.700 1290.690 2209.760 ;
        RECT 509.750 2209.560 510.070 2209.620 ;
        RECT 588.410 2209.560 588.730 2209.620 ;
        RECT 509.750 2209.420 588.730 2209.560 ;
        RECT 509.750 2209.360 510.070 2209.420 ;
        RECT 588.410 2209.360 588.730 2209.420 ;
        RECT 1018.510 2209.560 1018.830 2209.620 ;
        RECT 1045.190 2209.560 1045.510 2209.620 ;
        RECT 1018.510 2209.420 1045.510 2209.560 ;
        RECT 1018.510 2209.360 1018.830 2209.420 ;
        RECT 1045.190 2209.360 1045.510 2209.420 ;
        RECT 1096.710 2209.560 1097.030 2209.620 ;
        RECT 1301.410 2209.560 1301.730 2209.620 ;
        RECT 1096.710 2209.420 1301.730 2209.560 ;
        RECT 1096.710 2209.360 1097.030 2209.420 ;
        RECT 1301.410 2209.360 1301.730 2209.420 ;
        RECT 517.110 2209.220 517.430 2209.280 ;
        RECT 599.450 2209.220 599.770 2209.280 ;
        RECT 517.110 2209.080 599.770 2209.220 ;
        RECT 517.110 2209.020 517.430 2209.080 ;
        RECT 599.450 2209.020 599.770 2209.080 ;
        RECT 1069.110 2209.220 1069.430 2209.280 ;
        RECT 1224.590 2209.220 1224.910 2209.280 ;
        RECT 1267.830 2209.220 1268.150 2209.280 ;
        RECT 1069.110 2209.080 1224.360 2209.220 ;
        RECT 1069.110 2209.020 1069.430 2209.080 ;
        RECT 455.010 2208.880 455.330 2208.940 ;
        RECT 475.250 2208.880 475.570 2208.940 ;
        RECT 455.010 2208.740 475.570 2208.880 ;
        RECT 455.010 2208.680 455.330 2208.740 ;
        RECT 475.250 2208.680 475.570 2208.740 ;
        RECT 503.310 2208.880 503.630 2208.940 ;
        RECT 565.870 2208.880 566.190 2208.940 ;
        RECT 503.310 2208.740 566.190 2208.880 ;
        RECT 503.310 2208.680 503.630 2208.740 ;
        RECT 565.870 2208.680 566.190 2208.740 ;
        RECT 1055.310 2208.880 1055.630 2208.940 ;
        RECT 1222.290 2208.880 1222.610 2208.940 ;
        RECT 1055.310 2208.740 1222.610 2208.880 ;
        RECT 1224.220 2208.880 1224.360 2209.080 ;
        RECT 1224.590 2209.080 1268.150 2209.220 ;
        RECT 1224.590 2209.020 1224.910 2209.080 ;
        RECT 1267.830 2209.020 1268.150 2209.080 ;
        RECT 1242.990 2208.880 1243.310 2208.940 ;
        RECT 1224.220 2208.740 1243.310 2208.880 ;
        RECT 1055.310 2208.680 1055.630 2208.740 ;
        RECT 1222.290 2208.680 1222.610 2208.740 ;
        RECT 1242.990 2208.680 1243.310 2208.740 ;
        RECT 1243.450 2208.880 1243.770 2208.940 ;
        RECT 1256.790 2208.880 1257.110 2208.940 ;
        RECT 1243.450 2208.740 1257.110 2208.880 ;
        RECT 1243.450 2208.680 1243.770 2208.740 ;
        RECT 1256.790 2208.680 1257.110 2208.740 ;
        RECT 510.210 2208.540 510.530 2208.600 ;
        RECT 576.910 2208.540 577.230 2208.600 ;
        RECT 510.210 2208.400 577.230 2208.540 ;
        RECT 510.210 2208.340 510.530 2208.400 ;
        RECT 576.910 2208.340 577.230 2208.400 ;
        RECT 1062.210 2208.540 1062.530 2208.600 ;
        RECT 1210.330 2208.540 1210.650 2208.600 ;
        RECT 1062.210 2208.400 1210.650 2208.540 ;
        RECT 1062.210 2208.340 1062.530 2208.400 ;
        RECT 1210.330 2208.340 1210.650 2208.400 ;
        RECT 496.410 2208.200 496.730 2208.260 ;
        RECT 554.370 2208.200 554.690 2208.260 ;
        RECT 496.410 2208.060 554.690 2208.200 ;
        RECT 496.410 2208.000 496.730 2208.060 ;
        RECT 554.370 2208.000 554.690 2208.060 ;
        RECT 1054.850 2208.200 1055.170 2208.260 ;
        RECT 1211.250 2208.200 1211.570 2208.260 ;
        RECT 1054.850 2208.060 1211.570 2208.200 ;
        RECT 1054.850 2208.000 1055.170 2208.060 ;
        RECT 1211.250 2208.000 1211.570 2208.060 ;
        RECT 1225.510 2208.200 1225.830 2208.260 ;
        RECT 1278.870 2208.200 1279.190 2208.260 ;
        RECT 1225.510 2208.060 1279.190 2208.200 ;
        RECT 1225.510 2208.000 1225.830 2208.060 ;
        RECT 1278.870 2208.000 1279.190 2208.060 ;
      LAYER met1 ;
        RECT 305.130 1004.460 1494.550 2189.280 ;
      LAYER met1 ;
        RECT 1513.930 2187.120 1514.250 2187.180 ;
        RECT 2335.490 2187.120 2335.810 2187.180 ;
        RECT 1513.930 2186.980 2335.810 2187.120 ;
        RECT 1513.930 2186.920 1514.250 2186.980 ;
        RECT 2335.490 2186.920 2335.810 2186.980 ;
        RECT 1513.930 2173.520 1514.250 2173.580 ;
        RECT 1617.430 2173.520 1617.750 2173.580 ;
        RECT 1513.930 2173.380 1617.750 2173.520 ;
        RECT 1513.930 2173.320 1514.250 2173.380 ;
        RECT 1617.430 2173.320 1617.750 2173.380 ;
        RECT 1637.670 2173.520 1637.990 2173.580 ;
        RECT 1638.130 2173.520 1638.450 2173.580 ;
        RECT 1637.670 2173.380 1638.450 2173.520 ;
        RECT 1637.670 2173.320 1637.990 2173.380 ;
        RECT 1638.130 2173.320 1638.450 2173.380 ;
        RECT 1638.590 2173.520 1638.910 2173.580 ;
        RECT 2328.590 2173.520 2328.910 2173.580 ;
        RECT 1638.590 2173.380 2328.910 2173.520 ;
        RECT 1638.590 2173.320 1638.910 2173.380 ;
        RECT 2328.590 2173.320 2328.910 2173.380 ;
        RECT 1617.430 2172.500 1617.750 2172.560 ;
        RECT 1638.590 2172.500 1638.910 2172.560 ;
        RECT 1617.430 2172.360 1638.910 2172.500 ;
        RECT 1617.430 2172.300 1617.750 2172.360 ;
        RECT 1638.590 2172.300 1638.910 2172.360 ;
        RECT 1513.930 2166.380 1514.250 2166.440 ;
        RECT 2321.690 2166.380 2322.010 2166.440 ;
        RECT 1513.930 2166.240 2322.010 2166.380 ;
        RECT 1513.930 2166.180 1514.250 2166.240 ;
        RECT 2321.690 2166.180 2322.010 2166.240 ;
        RECT 1513.930 2152.780 1514.250 2152.840 ;
        RECT 1770.150 2152.780 1770.470 2152.840 ;
        RECT 1513.930 2152.640 1770.470 2152.780 ;
        RECT 1513.930 2152.580 1514.250 2152.640 ;
        RECT 1770.150 2152.580 1770.470 2152.640 ;
        RECT 1513.930 2145.640 1514.250 2145.700 ;
        RECT 1769.690 2145.640 1770.010 2145.700 ;
        RECT 1513.930 2145.500 1770.010 2145.640 ;
        RECT 1513.930 2145.440 1514.250 2145.500 ;
        RECT 1769.690 2145.440 1770.010 2145.500 ;
        RECT 1513.930 2132.040 1514.250 2132.100 ;
        RECT 1763.710 2132.040 1764.030 2132.100 ;
        RECT 1513.930 2131.900 1764.030 2132.040 ;
        RECT 1513.930 2131.840 1514.250 2131.900 ;
        RECT 1763.710 2131.840 1764.030 2131.900 ;
        RECT 1637.670 2118.440 1637.990 2118.500 ;
        RECT 1638.130 2118.440 1638.450 2118.500 ;
        RECT 1637.670 2118.300 1638.450 2118.440 ;
        RECT 1637.670 2118.240 1637.990 2118.300 ;
        RECT 1638.130 2118.240 1638.450 2118.300 ;
        RECT 1513.930 2118.100 1514.250 2118.160 ;
        RECT 1763.250 2118.100 1763.570 2118.160 ;
        RECT 1513.930 2117.960 1763.570 2118.100 ;
        RECT 1513.930 2117.900 1514.250 2117.960 ;
        RECT 1763.250 2117.900 1763.570 2117.960 ;
        RECT 1513.930 2111.300 1514.250 2111.360 ;
        RECT 1762.790 2111.300 1763.110 2111.360 ;
        RECT 1513.930 2111.160 1763.110 2111.300 ;
        RECT 1513.930 2111.100 1514.250 2111.160 ;
        RECT 1762.790 2111.100 1763.110 2111.160 ;
        RECT 1513.930 2097.360 1514.250 2097.420 ;
        RECT 1755.890 2097.360 1756.210 2097.420 ;
        RECT 1513.930 2097.220 1756.210 2097.360 ;
        RECT 1513.930 2097.160 1514.250 2097.220 ;
        RECT 1755.890 2097.160 1756.210 2097.220 ;
        RECT 1513.930 2090.560 1514.250 2090.620 ;
        RECT 1748.990 2090.560 1749.310 2090.620 ;
        RECT 1513.930 2090.420 1749.310 2090.560 ;
        RECT 1513.930 2090.360 1514.250 2090.420 ;
        RECT 1748.990 2090.360 1749.310 2090.420 ;
        RECT 1513.930 2076.960 1514.250 2077.020 ;
        RECT 1735.190 2076.960 1735.510 2077.020 ;
        RECT 1513.930 2076.820 1735.510 2076.960 ;
        RECT 1513.930 2076.760 1514.250 2076.820 ;
        RECT 1735.190 2076.760 1735.510 2076.820 ;
        RECT 1637.670 2069.820 1637.990 2069.880 ;
        RECT 1638.590 2069.820 1638.910 2069.880 ;
        RECT 1637.670 2069.680 1638.910 2069.820 ;
        RECT 1637.670 2069.620 1637.990 2069.680 ;
        RECT 1638.590 2069.620 1638.910 2069.680 ;
        RECT 1513.930 2063.020 1514.250 2063.080 ;
        RECT 2381.030 2063.020 2381.350 2063.080 ;
        RECT 1513.930 2062.880 2381.350 2063.020 ;
        RECT 1513.930 2062.820 1514.250 2062.880 ;
        RECT 2381.030 2062.820 2381.350 2062.880 ;
        RECT 1513.930 2056.220 1514.250 2056.280 ;
        RECT 2373.670 2056.220 2373.990 2056.280 ;
        RECT 1513.930 2056.080 2373.990 2056.220 ;
        RECT 1513.930 2056.020 1514.250 2056.080 ;
        RECT 2373.670 2056.020 2373.990 2056.080 ;
        RECT 1513.930 2042.280 1514.250 2042.340 ;
        RECT 2366.770 2042.280 2367.090 2042.340 ;
        RECT 1513.930 2042.140 2367.090 2042.280 ;
        RECT 1513.930 2042.080 1514.250 2042.140 ;
        RECT 2366.770 2042.080 2367.090 2042.140 ;
        RECT 1513.930 2035.480 1514.250 2035.540 ;
        RECT 2359.870 2035.480 2360.190 2035.540 ;
        RECT 1513.930 2035.340 2360.190 2035.480 ;
        RECT 1513.930 2035.280 1514.250 2035.340 ;
        RECT 2359.870 2035.280 2360.190 2035.340 ;
        RECT 1637.670 2021.880 1637.990 2021.940 ;
        RECT 1638.590 2021.880 1638.910 2021.940 ;
        RECT 1637.670 2021.740 1638.910 2021.880 ;
        RECT 1637.670 2021.680 1637.990 2021.740 ;
        RECT 1638.590 2021.680 1638.910 2021.740 ;
        RECT 1513.470 2021.540 1513.790 2021.600 ;
        RECT 2352.970 2021.540 2353.290 2021.600 ;
        RECT 1513.470 2021.400 2353.290 2021.540 ;
        RECT 1513.470 2021.340 1513.790 2021.400 ;
        RECT 2352.970 2021.340 2353.290 2021.400 ;
        RECT 1513.930 2007.940 1514.250 2008.000 ;
        RECT 2346.070 2007.940 2346.390 2008.000 ;
        RECT 1513.930 2007.800 2346.390 2007.940 ;
        RECT 1513.930 2007.740 1514.250 2007.800 ;
        RECT 2346.070 2007.740 2346.390 2007.800 ;
        RECT 1513.930 2000.800 1514.250 2000.860 ;
        RECT 2339.630 2000.800 2339.950 2000.860 ;
        RECT 1513.930 2000.660 2339.950 2000.800 ;
        RECT 1513.930 2000.600 1514.250 2000.660 ;
        RECT 2339.630 2000.600 2339.950 2000.660 ;
        RECT 1513.930 1987.200 1514.250 1987.260 ;
        RECT 2339.170 1987.200 2339.490 1987.260 ;
        RECT 1513.930 1987.060 2339.490 1987.200 ;
        RECT 1513.930 1987.000 1514.250 1987.060 ;
        RECT 2339.170 1987.000 2339.490 1987.060 ;
        RECT 1512.550 1980.060 1512.870 1980.120 ;
        RECT 2332.270 1980.060 2332.590 1980.120 ;
        RECT 1512.550 1979.920 2332.590 1980.060 ;
        RECT 1512.550 1979.860 1512.870 1979.920 ;
        RECT 2332.270 1979.860 2332.590 1979.920 ;
        RECT 1637.670 1973.260 1637.990 1973.320 ;
        RECT 1638.130 1973.260 1638.450 1973.320 ;
        RECT 1637.670 1973.120 1638.450 1973.260 ;
        RECT 1637.670 1973.060 1637.990 1973.120 ;
        RECT 1638.130 1973.060 1638.450 1973.120 ;
        RECT 1513.470 1966.460 1513.790 1966.520 ;
        RECT 2325.370 1966.460 2325.690 1966.520 ;
        RECT 1513.470 1966.320 2325.690 1966.460 ;
        RECT 1513.470 1966.260 1513.790 1966.320 ;
        RECT 2325.370 1966.260 2325.690 1966.320 ;
        RECT 1513.930 1952.520 1514.250 1952.580 ;
        RECT 2318.470 1952.520 2318.790 1952.580 ;
        RECT 1513.930 1952.380 2318.790 1952.520 ;
        RECT 1513.930 1952.320 1514.250 1952.380 ;
        RECT 2318.470 1952.320 2318.790 1952.380 ;
        RECT 1513.930 1945.720 1514.250 1945.780 ;
        RECT 2311.570 1945.720 2311.890 1945.780 ;
        RECT 1513.930 1945.580 2311.890 1945.720 ;
        RECT 1513.930 1945.520 1514.250 1945.580 ;
        RECT 2311.570 1945.520 2311.890 1945.580 ;
        RECT 1512.550 1931.780 1512.870 1931.840 ;
        RECT 2305.130 1931.780 2305.450 1931.840 ;
        RECT 1512.550 1931.640 2305.450 1931.780 ;
        RECT 1512.550 1931.580 1512.870 1931.640 ;
        RECT 2305.130 1931.580 2305.450 1931.640 ;
        RECT 1638.130 1925.320 1638.450 1925.380 ;
        RECT 1639.050 1925.320 1639.370 1925.380 ;
        RECT 1638.130 1925.180 1639.370 1925.320 ;
        RECT 1638.130 1925.120 1638.450 1925.180 ;
        RECT 1639.050 1925.120 1639.370 1925.180 ;
        RECT 1512.550 1924.980 1512.870 1925.040 ;
        RECT 2304.670 1924.980 2304.990 1925.040 ;
        RECT 1512.550 1924.840 2304.990 1924.980 ;
        RECT 1512.550 1924.780 1512.870 1924.840 ;
        RECT 2304.670 1924.780 2304.990 1924.840 ;
        RECT 1513.930 1911.040 1514.250 1911.100 ;
        RECT 2218.190 1911.040 2218.510 1911.100 ;
        RECT 1513.930 1910.900 2218.510 1911.040 ;
        RECT 1513.930 1910.840 1514.250 1910.900 ;
        RECT 2218.190 1910.840 2218.510 1910.900 ;
        RECT 1513.010 1904.240 1513.330 1904.300 ;
        RECT 1797.290 1904.240 1797.610 1904.300 ;
        RECT 1513.010 1904.100 1797.610 1904.240 ;
        RECT 1513.010 1904.040 1513.330 1904.100 ;
        RECT 1797.290 1904.040 1797.610 1904.100 ;
        RECT 1513.930 1890.640 1514.250 1890.700 ;
        RECT 1790.390 1890.640 1790.710 1890.700 ;
        RECT 1513.930 1890.500 1790.710 1890.640 ;
        RECT 1513.930 1890.440 1514.250 1890.500 ;
        RECT 1790.390 1890.440 1790.710 1890.500 ;
        RECT 1638.130 1883.840 1638.450 1883.900 ;
        RECT 1639.050 1883.840 1639.370 1883.900 ;
        RECT 1638.130 1883.700 1639.370 1883.840 ;
        RECT 1638.130 1883.640 1638.450 1883.700 ;
        RECT 1639.050 1883.640 1639.370 1883.700 ;
        RECT 1513.930 1876.700 1514.250 1876.760 ;
        RECT 1783.490 1876.700 1783.810 1876.760 ;
        RECT 1513.930 1876.560 1783.810 1876.700 ;
        RECT 1513.930 1876.500 1514.250 1876.560 ;
        RECT 1783.490 1876.500 1783.810 1876.560 ;
        RECT 1513.930 1869.900 1514.250 1869.960 ;
        RECT 1776.590 1869.900 1776.910 1869.960 ;
        RECT 1513.930 1869.760 1776.910 1869.900 ;
        RECT 1513.930 1869.700 1514.250 1869.760 ;
        RECT 1776.590 1869.700 1776.910 1869.760 ;
        RECT 1511.630 1855.960 1511.950 1856.020 ;
        RECT 1714.490 1855.960 1714.810 1856.020 ;
        RECT 1511.630 1855.820 1714.810 1855.960 ;
        RECT 1511.630 1855.760 1511.950 1855.820 ;
        RECT 1714.490 1855.760 1714.810 1855.820 ;
        RECT 1513.010 1849.160 1513.330 1849.220 ;
        RECT 2263.730 1849.160 2264.050 1849.220 ;
        RECT 1513.010 1849.020 2264.050 1849.160 ;
        RECT 1513.010 1848.960 1513.330 1849.020 ;
        RECT 2263.730 1848.960 2264.050 1849.020 ;
        RECT 1513.930 1835.220 1514.250 1835.280 ;
        RECT 1652.390 1835.220 1652.710 1835.280 ;
        RECT 1513.930 1835.080 1652.710 1835.220 ;
        RECT 1513.930 1835.020 1514.250 1835.080 ;
        RECT 1652.390 1835.020 1652.710 1835.080 ;
        RECT 1512.550 1821.620 1512.870 1821.680 ;
        RECT 1646.410 1821.620 1646.730 1821.680 ;
        RECT 1512.550 1821.480 1646.730 1821.620 ;
        RECT 1512.550 1821.420 1512.870 1821.480 ;
        RECT 1646.410 1821.420 1646.730 1821.480 ;
        RECT 1512.090 1814.480 1512.410 1814.540 ;
        RECT 1645.490 1814.480 1645.810 1814.540 ;
        RECT 1512.090 1814.340 1645.810 1814.480 ;
        RECT 1512.090 1814.280 1512.410 1814.340 ;
        RECT 1645.490 1814.280 1645.810 1814.340 ;
        RECT 1511.630 1800.880 1511.950 1800.940 ;
        RECT 1640.430 1800.880 1640.750 1800.940 ;
        RECT 1511.630 1800.740 1640.750 1800.880 ;
        RECT 1511.630 1800.680 1511.950 1800.740 ;
        RECT 1640.430 1800.680 1640.750 1800.740 ;
        RECT 1512.550 1793.740 1512.870 1793.800 ;
        RECT 1631.690 1793.740 1632.010 1793.800 ;
        RECT 1512.550 1793.600 1632.010 1793.740 ;
        RECT 1512.550 1793.540 1512.870 1793.600 ;
        RECT 1631.690 1793.540 1632.010 1793.600 ;
        RECT 1513.930 1780.140 1514.250 1780.200 ;
        RECT 1624.790 1780.140 1625.110 1780.200 ;
        RECT 1513.930 1780.000 1625.110 1780.140 ;
        RECT 1513.930 1779.940 1514.250 1780.000 ;
        RECT 1624.790 1779.940 1625.110 1780.000 ;
        RECT 1513.930 1766.200 1514.250 1766.260 ;
        RECT 1617.890 1766.200 1618.210 1766.260 ;
        RECT 1513.930 1766.060 1618.210 1766.200 ;
        RECT 1513.930 1766.000 1514.250 1766.060 ;
        RECT 1617.890 1766.000 1618.210 1766.060 ;
        RECT 1512.090 1759.400 1512.410 1759.460 ;
        RECT 1610.990 1759.400 1611.310 1759.460 ;
        RECT 1512.090 1759.260 1611.310 1759.400 ;
        RECT 1512.090 1759.200 1512.410 1759.260 ;
        RECT 1610.990 1759.200 1611.310 1759.260 ;
        RECT 1513.470 1745.460 1513.790 1745.520 ;
        RECT 2301.910 1745.460 2302.230 1745.520 ;
        RECT 1513.470 1745.320 2302.230 1745.460 ;
        RECT 1513.470 1745.260 1513.790 1745.320 ;
        RECT 2301.910 1745.260 2302.230 1745.320 ;
        RECT 1512.550 1738.660 1512.870 1738.720 ;
        RECT 2300.990 1738.660 2301.310 1738.720 ;
        RECT 1512.550 1738.520 2301.310 1738.660 ;
        RECT 1512.550 1738.460 1512.870 1738.520 ;
        RECT 2300.990 1738.460 2301.310 1738.520 ;
        RECT 1513.930 1725.060 1514.250 1725.120 ;
        RECT 2294.090 1725.060 2294.410 1725.120 ;
        RECT 1513.930 1724.920 2294.410 1725.060 ;
        RECT 1513.930 1724.860 1514.250 1724.920 ;
        RECT 2294.090 1724.860 2294.410 1724.920 ;
        RECT 1513.930 1711.120 1514.250 1711.180 ;
        RECT 2287.190 1711.120 2287.510 1711.180 ;
        RECT 1513.930 1710.980 2287.510 1711.120 ;
        RECT 1513.930 1710.920 1514.250 1710.980 ;
        RECT 2287.190 1710.920 2287.510 1710.980 ;
        RECT 1512.090 1704.320 1512.410 1704.380 ;
        RECT 2280.290 1704.320 2280.610 1704.380 ;
        RECT 1512.090 1704.180 2280.610 1704.320 ;
        RECT 1512.090 1704.120 1512.410 1704.180 ;
        RECT 2280.290 1704.120 2280.610 1704.180 ;
        RECT 1513.470 1690.380 1513.790 1690.440 ;
        RECT 2273.390 1690.380 2273.710 1690.440 ;
        RECT 1513.470 1690.240 2273.710 1690.380 ;
        RECT 1513.470 1690.180 1513.790 1690.240 ;
        RECT 2273.390 1690.180 2273.710 1690.240 ;
        RECT 1512.550 1683.580 1512.870 1683.640 ;
        RECT 2267.410 1683.580 2267.730 1683.640 ;
        RECT 1512.550 1683.440 2267.730 1683.580 ;
        RECT 1512.550 1683.380 1512.870 1683.440 ;
        RECT 2267.410 1683.380 2267.730 1683.440 ;
        RECT 1513.930 1669.640 1514.250 1669.700 ;
        RECT 2266.490 1669.640 2266.810 1669.700 ;
        RECT 1513.930 1669.500 2266.810 1669.640 ;
        RECT 1513.930 1669.440 1514.250 1669.500 ;
        RECT 2266.490 1669.440 2266.810 1669.500 ;
        RECT 1512.550 1655.700 1512.870 1655.760 ;
        RECT 1529.110 1655.700 1529.430 1655.760 ;
        RECT 1512.550 1655.560 1529.430 1655.700 ;
        RECT 1512.550 1655.500 1512.870 1655.560 ;
        RECT 1529.110 1655.500 1529.430 1655.560 ;
        RECT 1511.630 1647.200 1511.950 1647.260 ;
        RECT 1522.210 1647.200 1522.530 1647.260 ;
        RECT 1511.630 1647.060 1522.530 1647.200 ;
        RECT 1511.630 1647.000 1511.950 1647.060 ;
        RECT 1522.210 1647.000 1522.530 1647.060 ;
        RECT 1512.550 1634.620 1512.870 1634.680 ;
        RECT 1528.650 1634.620 1528.970 1634.680 ;
        RECT 1512.550 1634.480 1528.970 1634.620 ;
        RECT 1512.550 1634.420 1512.870 1634.480 ;
        RECT 1528.650 1634.420 1528.970 1634.480 ;
        RECT 1511.630 1622.380 1511.950 1622.440 ;
        RECT 1521.750 1622.380 1522.070 1622.440 ;
        RECT 1511.630 1622.240 1522.070 1622.380 ;
        RECT 1511.630 1622.180 1511.950 1622.240 ;
        RECT 1521.750 1622.180 1522.070 1622.240 ;
        RECT 1511.630 1613.540 1511.950 1613.600 ;
        RECT 1528.190 1613.540 1528.510 1613.600 ;
        RECT 1511.630 1613.400 1528.510 1613.540 ;
        RECT 1511.630 1613.340 1511.950 1613.400 ;
        RECT 1528.190 1613.340 1528.510 1613.400 ;
        RECT 1511.630 1600.620 1511.950 1600.680 ;
        RECT 1521.290 1600.620 1521.610 1600.680 ;
        RECT 1511.630 1600.480 1521.610 1600.620 ;
        RECT 1511.630 1600.420 1511.950 1600.480 ;
        RECT 1521.290 1600.420 1521.610 1600.480 ;
        RECT 1513.470 1591.780 1513.790 1591.840 ;
        RECT 1535.090 1591.780 1535.410 1591.840 ;
        RECT 1513.470 1591.640 1535.410 1591.780 ;
        RECT 1513.470 1591.580 1513.790 1591.640 ;
        RECT 1535.090 1591.580 1535.410 1591.640 ;
        RECT 1513.930 1579.880 1514.250 1579.940 ;
        RECT 1580.170 1579.880 1580.490 1579.940 ;
        RECT 1513.930 1579.740 1580.490 1579.880 ;
        RECT 1513.930 1579.680 1514.250 1579.740 ;
        RECT 1580.170 1579.680 1580.490 1579.740 ;
        RECT 1513.930 1573.080 1514.250 1573.140 ;
        RECT 1997.390 1573.080 1997.710 1573.140 ;
        RECT 1513.930 1572.940 1997.710 1573.080 ;
        RECT 1513.930 1572.880 1514.250 1572.940 ;
        RECT 1997.390 1572.880 1997.710 1572.940 ;
        RECT 1513.470 1559.140 1513.790 1559.200 ;
        RECT 1990.490 1559.140 1990.810 1559.200 ;
        RECT 1513.470 1559.000 1990.810 1559.140 ;
        RECT 1513.470 1558.940 1513.790 1559.000 ;
        RECT 1990.490 1558.940 1990.810 1559.000 ;
        RECT 1513.930 1545.540 1514.250 1545.600 ;
        RECT 1976.690 1545.540 1977.010 1545.600 ;
        RECT 1513.930 1545.400 1977.010 1545.540 ;
        RECT 1513.930 1545.340 1514.250 1545.400 ;
        RECT 1976.690 1545.340 1977.010 1545.400 ;
        RECT 1513.930 1538.740 1514.250 1538.800 ;
        RECT 1969.790 1538.740 1970.110 1538.800 ;
        RECT 1513.930 1538.600 1970.110 1538.740 ;
        RECT 1513.930 1538.540 1514.250 1538.600 ;
        RECT 1969.790 1538.540 1970.110 1538.600 ;
        RECT 1513.930 1524.800 1514.250 1524.860 ;
        RECT 1962.890 1524.800 1963.210 1524.860 ;
        RECT 1513.930 1524.660 1963.210 1524.800 ;
        RECT 1513.930 1524.600 1514.250 1524.660 ;
        RECT 1962.890 1524.600 1963.210 1524.660 ;
        RECT 1513.930 1518.000 1514.250 1518.060 ;
        RECT 1955.990 1518.000 1956.310 1518.060 ;
        RECT 1513.930 1517.860 1956.310 1518.000 ;
        RECT 1513.930 1517.800 1514.250 1517.860 ;
        RECT 1955.990 1517.800 1956.310 1517.860 ;
        RECT 1513.470 1504.060 1513.790 1504.120 ;
        RECT 1942.190 1504.060 1942.510 1504.120 ;
        RECT 1513.470 1503.920 1942.510 1504.060 ;
        RECT 1513.470 1503.860 1513.790 1503.920 ;
        RECT 1942.190 1503.860 1942.510 1503.920 ;
        RECT 1513.930 1490.460 1514.250 1490.520 ;
        RECT 2228.770 1490.460 2229.090 1490.520 ;
        RECT 1513.930 1490.320 2229.090 1490.460 ;
        RECT 1513.930 1490.260 1514.250 1490.320 ;
        RECT 2228.770 1490.260 2229.090 1490.320 ;
        RECT 1513.010 1479.580 1513.330 1479.640 ;
        RECT 1529.570 1479.580 1529.890 1479.640 ;
        RECT 1513.010 1479.440 1529.890 1479.580 ;
        RECT 1513.010 1479.380 1513.330 1479.440 ;
        RECT 1529.570 1479.380 1529.890 1479.440 ;
        RECT 1513.930 1469.720 1514.250 1469.780 ;
        RECT 2011.190 1469.720 2011.510 1469.780 ;
        RECT 1513.930 1469.580 2011.510 1469.720 ;
        RECT 1513.930 1469.520 1514.250 1469.580 ;
        RECT 2011.190 1469.520 2011.510 1469.580 ;
        RECT 1512.550 1462.580 1512.870 1462.640 ;
        RECT 1601.330 1462.580 1601.650 1462.640 ;
        RECT 1512.550 1462.440 1601.650 1462.580 ;
        RECT 1512.550 1462.380 1512.870 1462.440 ;
        RECT 1601.330 1462.380 1601.650 1462.440 ;
        RECT 1513.470 1448.980 1513.790 1449.040 ;
        RECT 1600.870 1448.980 1601.190 1449.040 ;
        RECT 1513.470 1448.840 1601.190 1448.980 ;
        RECT 1513.470 1448.780 1513.790 1448.840 ;
        RECT 1600.870 1448.780 1601.190 1448.840 ;
        RECT 1513.930 1435.040 1514.250 1435.100 ;
        RECT 1593.970 1435.040 1594.290 1435.100 ;
        RECT 1513.930 1434.900 1594.290 1435.040 ;
        RECT 1513.930 1434.840 1514.250 1434.900 ;
        RECT 1593.970 1434.840 1594.290 1434.900 ;
        RECT 1513.470 1426.540 1513.790 1426.600 ;
        RECT 1541.990 1426.540 1542.310 1426.600 ;
        RECT 1513.470 1426.400 1542.310 1426.540 ;
        RECT 1513.470 1426.340 1513.790 1426.400 ;
        RECT 1541.990 1426.340 1542.310 1426.400 ;
        RECT 1512.550 1414.300 1512.870 1414.360 ;
        RECT 2252.690 1414.300 2253.010 1414.360 ;
        RECT 1512.550 1414.160 2253.010 1414.300 ;
        RECT 1512.550 1414.100 1512.870 1414.160 ;
        RECT 2252.690 1414.100 2253.010 1414.160 ;
        RECT 1512.550 1407.500 1512.870 1407.560 ;
        RECT 2245.790 1407.500 2246.110 1407.560 ;
        RECT 1512.550 1407.360 2246.110 1407.500 ;
        RECT 1512.550 1407.300 1512.870 1407.360 ;
        RECT 2245.790 1407.300 2246.110 1407.360 ;
        RECT 1511.630 1393.560 1511.950 1393.620 ;
        RECT 2238.890 1393.560 2239.210 1393.620 ;
        RECT 1511.630 1393.420 2239.210 1393.560 ;
        RECT 1511.630 1393.360 1511.950 1393.420 ;
        RECT 2238.890 1393.360 2239.210 1393.420 ;
        RECT 1513.010 1386.760 1513.330 1386.820 ;
        RECT 2231.990 1386.760 2232.310 1386.820 ;
        RECT 1513.010 1386.620 2232.310 1386.760 ;
        RECT 1513.010 1386.560 1513.330 1386.620 ;
        RECT 2231.990 1386.560 2232.310 1386.620 ;
        RECT 1513.930 1373.160 1514.250 1373.220 ;
        RECT 1794.070 1373.160 1794.390 1373.220 ;
        RECT 1513.930 1373.020 1794.390 1373.160 ;
        RECT 1513.930 1372.960 1514.250 1373.020 ;
        RECT 1794.070 1372.960 1794.390 1373.020 ;
        RECT 1512.550 1359.220 1512.870 1359.280 ;
        RECT 1787.170 1359.220 1787.490 1359.280 ;
        RECT 1512.550 1359.080 1787.490 1359.220 ;
        RECT 1512.550 1359.020 1512.870 1359.080 ;
        RECT 1787.170 1359.020 1787.490 1359.080 ;
        RECT 1512.550 1352.420 1512.870 1352.480 ;
        RECT 1780.270 1352.420 1780.590 1352.480 ;
        RECT 1512.550 1352.280 1780.590 1352.420 ;
        RECT 1512.550 1352.220 1512.870 1352.280 ;
        RECT 1780.270 1352.220 1780.590 1352.280 ;
        RECT 1511.630 1338.480 1511.950 1338.540 ;
        RECT 1773.370 1338.480 1773.690 1338.540 ;
        RECT 1511.630 1338.340 1773.690 1338.480 ;
        RECT 1511.630 1338.280 1511.950 1338.340 ;
        RECT 1773.370 1338.280 1773.690 1338.340 ;
        RECT 1513.010 1331.680 1513.330 1331.740 ;
        RECT 1766.470 1331.680 1766.790 1331.740 ;
        RECT 1513.010 1331.540 1766.790 1331.680 ;
        RECT 1513.010 1331.480 1513.330 1331.540 ;
        RECT 1766.470 1331.480 1766.790 1331.540 ;
        RECT 1513.930 1317.740 1514.250 1317.800 ;
        RECT 1760.030 1317.740 1760.350 1317.800 ;
        RECT 1513.930 1317.600 1760.350 1317.740 ;
        RECT 1513.930 1317.540 1514.250 1317.600 ;
        RECT 1760.030 1317.540 1760.350 1317.600 ;
        RECT 1512.550 1304.140 1512.870 1304.200 ;
        RECT 1759.570 1304.140 1759.890 1304.200 ;
        RECT 1512.550 1304.000 1759.890 1304.140 ;
        RECT 1512.550 1303.940 1512.870 1304.000 ;
        RECT 1759.570 1303.940 1759.890 1304.000 ;
        RECT 1512.090 1297.000 1512.410 1297.060 ;
        RECT 1752.670 1297.000 1752.990 1297.060 ;
        RECT 1512.090 1296.860 1752.990 1297.000 ;
        RECT 1512.090 1296.800 1512.410 1296.860 ;
        RECT 1752.670 1296.800 1752.990 1296.860 ;
        RECT 1511.630 1283.400 1511.950 1283.460 ;
        RECT 1745.770 1283.400 1746.090 1283.460 ;
        RECT 1511.630 1283.260 1746.090 1283.400 ;
        RECT 1511.630 1283.200 1511.950 1283.260 ;
        RECT 1745.770 1283.200 1746.090 1283.260 ;
        RECT 1512.550 1276.260 1512.870 1276.320 ;
        RECT 1738.870 1276.260 1739.190 1276.320 ;
        RECT 1512.550 1276.120 1739.190 1276.260 ;
        RECT 1512.550 1276.060 1512.870 1276.120 ;
        RECT 1738.870 1276.060 1739.190 1276.120 ;
        RECT 1513.930 1262.660 1514.250 1262.720 ;
        RECT 1731.970 1262.660 1732.290 1262.720 ;
        RECT 1513.930 1262.520 1732.290 1262.660 ;
        RECT 1513.930 1262.460 1514.250 1262.520 ;
        RECT 1731.970 1262.460 1732.290 1262.520 ;
        RECT 1513.930 1248.720 1514.250 1248.780 ;
        RECT 1725.070 1248.720 1725.390 1248.780 ;
        RECT 1513.930 1248.580 1725.390 1248.720 ;
        RECT 1513.930 1248.520 1514.250 1248.580 ;
        RECT 1725.070 1248.520 1725.390 1248.580 ;
        RECT 1512.090 1241.920 1512.410 1241.980 ;
        RECT 1718.630 1241.920 1718.950 1241.980 ;
        RECT 1512.090 1241.780 1718.950 1241.920 ;
        RECT 1512.090 1241.720 1512.410 1241.780 ;
        RECT 1718.630 1241.720 1718.950 1241.780 ;
        RECT 1513.470 1227.980 1513.790 1228.040 ;
        RECT 1718.170 1227.980 1718.490 1228.040 ;
        RECT 1513.470 1227.840 1718.490 1227.980 ;
        RECT 1513.470 1227.780 1513.790 1227.840 ;
        RECT 1718.170 1227.780 1718.490 1227.840 ;
        RECT 1512.550 1221.180 1512.870 1221.240 ;
        RECT 1711.270 1221.180 1711.590 1221.240 ;
        RECT 1512.550 1221.040 1711.590 1221.180 ;
        RECT 1512.550 1220.980 1512.870 1221.040 ;
        RECT 1711.270 1220.980 1711.590 1221.040 ;
        RECT 1513.930 1207.240 1514.250 1207.300 ;
        RECT 1704.370 1207.240 1704.690 1207.300 ;
        RECT 1513.930 1207.100 1704.690 1207.240 ;
        RECT 1513.930 1207.040 1514.250 1207.100 ;
        RECT 1704.370 1207.040 1704.690 1207.100 ;
        RECT 1513.930 1193.640 1514.250 1193.700 ;
        RECT 1697.470 1193.640 1697.790 1193.700 ;
        RECT 1513.930 1193.500 1697.790 1193.640 ;
        RECT 1513.930 1193.440 1514.250 1193.500 ;
        RECT 1697.470 1193.440 1697.790 1193.500 ;
        RECT 1512.090 1186.840 1512.410 1186.900 ;
        RECT 1690.570 1186.840 1690.890 1186.900 ;
        RECT 1512.090 1186.700 1690.890 1186.840 ;
        RECT 1512.090 1186.640 1512.410 1186.700 ;
        RECT 1690.570 1186.640 1690.890 1186.700 ;
        RECT 1513.470 1172.900 1513.790 1172.960 ;
        RECT 1684.130 1172.900 1684.450 1172.960 ;
        RECT 1513.470 1172.760 1684.450 1172.900 ;
        RECT 1513.470 1172.700 1513.790 1172.760 ;
        RECT 1684.130 1172.700 1684.450 1172.760 ;
        RECT 1512.550 1166.100 1512.870 1166.160 ;
        RECT 1683.670 1166.100 1683.990 1166.160 ;
        RECT 1512.550 1165.960 1683.990 1166.100 ;
        RECT 1512.550 1165.900 1512.870 1165.960 ;
        RECT 1683.670 1165.900 1683.990 1165.960 ;
        RECT 1513.930 1152.160 1514.250 1152.220 ;
        RECT 1676.770 1152.160 1677.090 1152.220 ;
        RECT 1513.930 1152.020 1677.090 1152.160 ;
        RECT 1513.930 1151.960 1514.250 1152.020 ;
        RECT 1676.770 1151.960 1677.090 1152.020 ;
        RECT 1513.930 1138.560 1514.250 1138.620 ;
        RECT 1669.870 1138.560 1670.190 1138.620 ;
        RECT 1513.930 1138.420 1670.190 1138.560 ;
        RECT 1513.930 1138.360 1514.250 1138.420 ;
        RECT 1669.870 1138.360 1670.190 1138.420 ;
        RECT 1513.930 1131.420 1514.250 1131.480 ;
        RECT 1662.970 1131.420 1663.290 1131.480 ;
        RECT 1513.930 1131.280 1663.290 1131.420 ;
        RECT 1513.930 1131.220 1514.250 1131.280 ;
        RECT 1662.970 1131.220 1663.290 1131.280 ;
        RECT 1513.470 1117.820 1513.790 1117.880 ;
        RECT 1548.890 1117.820 1549.210 1117.880 ;
        RECT 1513.470 1117.680 1549.210 1117.820 ;
        RECT 1513.470 1117.620 1513.790 1117.680 ;
        RECT 1548.890 1117.620 1549.210 1117.680 ;
        RECT 1513.930 1110.680 1514.250 1110.740 ;
        RECT 1649.630 1110.680 1649.950 1110.740 ;
        RECT 1513.930 1110.540 1649.950 1110.680 ;
        RECT 1513.930 1110.480 1514.250 1110.540 ;
        RECT 1649.630 1110.480 1649.950 1110.540 ;
        RECT 1513.930 1097.080 1514.250 1097.140 ;
        RECT 1562.690 1097.080 1563.010 1097.140 ;
        RECT 1513.930 1096.940 1563.010 1097.080 ;
        RECT 1513.930 1096.880 1514.250 1096.940 ;
        RECT 1562.690 1096.880 1563.010 1096.940 ;
        RECT 1513.930 1083.140 1514.250 1083.200 ;
        RECT 1576.490 1083.140 1576.810 1083.200 ;
        RECT 1513.930 1083.000 1576.810 1083.140 ;
        RECT 1513.930 1082.940 1514.250 1083.000 ;
        RECT 1576.490 1082.940 1576.810 1083.000 ;
        RECT 1513.930 1076.340 1514.250 1076.400 ;
        RECT 1635.370 1076.340 1635.690 1076.400 ;
        RECT 1513.930 1076.200 1635.690 1076.340 ;
        RECT 1513.930 1076.140 1514.250 1076.200 ;
        RECT 1635.370 1076.140 1635.690 1076.200 ;
        RECT 1513.010 1062.400 1513.330 1062.460 ;
        RECT 1628.470 1062.400 1628.790 1062.460 ;
        RECT 1513.010 1062.260 1628.790 1062.400 ;
        RECT 1513.010 1062.200 1513.330 1062.260 ;
        RECT 1628.470 1062.200 1628.790 1062.260 ;
        RECT 1513.930 1055.600 1514.250 1055.660 ;
        RECT 1583.390 1055.600 1583.710 1055.660 ;
        RECT 1513.930 1055.460 1583.710 1055.600 ;
        RECT 1513.930 1055.400 1514.250 1055.460 ;
        RECT 1583.390 1055.400 1583.710 1055.460 ;
        RECT 1513.930 1041.660 1514.250 1041.720 ;
        RECT 1614.670 1041.660 1614.990 1041.720 ;
        RECT 1513.930 1041.520 1614.990 1041.660 ;
        RECT 1513.930 1041.460 1514.250 1041.520 ;
        RECT 1614.670 1041.460 1614.990 1041.520 ;
        RECT 1513.930 1028.060 1514.250 1028.120 ;
        RECT 1607.770 1028.060 1608.090 1028.120 ;
        RECT 1513.930 1027.920 1608.090 1028.060 ;
        RECT 1513.930 1027.860 1514.250 1027.920 ;
        RECT 1607.770 1027.860 1608.090 1027.920 ;
      LAYER via ;
        RECT 1318.920 2770.020 1319.180 2770.280 ;
        RECT 1892.540 2770.020 1892.800 2770.280 ;
        RECT 2539.300 2770.020 2539.560 2770.280 ;
        RECT 2566.900 2770.020 2567.160 2770.280 ;
        RECT 668.480 2766.960 668.740 2767.220 ;
        RECT 697.920 2766.960 698.180 2767.220 ;
        RECT 1295.920 2766.960 1296.180 2767.220 ;
        RECT 1318.920 2766.960 1319.180 2767.220 ;
        RECT 1892.540 2766.960 1892.800 2767.220 ;
        RECT 1914.620 2766.960 1914.880 2767.220 ;
        RECT 1946.820 2766.960 1947.080 2767.220 ;
        RECT 2539.300 2766.960 2539.560 2767.220 ;
        RECT 697.000 2751.320 697.260 2751.580 ;
        RECT 1332.260 2751.320 1332.520 2751.580 ;
        RECT 1511.200 2751.320 1511.460 2751.580 ;
        RECT 1945.900 2751.320 1946.160 2751.580 ;
        RECT 2582.080 2751.320 2582.340 2751.580 ;
        RECT 751.740 2732.280 752.000 2732.540 ;
        RECT 938.500 2732.280 938.760 2732.540 ;
        RECT 737.940 2725.480 738.200 2725.740 ;
        RECT 938.500 2725.480 938.760 2725.740 ;
        RECT 724.140 2718.680 724.400 2718.940 ;
        RECT 938.500 2718.680 938.760 2718.940 ;
        RECT 717.240 2711.880 717.500 2712.140 ;
        RECT 938.500 2711.880 938.760 2712.140 ;
        RECT 703.440 2698.280 703.700 2698.540 ;
        RECT 938.960 2698.280 939.220 2698.540 ;
        RECT 696.540 2697.940 696.800 2698.200 ;
        RECT 938.500 2697.940 938.760 2698.200 ;
        RECT 1352.040 2746.220 1352.300 2746.480 ;
        RECT 1511.200 2746.220 1511.460 2746.480 ;
        RECT 1522.240 2725.480 1522.500 2725.740 ;
        RECT 1538.340 2725.480 1538.600 2725.740 ;
        RECT 1521.780 2711.880 1522.040 2712.140 ;
        RECT 1536.040 2711.880 1536.300 2712.140 ;
        RECT 1521.320 2697.940 1521.580 2698.200 ;
        RECT 1538.340 2697.940 1538.600 2698.200 ;
        RECT 1345.600 2421.860 1345.860 2422.120 ;
        RECT 1514.420 2421.860 1514.680 2422.120 ;
        RECT 1514.880 2387.520 1515.140 2387.780 ;
        RECT 1535.580 2387.520 1535.840 2387.780 ;
        RECT 1997.420 2732.280 1997.680 2732.540 ;
        RECT 2187.400 2732.280 2187.660 2732.540 ;
        RECT 1990.520 2725.480 1990.780 2725.740 ;
        RECT 2187.400 2725.480 2187.660 2725.740 ;
        RECT 1976.720 2718.680 1976.980 2718.940 ;
        RECT 2187.400 2718.680 2187.660 2718.940 ;
        RECT 1969.820 2711.880 1970.080 2712.140 ;
        RECT 2187.400 2711.880 2187.660 2712.140 ;
        RECT 1962.920 2698.280 1963.180 2698.540 ;
        RECT 2187.860 2698.280 2188.120 2698.540 ;
        RECT 1956.020 2697.940 1956.280 2698.200 ;
        RECT 2187.400 2697.940 2187.660 2698.200 ;
        RECT 1942.220 2684.000 1942.480 2684.260 ;
        RECT 2187.400 2684.000 2187.660 2684.260 ;
        RECT 2011.220 2401.120 2011.480 2401.380 ;
        RECT 2187.400 2401.120 2187.660 2401.380 ;
        RECT 944.480 2300.820 944.740 2301.080 ;
        RECT 1514.880 2300.820 1515.140 2301.080 ;
        RECT 299.100 2297.420 299.360 2297.680 ;
        RECT 944.480 2297.420 944.740 2297.680 ;
        RECT 1514.880 2297.420 1515.140 2297.680 ;
        RECT 2190.620 2297.420 2190.880 2297.680 ;
        RECT 1514.420 2297.080 1514.680 2297.340 ;
        RECT 1945.900 2297.080 1946.160 2297.340 ;
        RECT 386.500 2290.620 386.760 2290.880 ;
        RECT 431.580 2290.620 431.840 2290.880 ;
        RECT 434.340 2290.620 434.600 2290.880 ;
        RECT 496.900 2290.620 497.160 2290.880 ;
        RECT 526.800 2290.620 527.060 2290.880 ;
        RECT 613.740 2290.620 614.000 2290.880 ;
        RECT 635.360 2290.620 635.620 2290.880 ;
        RECT 710.340 2290.620 710.600 2290.880 ;
        RECT 734.720 2290.620 734.980 2290.880 ;
        RECT 806.940 2290.620 807.200 2290.880 ;
        RECT 952.300 2290.620 952.560 2290.880 ;
        RECT 1000.140 2290.620 1000.400 2290.880 ;
        RECT 1048.900 2290.620 1049.160 2290.880 ;
        RECT 1076.500 2290.620 1076.760 2290.880 ;
        RECT 1086.160 2290.620 1086.420 2290.880 ;
        RECT 1096.740 2290.620 1097.000 2290.880 ;
        RECT 1131.700 2290.620 1131.960 2290.880 ;
        RECT 1676.800 2290.620 1677.060 2290.880 ;
        RECT 1723.720 2290.620 1723.980 2290.880 ;
        RECT 1766.500 2290.620 1766.760 2290.880 ;
        RECT 1770.180 2290.620 1770.440 2290.880 ;
        RECT 2422.000 2290.620 2422.260 2290.880 ;
        RECT 399.840 2290.280 400.100 2290.540 ;
        RECT 445.380 2290.280 445.640 2290.540 ;
        RECT 455.500 2290.280 455.760 2290.540 ;
        RECT 502.880 2290.280 503.140 2290.540 ;
        RECT 538.300 2290.280 538.560 2290.540 ;
        RECT 1117.900 2290.280 1118.160 2290.540 ;
        RECT 1118.360 2290.280 1118.620 2290.540 ;
        RECT 1159.300 2290.280 1159.560 2290.540 ;
        RECT 1645.520 2290.280 1645.780 2290.540 ;
        RECT 1690.140 2290.280 1690.400 2290.540 ;
        RECT 1721.880 2290.280 1722.140 2290.540 ;
        RECT 1759.600 2290.280 1759.860 2290.540 ;
        RECT 1763.740 2290.280 1764.000 2290.540 ;
        RECT 2415.100 2290.280 2415.360 2290.540 ;
        RECT 379.140 2289.940 379.400 2290.200 ;
        RECT 421.000 2289.940 421.260 2290.200 ;
        RECT 467.920 2289.940 468.180 2290.200 ;
        RECT 513.920 2289.940 514.180 2290.200 ;
        RECT 531.400 2289.940 531.660 2290.200 ;
        RECT 1104.100 2289.940 1104.360 2290.200 ;
        RECT 1121.580 2289.940 1121.840 2290.200 ;
        RECT 1166.200 2289.940 1166.460 2290.200 ;
        RECT 1717.740 2289.940 1718.000 2290.200 ;
        RECT 1759.140 2289.940 1759.400 2290.200 ;
        RECT 1769.720 2289.940 1769.980 2290.200 ;
        RECT 2416.020 2289.940 2416.280 2290.200 ;
        RECT 434.340 2289.600 434.600 2289.860 ;
        RECT 478.960 2289.600 479.220 2289.860 ;
        RECT 496.900 2289.600 497.160 2289.860 ;
        RECT 543.820 2289.600 544.080 2289.860 ;
        RECT 613.740 2289.600 614.000 2289.860 ;
        RECT 635.360 2289.600 635.620 2289.860 ;
        RECT 710.340 2289.600 710.600 2289.860 ;
        RECT 734.720 2289.600 734.980 2289.860 ;
        RECT 806.940 2289.600 807.200 2289.860 ;
        RECT 952.300 2289.600 952.560 2289.860 ;
        RECT 1000.140 2289.600 1000.400 2289.860 ;
        RECT 1124.800 2289.600 1125.060 2289.860 ;
        RECT 1129.400 2289.600 1129.660 2289.860 ;
        RECT 1173.100 2289.600 1173.360 2289.860 ;
        RECT 1682.780 2289.600 1683.040 2289.860 ;
        RECT 1729.700 2289.600 1729.960 2289.860 ;
        RECT 1768.340 2289.600 1768.600 2289.860 ;
        RECT 2358.980 2289.600 2359.240 2289.860 ;
        RECT 2402.220 2289.600 2402.480 2289.860 ;
        RECT 406.740 2289.260 407.000 2289.520 ;
        RECT 450.900 2289.260 451.160 2289.520 ;
        RECT 497.360 2289.260 497.620 2289.520 ;
        RECT 1041.080 2289.260 1041.340 2289.520 ;
        RECT 1083.400 2289.260 1083.660 2289.520 ;
        RECT 1085.700 2289.260 1085.960 2289.520 ;
        RECT 1086.160 2289.260 1086.420 2289.520 ;
        RECT 1121.580 2289.260 1121.840 2289.520 ;
        RECT 1656.560 2289.260 1656.820 2289.520 ;
        RECT 1659.320 2289.260 1659.580 2289.520 ;
        RECT 1706.240 2289.260 1706.500 2289.520 ;
        RECT 1752.700 2289.260 1752.960 2289.520 ;
        RECT 1753.160 2289.260 1753.420 2289.520 ;
        RECT 1780.300 2289.260 1780.560 2289.520 ;
        RECT 2301.020 2289.260 2301.280 2289.520 ;
        RECT 2343.800 2289.260 2344.060 2289.520 ;
        RECT 2391.640 2289.260 2391.900 2289.520 ;
        RECT 2435.800 2289.260 2436.060 2289.520 ;
        RECT 392.940 2288.920 393.200 2289.180 ;
        RECT 439.400 2288.920 439.660 2289.180 ;
        RECT 485.860 2288.920 486.120 2289.180 ;
        RECT 489.540 2288.920 489.800 2289.180 ;
        RECT 1065.460 2288.920 1065.720 2289.180 ;
        RECT 1112.840 2288.920 1113.100 2289.180 ;
        RECT 1159.300 2288.920 1159.560 2289.180 ;
        RECT 1695.200 2288.920 1695.460 2289.180 ;
        RECT 1704.400 2288.920 1704.660 2289.180 ;
        RECT 2324.940 2288.920 2325.200 2289.180 ;
        RECT 445.380 2288.580 445.640 2288.840 ;
        RECT 492.760 2288.580 493.020 2288.840 ;
        RECT 538.300 2288.580 538.560 2288.840 ;
        RECT 1070.060 2288.580 1070.320 2288.840 ;
        RECT 1118.360 2288.580 1118.620 2288.840 ;
        RECT 1132.160 2288.580 1132.420 2288.840 ;
        RECT 1135.840 2288.580 1136.100 2288.840 ;
        RECT 1180.000 2288.580 1180.260 2288.840 ;
        RECT 1663.000 2288.580 1663.260 2288.840 ;
        RECT 1665.760 2288.580 1666.020 2288.840 ;
        RECT 1712.680 2288.580 1712.940 2288.840 ;
        RECT 1717.740 2288.580 1718.000 2288.840 ;
        RECT 1746.260 2288.580 1746.520 2288.840 ;
        RECT 365.340 2288.240 365.600 2288.500 ;
        RECT 409.500 2288.240 409.760 2288.500 ;
        RECT 455.500 2288.240 455.760 2288.500 ;
        RECT 489.540 2288.240 489.800 2288.500 ;
        RECT 531.400 2288.240 531.660 2288.500 ;
        RECT 882.840 2288.240 883.100 2288.500 ;
        RECT 1007.500 2288.240 1007.760 2288.500 ;
        RECT 1038.780 2288.240 1039.040 2288.500 ;
        RECT 1048.440 2288.240 1048.700 2288.500 ;
        RECT 1094.440 2288.240 1094.700 2288.500 ;
        RECT 1141.820 2288.240 1142.080 2288.500 ;
        RECT 1186.900 2288.240 1187.160 2288.500 ;
        RECT 1690.140 2288.240 1690.400 2288.500 ;
        RECT 1734.300 2288.240 1734.560 2288.500 ;
        RECT 1748.560 2288.580 1748.820 2288.840 ;
        RECT 2267.440 2288.580 2267.700 2288.840 ;
        RECT 2315.280 2288.580 2315.540 2288.840 ;
        RECT 2356.680 2288.580 2356.940 2288.840 ;
        RECT 2357.600 2288.920 2357.860 2289.180 ;
        RECT 2377.380 2288.920 2377.640 2289.180 ;
        RECT 2422.000 2288.920 2422.260 2289.180 ;
        RECT 2367.260 2288.580 2367.520 2288.840 ;
        RECT 2401.300 2288.580 2401.560 2288.840 ;
        RECT 370.860 2287.900 371.120 2288.160 ;
        RECT 414.100 2287.900 414.360 2288.160 ;
        RECT 462.400 2287.900 462.660 2288.160 ;
        RECT 509.320 2287.900 509.580 2288.160 ;
        RECT 875.940 2287.900 876.200 2288.160 ;
        RECT 1001.060 2287.900 1001.320 2288.160 ;
        RECT 1045.680 2287.900 1045.940 2288.160 ;
        RECT 1052.580 2287.900 1052.840 2288.160 ;
        RECT 1100.880 2287.900 1101.140 2288.160 ;
        RECT 1147.800 2287.900 1148.060 2288.160 ;
        RECT 1193.800 2287.900 1194.060 2288.160 ;
        RECT 1699.340 2287.900 1699.600 2288.160 ;
        RECT 1746.260 2287.900 1746.520 2288.160 ;
        RECT 1753.160 2287.900 1753.420 2288.160 ;
        RECT 1787.200 2288.240 1787.460 2288.500 ;
        RECT 1797.320 2288.240 1797.580 2288.500 ;
        RECT 2290.900 2288.240 2291.160 2288.500 ;
        RECT 2301.940 2288.240 2302.200 2288.500 ;
        RECT 2349.780 2288.240 2350.040 2288.500 ;
        RECT 2397.160 2288.240 2397.420 2288.500 ;
        RECT 2442.700 2288.240 2442.960 2288.500 ;
        RECT 1794.100 2287.900 1794.360 2288.160 ;
        RECT 2266.520 2287.900 2266.780 2288.160 ;
        RECT 2308.840 2287.900 2309.100 2288.160 ;
        RECT 2358.980 2287.900 2359.240 2288.160 ;
        RECT 386.040 2287.560 386.300 2287.820 ;
        RECT 427.440 2287.560 427.700 2287.820 ;
        RECT 473.900 2287.560 474.160 2287.820 ;
        RECT 521.280 2287.560 521.540 2287.820 ;
        RECT 862.140 2287.560 862.400 2287.820 ;
        RECT 993.700 2287.560 993.960 2287.820 ;
        RECT 1062.240 2287.560 1062.500 2287.820 ;
        RECT 1106.860 2287.560 1107.120 2287.820 ;
        RECT 1152.400 2287.560 1152.660 2287.820 ;
        RECT 1670.360 2287.560 1670.620 2287.820 ;
        RECT 1721.880 2287.560 1722.140 2287.820 ;
        RECT 1768.340 2287.560 1768.600 2287.820 ;
        RECT 1775.240 2287.560 1775.500 2287.820 ;
        RECT 1790.420 2287.560 1790.680 2287.820 ;
        RECT 2284.000 2287.560 2284.260 2287.820 ;
        RECT 2325.860 2287.560 2326.120 2287.820 ;
        RECT 2356.220 2287.560 2356.480 2287.820 ;
        RECT 2356.680 2287.560 2356.940 2287.820 ;
        RECT 2361.280 2287.900 2361.540 2288.160 ;
        RECT 2408.200 2287.900 2408.460 2288.160 ;
        RECT 2381.520 2287.560 2381.780 2287.820 ;
        RECT 2384.740 2287.560 2385.000 2287.820 ;
        RECT 2428.900 2287.560 2429.160 2287.820 ;
        RECT 2218.220 2287.220 2218.480 2287.480 ;
        RECT 2297.800 2287.220 2298.060 2287.480 ;
        RECT 2328.620 2287.220 2328.880 2287.480 ;
        RECT 2435.800 2287.220 2436.060 2287.480 ;
        RECT 855.240 2286.880 855.500 2287.140 ;
        RECT 986.800 2286.880 987.060 2287.140 ;
        RECT 1045.220 2286.880 1045.480 2287.140 ;
        RECT 668.940 2286.540 669.200 2286.800 ;
        RECT 979.900 2286.540 980.160 2286.800 ;
        RECT 1010.720 2286.540 1010.980 2286.800 ;
        RECT 1062.240 2286.540 1062.500 2286.800 ;
        RECT 1085.700 2286.880 1085.960 2287.140 ;
        RECT 1124.800 2286.880 1125.060 2287.140 ;
        RECT 1548.920 2286.880 1549.180 2287.140 ;
        RECT 1656.100 2286.880 1656.360 2287.140 ;
        RECT 1704.400 2286.880 1704.660 2287.140 ;
        RECT 1741.200 2286.880 1741.460 2287.140 ;
        RECT 1748.560 2286.880 1748.820 2287.140 ;
        RECT 1776.620 2286.880 1776.880 2287.140 ;
        RECT 2270.200 2286.880 2270.460 2287.140 ;
        RECT 2273.420 2286.880 2273.680 2287.140 ;
        RECT 2324.940 2286.880 2325.200 2287.140 ;
        RECT 2335.520 2286.880 2335.780 2287.140 ;
        RECT 2442.700 2286.880 2442.960 2287.140 ;
        RECT 1088.000 2286.540 1088.260 2286.800 ;
        RECT 1132.160 2286.540 1132.420 2286.800 ;
        RECT 1611.020 2286.540 1611.280 2286.800 ;
        RECT 1656.560 2286.540 1656.820 2286.800 ;
        RECT 1714.520 2286.540 1714.780 2286.800 ;
        RECT 2263.300 2286.540 2263.560 2286.800 ;
        RECT 2321.720 2286.540 2321.980 2286.800 ;
        RECT 2428.900 2286.540 2429.160 2286.800 ;
        RECT 502.880 2286.200 503.140 2286.460 ;
        RECT 1048.900 2286.200 1049.160 2286.460 ;
        RECT 1049.360 2286.200 1049.620 2286.460 ;
        RECT 1096.740 2286.200 1097.000 2286.460 ;
        RECT 1562.720 2286.200 1562.980 2286.460 ;
        RECT 1649.200 2286.200 1649.460 2286.460 ;
        RECT 1749.020 2286.200 1749.280 2286.460 ;
        RECT 2387.500 2286.200 2387.760 2286.460 ;
        RECT 2401.300 2286.200 2401.560 2286.460 ;
        RECT 2415.560 2286.200 2415.820 2286.460 ;
        RECT 509.320 2285.860 509.580 2286.120 ;
        RECT 1062.700 2285.860 1062.960 2286.120 ;
        RECT 1639.540 2285.860 1639.800 2286.120 ;
        RECT 1682.780 2285.860 1683.040 2286.120 ;
        RECT 1755.920 2285.860 1756.180 2286.120 ;
        RECT 2394.400 2285.860 2394.660 2286.120 ;
        RECT 317.040 2285.520 317.300 2285.780 ;
        RECT 365.800 2285.520 366.060 2285.780 ;
        RECT 513.920 2285.520 514.180 2285.780 ;
        RECT 1069.600 2285.520 1069.860 2285.780 ;
        RECT 1076.040 2285.520 1076.300 2285.780 ;
        RECT 1231.520 2285.520 1231.780 2285.780 ;
        RECT 1576.520 2285.520 1576.780 2285.780 ;
        RECT 1642.300 2285.520 1642.560 2285.780 ;
        RECT 1646.440 2285.520 1646.700 2285.780 ;
        RECT 1695.200 2285.520 1695.460 2285.780 ;
        RECT 1762.820 2285.520 1763.080 2285.780 ;
        RECT 2402.680 2285.520 2402.940 2285.780 ;
        RECT 351.540 2285.180 351.800 2285.440 ;
        RECT 386.500 2285.180 386.760 2285.440 ;
        RECT 521.280 2285.180 521.540 2285.440 ;
        RECT 1083.400 2285.180 1083.660 2285.440 ;
        RECT 1617.920 2285.180 1618.180 2285.440 ;
        RECT 1663.000 2285.180 1663.260 2285.440 ;
        RECT 1763.280 2285.180 1763.540 2285.440 ;
        RECT 2408.200 2285.180 2408.460 2285.440 ;
        RECT 344.640 2284.840 344.900 2285.100 ;
        RECT 379.600 2284.840 379.860 2285.100 ;
        RECT 526.800 2284.840 527.060 2285.100 ;
        RECT 1097.200 2284.840 1097.460 2285.100 ;
        RECT 1542.020 2284.840 1542.280 2285.100 ;
        RECT 1587.100 2284.840 1587.360 2285.100 ;
        RECT 1735.220 2284.840 1735.480 2285.100 ;
        RECT 2380.600 2284.840 2380.860 2285.100 ;
        RECT 330.840 2284.500 331.100 2284.760 ;
        RECT 373.620 2284.500 373.880 2284.760 ;
        RECT 1034.180 2284.500 1034.440 2284.760 ;
        RECT 1076.500 2284.500 1076.760 2284.760 ;
        RECT 1624.820 2284.500 1625.080 2284.760 ;
        RECT 1670.360 2284.500 1670.620 2284.760 ;
        RECT 2296.880 2284.500 2297.140 2284.760 ;
        RECT 2340.120 2284.500 2340.380 2284.760 ;
        RECT 2381.520 2284.500 2381.780 2284.760 ;
        RECT 365.340 2284.160 365.600 2284.420 ;
        RECT 393.860 2284.160 394.120 2284.420 ;
        RECT 1027.280 2284.160 1027.540 2284.420 ;
        RECT 1070.060 2284.160 1070.320 2284.420 ;
        RECT 1082.940 2284.160 1083.200 2284.420 ;
        RECT 1224.620 2284.160 1224.880 2284.420 ;
        RECT 1631.720 2284.160 1631.980 2284.420 ;
        RECT 1677.260 2284.160 1677.520 2284.420 ;
        RECT 1783.520 2284.160 1783.780 2284.420 ;
        RECT 2277.100 2284.160 2277.360 2284.420 ;
        RECT 2283.540 2284.160 2283.800 2284.420 ;
        RECT 2325.860 2284.160 2326.120 2284.420 ;
        RECT 310.140 2283.820 310.400 2284.080 ;
        RECT 358.900 2283.820 359.160 2284.080 ;
        RECT 382.820 2283.820 383.080 2284.080 ;
        RECT 393.400 2283.820 393.660 2284.080 ;
        RECT 1017.620 2283.820 1017.880 2284.080 ;
        RECT 1065.460 2283.820 1065.720 2284.080 ;
        RECT 1089.840 2283.820 1090.100 2284.080 ;
        RECT 1210.820 2283.820 1211.080 2284.080 ;
        RECT 1583.420 2283.820 1583.680 2284.080 ;
        RECT 1621.600 2283.820 1621.860 2284.080 ;
        RECT 1652.420 2283.820 1652.680 2284.080 ;
        RECT 1699.340 2283.820 1699.600 2284.080 ;
        RECT 2290.440 2283.820 2290.700 2284.080 ;
        RECT 2333.220 2284.160 2333.480 2284.420 ;
        RECT 2355.760 2284.160 2356.020 2284.420 ;
        RECT 2356.220 2284.160 2356.480 2284.420 ;
        RECT 2374.160 2284.160 2374.420 2284.420 ;
        RECT 2415.100 2284.160 2415.360 2284.420 ;
        RECT 1638.160 2221.940 1638.420 2222.200 ;
        RECT 1638.620 2221.940 1638.880 2222.200 ;
        RECT 1211.740 2216.160 1212.000 2216.420 ;
        RECT 1225.540 2216.160 1225.800 2216.420 ;
        RECT 305.540 2214.460 305.800 2214.720 ;
        RECT 310.140 2214.460 310.400 2214.720 ;
        RECT 339.120 2214.460 339.380 2214.720 ;
        RECT 344.640 2214.460 344.900 2214.720 ;
        RECT 373.160 2214.460 373.420 2214.720 ;
        RECT 382.820 2214.460 383.080 2214.720 ;
        RECT 384.660 2214.460 384.920 2214.720 ;
        RECT 400.300 2214.460 400.560 2214.720 ;
        RECT 407.200 2214.460 407.460 2214.720 ;
        RECT 414.100 2214.460 414.360 2214.720 ;
        RECT 434.340 2214.460 434.600 2214.720 ;
        RECT 439.860 2214.460 440.120 2214.720 ;
        RECT 441.240 2214.460 441.500 2214.720 ;
        RECT 452.280 2214.460 452.540 2214.720 ;
        RECT 461.940 2214.460 462.200 2214.720 ;
        RECT 486.320 2214.460 486.580 2214.720 ;
        RECT 489.540 2214.460 489.800 2214.720 ;
        RECT 542.900 2214.460 543.160 2214.720 ;
        RECT 551.640 2214.460 551.900 2214.720 ;
        RECT 656.520 2214.460 656.780 2214.720 ;
        RECT 690.100 2214.460 690.360 2214.720 ;
        RECT 696.540 2214.460 696.800 2214.720 ;
        RECT 697.000 2214.460 697.260 2214.720 ;
        RECT 941.720 2214.460 941.980 2214.720 ;
        RECT 1030.040 2214.460 1030.300 2214.720 ;
        RECT 1038.780 2214.460 1039.040 2214.720 ;
        RECT 1041.080 2214.460 1041.340 2214.720 ;
        RECT 1045.680 2214.460 1045.940 2214.720 ;
        RECT 1124.340 2214.460 1124.600 2214.720 ;
        RECT 1346.980 2214.460 1347.240 2214.720 ;
        RECT 337.740 2214.120 338.000 2214.380 ;
        RECT 712.640 2214.120 712.900 2214.380 ;
        RECT 713.100 2214.120 713.360 2214.380 ;
        RECT 717.240 2214.120 717.500 2214.380 ;
        RECT 746.680 2214.120 746.940 2214.380 ;
        RECT 751.740 2214.120 752.000 2214.380 ;
        RECT 1131.240 2214.120 1131.500 2214.380 ;
        RECT 1358.480 2214.120 1358.740 2214.380 ;
        RECT 285.300 2213.780 285.560 2214.040 ;
        RECT 769.680 2213.780 769.940 2214.040 ;
        RECT 1007.500 2213.780 1007.760 2214.040 ;
        RECT 1038.320 2213.780 1038.580 2214.040 ;
        RECT 1130.780 2213.780 1131.040 2214.040 ;
        RECT 1369.520 2213.780 1369.780 2214.040 ;
        RECT 285.760 2213.440 286.020 2213.700 ;
        RECT 780.720 2213.440 780.980 2213.700 ;
        RECT 1138.140 2213.440 1138.400 2213.700 ;
        RECT 1381.020 2213.440 1381.280 2213.700 ;
        RECT 283.920 2213.100 284.180 2213.360 ;
        RECT 792.220 2213.100 792.480 2213.360 ;
        RECT 996.000 2213.100 996.260 2213.360 ;
        RECT 1031.420 2213.100 1031.680 2213.360 ;
        RECT 1145.040 2213.100 1145.300 2213.360 ;
        RECT 1392.060 2213.100 1392.320 2213.360 ;
        RECT 286.680 2212.760 286.940 2213.020 ;
        RECT 803.260 2212.760 803.520 2213.020 ;
        RECT 939.420 2212.760 939.680 2213.020 ;
        RECT 944.940 2212.760 945.200 2213.020 ;
        RECT 1013.940 2212.760 1014.200 2213.020 ;
        RECT 1143.200 2212.760 1143.460 2213.020 ;
        RECT 1151.940 2212.760 1152.200 2213.020 ;
        RECT 1403.560 2212.760 1403.820 2213.020 ;
        RECT 344.180 2212.420 344.440 2212.680 ;
        RECT 893.880 2212.420 894.140 2212.680 ;
        RECT 1020.840 2212.420 1021.100 2212.680 ;
        RECT 1154.240 2212.420 1154.500 2212.680 ;
        RECT 1158.840 2212.420 1159.100 2212.680 ;
        RECT 1415.060 2212.420 1415.320 2212.680 ;
        RECT 350.620 2212.080 350.880 2212.340 ;
        RECT 905.380 2212.080 905.640 2212.340 ;
        RECT 1027.740 2212.080 1028.000 2212.340 ;
        RECT 1163.900 2212.080 1164.160 2212.340 ;
        RECT 1165.280 2212.080 1165.540 2212.340 ;
        RECT 1426.100 2212.080 1426.360 2212.340 ;
        RECT 351.080 2211.740 351.340 2212.000 ;
        RECT 916.880 2211.740 917.140 2212.000 ;
        RECT 973.460 2211.740 973.720 2212.000 ;
        RECT 1017.620 2211.740 1017.880 2212.000 ;
        RECT 1034.640 2211.740 1034.900 2212.000 ;
        RECT 1177.240 2211.740 1177.500 2212.000 ;
        RECT 1179.540 2211.740 1179.800 2212.000 ;
        RECT 1460.140 2211.740 1460.400 2212.000 ;
        RECT 358.440 2211.400 358.700 2211.660 ;
        RECT 927.920 2211.400 928.180 2211.660 ;
        RECT 984.500 2211.400 984.760 2211.660 ;
        RECT 1024.520 2211.400 1024.780 2211.660 ;
        RECT 1041.540 2211.400 1041.800 2211.660 ;
        RECT 1188.280 2211.400 1188.540 2211.660 ;
        RECT 1193.340 2211.400 1193.600 2211.660 ;
        RECT 1482.680 2211.400 1482.940 2211.660 ;
        RECT 284.840 2211.060 285.100 2211.320 ;
        RECT 950.460 2211.060 950.720 2211.320 ;
        RECT 961.960 2211.060 962.220 2211.320 ;
        RECT 1010.720 2211.060 1010.980 2211.320 ;
        RECT 1048.440 2211.060 1048.700 2211.320 ;
        RECT 1199.780 2211.060 1200.040 2211.320 ;
        RECT 1210.360 2211.060 1210.620 2211.320 ;
        RECT 1231.060 2211.060 1231.320 2211.320 ;
        RECT 1231.520 2211.060 1231.780 2211.320 ;
        RECT 1256.360 2211.060 1256.620 2211.320 ;
        RECT 1256.820 2211.060 1257.080 2211.320 ;
        RECT 1494.180 2211.060 1494.440 2211.320 ;
        RECT 395.700 2210.720 395.960 2210.980 ;
        RECT 406.740 2210.720 407.000 2210.980 ;
        RECT 448.140 2210.720 448.400 2210.980 ;
        RECT 463.780 2210.720 464.040 2210.980 ;
        RECT 482.640 2210.720 482.900 2210.980 ;
        RECT 531.860 2210.720 532.120 2210.980 ;
        RECT 544.740 2210.720 545.000 2210.980 ;
        RECT 645.020 2210.720 645.280 2210.980 ;
        RECT 679.060 2210.720 679.320 2210.980 ;
        RECT 697.000 2210.720 697.260 2210.980 ;
        RECT 712.640 2210.720 712.900 2210.980 ;
        RECT 758.180 2210.720 758.440 2210.980 ;
        RECT 871.340 2210.720 871.600 2210.980 ;
        RECT 875.940 2210.720 876.200 2210.980 ;
        RECT 1117.440 2210.720 1117.700 2210.980 ;
        RECT 1335.480 2210.720 1335.740 2210.980 ;
        RECT 475.740 2210.380 476.000 2210.640 ;
        RECT 520.360 2210.380 520.620 2210.640 ;
        RECT 530.940 2210.380 531.200 2210.640 ;
        RECT 622.480 2210.380 622.740 2210.640 ;
        RECT 1103.640 2210.380 1103.900 2210.640 ;
        RECT 1312.940 2210.380 1313.200 2210.640 ;
        RECT 468.380 2210.040 468.640 2210.300 ;
        RECT 509.320 2210.040 509.580 2210.300 ;
        RECT 537.840 2210.040 538.100 2210.300 ;
        RECT 633.520 2210.040 633.780 2210.300 ;
        RECT 1110.540 2210.040 1110.800 2210.300 ;
        RECT 1324.440 2210.040 1324.700 2210.300 ;
        RECT 468.840 2209.700 469.100 2209.960 ;
        RECT 497.820 2209.700 498.080 2209.960 ;
        RECT 524.040 2209.700 524.300 2209.960 ;
        RECT 610.980 2209.700 611.240 2209.960 ;
        RECT 848.800 2209.700 849.060 2209.960 ;
        RECT 855.240 2209.700 855.500 2209.960 ;
        RECT 1089.380 2209.700 1089.640 2209.960 ;
        RECT 1290.400 2209.700 1290.660 2209.960 ;
        RECT 509.780 2209.360 510.040 2209.620 ;
        RECT 588.440 2209.360 588.700 2209.620 ;
        RECT 1018.540 2209.360 1018.800 2209.620 ;
        RECT 1045.220 2209.360 1045.480 2209.620 ;
        RECT 1096.740 2209.360 1097.000 2209.620 ;
        RECT 1301.440 2209.360 1301.700 2209.620 ;
        RECT 517.140 2209.020 517.400 2209.280 ;
        RECT 599.480 2209.020 599.740 2209.280 ;
        RECT 1069.140 2209.020 1069.400 2209.280 ;
        RECT 455.040 2208.680 455.300 2208.940 ;
        RECT 475.280 2208.680 475.540 2208.940 ;
        RECT 503.340 2208.680 503.600 2208.940 ;
        RECT 565.900 2208.680 566.160 2208.940 ;
        RECT 1055.340 2208.680 1055.600 2208.940 ;
        RECT 1222.320 2208.680 1222.580 2208.940 ;
        RECT 1224.620 2209.020 1224.880 2209.280 ;
        RECT 1267.860 2209.020 1268.120 2209.280 ;
        RECT 1243.020 2208.680 1243.280 2208.940 ;
        RECT 1243.480 2208.680 1243.740 2208.940 ;
        RECT 1256.820 2208.680 1257.080 2208.940 ;
        RECT 510.240 2208.340 510.500 2208.600 ;
        RECT 576.940 2208.340 577.200 2208.600 ;
        RECT 1062.240 2208.340 1062.500 2208.600 ;
        RECT 1210.360 2208.340 1210.620 2208.600 ;
        RECT 496.440 2208.000 496.700 2208.260 ;
        RECT 554.400 2208.000 554.660 2208.260 ;
        RECT 1054.880 2208.000 1055.140 2208.260 ;
        RECT 1211.280 2208.000 1211.540 2208.260 ;
        RECT 1225.540 2208.000 1225.800 2208.260 ;
        RECT 1278.900 2208.000 1279.160 2208.260 ;
        RECT 1513.960 2186.920 1514.220 2187.180 ;
        RECT 2335.520 2186.920 2335.780 2187.180 ;
        RECT 1513.960 2173.320 1514.220 2173.580 ;
        RECT 1617.460 2173.320 1617.720 2173.580 ;
        RECT 1637.700 2173.320 1637.960 2173.580 ;
        RECT 1638.160 2173.320 1638.420 2173.580 ;
        RECT 1638.620 2173.320 1638.880 2173.580 ;
        RECT 2328.620 2173.320 2328.880 2173.580 ;
        RECT 1617.460 2172.300 1617.720 2172.560 ;
        RECT 1638.620 2172.300 1638.880 2172.560 ;
        RECT 1513.960 2166.180 1514.220 2166.440 ;
        RECT 2321.720 2166.180 2321.980 2166.440 ;
        RECT 1513.960 2152.580 1514.220 2152.840 ;
        RECT 1770.180 2152.580 1770.440 2152.840 ;
        RECT 1513.960 2145.440 1514.220 2145.700 ;
        RECT 1769.720 2145.440 1769.980 2145.700 ;
        RECT 1513.960 2131.840 1514.220 2132.100 ;
        RECT 1763.740 2131.840 1764.000 2132.100 ;
        RECT 1637.700 2118.240 1637.960 2118.500 ;
        RECT 1638.160 2118.240 1638.420 2118.500 ;
        RECT 1513.960 2117.900 1514.220 2118.160 ;
        RECT 1763.280 2117.900 1763.540 2118.160 ;
        RECT 1513.960 2111.100 1514.220 2111.360 ;
        RECT 1762.820 2111.100 1763.080 2111.360 ;
        RECT 1513.960 2097.160 1514.220 2097.420 ;
        RECT 1755.920 2097.160 1756.180 2097.420 ;
        RECT 1513.960 2090.360 1514.220 2090.620 ;
        RECT 1749.020 2090.360 1749.280 2090.620 ;
        RECT 1513.960 2076.760 1514.220 2077.020 ;
        RECT 1735.220 2076.760 1735.480 2077.020 ;
        RECT 1637.700 2069.620 1637.960 2069.880 ;
        RECT 1638.620 2069.620 1638.880 2069.880 ;
        RECT 1513.960 2062.820 1514.220 2063.080 ;
        RECT 2381.060 2062.820 2381.320 2063.080 ;
        RECT 1513.960 2056.020 1514.220 2056.280 ;
        RECT 2373.700 2056.020 2373.960 2056.280 ;
        RECT 1513.960 2042.080 1514.220 2042.340 ;
        RECT 2366.800 2042.080 2367.060 2042.340 ;
        RECT 1513.960 2035.280 1514.220 2035.540 ;
        RECT 2359.900 2035.280 2360.160 2035.540 ;
        RECT 1637.700 2021.680 1637.960 2021.940 ;
        RECT 1638.620 2021.680 1638.880 2021.940 ;
        RECT 1513.500 2021.340 1513.760 2021.600 ;
        RECT 2353.000 2021.340 2353.260 2021.600 ;
        RECT 1513.960 2007.740 1514.220 2008.000 ;
        RECT 2346.100 2007.740 2346.360 2008.000 ;
        RECT 1513.960 2000.600 1514.220 2000.860 ;
        RECT 2339.660 2000.600 2339.920 2000.860 ;
        RECT 1513.960 1987.000 1514.220 1987.260 ;
        RECT 2339.200 1987.000 2339.460 1987.260 ;
        RECT 1512.580 1979.860 1512.840 1980.120 ;
        RECT 2332.300 1979.860 2332.560 1980.120 ;
        RECT 1637.700 1973.060 1637.960 1973.320 ;
        RECT 1638.160 1973.060 1638.420 1973.320 ;
        RECT 1513.500 1966.260 1513.760 1966.520 ;
        RECT 2325.400 1966.260 2325.660 1966.520 ;
        RECT 1513.960 1952.320 1514.220 1952.580 ;
        RECT 2318.500 1952.320 2318.760 1952.580 ;
        RECT 1513.960 1945.520 1514.220 1945.780 ;
        RECT 2311.600 1945.520 2311.860 1945.780 ;
        RECT 1512.580 1931.580 1512.840 1931.840 ;
        RECT 2305.160 1931.580 2305.420 1931.840 ;
        RECT 1638.160 1925.120 1638.420 1925.380 ;
        RECT 1639.080 1925.120 1639.340 1925.380 ;
        RECT 1512.580 1924.780 1512.840 1925.040 ;
        RECT 2304.700 1924.780 2304.960 1925.040 ;
        RECT 1513.960 1910.840 1514.220 1911.100 ;
        RECT 2218.220 1910.840 2218.480 1911.100 ;
        RECT 1513.040 1904.040 1513.300 1904.300 ;
        RECT 1797.320 1904.040 1797.580 1904.300 ;
        RECT 1513.960 1890.440 1514.220 1890.700 ;
        RECT 1790.420 1890.440 1790.680 1890.700 ;
        RECT 1638.160 1883.640 1638.420 1883.900 ;
        RECT 1639.080 1883.640 1639.340 1883.900 ;
        RECT 1513.960 1876.500 1514.220 1876.760 ;
        RECT 1783.520 1876.500 1783.780 1876.760 ;
        RECT 1513.960 1869.700 1514.220 1869.960 ;
        RECT 1776.620 1869.700 1776.880 1869.960 ;
        RECT 1511.660 1855.760 1511.920 1856.020 ;
        RECT 1714.520 1855.760 1714.780 1856.020 ;
        RECT 1513.040 1848.960 1513.300 1849.220 ;
        RECT 2263.760 1848.960 2264.020 1849.220 ;
        RECT 1513.960 1835.020 1514.220 1835.280 ;
        RECT 1652.420 1835.020 1652.680 1835.280 ;
        RECT 1512.580 1821.420 1512.840 1821.680 ;
        RECT 1646.440 1821.420 1646.700 1821.680 ;
        RECT 1512.120 1814.280 1512.380 1814.540 ;
        RECT 1645.520 1814.280 1645.780 1814.540 ;
        RECT 1511.660 1800.680 1511.920 1800.940 ;
        RECT 1640.460 1800.680 1640.720 1800.940 ;
        RECT 1512.580 1793.540 1512.840 1793.800 ;
        RECT 1631.720 1793.540 1631.980 1793.800 ;
        RECT 1513.960 1779.940 1514.220 1780.200 ;
        RECT 1624.820 1779.940 1625.080 1780.200 ;
        RECT 1513.960 1766.000 1514.220 1766.260 ;
        RECT 1617.920 1766.000 1618.180 1766.260 ;
        RECT 1512.120 1759.200 1512.380 1759.460 ;
        RECT 1611.020 1759.200 1611.280 1759.460 ;
        RECT 1513.500 1745.260 1513.760 1745.520 ;
        RECT 2301.940 1745.260 2302.200 1745.520 ;
        RECT 1512.580 1738.460 1512.840 1738.720 ;
        RECT 2301.020 1738.460 2301.280 1738.720 ;
        RECT 1513.960 1724.860 1514.220 1725.120 ;
        RECT 2294.120 1724.860 2294.380 1725.120 ;
        RECT 1513.960 1710.920 1514.220 1711.180 ;
        RECT 2287.220 1710.920 2287.480 1711.180 ;
        RECT 1512.120 1704.120 1512.380 1704.380 ;
        RECT 2280.320 1704.120 2280.580 1704.380 ;
        RECT 1513.500 1690.180 1513.760 1690.440 ;
        RECT 2273.420 1690.180 2273.680 1690.440 ;
        RECT 1512.580 1683.380 1512.840 1683.640 ;
        RECT 2267.440 1683.380 2267.700 1683.640 ;
        RECT 1513.960 1669.440 1514.220 1669.700 ;
        RECT 2266.520 1669.440 2266.780 1669.700 ;
        RECT 1512.580 1655.500 1512.840 1655.760 ;
        RECT 1529.140 1655.500 1529.400 1655.760 ;
        RECT 1511.660 1647.000 1511.920 1647.260 ;
        RECT 1522.240 1647.000 1522.500 1647.260 ;
        RECT 1512.580 1634.420 1512.840 1634.680 ;
        RECT 1528.680 1634.420 1528.940 1634.680 ;
        RECT 1511.660 1622.180 1511.920 1622.440 ;
        RECT 1521.780 1622.180 1522.040 1622.440 ;
        RECT 1511.660 1613.340 1511.920 1613.600 ;
        RECT 1528.220 1613.340 1528.480 1613.600 ;
        RECT 1511.660 1600.420 1511.920 1600.680 ;
        RECT 1521.320 1600.420 1521.580 1600.680 ;
        RECT 1513.500 1591.580 1513.760 1591.840 ;
        RECT 1535.120 1591.580 1535.380 1591.840 ;
        RECT 1513.960 1579.680 1514.220 1579.940 ;
        RECT 1580.200 1579.680 1580.460 1579.940 ;
        RECT 1513.960 1572.880 1514.220 1573.140 ;
        RECT 1997.420 1572.880 1997.680 1573.140 ;
        RECT 1513.500 1558.940 1513.760 1559.200 ;
        RECT 1990.520 1558.940 1990.780 1559.200 ;
        RECT 1513.960 1545.340 1514.220 1545.600 ;
        RECT 1976.720 1545.340 1976.980 1545.600 ;
        RECT 1513.960 1538.540 1514.220 1538.800 ;
        RECT 1969.820 1538.540 1970.080 1538.800 ;
        RECT 1513.960 1524.600 1514.220 1524.860 ;
        RECT 1962.920 1524.600 1963.180 1524.860 ;
        RECT 1513.960 1517.800 1514.220 1518.060 ;
        RECT 1956.020 1517.800 1956.280 1518.060 ;
        RECT 1513.500 1503.860 1513.760 1504.120 ;
        RECT 1942.220 1503.860 1942.480 1504.120 ;
        RECT 1513.960 1490.260 1514.220 1490.520 ;
        RECT 2228.800 1490.260 2229.060 1490.520 ;
        RECT 1513.040 1479.380 1513.300 1479.640 ;
        RECT 1529.600 1479.380 1529.860 1479.640 ;
        RECT 1513.960 1469.520 1514.220 1469.780 ;
        RECT 2011.220 1469.520 2011.480 1469.780 ;
        RECT 1512.580 1462.380 1512.840 1462.640 ;
        RECT 1601.360 1462.380 1601.620 1462.640 ;
        RECT 1513.500 1448.780 1513.760 1449.040 ;
        RECT 1600.900 1448.780 1601.160 1449.040 ;
        RECT 1513.960 1434.840 1514.220 1435.100 ;
        RECT 1594.000 1434.840 1594.260 1435.100 ;
        RECT 1513.500 1426.340 1513.760 1426.600 ;
        RECT 1542.020 1426.340 1542.280 1426.600 ;
        RECT 1512.580 1414.100 1512.840 1414.360 ;
        RECT 2252.720 1414.100 2252.980 1414.360 ;
        RECT 1512.580 1407.300 1512.840 1407.560 ;
        RECT 2245.820 1407.300 2246.080 1407.560 ;
        RECT 1511.660 1393.360 1511.920 1393.620 ;
        RECT 2238.920 1393.360 2239.180 1393.620 ;
        RECT 1513.040 1386.560 1513.300 1386.820 ;
        RECT 2232.020 1386.560 2232.280 1386.820 ;
        RECT 1513.960 1372.960 1514.220 1373.220 ;
        RECT 1794.100 1372.960 1794.360 1373.220 ;
        RECT 1512.580 1359.020 1512.840 1359.280 ;
        RECT 1787.200 1359.020 1787.460 1359.280 ;
        RECT 1512.580 1352.220 1512.840 1352.480 ;
        RECT 1780.300 1352.220 1780.560 1352.480 ;
        RECT 1511.660 1338.280 1511.920 1338.540 ;
        RECT 1773.400 1338.280 1773.660 1338.540 ;
        RECT 1513.040 1331.480 1513.300 1331.740 ;
        RECT 1766.500 1331.480 1766.760 1331.740 ;
        RECT 1513.960 1317.540 1514.220 1317.800 ;
        RECT 1760.060 1317.540 1760.320 1317.800 ;
        RECT 1512.580 1303.940 1512.840 1304.200 ;
        RECT 1759.600 1303.940 1759.860 1304.200 ;
        RECT 1512.120 1296.800 1512.380 1297.060 ;
        RECT 1752.700 1296.800 1752.960 1297.060 ;
        RECT 1511.660 1283.200 1511.920 1283.460 ;
        RECT 1745.800 1283.200 1746.060 1283.460 ;
        RECT 1512.580 1276.060 1512.840 1276.320 ;
        RECT 1738.900 1276.060 1739.160 1276.320 ;
        RECT 1513.960 1262.460 1514.220 1262.720 ;
        RECT 1732.000 1262.460 1732.260 1262.720 ;
        RECT 1513.960 1248.520 1514.220 1248.780 ;
        RECT 1725.100 1248.520 1725.360 1248.780 ;
        RECT 1512.120 1241.720 1512.380 1241.980 ;
        RECT 1718.660 1241.720 1718.920 1241.980 ;
        RECT 1513.500 1227.780 1513.760 1228.040 ;
        RECT 1718.200 1227.780 1718.460 1228.040 ;
        RECT 1512.580 1220.980 1512.840 1221.240 ;
        RECT 1711.300 1220.980 1711.560 1221.240 ;
        RECT 1513.960 1207.040 1514.220 1207.300 ;
        RECT 1704.400 1207.040 1704.660 1207.300 ;
        RECT 1513.960 1193.440 1514.220 1193.700 ;
        RECT 1697.500 1193.440 1697.760 1193.700 ;
        RECT 1512.120 1186.640 1512.380 1186.900 ;
        RECT 1690.600 1186.640 1690.860 1186.900 ;
        RECT 1513.500 1172.700 1513.760 1172.960 ;
        RECT 1684.160 1172.700 1684.420 1172.960 ;
        RECT 1512.580 1165.900 1512.840 1166.160 ;
        RECT 1683.700 1165.900 1683.960 1166.160 ;
        RECT 1513.960 1151.960 1514.220 1152.220 ;
        RECT 1676.800 1151.960 1677.060 1152.220 ;
        RECT 1513.960 1138.360 1514.220 1138.620 ;
        RECT 1669.900 1138.360 1670.160 1138.620 ;
        RECT 1513.960 1131.220 1514.220 1131.480 ;
        RECT 1663.000 1131.220 1663.260 1131.480 ;
        RECT 1513.500 1117.620 1513.760 1117.880 ;
        RECT 1548.920 1117.620 1549.180 1117.880 ;
        RECT 1513.960 1110.480 1514.220 1110.740 ;
        RECT 1649.660 1110.480 1649.920 1110.740 ;
        RECT 1513.960 1096.880 1514.220 1097.140 ;
        RECT 1562.720 1096.880 1562.980 1097.140 ;
        RECT 1513.960 1082.940 1514.220 1083.200 ;
        RECT 1576.520 1082.940 1576.780 1083.200 ;
        RECT 1513.960 1076.140 1514.220 1076.400 ;
        RECT 1635.400 1076.140 1635.660 1076.400 ;
        RECT 1513.040 1062.200 1513.300 1062.460 ;
        RECT 1628.500 1062.200 1628.760 1062.460 ;
        RECT 1513.960 1055.400 1514.220 1055.660 ;
        RECT 1583.420 1055.400 1583.680 1055.660 ;
        RECT 1513.960 1041.460 1514.220 1041.720 ;
        RECT 1614.700 1041.460 1614.960 1041.720 ;
        RECT 1513.960 1027.860 1514.220 1028.120 ;
        RECT 1607.800 1027.860 1608.060 1028.120 ;
      LAYER met2 ;
        RECT 1318.920 2769.990 1319.180 2770.310 ;
        RECT 1892.540 2769.990 1892.800 2770.310 ;
        RECT 2539.300 2769.990 2539.560 2770.310 ;
        RECT 2566.900 2769.990 2567.160 2770.310 ;
        RECT 1318.980 2767.445 1319.120 2769.990 ;
        RECT 1892.600 2767.445 1892.740 2769.990 ;
        RECT 2539.360 2767.445 2539.500 2769.990 ;
        RECT 2566.960 2767.445 2567.100 2769.990 ;
        RECT 668.470 2767.075 668.750 2767.445 ;
        RECT 668.480 2766.930 668.740 2767.075 ;
        RECT 697.920 2766.930 698.180 2767.250 ;
        RECT 1295.910 2767.075 1296.190 2767.445 ;
        RECT 1318.910 2767.075 1319.190 2767.445 ;
        RECT 1892.530 2767.075 1892.810 2767.445 ;
        RECT 1914.610 2767.075 1914.890 2767.445 ;
        RECT 1295.920 2766.930 1296.180 2767.075 ;
        RECT 1318.920 2766.930 1319.180 2767.075 ;
        RECT 1892.540 2766.930 1892.800 2767.075 ;
        RECT 1914.620 2766.930 1914.880 2767.075 ;
        RECT 1946.820 2766.930 1947.080 2767.250 ;
        RECT 2539.290 2767.075 2539.570 2767.445 ;
        RECT 2566.890 2767.075 2567.170 2767.445 ;
        RECT 2539.300 2766.930 2539.560 2767.075 ;
        RECT 697.000 2751.290 697.260 2751.610 ;
        RECT 287.590 2732.395 287.870 2732.765 ;
        RECT 287.130 2725.595 287.410 2725.965 ;
        RECT 284.370 2718.795 284.650 2719.165 ;
        RECT 283.910 2701.795 284.190 2702.165 ;
        RECT 283.980 2213.390 284.120 2701.795 ;
        RECT 283.920 2213.070 284.180 2213.390 ;
        RECT 284.440 2212.565 284.580 2718.795 ;
        RECT 286.670 2711.995 286.950 2712.365 ;
        RECT 285.750 2697.715 286.030 2698.085 ;
        RECT 285.290 2687.515 285.570 2687.885 ;
        RECT 284.830 2401.235 285.110 2401.605 ;
        RECT 284.370 2212.195 284.650 2212.565 ;
        RECT 284.900 2211.350 285.040 2401.235 ;
        RECT 285.360 2214.070 285.500 2687.515 ;
        RECT 285.300 2213.750 285.560 2214.070 ;
        RECT 285.820 2213.730 285.960 2697.715 ;
        RECT 285.760 2213.410 286.020 2213.730 ;
        RECT 286.740 2213.050 286.880 2711.995 ;
        RECT 286.680 2212.730 286.940 2213.050 ;
        RECT 287.200 2211.885 287.340 2725.595 ;
        RECT 287.130 2211.515 287.410 2211.885 ;
        RECT 284.840 2211.030 285.100 2211.350 ;
        RECT 287.660 2211.205 287.800 2732.395 ;
        RECT 299.090 2392.590 299.370 2392.960 ;
        RECT 299.160 2297.710 299.300 2392.590 ;
      LAYER met2 ;
        RECT 305.000 2305.000 681.480 2751.235 ;
      LAYER met2 ;
        RECT 697.060 2749.765 697.200 2751.290 ;
        RECT 696.990 2749.395 697.270 2749.765 ;
        RECT 697.980 2748.970 698.120 2766.930 ;
        RECT 1318.980 2766.775 1319.120 2766.930 ;
        RECT 1892.600 2766.775 1892.740 2766.930 ;
        RECT 1332.260 2751.290 1332.520 2751.610 ;
        RECT 1511.200 2751.290 1511.460 2751.610 ;
        RECT 1945.900 2751.290 1946.160 2751.610 ;
        RECT 697.060 2748.830 698.120 2748.970 ;
        RECT 696.540 2697.910 696.800 2698.230 ;
        RECT 299.100 2297.390 299.360 2297.710 ;
        RECT 386.490 2297.195 386.770 2297.565 ;
        RECT 386.560 2290.910 386.700 2297.195 ;
        RECT 526.860 2290.910 527.000 2291.065 ;
        RECT 370.850 2290.395 371.130 2290.765 ;
        RECT 379.130 2290.395 379.410 2290.765 ;
        RECT 386.500 2290.590 386.760 2290.910 ;
        RECT 431.580 2290.765 431.840 2290.910 ;
        RECT 399.830 2290.395 400.110 2290.765 ;
        RECT 409.490 2290.395 409.770 2290.765 ;
        RECT 414.090 2290.395 414.370 2290.765 ;
        RECT 420.990 2290.395 421.270 2290.765 ;
        RECT 427.430 2290.395 427.710 2290.765 ;
        RECT 431.570 2290.395 431.850 2290.765 ;
        RECT 434.340 2290.590 434.600 2290.910 ;
        RECT 365.330 2288.355 365.610 2288.725 ;
        RECT 365.340 2288.210 365.600 2288.355 ;
        RECT 370.920 2288.190 371.060 2290.395 ;
        RECT 379.200 2290.230 379.340 2290.395 ;
        RECT 399.840 2290.250 400.100 2290.395 ;
        RECT 379.140 2289.910 379.400 2290.230 ;
        RECT 406.730 2289.715 407.010 2290.085 ;
        RECT 406.800 2289.550 406.940 2289.715 ;
        RECT 392.930 2289.035 393.210 2289.405 ;
        RECT 406.740 2289.230 407.000 2289.550 ;
        RECT 392.940 2288.890 393.200 2289.035 ;
        RECT 409.560 2288.530 409.700 2290.395 ;
        RECT 409.500 2288.210 409.760 2288.530 ;
        RECT 414.160 2288.190 414.300 2290.395 ;
        RECT 421.060 2290.230 421.200 2290.395 ;
        RECT 421.000 2289.910 421.260 2290.230 ;
        RECT 370.860 2287.870 371.120 2288.190 ;
        RECT 386.030 2287.675 386.310 2288.045 ;
        RECT 414.100 2287.870 414.360 2288.190 ;
        RECT 427.500 2287.850 427.640 2290.395 ;
        RECT 434.400 2289.890 434.540 2290.590 ;
        RECT 439.390 2290.395 439.670 2290.765 ;
        RECT 445.370 2290.395 445.650 2290.765 ;
        RECT 450.890 2290.395 451.170 2290.765 ;
        RECT 455.490 2290.395 455.770 2290.765 ;
        RECT 462.390 2290.395 462.670 2290.765 ;
        RECT 467.910 2290.395 468.190 2290.765 ;
        RECT 473.890 2290.395 474.170 2290.765 ;
        RECT 478.950 2290.395 479.230 2290.765 ;
        RECT 485.850 2290.395 486.130 2290.765 ;
        RECT 492.750 2290.395 493.030 2290.765 ;
        RECT 496.900 2290.590 497.160 2290.910 ;
        RECT 526.800 2290.765 527.060 2290.910 ;
        RECT 434.340 2289.570 434.600 2289.890 ;
        RECT 439.460 2289.210 439.600 2290.395 ;
        RECT 445.380 2290.250 445.640 2290.395 ;
        RECT 439.400 2288.890 439.660 2289.210 ;
        RECT 445.440 2288.870 445.580 2290.250 ;
        RECT 450.960 2289.550 451.100 2290.395 ;
        RECT 455.500 2290.250 455.760 2290.395 ;
        RECT 450.900 2289.230 451.160 2289.550 ;
        RECT 445.380 2288.550 445.640 2288.870 ;
        RECT 455.560 2288.530 455.700 2290.250 ;
        RECT 455.500 2288.210 455.760 2288.530 ;
        RECT 462.460 2288.190 462.600 2290.395 ;
        RECT 467.980 2290.230 468.120 2290.395 ;
        RECT 467.920 2289.910 468.180 2290.230 ;
        RECT 462.400 2287.870 462.660 2288.190 ;
        RECT 473.960 2287.850 474.100 2290.395 ;
        RECT 479.020 2289.890 479.160 2290.395 ;
        RECT 478.960 2289.570 479.220 2289.890 ;
        RECT 485.920 2289.210 486.060 2290.395 ;
        RECT 485.860 2288.890 486.120 2289.210 ;
        RECT 489.540 2288.890 489.800 2289.210 ;
        RECT 489.600 2288.530 489.740 2288.890 ;
        RECT 492.820 2288.870 492.960 2290.395 ;
        RECT 496.960 2289.890 497.100 2290.590 ;
        RECT 497.350 2290.395 497.630 2290.765 ;
        RECT 496.900 2289.570 497.160 2289.890 ;
        RECT 497.420 2289.550 497.560 2290.395 ;
        RECT 502.880 2290.250 503.140 2290.570 ;
        RECT 503.330 2290.395 503.610 2290.765 ;
        RECT 509.770 2290.395 510.050 2290.765 ;
        RECT 513.910 2290.395 514.190 2290.765 ;
        RECT 517.130 2290.395 517.410 2290.765 ;
        RECT 521.270 2290.395 521.550 2290.765 ;
        RECT 524.030 2290.395 524.310 2290.765 ;
        RECT 526.790 2290.395 527.070 2290.765 ;
        RECT 530.930 2290.395 531.210 2290.765 ;
        RECT 537.830 2290.395 538.110 2290.765 ;
        RECT 502.940 2290.085 503.080 2290.250 ;
        RECT 502.870 2289.715 503.150 2290.085 ;
        RECT 497.360 2289.230 497.620 2289.550 ;
        RECT 492.760 2288.550 493.020 2288.870 ;
        RECT 489.540 2288.210 489.800 2288.530 ;
        RECT 386.040 2287.530 386.300 2287.675 ;
        RECT 427.440 2287.530 427.700 2287.850 ;
        RECT 473.900 2287.530 474.160 2287.850 ;
        RECT 365.790 2286.995 366.070 2287.365 ;
        RECT 379.590 2286.995 379.870 2287.365 ;
        RECT 317.040 2285.490 317.300 2285.810 ;
        RECT 358.890 2285.635 359.170 2286.005 ;
        RECT 365.860 2285.810 366.000 2286.995 ;
        RECT 310.140 2283.790 310.400 2284.110 ;
        RECT 310.200 2214.750 310.340 2283.790 ;
        RECT 305.540 2214.430 305.800 2214.750 ;
        RECT 310.140 2214.430 310.400 2214.750 ;
        RECT 287.590 2210.835 287.870 2211.205 ;
        RECT 305.600 2200.000 305.740 2214.430 ;
        RECT 305.600 2199.460 305.890 2200.000 ;
        RECT 305.610 2196.000 305.890 2199.460 ;
        RECT 316.650 2199.530 316.930 2200.000 ;
        RECT 317.100 2199.530 317.240 2285.490 ;
        RECT 344.640 2284.810 344.900 2285.130 ;
        RECT 351.070 2284.955 351.350 2285.325 ;
        RECT 351.540 2285.150 351.800 2285.470 ;
        RECT 330.840 2284.470 331.100 2284.790 ;
        RECT 316.650 2199.390 317.240 2199.530 ;
        RECT 316.650 2196.000 316.930 2199.390 ;
        RECT 328.150 2198.850 328.430 2200.000 ;
        RECT 330.900 2198.850 331.040 2284.470 ;
        RECT 337.730 2284.275 338.010 2284.645 ;
        RECT 344.170 2284.275 344.450 2284.645 ;
        RECT 337.800 2214.410 337.940 2284.275 ;
        RECT 339.120 2214.430 339.380 2214.750 ;
        RECT 337.740 2214.090 338.000 2214.410 ;
        RECT 339.180 2200.000 339.320 2214.430 ;
        RECT 344.240 2212.710 344.380 2284.275 ;
        RECT 344.700 2214.750 344.840 2284.810 ;
        RECT 350.610 2284.275 350.890 2284.645 ;
        RECT 344.640 2214.430 344.900 2214.750 ;
        RECT 344.180 2212.390 344.440 2212.710 ;
        RECT 350.680 2212.370 350.820 2284.275 ;
        RECT 350.620 2212.050 350.880 2212.370 ;
        RECT 351.140 2212.030 351.280 2284.955 ;
        RECT 351.080 2211.710 351.340 2212.030 ;
        RECT 339.180 2199.460 339.470 2200.000 ;
        RECT 328.150 2198.710 331.040 2198.850 ;
        RECT 328.150 2196.000 328.430 2198.710 ;
        RECT 339.190 2196.000 339.470 2199.460 ;
        RECT 350.690 2199.530 350.970 2200.000 ;
        RECT 351.600 2199.530 351.740 2285.150 ;
        RECT 358.430 2284.275 358.710 2284.645 ;
        RECT 358.500 2211.690 358.640 2284.275 ;
        RECT 358.960 2284.110 359.100 2285.635 ;
        RECT 365.800 2285.490 366.060 2285.810 ;
        RECT 373.610 2284.955 373.890 2285.325 ;
        RECT 379.660 2285.130 379.800 2286.995 ;
        RECT 502.940 2286.490 503.080 2289.715 ;
        RECT 502.880 2286.170 503.140 2286.490 ;
        RECT 386.490 2285.635 386.770 2286.005 ;
        RECT 475.730 2285.635 476.010 2286.005 ;
        RECT 496.430 2285.635 496.710 2286.005 ;
        RECT 386.560 2285.470 386.700 2285.635 ;
        RECT 386.500 2285.150 386.760 2285.470 ;
        RECT 373.680 2284.790 373.820 2284.955 ;
        RECT 379.600 2284.810 379.860 2285.130 ;
        RECT 393.850 2284.955 394.130 2285.325 ;
        RECT 468.830 2284.955 469.110 2285.325 ;
        RECT 373.620 2284.470 373.880 2284.790 ;
        RECT 365.340 2284.130 365.600 2284.450 ;
        RECT 393.390 2284.275 393.670 2284.645 ;
        RECT 393.920 2284.450 394.060 2284.955 ;
        RECT 358.900 2283.790 359.160 2284.110 ;
        RECT 358.440 2211.370 358.700 2211.690 ;
        RECT 350.690 2199.390 351.740 2199.530 ;
        RECT 350.690 2196.000 350.970 2199.390 ;
        RECT 362.190 2198.850 362.470 2200.000 ;
        RECT 365.400 2198.850 365.540 2284.130 ;
        RECT 393.460 2284.110 393.600 2284.275 ;
        RECT 393.860 2284.130 394.120 2284.450 ;
        RECT 400.290 2284.275 400.570 2284.645 ;
        RECT 407.190 2284.275 407.470 2284.645 ;
        RECT 414.090 2284.275 414.370 2284.645 ;
        RECT 420.990 2284.275 421.270 2284.645 ;
        RECT 431.110 2284.275 431.390 2284.645 ;
        RECT 434.330 2284.275 434.610 2284.645 ;
        RECT 441.230 2284.275 441.510 2284.645 ;
        RECT 448.130 2284.275 448.410 2284.645 ;
        RECT 455.030 2284.275 455.310 2284.645 ;
        RECT 461.930 2284.275 462.210 2284.645 ;
        RECT 468.370 2284.275 468.650 2284.645 ;
        RECT 382.820 2283.790 383.080 2284.110 ;
        RECT 393.400 2283.790 393.660 2284.110 ;
        RECT 382.880 2214.750 383.020 2283.790 ;
        RECT 400.360 2214.750 400.500 2284.275 ;
        RECT 407.260 2215.170 407.400 2284.275 ;
        RECT 406.800 2215.030 407.400 2215.170 ;
        RECT 373.160 2214.430 373.420 2214.750 ;
        RECT 382.820 2214.430 383.080 2214.750 ;
        RECT 384.660 2214.430 384.920 2214.750 ;
        RECT 400.300 2214.430 400.560 2214.750 ;
        RECT 373.220 2200.000 373.360 2214.430 ;
        RECT 384.720 2200.000 384.860 2214.430 ;
        RECT 406.800 2211.010 406.940 2215.030 ;
        RECT 414.160 2214.750 414.300 2284.275 ;
        RECT 407.200 2214.430 407.460 2214.750 ;
        RECT 414.100 2214.430 414.360 2214.750 ;
        RECT 395.700 2210.690 395.960 2211.010 ;
        RECT 406.740 2210.690 407.000 2211.010 ;
        RECT 395.760 2200.000 395.900 2210.690 ;
        RECT 407.260 2200.000 407.400 2214.430 ;
        RECT 421.060 2208.370 421.200 2284.275 ;
        RECT 420.600 2208.230 421.200 2208.370 ;
        RECT 373.220 2199.460 373.510 2200.000 ;
        RECT 384.720 2199.460 385.010 2200.000 ;
        RECT 395.760 2199.460 396.050 2200.000 ;
        RECT 407.260 2199.460 407.550 2200.000 ;
        RECT 362.190 2198.710 365.540 2198.850 ;
        RECT 362.190 2196.000 362.470 2198.710 ;
        RECT 373.230 2196.000 373.510 2199.460 ;
        RECT 384.730 2196.000 385.010 2199.460 ;
        RECT 395.770 2196.000 396.050 2199.460 ;
        RECT 407.270 2196.000 407.550 2199.460 ;
        RECT 418.770 2199.530 419.050 2200.000 ;
        RECT 420.600 2199.530 420.740 2208.230 ;
        RECT 418.770 2199.390 420.740 2199.530 ;
        RECT 429.810 2199.530 430.090 2200.000 ;
        RECT 431.180 2199.530 431.320 2284.275 ;
        RECT 434.400 2214.750 434.540 2284.275 ;
        RECT 441.300 2214.750 441.440 2284.275 ;
        RECT 434.340 2214.430 434.600 2214.750 ;
        RECT 439.860 2214.430 440.120 2214.750 ;
        RECT 441.240 2214.430 441.500 2214.750 ;
        RECT 429.810 2199.390 431.320 2199.530 ;
        RECT 439.920 2199.530 440.060 2214.430 ;
        RECT 448.200 2211.010 448.340 2284.275 ;
        RECT 452.280 2214.430 452.540 2214.750 ;
        RECT 448.140 2210.690 448.400 2211.010 ;
        RECT 452.340 2200.000 452.480 2214.430 ;
        RECT 455.100 2208.970 455.240 2284.275 ;
        RECT 462.000 2214.750 462.140 2284.275 ;
        RECT 461.940 2214.430 462.200 2214.750 ;
        RECT 463.780 2210.690 464.040 2211.010 ;
        RECT 455.040 2208.650 455.300 2208.970 ;
        RECT 463.840 2200.000 463.980 2210.690 ;
        RECT 468.440 2210.330 468.580 2284.275 ;
        RECT 468.380 2210.010 468.640 2210.330 ;
        RECT 468.900 2209.990 469.040 2284.955 ;
        RECT 475.800 2210.670 475.940 2285.635 ;
        RECT 482.630 2284.275 482.910 2284.645 ;
        RECT 489.530 2284.275 489.810 2284.645 ;
        RECT 482.700 2211.010 482.840 2284.275 ;
        RECT 489.600 2214.750 489.740 2284.275 ;
        RECT 486.320 2214.430 486.580 2214.750 ;
        RECT 489.540 2214.430 489.800 2214.750 ;
        RECT 482.640 2210.690 482.900 2211.010 ;
        RECT 475.740 2210.350 476.000 2210.670 ;
        RECT 468.840 2209.670 469.100 2209.990 ;
        RECT 475.280 2208.650 475.540 2208.970 ;
        RECT 475.340 2200.000 475.480 2208.650 ;
        RECT 486.380 2200.000 486.520 2214.430 ;
        RECT 496.500 2208.290 496.640 2285.635 ;
        RECT 497.820 2209.670 498.080 2209.990 ;
        RECT 496.440 2207.970 496.700 2208.290 ;
        RECT 497.880 2200.000 498.020 2209.670 ;
        RECT 503.400 2208.970 503.540 2290.395 ;
        RECT 509.310 2289.035 509.590 2289.405 ;
        RECT 509.380 2288.190 509.520 2289.035 ;
        RECT 509.320 2287.870 509.580 2288.190 ;
        RECT 509.380 2286.150 509.520 2287.870 ;
        RECT 509.320 2285.830 509.580 2286.150 ;
        RECT 509.320 2210.010 509.580 2210.330 ;
        RECT 503.340 2208.650 503.600 2208.970 ;
        RECT 509.380 2200.000 509.520 2210.010 ;
        RECT 509.840 2209.650 509.980 2290.395 ;
        RECT 513.980 2290.230 514.120 2290.395 ;
        RECT 510.230 2289.715 510.510 2290.085 ;
        RECT 513.920 2289.910 514.180 2290.230 ;
        RECT 509.780 2209.330 510.040 2209.650 ;
        RECT 510.300 2208.630 510.440 2289.715 ;
        RECT 513.980 2285.810 514.120 2289.910 ;
        RECT 513.920 2285.490 514.180 2285.810 ;
        RECT 517.200 2209.310 517.340 2290.395 ;
        RECT 521.340 2287.850 521.480 2290.395 ;
        RECT 521.280 2287.530 521.540 2287.850 ;
        RECT 521.340 2285.470 521.480 2287.530 ;
        RECT 521.280 2285.150 521.540 2285.470 ;
        RECT 520.360 2210.350 520.620 2210.670 ;
        RECT 517.140 2208.990 517.400 2209.310 ;
        RECT 510.240 2208.310 510.500 2208.630 ;
        RECT 520.420 2200.000 520.560 2210.350 ;
        RECT 524.100 2209.990 524.240 2290.395 ;
        RECT 526.860 2285.130 527.000 2290.395 ;
        RECT 526.800 2284.810 527.060 2285.130 ;
        RECT 531.000 2210.670 531.140 2290.395 ;
        RECT 531.400 2290.085 531.660 2290.230 ;
        RECT 531.390 2289.715 531.670 2290.085 ;
        RECT 531.460 2288.530 531.600 2289.715 ;
        RECT 531.400 2288.210 531.660 2288.530 ;
        RECT 531.860 2210.690 532.120 2211.010 ;
        RECT 530.940 2210.350 531.200 2210.670 ;
        RECT 524.040 2209.670 524.300 2209.990 ;
        RECT 531.920 2200.000 532.060 2210.690 ;
        RECT 537.900 2210.330 538.040 2290.395 ;
        RECT 538.300 2290.250 538.560 2290.570 ;
        RECT 543.810 2290.395 544.090 2290.765 ;
        RECT 551.630 2290.395 551.910 2290.765 ;
        RECT 613.740 2290.590 614.000 2290.910 ;
        RECT 635.360 2290.590 635.620 2290.910 ;
        RECT 538.360 2290.085 538.500 2290.250 ;
        RECT 538.290 2289.715 538.570 2290.085 ;
        RECT 543.880 2289.890 544.020 2290.395 ;
        RECT 538.360 2288.870 538.500 2289.715 ;
        RECT 543.820 2289.570 544.080 2289.890 ;
        RECT 544.730 2289.715 545.010 2290.085 ;
        RECT 538.300 2288.550 538.560 2288.870 ;
        RECT 542.900 2214.430 543.160 2214.750 ;
        RECT 537.840 2210.010 538.100 2210.330 ;
        RECT 542.960 2200.000 543.100 2214.430 ;
        RECT 544.800 2211.010 544.940 2289.715 ;
        RECT 551.700 2214.750 551.840 2290.395 ;
        RECT 613.800 2289.890 613.940 2290.590 ;
        RECT 635.420 2289.890 635.560 2290.590 ;
        RECT 613.740 2289.570 614.000 2289.890 ;
        RECT 635.360 2289.570 635.620 2289.890 ;
        RECT 668.940 2286.510 669.200 2286.830 ;
        RECT 551.640 2214.430 551.900 2214.750 ;
        RECT 656.520 2214.430 656.780 2214.750 ;
        RECT 544.740 2210.690 545.000 2211.010 ;
        RECT 645.020 2210.690 645.280 2211.010 ;
        RECT 622.480 2210.350 622.740 2210.670 ;
        RECT 610.980 2209.670 611.240 2209.990 ;
        RECT 588.440 2209.330 588.700 2209.650 ;
        RECT 565.900 2208.650 566.160 2208.970 ;
        RECT 554.400 2207.970 554.660 2208.290 ;
        RECT 554.460 2200.000 554.600 2207.970 ;
        RECT 565.960 2200.000 566.100 2208.650 ;
        RECT 576.940 2208.310 577.200 2208.630 ;
        RECT 577.000 2200.000 577.140 2208.310 ;
        RECT 588.500 2200.000 588.640 2209.330 ;
        RECT 599.480 2208.990 599.740 2209.310 ;
        RECT 599.540 2200.000 599.680 2208.990 ;
        RECT 611.040 2200.000 611.180 2209.670 ;
        RECT 622.540 2200.000 622.680 2210.350 ;
        RECT 633.520 2210.010 633.780 2210.330 ;
        RECT 633.580 2200.000 633.720 2210.010 ;
        RECT 645.080 2200.000 645.220 2210.690 ;
        RECT 656.580 2200.000 656.720 2214.430 ;
        RECT 441.310 2199.530 441.590 2200.000 ;
        RECT 439.920 2199.390 441.590 2199.530 ;
        RECT 452.340 2199.460 452.630 2200.000 ;
        RECT 463.840 2199.460 464.130 2200.000 ;
        RECT 475.340 2199.460 475.630 2200.000 ;
        RECT 486.380 2199.460 486.670 2200.000 ;
        RECT 497.880 2199.460 498.170 2200.000 ;
        RECT 509.380 2199.460 509.670 2200.000 ;
        RECT 520.420 2199.460 520.710 2200.000 ;
        RECT 531.920 2199.460 532.210 2200.000 ;
        RECT 542.960 2199.460 543.250 2200.000 ;
        RECT 554.460 2199.460 554.750 2200.000 ;
        RECT 565.960 2199.460 566.250 2200.000 ;
        RECT 577.000 2199.460 577.290 2200.000 ;
        RECT 588.500 2199.460 588.790 2200.000 ;
        RECT 599.540 2199.460 599.830 2200.000 ;
        RECT 611.040 2199.460 611.330 2200.000 ;
        RECT 622.540 2199.460 622.830 2200.000 ;
        RECT 633.580 2199.460 633.870 2200.000 ;
        RECT 645.080 2199.460 645.370 2200.000 ;
        RECT 656.580 2199.460 656.870 2200.000 ;
        RECT 418.770 2196.000 419.050 2199.390 ;
        RECT 429.810 2196.000 430.090 2199.390 ;
        RECT 441.310 2196.000 441.590 2199.390 ;
        RECT 452.350 2196.000 452.630 2199.460 ;
        RECT 463.850 2196.000 464.130 2199.460 ;
        RECT 475.350 2196.000 475.630 2199.460 ;
        RECT 486.390 2196.000 486.670 2199.460 ;
        RECT 497.890 2196.000 498.170 2199.460 ;
        RECT 509.390 2196.000 509.670 2199.460 ;
        RECT 520.430 2196.000 520.710 2199.460 ;
        RECT 531.930 2196.000 532.210 2199.460 ;
        RECT 542.970 2196.000 543.250 2199.460 ;
        RECT 554.470 2196.000 554.750 2199.460 ;
        RECT 565.970 2196.000 566.250 2199.460 ;
        RECT 577.010 2196.000 577.290 2199.460 ;
        RECT 588.510 2196.000 588.790 2199.460 ;
        RECT 599.550 2196.000 599.830 2199.460 ;
        RECT 611.050 2196.000 611.330 2199.460 ;
        RECT 622.550 2196.000 622.830 2199.460 ;
        RECT 633.590 2196.000 633.870 2199.460 ;
        RECT 645.090 2196.000 645.370 2199.460 ;
        RECT 656.590 2196.000 656.870 2199.460 ;
        RECT 667.630 2199.530 667.910 2200.000 ;
        RECT 669.000 2199.530 669.140 2286.510 ;
        RECT 696.600 2214.750 696.740 2697.910 ;
        RECT 697.060 2447.845 697.200 2748.830 ;
        RECT 751.740 2732.250 752.000 2732.570 ;
        RECT 938.490 2732.395 938.770 2732.765 ;
        RECT 938.500 2732.250 938.760 2732.395 ;
        RECT 737.940 2725.450 738.200 2725.770 ;
        RECT 724.140 2718.650 724.400 2718.970 ;
        RECT 717.240 2711.850 717.500 2712.170 ;
        RECT 703.440 2698.250 703.700 2698.570 ;
        RECT 696.990 2447.475 697.270 2447.845 ;
        RECT 690.100 2214.430 690.360 2214.750 ;
        RECT 696.540 2214.430 696.800 2214.750 ;
        RECT 697.000 2214.430 697.260 2214.750 ;
        RECT 679.060 2210.690 679.320 2211.010 ;
        RECT 667.630 2199.390 669.140 2199.530 ;
        RECT 679.120 2200.000 679.260 2210.690 ;
        RECT 690.160 2200.000 690.300 2214.430 ;
        RECT 697.060 2211.010 697.200 2214.430 ;
        RECT 697.000 2210.690 697.260 2211.010 ;
        RECT 679.120 2199.460 679.410 2200.000 ;
        RECT 690.160 2199.460 690.450 2200.000 ;
        RECT 667.630 2196.000 667.910 2199.390 ;
        RECT 679.130 2196.000 679.410 2199.460 ;
        RECT 690.170 2196.000 690.450 2199.460 ;
        RECT 701.670 2199.530 701.950 2200.000 ;
        RECT 703.500 2199.530 703.640 2698.250 ;
        RECT 710.340 2290.590 710.600 2290.910 ;
        RECT 710.400 2289.890 710.540 2290.590 ;
        RECT 710.340 2289.570 710.600 2289.890 ;
        RECT 717.300 2214.410 717.440 2711.850 ;
        RECT 712.640 2214.090 712.900 2214.410 ;
        RECT 713.100 2214.090 713.360 2214.410 ;
        RECT 717.240 2214.090 717.500 2214.410 ;
        RECT 712.700 2211.010 712.840 2214.090 ;
        RECT 712.640 2210.690 712.900 2211.010 ;
        RECT 701.670 2199.390 703.640 2199.530 ;
        RECT 713.160 2200.000 713.300 2214.090 ;
        RECT 724.200 2200.000 724.340 2718.650 ;
        RECT 734.720 2290.590 734.980 2290.910 ;
        RECT 734.780 2289.890 734.920 2290.590 ;
        RECT 734.720 2289.570 734.980 2289.890 ;
        RECT 713.160 2199.460 713.450 2200.000 ;
        RECT 724.200 2199.460 724.490 2200.000 ;
        RECT 701.670 2196.000 701.950 2199.390 ;
        RECT 713.170 2196.000 713.450 2199.460 ;
        RECT 724.210 2196.000 724.490 2199.460 ;
        RECT 735.710 2199.530 735.990 2200.000 ;
        RECT 738.000 2199.530 738.140 2725.450 ;
        RECT 751.800 2214.410 751.940 2732.250 ;
        RECT 938.490 2725.595 938.770 2725.965 ;
        RECT 938.500 2725.450 938.760 2725.595 ;
        RECT 938.490 2718.795 938.770 2719.165 ;
        RECT 938.500 2718.650 938.760 2718.795 ;
        RECT 938.490 2712.675 938.770 2713.045 ;
        RECT 938.560 2712.170 938.700 2712.675 ;
        RECT 938.500 2711.850 938.760 2712.170 ;
        RECT 938.950 2701.795 939.230 2702.165 ;
        RECT 938.490 2699.075 938.770 2699.445 ;
        RECT 938.560 2698.230 938.700 2699.075 ;
        RECT 939.020 2698.570 939.160 2701.795 ;
        RECT 938.960 2698.250 939.220 2698.570 ;
        RECT 938.500 2697.910 938.760 2698.230 ;
        RECT 941.710 2687.515 941.990 2687.885 ;
        RECT 806.940 2290.590 807.200 2290.910 ;
        RECT 807.000 2289.890 807.140 2290.590 ;
        RECT 806.940 2289.570 807.200 2289.890 ;
        RECT 882.840 2288.210 883.100 2288.530 ;
        RECT 875.940 2287.870 876.200 2288.190 ;
        RECT 862.140 2287.530 862.400 2287.850 ;
        RECT 855.240 2286.850 855.500 2287.170 ;
        RECT 746.680 2214.090 746.940 2214.410 ;
        RECT 751.740 2214.090 752.000 2214.410 ;
        RECT 735.710 2199.390 738.140 2199.530 ;
        RECT 746.740 2200.000 746.880 2214.090 ;
        RECT 769.680 2213.750 769.940 2214.070 ;
        RECT 758.180 2210.690 758.440 2211.010 ;
        RECT 758.240 2200.000 758.380 2210.690 ;
        RECT 769.740 2200.000 769.880 2213.750 ;
        RECT 780.720 2213.410 780.980 2213.730 ;
        RECT 780.780 2200.000 780.920 2213.410 ;
        RECT 792.220 2213.070 792.480 2213.390 ;
        RECT 792.280 2200.000 792.420 2213.070 ;
        RECT 803.260 2212.730 803.520 2213.050 ;
        RECT 803.320 2200.000 803.460 2212.730 ;
        RECT 814.750 2212.195 815.030 2212.565 ;
        RECT 814.820 2200.000 814.960 2212.195 ;
        RECT 826.250 2211.515 826.530 2211.885 ;
        RECT 826.320 2200.000 826.460 2211.515 ;
        RECT 837.290 2210.835 837.570 2211.205 ;
        RECT 837.360 2200.000 837.500 2210.835 ;
        RECT 855.300 2209.990 855.440 2286.850 ;
        RECT 848.800 2209.670 849.060 2209.990 ;
        RECT 855.240 2209.670 855.500 2209.990 ;
        RECT 848.860 2200.000 849.000 2209.670 ;
        RECT 746.740 2199.460 747.030 2200.000 ;
        RECT 758.240 2199.460 758.530 2200.000 ;
        RECT 769.740 2199.460 770.030 2200.000 ;
        RECT 780.780 2199.460 781.070 2200.000 ;
        RECT 792.280 2199.460 792.570 2200.000 ;
        RECT 803.320 2199.460 803.610 2200.000 ;
        RECT 814.820 2199.460 815.110 2200.000 ;
        RECT 826.320 2199.460 826.610 2200.000 ;
        RECT 837.360 2199.460 837.650 2200.000 ;
        RECT 848.860 2199.460 849.150 2200.000 ;
        RECT 735.710 2196.000 735.990 2199.390 ;
        RECT 746.750 2196.000 747.030 2199.460 ;
        RECT 758.250 2196.000 758.530 2199.460 ;
        RECT 769.750 2196.000 770.030 2199.460 ;
        RECT 780.790 2196.000 781.070 2199.460 ;
        RECT 792.290 2196.000 792.570 2199.460 ;
        RECT 803.330 2196.000 803.610 2199.460 ;
        RECT 814.830 2196.000 815.110 2199.460 ;
        RECT 826.330 2196.000 826.610 2199.460 ;
        RECT 837.370 2196.000 837.650 2199.460 ;
        RECT 848.870 2196.000 849.150 2199.460 ;
        RECT 860.370 2199.530 860.650 2200.000 ;
        RECT 862.200 2199.530 862.340 2287.530 ;
        RECT 876.000 2211.010 876.140 2287.870 ;
        RECT 871.340 2210.690 871.600 2211.010 ;
        RECT 875.940 2210.690 876.200 2211.010 ;
        RECT 860.370 2199.390 862.340 2199.530 ;
        RECT 871.400 2200.000 871.540 2210.690 ;
        RECT 882.900 2200.000 883.040 2288.210 ;
        RECT 941.780 2214.750 941.920 2687.515 ;
        RECT 944.930 2401.235 945.210 2401.605 ;
        RECT 944.470 2389.675 944.750 2390.045 ;
        RECT 944.540 2301.110 944.680 2389.675 ;
        RECT 944.480 2300.790 944.740 2301.110 ;
        RECT 944.540 2297.710 944.680 2300.790 ;
        RECT 944.480 2297.390 944.740 2297.710 ;
        RECT 941.720 2214.430 941.980 2214.750 ;
        RECT 945.000 2213.050 945.140 2401.235 ;
      LAYER met2 ;
        RECT 955.000 2305.000 1331.480 2751.235 ;
      LAYER met2 ;
        RECT 1332.320 2749.765 1332.460 2751.290 ;
        RECT 1332.250 2749.395 1332.530 2749.765 ;
        RECT 1352.030 2746.675 1352.310 2747.045 ;
        RECT 1352.100 2746.510 1352.240 2746.675 ;
        RECT 1511.260 2746.510 1511.400 2751.290 ;
        RECT 1352.040 2746.190 1352.300 2746.510 ;
        RECT 1511.200 2746.190 1511.460 2746.510 ;
        RECT 1345.590 2422.315 1345.870 2422.685 ;
        RECT 1345.660 2422.150 1345.800 2422.315 ;
        RECT 1345.600 2421.830 1345.860 2422.150 ;
        RECT 1076.560 2290.910 1076.700 2291.065 ;
        RECT 952.300 2290.590 952.560 2290.910 ;
        RECT 1000.140 2290.590 1000.400 2290.910 ;
        RECT 952.360 2289.890 952.500 2290.590 ;
        RECT 952.300 2289.570 952.560 2289.890 ;
        RECT 986.790 2289.715 987.070 2290.085 ;
        RECT 993.690 2289.715 993.970 2290.085 ;
        RECT 1000.200 2289.890 1000.340 2290.590 ;
        RECT 1001.050 2290.395 1001.330 2290.765 ;
        RECT 1048.900 2290.650 1049.160 2290.910 ;
        RECT 1076.500 2290.765 1076.760 2290.910 ;
        RECT 1048.900 2290.590 1049.560 2290.650 ;
        RECT 1048.960 2290.510 1049.560 2290.590 ;
        RECT 979.890 2287.675 980.170 2288.045 ;
        RECT 979.960 2286.830 980.100 2287.675 ;
        RECT 986.860 2287.170 987.000 2289.715 ;
        RECT 993.760 2287.850 993.900 2289.715 ;
        RECT 1000.140 2289.570 1000.400 2289.890 ;
        RECT 1001.120 2288.190 1001.260 2290.395 ;
        RECT 1038.310 2289.715 1038.590 2290.085 ;
        RECT 1041.070 2289.715 1041.350 2290.085 ;
        RECT 1007.490 2288.355 1007.770 2288.725 ;
        RECT 1007.500 2288.210 1007.760 2288.355 ;
        RECT 1001.060 2287.870 1001.320 2288.190 ;
        RECT 993.700 2287.530 993.960 2287.850 ;
        RECT 986.800 2286.850 987.060 2287.170 ;
        RECT 979.900 2286.510 980.160 2286.830 ;
        RECT 1010.720 2286.510 1010.980 2286.830 ;
        RECT 1010.780 2286.005 1010.920 2286.510 ;
        RECT 1031.410 2286.315 1031.690 2286.685 ;
        RECT 1034.170 2286.315 1034.450 2286.685 ;
        RECT 1010.710 2285.635 1010.990 2286.005 ;
        RECT 1013.930 2285.635 1014.210 2286.005 ;
        RECT 1007.500 2213.750 1007.760 2214.070 ;
        RECT 996.000 2213.070 996.260 2213.390 ;
        RECT 939.420 2212.730 939.680 2213.050 ;
        RECT 944.940 2212.730 945.200 2213.050 ;
        RECT 893.880 2212.390 894.140 2212.710 ;
        RECT 893.940 2200.000 894.080 2212.390 ;
        RECT 905.380 2212.050 905.640 2212.370 ;
        RECT 905.440 2200.000 905.580 2212.050 ;
        RECT 916.880 2211.710 917.140 2212.030 ;
        RECT 916.940 2200.000 917.080 2211.710 ;
        RECT 927.920 2211.370 928.180 2211.690 ;
        RECT 927.980 2200.000 928.120 2211.370 ;
        RECT 939.480 2200.000 939.620 2212.730 ;
        RECT 973.460 2211.710 973.720 2212.030 ;
        RECT 950.460 2211.030 950.720 2211.350 ;
        RECT 961.960 2211.030 962.220 2211.350 ;
        RECT 950.520 2200.000 950.660 2211.030 ;
        RECT 962.020 2200.000 962.160 2211.030 ;
        RECT 973.520 2200.000 973.660 2211.710 ;
        RECT 984.500 2211.370 984.760 2211.690 ;
        RECT 984.560 2200.000 984.700 2211.370 ;
        RECT 996.060 2200.000 996.200 2213.070 ;
        RECT 1007.560 2200.000 1007.700 2213.750 ;
        RECT 1010.780 2211.350 1010.920 2285.635 ;
        RECT 1014.000 2213.050 1014.140 2285.635 ;
        RECT 1024.510 2284.955 1024.790 2285.325 ;
        RECT 1027.270 2284.955 1027.550 2285.325 ;
        RECT 1017.610 2284.275 1017.890 2284.645 ;
        RECT 1020.830 2284.275 1021.110 2284.645 ;
        RECT 1017.680 2284.110 1017.820 2284.275 ;
        RECT 1017.620 2283.790 1017.880 2284.110 ;
        RECT 1013.940 2212.730 1014.200 2213.050 ;
        RECT 1017.680 2212.030 1017.820 2283.790 ;
        RECT 1020.900 2212.710 1021.040 2284.275 ;
        RECT 1020.840 2212.390 1021.100 2212.710 ;
        RECT 1017.620 2211.710 1017.880 2212.030 ;
        RECT 1024.580 2211.690 1024.720 2284.955 ;
        RECT 1027.340 2284.450 1027.480 2284.955 ;
        RECT 1027.280 2284.130 1027.540 2284.450 ;
        RECT 1027.730 2284.275 1028.010 2284.645 ;
        RECT 1027.800 2212.370 1027.940 2284.275 ;
        RECT 1030.040 2214.430 1030.300 2214.750 ;
        RECT 1027.740 2212.050 1028.000 2212.370 ;
        RECT 1024.520 2211.370 1024.780 2211.690 ;
        RECT 1010.720 2211.030 1010.980 2211.350 ;
        RECT 1018.540 2209.330 1018.800 2209.650 ;
        RECT 1018.600 2200.000 1018.740 2209.330 ;
        RECT 1030.100 2200.000 1030.240 2214.430 ;
        RECT 1031.480 2213.390 1031.620 2286.315 ;
        RECT 1034.240 2284.790 1034.380 2286.315 ;
        RECT 1034.630 2285.635 1034.910 2286.005 ;
        RECT 1034.180 2284.470 1034.440 2284.790 ;
        RECT 1031.420 2213.070 1031.680 2213.390 ;
        RECT 1034.700 2212.030 1034.840 2285.635 ;
        RECT 1038.380 2214.070 1038.520 2289.715 ;
        RECT 1041.140 2289.550 1041.280 2289.715 ;
        RECT 1041.080 2289.230 1041.340 2289.550 ;
        RECT 1038.780 2288.210 1039.040 2288.530 ;
        RECT 1048.430 2288.355 1048.710 2288.725 ;
        RECT 1048.440 2288.210 1048.700 2288.355 ;
        RECT 1038.840 2214.750 1038.980 2288.210 ;
        RECT 1045.680 2287.870 1045.940 2288.190 ;
        RECT 1045.210 2286.995 1045.490 2287.365 ;
        RECT 1045.220 2286.850 1045.480 2286.995 ;
        RECT 1041.530 2284.275 1041.810 2284.645 ;
        RECT 1038.780 2214.430 1039.040 2214.750 ;
        RECT 1041.080 2214.430 1041.340 2214.750 ;
        RECT 1038.320 2213.750 1038.580 2214.070 ;
        RECT 1034.640 2211.710 1034.900 2212.030 ;
        RECT 1041.140 2200.000 1041.280 2214.430 ;
        RECT 1041.600 2211.690 1041.740 2284.275 ;
        RECT 1041.540 2211.370 1041.800 2211.690 ;
        RECT 1045.280 2209.650 1045.420 2286.850 ;
        RECT 1045.740 2214.750 1045.880 2287.870 ;
        RECT 1049.420 2286.490 1049.560 2290.510 ;
        RECT 1052.570 2290.395 1052.850 2290.765 ;
        RECT 1062.230 2290.395 1062.510 2290.765 ;
        RECT 1065.450 2290.395 1065.730 2290.765 ;
        RECT 1070.050 2290.395 1070.330 2290.765 ;
        RECT 1076.490 2290.395 1076.770 2290.765 ;
        RECT 1083.390 2290.395 1083.670 2290.765 ;
        RECT 1086.160 2290.590 1086.420 2290.910 ;
        RECT 1052.640 2288.190 1052.780 2290.395 ;
        RECT 1052.580 2287.870 1052.840 2288.190 ;
        RECT 1062.300 2287.850 1062.440 2290.395 ;
        RECT 1065.520 2289.210 1065.660 2290.395 ;
        RECT 1065.460 2288.890 1065.720 2289.210 ;
        RECT 1062.240 2287.530 1062.500 2287.850 ;
        RECT 1062.300 2286.830 1062.440 2287.530 ;
        RECT 1062.240 2286.510 1062.500 2286.830 ;
        RECT 1048.900 2286.170 1049.160 2286.490 ;
        RECT 1049.360 2286.170 1049.620 2286.490 ;
        RECT 1048.430 2284.275 1048.710 2284.645 ;
        RECT 1045.680 2214.430 1045.940 2214.750 ;
        RECT 1048.500 2211.350 1048.640 2284.275 ;
        RECT 1048.440 2211.030 1048.700 2211.350 ;
        RECT 1045.220 2209.330 1045.480 2209.650 ;
        RECT 1048.960 2202.250 1049.100 2286.170 ;
        RECT 1054.870 2285.635 1055.150 2286.005 ;
        RECT 1062.700 2285.830 1062.960 2286.150 ;
        RECT 1054.940 2208.290 1055.080 2285.635 ;
        RECT 1055.330 2284.275 1055.610 2284.645 ;
        RECT 1062.230 2284.275 1062.510 2284.645 ;
        RECT 1055.400 2208.970 1055.540 2284.275 ;
        RECT 1055.340 2208.650 1055.600 2208.970 ;
        RECT 1062.300 2208.630 1062.440 2284.275 ;
        RECT 1062.240 2208.310 1062.500 2208.630 ;
        RECT 1054.880 2207.970 1055.140 2208.290 ;
        RECT 1048.960 2202.110 1050.940 2202.250 ;
        RECT 871.400 2199.460 871.690 2200.000 ;
        RECT 882.900 2199.460 883.190 2200.000 ;
        RECT 893.940 2199.460 894.230 2200.000 ;
        RECT 905.440 2199.460 905.730 2200.000 ;
        RECT 916.940 2199.460 917.230 2200.000 ;
        RECT 927.980 2199.460 928.270 2200.000 ;
        RECT 939.480 2199.460 939.770 2200.000 ;
        RECT 950.520 2199.460 950.810 2200.000 ;
        RECT 962.020 2199.460 962.310 2200.000 ;
        RECT 973.520 2199.460 973.810 2200.000 ;
        RECT 984.560 2199.460 984.850 2200.000 ;
        RECT 996.060 2199.460 996.350 2200.000 ;
        RECT 1007.560 2199.460 1007.850 2200.000 ;
        RECT 1018.600 2199.460 1018.890 2200.000 ;
        RECT 1030.100 2199.460 1030.390 2200.000 ;
        RECT 1041.140 2199.460 1041.430 2200.000 ;
        RECT 860.370 2196.000 860.650 2199.390 ;
        RECT 871.410 2196.000 871.690 2199.460 ;
        RECT 882.910 2196.000 883.190 2199.460 ;
        RECT 893.950 2196.000 894.230 2199.460 ;
        RECT 905.450 2196.000 905.730 2199.460 ;
        RECT 916.950 2196.000 917.230 2199.460 ;
        RECT 927.990 2196.000 928.270 2199.460 ;
        RECT 939.490 2196.000 939.770 2199.460 ;
        RECT 950.530 2196.000 950.810 2199.460 ;
        RECT 962.030 2196.000 962.310 2199.460 ;
        RECT 973.530 2196.000 973.810 2199.460 ;
        RECT 984.570 2196.000 984.850 2199.460 ;
        RECT 996.070 2196.000 996.350 2199.460 ;
        RECT 1007.570 2196.000 1007.850 2199.460 ;
        RECT 1018.610 2196.000 1018.890 2199.460 ;
        RECT 1030.110 2196.000 1030.390 2199.460 ;
        RECT 1041.150 2196.000 1041.430 2199.460 ;
        RECT 1050.800 2199.530 1050.940 2202.110 ;
        RECT 1052.650 2199.530 1052.930 2200.000 ;
        RECT 1050.800 2199.390 1052.930 2199.530 ;
        RECT 1062.760 2199.530 1062.900 2285.830 ;
        RECT 1065.520 2284.110 1065.660 2288.890 ;
        RECT 1070.120 2288.870 1070.260 2290.395 ;
        RECT 1070.060 2288.550 1070.320 2288.870 ;
        RECT 1069.600 2285.490 1069.860 2285.810 ;
        RECT 1069.130 2284.275 1069.410 2284.645 ;
        RECT 1065.460 2283.790 1065.720 2284.110 ;
        RECT 1069.200 2209.310 1069.340 2284.275 ;
        RECT 1069.140 2208.990 1069.400 2209.310 ;
        RECT 1069.660 2202.250 1069.800 2285.490 ;
        RECT 1070.120 2284.450 1070.260 2288.550 ;
        RECT 1076.030 2285.635 1076.310 2286.005 ;
        RECT 1076.040 2285.490 1076.300 2285.635 ;
        RECT 1076.560 2284.790 1076.700 2290.395 ;
        RECT 1083.460 2289.550 1083.600 2290.395 ;
        RECT 1086.220 2289.550 1086.360 2290.590 ;
        RECT 1087.990 2290.395 1088.270 2290.765 ;
        RECT 1094.430 2290.395 1094.710 2290.765 ;
        RECT 1096.740 2290.590 1097.000 2290.910 ;
        RECT 1083.400 2289.230 1083.660 2289.550 ;
        RECT 1085.700 2289.230 1085.960 2289.550 ;
        RECT 1086.160 2289.230 1086.420 2289.550 ;
        RECT 1082.930 2286.995 1083.210 2287.365 ;
        RECT 1085.760 2287.170 1085.900 2289.230 ;
        RECT 1076.500 2284.470 1076.760 2284.790 ;
        RECT 1083.000 2284.450 1083.140 2286.995 ;
        RECT 1085.700 2286.850 1085.960 2287.170 ;
        RECT 1088.060 2286.830 1088.200 2290.395 ;
        RECT 1094.500 2288.530 1094.640 2290.395 ;
        RECT 1094.440 2288.210 1094.700 2288.530 ;
        RECT 1088.000 2286.510 1088.260 2286.830 ;
        RECT 1096.800 2286.490 1096.940 2290.590 ;
        RECT 1100.870 2290.395 1101.150 2290.765 ;
        RECT 1106.850 2290.395 1107.130 2290.765 ;
        RECT 1112.830 2290.395 1113.110 2290.765 ;
        RECT 1100.940 2288.190 1101.080 2290.395 ;
        RECT 1104.100 2289.910 1104.360 2290.230 ;
        RECT 1100.880 2287.870 1101.140 2288.190 ;
        RECT 1096.740 2286.170 1097.000 2286.490 ;
        RECT 1089.830 2285.635 1090.110 2286.005 ;
        RECT 1103.630 2285.635 1103.910 2286.005 ;
        RECT 1083.400 2285.150 1083.660 2285.470 ;
        RECT 1070.060 2284.130 1070.320 2284.450 ;
        RECT 1082.940 2284.130 1083.200 2284.450 ;
        RECT 1083.460 2202.250 1083.600 2285.150 ;
        RECT 1089.370 2284.275 1089.650 2284.645 ;
        RECT 1089.440 2209.990 1089.580 2284.275 ;
        RECT 1089.900 2284.110 1090.040 2285.635 ;
        RECT 1097.200 2284.810 1097.460 2285.130 ;
        RECT 1096.730 2284.275 1097.010 2284.645 ;
        RECT 1089.840 2283.790 1090.100 2284.110 ;
        RECT 1089.380 2209.670 1089.640 2209.990 ;
        RECT 1096.800 2209.650 1096.940 2284.275 ;
        RECT 1096.740 2209.330 1097.000 2209.650 ;
        RECT 1069.660 2202.110 1073.940 2202.250 ;
        RECT 1083.460 2202.110 1084.980 2202.250 ;
        RECT 1064.150 2199.530 1064.430 2200.000 ;
        RECT 1062.760 2199.390 1064.430 2199.530 ;
        RECT 1073.800 2199.530 1073.940 2202.110 ;
        RECT 1075.190 2199.530 1075.470 2200.000 ;
        RECT 1073.800 2199.390 1075.470 2199.530 ;
        RECT 1084.840 2199.530 1084.980 2202.110 ;
        RECT 1086.690 2199.530 1086.970 2200.000 ;
        RECT 1084.840 2199.390 1086.970 2199.530 ;
        RECT 1097.260 2199.530 1097.400 2284.810 ;
        RECT 1103.700 2210.670 1103.840 2285.635 ;
        RECT 1103.640 2210.350 1103.900 2210.670 ;
        RECT 1104.160 2202.250 1104.300 2289.910 ;
        RECT 1106.920 2287.850 1107.060 2290.395 ;
        RECT 1112.900 2289.210 1113.040 2290.395 ;
        RECT 1117.900 2290.250 1118.160 2290.570 ;
        RECT 1118.350 2290.395 1118.630 2290.765 ;
        RECT 1121.570 2290.395 1121.850 2290.765 ;
        RECT 1129.390 2290.395 1129.670 2290.765 ;
        RECT 1131.700 2290.590 1131.960 2290.910 ;
        RECT 1118.360 2290.250 1118.620 2290.395 ;
        RECT 1112.840 2288.890 1113.100 2289.210 ;
        RECT 1106.860 2287.530 1107.120 2287.850 ;
        RECT 1110.530 2284.275 1110.810 2284.645 ;
        RECT 1117.430 2284.275 1117.710 2284.645 ;
        RECT 1110.600 2210.330 1110.740 2284.275 ;
        RECT 1117.500 2211.010 1117.640 2284.275 ;
        RECT 1117.440 2210.690 1117.700 2211.010 ;
        RECT 1110.540 2210.010 1110.800 2210.330 ;
        RECT 1117.960 2202.250 1118.100 2290.250 ;
        RECT 1118.420 2288.870 1118.560 2290.250 ;
        RECT 1121.640 2290.230 1121.780 2290.395 ;
        RECT 1121.580 2289.910 1121.840 2290.230 ;
        RECT 1121.640 2289.550 1121.780 2289.910 ;
        RECT 1129.460 2289.890 1129.600 2290.395 ;
        RECT 1124.800 2289.570 1125.060 2289.890 ;
        RECT 1129.400 2289.570 1129.660 2289.890 ;
        RECT 1121.580 2289.230 1121.840 2289.550 ;
        RECT 1118.360 2288.550 1118.620 2288.870 ;
        RECT 1124.860 2287.170 1125.000 2289.570 ;
        RECT 1124.800 2286.850 1125.060 2287.170 ;
        RECT 1131.230 2284.955 1131.510 2285.325 ;
        RECT 1124.330 2284.275 1124.610 2284.645 ;
        RECT 1130.770 2284.275 1131.050 2284.645 ;
        RECT 1124.400 2214.750 1124.540 2284.275 ;
        RECT 1124.340 2214.430 1124.600 2214.750 ;
        RECT 1130.840 2214.070 1130.980 2284.275 ;
        RECT 1131.300 2214.410 1131.440 2284.955 ;
        RECT 1131.240 2214.090 1131.500 2214.410 ;
        RECT 1130.780 2213.750 1131.040 2214.070 ;
        RECT 1104.160 2202.110 1107.980 2202.250 ;
        RECT 1117.960 2202.110 1119.020 2202.250 ;
        RECT 1097.730 2199.530 1098.010 2200.000 ;
        RECT 1097.260 2199.390 1098.010 2199.530 ;
        RECT 1107.840 2199.530 1107.980 2202.110 ;
        RECT 1109.230 2199.530 1109.510 2200.000 ;
        RECT 1107.840 2199.390 1109.510 2199.530 ;
        RECT 1118.880 2199.530 1119.020 2202.110 ;
        RECT 1131.760 2200.000 1131.900 2290.590 ;
        RECT 1135.830 2290.395 1136.110 2290.765 ;
        RECT 1141.810 2290.395 1142.090 2290.765 ;
        RECT 1147.790 2290.395 1148.070 2290.765 ;
        RECT 1159.290 2290.395 1159.570 2290.765 ;
        RECT 1166.190 2290.395 1166.470 2290.765 ;
        RECT 1135.900 2288.870 1136.040 2290.395 ;
        RECT 1132.160 2288.550 1132.420 2288.870 ;
        RECT 1135.840 2288.550 1136.100 2288.870 ;
        RECT 1132.220 2286.830 1132.360 2288.550 ;
        RECT 1141.880 2288.530 1142.020 2290.395 ;
        RECT 1141.820 2288.210 1142.080 2288.530 ;
        RECT 1147.860 2288.190 1148.000 2290.395 ;
        RECT 1159.300 2290.250 1159.560 2290.395 ;
        RECT 1166.260 2290.230 1166.400 2290.395 ;
        RECT 1166.200 2289.910 1166.460 2290.230 ;
        RECT 1173.090 2289.715 1173.370 2290.085 ;
        RECT 1173.100 2289.570 1173.360 2289.715 ;
        RECT 1159.290 2289.035 1159.570 2289.405 ;
        RECT 1179.990 2289.035 1180.270 2289.405 ;
        RECT 1159.300 2288.890 1159.560 2289.035 ;
        RECT 1180.060 2288.870 1180.200 2289.035 ;
        RECT 1180.000 2288.550 1180.260 2288.870 ;
        RECT 1186.890 2288.355 1187.170 2288.725 ;
        RECT 1193.790 2288.355 1194.070 2288.725 ;
        RECT 1186.900 2288.210 1187.160 2288.355 ;
        RECT 1193.860 2288.190 1194.000 2288.355 ;
        RECT 1147.800 2287.870 1148.060 2288.190 ;
        RECT 1152.390 2287.675 1152.670 2288.045 ;
        RECT 1193.800 2287.870 1194.060 2288.190 ;
        RECT 1152.400 2287.530 1152.660 2287.675 ;
        RECT 1132.160 2286.510 1132.420 2286.830 ;
        RECT 1231.520 2285.490 1231.780 2285.810 ;
        RECT 1165.270 2284.955 1165.550 2285.325 ;
        RECT 1138.130 2284.275 1138.410 2284.645 ;
        RECT 1145.030 2284.275 1145.310 2284.645 ;
        RECT 1151.930 2284.275 1152.210 2284.645 ;
        RECT 1158.830 2284.275 1159.110 2284.645 ;
        RECT 1138.200 2213.730 1138.340 2284.275 ;
        RECT 1138.140 2213.410 1138.400 2213.730 ;
        RECT 1145.100 2213.390 1145.240 2284.275 ;
        RECT 1145.040 2213.070 1145.300 2213.390 ;
        RECT 1152.000 2213.050 1152.140 2284.275 ;
        RECT 1143.200 2212.730 1143.460 2213.050 ;
        RECT 1151.940 2212.730 1152.200 2213.050 ;
        RECT 1143.260 2200.000 1143.400 2212.730 ;
        RECT 1158.900 2212.710 1159.040 2284.275 ;
        RECT 1154.240 2212.390 1154.500 2212.710 ;
        RECT 1158.840 2212.390 1159.100 2212.710 ;
        RECT 1154.300 2200.000 1154.440 2212.390 ;
        RECT 1165.340 2212.370 1165.480 2284.955 ;
        RECT 1165.730 2284.275 1166.010 2284.645 ;
        RECT 1172.630 2284.275 1172.910 2284.645 ;
        RECT 1179.530 2284.275 1179.810 2284.645 ;
        RECT 1186.430 2284.275 1186.710 2284.645 ;
        RECT 1193.330 2284.275 1193.610 2284.645 ;
        RECT 1200.230 2284.275 1200.510 2284.645 ;
        RECT 1165.800 2212.565 1165.940 2284.275 ;
        RECT 1163.900 2212.050 1164.160 2212.370 ;
        RECT 1165.280 2212.050 1165.540 2212.370 ;
        RECT 1165.730 2212.195 1166.010 2212.565 ;
        RECT 1120.730 2199.530 1121.010 2200.000 ;
        RECT 1118.880 2199.390 1121.010 2199.530 ;
        RECT 1131.760 2199.460 1132.050 2200.000 ;
        RECT 1143.260 2199.460 1143.550 2200.000 ;
        RECT 1154.300 2199.460 1154.590 2200.000 ;
        RECT 1052.650 2196.000 1052.930 2199.390 ;
        RECT 1064.150 2196.000 1064.430 2199.390 ;
        RECT 1075.190 2196.000 1075.470 2199.390 ;
        RECT 1086.690 2196.000 1086.970 2199.390 ;
        RECT 1097.730 2196.000 1098.010 2199.390 ;
        RECT 1109.230 2196.000 1109.510 2199.390 ;
        RECT 1120.730 2196.000 1121.010 2199.390 ;
        RECT 1131.770 2196.000 1132.050 2199.460 ;
        RECT 1143.270 2196.000 1143.550 2199.460 ;
        RECT 1154.310 2196.000 1154.590 2199.460 ;
        RECT 1163.960 2199.530 1164.100 2212.050 ;
        RECT 1172.700 2211.885 1172.840 2284.275 ;
        RECT 1179.600 2212.030 1179.740 2284.275 ;
        RECT 1172.630 2211.515 1172.910 2211.885 ;
        RECT 1177.240 2211.710 1177.500 2212.030 ;
        RECT 1179.540 2211.710 1179.800 2212.030 ;
        RECT 1177.300 2200.000 1177.440 2211.710 ;
        RECT 1186.500 2211.205 1186.640 2284.275 ;
        RECT 1193.400 2211.690 1193.540 2284.275 ;
        RECT 1188.280 2211.370 1188.540 2211.690 ;
        RECT 1193.340 2211.370 1193.600 2211.690 ;
        RECT 1186.430 2210.835 1186.710 2211.205 ;
        RECT 1188.340 2200.000 1188.480 2211.370 ;
        RECT 1199.780 2211.030 1200.040 2211.350 ;
        RECT 1199.840 2200.000 1199.980 2211.030 ;
        RECT 1200.300 2208.485 1200.440 2284.275 ;
        RECT 1224.620 2284.130 1224.880 2284.450 ;
        RECT 1210.820 2283.790 1211.080 2284.110 ;
        RECT 1210.880 2232.170 1211.020 2283.790 ;
        RECT 1210.880 2232.030 1211.940 2232.170 ;
        RECT 1211.800 2216.450 1211.940 2232.030 ;
        RECT 1211.740 2216.130 1212.000 2216.450 ;
        RECT 1210.360 2211.030 1210.620 2211.350 ;
        RECT 1210.420 2208.630 1210.560 2211.030 ;
        RECT 1224.680 2209.310 1224.820 2284.130 ;
        RECT 1225.540 2216.130 1225.800 2216.450 ;
        RECT 1224.620 2208.990 1224.880 2209.310 ;
        RECT 1222.320 2208.650 1222.580 2208.970 ;
        RECT 1200.230 2208.115 1200.510 2208.485 ;
        RECT 1210.360 2208.310 1210.620 2208.630 ;
        RECT 1211.280 2207.970 1211.540 2208.290 ;
        RECT 1211.340 2200.000 1211.480 2207.970 ;
        RECT 1222.380 2200.000 1222.520 2208.650 ;
        RECT 1225.600 2208.290 1225.740 2216.130 ;
        RECT 1231.580 2211.350 1231.720 2285.490 ;
        RECT 1346.980 2214.430 1347.240 2214.750 ;
        RECT 1231.060 2211.030 1231.320 2211.350 ;
        RECT 1231.520 2211.030 1231.780 2211.350 ;
        RECT 1256.360 2211.030 1256.620 2211.350 ;
        RECT 1256.820 2211.030 1257.080 2211.350 ;
        RECT 1225.540 2207.970 1225.800 2208.290 ;
        RECT 1165.810 2199.530 1166.090 2200.000 ;
        RECT 1163.960 2199.390 1166.090 2199.530 ;
        RECT 1177.300 2199.460 1177.590 2200.000 ;
        RECT 1188.340 2199.460 1188.630 2200.000 ;
        RECT 1199.840 2199.460 1200.130 2200.000 ;
        RECT 1211.340 2199.460 1211.630 2200.000 ;
        RECT 1222.380 2199.460 1222.670 2200.000 ;
        RECT 1165.810 2196.000 1166.090 2199.390 ;
        RECT 1177.310 2196.000 1177.590 2199.460 ;
        RECT 1188.350 2196.000 1188.630 2199.460 ;
        RECT 1199.850 2196.000 1200.130 2199.460 ;
        RECT 1211.350 2196.000 1211.630 2199.460 ;
        RECT 1222.390 2196.000 1222.670 2199.460 ;
        RECT 1231.120 2199.530 1231.260 2211.030 ;
        RECT 1243.020 2208.650 1243.280 2208.970 ;
        RECT 1243.480 2208.650 1243.740 2208.970 ;
        RECT 1233.890 2199.530 1234.170 2200.000 ;
        RECT 1231.120 2199.390 1234.170 2199.530 ;
        RECT 1243.080 2199.530 1243.220 2208.650 ;
        RECT 1243.540 2208.485 1243.680 2208.650 ;
        RECT 1243.470 2208.115 1243.750 2208.485 ;
        RECT 1256.420 2200.000 1256.560 2211.030 ;
        RECT 1256.880 2208.970 1257.020 2211.030 ;
        RECT 1335.480 2210.690 1335.740 2211.010 ;
        RECT 1312.940 2210.350 1313.200 2210.670 ;
        RECT 1290.400 2209.670 1290.660 2209.990 ;
        RECT 1267.860 2208.990 1268.120 2209.310 ;
        RECT 1256.820 2208.650 1257.080 2208.970 ;
        RECT 1267.920 2200.000 1268.060 2208.990 ;
        RECT 1278.900 2207.970 1279.160 2208.290 ;
        RECT 1278.960 2200.000 1279.100 2207.970 ;
        RECT 1290.460 2200.000 1290.600 2209.670 ;
        RECT 1301.440 2209.330 1301.700 2209.650 ;
        RECT 1301.500 2200.000 1301.640 2209.330 ;
        RECT 1313.000 2200.000 1313.140 2210.350 ;
        RECT 1324.440 2210.010 1324.700 2210.330 ;
        RECT 1324.500 2200.000 1324.640 2210.010 ;
        RECT 1335.540 2200.000 1335.680 2210.690 ;
        RECT 1347.040 2200.000 1347.180 2214.430 ;
        RECT 1358.480 2214.090 1358.740 2214.410 ;
        RECT 1358.540 2200.000 1358.680 2214.090 ;
        RECT 1369.520 2213.750 1369.780 2214.070 ;
        RECT 1369.580 2200.000 1369.720 2213.750 ;
        RECT 1381.020 2213.410 1381.280 2213.730 ;
        RECT 1381.080 2200.000 1381.220 2213.410 ;
        RECT 1392.060 2213.070 1392.320 2213.390 ;
        RECT 1392.120 2200.000 1392.260 2213.070 ;
        RECT 1403.560 2212.730 1403.820 2213.050 ;
        RECT 1403.620 2200.000 1403.760 2212.730 ;
        RECT 1415.060 2212.390 1415.320 2212.710 ;
        RECT 1415.120 2200.000 1415.260 2212.390 ;
        RECT 1426.100 2212.050 1426.360 2212.370 ;
        RECT 1437.590 2212.195 1437.870 2212.565 ;
        RECT 1426.160 2200.000 1426.300 2212.050 ;
        RECT 1437.660 2200.000 1437.800 2212.195 ;
        RECT 1448.630 2211.515 1448.910 2211.885 ;
        RECT 1460.140 2211.710 1460.400 2212.030 ;
        RECT 1448.700 2200.000 1448.840 2211.515 ;
        RECT 1460.200 2200.000 1460.340 2211.710 ;
        RECT 1482.680 2211.370 1482.940 2211.690 ;
        RECT 1471.630 2210.835 1471.910 2211.205 ;
        RECT 1471.700 2200.000 1471.840 2210.835 ;
        RECT 1482.740 2200.000 1482.880 2211.370 ;
        RECT 1494.180 2211.030 1494.440 2211.350 ;
        RECT 1494.240 2200.000 1494.380 2211.030 ;
        RECT 1244.930 2199.530 1245.210 2200.000 ;
        RECT 1243.080 2199.390 1245.210 2199.530 ;
        RECT 1256.420 2199.460 1256.710 2200.000 ;
        RECT 1267.920 2199.460 1268.210 2200.000 ;
        RECT 1278.960 2199.460 1279.250 2200.000 ;
        RECT 1290.460 2199.460 1290.750 2200.000 ;
        RECT 1301.500 2199.460 1301.790 2200.000 ;
        RECT 1313.000 2199.460 1313.290 2200.000 ;
        RECT 1324.500 2199.460 1324.790 2200.000 ;
        RECT 1335.540 2199.460 1335.830 2200.000 ;
        RECT 1347.040 2199.460 1347.330 2200.000 ;
        RECT 1358.540 2199.460 1358.830 2200.000 ;
        RECT 1369.580 2199.460 1369.870 2200.000 ;
        RECT 1381.080 2199.460 1381.370 2200.000 ;
        RECT 1392.120 2199.460 1392.410 2200.000 ;
        RECT 1403.620 2199.460 1403.910 2200.000 ;
        RECT 1415.120 2199.460 1415.410 2200.000 ;
        RECT 1426.160 2199.460 1426.450 2200.000 ;
        RECT 1437.660 2199.460 1437.950 2200.000 ;
        RECT 1448.700 2199.460 1448.990 2200.000 ;
        RECT 1460.200 2199.460 1460.490 2200.000 ;
        RECT 1471.700 2199.460 1471.990 2200.000 ;
        RECT 1482.740 2199.460 1483.030 2200.000 ;
        RECT 1494.240 2199.460 1494.530 2200.000 ;
        RECT 1233.890 2196.000 1234.170 2199.390 ;
        RECT 1244.930 2196.000 1245.210 2199.390 ;
        RECT 1256.430 2196.000 1256.710 2199.460 ;
        RECT 1267.930 2196.000 1268.210 2199.460 ;
        RECT 1278.970 2196.000 1279.250 2199.460 ;
        RECT 1290.470 2196.000 1290.750 2199.460 ;
        RECT 1301.510 2196.000 1301.790 2199.460 ;
        RECT 1313.010 2196.000 1313.290 2199.460 ;
        RECT 1324.510 2196.000 1324.790 2199.460 ;
        RECT 1335.550 2196.000 1335.830 2199.460 ;
        RECT 1347.050 2196.000 1347.330 2199.460 ;
        RECT 1358.550 2196.000 1358.830 2199.460 ;
        RECT 1369.590 2196.000 1369.870 2199.460 ;
        RECT 1381.090 2196.000 1381.370 2199.460 ;
        RECT 1392.130 2196.000 1392.410 2199.460 ;
        RECT 1403.630 2196.000 1403.910 2199.460 ;
        RECT 1415.130 2196.000 1415.410 2199.460 ;
        RECT 1426.170 2196.000 1426.450 2199.460 ;
        RECT 1437.670 2196.000 1437.950 2199.460 ;
        RECT 1448.710 2196.000 1448.990 2199.460 ;
        RECT 1460.210 2196.000 1460.490 2199.460 ;
        RECT 1471.710 2196.000 1471.990 2199.460 ;
        RECT 1482.750 2196.000 1483.030 2199.460 ;
        RECT 1494.250 2196.000 1494.530 2199.460 ;
      LAYER met2 ;
        RECT 305.160 2195.720 305.330 2196.000 ;
        RECT 306.170 2195.720 316.370 2196.000 ;
        RECT 317.210 2195.720 327.870 2196.000 ;
        RECT 328.710 2195.720 338.910 2196.000 ;
        RECT 339.750 2195.720 350.410 2196.000 ;
        RECT 351.250 2195.720 361.910 2196.000 ;
        RECT 362.750 2195.720 372.950 2196.000 ;
        RECT 373.790 2195.720 384.450 2196.000 ;
        RECT 385.290 2195.720 395.490 2196.000 ;
        RECT 396.330 2195.720 406.990 2196.000 ;
        RECT 407.830 2195.720 418.490 2196.000 ;
        RECT 419.330 2195.720 429.530 2196.000 ;
        RECT 430.370 2195.720 441.030 2196.000 ;
        RECT 441.870 2195.720 452.070 2196.000 ;
        RECT 452.910 2195.720 463.570 2196.000 ;
        RECT 464.410 2195.720 475.070 2196.000 ;
        RECT 475.910 2195.720 486.110 2196.000 ;
        RECT 486.950 2195.720 497.610 2196.000 ;
        RECT 498.450 2195.720 509.110 2196.000 ;
        RECT 509.950 2195.720 520.150 2196.000 ;
        RECT 520.990 2195.720 531.650 2196.000 ;
        RECT 532.490 2195.720 542.690 2196.000 ;
        RECT 543.530 2195.720 554.190 2196.000 ;
        RECT 555.030 2195.720 565.690 2196.000 ;
        RECT 566.530 2195.720 576.730 2196.000 ;
        RECT 577.570 2195.720 588.230 2196.000 ;
        RECT 589.070 2195.720 599.270 2196.000 ;
        RECT 600.110 2195.720 610.770 2196.000 ;
        RECT 611.610 2195.720 622.270 2196.000 ;
        RECT 623.110 2195.720 633.310 2196.000 ;
        RECT 634.150 2195.720 644.810 2196.000 ;
        RECT 645.650 2195.720 656.310 2196.000 ;
        RECT 657.150 2195.720 667.350 2196.000 ;
        RECT 668.190 2195.720 678.850 2196.000 ;
        RECT 679.690 2195.720 689.890 2196.000 ;
        RECT 690.730 2195.720 701.390 2196.000 ;
        RECT 702.230 2195.720 712.890 2196.000 ;
        RECT 713.730 2195.720 723.930 2196.000 ;
        RECT 724.770 2195.720 735.430 2196.000 ;
        RECT 736.270 2195.720 746.470 2196.000 ;
        RECT 747.310 2195.720 757.970 2196.000 ;
        RECT 758.810 2195.720 769.470 2196.000 ;
        RECT 770.310 2195.720 780.510 2196.000 ;
        RECT 781.350 2195.720 792.010 2196.000 ;
        RECT 792.850 2195.720 803.050 2196.000 ;
        RECT 803.890 2195.720 814.550 2196.000 ;
        RECT 815.390 2195.720 826.050 2196.000 ;
        RECT 826.890 2195.720 837.090 2196.000 ;
        RECT 837.930 2195.720 848.590 2196.000 ;
        RECT 849.430 2195.720 860.090 2196.000 ;
        RECT 860.930 2195.720 871.130 2196.000 ;
        RECT 871.970 2195.720 882.630 2196.000 ;
        RECT 883.470 2195.720 893.670 2196.000 ;
        RECT 894.510 2195.720 905.170 2196.000 ;
        RECT 906.010 2195.720 916.670 2196.000 ;
        RECT 917.510 2195.720 927.710 2196.000 ;
        RECT 928.550 2195.720 939.210 2196.000 ;
        RECT 940.050 2195.720 950.250 2196.000 ;
        RECT 951.090 2195.720 961.750 2196.000 ;
        RECT 962.590 2195.720 973.250 2196.000 ;
        RECT 974.090 2195.720 984.290 2196.000 ;
        RECT 985.130 2195.720 995.790 2196.000 ;
        RECT 996.630 2195.720 1007.290 2196.000 ;
        RECT 1008.130 2195.720 1018.330 2196.000 ;
        RECT 1019.170 2195.720 1029.830 2196.000 ;
        RECT 1030.670 2195.720 1040.870 2196.000 ;
        RECT 1041.710 2195.720 1052.370 2196.000 ;
        RECT 1053.210 2195.720 1063.870 2196.000 ;
        RECT 1064.710 2195.720 1074.910 2196.000 ;
        RECT 1075.750 2195.720 1086.410 2196.000 ;
        RECT 1087.250 2195.720 1097.450 2196.000 ;
        RECT 1098.290 2195.720 1108.950 2196.000 ;
        RECT 1109.790 2195.720 1120.450 2196.000 ;
        RECT 1121.290 2195.720 1131.490 2196.000 ;
        RECT 1132.330 2195.720 1142.990 2196.000 ;
        RECT 1143.830 2195.720 1154.030 2196.000 ;
        RECT 1154.870 2195.720 1165.530 2196.000 ;
        RECT 1166.370 2195.720 1177.030 2196.000 ;
        RECT 1177.870 2195.720 1188.070 2196.000 ;
        RECT 1188.910 2195.720 1199.570 2196.000 ;
        RECT 1200.410 2195.720 1211.070 2196.000 ;
        RECT 1211.910 2195.720 1222.110 2196.000 ;
        RECT 1222.950 2195.720 1233.610 2196.000 ;
        RECT 1234.450 2195.720 1244.650 2196.000 ;
        RECT 1245.490 2195.720 1256.150 2196.000 ;
        RECT 1256.990 2195.720 1267.650 2196.000 ;
        RECT 1268.490 2195.720 1278.690 2196.000 ;
        RECT 1279.530 2195.720 1290.190 2196.000 ;
        RECT 1291.030 2195.720 1301.230 2196.000 ;
        RECT 1302.070 2195.720 1312.730 2196.000 ;
        RECT 1313.570 2195.720 1324.230 2196.000 ;
        RECT 1325.070 2195.720 1335.270 2196.000 ;
        RECT 1336.110 2195.720 1346.770 2196.000 ;
        RECT 1347.610 2195.720 1358.270 2196.000 ;
        RECT 1359.110 2195.720 1369.310 2196.000 ;
        RECT 1370.150 2195.720 1380.810 2196.000 ;
        RECT 1381.650 2195.720 1391.850 2196.000 ;
        RECT 1392.690 2195.720 1403.350 2196.000 ;
        RECT 1404.190 2195.720 1414.850 2196.000 ;
        RECT 1415.690 2195.720 1425.890 2196.000 ;
        RECT 1426.730 2195.720 1437.390 2196.000 ;
        RECT 1438.230 2195.720 1448.430 2196.000 ;
        RECT 1449.270 2195.720 1459.930 2196.000 ;
        RECT 1460.770 2195.720 1471.430 2196.000 ;
        RECT 1472.270 2195.720 1482.470 2196.000 ;
        RECT 1483.310 2195.720 1493.970 2196.000 ;
        RECT 305.160 1004.280 1494.520 2195.720 ;
      LAYER met2 ;
        RECT 1511.260 1017.125 1511.400 2746.190 ;
        RECT 1529.130 2732.395 1529.410 2732.765 ;
        RECT 1522.240 2725.450 1522.500 2725.770 ;
        RECT 1521.780 2711.850 1522.040 2712.170 ;
        RECT 1521.320 2697.910 1521.580 2698.230 ;
        RECT 1514.420 2421.830 1514.680 2422.150 ;
        RECT 1514.480 2297.370 1514.620 2421.830 ;
        RECT 1514.880 2387.490 1515.140 2387.810 ;
        RECT 1514.940 2301.110 1515.080 2387.490 ;
        RECT 1514.880 2300.790 1515.140 2301.110 ;
        RECT 1514.940 2297.710 1515.080 2300.790 ;
        RECT 1514.880 2297.390 1515.140 2297.710 ;
        RECT 1514.420 2297.050 1514.680 2297.370 ;
        RECT 1513.960 2186.890 1514.220 2187.210 ;
        RECT 1514.020 2184.005 1514.160 2186.890 ;
        RECT 1513.950 2183.635 1514.230 2184.005 ;
        RECT 1513.960 2173.290 1514.220 2173.610 ;
        RECT 1514.020 2173.125 1514.160 2173.290 ;
        RECT 1513.950 2172.755 1514.230 2173.125 ;
        RECT 1513.960 2166.150 1514.220 2166.470 ;
        RECT 1514.020 2162.245 1514.160 2166.150 ;
        RECT 1513.950 2161.875 1514.230 2162.245 ;
        RECT 1513.960 2152.550 1514.220 2152.870 ;
        RECT 1514.020 2151.365 1514.160 2152.550 ;
        RECT 1513.950 2150.995 1514.230 2151.365 ;
        RECT 1513.960 2145.410 1514.220 2145.730 ;
        RECT 1514.020 2139.805 1514.160 2145.410 ;
        RECT 1513.950 2139.435 1514.230 2139.805 ;
        RECT 1513.960 2131.810 1514.220 2132.130 ;
        RECT 1514.020 2128.925 1514.160 2131.810 ;
        RECT 1513.950 2128.555 1514.230 2128.925 ;
        RECT 1513.960 2118.045 1514.220 2118.190 ;
        RECT 1513.950 2117.675 1514.230 2118.045 ;
        RECT 1513.960 2111.070 1514.220 2111.390 ;
        RECT 1514.020 2107.165 1514.160 2111.070 ;
        RECT 1513.950 2106.795 1514.230 2107.165 ;
        RECT 1513.960 2097.130 1514.220 2097.450 ;
        RECT 1514.020 2096.285 1514.160 2097.130 ;
        RECT 1513.950 2095.915 1514.230 2096.285 ;
        RECT 1513.960 2090.330 1514.220 2090.650 ;
        RECT 1514.020 2084.725 1514.160 2090.330 ;
        RECT 1513.950 2084.355 1514.230 2084.725 ;
        RECT 1513.960 2076.730 1514.220 2077.050 ;
        RECT 1514.020 2073.845 1514.160 2076.730 ;
        RECT 1513.950 2073.475 1514.230 2073.845 ;
        RECT 1513.960 2062.965 1514.220 2063.110 ;
        RECT 1513.950 2062.595 1514.230 2062.965 ;
        RECT 1513.960 2055.990 1514.220 2056.310 ;
        RECT 1514.020 2052.085 1514.160 2055.990 ;
        RECT 1513.950 2051.715 1514.230 2052.085 ;
        RECT 1513.960 2042.050 1514.220 2042.370 ;
        RECT 1514.020 2041.205 1514.160 2042.050 ;
        RECT 1513.950 2040.835 1514.230 2041.205 ;
        RECT 1513.960 2035.250 1514.220 2035.570 ;
        RECT 1514.020 2029.645 1514.160 2035.250 ;
        RECT 1513.950 2029.275 1514.230 2029.645 ;
        RECT 1513.500 2021.310 1513.760 2021.630 ;
        RECT 1513.560 2018.765 1513.700 2021.310 ;
        RECT 1513.490 2018.395 1513.770 2018.765 ;
        RECT 1513.960 2007.885 1514.220 2008.030 ;
        RECT 1513.950 2007.515 1514.230 2007.885 ;
        RECT 1513.960 2000.570 1514.220 2000.890 ;
        RECT 1514.020 1997.005 1514.160 2000.570 ;
        RECT 1513.950 1996.635 1514.230 1997.005 ;
        RECT 1513.960 1986.970 1514.220 1987.290 ;
        RECT 1514.020 1986.125 1514.160 1986.970 ;
        RECT 1513.950 1985.755 1514.230 1986.125 ;
        RECT 1512.580 1979.830 1512.840 1980.150 ;
        RECT 1512.640 1974.565 1512.780 1979.830 ;
        RECT 1512.570 1974.195 1512.850 1974.565 ;
        RECT 1513.500 1966.230 1513.760 1966.550 ;
        RECT 1513.560 1963.685 1513.700 1966.230 ;
        RECT 1513.490 1963.315 1513.770 1963.685 ;
        RECT 1513.950 1952.435 1514.230 1952.805 ;
        RECT 1513.960 1952.290 1514.220 1952.435 ;
        RECT 1513.960 1945.490 1514.220 1945.810 ;
        RECT 1514.020 1941.925 1514.160 1945.490 ;
        RECT 1513.950 1941.555 1514.230 1941.925 ;
        RECT 1512.580 1931.550 1512.840 1931.870 ;
        RECT 1512.640 1931.045 1512.780 1931.550 ;
        RECT 1512.570 1930.675 1512.850 1931.045 ;
        RECT 1512.580 1924.750 1512.840 1925.070 ;
        RECT 1512.640 1919.485 1512.780 1924.750 ;
        RECT 1512.570 1919.115 1512.850 1919.485 ;
        RECT 1513.960 1910.810 1514.220 1911.130 ;
        RECT 1514.020 1908.605 1514.160 1910.810 ;
        RECT 1513.950 1908.235 1514.230 1908.605 ;
        RECT 1513.040 1904.010 1513.300 1904.330 ;
        RECT 1513.100 1897.725 1513.240 1904.010 ;
        RECT 1513.030 1897.355 1513.310 1897.725 ;
        RECT 1513.960 1890.410 1514.220 1890.730 ;
        RECT 1514.020 1886.845 1514.160 1890.410 ;
        RECT 1513.950 1886.475 1514.230 1886.845 ;
        RECT 1513.960 1876.470 1514.220 1876.790 ;
        RECT 1514.020 1875.965 1514.160 1876.470 ;
        RECT 1513.950 1875.595 1514.230 1875.965 ;
        RECT 1513.960 1869.670 1514.220 1869.990 ;
        RECT 1514.020 1865.085 1514.160 1869.670 ;
        RECT 1513.950 1864.715 1514.230 1865.085 ;
        RECT 1511.660 1855.730 1511.920 1856.050 ;
        RECT 1511.720 1853.525 1511.860 1855.730 ;
        RECT 1511.650 1853.155 1511.930 1853.525 ;
        RECT 1513.040 1848.930 1513.300 1849.250 ;
        RECT 1513.100 1842.645 1513.240 1848.930 ;
        RECT 1513.030 1842.275 1513.310 1842.645 ;
        RECT 1513.960 1834.990 1514.220 1835.310 ;
        RECT 1514.020 1831.765 1514.160 1834.990 ;
        RECT 1513.950 1831.395 1514.230 1831.765 ;
        RECT 1512.580 1821.390 1512.840 1821.710 ;
        RECT 1512.640 1820.885 1512.780 1821.390 ;
        RECT 1512.570 1820.515 1512.850 1820.885 ;
        RECT 1512.120 1814.250 1512.380 1814.570 ;
        RECT 1512.180 1810.005 1512.320 1814.250 ;
        RECT 1512.110 1809.635 1512.390 1810.005 ;
        RECT 1511.660 1800.650 1511.920 1800.970 ;
        RECT 1511.720 1798.445 1511.860 1800.650 ;
        RECT 1511.650 1798.075 1511.930 1798.445 ;
        RECT 1512.580 1793.510 1512.840 1793.830 ;
        RECT 1512.640 1787.565 1512.780 1793.510 ;
        RECT 1512.570 1787.195 1512.850 1787.565 ;
        RECT 1513.960 1779.910 1514.220 1780.230 ;
        RECT 1514.020 1776.685 1514.160 1779.910 ;
        RECT 1513.950 1776.315 1514.230 1776.685 ;
        RECT 1513.960 1765.970 1514.220 1766.290 ;
        RECT 1514.020 1765.805 1514.160 1765.970 ;
        RECT 1513.950 1765.435 1514.230 1765.805 ;
        RECT 1512.120 1759.170 1512.380 1759.490 ;
        RECT 1512.180 1754.925 1512.320 1759.170 ;
        RECT 1512.110 1754.555 1512.390 1754.925 ;
        RECT 1513.500 1745.230 1513.760 1745.550 ;
        RECT 1513.560 1743.365 1513.700 1745.230 ;
        RECT 1513.490 1742.995 1513.770 1743.365 ;
        RECT 1512.580 1738.430 1512.840 1738.750 ;
        RECT 1512.640 1732.485 1512.780 1738.430 ;
        RECT 1512.570 1732.115 1512.850 1732.485 ;
        RECT 1513.960 1724.830 1514.220 1725.150 ;
        RECT 1514.020 1721.605 1514.160 1724.830 ;
        RECT 1513.950 1721.235 1514.230 1721.605 ;
        RECT 1513.960 1710.890 1514.220 1711.210 ;
        RECT 1514.020 1710.725 1514.160 1710.890 ;
        RECT 1513.950 1710.355 1514.230 1710.725 ;
        RECT 1512.120 1704.090 1512.380 1704.410 ;
        RECT 1512.180 1699.845 1512.320 1704.090 ;
        RECT 1512.110 1699.475 1512.390 1699.845 ;
        RECT 1513.500 1690.150 1513.760 1690.470 ;
        RECT 1513.560 1688.285 1513.700 1690.150 ;
        RECT 1513.490 1687.915 1513.770 1688.285 ;
        RECT 1512.580 1683.350 1512.840 1683.670 ;
        RECT 1512.640 1677.405 1512.780 1683.350 ;
        RECT 1512.570 1677.035 1512.850 1677.405 ;
        RECT 1513.960 1669.410 1514.220 1669.730 ;
        RECT 1514.020 1666.525 1514.160 1669.410 ;
        RECT 1513.950 1666.155 1514.230 1666.525 ;
        RECT 1512.580 1655.645 1512.840 1655.790 ;
        RECT 1512.570 1655.275 1512.850 1655.645 ;
        RECT 1511.660 1646.970 1511.920 1647.290 ;
        RECT 1511.720 1644.765 1511.860 1646.970 ;
        RECT 1511.650 1644.395 1511.930 1644.765 ;
        RECT 1512.580 1634.390 1512.840 1634.710 ;
        RECT 1512.640 1633.205 1512.780 1634.390 ;
        RECT 1512.570 1632.835 1512.850 1633.205 ;
        RECT 1511.660 1622.325 1511.920 1622.470 ;
        RECT 1511.650 1621.955 1511.930 1622.325 ;
        RECT 1511.660 1613.310 1511.920 1613.630 ;
        RECT 1511.720 1611.445 1511.860 1613.310 ;
        RECT 1511.650 1611.075 1511.930 1611.445 ;
        RECT 1511.660 1600.565 1511.920 1600.710 ;
        RECT 1511.650 1600.195 1511.930 1600.565 ;
        RECT 1513.500 1591.550 1513.760 1591.870 ;
        RECT 1513.560 1589.685 1513.700 1591.550 ;
        RECT 1513.490 1589.315 1513.770 1589.685 ;
        RECT 1513.960 1579.650 1514.220 1579.970 ;
        RECT 1514.020 1578.805 1514.160 1579.650 ;
        RECT 1513.950 1578.435 1514.230 1578.805 ;
        RECT 1513.960 1572.850 1514.220 1573.170 ;
        RECT 1514.020 1567.245 1514.160 1572.850 ;
        RECT 1513.950 1566.875 1514.230 1567.245 ;
        RECT 1513.500 1558.910 1513.760 1559.230 ;
        RECT 1513.560 1556.365 1513.700 1558.910 ;
        RECT 1513.490 1555.995 1513.770 1556.365 ;
        RECT 1513.960 1545.485 1514.220 1545.630 ;
        RECT 1513.950 1545.115 1514.230 1545.485 ;
        RECT 1513.960 1538.510 1514.220 1538.830 ;
        RECT 1514.020 1534.605 1514.160 1538.510 ;
        RECT 1513.950 1534.235 1514.230 1534.605 ;
        RECT 1513.960 1524.570 1514.220 1524.890 ;
        RECT 1514.020 1523.725 1514.160 1524.570 ;
        RECT 1513.950 1523.355 1514.230 1523.725 ;
        RECT 1513.960 1517.770 1514.220 1518.090 ;
        RECT 1514.020 1512.165 1514.160 1517.770 ;
        RECT 1513.950 1511.795 1514.230 1512.165 ;
        RECT 1513.500 1503.830 1513.760 1504.150 ;
        RECT 1513.560 1501.285 1513.700 1503.830 ;
        RECT 1513.490 1500.915 1513.770 1501.285 ;
        RECT 1513.960 1490.405 1514.220 1490.550 ;
        RECT 1513.950 1490.035 1514.230 1490.405 ;
        RECT 1513.040 1479.525 1513.300 1479.670 ;
        RECT 1513.030 1479.155 1513.310 1479.525 ;
        RECT 1513.960 1469.490 1514.220 1469.810 ;
        RECT 1514.020 1468.645 1514.160 1469.490 ;
        RECT 1513.950 1468.275 1514.230 1468.645 ;
        RECT 1512.580 1462.350 1512.840 1462.670 ;
        RECT 1512.640 1457.085 1512.780 1462.350 ;
        RECT 1512.570 1456.715 1512.850 1457.085 ;
        RECT 1513.500 1448.750 1513.760 1449.070 ;
        RECT 1513.560 1446.205 1513.700 1448.750 ;
        RECT 1513.490 1445.835 1513.770 1446.205 ;
        RECT 1513.950 1434.955 1514.230 1435.325 ;
        RECT 1513.960 1434.810 1514.220 1434.955 ;
        RECT 1513.500 1426.310 1513.760 1426.630 ;
        RECT 1513.560 1424.445 1513.700 1426.310 ;
        RECT 1513.490 1424.075 1513.770 1424.445 ;
        RECT 1512.580 1414.070 1512.840 1414.390 ;
        RECT 1512.640 1413.565 1512.780 1414.070 ;
        RECT 1512.570 1413.195 1512.850 1413.565 ;
        RECT 1512.580 1407.270 1512.840 1407.590 ;
        RECT 1512.640 1402.005 1512.780 1407.270 ;
        RECT 1512.570 1401.635 1512.850 1402.005 ;
        RECT 1511.660 1393.330 1511.920 1393.650 ;
        RECT 1511.720 1391.125 1511.860 1393.330 ;
        RECT 1511.650 1390.755 1511.930 1391.125 ;
        RECT 1513.040 1386.530 1513.300 1386.850 ;
        RECT 1513.100 1380.245 1513.240 1386.530 ;
        RECT 1513.030 1379.875 1513.310 1380.245 ;
        RECT 1513.960 1372.930 1514.220 1373.250 ;
        RECT 1514.020 1369.365 1514.160 1372.930 ;
        RECT 1513.950 1368.995 1514.230 1369.365 ;
        RECT 1512.580 1358.990 1512.840 1359.310 ;
        RECT 1512.640 1358.485 1512.780 1358.990 ;
        RECT 1512.570 1358.115 1512.850 1358.485 ;
        RECT 1512.580 1352.190 1512.840 1352.510 ;
        RECT 1512.640 1346.925 1512.780 1352.190 ;
        RECT 1512.570 1346.555 1512.850 1346.925 ;
        RECT 1511.660 1338.250 1511.920 1338.570 ;
        RECT 1511.720 1336.045 1511.860 1338.250 ;
        RECT 1511.650 1335.675 1511.930 1336.045 ;
        RECT 1513.040 1331.450 1513.300 1331.770 ;
        RECT 1513.100 1325.165 1513.240 1331.450 ;
        RECT 1513.030 1324.795 1513.310 1325.165 ;
        RECT 1513.960 1317.510 1514.220 1317.830 ;
        RECT 1514.020 1314.285 1514.160 1317.510 ;
        RECT 1513.950 1313.915 1514.230 1314.285 ;
        RECT 1512.580 1303.910 1512.840 1304.230 ;
        RECT 1512.640 1303.405 1512.780 1303.910 ;
        RECT 1512.570 1303.035 1512.850 1303.405 ;
        RECT 1512.120 1296.770 1512.380 1297.090 ;
        RECT 1512.180 1292.525 1512.320 1296.770 ;
        RECT 1512.110 1292.155 1512.390 1292.525 ;
        RECT 1511.660 1283.170 1511.920 1283.490 ;
        RECT 1511.720 1280.965 1511.860 1283.170 ;
        RECT 1511.650 1280.595 1511.930 1280.965 ;
        RECT 1512.580 1276.030 1512.840 1276.350 ;
        RECT 1512.640 1270.085 1512.780 1276.030 ;
        RECT 1512.570 1269.715 1512.850 1270.085 ;
        RECT 1513.960 1262.430 1514.220 1262.750 ;
        RECT 1514.020 1259.205 1514.160 1262.430 ;
        RECT 1513.950 1258.835 1514.230 1259.205 ;
        RECT 1513.960 1248.490 1514.220 1248.810 ;
        RECT 1514.020 1248.325 1514.160 1248.490 ;
        RECT 1513.950 1247.955 1514.230 1248.325 ;
        RECT 1512.120 1241.690 1512.380 1242.010 ;
        RECT 1512.180 1237.445 1512.320 1241.690 ;
        RECT 1512.110 1237.075 1512.390 1237.445 ;
        RECT 1513.500 1227.750 1513.760 1228.070 ;
        RECT 1513.560 1225.885 1513.700 1227.750 ;
        RECT 1513.490 1225.515 1513.770 1225.885 ;
        RECT 1512.580 1220.950 1512.840 1221.270 ;
        RECT 1512.640 1215.005 1512.780 1220.950 ;
        RECT 1512.570 1214.635 1512.850 1215.005 ;
        RECT 1513.960 1207.010 1514.220 1207.330 ;
        RECT 1514.020 1204.125 1514.160 1207.010 ;
        RECT 1513.950 1203.755 1514.230 1204.125 ;
        RECT 1513.960 1193.410 1514.220 1193.730 ;
        RECT 1514.020 1193.245 1514.160 1193.410 ;
        RECT 1513.950 1192.875 1514.230 1193.245 ;
        RECT 1512.120 1186.610 1512.380 1186.930 ;
        RECT 1512.180 1182.365 1512.320 1186.610 ;
        RECT 1512.110 1181.995 1512.390 1182.365 ;
        RECT 1513.500 1172.670 1513.760 1172.990 ;
        RECT 1513.560 1170.805 1513.700 1172.670 ;
        RECT 1513.490 1170.435 1513.770 1170.805 ;
        RECT 1512.580 1165.870 1512.840 1166.190 ;
        RECT 1512.640 1159.925 1512.780 1165.870 ;
        RECT 1512.570 1159.555 1512.850 1159.925 ;
        RECT 1513.960 1151.930 1514.220 1152.250 ;
        RECT 1514.020 1149.045 1514.160 1151.930 ;
        RECT 1513.950 1148.675 1514.230 1149.045 ;
        RECT 1513.960 1138.330 1514.220 1138.650 ;
        RECT 1514.020 1138.165 1514.160 1138.330 ;
        RECT 1513.950 1137.795 1514.230 1138.165 ;
        RECT 1513.960 1131.190 1514.220 1131.510 ;
        RECT 1514.020 1127.285 1514.160 1131.190 ;
        RECT 1513.950 1126.915 1514.230 1127.285 ;
        RECT 1513.500 1117.590 1513.760 1117.910 ;
        RECT 1513.560 1115.725 1513.700 1117.590 ;
        RECT 1513.490 1115.355 1513.770 1115.725 ;
        RECT 1513.960 1110.450 1514.220 1110.770 ;
        RECT 1514.020 1104.845 1514.160 1110.450 ;
        RECT 1513.950 1104.475 1514.230 1104.845 ;
        RECT 1513.960 1096.850 1514.220 1097.170 ;
        RECT 1514.020 1093.965 1514.160 1096.850 ;
        RECT 1513.950 1093.595 1514.230 1093.965 ;
        RECT 1513.960 1083.085 1514.220 1083.230 ;
        RECT 1513.950 1082.715 1514.230 1083.085 ;
        RECT 1513.960 1076.110 1514.220 1076.430 ;
        RECT 1514.020 1072.205 1514.160 1076.110 ;
        RECT 1513.950 1071.835 1514.230 1072.205 ;
        RECT 1513.040 1062.170 1513.300 1062.490 ;
        RECT 1513.100 1060.645 1513.240 1062.170 ;
        RECT 1513.030 1060.275 1513.310 1060.645 ;
        RECT 1513.960 1055.370 1514.220 1055.690 ;
        RECT 1514.020 1049.765 1514.160 1055.370 ;
        RECT 1513.950 1049.395 1514.230 1049.765 ;
        RECT 1513.960 1041.430 1514.220 1041.750 ;
        RECT 1514.020 1038.885 1514.160 1041.430 ;
        RECT 1513.950 1038.515 1514.230 1038.885 ;
        RECT 1513.960 1028.005 1514.220 1028.150 ;
        RECT 1513.950 1027.635 1514.230 1028.005 ;
        RECT 1511.190 1016.755 1511.470 1017.125 ;
        RECT 1514.480 1006.245 1514.620 2297.050 ;
        RECT 1514.940 2194.885 1515.080 2297.390 ;
        RECT 1514.870 2194.515 1515.150 2194.885 ;
        RECT 1521.380 1600.710 1521.520 2697.910 ;
        RECT 1521.840 1622.470 1521.980 2711.850 ;
        RECT 1522.300 1647.290 1522.440 2725.450 ;
        RECT 1528.670 2718.795 1528.950 2719.165 ;
        RECT 1528.210 2697.715 1528.490 2698.085 ;
        RECT 1522.240 1646.970 1522.500 1647.290 ;
        RECT 1521.780 1622.150 1522.040 1622.470 ;
        RECT 1528.280 1613.630 1528.420 2697.715 ;
        RECT 1528.740 1634.710 1528.880 2718.795 ;
        RECT 1529.200 1655.790 1529.340 2732.395 ;
        RECT 1538.330 2725.595 1538.610 2725.965 ;
        RECT 1538.340 2725.450 1538.600 2725.595 ;
        RECT 1536.030 2711.995 1536.310 2712.365 ;
        RECT 1536.040 2711.850 1536.300 2711.995 ;
        RECT 1536.490 2701.795 1536.770 2702.165 ;
        RECT 1536.560 2698.085 1536.700 2701.795 ;
        RECT 1538.330 2699.075 1538.610 2699.445 ;
        RECT 1538.400 2698.230 1538.540 2699.075 ;
        RECT 1536.490 2697.715 1536.770 2698.085 ;
        RECT 1538.340 2697.910 1538.600 2698.230 ;
        RECT 1535.110 2687.515 1535.390 2687.885 ;
        RECT 1529.590 2401.235 1529.870 2401.605 ;
        RECT 1529.140 1655.470 1529.400 1655.790 ;
        RECT 1528.680 1634.390 1528.940 1634.710 ;
        RECT 1528.220 1613.310 1528.480 1613.630 ;
        RECT 1521.320 1600.390 1521.580 1600.710 ;
        RECT 1529.660 1479.670 1529.800 2401.235 ;
        RECT 1535.180 1591.870 1535.320 2687.515 ;
        RECT 1535.570 2390.355 1535.850 2390.725 ;
        RECT 1535.640 2387.810 1535.780 2390.355 ;
        RECT 1535.580 2387.490 1535.840 2387.810 ;
      LAYER met2 ;
        RECT 1555.000 2305.000 1931.480 2751.235 ;
      LAYER met2 ;
        RECT 1945.960 2749.765 1946.100 2751.290 ;
        RECT 1945.890 2749.395 1946.170 2749.765 ;
        RECT 1946.880 2739.450 1947.020 2766.930 ;
        RECT 2539.360 2766.775 2539.500 2766.930 ;
        RECT 2594.490 2753.475 2594.770 2753.845 ;
        RECT 2582.080 2751.290 2582.340 2751.610 ;
        RECT 1945.960 2739.310 1947.020 2739.450 ;
        RECT 1942.220 2683.970 1942.480 2684.290 ;
        RECT 1759.130 2297.875 1759.410 2298.245 ;
        RECT 1639.530 2297.195 1639.810 2297.565 ;
        RECT 1607.790 2290.395 1608.070 2290.765 ;
        RECT 1614.690 2290.395 1614.970 2290.765 ;
        RECT 1628.490 2290.395 1628.770 2290.765 ;
        RECT 1635.390 2290.395 1635.670 2290.765 ;
        RECT 1587.090 2289.035 1587.370 2289.405 ;
        RECT 1548.920 2286.850 1549.180 2287.170 ;
        RECT 1542.020 2284.810 1542.280 2285.130 ;
        RECT 1535.120 1591.550 1535.380 1591.870 ;
        RECT 1529.600 1479.350 1529.860 1479.670 ;
        RECT 1542.080 1426.630 1542.220 2284.810 ;
        RECT 1542.020 1426.310 1542.280 1426.630 ;
        RECT 1548.980 1117.910 1549.120 2286.850 ;
        RECT 1562.720 2286.170 1562.980 2286.490 ;
        RECT 1548.920 1117.590 1549.180 1117.910 ;
        RECT 1562.780 1097.170 1562.920 2286.170 ;
        RECT 1576.520 2285.490 1576.780 2285.810 ;
        RECT 1562.720 1096.850 1562.980 1097.170 ;
        RECT 1576.580 1083.230 1576.720 2285.490 ;
        RECT 1587.160 2285.130 1587.300 2289.035 ;
        RECT 1587.100 2284.810 1587.360 2285.130 ;
        RECT 1601.350 2284.955 1601.630 2285.325 ;
        RECT 1580.190 2284.275 1580.470 2284.645 ;
        RECT 1593.990 2284.275 1594.270 2284.645 ;
        RECT 1600.890 2284.275 1601.170 2284.645 ;
        RECT 1580.260 1579.970 1580.400 2284.275 ;
        RECT 1583.420 2283.790 1583.680 2284.110 ;
        RECT 1580.200 1579.650 1580.460 1579.970 ;
        RECT 1576.520 1082.910 1576.780 1083.230 ;
        RECT 1583.480 1055.690 1583.620 2283.790 ;
        RECT 1594.060 1435.130 1594.200 2284.275 ;
        RECT 1600.960 1449.070 1601.100 2284.275 ;
        RECT 1601.420 1462.670 1601.560 2284.955 ;
        RECT 1601.360 1462.350 1601.620 1462.670 ;
        RECT 1600.900 1448.750 1601.160 1449.070 ;
        RECT 1594.000 1434.810 1594.260 1435.130 ;
        RECT 1583.420 1055.370 1583.680 1055.690 ;
        RECT 1607.860 1028.150 1608.000 2290.395 ;
        RECT 1611.010 2289.715 1611.290 2290.085 ;
        RECT 1611.080 2286.830 1611.220 2289.715 ;
        RECT 1611.020 2286.510 1611.280 2286.830 ;
        RECT 1611.080 1759.490 1611.220 2286.510 ;
        RECT 1611.020 1759.170 1611.280 1759.490 ;
        RECT 1614.760 1041.750 1614.900 2290.395 ;
        RECT 1617.910 2289.715 1618.190 2290.085 ;
        RECT 1617.980 2285.470 1618.120 2289.715 ;
        RECT 1624.810 2289.035 1625.090 2289.405 ;
        RECT 1621.590 2285.635 1621.870 2286.005 ;
        RECT 1617.920 2285.150 1618.180 2285.470 ;
        RECT 1617.460 2173.290 1617.720 2173.610 ;
        RECT 1617.520 2172.590 1617.660 2173.290 ;
        RECT 1617.460 2172.270 1617.720 2172.590 ;
        RECT 1617.980 1766.290 1618.120 2285.150 ;
        RECT 1621.660 2284.110 1621.800 2285.635 ;
        RECT 1624.880 2284.790 1625.020 2289.035 ;
        RECT 1624.820 2284.470 1625.080 2284.790 ;
        RECT 1621.600 2283.790 1621.860 2284.110 ;
        RECT 1624.880 1780.230 1625.020 2284.470 ;
        RECT 1624.820 1779.910 1625.080 1780.230 ;
        RECT 1617.920 1765.970 1618.180 1766.290 ;
        RECT 1628.560 1062.490 1628.700 2290.395 ;
        RECT 1631.710 2289.035 1631.990 2289.405 ;
        RECT 1631.780 2284.450 1631.920 2289.035 ;
        RECT 1631.720 2284.130 1631.980 2284.450 ;
        RECT 1631.780 1793.830 1631.920 2284.130 ;
        RECT 1631.720 1793.510 1631.980 1793.830 ;
        RECT 1635.460 1076.430 1635.600 2290.395 ;
        RECT 1639.600 2286.150 1639.740 2297.195 ;
        RECT 1676.800 2290.765 1677.060 2290.910 ;
        RECT 1723.720 2290.765 1723.980 2290.910 ;
        RECT 1645.510 2290.395 1645.790 2290.765 ;
        RECT 1649.650 2290.395 1649.930 2290.765 ;
        RECT 1659.310 2290.395 1659.590 2290.765 ;
        RECT 1665.750 2290.395 1666.030 2290.765 ;
        RECT 1670.350 2290.395 1670.630 2290.765 ;
        RECT 1676.790 2290.650 1677.070 2290.765 ;
        RECT 1676.790 2290.510 1677.460 2290.650 ;
        RECT 1676.790 2290.395 1677.070 2290.510 ;
        RECT 1645.520 2290.250 1645.780 2290.395 ;
        RECT 1639.540 2285.830 1639.800 2286.150 ;
        RECT 1639.600 2270.365 1639.740 2285.830 ;
        RECT 1642.290 2285.635 1642.570 2286.005 ;
        RECT 1642.300 2285.490 1642.560 2285.635 ;
        RECT 1638.610 2269.995 1638.890 2270.365 ;
        RECT 1639.530 2269.995 1639.810 2270.365 ;
        RECT 1638.680 2222.230 1638.820 2269.995 ;
        RECT 1638.160 2221.970 1638.420 2222.230 ;
        RECT 1637.760 2221.910 1638.420 2221.970 ;
        RECT 1638.620 2221.910 1638.880 2222.230 ;
        RECT 1637.760 2221.830 1638.360 2221.910 ;
        RECT 1637.760 2187.970 1637.900 2221.830 ;
        RECT 1637.760 2187.830 1638.360 2187.970 ;
        RECT 1638.220 2187.290 1638.360 2187.830 ;
        RECT 1637.760 2187.150 1638.360 2187.290 ;
        RECT 1637.760 2173.610 1637.900 2187.150 ;
        RECT 1637.700 2173.290 1637.960 2173.610 ;
        RECT 1638.160 2173.290 1638.420 2173.610 ;
        RECT 1638.620 2173.290 1638.880 2173.610 ;
        RECT 1638.220 2118.530 1638.360 2173.290 ;
        RECT 1638.680 2172.590 1638.820 2173.290 ;
        RECT 1638.620 2172.270 1638.880 2172.590 ;
        RECT 1637.700 2118.210 1637.960 2118.530 ;
        RECT 1638.160 2118.210 1638.420 2118.530 ;
        RECT 1637.760 2069.910 1637.900 2118.210 ;
        RECT 1637.700 2069.590 1637.960 2069.910 ;
        RECT 1638.620 2069.590 1638.880 2069.910 ;
        RECT 1638.680 2021.970 1638.820 2069.590 ;
        RECT 1637.700 2021.650 1637.960 2021.970 ;
        RECT 1638.620 2021.650 1638.880 2021.970 ;
        RECT 1637.760 1973.350 1637.900 2021.650 ;
        RECT 1637.700 1973.030 1637.960 1973.350 ;
        RECT 1638.160 1973.030 1638.420 1973.350 ;
        RECT 1638.220 1925.410 1638.360 1973.030 ;
        RECT 1638.160 1925.090 1638.420 1925.410 ;
        RECT 1639.080 1925.090 1639.340 1925.410 ;
        RECT 1639.140 1883.930 1639.280 1925.090 ;
        RECT 1638.160 1883.610 1638.420 1883.930 ;
        RECT 1639.080 1883.610 1639.340 1883.930 ;
        RECT 1638.220 1849.330 1638.360 1883.610 ;
        RECT 1638.220 1849.190 1639.280 1849.330 ;
        RECT 1639.140 1835.165 1639.280 1849.190 ;
        RECT 1639.070 1834.795 1639.350 1835.165 ;
        RECT 1640.450 1834.795 1640.730 1835.165 ;
        RECT 1640.520 1800.970 1640.660 1834.795 ;
        RECT 1645.580 1814.570 1645.720 2290.250 ;
        RECT 1646.430 2289.715 1646.710 2290.085 ;
        RECT 1646.500 2285.810 1646.640 2289.715 ;
        RECT 1649.190 2286.315 1649.470 2286.685 ;
        RECT 1649.200 2286.170 1649.460 2286.315 ;
        RECT 1646.440 2285.490 1646.700 2285.810 ;
        RECT 1646.500 1821.710 1646.640 2285.490 ;
        RECT 1646.440 1821.390 1646.700 1821.710 ;
        RECT 1645.520 1814.250 1645.780 1814.570 ;
        RECT 1640.460 1800.650 1640.720 1800.970 ;
        RECT 1649.720 1110.770 1649.860 2290.395 ;
        RECT 1659.380 2289.550 1659.520 2290.395 ;
        RECT 1652.410 2289.035 1652.690 2289.405 ;
        RECT 1656.560 2289.230 1656.820 2289.550 ;
        RECT 1659.320 2289.230 1659.580 2289.550 ;
        RECT 1652.480 2284.110 1652.620 2289.035 ;
        RECT 1656.090 2288.355 1656.370 2288.725 ;
        RECT 1656.160 2287.170 1656.300 2288.355 ;
        RECT 1656.100 2286.850 1656.360 2287.170 ;
        RECT 1656.620 2286.830 1656.760 2289.230 ;
        RECT 1665.820 2288.870 1665.960 2290.395 ;
        RECT 1663.000 2288.550 1663.260 2288.870 ;
        RECT 1665.760 2288.550 1666.020 2288.870 ;
        RECT 1656.560 2286.510 1656.820 2286.830 ;
        RECT 1663.060 2285.470 1663.200 2288.550 ;
        RECT 1670.420 2287.850 1670.560 2290.395 ;
        RECT 1670.360 2287.530 1670.620 2287.850 ;
        RECT 1663.000 2285.150 1663.260 2285.470 ;
        RECT 1670.420 2284.790 1670.560 2287.530 ;
        RECT 1676.790 2285.635 1677.070 2286.005 ;
        RECT 1662.990 2284.275 1663.270 2284.645 ;
        RECT 1669.890 2284.275 1670.170 2284.645 ;
        RECT 1670.360 2284.470 1670.620 2284.790 ;
        RECT 1652.420 2283.790 1652.680 2284.110 ;
        RECT 1652.480 1835.310 1652.620 2283.790 ;
        RECT 1652.420 1834.990 1652.680 1835.310 ;
        RECT 1663.060 1131.510 1663.200 2284.275 ;
        RECT 1669.960 1138.650 1670.100 2284.275 ;
        RECT 1676.860 1152.250 1677.000 2285.635 ;
        RECT 1677.320 2284.450 1677.460 2290.510 ;
        RECT 1682.770 2290.395 1683.050 2290.765 ;
        RECT 1690.130 2290.395 1690.410 2290.765 ;
        RECT 1695.190 2290.395 1695.470 2290.765 ;
        RECT 1699.330 2290.395 1699.610 2290.765 ;
        RECT 1706.230 2290.395 1706.510 2290.765 ;
        RECT 1711.290 2290.395 1711.570 2290.765 ;
        RECT 1718.190 2290.395 1718.470 2290.765 ;
        RECT 1682.840 2289.890 1682.980 2290.395 ;
        RECT 1690.140 2290.250 1690.400 2290.395 ;
        RECT 1682.780 2289.570 1683.040 2289.890 ;
        RECT 1682.840 2286.150 1682.980 2289.570 ;
        RECT 1690.200 2288.530 1690.340 2290.250 ;
        RECT 1695.260 2289.210 1695.400 2290.395 ;
        RECT 1695.200 2288.890 1695.460 2289.210 ;
        RECT 1690.140 2288.210 1690.400 2288.530 ;
        RECT 1682.780 2285.830 1683.040 2286.150 ;
        RECT 1695.260 2285.810 1695.400 2288.890 ;
        RECT 1699.400 2288.190 1699.540 2290.395 ;
        RECT 1706.300 2289.550 1706.440 2290.395 ;
        RECT 1706.240 2289.230 1706.500 2289.550 ;
        RECT 1704.400 2288.890 1704.660 2289.210 ;
        RECT 1699.340 2287.870 1699.600 2288.190 ;
        RECT 1695.200 2285.490 1695.460 2285.810 ;
        RECT 1684.150 2284.955 1684.430 2285.325 ;
        RECT 1677.260 2284.130 1677.520 2284.450 ;
        RECT 1683.690 2284.275 1683.970 2284.645 ;
        RECT 1683.760 1166.190 1683.900 2284.275 ;
        RECT 1684.220 1172.990 1684.360 2284.955 ;
        RECT 1690.590 2284.275 1690.870 2284.645 ;
        RECT 1697.490 2284.275 1697.770 2284.645 ;
        RECT 1690.660 1186.930 1690.800 2284.275 ;
        RECT 1697.560 1193.730 1697.700 2284.275 ;
        RECT 1699.400 2284.110 1699.540 2287.870 ;
        RECT 1704.460 2287.170 1704.600 2288.890 ;
        RECT 1704.400 2286.850 1704.660 2287.170 ;
        RECT 1704.390 2285.635 1704.670 2286.005 ;
        RECT 1699.340 2283.790 1699.600 2284.110 ;
        RECT 1704.460 1207.330 1704.600 2285.635 ;
        RECT 1711.360 1221.270 1711.500 2290.395 ;
        RECT 1712.670 2289.715 1712.950 2290.085 ;
        RECT 1717.740 2289.910 1718.000 2290.230 ;
        RECT 1712.740 2288.870 1712.880 2289.715 ;
        RECT 1717.800 2288.870 1717.940 2289.910 ;
        RECT 1712.680 2288.550 1712.940 2288.870 ;
        RECT 1717.740 2288.550 1718.000 2288.870 ;
        RECT 1714.520 2286.510 1714.780 2286.830 ;
        RECT 1714.580 1856.050 1714.720 2286.510 ;
        RECT 1714.520 1855.730 1714.780 1856.050 ;
        RECT 1718.260 1228.070 1718.400 2290.395 ;
        RECT 1721.880 2290.250 1722.140 2290.570 ;
        RECT 1723.710 2290.395 1723.990 2290.765 ;
        RECT 1725.090 2290.395 1725.370 2290.765 ;
        RECT 1731.990 2290.395 1732.270 2290.765 ;
        RECT 1738.890 2290.395 1739.170 2290.765 ;
        RECT 1745.790 2290.395 1746.070 2290.765 ;
        RECT 1721.940 2290.085 1722.080 2290.250 ;
        RECT 1721.870 2289.715 1722.150 2290.085 ;
        RECT 1718.650 2288.355 1718.930 2288.725 ;
        RECT 1718.720 1242.010 1718.860 2288.355 ;
        RECT 1721.940 2287.850 1722.080 2289.715 ;
        RECT 1721.880 2287.530 1722.140 2287.850 ;
        RECT 1725.160 1248.810 1725.300 2290.395 ;
        RECT 1729.690 2289.715 1729.970 2290.085 ;
        RECT 1729.700 2289.570 1729.960 2289.715 ;
        RECT 1732.060 1262.750 1732.200 2290.395 ;
        RECT 1734.290 2289.715 1734.570 2290.085 ;
        RECT 1734.360 2288.530 1734.500 2289.715 ;
        RECT 1734.300 2288.210 1734.560 2288.530 ;
        RECT 1735.220 2284.810 1735.480 2285.130 ;
        RECT 1735.280 2077.050 1735.420 2284.810 ;
        RECT 1735.220 2076.730 1735.480 2077.050 ;
        RECT 1738.960 1276.350 1739.100 2290.395 ;
        RECT 1741.190 2289.715 1741.470 2290.085 ;
        RECT 1741.260 2287.170 1741.400 2289.715 ;
        RECT 1741.200 2286.850 1741.460 2287.170 ;
        RECT 1745.860 1283.490 1746.000 2290.395 ;
        RECT 1759.200 2290.230 1759.340 2297.875 ;
        RECT 1794.090 2297.195 1794.370 2297.565 ;
        RECT 1766.500 2290.765 1766.760 2290.910 ;
        RECT 1759.590 2290.395 1759.870 2290.765 ;
        RECT 1759.600 2290.250 1759.860 2290.395 ;
        RECT 1763.740 2290.250 1764.000 2290.570 ;
        RECT 1766.490 2290.395 1766.770 2290.765 ;
        RECT 1770.180 2290.590 1770.440 2290.910 ;
        RECT 1746.250 2289.715 1746.530 2290.085 ;
        RECT 1752.690 2289.715 1752.970 2290.085 ;
        RECT 1759.140 2289.910 1759.400 2290.230 ;
        RECT 1746.320 2288.870 1746.460 2289.715 ;
        RECT 1752.760 2289.550 1752.900 2289.715 ;
        RECT 1752.700 2289.230 1752.960 2289.550 ;
        RECT 1753.160 2289.230 1753.420 2289.550 ;
        RECT 1746.260 2288.550 1746.520 2288.870 ;
        RECT 1748.560 2288.550 1748.820 2288.870 ;
        RECT 1746.320 2288.190 1746.460 2288.550 ;
        RECT 1746.260 2287.870 1746.520 2288.190 ;
        RECT 1748.620 2287.170 1748.760 2288.550 ;
        RECT 1753.220 2288.190 1753.360 2289.230 ;
        RECT 1753.160 2287.870 1753.420 2288.190 ;
        RECT 1748.560 2286.850 1748.820 2287.170 ;
        RECT 1749.020 2286.170 1749.280 2286.490 ;
        RECT 1749.080 2090.650 1749.220 2286.170 ;
        RECT 1755.920 2285.830 1756.180 2286.150 ;
        RECT 1752.690 2284.275 1752.970 2284.645 ;
        RECT 1749.020 2090.330 1749.280 2090.650 ;
        RECT 1752.760 1297.090 1752.900 2284.275 ;
        RECT 1755.980 2097.450 1756.120 2285.830 ;
        RECT 1762.820 2285.490 1763.080 2285.810 ;
        RECT 1760.050 2284.955 1760.330 2285.325 ;
        RECT 1759.590 2284.275 1759.870 2284.645 ;
        RECT 1755.920 2097.130 1756.180 2097.450 ;
        RECT 1759.660 1304.230 1759.800 2284.275 ;
        RECT 1760.120 1317.830 1760.260 2284.955 ;
        RECT 1762.880 2111.390 1763.020 2285.490 ;
        RECT 1763.280 2285.150 1763.540 2285.470 ;
        RECT 1763.340 2118.190 1763.480 2285.150 ;
        RECT 1763.800 2132.130 1763.940 2290.250 ;
        RECT 1769.720 2289.910 1769.980 2290.230 ;
        RECT 1768.340 2289.570 1768.600 2289.890 ;
        RECT 1768.400 2287.850 1768.540 2289.570 ;
        RECT 1768.340 2287.530 1768.600 2287.850 ;
        RECT 1766.490 2285.635 1766.770 2286.005 ;
        RECT 1763.740 2131.810 1764.000 2132.130 ;
        RECT 1763.280 2117.870 1763.540 2118.190 ;
        RECT 1762.820 2111.070 1763.080 2111.390 ;
        RECT 1766.560 1331.770 1766.700 2285.635 ;
        RECT 1769.780 2145.730 1769.920 2289.910 ;
        RECT 1770.240 2152.870 1770.380 2290.590 ;
        RECT 1780.290 2289.715 1780.570 2290.085 ;
        RECT 1780.360 2289.550 1780.500 2289.715 ;
        RECT 1775.230 2289.035 1775.510 2289.405 ;
        RECT 1780.300 2289.230 1780.560 2289.550 ;
        RECT 1775.300 2287.850 1775.440 2289.035 ;
        RECT 1787.190 2288.355 1787.470 2288.725 ;
        RECT 1787.200 2288.210 1787.460 2288.355 ;
        RECT 1794.160 2288.190 1794.300 2297.195 ;
        RECT 1797.320 2288.210 1797.580 2288.530 ;
        RECT 1794.100 2287.870 1794.360 2288.190 ;
        RECT 1775.240 2287.530 1775.500 2287.850 ;
        RECT 1790.420 2287.530 1790.680 2287.850 ;
        RECT 1776.620 2286.850 1776.880 2287.170 ;
        RECT 1773.390 2284.275 1773.670 2284.645 ;
        RECT 1770.180 2152.550 1770.440 2152.870 ;
        RECT 1769.720 2145.410 1769.980 2145.730 ;
        RECT 1773.460 1338.570 1773.600 2284.275 ;
        RECT 1776.680 1869.990 1776.820 2286.850 ;
        RECT 1780.290 2284.275 1780.570 2284.645 ;
        RECT 1776.620 1869.670 1776.880 1869.990 ;
        RECT 1780.360 1352.510 1780.500 2284.275 ;
        RECT 1783.520 2284.130 1783.780 2284.450 ;
        RECT 1787.190 2284.275 1787.470 2284.645 ;
        RECT 1783.580 1876.790 1783.720 2284.130 ;
        RECT 1783.520 1876.470 1783.780 1876.790 ;
        RECT 1787.260 1359.310 1787.400 2284.275 ;
        RECT 1790.480 1890.730 1790.620 2287.530 ;
        RECT 1794.090 2284.275 1794.370 2284.645 ;
        RECT 1790.420 1890.410 1790.680 1890.730 ;
        RECT 1794.160 1373.250 1794.300 2284.275 ;
        RECT 1797.380 1904.330 1797.520 2288.210 ;
        RECT 1797.320 1904.010 1797.580 1904.330 ;
        RECT 1942.280 1504.150 1942.420 2683.970 ;
        RECT 1945.960 2447.845 1946.100 2739.310 ;
        RECT 1997.420 2732.250 1997.680 2732.570 ;
        RECT 2187.390 2732.395 2187.670 2732.765 ;
        RECT 2187.400 2732.250 2187.660 2732.395 ;
        RECT 1990.520 2725.450 1990.780 2725.770 ;
        RECT 1976.720 2718.650 1976.980 2718.970 ;
        RECT 1969.820 2711.850 1970.080 2712.170 ;
        RECT 1962.920 2698.250 1963.180 2698.570 ;
        RECT 1956.020 2697.910 1956.280 2698.230 ;
        RECT 1945.890 2447.475 1946.170 2447.845 ;
        RECT 1945.890 2404.635 1946.170 2405.005 ;
        RECT 1945.960 2297.370 1946.100 2404.635 ;
        RECT 1945.900 2297.050 1946.160 2297.370 ;
        RECT 1956.080 1518.090 1956.220 2697.910 ;
        RECT 1962.980 1524.890 1963.120 2698.250 ;
        RECT 1969.880 1538.830 1970.020 2711.850 ;
        RECT 1976.780 1545.630 1976.920 2718.650 ;
        RECT 1990.580 1559.230 1990.720 2725.450 ;
        RECT 1997.480 1573.170 1997.620 2732.250 ;
        RECT 2187.390 2725.595 2187.670 2725.965 ;
        RECT 2187.400 2725.450 2187.660 2725.595 ;
        RECT 2187.390 2718.795 2187.670 2719.165 ;
        RECT 2187.400 2718.650 2187.660 2718.795 ;
        RECT 2187.390 2711.995 2187.670 2712.365 ;
        RECT 2187.400 2711.850 2187.660 2711.995 ;
        RECT 2187.850 2701.795 2188.130 2702.165 ;
        RECT 2187.390 2699.075 2187.670 2699.445 ;
        RECT 2187.460 2698.230 2187.600 2699.075 ;
        RECT 2187.920 2698.570 2188.060 2701.795 ;
        RECT 2187.860 2698.250 2188.120 2698.570 ;
        RECT 2187.400 2697.910 2187.660 2698.230 ;
        RECT 2187.390 2687.515 2187.670 2687.885 ;
        RECT 2187.460 2684.290 2187.600 2687.515 ;
        RECT 2187.400 2683.970 2187.660 2684.290 ;
        RECT 2011.220 2401.090 2011.480 2401.410 ;
        RECT 2187.390 2401.235 2187.670 2401.605 ;
        RECT 2187.400 2401.090 2187.660 2401.235 ;
        RECT 1997.420 1572.850 1997.680 1573.170 ;
        RECT 1990.520 1558.910 1990.780 1559.230 ;
        RECT 1976.720 1545.310 1976.980 1545.630 ;
        RECT 1969.820 1538.510 1970.080 1538.830 ;
        RECT 1962.920 1524.570 1963.180 1524.890 ;
        RECT 1956.020 1517.770 1956.280 1518.090 ;
        RECT 1942.220 1503.830 1942.480 1504.150 ;
        RECT 2011.280 1469.810 2011.420 2401.090 ;
        RECT 2190.610 2389.675 2190.890 2390.045 ;
        RECT 2190.680 2297.710 2190.820 2389.675 ;
      LAYER met2 ;
        RECT 2205.000 2305.000 2581.480 2751.235 ;
      LAYER met2 ;
        RECT 2582.140 2749.765 2582.280 2751.290 ;
        RECT 2582.070 2749.395 2582.350 2749.765 ;
        RECT 2594.560 2447.845 2594.700 2753.475 ;
        RECT 2594.490 2447.475 2594.770 2447.845 ;
        RECT 2190.620 2297.390 2190.880 2297.710 ;
        RECT 2415.090 2297.450 2415.370 2297.565 ;
        RECT 2415.090 2297.310 2415.760 2297.450 ;
        RECT 2415.090 2297.195 2415.370 2297.310 ;
        RECT 2308.830 2290.395 2309.110 2290.765 ;
        RECT 2315.270 2290.395 2315.550 2290.765 ;
        RECT 2324.930 2290.395 2325.210 2290.765 ;
        RECT 2325.850 2290.395 2326.130 2290.765 ;
        RECT 2343.790 2290.395 2344.070 2290.765 ;
        RECT 2349.770 2290.395 2350.050 2290.765 ;
        RECT 2358.970 2290.395 2359.250 2290.765 ;
        RECT 2361.270 2290.395 2361.550 2290.765 ;
        RECT 2367.250 2290.395 2367.530 2290.765 ;
        RECT 2374.150 2290.395 2374.430 2290.765 ;
        RECT 2377.370 2290.395 2377.650 2290.765 ;
        RECT 2384.730 2290.395 2385.010 2290.765 ;
        RECT 2391.630 2290.395 2391.910 2290.765 ;
        RECT 2397.150 2290.395 2397.430 2290.765 ;
        RECT 2415.090 2290.395 2415.370 2290.765 ;
        RECT 2301.010 2289.715 2301.290 2290.085 ;
        RECT 2301.080 2289.550 2301.220 2289.715 ;
        RECT 2290.890 2289.035 2291.170 2289.405 ;
        RECT 2301.020 2289.230 2301.280 2289.550 ;
        RECT 2267.440 2288.550 2267.700 2288.870 ;
        RECT 2266.520 2287.870 2266.780 2288.190 ;
        RECT 2218.220 2287.190 2218.480 2287.510 ;
        RECT 2218.280 1911.130 2218.420 2287.190 ;
        RECT 2263.290 2286.995 2263.570 2287.365 ;
        RECT 2263.360 2286.830 2263.500 2286.995 ;
        RECT 2263.300 2286.510 2263.560 2286.830 ;
        RECT 2252.710 2285.635 2252.990 2286.005 ;
        RECT 2232.010 2284.955 2232.290 2285.325 ;
        RECT 2228.790 2284.275 2229.070 2284.645 ;
        RECT 2218.220 1910.810 2218.480 1911.130 ;
        RECT 2228.860 1490.550 2229.000 2284.275 ;
        RECT 2228.800 1490.230 2229.060 1490.550 ;
        RECT 2011.220 1469.490 2011.480 1469.810 ;
        RECT 2232.080 1386.850 2232.220 2284.955 ;
        RECT 2238.910 2284.275 2239.190 2284.645 ;
        RECT 2245.810 2284.275 2246.090 2284.645 ;
        RECT 2238.980 1393.650 2239.120 2284.275 ;
        RECT 2245.880 1407.590 2246.020 2284.275 ;
        RECT 2252.780 1414.390 2252.920 2285.635 ;
        RECT 2266.580 2284.645 2266.720 2287.870 ;
        RECT 2267.500 2284.645 2267.640 2288.550 ;
        RECT 2290.960 2288.530 2291.100 2289.035 ;
        RECT 2290.900 2288.210 2291.160 2288.530 ;
        RECT 2283.990 2287.675 2284.270 2288.045 ;
        RECT 2297.790 2287.675 2298.070 2288.045 ;
        RECT 2284.000 2287.530 2284.260 2287.675 ;
        RECT 2297.860 2287.510 2298.000 2287.675 ;
        RECT 2270.190 2286.995 2270.470 2287.365 ;
        RECT 2297.800 2287.190 2298.060 2287.510 ;
        RECT 2270.200 2286.850 2270.460 2286.995 ;
        RECT 2273.420 2286.850 2273.680 2287.170 ;
        RECT 2273.480 2286.005 2273.620 2286.850 ;
        RECT 2273.410 2285.635 2273.690 2286.005 ;
        RECT 2294.110 2285.635 2294.390 2286.005 ;
        RECT 2296.870 2285.635 2297.150 2286.005 ;
        RECT 2263.750 2284.275 2264.030 2284.645 ;
        RECT 2266.510 2284.275 2266.790 2284.645 ;
        RECT 2267.430 2284.275 2267.710 2284.645 ;
        RECT 2263.820 1849.250 2263.960 2284.275 ;
        RECT 2263.760 1848.930 2264.020 1849.250 ;
        RECT 2266.580 1669.730 2266.720 2284.275 ;
        RECT 2267.500 1683.670 2267.640 2284.275 ;
        RECT 2273.480 1690.470 2273.620 2285.635 ;
        RECT 2280.310 2284.955 2280.590 2285.325 ;
        RECT 2283.530 2284.955 2283.810 2285.325 ;
        RECT 2277.090 2284.275 2277.370 2284.645 ;
        RECT 2277.100 2284.130 2277.360 2284.275 ;
        RECT 2280.380 1704.410 2280.520 2284.955 ;
        RECT 2283.600 2284.450 2283.740 2284.955 ;
        RECT 2283.540 2284.130 2283.800 2284.450 ;
        RECT 2287.210 2284.275 2287.490 2284.645 ;
        RECT 2290.430 2284.275 2290.710 2284.645 ;
        RECT 2287.280 1711.210 2287.420 2284.275 ;
        RECT 2290.500 2284.110 2290.640 2284.275 ;
        RECT 2290.440 2283.790 2290.700 2284.110 ;
        RECT 2294.180 1725.150 2294.320 2285.635 ;
        RECT 2296.940 2284.790 2297.080 2285.635 ;
        RECT 2296.880 2284.470 2297.140 2284.790 ;
        RECT 2301.080 1738.750 2301.220 2289.230 ;
        RECT 2301.930 2288.355 2302.210 2288.725 ;
        RECT 2301.940 2288.210 2302.200 2288.355 ;
        RECT 2302.000 1745.550 2302.140 2288.210 ;
        RECT 2308.900 2288.190 2309.040 2290.395 ;
        RECT 2315.340 2288.870 2315.480 2290.395 ;
        RECT 2325.000 2289.210 2325.140 2290.395 ;
        RECT 2324.940 2288.890 2325.200 2289.210 ;
        RECT 2315.280 2288.550 2315.540 2288.870 ;
        RECT 2308.840 2287.870 2309.100 2288.190 ;
        RECT 2325.000 2287.170 2325.140 2288.890 ;
        RECT 2325.920 2287.850 2326.060 2290.395 ;
        RECT 2340.110 2289.715 2340.390 2290.085 ;
        RECT 2333.210 2289.035 2333.490 2289.405 ;
        RECT 2325.860 2287.530 2326.120 2287.850 ;
        RECT 2324.940 2286.850 2325.200 2287.170 ;
        RECT 2321.720 2286.510 2321.980 2286.830 ;
        RECT 2305.150 2285.635 2305.430 2286.005 ;
        RECT 2304.690 2284.275 2304.970 2284.645 ;
        RECT 2304.760 1925.070 2304.900 2284.275 ;
        RECT 2305.220 1931.870 2305.360 2285.635 ;
        RECT 2311.590 2284.275 2311.870 2284.645 ;
        RECT 2318.490 2284.275 2318.770 2284.645 ;
        RECT 2311.660 1945.810 2311.800 2284.275 ;
        RECT 2318.560 1952.610 2318.700 2284.275 ;
        RECT 2321.780 2166.470 2321.920 2286.510 ;
        RECT 2325.390 2284.275 2325.670 2284.645 ;
        RECT 2325.920 2284.450 2326.060 2287.530 ;
        RECT 2328.620 2287.190 2328.880 2287.510 ;
        RECT 2321.720 2166.150 2321.980 2166.470 ;
        RECT 2325.460 1966.550 2325.600 2284.275 ;
        RECT 2325.860 2284.130 2326.120 2284.450 ;
        RECT 2328.680 2173.610 2328.820 2287.190 ;
        RECT 2332.290 2284.275 2332.570 2284.645 ;
        RECT 2333.280 2284.450 2333.420 2289.035 ;
        RECT 2335.520 2286.850 2335.780 2287.170 ;
        RECT 2328.620 2173.290 2328.880 2173.610 ;
        RECT 2332.360 1980.150 2332.500 2284.275 ;
        RECT 2333.220 2284.130 2333.480 2284.450 ;
        RECT 2335.580 2187.210 2335.720 2286.850 ;
        RECT 2339.650 2285.635 2339.930 2286.005 ;
        RECT 2339.190 2284.275 2339.470 2284.645 ;
        RECT 2335.520 2186.890 2335.780 2187.210 ;
        RECT 2339.260 1987.290 2339.400 2284.275 ;
        RECT 2339.720 2000.890 2339.860 2285.635 ;
        RECT 2340.180 2284.790 2340.320 2289.715 ;
        RECT 2343.860 2289.550 2344.000 2290.395 ;
        RECT 2343.800 2289.230 2344.060 2289.550 ;
        RECT 2349.840 2288.530 2349.980 2290.395 ;
        RECT 2359.040 2289.890 2359.180 2290.395 ;
        RECT 2358.980 2289.570 2359.240 2289.890 ;
        RECT 2355.820 2289.210 2357.800 2289.290 ;
        RECT 2355.820 2289.150 2357.860 2289.210 ;
        RECT 2349.780 2288.210 2350.040 2288.530 ;
        RECT 2340.120 2284.470 2340.380 2284.790 ;
        RECT 2346.090 2284.275 2346.370 2284.645 ;
        RECT 2352.990 2284.275 2353.270 2284.645 ;
        RECT 2355.820 2284.450 2355.960 2289.150 ;
        RECT 2357.600 2288.890 2357.860 2289.150 ;
        RECT 2356.680 2288.550 2356.940 2288.870 ;
        RECT 2356.740 2287.850 2356.880 2288.550 ;
        RECT 2359.040 2288.190 2359.180 2289.570 ;
        RECT 2361.340 2288.190 2361.480 2290.395 ;
        RECT 2367.320 2288.870 2367.460 2290.395 ;
        RECT 2367.260 2288.550 2367.520 2288.870 ;
        RECT 2358.980 2287.870 2359.240 2288.190 ;
        RECT 2361.280 2287.870 2361.540 2288.190 ;
        RECT 2356.220 2287.530 2356.480 2287.850 ;
        RECT 2356.680 2287.530 2356.940 2287.850 ;
        RECT 2356.280 2284.450 2356.420 2287.530 ;
        RECT 2359.890 2285.635 2360.170 2286.005 ;
        RECT 2346.160 2008.030 2346.300 2284.275 ;
        RECT 2353.060 2021.630 2353.200 2284.275 ;
        RECT 2355.760 2284.130 2356.020 2284.450 ;
        RECT 2356.220 2284.130 2356.480 2284.450 ;
        RECT 2359.960 2035.570 2360.100 2285.635 ;
        RECT 2366.790 2284.275 2367.070 2284.645 ;
        RECT 2373.690 2284.275 2373.970 2284.645 ;
        RECT 2374.220 2284.450 2374.360 2290.395 ;
        RECT 2377.440 2289.210 2377.580 2290.395 ;
        RECT 2377.380 2288.890 2377.640 2289.210 ;
        RECT 2384.800 2287.850 2384.940 2290.395 ;
        RECT 2391.700 2289.550 2391.840 2290.395 ;
        RECT 2391.640 2289.230 2391.900 2289.550 ;
        RECT 2394.390 2289.035 2394.670 2289.405 ;
        RECT 2381.520 2287.530 2381.780 2287.850 ;
        RECT 2384.740 2287.530 2385.000 2287.850 ;
        RECT 2380.590 2286.315 2380.870 2286.685 ;
        RECT 2380.660 2285.130 2380.800 2286.315 ;
        RECT 2381.050 2285.635 2381.330 2286.005 ;
        RECT 2380.600 2284.810 2380.860 2285.130 ;
        RECT 2366.860 2042.370 2367.000 2284.275 ;
        RECT 2373.760 2056.310 2373.900 2284.275 ;
        RECT 2374.160 2284.130 2374.420 2284.450 ;
        RECT 2381.120 2063.110 2381.260 2285.635 ;
        RECT 2381.580 2284.790 2381.720 2287.530 ;
        RECT 2387.490 2286.315 2387.770 2286.685 ;
        RECT 2387.500 2286.170 2387.760 2286.315 ;
        RECT 2394.460 2286.150 2394.600 2289.035 ;
        RECT 2397.220 2288.530 2397.360 2290.395 ;
        RECT 2415.100 2290.250 2415.360 2290.395 ;
        RECT 2402.210 2289.715 2402.490 2290.085 ;
        RECT 2402.220 2289.570 2402.480 2289.715 ;
        RECT 2402.670 2289.035 2402.950 2289.405 ;
        RECT 2401.300 2288.550 2401.560 2288.870 ;
        RECT 2397.160 2288.210 2397.420 2288.530 ;
        RECT 2401.360 2286.490 2401.500 2288.550 ;
        RECT 2401.300 2286.170 2401.560 2286.490 ;
        RECT 2394.400 2285.830 2394.660 2286.150 ;
        RECT 2402.740 2285.810 2402.880 2289.035 ;
        RECT 2408.190 2288.355 2408.470 2288.725 ;
        RECT 2408.260 2288.190 2408.400 2288.355 ;
        RECT 2408.200 2287.870 2408.460 2288.190 ;
        RECT 2415.090 2286.995 2415.370 2287.365 ;
        RECT 2402.680 2285.490 2402.940 2285.810 ;
        RECT 2408.190 2285.635 2408.470 2286.005 ;
        RECT 2408.260 2285.470 2408.400 2285.635 ;
        RECT 2408.200 2285.150 2408.460 2285.470 ;
        RECT 2381.520 2284.470 2381.780 2284.790 ;
        RECT 2415.160 2284.450 2415.300 2286.995 ;
        RECT 2415.620 2286.490 2415.760 2297.310 ;
        RECT 2422.000 2290.765 2422.260 2290.910 ;
        RECT 2416.010 2290.395 2416.290 2290.765 ;
        RECT 2421.990 2290.395 2422.270 2290.765 ;
        RECT 2416.080 2290.230 2416.220 2290.395 ;
        RECT 2416.020 2289.910 2416.280 2290.230 ;
        RECT 2435.790 2289.715 2436.070 2290.085 ;
        RECT 2435.860 2289.550 2436.000 2289.715 ;
        RECT 2421.990 2289.035 2422.270 2289.405 ;
        RECT 2435.800 2289.230 2436.060 2289.550 ;
        RECT 2422.000 2288.890 2422.260 2289.035 ;
        RECT 2428.890 2288.355 2429.170 2288.725 ;
        RECT 2442.690 2288.355 2442.970 2288.725 ;
        RECT 2428.960 2287.850 2429.100 2288.355 ;
        RECT 2442.700 2288.210 2442.960 2288.355 ;
        RECT 2428.900 2287.530 2429.160 2287.850 ;
        RECT 2435.790 2287.675 2436.070 2288.045 ;
        RECT 2435.860 2287.510 2436.000 2287.675 ;
        RECT 2428.890 2286.995 2429.170 2287.365 ;
        RECT 2435.800 2287.190 2436.060 2287.510 ;
        RECT 2442.690 2286.995 2442.970 2287.365 ;
        RECT 2428.960 2286.830 2429.100 2286.995 ;
        RECT 2442.700 2286.850 2442.960 2286.995 ;
        RECT 2428.900 2286.510 2429.160 2286.830 ;
        RECT 2415.560 2286.170 2415.820 2286.490 ;
        RECT 2415.100 2284.130 2415.360 2284.450 ;
        RECT 2381.060 2062.790 2381.320 2063.110 ;
        RECT 2373.700 2055.990 2373.960 2056.310 ;
        RECT 2366.800 2042.050 2367.060 2042.370 ;
        RECT 2359.900 2035.250 2360.160 2035.570 ;
        RECT 2353.000 2021.310 2353.260 2021.630 ;
        RECT 2346.100 2007.710 2346.360 2008.030 ;
        RECT 2339.660 2000.570 2339.920 2000.890 ;
        RECT 2339.200 1986.970 2339.460 1987.290 ;
        RECT 2332.300 1979.830 2332.560 1980.150 ;
        RECT 2325.400 1966.230 2325.660 1966.550 ;
        RECT 2318.500 1952.290 2318.760 1952.610 ;
        RECT 2311.600 1945.490 2311.860 1945.810 ;
        RECT 2305.160 1931.550 2305.420 1931.870 ;
        RECT 2304.700 1924.750 2304.960 1925.070 ;
        RECT 2301.940 1745.230 2302.200 1745.550 ;
        RECT 2301.020 1738.430 2301.280 1738.750 ;
        RECT 2294.120 1724.830 2294.380 1725.150 ;
        RECT 2287.220 1710.890 2287.480 1711.210 ;
        RECT 2280.320 1704.090 2280.580 1704.410 ;
        RECT 2273.420 1690.150 2273.680 1690.470 ;
        RECT 2267.440 1683.350 2267.700 1683.670 ;
        RECT 2266.520 1669.410 2266.780 1669.730 ;
        RECT 2252.720 1414.070 2252.980 1414.390 ;
        RECT 2245.820 1407.270 2246.080 1407.590 ;
        RECT 2238.920 1393.330 2239.180 1393.650 ;
        RECT 2232.020 1386.530 2232.280 1386.850 ;
        RECT 1794.100 1372.930 1794.360 1373.250 ;
        RECT 1787.200 1358.990 1787.460 1359.310 ;
        RECT 1780.300 1352.190 1780.560 1352.510 ;
        RECT 1773.400 1338.250 1773.660 1338.570 ;
        RECT 1766.500 1331.450 1766.760 1331.770 ;
        RECT 1760.060 1317.510 1760.320 1317.830 ;
        RECT 1759.600 1303.910 1759.860 1304.230 ;
        RECT 1752.700 1296.770 1752.960 1297.090 ;
        RECT 1745.800 1283.170 1746.060 1283.490 ;
        RECT 1738.900 1276.030 1739.160 1276.350 ;
        RECT 1732.000 1262.430 1732.260 1262.750 ;
        RECT 1725.100 1248.490 1725.360 1248.810 ;
        RECT 1718.660 1241.690 1718.920 1242.010 ;
        RECT 1718.200 1227.750 1718.460 1228.070 ;
        RECT 1711.300 1220.950 1711.560 1221.270 ;
        RECT 1704.400 1207.010 1704.660 1207.330 ;
        RECT 1697.500 1193.410 1697.760 1193.730 ;
        RECT 1690.600 1186.610 1690.860 1186.930 ;
        RECT 1684.160 1172.670 1684.420 1172.990 ;
        RECT 1683.700 1165.870 1683.960 1166.190 ;
        RECT 1676.800 1151.930 1677.060 1152.250 ;
        RECT 1669.900 1138.330 1670.160 1138.650 ;
        RECT 1663.000 1131.190 1663.260 1131.510 ;
        RECT 1649.660 1110.450 1649.920 1110.770 ;
        RECT 1635.400 1076.110 1635.660 1076.430 ;
        RECT 1628.500 1062.170 1628.760 1062.490 ;
        RECT 1614.700 1041.430 1614.960 1041.750 ;
        RECT 1607.800 1027.830 1608.060 1028.150 ;
        RECT 1514.410 1005.875 1514.690 1006.245 ;
      LAYER met2 ;
        RECT 305.710 1004.000 315.450 1004.280 ;
        RECT 316.290 1004.000 326.030 1004.280 ;
        RECT 326.870 1004.000 336.610 1004.280 ;
        RECT 337.450 1004.000 347.190 1004.280 ;
        RECT 348.030 1004.000 357.770 1004.280 ;
        RECT 358.610 1004.000 368.350 1004.280 ;
        RECT 369.190 1004.000 378.930 1004.280 ;
        RECT 379.770 1004.000 389.510 1004.280 ;
        RECT 390.350 1004.000 400.090 1004.280 ;
        RECT 400.930 1004.000 410.670 1004.280 ;
        RECT 411.510 1004.000 421.250 1004.280 ;
        RECT 422.090 1004.000 432.290 1004.280 ;
        RECT 433.130 1004.000 442.870 1004.280 ;
        RECT 443.710 1004.000 453.450 1004.280 ;
        RECT 454.290 1004.000 464.030 1004.280 ;
        RECT 464.870 1004.000 474.610 1004.280 ;
        RECT 475.450 1004.000 485.190 1004.280 ;
        RECT 486.030 1004.000 495.770 1004.280 ;
        RECT 496.610 1004.000 506.350 1004.280 ;
        RECT 507.190 1004.000 516.930 1004.280 ;
        RECT 517.770 1004.000 527.510 1004.280 ;
        RECT 528.350 1004.000 538.090 1004.280 ;
        RECT 538.930 1004.000 549.130 1004.280 ;
        RECT 549.970 1004.000 559.710 1004.280 ;
        RECT 560.550 1004.000 570.290 1004.280 ;
        RECT 571.130 1004.000 580.870 1004.280 ;
        RECT 581.710 1004.000 591.450 1004.280 ;
        RECT 592.290 1004.000 602.030 1004.280 ;
        RECT 602.870 1004.000 612.610 1004.280 ;
        RECT 613.450 1004.000 623.190 1004.280 ;
        RECT 624.030 1004.000 633.770 1004.280 ;
        RECT 634.610 1004.000 644.350 1004.280 ;
        RECT 645.190 1004.000 654.930 1004.280 ;
        RECT 655.770 1004.000 665.970 1004.280 ;
        RECT 666.810 1004.000 676.550 1004.280 ;
        RECT 677.390 1004.000 687.130 1004.280 ;
        RECT 687.970 1004.000 697.710 1004.280 ;
        RECT 698.550 1004.000 708.290 1004.280 ;
        RECT 709.130 1004.000 718.870 1004.280 ;
        RECT 719.710 1004.000 729.450 1004.280 ;
        RECT 730.290 1004.000 740.030 1004.280 ;
        RECT 740.870 1004.000 750.610 1004.280 ;
        RECT 751.450 1004.000 761.190 1004.280 ;
        RECT 762.030 1004.000 771.770 1004.280 ;
        RECT 772.610 1004.000 782.350 1004.280 ;
        RECT 783.190 1004.000 793.390 1004.280 ;
        RECT 794.230 1004.000 803.970 1004.280 ;
        RECT 804.810 1004.000 814.550 1004.280 ;
        RECT 815.390 1004.000 825.130 1004.280 ;
        RECT 825.970 1004.000 835.710 1004.280 ;
        RECT 836.550 1004.000 846.290 1004.280 ;
        RECT 847.130 1004.000 856.870 1004.280 ;
        RECT 857.710 1004.000 867.450 1004.280 ;
        RECT 868.290 1004.000 878.030 1004.280 ;
        RECT 878.870 1004.000 888.610 1004.280 ;
        RECT 889.450 1004.000 899.190 1004.280 ;
        RECT 900.030 1004.000 910.230 1004.280 ;
        RECT 911.070 1004.000 920.810 1004.280 ;
        RECT 921.650 1004.000 931.390 1004.280 ;
        RECT 932.230 1004.000 941.970 1004.280 ;
        RECT 942.810 1004.000 952.550 1004.280 ;
        RECT 953.390 1004.000 963.130 1004.280 ;
        RECT 963.970 1004.000 973.710 1004.280 ;
        RECT 974.550 1004.000 984.290 1004.280 ;
        RECT 985.130 1004.000 994.870 1004.280 ;
        RECT 995.710 1004.000 1005.450 1004.280 ;
        RECT 1006.290 1004.000 1016.030 1004.280 ;
        RECT 1016.870 1004.000 1027.070 1004.280 ;
        RECT 1027.910 1004.000 1037.650 1004.280 ;
        RECT 1038.490 1004.000 1048.230 1004.280 ;
        RECT 1049.070 1004.000 1058.810 1004.280 ;
        RECT 1059.650 1004.000 1069.390 1004.280 ;
        RECT 1070.230 1004.000 1079.970 1004.280 ;
        RECT 1080.810 1004.000 1090.550 1004.280 ;
        RECT 1091.390 1004.000 1101.130 1004.280 ;
        RECT 1101.970 1004.000 1111.710 1004.280 ;
        RECT 1112.550 1004.000 1122.290 1004.280 ;
        RECT 1123.130 1004.000 1132.870 1004.280 ;
        RECT 1133.710 1004.000 1143.450 1004.280 ;
        RECT 1144.290 1004.000 1154.490 1004.280 ;
        RECT 1155.330 1004.000 1165.070 1004.280 ;
        RECT 1165.910 1004.000 1175.650 1004.280 ;
        RECT 1176.490 1004.000 1186.230 1004.280 ;
        RECT 1187.070 1004.000 1196.810 1004.280 ;
        RECT 1197.650 1004.000 1207.390 1004.280 ;
        RECT 1208.230 1004.000 1217.970 1004.280 ;
        RECT 1218.810 1004.000 1228.550 1004.280 ;
        RECT 1229.390 1004.000 1239.130 1004.280 ;
        RECT 1239.970 1004.000 1249.710 1004.280 ;
        RECT 1250.550 1004.000 1260.290 1004.280 ;
        RECT 1261.130 1004.000 1271.330 1004.280 ;
        RECT 1272.170 1004.000 1281.910 1004.280 ;
        RECT 1282.750 1004.000 1292.490 1004.280 ;
        RECT 1293.330 1004.000 1303.070 1004.280 ;
        RECT 1303.910 1004.000 1313.650 1004.280 ;
        RECT 1314.490 1004.000 1324.230 1004.280 ;
        RECT 1325.070 1004.000 1334.810 1004.280 ;
        RECT 1335.650 1004.000 1345.390 1004.280 ;
        RECT 1346.230 1004.000 1355.970 1004.280 ;
        RECT 1356.810 1004.000 1366.550 1004.280 ;
        RECT 1367.390 1004.000 1377.130 1004.280 ;
        RECT 1377.970 1004.000 1388.170 1004.280 ;
        RECT 1389.010 1004.000 1398.750 1004.280 ;
        RECT 1399.590 1004.000 1409.330 1004.280 ;
        RECT 1410.170 1004.000 1419.910 1004.280 ;
        RECT 1420.750 1004.000 1430.490 1004.280 ;
        RECT 1431.330 1004.000 1441.070 1004.280 ;
        RECT 1441.910 1004.000 1451.650 1004.280 ;
        RECT 1452.490 1004.000 1462.230 1004.280 ;
        RECT 1463.070 1004.000 1472.810 1004.280 ;
        RECT 1473.650 1004.000 1483.390 1004.280 ;
        RECT 1484.230 1004.000 1493.970 1004.280 ;
      LAYER via2 ;
        RECT 668.470 2767.120 668.750 2767.400 ;
        RECT 1295.910 2767.120 1296.190 2767.400 ;
        RECT 1318.910 2767.120 1319.190 2767.400 ;
        RECT 1892.530 2767.120 1892.810 2767.400 ;
        RECT 1914.610 2767.120 1914.890 2767.400 ;
        RECT 2539.290 2767.120 2539.570 2767.400 ;
        RECT 2566.890 2767.120 2567.170 2767.400 ;
        RECT 287.590 2732.440 287.870 2732.720 ;
        RECT 287.130 2725.640 287.410 2725.920 ;
        RECT 284.370 2718.840 284.650 2719.120 ;
        RECT 283.910 2701.840 284.190 2702.120 ;
        RECT 286.670 2712.040 286.950 2712.320 ;
        RECT 285.750 2697.760 286.030 2698.040 ;
        RECT 285.290 2687.560 285.570 2687.840 ;
        RECT 284.830 2401.280 285.110 2401.560 ;
        RECT 284.370 2212.240 284.650 2212.520 ;
        RECT 287.130 2211.560 287.410 2211.840 ;
        RECT 299.090 2392.635 299.370 2392.915 ;
        RECT 696.990 2749.440 697.270 2749.720 ;
        RECT 386.490 2297.240 386.770 2297.520 ;
        RECT 370.850 2290.440 371.130 2290.720 ;
        RECT 379.130 2290.440 379.410 2290.720 ;
        RECT 399.830 2290.440 400.110 2290.720 ;
        RECT 409.490 2290.440 409.770 2290.720 ;
        RECT 414.090 2290.440 414.370 2290.720 ;
        RECT 420.990 2290.440 421.270 2290.720 ;
        RECT 427.430 2290.440 427.710 2290.720 ;
        RECT 431.570 2290.440 431.850 2290.720 ;
        RECT 365.330 2288.400 365.610 2288.680 ;
        RECT 406.730 2289.760 407.010 2290.040 ;
        RECT 392.930 2289.080 393.210 2289.360 ;
        RECT 386.030 2287.720 386.310 2288.000 ;
        RECT 439.390 2290.440 439.670 2290.720 ;
        RECT 445.370 2290.440 445.650 2290.720 ;
        RECT 450.890 2290.440 451.170 2290.720 ;
        RECT 455.490 2290.440 455.770 2290.720 ;
        RECT 462.390 2290.440 462.670 2290.720 ;
        RECT 467.910 2290.440 468.190 2290.720 ;
        RECT 473.890 2290.440 474.170 2290.720 ;
        RECT 478.950 2290.440 479.230 2290.720 ;
        RECT 485.850 2290.440 486.130 2290.720 ;
        RECT 492.750 2290.440 493.030 2290.720 ;
        RECT 497.350 2290.440 497.630 2290.720 ;
        RECT 503.330 2290.440 503.610 2290.720 ;
        RECT 509.770 2290.440 510.050 2290.720 ;
        RECT 513.910 2290.440 514.190 2290.720 ;
        RECT 517.130 2290.440 517.410 2290.720 ;
        RECT 521.270 2290.440 521.550 2290.720 ;
        RECT 524.030 2290.440 524.310 2290.720 ;
        RECT 526.790 2290.440 527.070 2290.720 ;
        RECT 530.930 2290.440 531.210 2290.720 ;
        RECT 537.830 2290.440 538.110 2290.720 ;
        RECT 502.870 2289.760 503.150 2290.040 ;
        RECT 365.790 2287.040 366.070 2287.320 ;
        RECT 379.590 2287.040 379.870 2287.320 ;
        RECT 358.890 2285.680 359.170 2285.960 ;
        RECT 287.590 2210.880 287.870 2211.160 ;
        RECT 351.070 2285.000 351.350 2285.280 ;
        RECT 337.730 2284.320 338.010 2284.600 ;
        RECT 344.170 2284.320 344.450 2284.600 ;
        RECT 350.610 2284.320 350.890 2284.600 ;
        RECT 358.430 2284.320 358.710 2284.600 ;
        RECT 373.610 2285.000 373.890 2285.280 ;
        RECT 386.490 2285.680 386.770 2285.960 ;
        RECT 475.730 2285.680 476.010 2285.960 ;
        RECT 496.430 2285.680 496.710 2285.960 ;
        RECT 393.850 2285.000 394.130 2285.280 ;
        RECT 468.830 2285.000 469.110 2285.280 ;
        RECT 393.390 2284.320 393.670 2284.600 ;
        RECT 400.290 2284.320 400.570 2284.600 ;
        RECT 407.190 2284.320 407.470 2284.600 ;
        RECT 414.090 2284.320 414.370 2284.600 ;
        RECT 420.990 2284.320 421.270 2284.600 ;
        RECT 431.110 2284.320 431.390 2284.600 ;
        RECT 434.330 2284.320 434.610 2284.600 ;
        RECT 441.230 2284.320 441.510 2284.600 ;
        RECT 448.130 2284.320 448.410 2284.600 ;
        RECT 455.030 2284.320 455.310 2284.600 ;
        RECT 461.930 2284.320 462.210 2284.600 ;
        RECT 468.370 2284.320 468.650 2284.600 ;
        RECT 482.630 2284.320 482.910 2284.600 ;
        RECT 489.530 2284.320 489.810 2284.600 ;
        RECT 509.310 2289.080 509.590 2289.360 ;
        RECT 510.230 2289.760 510.510 2290.040 ;
        RECT 531.390 2289.760 531.670 2290.040 ;
        RECT 543.810 2290.440 544.090 2290.720 ;
        RECT 551.630 2290.440 551.910 2290.720 ;
        RECT 538.290 2289.760 538.570 2290.040 ;
        RECT 544.730 2289.760 545.010 2290.040 ;
        RECT 938.490 2732.440 938.770 2732.720 ;
        RECT 696.990 2447.520 697.270 2447.800 ;
        RECT 938.490 2725.640 938.770 2725.920 ;
        RECT 938.490 2718.840 938.770 2719.120 ;
        RECT 938.490 2712.720 938.770 2713.000 ;
        RECT 938.950 2701.840 939.230 2702.120 ;
        RECT 938.490 2699.120 938.770 2699.400 ;
        RECT 941.710 2687.560 941.990 2687.840 ;
        RECT 814.750 2212.240 815.030 2212.520 ;
        RECT 826.250 2211.560 826.530 2211.840 ;
        RECT 837.290 2210.880 837.570 2211.160 ;
        RECT 944.930 2401.280 945.210 2401.560 ;
        RECT 944.470 2389.720 944.750 2390.000 ;
        RECT 1332.250 2749.440 1332.530 2749.720 ;
        RECT 1352.030 2746.720 1352.310 2747.000 ;
        RECT 1345.590 2422.360 1345.870 2422.640 ;
        RECT 986.790 2289.760 987.070 2290.040 ;
        RECT 993.690 2289.760 993.970 2290.040 ;
        RECT 1001.050 2290.440 1001.330 2290.720 ;
        RECT 979.890 2287.720 980.170 2288.000 ;
        RECT 1038.310 2289.760 1038.590 2290.040 ;
        RECT 1041.070 2289.760 1041.350 2290.040 ;
        RECT 1007.490 2288.400 1007.770 2288.680 ;
        RECT 1031.410 2286.360 1031.690 2286.640 ;
        RECT 1034.170 2286.360 1034.450 2286.640 ;
        RECT 1010.710 2285.680 1010.990 2285.960 ;
        RECT 1013.930 2285.680 1014.210 2285.960 ;
        RECT 1024.510 2285.000 1024.790 2285.280 ;
        RECT 1027.270 2285.000 1027.550 2285.280 ;
        RECT 1017.610 2284.320 1017.890 2284.600 ;
        RECT 1020.830 2284.320 1021.110 2284.600 ;
        RECT 1027.730 2284.320 1028.010 2284.600 ;
        RECT 1034.630 2285.680 1034.910 2285.960 ;
        RECT 1048.430 2288.400 1048.710 2288.680 ;
        RECT 1045.210 2287.040 1045.490 2287.320 ;
        RECT 1041.530 2284.320 1041.810 2284.600 ;
        RECT 1052.570 2290.440 1052.850 2290.720 ;
        RECT 1062.230 2290.440 1062.510 2290.720 ;
        RECT 1065.450 2290.440 1065.730 2290.720 ;
        RECT 1070.050 2290.440 1070.330 2290.720 ;
        RECT 1076.490 2290.440 1076.770 2290.720 ;
        RECT 1083.390 2290.440 1083.670 2290.720 ;
        RECT 1048.430 2284.320 1048.710 2284.600 ;
        RECT 1054.870 2285.680 1055.150 2285.960 ;
        RECT 1055.330 2284.320 1055.610 2284.600 ;
        RECT 1062.230 2284.320 1062.510 2284.600 ;
        RECT 1069.130 2284.320 1069.410 2284.600 ;
        RECT 1076.030 2285.680 1076.310 2285.960 ;
        RECT 1087.990 2290.440 1088.270 2290.720 ;
        RECT 1094.430 2290.440 1094.710 2290.720 ;
        RECT 1082.930 2287.040 1083.210 2287.320 ;
        RECT 1100.870 2290.440 1101.150 2290.720 ;
        RECT 1106.850 2290.440 1107.130 2290.720 ;
        RECT 1112.830 2290.440 1113.110 2290.720 ;
        RECT 1089.830 2285.680 1090.110 2285.960 ;
        RECT 1103.630 2285.680 1103.910 2285.960 ;
        RECT 1089.370 2284.320 1089.650 2284.600 ;
        RECT 1096.730 2284.320 1097.010 2284.600 ;
        RECT 1118.350 2290.440 1118.630 2290.720 ;
        RECT 1121.570 2290.440 1121.850 2290.720 ;
        RECT 1129.390 2290.440 1129.670 2290.720 ;
        RECT 1110.530 2284.320 1110.810 2284.600 ;
        RECT 1117.430 2284.320 1117.710 2284.600 ;
        RECT 1131.230 2285.000 1131.510 2285.280 ;
        RECT 1124.330 2284.320 1124.610 2284.600 ;
        RECT 1130.770 2284.320 1131.050 2284.600 ;
        RECT 1135.830 2290.440 1136.110 2290.720 ;
        RECT 1141.810 2290.440 1142.090 2290.720 ;
        RECT 1147.790 2290.440 1148.070 2290.720 ;
        RECT 1159.290 2290.440 1159.570 2290.720 ;
        RECT 1166.190 2290.440 1166.470 2290.720 ;
        RECT 1173.090 2289.760 1173.370 2290.040 ;
        RECT 1159.290 2289.080 1159.570 2289.360 ;
        RECT 1179.990 2289.080 1180.270 2289.360 ;
        RECT 1186.890 2288.400 1187.170 2288.680 ;
        RECT 1193.790 2288.400 1194.070 2288.680 ;
        RECT 1152.390 2287.720 1152.670 2288.000 ;
        RECT 1165.270 2285.000 1165.550 2285.280 ;
        RECT 1138.130 2284.320 1138.410 2284.600 ;
        RECT 1145.030 2284.320 1145.310 2284.600 ;
        RECT 1151.930 2284.320 1152.210 2284.600 ;
        RECT 1158.830 2284.320 1159.110 2284.600 ;
        RECT 1165.730 2284.320 1166.010 2284.600 ;
        RECT 1172.630 2284.320 1172.910 2284.600 ;
        RECT 1179.530 2284.320 1179.810 2284.600 ;
        RECT 1186.430 2284.320 1186.710 2284.600 ;
        RECT 1193.330 2284.320 1193.610 2284.600 ;
        RECT 1200.230 2284.320 1200.510 2284.600 ;
        RECT 1165.730 2212.240 1166.010 2212.520 ;
        RECT 1172.630 2211.560 1172.910 2211.840 ;
        RECT 1186.430 2210.880 1186.710 2211.160 ;
        RECT 1200.230 2208.160 1200.510 2208.440 ;
        RECT 1243.470 2208.160 1243.750 2208.440 ;
        RECT 1437.590 2212.240 1437.870 2212.520 ;
        RECT 1448.630 2211.560 1448.910 2211.840 ;
        RECT 1471.630 2210.880 1471.910 2211.160 ;
        RECT 1529.130 2732.440 1529.410 2732.720 ;
        RECT 1513.950 2183.680 1514.230 2183.960 ;
        RECT 1513.950 2172.800 1514.230 2173.080 ;
        RECT 1513.950 2161.920 1514.230 2162.200 ;
        RECT 1513.950 2151.040 1514.230 2151.320 ;
        RECT 1513.950 2139.480 1514.230 2139.760 ;
        RECT 1513.950 2128.600 1514.230 2128.880 ;
        RECT 1513.950 2117.720 1514.230 2118.000 ;
        RECT 1513.950 2106.840 1514.230 2107.120 ;
        RECT 1513.950 2095.960 1514.230 2096.240 ;
        RECT 1513.950 2084.400 1514.230 2084.680 ;
        RECT 1513.950 2073.520 1514.230 2073.800 ;
        RECT 1513.950 2062.640 1514.230 2062.920 ;
        RECT 1513.950 2051.760 1514.230 2052.040 ;
        RECT 1513.950 2040.880 1514.230 2041.160 ;
        RECT 1513.950 2029.320 1514.230 2029.600 ;
        RECT 1513.490 2018.440 1513.770 2018.720 ;
        RECT 1513.950 2007.560 1514.230 2007.840 ;
        RECT 1513.950 1996.680 1514.230 1996.960 ;
        RECT 1513.950 1985.800 1514.230 1986.080 ;
        RECT 1512.570 1974.240 1512.850 1974.520 ;
        RECT 1513.490 1963.360 1513.770 1963.640 ;
        RECT 1513.950 1952.480 1514.230 1952.760 ;
        RECT 1513.950 1941.600 1514.230 1941.880 ;
        RECT 1512.570 1930.720 1512.850 1931.000 ;
        RECT 1512.570 1919.160 1512.850 1919.440 ;
        RECT 1513.950 1908.280 1514.230 1908.560 ;
        RECT 1513.030 1897.400 1513.310 1897.680 ;
        RECT 1513.950 1886.520 1514.230 1886.800 ;
        RECT 1513.950 1875.640 1514.230 1875.920 ;
        RECT 1513.950 1864.760 1514.230 1865.040 ;
        RECT 1511.650 1853.200 1511.930 1853.480 ;
        RECT 1513.030 1842.320 1513.310 1842.600 ;
        RECT 1513.950 1831.440 1514.230 1831.720 ;
        RECT 1512.570 1820.560 1512.850 1820.840 ;
        RECT 1512.110 1809.680 1512.390 1809.960 ;
        RECT 1511.650 1798.120 1511.930 1798.400 ;
        RECT 1512.570 1787.240 1512.850 1787.520 ;
        RECT 1513.950 1776.360 1514.230 1776.640 ;
        RECT 1513.950 1765.480 1514.230 1765.760 ;
        RECT 1512.110 1754.600 1512.390 1754.880 ;
        RECT 1513.490 1743.040 1513.770 1743.320 ;
        RECT 1512.570 1732.160 1512.850 1732.440 ;
        RECT 1513.950 1721.280 1514.230 1721.560 ;
        RECT 1513.950 1710.400 1514.230 1710.680 ;
        RECT 1512.110 1699.520 1512.390 1699.800 ;
        RECT 1513.490 1687.960 1513.770 1688.240 ;
        RECT 1512.570 1677.080 1512.850 1677.360 ;
        RECT 1513.950 1666.200 1514.230 1666.480 ;
        RECT 1512.570 1655.320 1512.850 1655.600 ;
        RECT 1511.650 1644.440 1511.930 1644.720 ;
        RECT 1512.570 1632.880 1512.850 1633.160 ;
        RECT 1511.650 1622.000 1511.930 1622.280 ;
        RECT 1511.650 1611.120 1511.930 1611.400 ;
        RECT 1511.650 1600.240 1511.930 1600.520 ;
        RECT 1513.490 1589.360 1513.770 1589.640 ;
        RECT 1513.950 1578.480 1514.230 1578.760 ;
        RECT 1513.950 1566.920 1514.230 1567.200 ;
        RECT 1513.490 1556.040 1513.770 1556.320 ;
        RECT 1513.950 1545.160 1514.230 1545.440 ;
        RECT 1513.950 1534.280 1514.230 1534.560 ;
        RECT 1513.950 1523.400 1514.230 1523.680 ;
        RECT 1513.950 1511.840 1514.230 1512.120 ;
        RECT 1513.490 1500.960 1513.770 1501.240 ;
        RECT 1513.950 1490.080 1514.230 1490.360 ;
        RECT 1513.030 1479.200 1513.310 1479.480 ;
        RECT 1513.950 1468.320 1514.230 1468.600 ;
        RECT 1512.570 1456.760 1512.850 1457.040 ;
        RECT 1513.490 1445.880 1513.770 1446.160 ;
        RECT 1513.950 1435.000 1514.230 1435.280 ;
        RECT 1513.490 1424.120 1513.770 1424.400 ;
        RECT 1512.570 1413.240 1512.850 1413.520 ;
        RECT 1512.570 1401.680 1512.850 1401.960 ;
        RECT 1511.650 1390.800 1511.930 1391.080 ;
        RECT 1513.030 1379.920 1513.310 1380.200 ;
        RECT 1513.950 1369.040 1514.230 1369.320 ;
        RECT 1512.570 1358.160 1512.850 1358.440 ;
        RECT 1512.570 1346.600 1512.850 1346.880 ;
        RECT 1511.650 1335.720 1511.930 1336.000 ;
        RECT 1513.030 1324.840 1513.310 1325.120 ;
        RECT 1513.950 1313.960 1514.230 1314.240 ;
        RECT 1512.570 1303.080 1512.850 1303.360 ;
        RECT 1512.110 1292.200 1512.390 1292.480 ;
        RECT 1511.650 1280.640 1511.930 1280.920 ;
        RECT 1512.570 1269.760 1512.850 1270.040 ;
        RECT 1513.950 1258.880 1514.230 1259.160 ;
        RECT 1513.950 1248.000 1514.230 1248.280 ;
        RECT 1512.110 1237.120 1512.390 1237.400 ;
        RECT 1513.490 1225.560 1513.770 1225.840 ;
        RECT 1512.570 1214.680 1512.850 1214.960 ;
        RECT 1513.950 1203.800 1514.230 1204.080 ;
        RECT 1513.950 1192.920 1514.230 1193.200 ;
        RECT 1512.110 1182.040 1512.390 1182.320 ;
        RECT 1513.490 1170.480 1513.770 1170.760 ;
        RECT 1512.570 1159.600 1512.850 1159.880 ;
        RECT 1513.950 1148.720 1514.230 1149.000 ;
        RECT 1513.950 1137.840 1514.230 1138.120 ;
        RECT 1513.950 1126.960 1514.230 1127.240 ;
        RECT 1513.490 1115.400 1513.770 1115.680 ;
        RECT 1513.950 1104.520 1514.230 1104.800 ;
        RECT 1513.950 1093.640 1514.230 1093.920 ;
        RECT 1513.950 1082.760 1514.230 1083.040 ;
        RECT 1513.950 1071.880 1514.230 1072.160 ;
        RECT 1513.030 1060.320 1513.310 1060.600 ;
        RECT 1513.950 1049.440 1514.230 1049.720 ;
        RECT 1513.950 1038.560 1514.230 1038.840 ;
        RECT 1513.950 1027.680 1514.230 1027.960 ;
        RECT 1511.190 1016.800 1511.470 1017.080 ;
        RECT 1514.870 2194.560 1515.150 2194.840 ;
        RECT 1528.670 2718.840 1528.950 2719.120 ;
        RECT 1528.210 2697.760 1528.490 2698.040 ;
        RECT 1538.330 2725.640 1538.610 2725.920 ;
        RECT 1536.030 2712.040 1536.310 2712.320 ;
        RECT 1536.490 2701.840 1536.770 2702.120 ;
        RECT 1538.330 2699.120 1538.610 2699.400 ;
        RECT 1536.490 2697.760 1536.770 2698.040 ;
        RECT 1535.110 2687.560 1535.390 2687.840 ;
        RECT 1529.590 2401.280 1529.870 2401.560 ;
        RECT 1535.570 2390.400 1535.850 2390.680 ;
        RECT 1945.890 2749.440 1946.170 2749.720 ;
        RECT 2594.490 2753.520 2594.770 2753.800 ;
        RECT 1759.130 2297.920 1759.410 2298.200 ;
        RECT 1639.530 2297.240 1639.810 2297.520 ;
        RECT 1607.790 2290.440 1608.070 2290.720 ;
        RECT 1614.690 2290.440 1614.970 2290.720 ;
        RECT 1628.490 2290.440 1628.770 2290.720 ;
        RECT 1635.390 2290.440 1635.670 2290.720 ;
        RECT 1587.090 2289.080 1587.370 2289.360 ;
        RECT 1601.350 2285.000 1601.630 2285.280 ;
        RECT 1580.190 2284.320 1580.470 2284.600 ;
        RECT 1593.990 2284.320 1594.270 2284.600 ;
        RECT 1600.890 2284.320 1601.170 2284.600 ;
        RECT 1611.010 2289.760 1611.290 2290.040 ;
        RECT 1617.910 2289.760 1618.190 2290.040 ;
        RECT 1624.810 2289.080 1625.090 2289.360 ;
        RECT 1621.590 2285.680 1621.870 2285.960 ;
        RECT 1631.710 2289.080 1631.990 2289.360 ;
        RECT 1645.510 2290.440 1645.790 2290.720 ;
        RECT 1649.650 2290.440 1649.930 2290.720 ;
        RECT 1659.310 2290.440 1659.590 2290.720 ;
        RECT 1665.750 2290.440 1666.030 2290.720 ;
        RECT 1670.350 2290.440 1670.630 2290.720 ;
        RECT 1676.790 2290.440 1677.070 2290.720 ;
        RECT 1642.290 2285.680 1642.570 2285.960 ;
        RECT 1638.610 2270.040 1638.890 2270.320 ;
        RECT 1639.530 2270.040 1639.810 2270.320 ;
        RECT 1639.070 1834.840 1639.350 1835.120 ;
        RECT 1640.450 1834.840 1640.730 1835.120 ;
        RECT 1646.430 2289.760 1646.710 2290.040 ;
        RECT 1649.190 2286.360 1649.470 2286.640 ;
        RECT 1652.410 2289.080 1652.690 2289.360 ;
        RECT 1656.090 2288.400 1656.370 2288.680 ;
        RECT 1676.790 2285.680 1677.070 2285.960 ;
        RECT 1662.990 2284.320 1663.270 2284.600 ;
        RECT 1669.890 2284.320 1670.170 2284.600 ;
        RECT 1682.770 2290.440 1683.050 2290.720 ;
        RECT 1690.130 2290.440 1690.410 2290.720 ;
        RECT 1695.190 2290.440 1695.470 2290.720 ;
        RECT 1699.330 2290.440 1699.610 2290.720 ;
        RECT 1706.230 2290.440 1706.510 2290.720 ;
        RECT 1711.290 2290.440 1711.570 2290.720 ;
        RECT 1718.190 2290.440 1718.470 2290.720 ;
        RECT 1684.150 2285.000 1684.430 2285.280 ;
        RECT 1683.690 2284.320 1683.970 2284.600 ;
        RECT 1690.590 2284.320 1690.870 2284.600 ;
        RECT 1697.490 2284.320 1697.770 2284.600 ;
        RECT 1704.390 2285.680 1704.670 2285.960 ;
        RECT 1712.670 2289.760 1712.950 2290.040 ;
        RECT 1723.710 2290.440 1723.990 2290.720 ;
        RECT 1725.090 2290.440 1725.370 2290.720 ;
        RECT 1731.990 2290.440 1732.270 2290.720 ;
        RECT 1738.890 2290.440 1739.170 2290.720 ;
        RECT 1745.790 2290.440 1746.070 2290.720 ;
        RECT 1721.870 2289.760 1722.150 2290.040 ;
        RECT 1718.650 2288.400 1718.930 2288.680 ;
        RECT 1729.690 2289.760 1729.970 2290.040 ;
        RECT 1734.290 2289.760 1734.570 2290.040 ;
        RECT 1741.190 2289.760 1741.470 2290.040 ;
        RECT 1794.090 2297.240 1794.370 2297.520 ;
        RECT 1759.590 2290.440 1759.870 2290.720 ;
        RECT 1766.490 2290.440 1766.770 2290.720 ;
        RECT 1746.250 2289.760 1746.530 2290.040 ;
        RECT 1752.690 2289.760 1752.970 2290.040 ;
        RECT 1752.690 2284.320 1752.970 2284.600 ;
        RECT 1760.050 2285.000 1760.330 2285.280 ;
        RECT 1759.590 2284.320 1759.870 2284.600 ;
        RECT 1766.490 2285.680 1766.770 2285.960 ;
        RECT 1780.290 2289.760 1780.570 2290.040 ;
        RECT 1775.230 2289.080 1775.510 2289.360 ;
        RECT 1787.190 2288.400 1787.470 2288.680 ;
        RECT 1773.390 2284.320 1773.670 2284.600 ;
        RECT 1780.290 2284.320 1780.570 2284.600 ;
        RECT 1787.190 2284.320 1787.470 2284.600 ;
        RECT 1794.090 2284.320 1794.370 2284.600 ;
        RECT 2187.390 2732.440 2187.670 2732.720 ;
        RECT 1945.890 2447.520 1946.170 2447.800 ;
        RECT 1945.890 2404.680 1946.170 2404.960 ;
        RECT 2187.390 2725.640 2187.670 2725.920 ;
        RECT 2187.390 2718.840 2187.670 2719.120 ;
        RECT 2187.390 2712.040 2187.670 2712.320 ;
        RECT 2187.850 2701.840 2188.130 2702.120 ;
        RECT 2187.390 2699.120 2187.670 2699.400 ;
        RECT 2187.390 2687.560 2187.670 2687.840 ;
        RECT 2187.390 2401.280 2187.670 2401.560 ;
        RECT 2190.610 2389.720 2190.890 2390.000 ;
        RECT 2582.070 2749.440 2582.350 2749.720 ;
        RECT 2594.490 2447.520 2594.770 2447.800 ;
        RECT 2415.090 2297.240 2415.370 2297.520 ;
        RECT 2308.830 2290.440 2309.110 2290.720 ;
        RECT 2315.270 2290.440 2315.550 2290.720 ;
        RECT 2324.930 2290.440 2325.210 2290.720 ;
        RECT 2325.850 2290.440 2326.130 2290.720 ;
        RECT 2343.790 2290.440 2344.070 2290.720 ;
        RECT 2349.770 2290.440 2350.050 2290.720 ;
        RECT 2358.970 2290.440 2359.250 2290.720 ;
        RECT 2361.270 2290.440 2361.550 2290.720 ;
        RECT 2367.250 2290.440 2367.530 2290.720 ;
        RECT 2374.150 2290.440 2374.430 2290.720 ;
        RECT 2377.370 2290.440 2377.650 2290.720 ;
        RECT 2384.730 2290.440 2385.010 2290.720 ;
        RECT 2391.630 2290.440 2391.910 2290.720 ;
        RECT 2397.150 2290.440 2397.430 2290.720 ;
        RECT 2415.090 2290.440 2415.370 2290.720 ;
        RECT 2301.010 2289.760 2301.290 2290.040 ;
        RECT 2290.890 2289.080 2291.170 2289.360 ;
        RECT 2263.290 2287.040 2263.570 2287.320 ;
        RECT 2252.710 2285.680 2252.990 2285.960 ;
        RECT 2232.010 2285.000 2232.290 2285.280 ;
        RECT 2228.790 2284.320 2229.070 2284.600 ;
        RECT 2238.910 2284.320 2239.190 2284.600 ;
        RECT 2245.810 2284.320 2246.090 2284.600 ;
        RECT 2283.990 2287.720 2284.270 2288.000 ;
        RECT 2297.790 2287.720 2298.070 2288.000 ;
        RECT 2270.190 2287.040 2270.470 2287.320 ;
        RECT 2273.410 2285.680 2273.690 2285.960 ;
        RECT 2294.110 2285.680 2294.390 2285.960 ;
        RECT 2296.870 2285.680 2297.150 2285.960 ;
        RECT 2263.750 2284.320 2264.030 2284.600 ;
        RECT 2266.510 2284.320 2266.790 2284.600 ;
        RECT 2267.430 2284.320 2267.710 2284.600 ;
        RECT 2280.310 2285.000 2280.590 2285.280 ;
        RECT 2283.530 2285.000 2283.810 2285.280 ;
        RECT 2277.090 2284.320 2277.370 2284.600 ;
        RECT 2287.210 2284.320 2287.490 2284.600 ;
        RECT 2290.430 2284.320 2290.710 2284.600 ;
        RECT 2301.930 2288.400 2302.210 2288.680 ;
        RECT 2340.110 2289.760 2340.390 2290.040 ;
        RECT 2333.210 2289.080 2333.490 2289.360 ;
        RECT 2305.150 2285.680 2305.430 2285.960 ;
        RECT 2304.690 2284.320 2304.970 2284.600 ;
        RECT 2311.590 2284.320 2311.870 2284.600 ;
        RECT 2318.490 2284.320 2318.770 2284.600 ;
        RECT 2325.390 2284.320 2325.670 2284.600 ;
        RECT 2332.290 2284.320 2332.570 2284.600 ;
        RECT 2339.650 2285.680 2339.930 2285.960 ;
        RECT 2339.190 2284.320 2339.470 2284.600 ;
        RECT 2346.090 2284.320 2346.370 2284.600 ;
        RECT 2352.990 2284.320 2353.270 2284.600 ;
        RECT 2359.890 2285.680 2360.170 2285.960 ;
        RECT 2366.790 2284.320 2367.070 2284.600 ;
        RECT 2373.690 2284.320 2373.970 2284.600 ;
        RECT 2394.390 2289.080 2394.670 2289.360 ;
        RECT 2380.590 2286.360 2380.870 2286.640 ;
        RECT 2381.050 2285.680 2381.330 2285.960 ;
        RECT 2387.490 2286.360 2387.770 2286.640 ;
        RECT 2402.210 2289.760 2402.490 2290.040 ;
        RECT 2402.670 2289.080 2402.950 2289.360 ;
        RECT 2408.190 2288.400 2408.470 2288.680 ;
        RECT 2415.090 2287.040 2415.370 2287.320 ;
        RECT 2408.190 2285.680 2408.470 2285.960 ;
        RECT 2416.010 2290.440 2416.290 2290.720 ;
        RECT 2421.990 2290.440 2422.270 2290.720 ;
        RECT 2435.790 2289.760 2436.070 2290.040 ;
        RECT 2421.990 2289.080 2422.270 2289.360 ;
        RECT 2428.890 2288.400 2429.170 2288.680 ;
        RECT 2442.690 2288.400 2442.970 2288.680 ;
        RECT 2435.790 2287.720 2436.070 2288.000 ;
        RECT 2428.890 2287.040 2429.170 2287.320 ;
        RECT 2442.690 2287.040 2442.970 2287.320 ;
        RECT 1514.410 1005.920 1514.690 1006.200 ;
      LAYER met3 ;
        RECT 668.445 2767.420 668.775 2767.425 ;
        RECT 1295.885 2767.420 1296.215 2767.425 ;
        RECT 1318.885 2767.420 1319.215 2767.425 ;
        RECT 668.190 2767.410 668.775 2767.420 ;
        RECT 1295.630 2767.410 1296.215 2767.420 ;
        RECT 1318.630 2767.410 1319.215 2767.420 ;
        RECT 667.990 2767.110 668.775 2767.410 ;
        RECT 1295.430 2767.110 1296.215 2767.410 ;
        RECT 1318.430 2767.110 1319.215 2767.410 ;
        RECT 668.190 2767.100 668.775 2767.110 ;
        RECT 1295.630 2767.100 1296.215 2767.110 ;
        RECT 1318.630 2767.100 1319.215 2767.110 ;
        RECT 668.445 2767.095 668.775 2767.100 ;
        RECT 1295.885 2767.095 1296.215 2767.100 ;
        RECT 1318.885 2767.095 1319.215 2767.100 ;
        RECT 1892.505 2767.420 1892.835 2767.425 ;
        RECT 1914.585 2767.420 1914.915 2767.425 ;
        RECT 2539.265 2767.420 2539.595 2767.425 ;
        RECT 2566.865 2767.420 2567.195 2767.425 ;
        RECT 1892.505 2767.410 1893.090 2767.420 ;
        RECT 1914.585 2767.410 1915.170 2767.420 ;
        RECT 2539.265 2767.410 2539.850 2767.420 ;
        RECT 2566.865 2767.410 2567.450 2767.420 ;
        RECT 1892.505 2767.110 1893.290 2767.410 ;
        RECT 1914.585 2767.110 1915.370 2767.410 ;
        RECT 2539.265 2767.110 2540.050 2767.410 ;
        RECT 2566.865 2767.110 2567.650 2767.410 ;
        RECT 1892.505 2767.100 1893.090 2767.110 ;
        RECT 1914.585 2767.100 1915.170 2767.110 ;
        RECT 2539.265 2767.100 2539.850 2767.110 ;
        RECT 2566.865 2767.100 2567.450 2767.110 ;
        RECT 1892.505 2767.095 1892.835 2767.100 ;
        RECT 1914.585 2767.095 1914.915 2767.100 ;
        RECT 2539.265 2767.095 2539.595 2767.100 ;
        RECT 2566.865 2767.095 2567.195 2767.100 ;
        RECT 646.110 2755.850 646.490 2755.860 ;
        RECT 664.510 2755.850 664.890 2755.860 ;
        RECT 646.110 2755.550 664.890 2755.850 ;
        RECT 646.110 2755.540 646.490 2755.550 ;
        RECT 664.510 2755.540 664.890 2755.550 ;
        RECT 2570.750 2753.810 2571.130 2753.820 ;
        RECT 2594.465 2753.810 2594.795 2753.825 ;
        RECT 2570.750 2753.510 2594.795 2753.810 ;
        RECT 2570.750 2753.500 2571.130 2753.510 ;
        RECT 2594.465 2753.495 2594.795 2753.510 ;
        RECT 659.280 2751.235 661.020 2752.140 ;
        RECT 1309.280 2751.235 1311.020 2752.140 ;
        RECT 1909.280 2751.235 1911.020 2752.140 ;
        RECT 2559.280 2751.235 2561.020 2752.140 ;
        RECT 297.470 2732.785 304.600 2733.085 ;
        RECT 287.565 2732.730 287.895 2732.745 ;
        RECT 297.470 2732.730 297.770 2732.785 ;
        RECT 287.565 2732.430 297.770 2732.730 ;
        RECT 287.565 2732.415 287.895 2732.430 ;
        RECT 300.000 2727.145 304.600 2727.445 ;
        RECT 287.105 2725.930 287.435 2725.945 ;
        RECT 300.230 2725.930 300.530 2727.145 ;
        RECT 287.105 2725.630 300.530 2725.930 ;
        RECT 287.105 2725.615 287.435 2725.630 ;
        RECT 284.345 2719.130 284.675 2719.145 ;
        RECT 284.345 2718.945 300.530 2719.130 ;
        RECT 284.345 2718.830 304.600 2718.945 ;
        RECT 284.345 2718.815 284.675 2718.830 ;
        RECT 300.000 2718.645 304.600 2718.830 ;
        RECT 300.000 2713.005 304.600 2713.305 ;
        RECT 286.645 2712.330 286.975 2712.345 ;
        RECT 300.230 2712.330 300.530 2713.005 ;
        RECT 286.645 2712.030 300.530 2712.330 ;
        RECT 286.645 2712.015 286.975 2712.030 ;
        RECT 300.000 2704.505 304.600 2704.805 ;
        RECT 283.885 2702.130 284.215 2702.145 ;
        RECT 300.230 2702.130 300.530 2704.505 ;
        RECT 283.885 2701.830 300.530 2702.130 ;
        RECT 283.885 2701.815 284.215 2701.830 ;
        RECT 300.000 2698.865 304.600 2699.165 ;
        RECT 285.725 2698.050 286.055 2698.065 ;
        RECT 300.230 2698.050 300.530 2698.865 ;
        RECT 285.725 2697.750 300.530 2698.050 ;
        RECT 285.725 2697.735 286.055 2697.750 ;
        RECT 300.000 2690.365 304.600 2690.665 ;
        RECT 285.265 2687.850 285.595 2687.865 ;
        RECT 300.230 2687.850 300.530 2690.365 ;
        RECT 285.265 2687.550 300.530 2687.850 ;
        RECT 285.265 2687.535 285.595 2687.550 ;
        RECT 284.805 2401.570 285.135 2401.585 ;
        RECT 284.805 2401.425 300.530 2401.570 ;
        RECT 284.805 2401.270 304.600 2401.425 ;
        RECT 284.805 2401.255 285.135 2401.270 ;
        RECT 300.000 2401.125 304.600 2401.270 ;
        RECT 299.065 2392.925 299.395 2392.940 ;
        RECT 299.065 2392.625 304.600 2392.925 ;
        RECT 299.065 2392.610 299.395 2392.625 ;
      LAYER met3 ;
        RECT 305.000 2305.000 681.480 2751.235 ;
      LAYER met3 ;
        RECT 696.965 2749.730 697.295 2749.745 ;
        RECT 685.710 2749.430 697.295 2749.730 ;
        RECT 685.710 2748.565 686.010 2749.430 ;
        RECT 696.965 2749.415 697.295 2749.430 ;
        RECT 681.880 2748.265 686.480 2748.565 ;
        RECT 947.910 2732.785 954.600 2733.085 ;
        RECT 938.465 2732.730 938.795 2732.745 ;
        RECT 947.910 2732.730 948.210 2732.785 ;
        RECT 938.465 2732.430 948.210 2732.730 ;
        RECT 938.465 2732.415 938.795 2732.430 ;
        RECT 950.000 2727.145 954.600 2727.445 ;
        RECT 938.465 2725.930 938.795 2725.945 ;
        RECT 950.670 2725.930 950.970 2727.145 ;
        RECT 938.465 2725.630 950.970 2725.930 ;
        RECT 938.465 2725.615 938.795 2725.630 ;
        RECT 938.465 2719.130 938.795 2719.145 ;
        RECT 938.465 2718.945 950.970 2719.130 ;
        RECT 938.465 2718.830 954.600 2718.945 ;
        RECT 938.465 2718.815 938.795 2718.830 ;
        RECT 950.000 2718.645 954.600 2718.830 ;
        RECT 938.465 2713.010 938.795 2713.025 ;
        RECT 950.000 2713.010 954.600 2713.305 ;
        RECT 938.465 2713.005 954.600 2713.010 ;
        RECT 938.465 2712.710 950.970 2713.005 ;
        RECT 938.465 2712.695 938.795 2712.710 ;
        RECT 950.000 2704.505 954.600 2704.805 ;
        RECT 938.925 2702.130 939.255 2702.145 ;
        RECT 950.670 2702.130 950.970 2704.505 ;
        RECT 938.925 2701.830 950.970 2702.130 ;
        RECT 938.925 2701.815 939.255 2701.830 ;
        RECT 938.465 2699.410 938.795 2699.425 ;
        RECT 938.465 2699.165 950.970 2699.410 ;
        RECT 938.465 2699.110 954.600 2699.165 ;
        RECT 938.465 2699.095 938.795 2699.110 ;
        RECT 950.000 2698.865 954.600 2699.110 ;
        RECT 950.000 2690.365 954.600 2690.665 ;
        RECT 941.685 2687.850 942.015 2687.865 ;
        RECT 950.670 2687.850 950.970 2690.365 ;
        RECT 941.685 2687.550 950.970 2687.850 ;
        RECT 941.685 2687.535 942.015 2687.550 ;
        RECT 696.965 2447.810 697.295 2447.825 ;
        RECT 685.710 2447.510 697.295 2447.810 ;
        RECT 685.710 2447.210 686.010 2447.510 ;
        RECT 696.965 2447.495 697.295 2447.510 ;
        RECT 681.880 2446.910 686.480 2447.210 ;
        RECT 685.710 2438.710 686.010 2446.910 ;
        RECT 681.880 2438.410 686.480 2438.710 ;
        RECT 685.710 2433.070 686.010 2438.410 ;
        RECT 681.880 2432.770 686.480 2433.070 ;
        RECT 685.710 2424.570 686.010 2432.770 ;
        RECT 681.880 2424.270 686.480 2424.570 ;
        RECT 685.710 2418.930 686.010 2424.270 ;
        RECT 681.880 2418.630 686.480 2418.930 ;
        RECT 685.710 2410.430 686.010 2418.630 ;
        RECT 681.880 2410.130 686.480 2410.430 ;
        RECT 685.710 2404.790 686.010 2410.130 ;
        RECT 681.880 2404.490 686.480 2404.790 ;
        RECT 944.905 2401.570 945.235 2401.585 ;
        RECT 944.905 2401.425 950.970 2401.570 ;
        RECT 944.905 2401.270 954.600 2401.425 ;
        RECT 944.905 2401.255 945.235 2401.270 ;
        RECT 950.000 2401.125 954.600 2401.270 ;
        RECT 950.000 2392.625 954.600 2392.925 ;
        RECT 944.445 2390.010 944.775 2390.025 ;
        RECT 950.670 2390.010 950.970 2392.625 ;
        RECT 944.445 2389.710 950.970 2390.010 ;
        RECT 944.445 2389.695 944.775 2389.710 ;
      LAYER met3 ;
        RECT 955.000 2305.000 1331.480 2751.235 ;
      LAYER met3 ;
        RECT 1332.225 2749.730 1332.555 2749.745 ;
        RECT 1332.225 2749.415 1332.770 2749.730 ;
        RECT 1332.470 2748.565 1332.770 2749.415 ;
        RECT 1331.880 2748.265 1336.480 2748.565 ;
        RECT 1332.470 2747.010 1332.770 2748.265 ;
        RECT 1352.005 2747.010 1352.335 2747.025 ;
        RECT 1332.470 2746.710 1352.335 2747.010 ;
        RECT 1352.005 2746.695 1352.335 2746.710 ;
        RECT 1547.750 2732.785 1554.600 2733.085 ;
        RECT 1529.105 2732.730 1529.435 2732.745 ;
        RECT 1547.750 2732.730 1548.050 2732.785 ;
        RECT 1529.105 2732.430 1548.050 2732.730 ;
        RECT 1529.105 2732.415 1529.435 2732.430 ;
        RECT 1550.000 2727.145 1554.600 2727.445 ;
        RECT 1538.305 2725.930 1538.635 2725.945 ;
        RECT 1550.510 2725.930 1550.810 2727.145 ;
        RECT 1538.305 2725.630 1550.810 2725.930 ;
        RECT 1538.305 2725.615 1538.635 2725.630 ;
        RECT 1528.645 2719.130 1528.975 2719.145 ;
        RECT 1528.645 2718.945 1550.810 2719.130 ;
        RECT 1528.645 2718.830 1554.600 2718.945 ;
        RECT 1528.645 2718.815 1528.975 2718.830 ;
        RECT 1550.000 2718.645 1554.600 2718.830 ;
        RECT 1550.000 2713.005 1554.600 2713.305 ;
        RECT 1536.005 2712.330 1536.335 2712.345 ;
        RECT 1550.510 2712.330 1550.810 2713.005 ;
        RECT 1536.005 2712.030 1550.810 2712.330 ;
        RECT 1536.005 2712.015 1536.335 2712.030 ;
        RECT 1550.000 2704.505 1554.600 2704.805 ;
        RECT 1536.465 2702.130 1536.795 2702.145 ;
        RECT 1550.510 2702.130 1550.810 2704.505 ;
        RECT 1536.465 2701.830 1550.810 2702.130 ;
        RECT 1536.465 2701.815 1536.795 2701.830 ;
        RECT 1538.305 2699.410 1538.635 2699.425 ;
        RECT 1538.305 2699.165 1550.810 2699.410 ;
        RECT 1538.305 2699.110 1554.600 2699.165 ;
        RECT 1538.305 2699.095 1538.635 2699.110 ;
        RECT 1550.000 2698.865 1554.600 2699.110 ;
        RECT 1528.185 2698.050 1528.515 2698.065 ;
        RECT 1536.465 2698.050 1536.795 2698.065 ;
        RECT 1528.185 2697.750 1536.795 2698.050 ;
        RECT 1528.185 2697.735 1528.515 2697.750 ;
        RECT 1536.465 2697.735 1536.795 2697.750 ;
        RECT 1550.000 2690.365 1554.600 2690.665 ;
        RECT 1535.085 2687.850 1535.415 2687.865 ;
        RECT 1550.510 2687.850 1550.810 2690.365 ;
        RECT 1535.085 2687.550 1550.810 2687.850 ;
        RECT 1535.085 2687.535 1535.415 2687.550 ;
        RECT 1331.880 2446.910 1336.480 2447.210 ;
        RECT 1333.390 2438.710 1333.690 2446.910 ;
        RECT 1331.880 2438.410 1336.480 2438.710 ;
        RECT 1333.390 2433.070 1333.690 2438.410 ;
        RECT 1331.880 2432.770 1336.480 2433.070 ;
        RECT 1333.390 2424.570 1333.690 2432.770 ;
        RECT 1331.880 2424.270 1336.480 2424.570 ;
        RECT 1336.150 2422.650 1336.450 2424.270 ;
        RECT 1345.565 2422.650 1345.895 2422.665 ;
        RECT 1336.150 2422.350 1345.895 2422.650 ;
        RECT 1336.150 2418.930 1336.450 2422.350 ;
        RECT 1345.565 2422.335 1345.895 2422.350 ;
        RECT 1331.880 2418.630 1336.480 2418.930 ;
        RECT 1336.150 2410.430 1336.450 2418.630 ;
        RECT 1331.880 2410.130 1336.480 2410.430 ;
        RECT 1336.150 2404.790 1336.450 2410.130 ;
        RECT 1331.880 2404.490 1336.480 2404.790 ;
        RECT 1529.565 2401.570 1529.895 2401.585 ;
        RECT 1529.565 2401.425 1550.810 2401.570 ;
        RECT 1529.565 2401.270 1554.600 2401.425 ;
        RECT 1529.565 2401.255 1529.895 2401.270 ;
        RECT 1550.000 2401.125 1554.600 2401.270 ;
        RECT 1550.000 2392.625 1554.600 2392.925 ;
        RECT 1535.545 2390.690 1535.875 2390.705 ;
        RECT 1550.510 2390.690 1550.810 2392.625 ;
        RECT 1535.545 2390.390 1550.810 2390.690 ;
        RECT 1535.545 2390.375 1535.875 2390.390 ;
      LAYER met3 ;
        RECT 1555.000 2305.000 1931.480 2751.235 ;
      LAYER met3 ;
        RECT 1945.865 2749.730 1946.195 2749.745 ;
        RECT 1935.990 2749.430 1946.195 2749.730 ;
        RECT 1935.990 2748.565 1936.290 2749.430 ;
        RECT 1945.865 2749.415 1946.195 2749.430 ;
        RECT 1931.880 2748.265 1936.480 2748.565 ;
        RECT 2197.270 2732.785 2204.600 2733.085 ;
        RECT 2187.365 2732.730 2187.695 2732.745 ;
        RECT 2197.270 2732.730 2197.570 2732.785 ;
        RECT 2187.365 2732.430 2197.570 2732.730 ;
        RECT 2187.365 2732.415 2187.695 2732.430 ;
        RECT 2200.000 2727.145 2204.600 2727.445 ;
        RECT 2187.365 2725.930 2187.695 2725.945 ;
        RECT 2200.030 2725.930 2200.330 2727.145 ;
        RECT 2187.365 2725.630 2200.330 2725.930 ;
        RECT 2187.365 2725.615 2187.695 2725.630 ;
        RECT 2187.365 2719.130 2187.695 2719.145 ;
        RECT 2187.365 2718.945 2200.330 2719.130 ;
        RECT 2187.365 2718.830 2204.600 2718.945 ;
        RECT 2187.365 2718.815 2187.695 2718.830 ;
        RECT 2200.000 2718.645 2204.600 2718.830 ;
        RECT 2200.000 2713.005 2204.600 2713.305 ;
        RECT 2187.365 2712.330 2187.695 2712.345 ;
        RECT 2200.030 2712.330 2200.330 2713.005 ;
        RECT 2187.365 2712.030 2200.330 2712.330 ;
        RECT 2187.365 2712.015 2187.695 2712.030 ;
        RECT 2200.000 2704.505 2204.600 2704.805 ;
        RECT 2187.825 2702.130 2188.155 2702.145 ;
        RECT 2200.030 2702.130 2200.330 2704.505 ;
        RECT 2187.825 2701.830 2200.330 2702.130 ;
        RECT 2187.825 2701.815 2188.155 2701.830 ;
        RECT 2187.365 2699.410 2187.695 2699.425 ;
        RECT 2187.365 2699.165 2200.330 2699.410 ;
        RECT 2187.365 2699.110 2204.600 2699.165 ;
        RECT 2187.365 2699.095 2187.695 2699.110 ;
        RECT 2200.000 2698.865 2204.600 2699.110 ;
        RECT 2200.000 2690.365 2204.600 2690.665 ;
        RECT 2187.365 2687.850 2187.695 2687.865 ;
        RECT 2200.030 2687.850 2200.330 2690.365 ;
        RECT 2187.365 2687.550 2200.330 2687.850 ;
        RECT 2187.365 2687.535 2187.695 2687.550 ;
        RECT 1945.865 2447.810 1946.195 2447.825 ;
        RECT 1935.990 2447.510 1946.195 2447.810 ;
        RECT 1935.990 2447.210 1936.290 2447.510 ;
        RECT 1945.865 2447.495 1946.195 2447.510 ;
        RECT 1931.880 2446.910 1936.480 2447.210 ;
        RECT 1935.990 2438.710 1936.290 2446.910 ;
        RECT 1931.880 2438.410 1936.480 2438.710 ;
        RECT 1935.990 2433.070 1936.290 2438.410 ;
        RECT 1931.880 2432.770 1936.480 2433.070 ;
        RECT 1935.990 2424.570 1936.290 2432.770 ;
        RECT 1931.880 2424.270 1936.480 2424.570 ;
        RECT 1935.990 2418.930 1936.290 2424.270 ;
        RECT 1931.880 2418.630 1936.480 2418.930 ;
        RECT 1935.990 2410.430 1936.290 2418.630 ;
        RECT 1931.880 2410.130 1936.480 2410.430 ;
        RECT 1935.990 2404.970 1936.290 2410.130 ;
        RECT 1945.865 2404.970 1946.195 2404.985 ;
        RECT 1935.990 2404.790 1946.195 2404.970 ;
        RECT 1931.880 2404.670 1946.195 2404.790 ;
        RECT 1931.880 2404.490 1936.480 2404.670 ;
        RECT 1945.865 2404.655 1946.195 2404.670 ;
        RECT 2187.365 2401.570 2187.695 2401.585 ;
        RECT 2187.365 2401.425 2200.330 2401.570 ;
        RECT 2187.365 2401.270 2204.600 2401.425 ;
        RECT 2187.365 2401.255 2187.695 2401.270 ;
        RECT 2200.000 2401.125 2204.600 2401.270 ;
        RECT 2200.000 2392.625 2204.600 2392.925 ;
        RECT 2190.585 2390.010 2190.915 2390.025 ;
        RECT 2200.030 2390.010 2200.330 2392.625 ;
        RECT 2190.585 2389.710 2200.330 2390.010 ;
        RECT 2190.585 2389.695 2190.915 2389.710 ;
      LAYER met3 ;
        RECT 2205.000 2305.000 2581.480 2751.235 ;
      LAYER met3 ;
        RECT 2582.045 2749.730 2582.375 2749.745 ;
        RECT 2582.045 2749.430 2583.050 2749.730 ;
        RECT 2582.045 2749.415 2582.375 2749.430 ;
        RECT 2582.750 2748.565 2583.050 2749.430 ;
        RECT 2581.880 2748.265 2586.480 2748.565 ;
        RECT 2594.465 2447.810 2594.795 2447.825 ;
        RECT 2585.510 2447.510 2594.795 2447.810 ;
        RECT 2585.510 2447.210 2585.810 2447.510 ;
        RECT 2594.465 2447.495 2594.795 2447.510 ;
        RECT 2581.880 2446.910 2586.480 2447.210 ;
        RECT 2585.510 2438.710 2585.810 2446.910 ;
        RECT 2581.880 2438.410 2586.480 2438.710 ;
        RECT 2585.510 2433.070 2585.810 2438.410 ;
        RECT 2581.880 2432.770 2586.480 2433.070 ;
        RECT 2585.510 2424.570 2585.810 2432.770 ;
        RECT 2581.880 2424.270 2586.480 2424.570 ;
        RECT 2582.750 2418.930 2583.050 2424.270 ;
        RECT 2581.880 2418.630 2586.480 2418.930 ;
        RECT 2582.750 2410.430 2583.050 2418.630 ;
        RECT 2581.880 2410.130 2586.480 2410.430 ;
        RECT 2582.750 2404.790 2583.050 2410.130 ;
        RECT 2581.880 2404.490 2586.480 2404.790 ;
        RECT 1759.105 2298.220 1759.435 2298.225 ;
        RECT 1759.105 2298.210 1759.550 2298.220 ;
        RECT 1758.740 2297.910 1759.550 2298.210 ;
        RECT 1759.105 2297.900 1759.550 2297.910 ;
        RECT 1759.105 2297.895 1759.435 2297.900 ;
        RECT 386.465 2297.540 386.795 2297.545 ;
        RECT 386.465 2297.530 386.910 2297.540 ;
        RECT 386.100 2297.230 386.910 2297.530 ;
        RECT 386.465 2297.220 386.910 2297.230 ;
        RECT 1636.530 2297.530 1636.910 2297.540 ;
        RECT 1639.505 2297.530 1639.835 2297.545 ;
        RECT 1794.065 2297.540 1794.395 2297.545 ;
        RECT 2415.065 2297.540 2415.395 2297.545 ;
        RECT 1636.530 2297.230 1639.835 2297.530 ;
        RECT 1636.530 2297.220 1636.910 2297.230 ;
        RECT 386.465 2297.215 386.795 2297.220 ;
        RECT 1639.505 2297.215 1639.835 2297.230 ;
        RECT 1642.370 2297.530 1642.750 2297.540 ;
        RECT 1644.310 2297.530 1644.690 2297.540 ;
        RECT 1794.065 2297.530 1794.590 2297.540 ;
        RECT 1642.370 2297.230 1644.690 2297.530 ;
        RECT 1793.780 2297.230 1794.590 2297.530 ;
        RECT 1642.370 2297.220 1642.750 2297.230 ;
        RECT 1644.310 2297.220 1644.690 2297.230 ;
        RECT 1794.065 2297.220 1794.590 2297.230 ;
        RECT 2263.170 2297.530 2263.550 2297.540 ;
        RECT 2265.310 2297.530 2265.690 2297.540 ;
        RECT 2263.170 2297.230 2265.690 2297.530 ;
        RECT 2263.170 2297.220 2263.550 2297.230 ;
        RECT 2265.310 2297.220 2265.690 2297.230 ;
        RECT 2415.010 2297.530 2415.395 2297.540 ;
        RECT 2415.010 2297.230 2415.820 2297.530 ;
        RECT 2415.010 2297.220 2415.395 2297.230 ;
        RECT 1794.065 2297.215 1794.395 2297.220 ;
        RECT 2415.065 2297.215 2415.395 2297.220 ;
        RECT 369.190 2290.730 369.570 2290.740 ;
        RECT 370.825 2290.730 371.155 2290.745 ;
        RECT 369.190 2290.430 371.155 2290.730 ;
        RECT 369.190 2290.420 369.570 2290.430 ;
        RECT 370.825 2290.415 371.155 2290.430 ;
        RECT 374.710 2290.730 375.090 2290.740 ;
        RECT 379.105 2290.730 379.435 2290.745 ;
        RECT 374.710 2290.430 379.435 2290.730 ;
        RECT 374.710 2290.420 375.090 2290.430 ;
        RECT 379.105 2290.415 379.435 2290.430 ;
        RECT 396.790 2290.730 397.170 2290.740 ;
        RECT 399.805 2290.730 400.135 2290.745 ;
        RECT 396.790 2290.430 400.135 2290.730 ;
        RECT 396.790 2290.420 397.170 2290.430 ;
        RECT 399.805 2290.415 400.135 2290.430 ;
        RECT 409.465 2290.740 409.795 2290.745 ;
        RECT 414.065 2290.740 414.395 2290.745 ;
        RECT 420.965 2290.740 421.295 2290.745 ;
        RECT 427.405 2290.740 427.735 2290.745 ;
        RECT 409.465 2290.730 410.050 2290.740 ;
        RECT 414.065 2290.730 414.650 2290.740 ;
        RECT 420.710 2290.730 421.295 2290.740 ;
        RECT 427.150 2290.730 427.735 2290.740 ;
        RECT 409.465 2290.430 410.250 2290.730 ;
        RECT 414.065 2290.430 414.850 2290.730 ;
        RECT 420.710 2290.430 421.520 2290.730 ;
        RECT 426.950 2290.430 427.735 2290.730 ;
        RECT 409.465 2290.420 410.050 2290.430 ;
        RECT 414.065 2290.420 414.650 2290.430 ;
        RECT 420.710 2290.420 421.295 2290.430 ;
        RECT 427.150 2290.420 427.735 2290.430 ;
        RECT 409.465 2290.415 409.795 2290.420 ;
        RECT 414.065 2290.415 414.395 2290.420 ;
        RECT 420.965 2290.415 421.295 2290.420 ;
        RECT 427.405 2290.415 427.735 2290.420 ;
        RECT 431.545 2290.740 431.875 2290.745 ;
        RECT 439.365 2290.740 439.695 2290.745 ;
        RECT 431.545 2290.730 432.130 2290.740 ;
        RECT 439.110 2290.730 439.695 2290.740 ;
        RECT 431.545 2290.430 432.330 2290.730 ;
        RECT 438.910 2290.430 439.695 2290.730 ;
        RECT 431.545 2290.420 432.130 2290.430 ;
        RECT 439.110 2290.420 439.695 2290.430 ;
        RECT 444.630 2290.730 445.010 2290.740 ;
        RECT 445.345 2290.730 445.675 2290.745 ;
        RECT 444.630 2290.430 445.675 2290.730 ;
        RECT 444.630 2290.420 445.010 2290.430 ;
        RECT 431.545 2290.415 431.875 2290.420 ;
        RECT 439.365 2290.415 439.695 2290.420 ;
        RECT 445.345 2290.415 445.675 2290.430 ;
        RECT 450.865 2290.740 451.195 2290.745 ;
        RECT 450.865 2290.730 451.450 2290.740 ;
        RECT 455.465 2290.730 455.795 2290.745 ;
        RECT 462.365 2290.740 462.695 2290.745 ;
        RECT 467.885 2290.740 468.215 2290.745 ;
        RECT 456.590 2290.730 456.970 2290.740 ;
        RECT 462.110 2290.730 462.695 2290.740 ;
        RECT 450.865 2290.430 451.650 2290.730 ;
        RECT 455.465 2290.430 456.970 2290.730 ;
        RECT 461.910 2290.430 462.695 2290.730 ;
        RECT 450.865 2290.420 451.450 2290.430 ;
        RECT 450.865 2290.415 451.195 2290.420 ;
        RECT 455.465 2290.415 455.795 2290.430 ;
        RECT 456.590 2290.420 456.970 2290.430 ;
        RECT 462.110 2290.420 462.695 2290.430 ;
        RECT 467.630 2290.730 468.215 2290.740 ;
        RECT 473.865 2290.740 474.195 2290.745 ;
        RECT 478.925 2290.740 479.255 2290.745 ;
        RECT 473.865 2290.730 474.450 2290.740 ;
        RECT 478.670 2290.730 479.255 2290.740 ;
        RECT 467.630 2290.430 468.440 2290.730 ;
        RECT 473.865 2290.430 474.650 2290.730 ;
        RECT 478.470 2290.430 479.255 2290.730 ;
        RECT 467.630 2290.420 468.215 2290.430 ;
        RECT 462.365 2290.415 462.695 2290.420 ;
        RECT 467.885 2290.415 468.215 2290.420 ;
        RECT 473.865 2290.420 474.450 2290.430 ;
        RECT 478.670 2290.420 479.255 2290.430 ;
        RECT 473.865 2290.415 474.195 2290.420 ;
        RECT 478.925 2290.415 479.255 2290.420 ;
        RECT 485.825 2290.740 486.155 2290.745 ;
        RECT 485.825 2290.730 486.410 2290.740 ;
        RECT 491.550 2290.730 491.930 2290.740 ;
        RECT 492.725 2290.730 493.055 2290.745 ;
        RECT 497.325 2290.740 497.655 2290.745 ;
        RECT 497.070 2290.730 497.655 2290.740 ;
        RECT 485.825 2290.430 486.610 2290.730 ;
        RECT 491.550 2290.430 493.055 2290.730 ;
        RECT 496.870 2290.430 497.655 2290.730 ;
        RECT 485.825 2290.420 486.410 2290.430 ;
        RECT 491.550 2290.420 491.930 2290.430 ;
        RECT 485.825 2290.415 486.155 2290.420 ;
        RECT 492.725 2290.415 493.055 2290.430 ;
        RECT 497.070 2290.420 497.655 2290.430 ;
        RECT 500.750 2290.730 501.130 2290.740 ;
        RECT 503.305 2290.730 503.635 2290.745 ;
        RECT 509.745 2290.740 510.075 2290.745 ;
        RECT 513.885 2290.740 514.215 2290.745 ;
        RECT 509.745 2290.730 510.330 2290.740 ;
        RECT 513.630 2290.730 514.215 2290.740 ;
        RECT 500.750 2290.430 503.635 2290.730 ;
        RECT 509.520 2290.430 510.330 2290.730 ;
        RECT 513.430 2290.430 514.215 2290.730 ;
        RECT 500.750 2290.420 501.130 2290.430 ;
        RECT 497.325 2290.415 497.655 2290.420 ;
        RECT 503.305 2290.415 503.635 2290.430 ;
        RECT 509.745 2290.420 510.330 2290.430 ;
        RECT 513.630 2290.420 514.215 2290.430 ;
        RECT 515.470 2290.730 515.850 2290.740 ;
        RECT 517.105 2290.730 517.435 2290.745 ;
        RECT 521.245 2290.740 521.575 2290.745 ;
        RECT 524.005 2290.740 524.335 2290.745 ;
        RECT 526.765 2290.740 527.095 2290.745 ;
        RECT 520.990 2290.730 521.575 2290.740 ;
        RECT 515.470 2290.430 517.435 2290.730 ;
        RECT 520.790 2290.430 521.575 2290.730 ;
        RECT 515.470 2290.420 515.850 2290.430 ;
        RECT 509.745 2290.415 510.075 2290.420 ;
        RECT 513.885 2290.415 514.215 2290.420 ;
        RECT 517.105 2290.415 517.435 2290.430 ;
        RECT 520.990 2290.420 521.575 2290.430 ;
        RECT 523.750 2290.730 524.335 2290.740 ;
        RECT 526.510 2290.730 527.095 2290.740 ;
        RECT 523.750 2290.430 524.560 2290.730 ;
        RECT 526.310 2290.430 527.095 2290.730 ;
        RECT 523.750 2290.420 524.335 2290.430 ;
        RECT 526.510 2290.420 527.095 2290.430 ;
        RECT 527.430 2290.730 527.810 2290.740 ;
        RECT 530.905 2290.730 531.235 2290.745 ;
        RECT 527.430 2290.430 531.235 2290.730 ;
        RECT 527.430 2290.420 527.810 2290.430 ;
        RECT 521.245 2290.415 521.575 2290.420 ;
        RECT 524.005 2290.415 524.335 2290.420 ;
        RECT 526.765 2290.415 527.095 2290.420 ;
        RECT 530.905 2290.415 531.235 2290.430 ;
        RECT 535.710 2290.730 536.090 2290.740 ;
        RECT 537.805 2290.730 538.135 2290.745 ;
        RECT 543.785 2290.740 544.115 2290.745 ;
        RECT 543.785 2290.730 544.370 2290.740 ;
        RECT 535.710 2290.430 538.135 2290.730 ;
        RECT 543.560 2290.430 544.370 2290.730 ;
        RECT 535.710 2290.420 536.090 2290.430 ;
        RECT 537.805 2290.415 538.135 2290.430 ;
        RECT 543.785 2290.420 544.370 2290.430 ;
        RECT 544.910 2290.730 545.290 2290.740 ;
        RECT 551.605 2290.730 551.935 2290.745 ;
        RECT 1001.025 2290.740 1001.355 2290.745 ;
        RECT 1052.545 2290.740 1052.875 2290.745 ;
        RECT 1001.025 2290.730 1001.610 2290.740 ;
        RECT 544.910 2290.430 551.935 2290.730 ;
        RECT 1000.800 2290.430 1001.610 2290.730 ;
        RECT 544.910 2290.420 545.290 2290.430 ;
        RECT 543.785 2290.415 544.115 2290.420 ;
        RECT 551.605 2290.415 551.935 2290.430 ;
        RECT 1001.025 2290.420 1001.610 2290.430 ;
        RECT 1052.545 2290.730 1053.130 2290.740 ;
        RECT 1060.110 2290.730 1060.490 2290.740 ;
        RECT 1062.205 2290.730 1062.535 2290.745 ;
        RECT 1052.545 2290.430 1053.330 2290.730 ;
        RECT 1060.110 2290.430 1062.535 2290.730 ;
        RECT 1052.545 2290.420 1053.130 2290.430 ;
        RECT 1060.110 2290.420 1060.490 2290.430 ;
        RECT 1001.025 2290.415 1001.355 2290.420 ;
        RECT 1052.545 2290.415 1052.875 2290.420 ;
        RECT 1062.205 2290.415 1062.535 2290.430 ;
        RECT 1065.425 2290.740 1065.755 2290.745 ;
        RECT 1070.025 2290.740 1070.355 2290.745 ;
        RECT 1076.465 2290.740 1076.795 2290.745 ;
        RECT 1083.365 2290.740 1083.695 2290.745 ;
        RECT 1087.965 2290.740 1088.295 2290.745 ;
        RECT 1094.405 2290.740 1094.735 2290.745 ;
        RECT 1100.845 2290.740 1101.175 2290.745 ;
        RECT 1065.425 2290.730 1066.010 2290.740 ;
        RECT 1070.025 2290.730 1070.610 2290.740 ;
        RECT 1076.465 2290.730 1077.050 2290.740 ;
        RECT 1083.110 2290.730 1083.695 2290.740 ;
        RECT 1087.710 2290.730 1088.295 2290.740 ;
        RECT 1094.150 2290.730 1094.735 2290.740 ;
        RECT 1100.590 2290.730 1101.175 2290.740 ;
        RECT 1065.425 2290.430 1066.210 2290.730 ;
        RECT 1070.025 2290.430 1070.810 2290.730 ;
        RECT 1076.465 2290.430 1077.250 2290.730 ;
        RECT 1082.910 2290.430 1083.695 2290.730 ;
        RECT 1087.510 2290.430 1088.295 2290.730 ;
        RECT 1093.950 2290.430 1094.735 2290.730 ;
        RECT 1100.390 2290.430 1101.175 2290.730 ;
        RECT 1065.425 2290.420 1066.010 2290.430 ;
        RECT 1070.025 2290.420 1070.610 2290.430 ;
        RECT 1076.465 2290.420 1077.050 2290.430 ;
        RECT 1083.110 2290.420 1083.695 2290.430 ;
        RECT 1087.710 2290.420 1088.295 2290.430 ;
        RECT 1094.150 2290.420 1094.735 2290.430 ;
        RECT 1100.590 2290.420 1101.175 2290.430 ;
        RECT 1065.425 2290.415 1065.755 2290.420 ;
        RECT 1070.025 2290.415 1070.355 2290.420 ;
        RECT 1076.465 2290.415 1076.795 2290.420 ;
        RECT 1083.365 2290.415 1083.695 2290.420 ;
        RECT 1087.965 2290.415 1088.295 2290.420 ;
        RECT 1094.405 2290.415 1094.735 2290.420 ;
        RECT 1100.845 2290.415 1101.175 2290.420 ;
        RECT 1106.825 2290.740 1107.155 2290.745 ;
        RECT 1112.805 2290.740 1113.135 2290.745 ;
        RECT 1118.325 2290.740 1118.655 2290.745 ;
        RECT 1106.825 2290.730 1107.410 2290.740 ;
        RECT 1112.550 2290.730 1113.135 2290.740 ;
        RECT 1118.070 2290.730 1118.655 2290.740 ;
        RECT 1106.825 2290.430 1107.610 2290.730 ;
        RECT 1112.350 2290.430 1113.135 2290.730 ;
        RECT 1117.870 2290.430 1118.655 2290.730 ;
        RECT 1106.825 2290.420 1107.410 2290.430 ;
        RECT 1112.550 2290.420 1113.135 2290.430 ;
        RECT 1118.070 2290.420 1118.655 2290.430 ;
        RECT 1106.825 2290.415 1107.155 2290.420 ;
        RECT 1112.805 2290.415 1113.135 2290.420 ;
        RECT 1118.325 2290.415 1118.655 2290.420 ;
        RECT 1121.545 2290.740 1121.875 2290.745 ;
        RECT 1129.365 2290.740 1129.695 2290.745 ;
        RECT 1135.805 2290.740 1136.135 2290.745 ;
        RECT 1121.545 2290.730 1122.130 2290.740 ;
        RECT 1129.110 2290.730 1129.695 2290.740 ;
        RECT 1135.550 2290.730 1136.135 2290.740 ;
        RECT 1121.545 2290.430 1122.330 2290.730 ;
        RECT 1128.910 2290.430 1129.695 2290.730 ;
        RECT 1135.350 2290.430 1136.135 2290.730 ;
        RECT 1121.545 2290.420 1122.130 2290.430 ;
        RECT 1129.110 2290.420 1129.695 2290.430 ;
        RECT 1135.550 2290.420 1136.135 2290.430 ;
        RECT 1121.545 2290.415 1121.875 2290.420 ;
        RECT 1129.365 2290.415 1129.695 2290.420 ;
        RECT 1135.805 2290.415 1136.135 2290.420 ;
        RECT 1141.785 2290.740 1142.115 2290.745 ;
        RECT 1147.765 2290.740 1148.095 2290.745 ;
        RECT 1141.785 2290.730 1142.370 2290.740 ;
        RECT 1147.510 2290.730 1148.095 2290.740 ;
        RECT 1141.785 2290.430 1142.570 2290.730 ;
        RECT 1147.310 2290.430 1148.095 2290.730 ;
        RECT 1141.785 2290.420 1142.370 2290.430 ;
        RECT 1147.510 2290.420 1148.095 2290.430 ;
        RECT 1141.785 2290.415 1142.115 2290.420 ;
        RECT 1147.765 2290.415 1148.095 2290.420 ;
        RECT 1159.265 2290.730 1159.595 2290.745 ;
        RECT 1164.070 2290.730 1164.450 2290.740 ;
        RECT 1159.265 2290.430 1164.450 2290.730 ;
        RECT 1159.265 2290.415 1159.595 2290.430 ;
        RECT 1164.070 2290.420 1164.450 2290.430 ;
        RECT 1166.165 2290.730 1166.495 2290.745 ;
        RECT 1167.750 2290.730 1168.130 2290.740 ;
        RECT 1166.165 2290.430 1168.130 2290.730 ;
        RECT 1166.165 2290.415 1166.495 2290.430 ;
        RECT 1167.750 2290.420 1168.130 2290.430 ;
        RECT 1607.765 2290.730 1608.095 2290.745 ;
        RECT 1613.950 2290.730 1614.330 2290.740 ;
        RECT 1607.765 2290.430 1614.330 2290.730 ;
        RECT 1607.765 2290.415 1608.095 2290.430 ;
        RECT 1613.950 2290.420 1614.330 2290.430 ;
        RECT 1614.665 2290.730 1614.995 2290.745 ;
        RECT 1619.470 2290.730 1619.850 2290.740 ;
        RECT 1614.665 2290.430 1619.850 2290.730 ;
        RECT 1614.665 2290.415 1614.995 2290.430 ;
        RECT 1619.470 2290.420 1619.850 2290.430 ;
        RECT 1628.465 2290.730 1628.795 2290.745 ;
        RECT 1631.430 2290.730 1631.810 2290.740 ;
        RECT 1628.465 2290.430 1631.810 2290.730 ;
        RECT 1628.465 2290.415 1628.795 2290.430 ;
        RECT 1631.430 2290.420 1631.810 2290.430 ;
        RECT 1635.365 2290.730 1635.695 2290.745 ;
        RECT 1636.950 2290.730 1637.330 2290.740 ;
        RECT 1635.365 2290.430 1637.330 2290.730 ;
        RECT 1635.365 2290.415 1635.695 2290.430 ;
        RECT 1636.950 2290.420 1637.330 2290.430 ;
        RECT 1644.310 2290.730 1644.690 2290.740 ;
        RECT 1645.485 2290.730 1645.815 2290.745 ;
        RECT 1644.310 2290.430 1645.815 2290.730 ;
        RECT 1644.310 2290.420 1644.690 2290.430 ;
        RECT 1645.485 2290.415 1645.815 2290.430 ;
        RECT 1649.625 2290.730 1649.955 2290.745 ;
        RECT 1659.285 2290.740 1659.615 2290.745 ;
        RECT 1665.725 2290.740 1666.055 2290.745 ;
        RECT 1670.325 2290.740 1670.655 2290.745 ;
        RECT 1676.765 2290.740 1677.095 2290.745 ;
        RECT 1654.430 2290.730 1654.810 2290.740 ;
        RECT 1659.030 2290.730 1659.615 2290.740 ;
        RECT 1665.470 2290.730 1666.055 2290.740 ;
        RECT 1670.070 2290.730 1670.655 2290.740 ;
        RECT 1649.625 2290.430 1654.810 2290.730 ;
        RECT 1658.830 2290.430 1659.615 2290.730 ;
        RECT 1665.270 2290.430 1666.055 2290.730 ;
        RECT 1669.870 2290.430 1670.655 2290.730 ;
        RECT 1649.625 2290.415 1649.955 2290.430 ;
        RECT 1654.430 2290.420 1654.810 2290.430 ;
        RECT 1659.030 2290.420 1659.615 2290.430 ;
        RECT 1665.470 2290.420 1666.055 2290.430 ;
        RECT 1670.070 2290.420 1670.655 2290.430 ;
        RECT 1676.510 2290.730 1677.095 2290.740 ;
        RECT 1682.745 2290.740 1683.075 2290.745 ;
        RECT 1682.745 2290.730 1683.330 2290.740 ;
        RECT 1688.470 2290.730 1688.850 2290.740 ;
        RECT 1690.105 2290.730 1690.435 2290.745 ;
        RECT 1695.165 2290.740 1695.495 2290.745 ;
        RECT 1694.910 2290.730 1695.495 2290.740 ;
        RECT 1676.510 2290.430 1677.320 2290.730 ;
        RECT 1682.745 2290.430 1683.530 2290.730 ;
        RECT 1688.470 2290.430 1690.435 2290.730 ;
        RECT 1694.710 2290.430 1695.495 2290.730 ;
        RECT 1676.510 2290.420 1677.095 2290.430 ;
        RECT 1659.285 2290.415 1659.615 2290.420 ;
        RECT 1665.725 2290.415 1666.055 2290.420 ;
        RECT 1670.325 2290.415 1670.655 2290.420 ;
        RECT 1676.765 2290.415 1677.095 2290.420 ;
        RECT 1682.745 2290.420 1683.330 2290.430 ;
        RECT 1688.470 2290.420 1688.850 2290.430 ;
        RECT 1682.745 2290.415 1683.075 2290.420 ;
        RECT 1690.105 2290.415 1690.435 2290.430 ;
        RECT 1694.910 2290.420 1695.495 2290.430 ;
        RECT 1695.165 2290.415 1695.495 2290.420 ;
        RECT 1699.305 2290.740 1699.635 2290.745 ;
        RECT 1706.205 2290.740 1706.535 2290.745 ;
        RECT 1699.305 2290.730 1699.890 2290.740 ;
        RECT 1705.950 2290.730 1706.535 2290.740 ;
        RECT 1699.305 2290.430 1700.090 2290.730 ;
        RECT 1705.750 2290.430 1706.535 2290.730 ;
        RECT 1699.305 2290.420 1699.890 2290.430 ;
        RECT 1705.950 2290.420 1706.535 2290.430 ;
        RECT 1699.305 2290.415 1699.635 2290.420 ;
        RECT 1706.205 2290.415 1706.535 2290.420 ;
        RECT 1711.265 2290.730 1711.595 2290.745 ;
        RECT 1713.310 2290.730 1713.690 2290.740 ;
        RECT 1711.265 2290.430 1713.690 2290.730 ;
        RECT 1711.265 2290.415 1711.595 2290.430 ;
        RECT 1713.310 2290.420 1713.690 2290.430 ;
        RECT 1718.165 2290.730 1718.495 2290.745 ;
        RECT 1723.685 2290.740 1724.015 2290.745 ;
        RECT 1719.750 2290.730 1720.130 2290.740 ;
        RECT 1723.430 2290.730 1724.015 2290.740 ;
        RECT 1718.165 2290.430 1720.130 2290.730 ;
        RECT 1723.230 2290.430 1724.015 2290.730 ;
        RECT 1718.165 2290.415 1718.495 2290.430 ;
        RECT 1719.750 2290.420 1720.130 2290.430 ;
        RECT 1723.430 2290.420 1724.015 2290.430 ;
        RECT 1723.685 2290.415 1724.015 2290.420 ;
        RECT 1725.065 2290.730 1725.395 2290.745 ;
        RECT 1730.790 2290.730 1731.170 2290.740 ;
        RECT 1725.065 2290.430 1731.170 2290.730 ;
        RECT 1725.065 2290.415 1725.395 2290.430 ;
        RECT 1730.790 2290.420 1731.170 2290.430 ;
        RECT 1731.965 2290.730 1732.295 2290.745 ;
        RECT 1736.310 2290.730 1736.690 2290.740 ;
        RECT 1731.965 2290.430 1736.690 2290.730 ;
        RECT 1731.965 2290.415 1732.295 2290.430 ;
        RECT 1736.310 2290.420 1736.690 2290.430 ;
        RECT 1738.865 2290.730 1739.195 2290.745 ;
        RECT 1741.830 2290.730 1742.210 2290.740 ;
        RECT 1738.865 2290.430 1742.210 2290.730 ;
        RECT 1738.865 2290.415 1739.195 2290.430 ;
        RECT 1741.830 2290.420 1742.210 2290.430 ;
        RECT 1745.765 2290.730 1746.095 2290.745 ;
        RECT 1748.270 2290.730 1748.650 2290.740 ;
        RECT 1745.765 2290.430 1748.650 2290.730 ;
        RECT 1745.765 2290.415 1746.095 2290.430 ;
        RECT 1748.270 2290.420 1748.650 2290.430 ;
        RECT 1759.565 2290.730 1759.895 2290.745 ;
        RECT 1764.830 2290.730 1765.210 2290.740 ;
        RECT 1759.565 2290.430 1765.210 2290.730 ;
        RECT 1759.565 2290.415 1759.895 2290.430 ;
        RECT 1764.830 2290.420 1765.210 2290.430 ;
        RECT 1766.465 2290.730 1766.795 2290.745 ;
        RECT 2308.805 2290.740 2309.135 2290.745 ;
        RECT 2315.245 2290.740 2315.575 2290.745 ;
        RECT 1767.590 2290.730 1767.970 2290.740 ;
        RECT 2308.550 2290.730 2309.135 2290.740 ;
        RECT 2314.990 2290.730 2315.575 2290.740 ;
        RECT 1766.465 2290.430 1767.970 2290.730 ;
        RECT 2308.350 2290.430 2309.135 2290.730 ;
        RECT 2314.790 2290.430 2315.575 2290.730 ;
        RECT 1766.465 2290.415 1766.795 2290.430 ;
        RECT 1767.590 2290.420 1767.970 2290.430 ;
        RECT 2308.550 2290.420 2309.135 2290.430 ;
        RECT 2314.990 2290.420 2315.575 2290.430 ;
        RECT 2321.430 2290.730 2321.810 2290.740 ;
        RECT 2324.905 2290.730 2325.235 2290.745 ;
        RECT 2321.430 2290.430 2325.235 2290.730 ;
        RECT 2321.430 2290.420 2321.810 2290.430 ;
        RECT 2308.805 2290.415 2309.135 2290.420 ;
        RECT 2315.245 2290.415 2315.575 2290.420 ;
        RECT 2324.905 2290.415 2325.235 2290.430 ;
        RECT 2325.825 2290.740 2326.155 2290.745 ;
        RECT 2343.765 2290.740 2344.095 2290.745 ;
        RECT 2325.825 2290.730 2326.410 2290.740 ;
        RECT 2343.510 2290.730 2344.095 2290.740 ;
        RECT 2325.825 2290.430 2326.610 2290.730 ;
        RECT 2343.310 2290.430 2344.095 2290.730 ;
        RECT 2325.825 2290.420 2326.410 2290.430 ;
        RECT 2343.510 2290.420 2344.095 2290.430 ;
        RECT 2325.825 2290.415 2326.155 2290.420 ;
        RECT 2343.765 2290.415 2344.095 2290.420 ;
        RECT 2349.745 2290.740 2350.075 2290.745 ;
        RECT 2349.745 2290.730 2350.330 2290.740 ;
        RECT 2356.390 2290.730 2356.770 2290.740 ;
        RECT 2358.945 2290.730 2359.275 2290.745 ;
        RECT 2361.245 2290.740 2361.575 2290.745 ;
        RECT 2360.990 2290.730 2361.575 2290.740 ;
        RECT 2349.745 2290.430 2350.530 2290.730 ;
        RECT 2356.390 2290.430 2359.275 2290.730 ;
        RECT 2360.790 2290.430 2361.575 2290.730 ;
        RECT 2349.745 2290.420 2350.330 2290.430 ;
        RECT 2356.390 2290.420 2356.770 2290.430 ;
        RECT 2349.745 2290.415 2350.075 2290.420 ;
        RECT 2358.945 2290.415 2359.275 2290.430 ;
        RECT 2360.990 2290.420 2361.575 2290.430 ;
        RECT 2361.245 2290.415 2361.575 2290.420 ;
        RECT 2367.225 2290.740 2367.555 2290.745 ;
        RECT 2374.125 2290.740 2374.455 2290.745 ;
        RECT 2367.225 2290.730 2367.810 2290.740 ;
        RECT 2373.870 2290.730 2374.455 2290.740 ;
        RECT 2367.225 2290.430 2368.010 2290.730 ;
        RECT 2373.670 2290.430 2374.455 2290.730 ;
        RECT 2367.225 2290.420 2367.810 2290.430 ;
        RECT 2373.870 2290.420 2374.455 2290.430 ;
        RECT 2367.225 2290.415 2367.555 2290.420 ;
        RECT 2374.125 2290.415 2374.455 2290.420 ;
        RECT 2377.345 2290.740 2377.675 2290.745 ;
        RECT 2384.705 2290.740 2385.035 2290.745 ;
        RECT 2391.605 2290.740 2391.935 2290.745 ;
        RECT 2397.125 2290.740 2397.455 2290.745 ;
        RECT 2377.345 2290.730 2377.930 2290.740 ;
        RECT 2384.705 2290.730 2385.290 2290.740 ;
        RECT 2391.350 2290.730 2391.935 2290.740 ;
        RECT 2396.870 2290.730 2397.455 2290.740 ;
        RECT 2415.065 2290.740 2415.395 2290.745 ;
        RECT 2415.065 2290.730 2415.650 2290.740 ;
        RECT 2377.345 2290.430 2378.130 2290.730 ;
        RECT 2384.705 2290.430 2385.490 2290.730 ;
        RECT 2391.150 2290.430 2391.935 2290.730 ;
        RECT 2396.670 2290.430 2397.455 2290.730 ;
        RECT 2414.840 2290.430 2415.650 2290.730 ;
        RECT 2377.345 2290.420 2377.930 2290.430 ;
        RECT 2384.705 2290.420 2385.290 2290.430 ;
        RECT 2391.350 2290.420 2391.935 2290.430 ;
        RECT 2396.870 2290.420 2397.455 2290.430 ;
        RECT 2377.345 2290.415 2377.675 2290.420 ;
        RECT 2384.705 2290.415 2385.035 2290.420 ;
        RECT 2391.605 2290.415 2391.935 2290.420 ;
        RECT 2397.125 2290.415 2397.455 2290.420 ;
        RECT 2415.065 2290.420 2415.650 2290.430 ;
        RECT 2415.985 2290.730 2416.315 2290.745 ;
        RECT 2420.790 2290.730 2421.170 2290.740 ;
        RECT 2415.985 2290.430 2421.170 2290.730 ;
        RECT 2415.065 2290.415 2415.395 2290.420 ;
        RECT 2415.985 2290.415 2416.315 2290.430 ;
        RECT 2420.790 2290.420 2421.170 2290.430 ;
        RECT 2421.965 2290.730 2422.295 2290.745 ;
        RECT 2427.230 2290.730 2427.610 2290.740 ;
        RECT 2421.965 2290.430 2427.610 2290.730 ;
        RECT 2421.965 2290.415 2422.295 2290.430 ;
        RECT 2427.230 2290.420 2427.610 2290.430 ;
        RECT 403.230 2290.050 403.610 2290.060 ;
        RECT 406.705 2290.050 407.035 2290.065 ;
        RECT 502.845 2290.060 503.175 2290.065 ;
        RECT 502.590 2290.050 503.175 2290.060 ;
        RECT 403.230 2289.750 407.035 2290.050 ;
        RECT 502.390 2289.750 503.175 2290.050 ;
        RECT 403.230 2289.740 403.610 2289.750 ;
        RECT 406.705 2289.735 407.035 2289.750 ;
        RECT 502.590 2289.740 503.175 2289.750 ;
        RECT 507.190 2290.050 507.570 2290.060 ;
        RECT 510.205 2290.050 510.535 2290.065 ;
        RECT 507.190 2289.750 510.535 2290.050 ;
        RECT 507.190 2289.740 507.570 2289.750 ;
        RECT 502.845 2289.735 503.175 2289.740 ;
        RECT 510.205 2289.735 510.535 2289.750 ;
        RECT 531.365 2290.050 531.695 2290.065 ;
        RECT 538.265 2290.060 538.595 2290.065 ;
        RECT 532.030 2290.050 532.410 2290.060 ;
        RECT 531.365 2289.750 532.410 2290.050 ;
        RECT 531.365 2289.735 531.695 2289.750 ;
        RECT 532.030 2289.740 532.410 2289.750 ;
        RECT 538.265 2290.050 538.850 2290.060 ;
        RECT 542.150 2290.050 542.530 2290.060 ;
        RECT 544.705 2290.050 545.035 2290.065 ;
        RECT 538.265 2289.750 539.050 2290.050 ;
        RECT 542.150 2289.750 545.035 2290.050 ;
        RECT 538.265 2289.740 538.850 2289.750 ;
        RECT 542.150 2289.740 542.530 2289.750 ;
        RECT 538.265 2289.735 538.595 2289.740 ;
        RECT 544.705 2289.735 545.035 2289.750 ;
        RECT 986.765 2290.050 987.095 2290.065 ;
        RECT 987.430 2290.050 987.810 2290.060 ;
        RECT 986.765 2289.750 987.810 2290.050 ;
        RECT 986.765 2289.735 987.095 2289.750 ;
        RECT 987.430 2289.740 987.810 2289.750 ;
        RECT 993.665 2290.050 993.995 2290.065 ;
        RECT 995.710 2290.050 996.090 2290.060 ;
        RECT 993.665 2289.750 996.090 2290.050 ;
        RECT 993.665 2289.735 993.995 2289.750 ;
        RECT 995.710 2289.740 996.090 2289.750 ;
        RECT 1035.270 2290.050 1035.650 2290.060 ;
        RECT 1038.285 2290.050 1038.615 2290.065 ;
        RECT 1041.045 2290.050 1041.375 2290.065 ;
        RECT 1173.065 2290.060 1173.395 2290.065 ;
        RECT 1173.065 2290.050 1173.650 2290.060 ;
        RECT 1035.270 2289.750 1041.375 2290.050 ;
        RECT 1172.840 2289.750 1173.650 2290.050 ;
        RECT 1035.270 2289.740 1035.650 2289.750 ;
        RECT 1038.285 2289.735 1038.615 2289.750 ;
        RECT 1041.045 2289.735 1041.375 2289.750 ;
        RECT 1173.065 2289.740 1173.650 2289.750 ;
        RECT 1610.985 2290.050 1611.315 2290.065 ;
        RECT 1617.885 2290.060 1618.215 2290.065 ;
        RECT 1613.030 2290.050 1613.410 2290.060 ;
        RECT 1617.630 2290.050 1618.215 2290.060 ;
        RECT 1610.985 2289.750 1613.410 2290.050 ;
        RECT 1617.430 2289.750 1618.215 2290.050 ;
        RECT 1173.065 2289.735 1173.395 2289.740 ;
        RECT 1610.985 2289.735 1611.315 2289.750 ;
        RECT 1613.030 2289.740 1613.410 2289.750 ;
        RECT 1617.630 2289.740 1618.215 2289.750 ;
        RECT 1617.885 2289.735 1618.215 2289.740 ;
        RECT 1646.405 2290.050 1646.735 2290.065 ;
        RECT 1712.645 2290.060 1712.975 2290.065 ;
        RECT 1647.990 2290.050 1648.370 2290.060 ;
        RECT 1712.390 2290.050 1712.975 2290.060 ;
        RECT 1646.405 2289.750 1648.370 2290.050 ;
        RECT 1712.190 2289.750 1712.975 2290.050 ;
        RECT 1646.405 2289.735 1646.735 2289.750 ;
        RECT 1647.990 2289.740 1648.370 2289.750 ;
        RECT 1712.390 2289.740 1712.975 2289.750 ;
        RECT 1717.910 2290.050 1718.290 2290.060 ;
        RECT 1721.845 2290.050 1722.175 2290.065 ;
        RECT 1717.910 2289.750 1722.175 2290.050 ;
        RECT 1717.910 2289.740 1718.290 2289.750 ;
        RECT 1712.645 2289.735 1712.975 2289.740 ;
        RECT 1721.845 2289.735 1722.175 2289.750 ;
        RECT 1729.665 2290.060 1729.995 2290.065 ;
        RECT 1734.265 2290.060 1734.595 2290.065 ;
        RECT 1741.165 2290.060 1741.495 2290.065 ;
        RECT 1729.665 2290.050 1730.250 2290.060 ;
        RECT 1734.265 2290.050 1734.850 2290.060 ;
        RECT 1740.910 2290.050 1741.495 2290.060 ;
        RECT 1729.665 2289.750 1730.450 2290.050 ;
        RECT 1734.265 2289.750 1735.050 2290.050 ;
        RECT 1740.710 2289.750 1741.495 2290.050 ;
        RECT 1729.665 2289.740 1730.250 2289.750 ;
        RECT 1734.265 2289.740 1734.850 2289.750 ;
        RECT 1740.910 2289.740 1741.495 2289.750 ;
        RECT 1729.665 2289.735 1729.995 2289.740 ;
        RECT 1734.265 2289.735 1734.595 2289.740 ;
        RECT 1741.165 2289.735 1741.495 2289.740 ;
        RECT 1746.225 2290.050 1746.555 2290.065 ;
        RECT 1752.665 2290.060 1752.995 2290.065 ;
        RECT 1747.350 2290.050 1747.730 2290.060 ;
        RECT 1752.665 2290.050 1753.250 2290.060 ;
        RECT 1746.225 2289.750 1747.730 2290.050 ;
        RECT 1752.440 2289.750 1753.250 2290.050 ;
        RECT 1746.225 2289.735 1746.555 2289.750 ;
        RECT 1747.350 2289.740 1747.730 2289.750 ;
        RECT 1752.665 2289.740 1753.250 2289.750 ;
        RECT 1780.265 2290.050 1780.595 2290.065 ;
        RECT 1782.310 2290.050 1782.690 2290.060 ;
        RECT 1780.265 2289.750 1782.690 2290.050 ;
        RECT 1752.665 2289.735 1752.995 2289.740 ;
        RECT 1780.265 2289.735 1780.595 2289.750 ;
        RECT 1782.310 2289.740 1782.690 2289.750 ;
        RECT 2297.510 2290.050 2297.890 2290.060 ;
        RECT 2300.985 2290.050 2301.315 2290.065 ;
        RECT 2297.510 2289.750 2301.315 2290.050 ;
        RECT 2297.510 2289.740 2297.890 2289.750 ;
        RECT 2300.985 2289.735 2301.315 2289.750 ;
        RECT 2338.910 2290.050 2339.290 2290.060 ;
        RECT 2340.085 2290.050 2340.415 2290.065 ;
        RECT 2338.910 2289.750 2340.415 2290.050 ;
        RECT 2338.910 2289.740 2339.290 2289.750 ;
        RECT 2340.085 2289.735 2340.415 2289.750 ;
        RECT 2402.185 2290.050 2402.515 2290.065 ;
        RECT 2403.310 2290.050 2403.690 2290.060 ;
        RECT 2402.185 2289.750 2403.690 2290.050 ;
        RECT 2402.185 2289.735 2402.515 2289.750 ;
        RECT 2403.310 2289.740 2403.690 2289.750 ;
        RECT 2435.765 2290.050 2436.095 2290.065 ;
        RECT 2438.270 2290.050 2438.650 2290.060 ;
        RECT 2435.765 2289.750 2438.650 2290.050 ;
        RECT 2435.765 2289.735 2436.095 2289.750 ;
        RECT 2438.270 2289.740 2438.650 2289.750 ;
        RECT 392.190 2289.370 392.570 2289.380 ;
        RECT 392.905 2289.370 393.235 2289.385 ;
        RECT 509.285 2289.380 509.615 2289.385 ;
        RECT 509.030 2289.370 509.615 2289.380 ;
        RECT 1159.265 2289.380 1159.595 2289.385 ;
        RECT 1159.265 2289.370 1159.850 2289.380 ;
        RECT 392.190 2289.070 393.235 2289.370 ;
        RECT 508.830 2289.070 509.615 2289.370 ;
        RECT 1159.040 2289.070 1159.850 2289.370 ;
        RECT 392.190 2289.060 392.570 2289.070 ;
        RECT 392.905 2289.055 393.235 2289.070 ;
        RECT 509.030 2289.060 509.615 2289.070 ;
        RECT 509.285 2289.055 509.615 2289.060 ;
        RECT 1159.265 2289.060 1159.850 2289.070 ;
        RECT 1179.965 2289.370 1180.295 2289.385 ;
        RECT 1587.065 2289.380 1587.395 2289.385 ;
        RECT 1182.470 2289.370 1182.850 2289.380 ;
        RECT 1587.065 2289.370 1587.650 2289.380 ;
        RECT 1179.965 2289.070 1182.850 2289.370 ;
        RECT 1586.840 2289.070 1587.650 2289.370 ;
        RECT 1159.265 2289.055 1159.595 2289.060 ;
        RECT 1179.965 2289.055 1180.295 2289.070 ;
        RECT 1182.470 2289.060 1182.850 2289.070 ;
        RECT 1587.065 2289.060 1587.650 2289.070 ;
        RECT 1624.070 2289.370 1624.450 2289.380 ;
        RECT 1624.785 2289.370 1625.115 2289.385 ;
        RECT 1624.070 2289.070 1625.115 2289.370 ;
        RECT 1624.070 2289.060 1624.450 2289.070 ;
        RECT 1587.065 2289.055 1587.395 2289.060 ;
        RECT 1624.785 2289.055 1625.115 2289.070 ;
        RECT 1630.510 2289.370 1630.890 2289.380 ;
        RECT 1631.685 2289.370 1632.015 2289.385 ;
        RECT 1652.385 2289.380 1652.715 2289.385 ;
        RECT 1652.385 2289.370 1652.970 2289.380 ;
        RECT 1630.510 2289.070 1632.015 2289.370 ;
        RECT 1652.160 2289.070 1652.970 2289.370 ;
        RECT 1630.510 2289.060 1630.890 2289.070 ;
        RECT 1631.685 2289.055 1632.015 2289.070 ;
        RECT 1652.385 2289.060 1652.970 2289.070 ;
        RECT 1775.205 2289.370 1775.535 2289.385 ;
        RECT 1775.870 2289.370 1776.250 2289.380 ;
        RECT 1775.205 2289.070 1776.250 2289.370 ;
        RECT 1652.385 2289.055 1652.715 2289.060 ;
        RECT 1775.205 2289.055 1775.535 2289.070 ;
        RECT 1775.870 2289.060 1776.250 2289.070 ;
        RECT 2290.865 2289.370 2291.195 2289.385 ;
        RECT 2292.910 2289.370 2293.290 2289.380 ;
        RECT 2290.865 2289.070 2293.290 2289.370 ;
        RECT 2290.865 2289.055 2291.195 2289.070 ;
        RECT 2292.910 2289.060 2293.290 2289.070 ;
        RECT 2332.470 2289.370 2332.850 2289.380 ;
        RECT 2333.185 2289.370 2333.515 2289.385 ;
        RECT 2332.470 2289.070 2333.515 2289.370 ;
        RECT 2332.470 2289.060 2332.850 2289.070 ;
        RECT 2333.185 2289.055 2333.515 2289.070 ;
        RECT 2394.365 2289.370 2394.695 2289.385 ;
        RECT 2397.790 2289.370 2398.170 2289.380 ;
        RECT 2394.365 2289.070 2398.170 2289.370 ;
        RECT 2394.365 2289.055 2394.695 2289.070 ;
        RECT 2397.790 2289.060 2398.170 2289.070 ;
        RECT 2402.645 2289.370 2402.975 2289.385 ;
        RECT 2404.230 2289.370 2404.610 2289.380 ;
        RECT 2402.645 2289.070 2404.610 2289.370 ;
        RECT 2402.645 2289.055 2402.975 2289.070 ;
        RECT 2404.230 2289.060 2404.610 2289.070 ;
        RECT 2421.965 2289.370 2422.295 2289.385 ;
        RECT 2423.550 2289.370 2423.930 2289.380 ;
        RECT 2421.965 2289.070 2423.930 2289.370 ;
        RECT 2421.965 2289.055 2422.295 2289.070 ;
        RECT 2423.550 2289.060 2423.930 2289.070 ;
        RECT 363.670 2288.690 364.050 2288.700 ;
        RECT 365.305 2288.690 365.635 2288.705 ;
        RECT 1007.465 2288.700 1007.795 2288.705 ;
        RECT 1048.405 2288.700 1048.735 2288.705 ;
        RECT 1007.465 2288.690 1008.050 2288.700 ;
        RECT 1048.150 2288.690 1048.735 2288.700 ;
        RECT 1186.865 2288.700 1187.195 2288.705 ;
        RECT 1186.865 2288.690 1187.450 2288.700 ;
        RECT 363.670 2288.390 365.635 2288.690 ;
        RECT 1007.240 2288.390 1008.050 2288.690 ;
        RECT 1047.950 2288.390 1048.735 2288.690 ;
        RECT 1186.640 2288.390 1187.450 2288.690 ;
        RECT 363.670 2288.380 364.050 2288.390 ;
        RECT 365.305 2288.375 365.635 2288.390 ;
        RECT 1007.465 2288.380 1008.050 2288.390 ;
        RECT 1048.150 2288.380 1048.735 2288.390 ;
        RECT 1007.465 2288.375 1007.795 2288.380 ;
        RECT 1048.405 2288.375 1048.735 2288.380 ;
        RECT 1186.865 2288.380 1187.450 2288.390 ;
        RECT 1193.765 2288.690 1194.095 2288.705 ;
        RECT 1194.430 2288.690 1194.810 2288.700 ;
        RECT 1193.765 2288.390 1194.810 2288.690 ;
        RECT 1186.865 2288.375 1187.195 2288.380 ;
        RECT 1193.765 2288.375 1194.095 2288.390 ;
        RECT 1194.430 2288.380 1194.810 2288.390 ;
        RECT 1656.065 2288.690 1656.395 2288.705 ;
        RECT 1659.950 2288.690 1660.330 2288.700 ;
        RECT 1656.065 2288.390 1660.330 2288.690 ;
        RECT 1656.065 2288.375 1656.395 2288.390 ;
        RECT 1659.950 2288.380 1660.330 2288.390 ;
        RECT 1718.625 2288.690 1718.955 2288.705 ;
        RECT 1787.165 2288.700 1787.495 2288.705 ;
        RECT 1724.350 2288.690 1724.730 2288.700 ;
        RECT 1718.625 2288.390 1724.730 2288.690 ;
        RECT 1718.625 2288.375 1718.955 2288.390 ;
        RECT 1724.350 2288.380 1724.730 2288.390 ;
        RECT 1786.910 2288.690 1787.495 2288.700 ;
        RECT 2301.905 2288.690 2302.235 2288.705 ;
        RECT 2408.165 2288.700 2408.495 2288.705 ;
        RECT 2303.950 2288.690 2304.330 2288.700 ;
        RECT 1786.910 2288.390 1787.720 2288.690 ;
        RECT 2301.905 2288.390 2304.330 2288.690 ;
        RECT 1786.910 2288.380 1787.495 2288.390 ;
        RECT 1787.165 2288.375 1787.495 2288.380 ;
        RECT 2301.905 2288.375 2302.235 2288.390 ;
        RECT 2303.950 2288.380 2304.330 2288.390 ;
        RECT 2407.910 2288.690 2408.495 2288.700 ;
        RECT 2428.865 2288.690 2429.195 2288.705 ;
        RECT 2442.665 2288.700 2442.995 2288.705 ;
        RECT 2429.990 2288.690 2430.370 2288.700 ;
        RECT 2442.665 2288.690 2443.250 2288.700 ;
        RECT 2407.910 2288.390 2408.720 2288.690 ;
        RECT 2428.865 2288.390 2430.370 2288.690 ;
        RECT 2442.440 2288.390 2443.250 2288.690 ;
        RECT 2407.910 2288.380 2408.495 2288.390 ;
        RECT 2408.165 2288.375 2408.495 2288.380 ;
        RECT 2428.865 2288.375 2429.195 2288.390 ;
        RECT 2429.990 2288.380 2430.370 2288.390 ;
        RECT 2442.665 2288.380 2443.250 2288.390 ;
        RECT 2442.665 2288.375 2442.995 2288.380 ;
        RECT 379.310 2288.010 379.690 2288.020 ;
        RECT 386.005 2288.010 386.335 2288.025 ;
        RECT 379.310 2287.710 386.335 2288.010 ;
        RECT 379.310 2287.700 379.690 2287.710 ;
        RECT 386.005 2287.695 386.335 2287.710 ;
        RECT 979.865 2288.010 980.195 2288.025 ;
        RECT 983.750 2288.010 984.130 2288.020 ;
        RECT 979.865 2287.710 984.130 2288.010 ;
        RECT 979.865 2287.695 980.195 2287.710 ;
        RECT 983.750 2287.700 984.130 2287.710 ;
        RECT 1152.365 2288.010 1152.695 2288.025 ;
        RECT 1153.030 2288.010 1153.410 2288.020 ;
        RECT 1152.365 2287.710 1153.410 2288.010 ;
        RECT 1152.365 2287.695 1152.695 2287.710 ;
        RECT 1153.030 2287.700 1153.410 2287.710 ;
        RECT 2283.965 2288.010 2284.295 2288.025 ;
        RECT 2287.390 2288.010 2287.770 2288.020 ;
        RECT 2283.965 2287.710 2287.770 2288.010 ;
        RECT 2283.965 2287.695 2284.295 2287.710 ;
        RECT 2287.390 2287.700 2287.770 2287.710 ;
        RECT 2297.765 2288.010 2298.095 2288.025 ;
        RECT 2298.430 2288.010 2298.810 2288.020 ;
        RECT 2297.765 2287.710 2298.810 2288.010 ;
        RECT 2297.765 2287.695 2298.095 2287.710 ;
        RECT 2298.430 2287.700 2298.810 2287.710 ;
        RECT 2435.765 2288.010 2436.095 2288.025 ;
        RECT 2439.190 2288.010 2439.570 2288.020 ;
        RECT 2435.765 2287.710 2439.570 2288.010 ;
        RECT 2435.765 2287.695 2436.095 2287.710 ;
        RECT 2439.190 2287.700 2439.570 2287.710 ;
        RECT 365.765 2287.330 366.095 2287.345 ;
        RECT 371.030 2287.330 371.410 2287.340 ;
        RECT 365.765 2287.030 371.410 2287.330 ;
        RECT 365.765 2287.015 366.095 2287.030 ;
        RECT 371.030 2287.020 371.410 2287.030 ;
        RECT 379.565 2287.330 379.895 2287.345 ;
        RECT 381.150 2287.330 381.530 2287.340 ;
        RECT 379.565 2287.030 381.530 2287.330 ;
        RECT 379.565 2287.015 379.895 2287.030 ;
        RECT 381.150 2287.020 381.530 2287.030 ;
        RECT 1042.630 2287.330 1043.010 2287.340 ;
        RECT 1045.185 2287.330 1045.515 2287.345 ;
        RECT 1042.630 2287.030 1045.515 2287.330 ;
        RECT 1042.630 2287.020 1043.010 2287.030 ;
        RECT 1045.185 2287.015 1045.515 2287.030 ;
        RECT 1081.270 2287.330 1081.650 2287.340 ;
        RECT 1082.905 2287.330 1083.235 2287.345 ;
        RECT 1081.270 2287.030 1083.235 2287.330 ;
        RECT 1081.270 2287.020 1081.650 2287.030 ;
        RECT 1082.905 2287.015 1083.235 2287.030 ;
        RECT 2263.265 2287.330 2263.595 2287.345 ;
        RECT 2268.990 2287.330 2269.370 2287.340 ;
        RECT 2263.265 2287.030 2269.370 2287.330 ;
        RECT 2263.265 2287.015 2263.595 2287.030 ;
        RECT 2268.990 2287.020 2269.370 2287.030 ;
        RECT 2270.165 2287.330 2270.495 2287.345 ;
        RECT 2275.430 2287.330 2275.810 2287.340 ;
        RECT 2270.165 2287.030 2275.810 2287.330 ;
        RECT 2270.165 2287.015 2270.495 2287.030 ;
        RECT 2275.430 2287.020 2275.810 2287.030 ;
        RECT 2415.065 2287.330 2415.395 2287.345 ;
        RECT 2418.030 2287.330 2418.410 2287.340 ;
        RECT 2415.065 2287.030 2418.410 2287.330 ;
        RECT 2415.065 2287.015 2415.395 2287.030 ;
        RECT 2418.030 2287.020 2418.410 2287.030 ;
        RECT 2428.865 2287.330 2429.195 2287.345 ;
        RECT 2432.750 2287.330 2433.130 2287.340 ;
        RECT 2428.865 2287.030 2433.130 2287.330 ;
        RECT 2428.865 2287.015 2429.195 2287.030 ;
        RECT 2432.750 2287.020 2433.130 2287.030 ;
        RECT 2442.665 2287.330 2442.995 2287.345 ;
        RECT 2444.710 2287.330 2445.090 2287.340 ;
        RECT 2442.665 2287.030 2445.090 2287.330 ;
        RECT 2442.665 2287.015 2442.995 2287.030 ;
        RECT 2444.710 2287.020 2445.090 2287.030 ;
        RECT 1030.670 2286.650 1031.050 2286.660 ;
        RECT 1031.385 2286.650 1031.715 2286.665 ;
        RECT 1034.145 2286.650 1034.475 2286.665 ;
        RECT 1649.165 2286.660 1649.495 2286.665 ;
        RECT 1030.670 2286.350 1034.475 2286.650 ;
        RECT 1030.670 2286.340 1031.050 2286.350 ;
        RECT 1031.385 2286.335 1031.715 2286.350 ;
        RECT 1034.145 2286.335 1034.475 2286.350 ;
        RECT 1648.910 2286.650 1649.495 2286.660 ;
        RECT 2380.565 2286.650 2380.895 2286.665 ;
        RECT 2385.830 2286.650 2386.210 2286.660 ;
        RECT 1648.910 2286.350 1649.720 2286.650 ;
        RECT 2380.565 2286.350 2386.210 2286.650 ;
        RECT 1648.910 2286.340 1649.495 2286.350 ;
        RECT 1649.165 2286.335 1649.495 2286.340 ;
        RECT 2380.565 2286.335 2380.895 2286.350 ;
        RECT 2385.830 2286.340 2386.210 2286.350 ;
        RECT 2387.465 2286.650 2387.795 2286.665 ;
        RECT 2392.270 2286.650 2392.650 2286.660 ;
        RECT 2387.465 2286.350 2392.650 2286.650 ;
        RECT 2387.465 2286.335 2387.795 2286.350 ;
        RECT 2392.270 2286.340 2392.650 2286.350 ;
        RECT 358.865 2285.970 359.195 2285.985 ;
        RECT 386.465 2285.980 386.795 2285.985 ;
        RECT 364.590 2285.970 364.970 2285.980 ;
        RECT 386.465 2285.970 387.050 2285.980 ;
        RECT 358.865 2285.670 364.970 2285.970 ;
        RECT 386.240 2285.670 387.050 2285.970 ;
        RECT 358.865 2285.655 359.195 2285.670 ;
        RECT 364.590 2285.660 364.970 2285.670 ;
        RECT 386.465 2285.660 387.050 2285.670 ;
        RECT 474.990 2285.970 475.370 2285.980 ;
        RECT 475.705 2285.970 476.035 2285.985 ;
        RECT 474.990 2285.670 476.035 2285.970 ;
        RECT 474.990 2285.660 475.370 2285.670 ;
        RECT 386.465 2285.655 386.795 2285.660 ;
        RECT 475.705 2285.655 476.035 2285.670 ;
        RECT 492.470 2285.970 492.850 2285.980 ;
        RECT 496.405 2285.970 496.735 2285.985 ;
        RECT 492.470 2285.670 496.735 2285.970 ;
        RECT 492.470 2285.660 492.850 2285.670 ;
        RECT 496.405 2285.655 496.735 2285.670 ;
        RECT 1010.685 2285.970 1011.015 2285.985 ;
        RECT 1012.270 2285.970 1012.650 2285.980 ;
        RECT 1010.685 2285.670 1012.650 2285.970 ;
        RECT 1010.685 2285.655 1011.015 2285.670 ;
        RECT 1012.270 2285.660 1012.650 2285.670 ;
        RECT 1013.190 2285.970 1013.570 2285.980 ;
        RECT 1013.905 2285.970 1014.235 2285.985 ;
        RECT 1013.190 2285.670 1014.235 2285.970 ;
        RECT 1013.190 2285.660 1013.570 2285.670 ;
        RECT 1013.905 2285.655 1014.235 2285.670 ;
        RECT 1031.590 2285.970 1031.970 2285.980 ;
        RECT 1034.605 2285.970 1034.935 2285.985 ;
        RECT 1031.590 2285.670 1034.935 2285.970 ;
        RECT 1031.590 2285.660 1031.970 2285.670 ;
        RECT 1034.605 2285.655 1034.935 2285.670 ;
        RECT 1049.070 2285.970 1049.450 2285.980 ;
        RECT 1054.845 2285.970 1055.175 2285.985 ;
        RECT 1049.070 2285.670 1055.175 2285.970 ;
        RECT 1049.070 2285.660 1049.450 2285.670 ;
        RECT 1054.845 2285.655 1055.175 2285.670 ;
        RECT 1072.070 2285.970 1072.450 2285.980 ;
        RECT 1076.005 2285.970 1076.335 2285.985 ;
        RECT 1072.070 2285.670 1076.335 2285.970 ;
        RECT 1072.070 2285.660 1072.450 2285.670 ;
        RECT 1076.005 2285.655 1076.335 2285.670 ;
        RECT 1084.030 2285.970 1084.410 2285.980 ;
        RECT 1089.805 2285.970 1090.135 2285.985 ;
        RECT 1084.030 2285.670 1090.135 2285.970 ;
        RECT 1084.030 2285.660 1084.410 2285.670 ;
        RECT 1089.805 2285.655 1090.135 2285.670 ;
        RECT 1101.510 2285.970 1101.890 2285.980 ;
        RECT 1103.605 2285.970 1103.935 2285.985 ;
        RECT 1101.510 2285.670 1103.935 2285.970 ;
        RECT 1101.510 2285.660 1101.890 2285.670 ;
        RECT 1103.605 2285.655 1103.935 2285.670 ;
        RECT 1621.565 2285.970 1621.895 2285.985 ;
        RECT 1642.265 2285.980 1642.595 2285.985 ;
        RECT 1624.990 2285.970 1625.370 2285.980 ;
        RECT 1642.265 2285.970 1642.850 2285.980 ;
        RECT 1621.565 2285.670 1625.370 2285.970 ;
        RECT 1642.040 2285.670 1642.850 2285.970 ;
        RECT 1621.565 2285.655 1621.895 2285.670 ;
        RECT 1624.990 2285.660 1625.370 2285.670 ;
        RECT 1642.265 2285.660 1642.850 2285.670 ;
        RECT 1676.765 2285.970 1677.095 2285.985 ;
        RECT 1677.430 2285.970 1677.810 2285.980 ;
        RECT 1676.765 2285.670 1677.810 2285.970 ;
        RECT 1642.265 2285.655 1642.595 2285.660 ;
        RECT 1676.765 2285.655 1677.095 2285.670 ;
        RECT 1677.430 2285.660 1677.810 2285.670 ;
        RECT 1704.365 2285.970 1704.695 2285.985 ;
        RECT 1706.870 2285.970 1707.250 2285.980 ;
        RECT 1704.365 2285.670 1707.250 2285.970 ;
        RECT 1704.365 2285.655 1704.695 2285.670 ;
        RECT 1706.870 2285.660 1707.250 2285.670 ;
        RECT 1766.465 2285.970 1766.795 2285.985 ;
        RECT 1771.270 2285.970 1771.650 2285.980 ;
        RECT 1766.465 2285.670 1771.650 2285.970 ;
        RECT 1766.465 2285.655 1766.795 2285.670 ;
        RECT 1771.270 2285.660 1771.650 2285.670 ;
        RECT 2252.685 2285.970 2253.015 2285.985 ;
        RECT 2273.385 2285.980 2273.715 2285.985 ;
        RECT 2257.030 2285.970 2257.410 2285.980 ;
        RECT 2252.685 2285.670 2257.410 2285.970 ;
        RECT 2252.685 2285.655 2253.015 2285.670 ;
        RECT 2257.030 2285.660 2257.410 2285.670 ;
        RECT 2273.385 2285.970 2273.970 2285.980 ;
        RECT 2291.070 2285.970 2291.450 2285.980 ;
        RECT 2294.085 2285.970 2294.415 2285.985 ;
        RECT 2296.845 2285.970 2297.175 2285.985 ;
        RECT 2273.385 2285.670 2274.170 2285.970 ;
        RECT 2291.070 2285.670 2297.175 2285.970 ;
        RECT 2273.385 2285.660 2273.970 2285.670 ;
        RECT 2291.070 2285.660 2291.450 2285.670 ;
        RECT 2273.385 2285.655 2273.715 2285.660 ;
        RECT 2294.085 2285.655 2294.415 2285.670 ;
        RECT 2296.845 2285.655 2297.175 2285.670 ;
        RECT 2305.125 2285.970 2305.455 2285.985 ;
        RECT 2310.390 2285.970 2310.770 2285.980 ;
        RECT 2305.125 2285.670 2310.770 2285.970 ;
        RECT 2305.125 2285.655 2305.455 2285.670 ;
        RECT 2310.390 2285.660 2310.770 2285.670 ;
        RECT 2339.625 2285.970 2339.955 2285.985 ;
        RECT 2345.350 2285.970 2345.730 2285.980 ;
        RECT 2339.625 2285.670 2345.730 2285.970 ;
        RECT 2339.625 2285.655 2339.955 2285.670 ;
        RECT 2345.350 2285.660 2345.730 2285.670 ;
        RECT 2359.865 2285.970 2360.195 2285.985 ;
        RECT 2362.830 2285.970 2363.210 2285.980 ;
        RECT 2359.865 2285.670 2363.210 2285.970 ;
        RECT 2359.865 2285.655 2360.195 2285.670 ;
        RECT 2362.830 2285.660 2363.210 2285.670 ;
        RECT 2380.310 2285.970 2380.690 2285.980 ;
        RECT 2381.025 2285.970 2381.355 2285.985 ;
        RECT 2380.310 2285.670 2381.355 2285.970 ;
        RECT 2380.310 2285.660 2380.690 2285.670 ;
        RECT 2381.025 2285.655 2381.355 2285.670 ;
        RECT 2408.165 2285.970 2408.495 2285.985 ;
        RECT 2409.750 2285.970 2410.130 2285.980 ;
        RECT 2408.165 2285.670 2410.130 2285.970 ;
        RECT 2408.165 2285.655 2408.495 2285.670 ;
        RECT 2409.750 2285.660 2410.130 2285.670 ;
        RECT 351.045 2285.300 351.375 2285.305 ;
        RECT 350.790 2285.290 351.375 2285.300 ;
        RECT 373.585 2285.290 373.915 2285.305 ;
        RECT 375.630 2285.290 376.010 2285.300 ;
        RECT 350.790 2284.990 351.600 2285.290 ;
        RECT 373.585 2284.990 376.010 2285.290 ;
        RECT 350.790 2284.980 351.375 2284.990 ;
        RECT 351.045 2284.975 351.375 2284.980 ;
        RECT 373.585 2284.975 373.915 2284.990 ;
        RECT 375.630 2284.980 376.010 2284.990 ;
        RECT 393.110 2285.290 393.490 2285.300 ;
        RECT 393.825 2285.290 394.155 2285.305 ;
        RECT 393.110 2284.990 394.155 2285.290 ;
        RECT 393.110 2284.980 393.490 2284.990 ;
        RECT 393.825 2284.975 394.155 2284.990 ;
        RECT 465.790 2285.290 466.170 2285.300 ;
        RECT 468.805 2285.290 469.135 2285.305 ;
        RECT 465.790 2284.990 469.135 2285.290 ;
        RECT 465.790 2284.980 466.170 2284.990 ;
        RECT 468.805 2284.975 469.135 2284.990 ;
        RECT 1024.485 2285.290 1024.815 2285.305 ;
        RECT 1025.150 2285.290 1025.530 2285.300 ;
        RECT 1027.245 2285.290 1027.575 2285.305 ;
        RECT 1024.485 2284.990 1027.575 2285.290 ;
        RECT 1024.485 2284.975 1024.815 2284.990 ;
        RECT 1025.150 2284.980 1025.530 2284.990 ;
        RECT 1027.245 2284.975 1027.575 2284.990 ;
        RECT 1128.190 2285.290 1128.570 2285.300 ;
        RECT 1131.205 2285.290 1131.535 2285.305 ;
        RECT 1128.190 2284.990 1131.535 2285.290 ;
        RECT 1128.190 2284.980 1128.570 2284.990 ;
        RECT 1131.205 2284.975 1131.535 2284.990 ;
        RECT 1163.150 2285.290 1163.530 2285.300 ;
        RECT 1165.245 2285.290 1165.575 2285.305 ;
        RECT 1163.150 2284.990 1165.575 2285.290 ;
        RECT 1163.150 2284.980 1163.530 2284.990 ;
        RECT 1165.245 2284.975 1165.575 2284.990 ;
        RECT 1601.325 2285.290 1601.655 2285.305 ;
        RECT 1604.750 2285.290 1605.130 2285.300 ;
        RECT 1601.325 2284.990 1605.130 2285.290 ;
        RECT 1601.325 2284.975 1601.655 2284.990 ;
        RECT 1604.750 2284.980 1605.130 2284.990 ;
        RECT 1684.125 2285.290 1684.455 2285.305 ;
        RECT 1689.390 2285.290 1689.770 2285.300 ;
        RECT 1684.125 2284.990 1689.770 2285.290 ;
        RECT 1684.125 2284.975 1684.455 2284.990 ;
        RECT 1689.390 2284.980 1689.770 2284.990 ;
        RECT 1760.025 2285.290 1760.355 2285.305 ;
        RECT 1765.750 2285.290 1766.130 2285.300 ;
        RECT 1760.025 2284.990 1766.130 2285.290 ;
        RECT 1760.025 2284.975 1760.355 2284.990 ;
        RECT 1765.750 2284.980 1766.130 2284.990 ;
        RECT 2231.985 2285.290 2232.315 2285.305 ;
        RECT 2280.285 2285.300 2280.615 2285.305 ;
        RECT 2239.550 2285.290 2239.930 2285.300 ;
        RECT 2280.030 2285.290 2280.615 2285.300 ;
        RECT 2283.505 2285.290 2283.835 2285.305 ;
        RECT 2231.985 2284.990 2239.930 2285.290 ;
        RECT 2279.650 2284.990 2283.835 2285.290 ;
        RECT 2231.985 2284.975 2232.315 2284.990 ;
        RECT 2239.550 2284.980 2239.930 2284.990 ;
        RECT 2280.030 2284.980 2280.615 2284.990 ;
        RECT 2280.285 2284.975 2280.615 2284.980 ;
        RECT 2283.505 2284.975 2283.835 2284.990 ;
        RECT 334.230 2284.610 334.610 2284.620 ;
        RECT 337.705 2284.610 338.035 2284.625 ;
        RECT 334.230 2284.310 338.035 2284.610 ;
        RECT 334.230 2284.300 334.610 2284.310 ;
        RECT 337.705 2284.295 338.035 2284.310 ;
        RECT 339.750 2284.610 340.130 2284.620 ;
        RECT 344.145 2284.610 344.475 2284.625 ;
        RECT 339.750 2284.310 344.475 2284.610 ;
        RECT 339.750 2284.300 340.130 2284.310 ;
        RECT 344.145 2284.295 344.475 2284.310 ;
        RECT 348.950 2284.610 349.330 2284.620 ;
        RECT 350.585 2284.610 350.915 2284.625 ;
        RECT 348.950 2284.310 350.915 2284.610 ;
        RECT 348.950 2284.300 349.330 2284.310 ;
        RECT 350.585 2284.295 350.915 2284.310 ;
        RECT 357.230 2284.610 357.610 2284.620 ;
        RECT 358.405 2284.610 358.735 2284.625 ;
        RECT 357.230 2284.310 358.735 2284.610 ;
        RECT 357.230 2284.300 357.610 2284.310 ;
        RECT 358.405 2284.295 358.735 2284.310 ;
        RECT 393.365 2284.610 393.695 2284.625 ;
        RECT 398.630 2284.610 399.010 2284.620 ;
        RECT 393.365 2284.310 399.010 2284.610 ;
        RECT 393.365 2284.295 393.695 2284.310 ;
        RECT 398.630 2284.300 399.010 2284.310 ;
        RECT 400.265 2284.610 400.595 2284.625 ;
        RECT 404.150 2284.610 404.530 2284.620 ;
        RECT 400.265 2284.310 404.530 2284.610 ;
        RECT 400.265 2284.295 400.595 2284.310 ;
        RECT 404.150 2284.300 404.530 2284.310 ;
        RECT 407.165 2284.610 407.495 2284.625 ;
        RECT 410.590 2284.610 410.970 2284.620 ;
        RECT 407.165 2284.310 410.970 2284.610 ;
        RECT 407.165 2284.295 407.495 2284.310 ;
        RECT 410.590 2284.300 410.970 2284.310 ;
        RECT 414.065 2284.610 414.395 2284.625 ;
        RECT 416.110 2284.610 416.490 2284.620 ;
        RECT 414.065 2284.310 416.490 2284.610 ;
        RECT 414.065 2284.295 414.395 2284.310 ;
        RECT 416.110 2284.300 416.490 2284.310 ;
        RECT 420.965 2284.610 421.295 2284.625 ;
        RECT 421.630 2284.610 422.010 2284.620 ;
        RECT 420.965 2284.310 422.010 2284.610 ;
        RECT 420.965 2284.295 421.295 2284.310 ;
        RECT 421.630 2284.300 422.010 2284.310 ;
        RECT 428.070 2284.610 428.450 2284.620 ;
        RECT 431.085 2284.610 431.415 2284.625 ;
        RECT 428.070 2284.310 431.415 2284.610 ;
        RECT 428.070 2284.300 428.450 2284.310 ;
        RECT 431.085 2284.295 431.415 2284.310 ;
        RECT 433.590 2284.610 433.970 2284.620 ;
        RECT 434.305 2284.610 434.635 2284.625 ;
        RECT 433.590 2284.310 434.635 2284.610 ;
        RECT 433.590 2284.300 433.970 2284.310 ;
        RECT 434.305 2284.295 434.635 2284.310 ;
        RECT 440.030 2284.610 440.410 2284.620 ;
        RECT 441.205 2284.610 441.535 2284.625 ;
        RECT 440.030 2284.310 441.535 2284.610 ;
        RECT 440.030 2284.300 440.410 2284.310 ;
        RECT 441.205 2284.295 441.535 2284.310 ;
        RECT 445.550 2284.610 445.930 2284.620 ;
        RECT 448.105 2284.610 448.435 2284.625 ;
        RECT 445.550 2284.310 448.435 2284.610 ;
        RECT 445.550 2284.300 445.930 2284.310 ;
        RECT 448.105 2284.295 448.435 2284.310 ;
        RECT 452.910 2284.610 453.290 2284.620 ;
        RECT 455.005 2284.610 455.335 2284.625 ;
        RECT 452.910 2284.310 455.335 2284.610 ;
        RECT 452.910 2284.300 453.290 2284.310 ;
        RECT 455.005 2284.295 455.335 2284.310 ;
        RECT 457.510 2284.610 457.890 2284.620 ;
        RECT 461.905 2284.610 462.235 2284.625 ;
        RECT 468.345 2284.620 468.675 2284.625 ;
        RECT 468.345 2284.610 468.930 2284.620 ;
        RECT 457.510 2284.310 462.235 2284.610 ;
        RECT 468.120 2284.310 468.930 2284.610 ;
        RECT 457.510 2284.300 457.890 2284.310 ;
        RECT 461.905 2284.295 462.235 2284.310 ;
        RECT 468.345 2284.300 468.930 2284.310 ;
        RECT 480.510 2284.610 480.890 2284.620 ;
        RECT 482.605 2284.610 482.935 2284.625 ;
        RECT 480.510 2284.310 482.935 2284.610 ;
        RECT 480.510 2284.300 480.890 2284.310 ;
        RECT 468.345 2284.295 468.675 2284.300 ;
        RECT 482.605 2284.295 482.935 2284.310 ;
        RECT 488.790 2284.610 489.170 2284.620 ;
        RECT 489.505 2284.610 489.835 2284.625 ;
        RECT 488.790 2284.310 489.835 2284.610 ;
        RECT 488.790 2284.300 489.170 2284.310 ;
        RECT 489.505 2284.295 489.835 2284.310 ;
        RECT 1017.585 2284.610 1017.915 2284.625 ;
        RECT 1018.710 2284.610 1019.090 2284.620 ;
        RECT 1017.585 2284.310 1019.090 2284.610 ;
        RECT 1017.585 2284.295 1017.915 2284.310 ;
        RECT 1018.710 2284.300 1019.090 2284.310 ;
        RECT 1019.630 2284.610 1020.010 2284.620 ;
        RECT 1020.805 2284.610 1021.135 2284.625 ;
        RECT 1019.630 2284.310 1021.135 2284.610 ;
        RECT 1019.630 2284.300 1020.010 2284.310 ;
        RECT 1020.805 2284.295 1021.135 2284.310 ;
        RECT 1026.990 2284.610 1027.370 2284.620 ;
        RECT 1027.705 2284.610 1028.035 2284.625 ;
        RECT 1026.990 2284.310 1028.035 2284.610 ;
        RECT 1026.990 2284.300 1027.370 2284.310 ;
        RECT 1027.705 2284.295 1028.035 2284.310 ;
        RECT 1037.110 2284.610 1037.490 2284.620 ;
        RECT 1041.505 2284.610 1041.835 2284.625 ;
        RECT 1037.110 2284.310 1041.835 2284.610 ;
        RECT 1037.110 2284.300 1037.490 2284.310 ;
        RECT 1041.505 2284.295 1041.835 2284.310 ;
        RECT 1046.310 2284.610 1046.690 2284.620 ;
        RECT 1048.405 2284.610 1048.735 2284.625 ;
        RECT 1046.310 2284.310 1048.735 2284.610 ;
        RECT 1046.310 2284.300 1046.690 2284.310 ;
        RECT 1048.405 2284.295 1048.735 2284.310 ;
        RECT 1054.590 2284.610 1054.970 2284.620 ;
        RECT 1055.305 2284.610 1055.635 2284.625 ;
        RECT 1062.205 2284.620 1062.535 2284.625 ;
        RECT 1054.590 2284.310 1055.635 2284.610 ;
        RECT 1054.590 2284.300 1054.970 2284.310 ;
        RECT 1055.305 2284.295 1055.635 2284.310 ;
        RECT 1061.950 2284.610 1062.535 2284.620 ;
        RECT 1066.550 2284.610 1066.930 2284.620 ;
        RECT 1069.105 2284.610 1069.435 2284.625 ;
        RECT 1089.345 2284.620 1089.675 2284.625 ;
        RECT 1089.345 2284.610 1089.930 2284.620 ;
        RECT 1061.950 2284.310 1062.760 2284.610 ;
        RECT 1066.550 2284.310 1069.435 2284.610 ;
        RECT 1089.120 2284.310 1089.930 2284.610 ;
        RECT 1061.950 2284.300 1062.535 2284.310 ;
        RECT 1066.550 2284.300 1066.930 2284.310 ;
        RECT 1062.205 2284.295 1062.535 2284.300 ;
        RECT 1069.105 2284.295 1069.435 2284.310 ;
        RECT 1089.345 2284.300 1089.930 2284.310 ;
        RECT 1095.990 2284.610 1096.370 2284.620 ;
        RECT 1096.705 2284.610 1097.035 2284.625 ;
        RECT 1095.990 2284.310 1097.035 2284.610 ;
        RECT 1095.990 2284.300 1096.370 2284.310 ;
        RECT 1089.345 2284.295 1089.675 2284.300 ;
        RECT 1096.705 2284.295 1097.035 2284.310 ;
        RECT 1109.790 2284.610 1110.170 2284.620 ;
        RECT 1110.505 2284.610 1110.835 2284.625 ;
        RECT 1109.790 2284.310 1110.835 2284.610 ;
        RECT 1109.790 2284.300 1110.170 2284.310 ;
        RECT 1110.505 2284.295 1110.835 2284.310 ;
        RECT 1116.230 2284.610 1116.610 2284.620 ;
        RECT 1117.405 2284.610 1117.735 2284.625 ;
        RECT 1116.230 2284.310 1117.735 2284.610 ;
        RECT 1116.230 2284.300 1116.610 2284.310 ;
        RECT 1117.405 2284.295 1117.735 2284.310 ;
        RECT 1118.990 2284.610 1119.370 2284.620 ;
        RECT 1124.305 2284.610 1124.635 2284.625 ;
        RECT 1130.745 2284.620 1131.075 2284.625 ;
        RECT 1130.745 2284.610 1131.330 2284.620 ;
        RECT 1118.990 2284.310 1124.635 2284.610 ;
        RECT 1130.520 2284.310 1131.330 2284.610 ;
        RECT 1118.990 2284.300 1119.370 2284.310 ;
        RECT 1124.305 2284.295 1124.635 2284.310 ;
        RECT 1130.745 2284.300 1131.330 2284.310 ;
        RECT 1136.470 2284.610 1136.850 2284.620 ;
        RECT 1138.105 2284.610 1138.435 2284.625 ;
        RECT 1145.005 2284.620 1145.335 2284.625 ;
        RECT 1144.750 2284.610 1145.335 2284.620 ;
        RECT 1136.470 2284.310 1138.435 2284.610 ;
        RECT 1144.550 2284.310 1145.335 2284.610 ;
        RECT 1136.470 2284.300 1136.850 2284.310 ;
        RECT 1130.745 2284.295 1131.075 2284.300 ;
        RECT 1138.105 2284.295 1138.435 2284.310 ;
        RECT 1144.750 2284.300 1145.335 2284.310 ;
        RECT 1148.430 2284.610 1148.810 2284.620 ;
        RECT 1151.905 2284.610 1152.235 2284.625 ;
        RECT 1148.430 2284.310 1152.235 2284.610 ;
        RECT 1148.430 2284.300 1148.810 2284.310 ;
        RECT 1145.005 2284.295 1145.335 2284.300 ;
        RECT 1151.905 2284.295 1152.235 2284.310 ;
        RECT 1153.950 2284.610 1154.330 2284.620 ;
        RECT 1158.805 2284.610 1159.135 2284.625 ;
        RECT 1153.950 2284.310 1159.135 2284.610 ;
        RECT 1153.950 2284.300 1154.330 2284.310 ;
        RECT 1158.805 2284.295 1159.135 2284.310 ;
        RECT 1164.990 2284.610 1165.370 2284.620 ;
        RECT 1165.705 2284.610 1166.035 2284.625 ;
        RECT 1164.990 2284.310 1166.035 2284.610 ;
        RECT 1164.990 2284.300 1165.370 2284.310 ;
        RECT 1165.705 2284.295 1166.035 2284.310 ;
        RECT 1171.430 2284.610 1171.810 2284.620 ;
        RECT 1172.605 2284.610 1172.935 2284.625 ;
        RECT 1171.430 2284.310 1172.935 2284.610 ;
        RECT 1171.430 2284.300 1171.810 2284.310 ;
        RECT 1172.605 2284.295 1172.935 2284.310 ;
        RECT 1178.790 2284.610 1179.170 2284.620 ;
        RECT 1179.505 2284.610 1179.835 2284.625 ;
        RECT 1178.790 2284.310 1179.835 2284.610 ;
        RECT 1178.790 2284.300 1179.170 2284.310 ;
        RECT 1179.505 2284.295 1179.835 2284.310 ;
        RECT 1183.390 2284.610 1183.770 2284.620 ;
        RECT 1186.405 2284.610 1186.735 2284.625 ;
        RECT 1183.390 2284.310 1186.735 2284.610 ;
        RECT 1183.390 2284.300 1183.770 2284.310 ;
        RECT 1186.405 2284.295 1186.735 2284.310 ;
        RECT 1188.910 2284.610 1189.290 2284.620 ;
        RECT 1193.305 2284.610 1193.635 2284.625 ;
        RECT 1188.910 2284.310 1193.635 2284.610 ;
        RECT 1188.910 2284.300 1189.290 2284.310 ;
        RECT 1193.305 2284.295 1193.635 2284.310 ;
        RECT 1198.110 2284.610 1198.490 2284.620 ;
        RECT 1200.205 2284.610 1200.535 2284.625 ;
        RECT 1198.110 2284.310 1200.535 2284.610 ;
        RECT 1198.110 2284.300 1198.490 2284.310 ;
        RECT 1200.205 2284.295 1200.535 2284.310 ;
        RECT 1580.165 2284.610 1580.495 2284.625 ;
        RECT 1580.830 2284.610 1581.210 2284.620 ;
        RECT 1580.165 2284.310 1581.210 2284.610 ;
        RECT 1580.165 2284.295 1580.495 2284.310 ;
        RECT 1580.830 2284.300 1581.210 2284.310 ;
        RECT 1593.965 2284.610 1594.295 2284.625 ;
        RECT 1600.865 2284.620 1601.195 2284.625 ;
        RECT 1595.550 2284.610 1595.930 2284.620 ;
        RECT 1600.865 2284.610 1601.450 2284.620 ;
        RECT 1593.965 2284.310 1595.930 2284.610 ;
        RECT 1600.640 2284.310 1601.450 2284.610 ;
        RECT 1593.965 2284.295 1594.295 2284.310 ;
        RECT 1595.550 2284.300 1595.930 2284.310 ;
        RECT 1600.865 2284.300 1601.450 2284.310 ;
        RECT 1662.965 2284.610 1663.295 2284.625 ;
        RECT 1666.390 2284.610 1666.770 2284.620 ;
        RECT 1662.965 2284.310 1666.770 2284.610 ;
        RECT 1600.865 2284.295 1601.195 2284.300 ;
        RECT 1662.965 2284.295 1663.295 2284.310 ;
        RECT 1666.390 2284.300 1666.770 2284.310 ;
        RECT 1669.865 2284.610 1670.195 2284.625 ;
        RECT 1683.665 2284.620 1683.995 2284.625 ;
        RECT 1671.910 2284.610 1672.290 2284.620 ;
        RECT 1683.665 2284.610 1684.250 2284.620 ;
        RECT 1669.865 2284.310 1672.290 2284.610 ;
        RECT 1683.440 2284.310 1684.250 2284.610 ;
        RECT 1669.865 2284.295 1670.195 2284.310 ;
        RECT 1671.910 2284.300 1672.290 2284.310 ;
        RECT 1683.665 2284.300 1684.250 2284.310 ;
        RECT 1690.565 2284.610 1690.895 2284.625 ;
        RECT 1695.830 2284.610 1696.210 2284.620 ;
        RECT 1690.565 2284.310 1696.210 2284.610 ;
        RECT 1683.665 2284.295 1683.995 2284.300 ;
        RECT 1690.565 2284.295 1690.895 2284.310 ;
        RECT 1695.830 2284.300 1696.210 2284.310 ;
        RECT 1697.465 2284.610 1697.795 2284.625 ;
        RECT 1701.350 2284.610 1701.730 2284.620 ;
        RECT 1697.465 2284.310 1701.730 2284.610 ;
        RECT 1697.465 2284.295 1697.795 2284.310 ;
        RECT 1701.350 2284.300 1701.730 2284.310 ;
        RECT 1752.665 2284.610 1752.995 2284.625 ;
        RECT 1759.565 2284.620 1759.895 2284.625 ;
        RECT 1754.710 2284.610 1755.090 2284.620 ;
        RECT 1752.665 2284.310 1755.090 2284.610 ;
        RECT 1752.665 2284.295 1752.995 2284.310 ;
        RECT 1754.710 2284.300 1755.090 2284.310 ;
        RECT 1759.310 2284.610 1759.895 2284.620 ;
        RECT 1773.365 2284.610 1773.695 2284.625 ;
        RECT 1776.790 2284.610 1777.170 2284.620 ;
        RECT 1759.310 2284.310 1760.120 2284.610 ;
        RECT 1773.365 2284.310 1777.170 2284.610 ;
        RECT 1759.310 2284.300 1759.895 2284.310 ;
        RECT 1759.565 2284.295 1759.895 2284.300 ;
        RECT 1773.365 2284.295 1773.695 2284.310 ;
        RECT 1776.790 2284.300 1777.170 2284.310 ;
        RECT 1780.265 2284.610 1780.595 2284.625 ;
        RECT 1783.230 2284.610 1783.610 2284.620 ;
        RECT 1780.265 2284.310 1783.610 2284.610 ;
        RECT 1780.265 2284.295 1780.595 2284.310 ;
        RECT 1783.230 2284.300 1783.610 2284.310 ;
        RECT 1787.165 2284.610 1787.495 2284.625 ;
        RECT 1794.065 2284.620 1794.395 2284.625 ;
        RECT 1788.750 2284.610 1789.130 2284.620 ;
        RECT 1794.065 2284.610 1794.650 2284.620 ;
        RECT 1787.165 2284.310 1789.130 2284.610 ;
        RECT 1793.840 2284.310 1794.650 2284.610 ;
        RECT 1787.165 2284.295 1787.495 2284.310 ;
        RECT 1788.750 2284.300 1789.130 2284.310 ;
        RECT 1794.065 2284.300 1794.650 2284.310 ;
        RECT 2228.765 2284.610 2229.095 2284.625 ;
        RECT 2234.030 2284.610 2234.410 2284.620 ;
        RECT 2228.765 2284.310 2234.410 2284.610 ;
        RECT 1794.065 2284.295 1794.395 2284.300 ;
        RECT 2228.765 2284.295 2229.095 2284.310 ;
        RECT 2234.030 2284.300 2234.410 2284.310 ;
        RECT 2238.885 2284.610 2239.215 2284.625 ;
        RECT 2242.310 2284.610 2242.690 2284.620 ;
        RECT 2238.885 2284.310 2242.690 2284.610 ;
        RECT 2238.885 2284.295 2239.215 2284.310 ;
        RECT 2242.310 2284.300 2242.690 2284.310 ;
        RECT 2245.785 2284.610 2246.115 2284.625 ;
        RECT 2263.725 2284.620 2264.055 2284.625 ;
        RECT 2251.510 2284.610 2251.890 2284.620 ;
        RECT 2245.785 2284.310 2251.890 2284.610 ;
        RECT 2245.785 2284.295 2246.115 2284.310 ;
        RECT 2251.510 2284.300 2251.890 2284.310 ;
        RECT 2263.470 2284.610 2264.055 2284.620 ;
        RECT 2265.310 2284.610 2265.690 2284.620 ;
        RECT 2266.485 2284.610 2266.815 2284.625 ;
        RECT 2263.470 2284.310 2264.280 2284.610 ;
        RECT 2265.310 2284.310 2266.815 2284.610 ;
        RECT 2263.470 2284.300 2264.055 2284.310 ;
        RECT 2265.310 2284.300 2265.690 2284.310 ;
        RECT 2263.725 2284.295 2264.055 2284.300 ;
        RECT 2266.485 2284.295 2266.815 2284.310 ;
        RECT 2267.405 2284.610 2267.735 2284.625 ;
        RECT 2268.070 2284.610 2268.450 2284.620 ;
        RECT 2267.405 2284.310 2268.450 2284.610 ;
        RECT 2267.405 2284.295 2267.735 2284.310 ;
        RECT 2268.070 2284.300 2268.450 2284.310 ;
        RECT 2277.065 2284.610 2277.395 2284.625 ;
        RECT 2280.950 2284.610 2281.330 2284.620 ;
        RECT 2277.065 2284.310 2281.330 2284.610 ;
        RECT 2277.065 2284.295 2277.395 2284.310 ;
        RECT 2280.950 2284.300 2281.330 2284.310 ;
        RECT 2286.470 2284.610 2286.850 2284.620 ;
        RECT 2287.185 2284.610 2287.515 2284.625 ;
        RECT 2290.405 2284.610 2290.735 2284.625 ;
        RECT 2286.470 2284.310 2290.735 2284.610 ;
        RECT 2286.470 2284.300 2286.850 2284.310 ;
        RECT 2287.185 2284.295 2287.515 2284.310 ;
        RECT 2290.405 2284.295 2290.735 2284.310 ;
        RECT 2304.665 2284.620 2304.995 2284.625 ;
        RECT 2304.665 2284.610 2305.250 2284.620 ;
        RECT 2311.565 2284.610 2311.895 2284.625 ;
        RECT 2315.910 2284.610 2316.290 2284.620 ;
        RECT 2304.665 2284.310 2305.450 2284.610 ;
        RECT 2311.565 2284.310 2316.290 2284.610 ;
        RECT 2304.665 2284.300 2305.250 2284.310 ;
        RECT 2304.665 2284.295 2304.995 2284.300 ;
        RECT 2311.565 2284.295 2311.895 2284.310 ;
        RECT 2315.910 2284.300 2316.290 2284.310 ;
        RECT 2318.465 2284.610 2318.795 2284.625 ;
        RECT 2322.350 2284.610 2322.730 2284.620 ;
        RECT 2318.465 2284.310 2322.730 2284.610 ;
        RECT 2318.465 2284.295 2318.795 2284.310 ;
        RECT 2322.350 2284.300 2322.730 2284.310 ;
        RECT 2325.365 2284.610 2325.695 2284.625 ;
        RECT 2327.870 2284.610 2328.250 2284.620 ;
        RECT 2325.365 2284.310 2328.250 2284.610 ;
        RECT 2325.365 2284.295 2325.695 2284.310 ;
        RECT 2327.870 2284.300 2328.250 2284.310 ;
        RECT 2332.265 2284.610 2332.595 2284.625 ;
        RECT 2333.390 2284.610 2333.770 2284.620 ;
        RECT 2332.265 2284.310 2333.770 2284.610 ;
        RECT 2332.265 2284.295 2332.595 2284.310 ;
        RECT 2333.390 2284.300 2333.770 2284.310 ;
        RECT 2339.165 2284.610 2339.495 2284.625 ;
        RECT 2339.830 2284.610 2340.210 2284.620 ;
        RECT 2339.165 2284.310 2340.210 2284.610 ;
        RECT 2339.165 2284.295 2339.495 2284.310 ;
        RECT 2339.830 2284.300 2340.210 2284.310 ;
        RECT 2346.065 2284.610 2346.395 2284.625 ;
        RECT 2350.870 2284.610 2351.250 2284.620 ;
        RECT 2346.065 2284.310 2351.250 2284.610 ;
        RECT 2346.065 2284.295 2346.395 2284.310 ;
        RECT 2350.870 2284.300 2351.250 2284.310 ;
        RECT 2352.965 2284.610 2353.295 2284.625 ;
        RECT 2357.310 2284.610 2357.690 2284.620 ;
        RECT 2352.965 2284.310 2357.690 2284.610 ;
        RECT 2352.965 2284.295 2353.295 2284.310 ;
        RECT 2357.310 2284.300 2357.690 2284.310 ;
        RECT 2366.765 2284.610 2367.095 2284.625 ;
        RECT 2368.350 2284.610 2368.730 2284.620 ;
        RECT 2366.765 2284.310 2368.730 2284.610 ;
        RECT 2366.765 2284.295 2367.095 2284.310 ;
        RECT 2368.350 2284.300 2368.730 2284.310 ;
        RECT 2373.665 2284.610 2373.995 2284.625 ;
        RECT 2374.790 2284.610 2375.170 2284.620 ;
        RECT 2373.665 2284.310 2375.170 2284.610 ;
        RECT 2373.665 2284.295 2373.995 2284.310 ;
        RECT 2374.790 2284.300 2375.170 2284.310 ;
        RECT 1638.585 2270.330 1638.915 2270.345 ;
        RECT 1639.505 2270.330 1639.835 2270.345 ;
        RECT 1638.585 2270.030 1639.835 2270.330 ;
        RECT 1638.585 2270.015 1638.915 2270.030 ;
        RECT 1639.505 2270.015 1639.835 2270.030 ;
        RECT 284.345 2212.530 284.675 2212.545 ;
        RECT 814.725 2212.530 815.055 2212.545 ;
        RECT 284.345 2212.230 815.055 2212.530 ;
        RECT 284.345 2212.215 284.675 2212.230 ;
        RECT 814.725 2212.215 815.055 2212.230 ;
        RECT 1165.705 2212.530 1166.035 2212.545 ;
        RECT 1437.565 2212.530 1437.895 2212.545 ;
        RECT 1165.705 2212.230 1437.895 2212.530 ;
        RECT 1165.705 2212.215 1166.035 2212.230 ;
        RECT 1437.565 2212.215 1437.895 2212.230 ;
        RECT 287.105 2211.850 287.435 2211.865 ;
        RECT 826.225 2211.850 826.555 2211.865 ;
        RECT 287.105 2211.550 826.555 2211.850 ;
        RECT 287.105 2211.535 287.435 2211.550 ;
        RECT 826.225 2211.535 826.555 2211.550 ;
        RECT 1172.605 2211.850 1172.935 2211.865 ;
        RECT 1448.605 2211.850 1448.935 2211.865 ;
        RECT 1172.605 2211.550 1448.935 2211.850 ;
        RECT 1172.605 2211.535 1172.935 2211.550 ;
        RECT 1448.605 2211.535 1448.935 2211.550 ;
        RECT 287.565 2211.170 287.895 2211.185 ;
        RECT 837.265 2211.170 837.595 2211.185 ;
        RECT 287.565 2210.870 837.595 2211.170 ;
        RECT 287.565 2210.855 287.895 2210.870 ;
        RECT 837.265 2210.855 837.595 2210.870 ;
        RECT 1186.405 2211.170 1186.735 2211.185 ;
        RECT 1471.605 2211.170 1471.935 2211.185 ;
        RECT 1186.405 2210.870 1471.935 2211.170 ;
        RECT 1186.405 2210.855 1186.735 2210.870 ;
        RECT 1471.605 2210.855 1471.935 2210.870 ;
        RECT 1200.205 2208.450 1200.535 2208.465 ;
        RECT 1243.445 2208.450 1243.775 2208.465 ;
        RECT 1200.205 2208.150 1243.775 2208.450 ;
        RECT 1200.205 2208.135 1200.535 2208.150 ;
        RECT 1243.445 2208.135 1243.775 2208.150 ;
        RECT 1514.845 2194.850 1515.175 2194.865 ;
        RECT 1499.140 2194.720 1515.175 2194.850 ;
      LAYER met3 ;
        RECT 304.400 2193.720 1495.600 2194.585 ;
      LAYER met3 ;
        RECT 1496.000 2194.550 1515.175 2194.720 ;
        RECT 1496.000 2194.120 1500.000 2194.550 ;
        RECT 1514.845 2194.535 1515.175 2194.550 ;
      LAYER met3 ;
        RECT 304.000 2184.920 1496.000 2193.720 ;
        RECT 304.400 2184.240 1496.000 2184.920 ;
        RECT 304.400 2183.520 1495.600 2184.240 ;
      LAYER met3 ;
        RECT 1513.925 2183.970 1514.255 2183.985 ;
        RECT 1499.140 2183.840 1514.255 2183.970 ;
      LAYER met3 ;
        RECT 304.000 2182.840 1495.600 2183.520 ;
      LAYER met3 ;
        RECT 1496.000 2183.670 1514.255 2183.840 ;
        RECT 1496.000 2183.240 1500.000 2183.670 ;
        RECT 1513.925 2183.655 1514.255 2183.670 ;
      LAYER met3 ;
        RECT 304.000 2174.040 1496.000 2182.840 ;
        RECT 304.400 2173.360 1496.000 2174.040 ;
        RECT 304.400 2172.640 1495.600 2173.360 ;
      LAYER met3 ;
        RECT 1513.925 2173.090 1514.255 2173.105 ;
        RECT 1499.140 2172.960 1514.255 2173.090 ;
      LAYER met3 ;
        RECT 304.000 2171.960 1495.600 2172.640 ;
      LAYER met3 ;
        RECT 1496.000 2172.790 1514.255 2172.960 ;
        RECT 1496.000 2172.360 1500.000 2172.790 ;
        RECT 1513.925 2172.775 1514.255 2172.790 ;
      LAYER met3 ;
        RECT 304.000 2163.840 1496.000 2171.960 ;
        RECT 304.400 2162.480 1496.000 2163.840 ;
        RECT 304.400 2162.440 1495.600 2162.480 ;
        RECT 304.000 2161.080 1495.600 2162.440 ;
      LAYER met3 ;
        RECT 1513.925 2162.210 1514.255 2162.225 ;
        RECT 1499.140 2162.080 1514.255 2162.210 ;
        RECT 1496.000 2161.910 1514.255 2162.080 ;
        RECT 1496.000 2161.480 1500.000 2161.910 ;
        RECT 1513.925 2161.895 1514.255 2161.910 ;
      LAYER met3 ;
        RECT 304.000 2152.960 1496.000 2161.080 ;
        RECT 304.400 2151.600 1496.000 2152.960 ;
        RECT 304.400 2151.560 1495.600 2151.600 ;
        RECT 304.000 2150.200 1495.600 2151.560 ;
      LAYER met3 ;
        RECT 1513.925 2151.330 1514.255 2151.345 ;
        RECT 1499.140 2151.200 1514.255 2151.330 ;
        RECT 1496.000 2151.030 1514.255 2151.200 ;
        RECT 1496.000 2150.600 1500.000 2151.030 ;
        RECT 1513.925 2151.015 1514.255 2151.030 ;
      LAYER met3 ;
        RECT 304.000 2142.760 1496.000 2150.200 ;
        RECT 304.400 2141.360 1496.000 2142.760 ;
        RECT 304.000 2140.040 1496.000 2141.360 ;
        RECT 304.000 2138.640 1495.600 2140.040 ;
      LAYER met3 ;
        RECT 1513.925 2139.770 1514.255 2139.785 ;
        RECT 1499.140 2139.640 1514.255 2139.770 ;
        RECT 1496.000 2139.470 1514.255 2139.640 ;
        RECT 1496.000 2139.040 1500.000 2139.470 ;
        RECT 1513.925 2139.455 1514.255 2139.470 ;
      LAYER met3 ;
        RECT 304.000 2131.880 1496.000 2138.640 ;
        RECT 304.400 2130.480 1496.000 2131.880 ;
        RECT 304.000 2129.160 1496.000 2130.480 ;
        RECT 304.000 2127.760 1495.600 2129.160 ;
      LAYER met3 ;
        RECT 1513.925 2128.890 1514.255 2128.905 ;
        RECT 1499.140 2128.760 1514.255 2128.890 ;
        RECT 1496.000 2128.590 1514.255 2128.760 ;
        RECT 1496.000 2128.160 1500.000 2128.590 ;
        RECT 1513.925 2128.575 1514.255 2128.590 ;
      LAYER met3 ;
        RECT 304.000 2121.680 1496.000 2127.760 ;
        RECT 304.400 2120.280 1496.000 2121.680 ;
        RECT 304.000 2118.280 1496.000 2120.280 ;
        RECT 304.000 2116.880 1495.600 2118.280 ;
      LAYER met3 ;
        RECT 1513.925 2118.010 1514.255 2118.025 ;
        RECT 1499.140 2117.880 1514.255 2118.010 ;
        RECT 1496.000 2117.710 1514.255 2117.880 ;
        RECT 1496.000 2117.280 1500.000 2117.710 ;
        RECT 1513.925 2117.695 1514.255 2117.710 ;
      LAYER met3 ;
        RECT 304.000 2110.800 1496.000 2116.880 ;
        RECT 304.400 2109.400 1496.000 2110.800 ;
        RECT 304.000 2107.400 1496.000 2109.400 ;
        RECT 304.000 2106.000 1495.600 2107.400 ;
      LAYER met3 ;
        RECT 1513.925 2107.130 1514.255 2107.145 ;
        RECT 1499.140 2107.000 1514.255 2107.130 ;
        RECT 1496.000 2106.830 1514.255 2107.000 ;
        RECT 1496.000 2106.400 1500.000 2106.830 ;
        RECT 1513.925 2106.815 1514.255 2106.830 ;
      LAYER met3 ;
        RECT 304.000 2100.600 1496.000 2106.000 ;
        RECT 304.400 2099.200 1496.000 2100.600 ;
        RECT 304.000 2096.520 1496.000 2099.200 ;
        RECT 304.000 2095.120 1495.600 2096.520 ;
      LAYER met3 ;
        RECT 1513.925 2096.250 1514.255 2096.265 ;
        RECT 1499.140 2096.120 1514.255 2096.250 ;
        RECT 1496.000 2095.950 1514.255 2096.120 ;
        RECT 1496.000 2095.520 1500.000 2095.950 ;
        RECT 1513.925 2095.935 1514.255 2095.950 ;
      LAYER met3 ;
        RECT 304.000 2089.720 1496.000 2095.120 ;
        RECT 304.400 2088.320 1496.000 2089.720 ;
        RECT 304.000 2084.960 1496.000 2088.320 ;
        RECT 304.000 2083.560 1495.600 2084.960 ;
      LAYER met3 ;
        RECT 1513.925 2084.690 1514.255 2084.705 ;
        RECT 1499.140 2084.560 1514.255 2084.690 ;
        RECT 1496.000 2084.390 1514.255 2084.560 ;
        RECT 1496.000 2083.960 1500.000 2084.390 ;
        RECT 1513.925 2084.375 1514.255 2084.390 ;
      LAYER met3 ;
        RECT 304.000 2079.520 1496.000 2083.560 ;
        RECT 304.400 2078.120 1496.000 2079.520 ;
        RECT 304.000 2074.080 1496.000 2078.120 ;
        RECT 304.000 2072.680 1495.600 2074.080 ;
      LAYER met3 ;
        RECT 1513.925 2073.810 1514.255 2073.825 ;
        RECT 1499.140 2073.680 1514.255 2073.810 ;
        RECT 1496.000 2073.510 1514.255 2073.680 ;
        RECT 1496.000 2073.080 1500.000 2073.510 ;
        RECT 1513.925 2073.495 1514.255 2073.510 ;
      LAYER met3 ;
        RECT 304.000 2068.640 1496.000 2072.680 ;
        RECT 304.400 2067.240 1496.000 2068.640 ;
        RECT 304.000 2063.200 1496.000 2067.240 ;
        RECT 304.000 2061.800 1495.600 2063.200 ;
      LAYER met3 ;
        RECT 1513.925 2062.930 1514.255 2062.945 ;
        RECT 1499.140 2062.800 1514.255 2062.930 ;
        RECT 1496.000 2062.630 1514.255 2062.800 ;
        RECT 1496.000 2062.200 1500.000 2062.630 ;
        RECT 1513.925 2062.615 1514.255 2062.630 ;
      LAYER met3 ;
        RECT 304.000 2058.440 1496.000 2061.800 ;
        RECT 304.400 2057.040 1496.000 2058.440 ;
        RECT 304.000 2052.320 1496.000 2057.040 ;
        RECT 304.000 2050.920 1495.600 2052.320 ;
      LAYER met3 ;
        RECT 1513.925 2052.050 1514.255 2052.065 ;
        RECT 1499.140 2051.920 1514.255 2052.050 ;
        RECT 1496.000 2051.750 1514.255 2051.920 ;
        RECT 1496.000 2051.320 1500.000 2051.750 ;
        RECT 1513.925 2051.735 1514.255 2051.750 ;
      LAYER met3 ;
        RECT 304.000 2047.560 1496.000 2050.920 ;
        RECT 304.400 2046.160 1496.000 2047.560 ;
        RECT 304.000 2041.440 1496.000 2046.160 ;
        RECT 304.000 2040.040 1495.600 2041.440 ;
      LAYER met3 ;
        RECT 1513.925 2041.170 1514.255 2041.185 ;
        RECT 1499.140 2041.040 1514.255 2041.170 ;
        RECT 1496.000 2040.870 1514.255 2041.040 ;
        RECT 1496.000 2040.440 1500.000 2040.870 ;
        RECT 1513.925 2040.855 1514.255 2040.870 ;
      LAYER met3 ;
        RECT 304.000 2037.360 1496.000 2040.040 ;
        RECT 304.400 2035.960 1496.000 2037.360 ;
        RECT 304.000 2029.880 1496.000 2035.960 ;
        RECT 304.000 2028.480 1495.600 2029.880 ;
      LAYER met3 ;
        RECT 1513.925 2029.610 1514.255 2029.625 ;
        RECT 1499.140 2029.480 1514.255 2029.610 ;
        RECT 1496.000 2029.310 1514.255 2029.480 ;
        RECT 1496.000 2028.880 1500.000 2029.310 ;
        RECT 1513.925 2029.295 1514.255 2029.310 ;
      LAYER met3 ;
        RECT 304.000 2026.480 1496.000 2028.480 ;
        RECT 304.400 2025.080 1496.000 2026.480 ;
        RECT 304.000 2019.000 1496.000 2025.080 ;
        RECT 304.000 2017.600 1495.600 2019.000 ;
      LAYER met3 ;
        RECT 1513.465 2018.730 1513.795 2018.745 ;
        RECT 1499.140 2018.600 1513.795 2018.730 ;
        RECT 1496.000 2018.430 1513.795 2018.600 ;
        RECT 1496.000 2018.000 1500.000 2018.430 ;
        RECT 1513.465 2018.415 1513.795 2018.430 ;
      LAYER met3 ;
        RECT 304.000 2016.280 1496.000 2017.600 ;
        RECT 304.400 2014.880 1496.000 2016.280 ;
        RECT 304.000 2008.120 1496.000 2014.880 ;
        RECT 304.000 2006.720 1495.600 2008.120 ;
      LAYER met3 ;
        RECT 1513.925 2007.850 1514.255 2007.865 ;
        RECT 1499.140 2007.720 1514.255 2007.850 ;
        RECT 1496.000 2007.550 1514.255 2007.720 ;
        RECT 1496.000 2007.120 1500.000 2007.550 ;
        RECT 1513.925 2007.535 1514.255 2007.550 ;
      LAYER met3 ;
        RECT 304.000 2005.400 1496.000 2006.720 ;
        RECT 304.400 2004.000 1496.000 2005.400 ;
        RECT 304.000 1997.240 1496.000 2004.000 ;
        RECT 304.000 1995.840 1495.600 1997.240 ;
      LAYER met3 ;
        RECT 1513.925 1996.970 1514.255 1996.985 ;
        RECT 1499.140 1996.840 1514.255 1996.970 ;
        RECT 1496.000 1996.670 1514.255 1996.840 ;
        RECT 1496.000 1996.240 1500.000 1996.670 ;
        RECT 1513.925 1996.655 1514.255 1996.670 ;
      LAYER met3 ;
        RECT 304.000 1995.200 1496.000 1995.840 ;
        RECT 304.400 1993.800 1496.000 1995.200 ;
        RECT 304.000 1986.360 1496.000 1993.800 ;
        RECT 304.000 1984.960 1495.600 1986.360 ;
      LAYER met3 ;
        RECT 1513.925 1986.090 1514.255 1986.105 ;
        RECT 1499.140 1985.960 1514.255 1986.090 ;
        RECT 1496.000 1985.790 1514.255 1985.960 ;
        RECT 1496.000 1985.360 1500.000 1985.790 ;
        RECT 1513.925 1985.775 1514.255 1985.790 ;
      LAYER met3 ;
        RECT 304.000 1984.320 1496.000 1984.960 ;
        RECT 304.400 1982.920 1496.000 1984.320 ;
        RECT 304.000 1974.800 1496.000 1982.920 ;
        RECT 304.000 1974.120 1495.600 1974.800 ;
      LAYER met3 ;
        RECT 1512.545 1974.530 1512.875 1974.545 ;
        RECT 1499.140 1974.400 1512.875 1974.530 ;
      LAYER met3 ;
        RECT 304.400 1973.400 1495.600 1974.120 ;
      LAYER met3 ;
        RECT 1496.000 1974.230 1512.875 1974.400 ;
        RECT 1496.000 1973.800 1500.000 1974.230 ;
        RECT 1512.545 1974.215 1512.875 1974.230 ;
      LAYER met3 ;
        RECT 304.400 1972.720 1496.000 1973.400 ;
        RECT 304.000 1963.920 1496.000 1972.720 ;
        RECT 304.000 1963.240 1495.600 1963.920 ;
      LAYER met3 ;
        RECT 1513.465 1963.650 1513.795 1963.665 ;
        RECT 1499.140 1963.520 1513.795 1963.650 ;
      LAYER met3 ;
        RECT 304.400 1962.520 1495.600 1963.240 ;
      LAYER met3 ;
        RECT 1496.000 1963.350 1513.795 1963.520 ;
        RECT 1496.000 1962.920 1500.000 1963.350 ;
        RECT 1513.465 1963.335 1513.795 1963.350 ;
      LAYER met3 ;
        RECT 304.400 1961.840 1496.000 1962.520 ;
        RECT 304.000 1953.040 1496.000 1961.840 ;
        RECT 304.400 1951.640 1495.600 1953.040 ;
      LAYER met3 ;
        RECT 1513.925 1952.770 1514.255 1952.785 ;
        RECT 1499.140 1952.640 1514.255 1952.770 ;
        RECT 1496.000 1952.470 1514.255 1952.640 ;
        RECT 1496.000 1952.040 1500.000 1952.470 ;
        RECT 1513.925 1952.455 1514.255 1952.470 ;
      LAYER met3 ;
        RECT 304.000 1942.160 1496.000 1951.640 ;
        RECT 304.400 1940.760 1495.600 1942.160 ;
      LAYER met3 ;
        RECT 1513.925 1941.890 1514.255 1941.905 ;
        RECT 1499.140 1941.760 1514.255 1941.890 ;
        RECT 1496.000 1941.590 1514.255 1941.760 ;
        RECT 1496.000 1941.160 1500.000 1941.590 ;
        RECT 1513.925 1941.575 1514.255 1941.590 ;
      LAYER met3 ;
        RECT 304.000 1931.960 1496.000 1940.760 ;
        RECT 304.400 1931.280 1496.000 1931.960 ;
        RECT 304.400 1930.560 1495.600 1931.280 ;
      LAYER met3 ;
        RECT 1512.545 1931.010 1512.875 1931.025 ;
        RECT 1499.140 1930.880 1512.875 1931.010 ;
      LAYER met3 ;
        RECT 304.000 1929.880 1495.600 1930.560 ;
      LAYER met3 ;
        RECT 1496.000 1930.710 1512.875 1930.880 ;
        RECT 1496.000 1930.280 1500.000 1930.710 ;
        RECT 1512.545 1930.695 1512.875 1930.710 ;
      LAYER met3 ;
        RECT 304.000 1921.080 1496.000 1929.880 ;
        RECT 304.400 1919.720 1496.000 1921.080 ;
        RECT 304.400 1919.680 1495.600 1919.720 ;
        RECT 304.000 1918.320 1495.600 1919.680 ;
      LAYER met3 ;
        RECT 1512.545 1919.450 1512.875 1919.465 ;
        RECT 1499.140 1919.320 1512.875 1919.450 ;
        RECT 1496.000 1919.150 1512.875 1919.320 ;
        RECT 1496.000 1918.720 1500.000 1919.150 ;
        RECT 1512.545 1919.135 1512.875 1919.150 ;
      LAYER met3 ;
        RECT 304.000 1910.880 1496.000 1918.320 ;
        RECT 304.400 1909.480 1496.000 1910.880 ;
        RECT 304.000 1908.840 1496.000 1909.480 ;
        RECT 304.000 1907.440 1495.600 1908.840 ;
      LAYER met3 ;
        RECT 1513.925 1908.570 1514.255 1908.585 ;
        RECT 1499.140 1908.440 1514.255 1908.570 ;
        RECT 1496.000 1908.270 1514.255 1908.440 ;
        RECT 1496.000 1907.840 1500.000 1908.270 ;
        RECT 1513.925 1908.255 1514.255 1908.270 ;
      LAYER met3 ;
        RECT 304.000 1900.680 1496.000 1907.440 ;
        RECT 304.400 1899.280 1496.000 1900.680 ;
        RECT 304.000 1897.960 1496.000 1899.280 ;
        RECT 304.000 1896.560 1495.600 1897.960 ;
      LAYER met3 ;
        RECT 1513.005 1897.690 1513.335 1897.705 ;
        RECT 1499.140 1897.560 1513.335 1897.690 ;
        RECT 1496.000 1897.390 1513.335 1897.560 ;
        RECT 1496.000 1896.960 1500.000 1897.390 ;
        RECT 1513.005 1897.375 1513.335 1897.390 ;
      LAYER met3 ;
        RECT 304.000 1889.800 1496.000 1896.560 ;
        RECT 304.400 1888.400 1496.000 1889.800 ;
        RECT 304.000 1887.080 1496.000 1888.400 ;
        RECT 304.000 1885.680 1495.600 1887.080 ;
      LAYER met3 ;
        RECT 1513.925 1886.810 1514.255 1886.825 ;
        RECT 1499.140 1886.680 1514.255 1886.810 ;
        RECT 1496.000 1886.510 1514.255 1886.680 ;
        RECT 1496.000 1886.080 1500.000 1886.510 ;
        RECT 1513.925 1886.495 1514.255 1886.510 ;
      LAYER met3 ;
        RECT 304.000 1879.600 1496.000 1885.680 ;
        RECT 304.400 1878.200 1496.000 1879.600 ;
        RECT 304.000 1876.200 1496.000 1878.200 ;
        RECT 304.000 1874.800 1495.600 1876.200 ;
      LAYER met3 ;
        RECT 1513.925 1875.930 1514.255 1875.945 ;
        RECT 1499.140 1875.800 1514.255 1875.930 ;
        RECT 1496.000 1875.630 1514.255 1875.800 ;
        RECT 1496.000 1875.200 1500.000 1875.630 ;
        RECT 1513.925 1875.615 1514.255 1875.630 ;
      LAYER met3 ;
        RECT 304.000 1868.720 1496.000 1874.800 ;
        RECT 304.400 1867.320 1496.000 1868.720 ;
        RECT 304.000 1865.320 1496.000 1867.320 ;
        RECT 304.000 1863.920 1495.600 1865.320 ;
      LAYER met3 ;
        RECT 1513.925 1865.050 1514.255 1865.065 ;
        RECT 1499.140 1864.920 1514.255 1865.050 ;
        RECT 1496.000 1864.750 1514.255 1864.920 ;
        RECT 1496.000 1864.320 1500.000 1864.750 ;
        RECT 1513.925 1864.735 1514.255 1864.750 ;
      LAYER met3 ;
        RECT 304.000 1858.520 1496.000 1863.920 ;
        RECT 304.400 1857.120 1496.000 1858.520 ;
        RECT 304.000 1853.760 1496.000 1857.120 ;
        RECT 304.000 1852.360 1495.600 1853.760 ;
      LAYER met3 ;
        RECT 1511.625 1853.490 1511.955 1853.505 ;
        RECT 1499.140 1853.360 1511.955 1853.490 ;
        RECT 1496.000 1853.190 1511.955 1853.360 ;
        RECT 1496.000 1852.760 1500.000 1853.190 ;
        RECT 1511.625 1853.175 1511.955 1853.190 ;
      LAYER met3 ;
        RECT 304.000 1847.640 1496.000 1852.360 ;
        RECT 304.400 1846.240 1496.000 1847.640 ;
        RECT 304.000 1842.880 1496.000 1846.240 ;
        RECT 304.000 1841.480 1495.600 1842.880 ;
      LAYER met3 ;
        RECT 1513.005 1842.610 1513.335 1842.625 ;
        RECT 1499.140 1842.480 1513.335 1842.610 ;
        RECT 1496.000 1842.310 1513.335 1842.480 ;
        RECT 1496.000 1841.880 1500.000 1842.310 ;
        RECT 1513.005 1842.295 1513.335 1842.310 ;
      LAYER met3 ;
        RECT 304.000 1837.440 1496.000 1841.480 ;
        RECT 304.400 1836.040 1496.000 1837.440 ;
        RECT 304.000 1832.000 1496.000 1836.040 ;
      LAYER met3 ;
        RECT 1639.045 1835.130 1639.375 1835.145 ;
        RECT 1640.425 1835.130 1640.755 1835.145 ;
        RECT 1639.045 1834.830 1640.755 1835.130 ;
        RECT 1639.045 1834.815 1639.375 1834.830 ;
        RECT 1640.425 1834.815 1640.755 1834.830 ;
      LAYER met3 ;
        RECT 304.000 1830.600 1495.600 1832.000 ;
      LAYER met3 ;
        RECT 1513.925 1831.730 1514.255 1831.745 ;
        RECT 1499.140 1831.600 1514.255 1831.730 ;
        RECT 1496.000 1831.430 1514.255 1831.600 ;
        RECT 1496.000 1831.000 1500.000 1831.430 ;
        RECT 1513.925 1831.415 1514.255 1831.430 ;
      LAYER met3 ;
        RECT 304.000 1826.560 1496.000 1830.600 ;
        RECT 304.400 1825.160 1496.000 1826.560 ;
        RECT 304.000 1821.120 1496.000 1825.160 ;
        RECT 304.000 1819.720 1495.600 1821.120 ;
      LAYER met3 ;
        RECT 1512.545 1820.850 1512.875 1820.865 ;
        RECT 1499.140 1820.720 1512.875 1820.850 ;
        RECT 1496.000 1820.550 1512.875 1820.720 ;
        RECT 1496.000 1820.120 1500.000 1820.550 ;
        RECT 1512.545 1820.535 1512.875 1820.550 ;
      LAYER met3 ;
        RECT 304.000 1816.360 1496.000 1819.720 ;
        RECT 304.400 1814.960 1496.000 1816.360 ;
        RECT 304.000 1810.240 1496.000 1814.960 ;
        RECT 304.000 1808.840 1495.600 1810.240 ;
      LAYER met3 ;
        RECT 1512.085 1809.970 1512.415 1809.985 ;
        RECT 1499.140 1809.840 1512.415 1809.970 ;
        RECT 1496.000 1809.670 1512.415 1809.840 ;
        RECT 1496.000 1809.240 1500.000 1809.670 ;
        RECT 1512.085 1809.655 1512.415 1809.670 ;
      LAYER met3 ;
        RECT 304.000 1805.480 1496.000 1808.840 ;
        RECT 304.400 1804.080 1496.000 1805.480 ;
        RECT 304.000 1798.680 1496.000 1804.080 ;
        RECT 304.000 1797.280 1495.600 1798.680 ;
      LAYER met3 ;
        RECT 1511.625 1798.410 1511.955 1798.425 ;
        RECT 1499.140 1798.280 1511.955 1798.410 ;
        RECT 1496.000 1798.110 1511.955 1798.280 ;
        RECT 1496.000 1797.680 1500.000 1798.110 ;
        RECT 1511.625 1798.095 1511.955 1798.110 ;
      LAYER met3 ;
        RECT 304.000 1795.280 1496.000 1797.280 ;
        RECT 304.400 1793.880 1496.000 1795.280 ;
        RECT 304.000 1787.800 1496.000 1793.880 ;
        RECT 304.000 1786.400 1495.600 1787.800 ;
      LAYER met3 ;
        RECT 1512.545 1787.530 1512.875 1787.545 ;
        RECT 1499.140 1787.400 1512.875 1787.530 ;
        RECT 1496.000 1787.230 1512.875 1787.400 ;
        RECT 1496.000 1786.800 1500.000 1787.230 ;
        RECT 1512.545 1787.215 1512.875 1787.230 ;
      LAYER met3 ;
        RECT 304.000 1784.400 1496.000 1786.400 ;
        RECT 304.400 1783.000 1496.000 1784.400 ;
        RECT 304.000 1776.920 1496.000 1783.000 ;
        RECT 304.000 1775.520 1495.600 1776.920 ;
      LAYER met3 ;
        RECT 1513.925 1776.650 1514.255 1776.665 ;
        RECT 1499.140 1776.520 1514.255 1776.650 ;
        RECT 1496.000 1776.350 1514.255 1776.520 ;
        RECT 1496.000 1775.920 1500.000 1776.350 ;
        RECT 1513.925 1776.335 1514.255 1776.350 ;
      LAYER met3 ;
        RECT 304.000 1774.200 1496.000 1775.520 ;
        RECT 304.400 1772.800 1496.000 1774.200 ;
        RECT 304.000 1766.040 1496.000 1772.800 ;
        RECT 304.000 1764.640 1495.600 1766.040 ;
      LAYER met3 ;
        RECT 1513.925 1765.770 1514.255 1765.785 ;
        RECT 1499.140 1765.640 1514.255 1765.770 ;
        RECT 1496.000 1765.470 1514.255 1765.640 ;
        RECT 1496.000 1765.040 1500.000 1765.470 ;
        RECT 1513.925 1765.455 1514.255 1765.470 ;
      LAYER met3 ;
        RECT 304.000 1763.320 1496.000 1764.640 ;
        RECT 304.400 1761.920 1496.000 1763.320 ;
        RECT 304.000 1755.160 1496.000 1761.920 ;
        RECT 304.000 1753.760 1495.600 1755.160 ;
      LAYER met3 ;
        RECT 1512.085 1754.890 1512.415 1754.905 ;
        RECT 1499.140 1754.760 1512.415 1754.890 ;
        RECT 1496.000 1754.590 1512.415 1754.760 ;
        RECT 1496.000 1754.160 1500.000 1754.590 ;
        RECT 1512.085 1754.575 1512.415 1754.590 ;
      LAYER met3 ;
        RECT 304.000 1753.120 1496.000 1753.760 ;
        RECT 304.400 1751.720 1496.000 1753.120 ;
        RECT 304.000 1743.600 1496.000 1751.720 ;
        RECT 304.000 1742.240 1495.600 1743.600 ;
      LAYER met3 ;
        RECT 1513.465 1743.330 1513.795 1743.345 ;
        RECT 1499.140 1743.200 1513.795 1743.330 ;
        RECT 1496.000 1743.030 1513.795 1743.200 ;
        RECT 1496.000 1742.600 1500.000 1743.030 ;
        RECT 1513.465 1743.015 1513.795 1743.030 ;
      LAYER met3 ;
        RECT 304.400 1742.200 1495.600 1742.240 ;
        RECT 304.400 1740.840 1496.000 1742.200 ;
        RECT 304.000 1732.720 1496.000 1740.840 ;
        RECT 304.000 1732.040 1495.600 1732.720 ;
      LAYER met3 ;
        RECT 1512.545 1732.450 1512.875 1732.465 ;
        RECT 1499.140 1732.320 1512.875 1732.450 ;
      LAYER met3 ;
        RECT 304.400 1731.320 1495.600 1732.040 ;
      LAYER met3 ;
        RECT 1496.000 1732.150 1512.875 1732.320 ;
        RECT 1496.000 1731.720 1500.000 1732.150 ;
        RECT 1512.545 1732.135 1512.875 1732.150 ;
      LAYER met3 ;
        RECT 304.400 1730.640 1496.000 1731.320 ;
        RECT 304.000 1721.840 1496.000 1730.640 ;
        RECT 304.000 1721.160 1495.600 1721.840 ;
      LAYER met3 ;
        RECT 1513.925 1721.570 1514.255 1721.585 ;
        RECT 1499.140 1721.440 1514.255 1721.570 ;
      LAYER met3 ;
        RECT 304.400 1720.440 1495.600 1721.160 ;
      LAYER met3 ;
        RECT 1496.000 1721.270 1514.255 1721.440 ;
        RECT 1496.000 1720.840 1500.000 1721.270 ;
        RECT 1513.925 1721.255 1514.255 1721.270 ;
      LAYER met3 ;
        RECT 304.400 1719.760 1496.000 1720.440 ;
        RECT 304.000 1710.960 1496.000 1719.760 ;
        RECT 304.400 1709.560 1495.600 1710.960 ;
      LAYER met3 ;
        RECT 1513.925 1710.690 1514.255 1710.705 ;
        RECT 1499.140 1710.560 1514.255 1710.690 ;
        RECT 1496.000 1710.390 1514.255 1710.560 ;
        RECT 1496.000 1709.960 1500.000 1710.390 ;
        RECT 1513.925 1710.375 1514.255 1710.390 ;
      LAYER met3 ;
        RECT 304.000 1700.080 1496.000 1709.560 ;
        RECT 304.400 1698.680 1495.600 1700.080 ;
      LAYER met3 ;
        RECT 1512.085 1699.810 1512.415 1699.825 ;
        RECT 1499.140 1699.680 1512.415 1699.810 ;
        RECT 1496.000 1699.510 1512.415 1699.680 ;
        RECT 1496.000 1699.080 1500.000 1699.510 ;
        RECT 1512.085 1699.495 1512.415 1699.510 ;
      LAYER met3 ;
        RECT 304.000 1689.880 1496.000 1698.680 ;
        RECT 304.400 1688.520 1496.000 1689.880 ;
        RECT 304.400 1688.480 1495.600 1688.520 ;
        RECT 304.000 1687.120 1495.600 1688.480 ;
      LAYER met3 ;
        RECT 1513.465 1688.250 1513.795 1688.265 ;
        RECT 1499.140 1688.120 1513.795 1688.250 ;
        RECT 1496.000 1687.950 1513.795 1688.120 ;
        RECT 1496.000 1687.520 1500.000 1687.950 ;
        RECT 1513.465 1687.935 1513.795 1687.950 ;
      LAYER met3 ;
        RECT 304.000 1679.000 1496.000 1687.120 ;
        RECT 304.400 1677.640 1496.000 1679.000 ;
        RECT 304.400 1677.600 1495.600 1677.640 ;
        RECT 304.000 1676.240 1495.600 1677.600 ;
      LAYER met3 ;
        RECT 1512.545 1677.370 1512.875 1677.385 ;
        RECT 1499.140 1677.240 1512.875 1677.370 ;
        RECT 1496.000 1677.070 1512.875 1677.240 ;
        RECT 1496.000 1676.640 1500.000 1677.070 ;
        RECT 1512.545 1677.055 1512.875 1677.070 ;
      LAYER met3 ;
        RECT 304.000 1668.800 1496.000 1676.240 ;
        RECT 304.400 1667.400 1496.000 1668.800 ;
        RECT 304.000 1666.760 1496.000 1667.400 ;
        RECT 304.000 1665.360 1495.600 1666.760 ;
      LAYER met3 ;
        RECT 1513.925 1666.490 1514.255 1666.505 ;
        RECT 1499.140 1666.360 1514.255 1666.490 ;
        RECT 1496.000 1666.190 1514.255 1666.360 ;
        RECT 1496.000 1665.760 1500.000 1666.190 ;
        RECT 1513.925 1666.175 1514.255 1666.190 ;
      LAYER met3 ;
        RECT 304.000 1657.920 1496.000 1665.360 ;
        RECT 304.400 1656.520 1496.000 1657.920 ;
        RECT 304.000 1655.880 1496.000 1656.520 ;
        RECT 304.000 1654.480 1495.600 1655.880 ;
      LAYER met3 ;
        RECT 1512.545 1655.610 1512.875 1655.625 ;
        RECT 1499.140 1655.480 1512.875 1655.610 ;
        RECT 1496.000 1655.310 1512.875 1655.480 ;
        RECT 1496.000 1654.880 1500.000 1655.310 ;
        RECT 1512.545 1655.295 1512.875 1655.310 ;
      LAYER met3 ;
        RECT 304.000 1647.720 1496.000 1654.480 ;
        RECT 304.400 1646.320 1496.000 1647.720 ;
        RECT 304.000 1645.000 1496.000 1646.320 ;
        RECT 304.000 1643.600 1495.600 1645.000 ;
      LAYER met3 ;
        RECT 1511.625 1644.730 1511.955 1644.745 ;
        RECT 1499.140 1644.600 1511.955 1644.730 ;
        RECT 1496.000 1644.430 1511.955 1644.600 ;
        RECT 1496.000 1644.000 1500.000 1644.430 ;
        RECT 1511.625 1644.415 1511.955 1644.430 ;
      LAYER met3 ;
        RECT 304.000 1636.840 1496.000 1643.600 ;
        RECT 304.400 1635.440 1496.000 1636.840 ;
        RECT 304.000 1633.440 1496.000 1635.440 ;
        RECT 304.000 1632.040 1495.600 1633.440 ;
      LAYER met3 ;
        RECT 1512.545 1633.170 1512.875 1633.185 ;
        RECT 1499.140 1633.040 1512.875 1633.170 ;
        RECT 1496.000 1632.870 1512.875 1633.040 ;
        RECT 1496.000 1632.440 1500.000 1632.870 ;
        RECT 1512.545 1632.855 1512.875 1632.870 ;
      LAYER met3 ;
        RECT 304.000 1626.640 1496.000 1632.040 ;
        RECT 304.400 1625.240 1496.000 1626.640 ;
        RECT 304.000 1622.560 1496.000 1625.240 ;
        RECT 304.000 1621.160 1495.600 1622.560 ;
      LAYER met3 ;
        RECT 1511.625 1622.290 1511.955 1622.305 ;
        RECT 1499.140 1622.160 1511.955 1622.290 ;
        RECT 1496.000 1621.990 1511.955 1622.160 ;
        RECT 1496.000 1621.560 1500.000 1621.990 ;
        RECT 1511.625 1621.975 1511.955 1621.990 ;
      LAYER met3 ;
        RECT 304.000 1615.760 1496.000 1621.160 ;
        RECT 304.400 1614.360 1496.000 1615.760 ;
        RECT 304.000 1611.680 1496.000 1614.360 ;
        RECT 304.000 1610.280 1495.600 1611.680 ;
      LAYER met3 ;
        RECT 1511.625 1611.410 1511.955 1611.425 ;
        RECT 1499.140 1611.280 1511.955 1611.410 ;
        RECT 1496.000 1611.110 1511.955 1611.280 ;
        RECT 1496.000 1610.680 1500.000 1611.110 ;
        RECT 1511.625 1611.095 1511.955 1611.110 ;
      LAYER met3 ;
        RECT 304.000 1605.560 1496.000 1610.280 ;
        RECT 304.400 1604.160 1496.000 1605.560 ;
        RECT 304.000 1600.800 1496.000 1604.160 ;
        RECT 304.000 1599.400 1495.600 1600.800 ;
      LAYER met3 ;
        RECT 1511.625 1600.530 1511.955 1600.545 ;
        RECT 1499.140 1600.400 1511.955 1600.530 ;
        RECT 1496.000 1600.230 1511.955 1600.400 ;
        RECT 1496.000 1599.800 1500.000 1600.230 ;
        RECT 1511.625 1600.215 1511.955 1600.230 ;
      LAYER met3 ;
        RECT 304.000 1595.360 1496.000 1599.400 ;
        RECT 304.400 1593.960 1496.000 1595.360 ;
        RECT 304.000 1589.920 1496.000 1593.960 ;
        RECT 304.000 1588.520 1495.600 1589.920 ;
      LAYER met3 ;
        RECT 1513.465 1589.650 1513.795 1589.665 ;
        RECT 1499.140 1589.520 1513.795 1589.650 ;
        RECT 1496.000 1589.350 1513.795 1589.520 ;
        RECT 1496.000 1588.920 1500.000 1589.350 ;
        RECT 1513.465 1589.335 1513.795 1589.350 ;
      LAYER met3 ;
        RECT 304.000 1584.480 1496.000 1588.520 ;
        RECT 304.400 1583.080 1496.000 1584.480 ;
        RECT 304.000 1579.040 1496.000 1583.080 ;
        RECT 304.000 1577.640 1495.600 1579.040 ;
      LAYER met3 ;
        RECT 1513.925 1578.770 1514.255 1578.785 ;
        RECT 1499.140 1578.640 1514.255 1578.770 ;
        RECT 1496.000 1578.470 1514.255 1578.640 ;
        RECT 1496.000 1578.040 1500.000 1578.470 ;
        RECT 1513.925 1578.455 1514.255 1578.470 ;
      LAYER met3 ;
        RECT 304.000 1574.280 1496.000 1577.640 ;
        RECT 304.400 1572.880 1496.000 1574.280 ;
        RECT 304.000 1567.480 1496.000 1572.880 ;
        RECT 304.000 1566.080 1495.600 1567.480 ;
      LAYER met3 ;
        RECT 1513.925 1567.210 1514.255 1567.225 ;
        RECT 1499.140 1567.080 1514.255 1567.210 ;
        RECT 1496.000 1566.910 1514.255 1567.080 ;
        RECT 1496.000 1566.480 1500.000 1566.910 ;
        RECT 1513.925 1566.895 1514.255 1566.910 ;
      LAYER met3 ;
        RECT 304.000 1563.400 1496.000 1566.080 ;
        RECT 304.400 1562.000 1496.000 1563.400 ;
        RECT 304.000 1556.600 1496.000 1562.000 ;
        RECT 304.000 1555.200 1495.600 1556.600 ;
      LAYER met3 ;
        RECT 1513.465 1556.330 1513.795 1556.345 ;
        RECT 1499.140 1556.200 1513.795 1556.330 ;
        RECT 1496.000 1556.030 1513.795 1556.200 ;
        RECT 1496.000 1555.600 1500.000 1556.030 ;
        RECT 1513.465 1556.015 1513.795 1556.030 ;
      LAYER met3 ;
        RECT 304.000 1553.200 1496.000 1555.200 ;
        RECT 304.400 1551.800 1496.000 1553.200 ;
        RECT 304.000 1545.720 1496.000 1551.800 ;
        RECT 304.000 1544.320 1495.600 1545.720 ;
      LAYER met3 ;
        RECT 1513.925 1545.450 1514.255 1545.465 ;
        RECT 1499.140 1545.320 1514.255 1545.450 ;
        RECT 1496.000 1545.150 1514.255 1545.320 ;
        RECT 1496.000 1544.720 1500.000 1545.150 ;
        RECT 1513.925 1545.135 1514.255 1545.150 ;
      LAYER met3 ;
        RECT 304.000 1542.320 1496.000 1544.320 ;
        RECT 304.400 1540.920 1496.000 1542.320 ;
        RECT 304.000 1534.840 1496.000 1540.920 ;
        RECT 304.000 1533.440 1495.600 1534.840 ;
      LAYER met3 ;
        RECT 1513.925 1534.570 1514.255 1534.585 ;
        RECT 1499.140 1534.440 1514.255 1534.570 ;
        RECT 1496.000 1534.270 1514.255 1534.440 ;
        RECT 1496.000 1533.840 1500.000 1534.270 ;
        RECT 1513.925 1534.255 1514.255 1534.270 ;
      LAYER met3 ;
        RECT 304.000 1532.120 1496.000 1533.440 ;
        RECT 304.400 1530.720 1496.000 1532.120 ;
        RECT 304.000 1523.960 1496.000 1530.720 ;
        RECT 304.000 1522.560 1495.600 1523.960 ;
      LAYER met3 ;
        RECT 1513.925 1523.690 1514.255 1523.705 ;
        RECT 1499.140 1523.560 1514.255 1523.690 ;
        RECT 1496.000 1523.390 1514.255 1523.560 ;
        RECT 1496.000 1522.960 1500.000 1523.390 ;
        RECT 1513.925 1523.375 1514.255 1523.390 ;
      LAYER met3 ;
        RECT 304.000 1521.240 1496.000 1522.560 ;
        RECT 304.400 1519.840 1496.000 1521.240 ;
        RECT 304.000 1512.400 1496.000 1519.840 ;
        RECT 304.000 1511.040 1495.600 1512.400 ;
      LAYER met3 ;
        RECT 1513.925 1512.130 1514.255 1512.145 ;
        RECT 1499.140 1512.000 1514.255 1512.130 ;
        RECT 1496.000 1511.830 1514.255 1512.000 ;
        RECT 1496.000 1511.400 1500.000 1511.830 ;
        RECT 1513.925 1511.815 1514.255 1511.830 ;
      LAYER met3 ;
        RECT 304.400 1511.000 1495.600 1511.040 ;
        RECT 304.400 1509.640 1496.000 1511.000 ;
        RECT 304.000 1501.520 1496.000 1509.640 ;
        RECT 304.000 1500.160 1495.600 1501.520 ;
      LAYER met3 ;
        RECT 1513.465 1501.250 1513.795 1501.265 ;
        RECT 1499.140 1501.120 1513.795 1501.250 ;
        RECT 1496.000 1500.950 1513.795 1501.120 ;
        RECT 1496.000 1500.520 1500.000 1500.950 ;
        RECT 1513.465 1500.935 1513.795 1500.950 ;
      LAYER met3 ;
        RECT 304.400 1500.120 1495.600 1500.160 ;
        RECT 304.400 1498.760 1496.000 1500.120 ;
        RECT 304.000 1490.640 1496.000 1498.760 ;
        RECT 304.000 1489.960 1495.600 1490.640 ;
      LAYER met3 ;
        RECT 1513.925 1490.370 1514.255 1490.385 ;
        RECT 1499.140 1490.240 1514.255 1490.370 ;
      LAYER met3 ;
        RECT 304.400 1489.240 1495.600 1489.960 ;
      LAYER met3 ;
        RECT 1496.000 1490.070 1514.255 1490.240 ;
        RECT 1496.000 1489.640 1500.000 1490.070 ;
        RECT 1513.925 1490.055 1514.255 1490.070 ;
      LAYER met3 ;
        RECT 304.400 1488.560 1496.000 1489.240 ;
        RECT 304.000 1479.760 1496.000 1488.560 ;
        RECT 304.000 1479.080 1495.600 1479.760 ;
      LAYER met3 ;
        RECT 1513.005 1479.490 1513.335 1479.505 ;
        RECT 1499.140 1479.360 1513.335 1479.490 ;
      LAYER met3 ;
        RECT 304.400 1478.360 1495.600 1479.080 ;
      LAYER met3 ;
        RECT 1496.000 1479.190 1513.335 1479.360 ;
        RECT 1496.000 1478.760 1500.000 1479.190 ;
        RECT 1513.005 1479.175 1513.335 1479.190 ;
      LAYER met3 ;
        RECT 304.400 1477.680 1496.000 1478.360 ;
        RECT 304.000 1468.880 1496.000 1477.680 ;
        RECT 304.400 1467.480 1495.600 1468.880 ;
      LAYER met3 ;
        RECT 1513.925 1468.610 1514.255 1468.625 ;
        RECT 1499.140 1468.480 1514.255 1468.610 ;
        RECT 1496.000 1468.310 1514.255 1468.480 ;
        RECT 1496.000 1467.880 1500.000 1468.310 ;
        RECT 1513.925 1468.295 1514.255 1468.310 ;
      LAYER met3 ;
        RECT 304.000 1458.000 1496.000 1467.480 ;
        RECT 304.400 1457.320 1496.000 1458.000 ;
        RECT 304.400 1456.600 1495.600 1457.320 ;
      LAYER met3 ;
        RECT 1512.545 1457.050 1512.875 1457.065 ;
        RECT 1499.140 1456.920 1512.875 1457.050 ;
      LAYER met3 ;
        RECT 304.000 1455.920 1495.600 1456.600 ;
      LAYER met3 ;
        RECT 1496.000 1456.750 1512.875 1456.920 ;
        RECT 1496.000 1456.320 1500.000 1456.750 ;
        RECT 1512.545 1456.735 1512.875 1456.750 ;
      LAYER met3 ;
        RECT 304.000 1447.800 1496.000 1455.920 ;
        RECT 304.400 1446.440 1496.000 1447.800 ;
        RECT 304.400 1446.400 1495.600 1446.440 ;
        RECT 304.000 1445.040 1495.600 1446.400 ;
      LAYER met3 ;
        RECT 1513.465 1446.170 1513.795 1446.185 ;
        RECT 1499.140 1446.040 1513.795 1446.170 ;
        RECT 1496.000 1445.870 1513.795 1446.040 ;
        RECT 1496.000 1445.440 1500.000 1445.870 ;
        RECT 1513.465 1445.855 1513.795 1445.870 ;
      LAYER met3 ;
        RECT 304.000 1436.920 1496.000 1445.040 ;
        RECT 304.400 1435.560 1496.000 1436.920 ;
        RECT 304.400 1435.520 1495.600 1435.560 ;
        RECT 304.000 1434.160 1495.600 1435.520 ;
      LAYER met3 ;
        RECT 1513.925 1435.290 1514.255 1435.305 ;
        RECT 1499.140 1435.160 1514.255 1435.290 ;
        RECT 1496.000 1434.990 1514.255 1435.160 ;
        RECT 1496.000 1434.560 1500.000 1434.990 ;
        RECT 1513.925 1434.975 1514.255 1434.990 ;
      LAYER met3 ;
        RECT 304.000 1426.720 1496.000 1434.160 ;
        RECT 304.400 1425.320 1496.000 1426.720 ;
        RECT 304.000 1424.680 1496.000 1425.320 ;
        RECT 304.000 1423.280 1495.600 1424.680 ;
      LAYER met3 ;
        RECT 1513.465 1424.410 1513.795 1424.425 ;
        RECT 1499.140 1424.280 1513.795 1424.410 ;
        RECT 1496.000 1424.110 1513.795 1424.280 ;
        RECT 1496.000 1423.680 1500.000 1424.110 ;
        RECT 1513.465 1424.095 1513.795 1424.110 ;
      LAYER met3 ;
        RECT 304.000 1415.840 1496.000 1423.280 ;
        RECT 304.400 1414.440 1496.000 1415.840 ;
        RECT 304.000 1413.800 1496.000 1414.440 ;
        RECT 304.000 1412.400 1495.600 1413.800 ;
      LAYER met3 ;
        RECT 1512.545 1413.530 1512.875 1413.545 ;
        RECT 1499.140 1413.400 1512.875 1413.530 ;
        RECT 1496.000 1413.230 1512.875 1413.400 ;
        RECT 1496.000 1412.800 1500.000 1413.230 ;
        RECT 1512.545 1413.215 1512.875 1413.230 ;
      LAYER met3 ;
        RECT 304.000 1405.640 1496.000 1412.400 ;
        RECT 304.400 1404.240 1496.000 1405.640 ;
        RECT 304.000 1402.240 1496.000 1404.240 ;
        RECT 304.000 1400.840 1495.600 1402.240 ;
      LAYER met3 ;
        RECT 1512.545 1401.970 1512.875 1401.985 ;
        RECT 1499.140 1401.840 1512.875 1401.970 ;
        RECT 1496.000 1401.670 1512.875 1401.840 ;
        RECT 1496.000 1401.240 1500.000 1401.670 ;
        RECT 1512.545 1401.655 1512.875 1401.670 ;
      LAYER met3 ;
        RECT 304.000 1394.760 1496.000 1400.840 ;
        RECT 304.400 1393.360 1496.000 1394.760 ;
        RECT 304.000 1391.360 1496.000 1393.360 ;
        RECT 304.000 1389.960 1495.600 1391.360 ;
      LAYER met3 ;
        RECT 1511.625 1391.090 1511.955 1391.105 ;
        RECT 1499.140 1390.960 1511.955 1391.090 ;
        RECT 1496.000 1390.790 1511.955 1390.960 ;
        RECT 1496.000 1390.360 1500.000 1390.790 ;
        RECT 1511.625 1390.775 1511.955 1390.790 ;
      LAYER met3 ;
        RECT 304.000 1384.560 1496.000 1389.960 ;
        RECT 304.400 1383.160 1496.000 1384.560 ;
        RECT 304.000 1380.480 1496.000 1383.160 ;
        RECT 304.000 1379.080 1495.600 1380.480 ;
      LAYER met3 ;
        RECT 1513.005 1380.210 1513.335 1380.225 ;
        RECT 1499.140 1380.080 1513.335 1380.210 ;
        RECT 1496.000 1379.910 1513.335 1380.080 ;
        RECT 1496.000 1379.480 1500.000 1379.910 ;
        RECT 1513.005 1379.895 1513.335 1379.910 ;
      LAYER met3 ;
        RECT 304.000 1373.680 1496.000 1379.080 ;
        RECT 304.400 1372.280 1496.000 1373.680 ;
        RECT 304.000 1369.600 1496.000 1372.280 ;
        RECT 304.000 1368.200 1495.600 1369.600 ;
      LAYER met3 ;
        RECT 1513.925 1369.330 1514.255 1369.345 ;
        RECT 1499.140 1369.200 1514.255 1369.330 ;
        RECT 1496.000 1369.030 1514.255 1369.200 ;
        RECT 1496.000 1368.600 1500.000 1369.030 ;
        RECT 1513.925 1369.015 1514.255 1369.030 ;
      LAYER met3 ;
        RECT 304.000 1363.480 1496.000 1368.200 ;
        RECT 304.400 1362.080 1496.000 1363.480 ;
        RECT 304.000 1358.720 1496.000 1362.080 ;
        RECT 304.000 1357.320 1495.600 1358.720 ;
      LAYER met3 ;
        RECT 1512.545 1358.450 1512.875 1358.465 ;
        RECT 1499.140 1358.320 1512.875 1358.450 ;
        RECT 1496.000 1358.150 1512.875 1358.320 ;
        RECT 1496.000 1357.720 1500.000 1358.150 ;
        RECT 1512.545 1358.135 1512.875 1358.150 ;
      LAYER met3 ;
        RECT 304.000 1352.600 1496.000 1357.320 ;
        RECT 304.400 1351.200 1496.000 1352.600 ;
        RECT 304.000 1347.160 1496.000 1351.200 ;
        RECT 304.000 1345.760 1495.600 1347.160 ;
      LAYER met3 ;
        RECT 1512.545 1346.890 1512.875 1346.905 ;
        RECT 1499.140 1346.760 1512.875 1346.890 ;
        RECT 1496.000 1346.590 1512.875 1346.760 ;
        RECT 1496.000 1346.160 1500.000 1346.590 ;
        RECT 1512.545 1346.575 1512.875 1346.590 ;
      LAYER met3 ;
        RECT 304.000 1342.400 1496.000 1345.760 ;
        RECT 304.400 1341.000 1496.000 1342.400 ;
        RECT 304.000 1336.280 1496.000 1341.000 ;
        RECT 304.000 1334.880 1495.600 1336.280 ;
      LAYER met3 ;
        RECT 1511.625 1336.010 1511.955 1336.025 ;
        RECT 1499.140 1335.880 1511.955 1336.010 ;
        RECT 1496.000 1335.710 1511.955 1335.880 ;
        RECT 1496.000 1335.280 1500.000 1335.710 ;
        RECT 1511.625 1335.695 1511.955 1335.710 ;
      LAYER met3 ;
        RECT 304.000 1331.520 1496.000 1334.880 ;
        RECT 304.400 1330.120 1496.000 1331.520 ;
        RECT 304.000 1325.400 1496.000 1330.120 ;
        RECT 304.000 1324.000 1495.600 1325.400 ;
      LAYER met3 ;
        RECT 1513.005 1325.130 1513.335 1325.145 ;
        RECT 1499.140 1325.000 1513.335 1325.130 ;
        RECT 1496.000 1324.830 1513.335 1325.000 ;
        RECT 1496.000 1324.400 1500.000 1324.830 ;
        RECT 1513.005 1324.815 1513.335 1324.830 ;
      LAYER met3 ;
        RECT 304.000 1321.320 1496.000 1324.000 ;
        RECT 304.400 1319.920 1496.000 1321.320 ;
        RECT 304.000 1314.520 1496.000 1319.920 ;
        RECT 304.000 1313.120 1495.600 1314.520 ;
      LAYER met3 ;
        RECT 1513.925 1314.250 1514.255 1314.265 ;
        RECT 1499.140 1314.120 1514.255 1314.250 ;
        RECT 1496.000 1313.950 1514.255 1314.120 ;
        RECT 1496.000 1313.520 1500.000 1313.950 ;
        RECT 1513.925 1313.935 1514.255 1313.950 ;
      LAYER met3 ;
        RECT 304.000 1310.440 1496.000 1313.120 ;
        RECT 304.400 1309.040 1496.000 1310.440 ;
        RECT 304.000 1303.640 1496.000 1309.040 ;
        RECT 304.000 1302.240 1495.600 1303.640 ;
      LAYER met3 ;
        RECT 1512.545 1303.370 1512.875 1303.385 ;
        RECT 1499.140 1303.240 1512.875 1303.370 ;
        RECT 1496.000 1303.070 1512.875 1303.240 ;
        RECT 1496.000 1302.640 1500.000 1303.070 ;
        RECT 1512.545 1303.055 1512.875 1303.070 ;
      LAYER met3 ;
        RECT 304.000 1300.240 1496.000 1302.240 ;
        RECT 304.400 1298.840 1496.000 1300.240 ;
        RECT 304.000 1292.760 1496.000 1298.840 ;
        RECT 304.000 1291.360 1495.600 1292.760 ;
      LAYER met3 ;
        RECT 1512.085 1292.490 1512.415 1292.505 ;
        RECT 1499.140 1292.360 1512.415 1292.490 ;
        RECT 1496.000 1292.190 1512.415 1292.360 ;
        RECT 1496.000 1291.760 1500.000 1292.190 ;
        RECT 1512.085 1292.175 1512.415 1292.190 ;
      LAYER met3 ;
        RECT 304.000 1290.040 1496.000 1291.360 ;
        RECT 304.400 1288.640 1496.000 1290.040 ;
        RECT 304.000 1281.200 1496.000 1288.640 ;
        RECT 304.000 1279.800 1495.600 1281.200 ;
      LAYER met3 ;
        RECT 1511.625 1280.930 1511.955 1280.945 ;
        RECT 1499.140 1280.800 1511.955 1280.930 ;
        RECT 1496.000 1280.630 1511.955 1280.800 ;
        RECT 1496.000 1280.200 1500.000 1280.630 ;
        RECT 1511.625 1280.615 1511.955 1280.630 ;
      LAYER met3 ;
        RECT 304.000 1279.160 1496.000 1279.800 ;
        RECT 304.400 1277.760 1496.000 1279.160 ;
        RECT 304.000 1270.320 1496.000 1277.760 ;
        RECT 304.000 1268.960 1495.600 1270.320 ;
      LAYER met3 ;
        RECT 1512.545 1270.050 1512.875 1270.065 ;
        RECT 1499.140 1269.920 1512.875 1270.050 ;
        RECT 1496.000 1269.750 1512.875 1269.920 ;
        RECT 1496.000 1269.320 1500.000 1269.750 ;
        RECT 1512.545 1269.735 1512.875 1269.750 ;
      LAYER met3 ;
        RECT 304.400 1268.920 1495.600 1268.960 ;
        RECT 304.400 1267.560 1496.000 1268.920 ;
        RECT 304.000 1259.440 1496.000 1267.560 ;
        RECT 304.000 1258.080 1495.600 1259.440 ;
      LAYER met3 ;
        RECT 1513.925 1259.170 1514.255 1259.185 ;
        RECT 1499.140 1259.040 1514.255 1259.170 ;
        RECT 1496.000 1258.870 1514.255 1259.040 ;
        RECT 1496.000 1258.440 1500.000 1258.870 ;
        RECT 1513.925 1258.855 1514.255 1258.870 ;
      LAYER met3 ;
        RECT 304.400 1258.040 1495.600 1258.080 ;
        RECT 304.400 1256.680 1496.000 1258.040 ;
        RECT 304.000 1248.560 1496.000 1256.680 ;
        RECT 304.000 1247.880 1495.600 1248.560 ;
      LAYER met3 ;
        RECT 1513.925 1248.290 1514.255 1248.305 ;
        RECT 1499.140 1248.160 1514.255 1248.290 ;
      LAYER met3 ;
        RECT 304.400 1247.160 1495.600 1247.880 ;
      LAYER met3 ;
        RECT 1496.000 1247.990 1514.255 1248.160 ;
        RECT 1496.000 1247.560 1500.000 1247.990 ;
        RECT 1513.925 1247.975 1514.255 1247.990 ;
      LAYER met3 ;
        RECT 304.400 1246.480 1496.000 1247.160 ;
        RECT 304.000 1237.680 1496.000 1246.480 ;
        RECT 304.000 1237.000 1495.600 1237.680 ;
      LAYER met3 ;
        RECT 1512.085 1237.410 1512.415 1237.425 ;
        RECT 1499.140 1237.280 1512.415 1237.410 ;
      LAYER met3 ;
        RECT 304.400 1236.280 1495.600 1237.000 ;
      LAYER met3 ;
        RECT 1496.000 1237.110 1512.415 1237.280 ;
        RECT 1496.000 1236.680 1500.000 1237.110 ;
        RECT 1512.085 1237.095 1512.415 1237.110 ;
      LAYER met3 ;
        RECT 304.400 1235.600 1496.000 1236.280 ;
        RECT 304.000 1226.800 1496.000 1235.600 ;
        RECT 304.400 1226.120 1496.000 1226.800 ;
        RECT 304.400 1225.400 1495.600 1226.120 ;
      LAYER met3 ;
        RECT 1513.465 1225.850 1513.795 1225.865 ;
        RECT 1499.140 1225.720 1513.795 1225.850 ;
      LAYER met3 ;
        RECT 304.000 1224.720 1495.600 1225.400 ;
      LAYER met3 ;
        RECT 1496.000 1225.550 1513.795 1225.720 ;
        RECT 1496.000 1225.120 1500.000 1225.550 ;
        RECT 1513.465 1225.535 1513.795 1225.550 ;
      LAYER met3 ;
        RECT 304.000 1215.920 1496.000 1224.720 ;
        RECT 304.400 1215.240 1496.000 1215.920 ;
        RECT 304.400 1214.520 1495.600 1215.240 ;
      LAYER met3 ;
        RECT 1512.545 1214.970 1512.875 1214.985 ;
        RECT 1499.140 1214.840 1512.875 1214.970 ;
      LAYER met3 ;
        RECT 304.000 1213.840 1495.600 1214.520 ;
      LAYER met3 ;
        RECT 1496.000 1214.670 1512.875 1214.840 ;
        RECT 1496.000 1214.240 1500.000 1214.670 ;
        RECT 1512.545 1214.655 1512.875 1214.670 ;
      LAYER met3 ;
        RECT 304.000 1205.720 1496.000 1213.840 ;
        RECT 304.400 1204.360 1496.000 1205.720 ;
        RECT 304.400 1204.320 1495.600 1204.360 ;
        RECT 304.000 1202.960 1495.600 1204.320 ;
      LAYER met3 ;
        RECT 1513.925 1204.090 1514.255 1204.105 ;
        RECT 1499.140 1203.960 1514.255 1204.090 ;
        RECT 1496.000 1203.790 1514.255 1203.960 ;
        RECT 1496.000 1203.360 1500.000 1203.790 ;
        RECT 1513.925 1203.775 1514.255 1203.790 ;
      LAYER met3 ;
        RECT 304.000 1194.840 1496.000 1202.960 ;
        RECT 304.400 1193.480 1496.000 1194.840 ;
        RECT 304.400 1193.440 1495.600 1193.480 ;
        RECT 304.000 1192.080 1495.600 1193.440 ;
      LAYER met3 ;
        RECT 1513.925 1193.210 1514.255 1193.225 ;
        RECT 1499.140 1193.080 1514.255 1193.210 ;
        RECT 1496.000 1192.910 1514.255 1193.080 ;
        RECT 1496.000 1192.480 1500.000 1192.910 ;
        RECT 1513.925 1192.895 1514.255 1192.910 ;
      LAYER met3 ;
        RECT 304.000 1184.640 1496.000 1192.080 ;
        RECT 304.400 1183.240 1496.000 1184.640 ;
        RECT 304.000 1182.600 1496.000 1183.240 ;
        RECT 304.000 1181.200 1495.600 1182.600 ;
      LAYER met3 ;
        RECT 1512.085 1182.330 1512.415 1182.345 ;
        RECT 1499.140 1182.200 1512.415 1182.330 ;
        RECT 1496.000 1182.030 1512.415 1182.200 ;
        RECT 1496.000 1181.600 1500.000 1182.030 ;
        RECT 1512.085 1182.015 1512.415 1182.030 ;
      LAYER met3 ;
        RECT 304.000 1173.760 1496.000 1181.200 ;
        RECT 304.400 1172.360 1496.000 1173.760 ;
        RECT 304.000 1171.040 1496.000 1172.360 ;
        RECT 304.000 1169.640 1495.600 1171.040 ;
      LAYER met3 ;
        RECT 1513.465 1170.770 1513.795 1170.785 ;
        RECT 1499.140 1170.640 1513.795 1170.770 ;
        RECT 1496.000 1170.470 1513.795 1170.640 ;
        RECT 1496.000 1170.040 1500.000 1170.470 ;
        RECT 1513.465 1170.455 1513.795 1170.470 ;
      LAYER met3 ;
        RECT 304.000 1163.560 1496.000 1169.640 ;
        RECT 304.400 1162.160 1496.000 1163.560 ;
        RECT 304.000 1160.160 1496.000 1162.160 ;
        RECT 304.000 1158.760 1495.600 1160.160 ;
      LAYER met3 ;
        RECT 1512.545 1159.890 1512.875 1159.905 ;
        RECT 1499.140 1159.760 1512.875 1159.890 ;
        RECT 1496.000 1159.590 1512.875 1159.760 ;
        RECT 1496.000 1159.160 1500.000 1159.590 ;
        RECT 1512.545 1159.575 1512.875 1159.590 ;
      LAYER met3 ;
        RECT 304.000 1152.680 1496.000 1158.760 ;
        RECT 304.400 1151.280 1496.000 1152.680 ;
        RECT 304.000 1149.280 1496.000 1151.280 ;
        RECT 304.000 1147.880 1495.600 1149.280 ;
      LAYER met3 ;
        RECT 1513.925 1149.010 1514.255 1149.025 ;
        RECT 1499.140 1148.880 1514.255 1149.010 ;
        RECT 1496.000 1148.710 1514.255 1148.880 ;
        RECT 1496.000 1148.280 1500.000 1148.710 ;
        RECT 1513.925 1148.695 1514.255 1148.710 ;
      LAYER met3 ;
        RECT 304.000 1142.480 1496.000 1147.880 ;
        RECT 304.400 1141.080 1496.000 1142.480 ;
        RECT 304.000 1138.400 1496.000 1141.080 ;
        RECT 304.000 1137.000 1495.600 1138.400 ;
      LAYER met3 ;
        RECT 1513.925 1138.130 1514.255 1138.145 ;
        RECT 1499.140 1138.000 1514.255 1138.130 ;
        RECT 1496.000 1137.830 1514.255 1138.000 ;
        RECT 1496.000 1137.400 1500.000 1137.830 ;
        RECT 1513.925 1137.815 1514.255 1137.830 ;
      LAYER met3 ;
        RECT 304.000 1131.600 1496.000 1137.000 ;
        RECT 304.400 1130.200 1496.000 1131.600 ;
        RECT 304.000 1127.520 1496.000 1130.200 ;
        RECT 304.000 1126.120 1495.600 1127.520 ;
      LAYER met3 ;
        RECT 1513.925 1127.250 1514.255 1127.265 ;
        RECT 1499.140 1127.120 1514.255 1127.250 ;
        RECT 1496.000 1126.950 1514.255 1127.120 ;
        RECT 1496.000 1126.520 1500.000 1126.950 ;
        RECT 1513.925 1126.935 1514.255 1126.950 ;
      LAYER met3 ;
        RECT 304.000 1121.400 1496.000 1126.120 ;
        RECT 304.400 1120.000 1496.000 1121.400 ;
        RECT 304.000 1115.960 1496.000 1120.000 ;
        RECT 304.000 1114.560 1495.600 1115.960 ;
      LAYER met3 ;
        RECT 1513.465 1115.690 1513.795 1115.705 ;
        RECT 1499.140 1115.560 1513.795 1115.690 ;
        RECT 1496.000 1115.390 1513.795 1115.560 ;
        RECT 1496.000 1114.960 1500.000 1115.390 ;
        RECT 1513.465 1115.375 1513.795 1115.390 ;
      LAYER met3 ;
        RECT 304.000 1110.520 1496.000 1114.560 ;
        RECT 304.400 1109.120 1496.000 1110.520 ;
        RECT 304.000 1105.080 1496.000 1109.120 ;
        RECT 304.000 1103.680 1495.600 1105.080 ;
      LAYER met3 ;
        RECT 1513.925 1104.810 1514.255 1104.825 ;
        RECT 1499.140 1104.680 1514.255 1104.810 ;
        RECT 1496.000 1104.510 1514.255 1104.680 ;
        RECT 1496.000 1104.080 1500.000 1104.510 ;
        RECT 1513.925 1104.495 1514.255 1104.510 ;
      LAYER met3 ;
        RECT 304.000 1100.320 1496.000 1103.680 ;
        RECT 304.400 1098.920 1496.000 1100.320 ;
        RECT 304.000 1094.200 1496.000 1098.920 ;
        RECT 304.000 1092.800 1495.600 1094.200 ;
      LAYER met3 ;
        RECT 1513.925 1093.930 1514.255 1093.945 ;
        RECT 1499.140 1093.800 1514.255 1093.930 ;
        RECT 1496.000 1093.630 1514.255 1093.800 ;
        RECT 1496.000 1093.200 1500.000 1093.630 ;
        RECT 1513.925 1093.615 1514.255 1093.630 ;
      LAYER met3 ;
        RECT 304.000 1089.440 1496.000 1092.800 ;
        RECT 304.400 1088.040 1496.000 1089.440 ;
        RECT 304.000 1083.320 1496.000 1088.040 ;
        RECT 304.000 1081.920 1495.600 1083.320 ;
      LAYER met3 ;
        RECT 1513.925 1083.050 1514.255 1083.065 ;
        RECT 1499.140 1082.920 1514.255 1083.050 ;
        RECT 1496.000 1082.750 1514.255 1082.920 ;
        RECT 1496.000 1082.320 1500.000 1082.750 ;
        RECT 1513.925 1082.735 1514.255 1082.750 ;
      LAYER met3 ;
        RECT 304.000 1079.240 1496.000 1081.920 ;
        RECT 304.400 1077.840 1496.000 1079.240 ;
        RECT 304.000 1072.440 1496.000 1077.840 ;
        RECT 304.000 1071.040 1495.600 1072.440 ;
      LAYER met3 ;
        RECT 1513.925 1072.170 1514.255 1072.185 ;
        RECT 1499.140 1072.040 1514.255 1072.170 ;
        RECT 1496.000 1071.870 1514.255 1072.040 ;
        RECT 1496.000 1071.440 1500.000 1071.870 ;
        RECT 1513.925 1071.855 1514.255 1071.870 ;
      LAYER met3 ;
        RECT 304.000 1068.360 1496.000 1071.040 ;
        RECT 304.400 1066.960 1496.000 1068.360 ;
        RECT 304.000 1060.880 1496.000 1066.960 ;
        RECT 304.000 1059.480 1495.600 1060.880 ;
      LAYER met3 ;
        RECT 1513.005 1060.610 1513.335 1060.625 ;
        RECT 1499.140 1060.480 1513.335 1060.610 ;
        RECT 1496.000 1060.310 1513.335 1060.480 ;
        RECT 1496.000 1059.880 1500.000 1060.310 ;
        RECT 1513.005 1060.295 1513.335 1060.310 ;
      LAYER met3 ;
        RECT 304.000 1058.160 1496.000 1059.480 ;
        RECT 304.400 1056.760 1496.000 1058.160 ;
        RECT 304.000 1050.000 1496.000 1056.760 ;
        RECT 304.000 1048.600 1495.600 1050.000 ;
      LAYER met3 ;
        RECT 1513.925 1049.730 1514.255 1049.745 ;
        RECT 1499.140 1049.600 1514.255 1049.730 ;
        RECT 1496.000 1049.430 1514.255 1049.600 ;
        RECT 1496.000 1049.000 1500.000 1049.430 ;
        RECT 1513.925 1049.415 1514.255 1049.430 ;
      LAYER met3 ;
        RECT 304.000 1047.280 1496.000 1048.600 ;
        RECT 304.400 1045.880 1496.000 1047.280 ;
        RECT 304.000 1039.120 1496.000 1045.880 ;
        RECT 304.000 1037.720 1495.600 1039.120 ;
      LAYER met3 ;
        RECT 1513.925 1038.850 1514.255 1038.865 ;
        RECT 1499.140 1038.720 1514.255 1038.850 ;
        RECT 1496.000 1038.550 1514.255 1038.720 ;
        RECT 1496.000 1038.120 1500.000 1038.550 ;
        RECT 1513.925 1038.535 1514.255 1038.550 ;
      LAYER met3 ;
        RECT 304.000 1037.080 1496.000 1037.720 ;
        RECT 304.400 1035.680 1496.000 1037.080 ;
        RECT 304.000 1028.240 1496.000 1035.680 ;
        RECT 304.000 1026.840 1495.600 1028.240 ;
      LAYER met3 ;
        RECT 1513.925 1027.970 1514.255 1027.985 ;
        RECT 1499.140 1027.840 1514.255 1027.970 ;
        RECT 1496.000 1027.670 1514.255 1027.840 ;
        RECT 1496.000 1027.240 1500.000 1027.670 ;
        RECT 1513.925 1027.655 1514.255 1027.670 ;
      LAYER met3 ;
        RECT 304.000 1026.200 1496.000 1026.840 ;
        RECT 304.400 1024.800 1496.000 1026.200 ;
        RECT 304.000 1017.360 1496.000 1024.800 ;
        RECT 304.000 1016.000 1495.600 1017.360 ;
      LAYER met3 ;
        RECT 1511.165 1017.090 1511.495 1017.105 ;
        RECT 1499.140 1016.960 1511.495 1017.090 ;
        RECT 1496.000 1016.790 1511.495 1016.960 ;
        RECT 1496.000 1016.360 1500.000 1016.790 ;
        RECT 1511.165 1016.775 1511.495 1016.790 ;
      LAYER met3 ;
        RECT 304.400 1015.960 1495.600 1016.000 ;
        RECT 304.400 1014.600 1496.000 1015.960 ;
        RECT 304.000 1006.480 1496.000 1014.600 ;
        RECT 304.000 1005.800 1495.600 1006.480 ;
      LAYER met3 ;
        RECT 1514.385 1006.210 1514.715 1006.225 ;
        RECT 1499.140 1006.080 1514.715 1006.210 ;
      LAYER met3 ;
        RECT 304.400 1005.080 1495.600 1005.800 ;
      LAYER met3 ;
        RECT 1496.000 1005.910 1514.715 1006.080 ;
        RECT 1496.000 1005.480 1500.000 1005.910 ;
        RECT 1514.385 1005.895 1514.715 1005.910 ;
      LAYER met3 ;
        RECT 304.400 1004.400 1496.000 1005.080 ;
        RECT 304.000 1004.255 1496.000 1004.400 ;
      LAYER via3 ;
        RECT 668.220 2767.100 668.540 2767.420 ;
        RECT 1295.660 2767.100 1295.980 2767.420 ;
        RECT 1318.660 2767.100 1318.980 2767.420 ;
        RECT 1892.740 2767.100 1893.060 2767.420 ;
        RECT 1914.820 2767.100 1915.140 2767.420 ;
        RECT 2539.500 2767.100 2539.820 2767.420 ;
        RECT 2567.100 2767.100 2567.420 2767.420 ;
        RECT 646.140 2755.540 646.460 2755.860 ;
        RECT 664.540 2755.540 664.860 2755.860 ;
        RECT 2570.780 2753.500 2571.100 2753.820 ;
        RECT 1759.200 2297.900 1759.520 2298.220 ;
        RECT 386.560 2297.220 386.880 2297.540 ;
        RECT 1636.560 2297.220 1636.880 2297.540 ;
        RECT 1642.400 2297.220 1642.720 2297.540 ;
        RECT 1644.340 2297.220 1644.660 2297.540 ;
        RECT 1794.240 2297.220 1794.560 2297.540 ;
        RECT 2263.200 2297.220 2263.520 2297.540 ;
        RECT 2265.340 2297.220 2265.660 2297.540 ;
        RECT 2415.040 2297.220 2415.360 2297.540 ;
        RECT 369.220 2290.420 369.540 2290.740 ;
        RECT 374.740 2290.420 375.060 2290.740 ;
        RECT 396.820 2290.420 397.140 2290.740 ;
        RECT 409.700 2290.420 410.020 2290.740 ;
        RECT 414.300 2290.420 414.620 2290.740 ;
        RECT 420.740 2290.420 421.060 2290.740 ;
        RECT 427.180 2290.420 427.500 2290.740 ;
        RECT 431.780 2290.420 432.100 2290.740 ;
        RECT 439.140 2290.420 439.460 2290.740 ;
        RECT 444.660 2290.420 444.980 2290.740 ;
        RECT 451.100 2290.420 451.420 2290.740 ;
        RECT 456.620 2290.420 456.940 2290.740 ;
        RECT 462.140 2290.420 462.460 2290.740 ;
        RECT 467.660 2290.420 467.980 2290.740 ;
        RECT 474.100 2290.420 474.420 2290.740 ;
        RECT 478.700 2290.420 479.020 2290.740 ;
        RECT 486.060 2290.420 486.380 2290.740 ;
        RECT 491.580 2290.420 491.900 2290.740 ;
        RECT 497.100 2290.420 497.420 2290.740 ;
        RECT 500.780 2290.420 501.100 2290.740 ;
        RECT 509.980 2290.420 510.300 2290.740 ;
        RECT 513.660 2290.420 513.980 2290.740 ;
        RECT 515.500 2290.420 515.820 2290.740 ;
        RECT 521.020 2290.420 521.340 2290.740 ;
        RECT 523.780 2290.420 524.100 2290.740 ;
        RECT 526.540 2290.420 526.860 2290.740 ;
        RECT 527.460 2290.420 527.780 2290.740 ;
        RECT 535.740 2290.420 536.060 2290.740 ;
        RECT 544.020 2290.420 544.340 2290.740 ;
        RECT 544.940 2290.420 545.260 2290.740 ;
        RECT 1001.260 2290.420 1001.580 2290.740 ;
        RECT 1052.780 2290.420 1053.100 2290.740 ;
        RECT 1060.140 2290.420 1060.460 2290.740 ;
        RECT 1065.660 2290.420 1065.980 2290.740 ;
        RECT 1070.260 2290.420 1070.580 2290.740 ;
        RECT 1076.700 2290.420 1077.020 2290.740 ;
        RECT 1083.140 2290.420 1083.460 2290.740 ;
        RECT 1087.740 2290.420 1088.060 2290.740 ;
        RECT 1094.180 2290.420 1094.500 2290.740 ;
        RECT 1100.620 2290.420 1100.940 2290.740 ;
        RECT 1107.060 2290.420 1107.380 2290.740 ;
        RECT 1112.580 2290.420 1112.900 2290.740 ;
        RECT 1118.100 2290.420 1118.420 2290.740 ;
        RECT 1121.780 2290.420 1122.100 2290.740 ;
        RECT 1129.140 2290.420 1129.460 2290.740 ;
        RECT 1135.580 2290.420 1135.900 2290.740 ;
        RECT 1142.020 2290.420 1142.340 2290.740 ;
        RECT 1147.540 2290.420 1147.860 2290.740 ;
        RECT 1164.100 2290.420 1164.420 2290.740 ;
        RECT 1167.780 2290.420 1168.100 2290.740 ;
        RECT 1613.980 2290.420 1614.300 2290.740 ;
        RECT 1619.500 2290.420 1619.820 2290.740 ;
        RECT 1631.460 2290.420 1631.780 2290.740 ;
        RECT 1636.980 2290.420 1637.300 2290.740 ;
        RECT 1644.340 2290.420 1644.660 2290.740 ;
        RECT 1654.460 2290.420 1654.780 2290.740 ;
        RECT 1659.060 2290.420 1659.380 2290.740 ;
        RECT 1665.500 2290.420 1665.820 2290.740 ;
        RECT 1670.100 2290.420 1670.420 2290.740 ;
        RECT 1676.540 2290.420 1676.860 2290.740 ;
        RECT 1682.980 2290.420 1683.300 2290.740 ;
        RECT 1688.500 2290.420 1688.820 2290.740 ;
        RECT 1694.940 2290.420 1695.260 2290.740 ;
        RECT 1699.540 2290.420 1699.860 2290.740 ;
        RECT 1705.980 2290.420 1706.300 2290.740 ;
        RECT 1713.340 2290.420 1713.660 2290.740 ;
        RECT 1719.780 2290.420 1720.100 2290.740 ;
        RECT 1723.460 2290.420 1723.780 2290.740 ;
        RECT 1730.820 2290.420 1731.140 2290.740 ;
        RECT 1736.340 2290.420 1736.660 2290.740 ;
        RECT 1741.860 2290.420 1742.180 2290.740 ;
        RECT 1748.300 2290.420 1748.620 2290.740 ;
        RECT 1764.860 2290.420 1765.180 2290.740 ;
        RECT 1767.620 2290.420 1767.940 2290.740 ;
        RECT 2308.580 2290.420 2308.900 2290.740 ;
        RECT 2315.020 2290.420 2315.340 2290.740 ;
        RECT 2321.460 2290.420 2321.780 2290.740 ;
        RECT 2326.060 2290.420 2326.380 2290.740 ;
        RECT 2343.540 2290.420 2343.860 2290.740 ;
        RECT 2349.980 2290.420 2350.300 2290.740 ;
        RECT 2356.420 2290.420 2356.740 2290.740 ;
        RECT 2361.020 2290.420 2361.340 2290.740 ;
        RECT 2367.460 2290.420 2367.780 2290.740 ;
        RECT 2373.900 2290.420 2374.220 2290.740 ;
        RECT 2377.580 2290.420 2377.900 2290.740 ;
        RECT 2384.940 2290.420 2385.260 2290.740 ;
        RECT 2391.380 2290.420 2391.700 2290.740 ;
        RECT 2396.900 2290.420 2397.220 2290.740 ;
        RECT 2415.300 2290.420 2415.620 2290.740 ;
        RECT 2420.820 2290.420 2421.140 2290.740 ;
        RECT 2427.260 2290.420 2427.580 2290.740 ;
        RECT 403.260 2289.740 403.580 2290.060 ;
        RECT 502.620 2289.740 502.940 2290.060 ;
        RECT 507.220 2289.740 507.540 2290.060 ;
        RECT 532.060 2289.740 532.380 2290.060 ;
        RECT 538.500 2289.740 538.820 2290.060 ;
        RECT 542.180 2289.740 542.500 2290.060 ;
        RECT 987.460 2289.740 987.780 2290.060 ;
        RECT 995.740 2289.740 996.060 2290.060 ;
        RECT 1035.300 2289.740 1035.620 2290.060 ;
        RECT 1173.300 2289.740 1173.620 2290.060 ;
        RECT 1613.060 2289.740 1613.380 2290.060 ;
        RECT 1617.660 2289.740 1617.980 2290.060 ;
        RECT 1648.020 2289.740 1648.340 2290.060 ;
        RECT 1712.420 2289.740 1712.740 2290.060 ;
        RECT 1717.940 2289.740 1718.260 2290.060 ;
        RECT 1729.900 2289.740 1730.220 2290.060 ;
        RECT 1734.500 2289.740 1734.820 2290.060 ;
        RECT 1740.940 2289.740 1741.260 2290.060 ;
        RECT 1747.380 2289.740 1747.700 2290.060 ;
        RECT 1752.900 2289.740 1753.220 2290.060 ;
        RECT 1782.340 2289.740 1782.660 2290.060 ;
        RECT 2297.540 2289.740 2297.860 2290.060 ;
        RECT 2338.940 2289.740 2339.260 2290.060 ;
        RECT 2403.340 2289.740 2403.660 2290.060 ;
        RECT 2438.300 2289.740 2438.620 2290.060 ;
        RECT 392.220 2289.060 392.540 2289.380 ;
        RECT 509.060 2289.060 509.380 2289.380 ;
        RECT 1159.500 2289.060 1159.820 2289.380 ;
        RECT 1182.500 2289.060 1182.820 2289.380 ;
        RECT 1587.300 2289.060 1587.620 2289.380 ;
        RECT 1624.100 2289.060 1624.420 2289.380 ;
        RECT 1630.540 2289.060 1630.860 2289.380 ;
        RECT 1652.620 2289.060 1652.940 2289.380 ;
        RECT 1775.900 2289.060 1776.220 2289.380 ;
        RECT 2292.940 2289.060 2293.260 2289.380 ;
        RECT 2332.500 2289.060 2332.820 2289.380 ;
        RECT 2397.820 2289.060 2398.140 2289.380 ;
        RECT 2404.260 2289.060 2404.580 2289.380 ;
        RECT 2423.580 2289.060 2423.900 2289.380 ;
        RECT 363.700 2288.380 364.020 2288.700 ;
        RECT 1007.700 2288.380 1008.020 2288.700 ;
        RECT 1048.180 2288.380 1048.500 2288.700 ;
        RECT 1187.100 2288.380 1187.420 2288.700 ;
        RECT 1194.460 2288.380 1194.780 2288.700 ;
        RECT 1659.980 2288.380 1660.300 2288.700 ;
        RECT 1724.380 2288.380 1724.700 2288.700 ;
        RECT 1786.940 2288.380 1787.260 2288.700 ;
        RECT 2303.980 2288.380 2304.300 2288.700 ;
        RECT 2407.940 2288.380 2408.260 2288.700 ;
        RECT 2430.020 2288.380 2430.340 2288.700 ;
        RECT 2442.900 2288.380 2443.220 2288.700 ;
        RECT 379.340 2287.700 379.660 2288.020 ;
        RECT 983.780 2287.700 984.100 2288.020 ;
        RECT 1153.060 2287.700 1153.380 2288.020 ;
        RECT 2287.420 2287.700 2287.740 2288.020 ;
        RECT 2298.460 2287.700 2298.780 2288.020 ;
        RECT 2439.220 2287.700 2439.540 2288.020 ;
        RECT 371.060 2287.020 371.380 2287.340 ;
        RECT 381.180 2287.020 381.500 2287.340 ;
        RECT 1042.660 2287.020 1042.980 2287.340 ;
        RECT 1081.300 2287.020 1081.620 2287.340 ;
        RECT 2269.020 2287.020 2269.340 2287.340 ;
        RECT 2275.460 2287.020 2275.780 2287.340 ;
        RECT 2418.060 2287.020 2418.380 2287.340 ;
        RECT 2432.780 2287.020 2433.100 2287.340 ;
        RECT 2444.740 2287.020 2445.060 2287.340 ;
        RECT 1030.700 2286.340 1031.020 2286.660 ;
        RECT 1648.940 2286.340 1649.260 2286.660 ;
        RECT 2385.860 2286.340 2386.180 2286.660 ;
        RECT 2392.300 2286.340 2392.620 2286.660 ;
        RECT 364.620 2285.660 364.940 2285.980 ;
        RECT 386.700 2285.660 387.020 2285.980 ;
        RECT 475.020 2285.660 475.340 2285.980 ;
        RECT 492.500 2285.660 492.820 2285.980 ;
        RECT 1012.300 2285.660 1012.620 2285.980 ;
        RECT 1013.220 2285.660 1013.540 2285.980 ;
        RECT 1031.620 2285.660 1031.940 2285.980 ;
        RECT 1049.100 2285.660 1049.420 2285.980 ;
        RECT 1072.100 2285.660 1072.420 2285.980 ;
        RECT 1084.060 2285.660 1084.380 2285.980 ;
        RECT 1101.540 2285.660 1101.860 2285.980 ;
        RECT 1625.020 2285.660 1625.340 2285.980 ;
        RECT 1642.500 2285.660 1642.820 2285.980 ;
        RECT 1677.460 2285.660 1677.780 2285.980 ;
        RECT 1706.900 2285.660 1707.220 2285.980 ;
        RECT 1771.300 2285.660 1771.620 2285.980 ;
        RECT 2257.060 2285.660 2257.380 2285.980 ;
        RECT 2273.620 2285.660 2273.940 2285.980 ;
        RECT 2291.100 2285.660 2291.420 2285.980 ;
        RECT 2310.420 2285.660 2310.740 2285.980 ;
        RECT 2345.380 2285.660 2345.700 2285.980 ;
        RECT 2362.860 2285.660 2363.180 2285.980 ;
        RECT 2380.340 2285.660 2380.660 2285.980 ;
        RECT 2409.780 2285.660 2410.100 2285.980 ;
        RECT 350.820 2284.980 351.140 2285.300 ;
        RECT 375.660 2284.980 375.980 2285.300 ;
        RECT 393.140 2284.980 393.460 2285.300 ;
        RECT 465.820 2284.980 466.140 2285.300 ;
        RECT 1025.180 2284.980 1025.500 2285.300 ;
        RECT 1128.220 2284.980 1128.540 2285.300 ;
        RECT 1163.180 2284.980 1163.500 2285.300 ;
        RECT 1604.780 2284.980 1605.100 2285.300 ;
        RECT 1689.420 2284.980 1689.740 2285.300 ;
        RECT 1765.780 2284.980 1766.100 2285.300 ;
        RECT 2239.580 2284.980 2239.900 2285.300 ;
        RECT 2280.060 2284.980 2280.380 2285.300 ;
        RECT 334.260 2284.300 334.580 2284.620 ;
        RECT 339.780 2284.300 340.100 2284.620 ;
        RECT 348.980 2284.300 349.300 2284.620 ;
        RECT 357.260 2284.300 357.580 2284.620 ;
        RECT 398.660 2284.300 398.980 2284.620 ;
        RECT 404.180 2284.300 404.500 2284.620 ;
        RECT 410.620 2284.300 410.940 2284.620 ;
        RECT 416.140 2284.300 416.460 2284.620 ;
        RECT 421.660 2284.300 421.980 2284.620 ;
        RECT 428.100 2284.300 428.420 2284.620 ;
        RECT 433.620 2284.300 433.940 2284.620 ;
        RECT 440.060 2284.300 440.380 2284.620 ;
        RECT 445.580 2284.300 445.900 2284.620 ;
        RECT 452.940 2284.300 453.260 2284.620 ;
        RECT 457.540 2284.300 457.860 2284.620 ;
        RECT 468.580 2284.300 468.900 2284.620 ;
        RECT 480.540 2284.300 480.860 2284.620 ;
        RECT 488.820 2284.300 489.140 2284.620 ;
        RECT 1018.740 2284.300 1019.060 2284.620 ;
        RECT 1019.660 2284.300 1019.980 2284.620 ;
        RECT 1027.020 2284.300 1027.340 2284.620 ;
        RECT 1037.140 2284.300 1037.460 2284.620 ;
        RECT 1046.340 2284.300 1046.660 2284.620 ;
        RECT 1054.620 2284.300 1054.940 2284.620 ;
        RECT 1061.980 2284.300 1062.300 2284.620 ;
        RECT 1066.580 2284.300 1066.900 2284.620 ;
        RECT 1089.580 2284.300 1089.900 2284.620 ;
        RECT 1096.020 2284.300 1096.340 2284.620 ;
        RECT 1109.820 2284.300 1110.140 2284.620 ;
        RECT 1116.260 2284.300 1116.580 2284.620 ;
        RECT 1119.020 2284.300 1119.340 2284.620 ;
        RECT 1130.980 2284.300 1131.300 2284.620 ;
        RECT 1136.500 2284.300 1136.820 2284.620 ;
        RECT 1144.780 2284.300 1145.100 2284.620 ;
        RECT 1148.460 2284.300 1148.780 2284.620 ;
        RECT 1153.980 2284.300 1154.300 2284.620 ;
        RECT 1165.020 2284.300 1165.340 2284.620 ;
        RECT 1171.460 2284.300 1171.780 2284.620 ;
        RECT 1178.820 2284.300 1179.140 2284.620 ;
        RECT 1183.420 2284.300 1183.740 2284.620 ;
        RECT 1188.940 2284.300 1189.260 2284.620 ;
        RECT 1198.140 2284.300 1198.460 2284.620 ;
        RECT 1580.860 2284.300 1581.180 2284.620 ;
        RECT 1595.580 2284.300 1595.900 2284.620 ;
        RECT 1601.100 2284.300 1601.420 2284.620 ;
        RECT 1666.420 2284.300 1666.740 2284.620 ;
        RECT 1671.940 2284.300 1672.260 2284.620 ;
        RECT 1683.900 2284.300 1684.220 2284.620 ;
        RECT 1695.860 2284.300 1696.180 2284.620 ;
        RECT 1701.380 2284.300 1701.700 2284.620 ;
        RECT 1754.740 2284.300 1755.060 2284.620 ;
        RECT 1759.340 2284.300 1759.660 2284.620 ;
        RECT 1776.820 2284.300 1777.140 2284.620 ;
        RECT 1783.260 2284.300 1783.580 2284.620 ;
        RECT 1788.780 2284.300 1789.100 2284.620 ;
        RECT 1794.300 2284.300 1794.620 2284.620 ;
        RECT 2234.060 2284.300 2234.380 2284.620 ;
        RECT 2242.340 2284.300 2242.660 2284.620 ;
        RECT 2251.540 2284.300 2251.860 2284.620 ;
        RECT 2263.500 2284.300 2263.820 2284.620 ;
        RECT 2265.340 2284.300 2265.660 2284.620 ;
        RECT 2268.100 2284.300 2268.420 2284.620 ;
        RECT 2280.980 2284.300 2281.300 2284.620 ;
        RECT 2286.500 2284.300 2286.820 2284.620 ;
        RECT 2304.900 2284.300 2305.220 2284.620 ;
        RECT 2315.940 2284.300 2316.260 2284.620 ;
        RECT 2322.380 2284.300 2322.700 2284.620 ;
        RECT 2327.900 2284.300 2328.220 2284.620 ;
        RECT 2333.420 2284.300 2333.740 2284.620 ;
        RECT 2339.860 2284.300 2340.180 2284.620 ;
        RECT 2350.900 2284.300 2351.220 2284.620 ;
        RECT 2357.340 2284.300 2357.660 2284.620 ;
        RECT 2368.380 2284.300 2368.700 2284.620 ;
        RECT 2374.820 2284.300 2375.140 2284.620 ;
      LAYER met4 ;
        RECT 668.215 2767.095 668.545 2767.425 ;
        RECT 1295.655 2767.095 1295.985 2767.425 ;
        RECT 1318.655 2767.095 1318.985 2767.425 ;
        RECT 1892.735 2767.095 1893.065 2767.425 ;
        RECT 1914.815 2767.095 1915.145 2767.425 ;
        RECT 2539.495 2767.095 2539.825 2767.425 ;
        RECT 2567.095 2767.095 2567.425 2767.425 ;
        RECT 668.230 2759.250 668.530 2767.095 ;
        RECT 667.865 2758.950 668.530 2759.250 ;
        RECT 394.025 2751.635 394.325 2756.235 ;
        RECT 400.265 2751.635 400.565 2756.235 ;
        RECT 406.505 2751.635 406.805 2756.235 ;
        RECT 412.745 2751.635 413.045 2756.235 ;
        RECT 418.985 2751.635 419.285 2756.235 ;
        RECT 425.225 2751.635 425.525 2756.235 ;
        RECT 431.465 2751.635 431.765 2756.235 ;
        RECT 437.705 2751.635 438.005 2756.235 ;
        RECT 443.945 2751.635 444.245 2756.235 ;
        RECT 450.185 2751.635 450.485 2756.235 ;
        RECT 456.425 2751.635 456.725 2756.235 ;
        RECT 462.665 2751.635 462.965 2756.235 ;
        RECT 468.905 2751.635 469.205 2756.235 ;
        RECT 475.145 2751.635 475.445 2756.235 ;
        RECT 481.385 2751.635 481.685 2756.235 ;
        RECT 487.625 2751.635 487.925 2756.235 ;
        RECT 493.865 2751.635 494.165 2756.235 ;
        RECT 500.105 2751.635 500.405 2756.235 ;
        RECT 506.345 2751.635 506.645 2756.235 ;
        RECT 512.585 2751.635 512.885 2756.235 ;
        RECT 518.825 2751.635 519.125 2756.235 ;
        RECT 525.065 2751.635 525.365 2756.235 ;
        RECT 531.305 2751.635 531.605 2756.235 ;
        RECT 537.545 2751.635 537.845 2756.235 ;
        RECT 543.785 2751.635 544.085 2756.235 ;
        RECT 550.025 2751.635 550.325 2756.235 ;
        RECT 556.265 2751.635 556.565 2756.235 ;
        RECT 562.505 2751.635 562.805 2756.235 ;
        RECT 568.745 2751.635 569.045 2756.235 ;
        RECT 574.985 2751.635 575.285 2756.235 ;
        RECT 581.225 2751.635 581.525 2756.235 ;
        RECT 587.465 2751.635 587.765 2756.235 ;
        RECT 642.890 2755.850 643.190 2756.235 ;
        RECT 646.135 2755.850 646.465 2755.865 ;
        RECT 642.890 2755.550 646.465 2755.850 ;
        RECT 642.890 2751.635 643.190 2755.550 ;
        RECT 646.135 2755.535 646.465 2755.550 ;
        RECT 664.535 2755.850 664.865 2755.865 ;
        RECT 667.865 2755.850 668.165 2758.950 ;
        RECT 664.535 2755.550 668.165 2755.850 ;
        RECT 664.535 2755.535 664.865 2755.550 ;
        RECT 667.865 2751.635 668.165 2755.550 ;
        RECT 1044.025 2751.635 1044.325 2756.235 ;
        RECT 1050.265 2751.635 1050.565 2756.235 ;
        RECT 1056.505 2751.635 1056.805 2756.235 ;
        RECT 1062.745 2751.635 1063.045 2756.235 ;
        RECT 1068.985 2751.635 1069.285 2756.235 ;
        RECT 1075.225 2751.635 1075.525 2756.235 ;
        RECT 1081.465 2751.635 1081.765 2756.235 ;
        RECT 1087.705 2751.635 1088.005 2756.235 ;
        RECT 1093.945 2751.635 1094.245 2756.235 ;
        RECT 1100.185 2751.635 1100.485 2756.235 ;
        RECT 1106.425 2751.635 1106.725 2756.235 ;
        RECT 1112.665 2751.635 1112.965 2756.235 ;
        RECT 1118.905 2751.635 1119.205 2756.235 ;
        RECT 1125.145 2751.635 1125.445 2756.235 ;
        RECT 1131.385 2751.635 1131.685 2756.235 ;
        RECT 1137.625 2751.635 1137.925 2756.235 ;
        RECT 1143.865 2751.635 1144.165 2756.235 ;
        RECT 1150.105 2751.635 1150.405 2756.235 ;
        RECT 1156.345 2751.635 1156.645 2756.235 ;
        RECT 1162.585 2751.635 1162.885 2756.235 ;
        RECT 1168.825 2751.635 1169.125 2756.235 ;
        RECT 1175.065 2751.635 1175.365 2756.235 ;
        RECT 1181.305 2751.635 1181.605 2756.235 ;
        RECT 1187.545 2751.635 1187.845 2756.235 ;
        RECT 1193.785 2751.635 1194.085 2756.235 ;
        RECT 1200.025 2751.635 1200.325 2756.235 ;
        RECT 1206.265 2751.635 1206.565 2756.235 ;
        RECT 1212.505 2751.635 1212.805 2756.235 ;
        RECT 1218.745 2751.635 1219.045 2756.235 ;
        RECT 1224.985 2751.635 1225.285 2756.235 ;
        RECT 1231.225 2751.635 1231.525 2756.235 ;
        RECT 1237.465 2751.635 1237.765 2756.235 ;
        RECT 1292.890 2755.850 1293.190 2756.235 ;
        RECT 1295.670 2755.850 1295.970 2767.095 ;
        RECT 1292.890 2755.550 1295.970 2755.850 ;
        RECT 1317.865 2755.850 1318.165 2756.235 ;
        RECT 1318.670 2755.850 1318.970 2767.095 ;
        RECT 1892.750 2756.235 1893.050 2767.095 ;
        RECT 1317.865 2755.550 1318.970 2755.850 ;
        RECT 1292.890 2751.635 1293.190 2755.550 ;
        RECT 1317.865 2751.635 1318.165 2755.550 ;
        RECT 1644.025 2751.635 1644.325 2756.235 ;
        RECT 1650.265 2751.635 1650.565 2756.235 ;
        RECT 1656.505 2751.635 1656.805 2756.235 ;
        RECT 1662.745 2751.635 1663.045 2756.235 ;
        RECT 1668.985 2751.635 1669.285 2756.235 ;
        RECT 1675.225 2751.635 1675.525 2756.235 ;
        RECT 1681.465 2751.635 1681.765 2756.235 ;
        RECT 1687.705 2751.635 1688.005 2756.235 ;
        RECT 1693.945 2751.635 1694.245 2756.235 ;
        RECT 1700.185 2751.635 1700.485 2756.235 ;
        RECT 1706.425 2751.635 1706.725 2756.235 ;
        RECT 1712.665 2751.635 1712.965 2756.235 ;
        RECT 1718.905 2751.635 1719.205 2756.235 ;
        RECT 1725.145 2751.635 1725.445 2756.235 ;
        RECT 1731.385 2751.635 1731.685 2756.235 ;
        RECT 1737.625 2751.635 1737.925 2756.235 ;
        RECT 1743.865 2751.635 1744.165 2756.235 ;
        RECT 1750.105 2751.635 1750.405 2756.235 ;
        RECT 1756.345 2751.635 1756.645 2756.235 ;
        RECT 1762.585 2751.635 1762.885 2756.235 ;
        RECT 1768.825 2751.635 1769.125 2756.235 ;
        RECT 1775.065 2751.635 1775.365 2756.235 ;
        RECT 1781.305 2751.635 1781.605 2756.235 ;
        RECT 1787.545 2751.635 1787.845 2756.235 ;
        RECT 1793.785 2751.635 1794.085 2756.235 ;
        RECT 1800.025 2751.635 1800.325 2756.235 ;
        RECT 1806.265 2751.635 1806.565 2756.235 ;
        RECT 1812.505 2751.635 1812.805 2756.235 ;
        RECT 1818.745 2751.635 1819.045 2756.235 ;
        RECT 1824.985 2751.635 1825.285 2756.235 ;
        RECT 1831.225 2751.635 1831.525 2756.235 ;
        RECT 1837.465 2751.635 1837.765 2756.235 ;
        RECT 1892.750 2755.550 1893.190 2756.235 ;
        RECT 1914.830 2755.850 1915.130 2767.095 ;
        RECT 1917.865 2755.850 1918.165 2756.235 ;
        RECT 1914.830 2755.550 1918.165 2755.850 ;
        RECT 1892.890 2751.635 1893.190 2755.550 ;
        RECT 1917.865 2751.635 1918.165 2755.550 ;
        RECT 2294.025 2751.635 2294.325 2756.235 ;
        RECT 2300.265 2751.635 2300.565 2756.235 ;
        RECT 2306.505 2751.635 2306.805 2756.235 ;
        RECT 2312.745 2751.635 2313.045 2756.235 ;
        RECT 2318.985 2751.635 2319.285 2756.235 ;
        RECT 2325.225 2751.635 2325.525 2756.235 ;
        RECT 2331.465 2751.635 2331.765 2756.235 ;
        RECT 2337.705 2751.635 2338.005 2756.235 ;
        RECT 2343.945 2751.635 2344.245 2756.235 ;
        RECT 2350.185 2751.635 2350.485 2756.235 ;
        RECT 2356.425 2751.635 2356.725 2756.235 ;
        RECT 2362.665 2751.635 2362.965 2756.235 ;
        RECT 2368.905 2751.635 2369.205 2756.235 ;
        RECT 2375.145 2751.635 2375.445 2756.235 ;
        RECT 2381.385 2751.635 2381.685 2756.235 ;
        RECT 2387.625 2751.635 2387.925 2756.235 ;
        RECT 2393.865 2751.635 2394.165 2756.235 ;
        RECT 2400.105 2751.635 2400.405 2756.235 ;
        RECT 2406.345 2751.635 2406.645 2756.235 ;
        RECT 2412.585 2751.635 2412.885 2756.235 ;
        RECT 2418.825 2751.635 2419.125 2756.235 ;
        RECT 2425.065 2751.635 2425.365 2756.235 ;
        RECT 2431.305 2751.635 2431.605 2756.235 ;
        RECT 2437.545 2751.635 2437.845 2756.235 ;
        RECT 2443.785 2751.635 2444.085 2756.235 ;
        RECT 2450.025 2751.635 2450.325 2756.235 ;
        RECT 2456.265 2751.635 2456.565 2756.235 ;
        RECT 2462.505 2751.635 2462.805 2756.235 ;
        RECT 2468.745 2751.635 2469.045 2756.235 ;
        RECT 2474.985 2751.635 2475.285 2756.235 ;
        RECT 2481.225 2751.635 2481.525 2756.235 ;
        RECT 2487.465 2751.635 2487.765 2756.235 ;
        RECT 2539.510 2755.850 2539.810 2767.095 ;
        RECT 2542.890 2755.850 2543.190 2756.235 ;
        RECT 2539.510 2755.550 2543.190 2755.850 ;
        RECT 2567.110 2755.850 2567.410 2767.095 ;
        RECT 2567.865 2755.850 2568.165 2756.235 ;
        RECT 2567.110 2755.550 2571.090 2755.850 ;
        RECT 2542.890 2751.635 2543.190 2755.550 ;
        RECT 2567.865 2751.635 2568.165 2755.550 ;
        RECT 2570.790 2753.825 2571.090 2755.550 ;
        RECT 2570.775 2753.495 2571.105 2753.825 ;
      LAYER met4 ;
        RECT 305.000 2305.000 681.480 2751.235 ;
        RECT 955.000 2305.000 1331.480 2751.235 ;
        RECT 1555.000 2305.000 1931.480 2751.235 ;
        RECT 2205.000 2305.000 2581.480 2751.235 ;
      LAYER met4 ;
        RECT 334.010 2296.850 334.310 2304.600 ;
        RECT 339.850 2296.850 340.150 2304.600 ;
        RECT 345.690 2301.950 345.990 2304.600 ;
        RECT 351.530 2301.950 351.830 2304.600 ;
        RECT 345.690 2301.650 349.290 2301.950 ;
        RECT 345.690 2300.000 345.990 2301.650 ;
        RECT 334.010 2296.550 334.570 2296.850 ;
        RECT 310.020 2215.000 313.020 2285.000 ;
        RECT 328.020 2215.000 331.020 2285.000 ;
        RECT 334.270 2284.625 334.570 2296.550 ;
        RECT 339.790 2296.550 340.150 2296.850 ;
        RECT 339.790 2284.625 340.090 2296.550 ;
        RECT 348.990 2284.625 349.290 2301.650 ;
        RECT 350.830 2301.650 351.830 2301.950 ;
        RECT 350.830 2285.305 351.130 2301.650 ;
        RECT 351.530 2300.000 351.830 2301.650 ;
        RECT 357.370 2296.850 357.670 2304.600 ;
        RECT 357.270 2296.550 357.670 2296.850 ;
        RECT 363.210 2296.850 363.510 2304.600 ;
        RECT 363.830 2301.950 364.130 2304.600 ;
        RECT 363.830 2301.650 364.930 2301.950 ;
        RECT 363.830 2300.000 364.130 2301.650 ;
        RECT 363.210 2296.550 364.010 2296.850 ;
        RECT 350.815 2284.975 351.145 2285.305 ;
        RECT 357.270 2284.625 357.570 2296.550 ;
        RECT 363.710 2288.705 364.010 2296.550 ;
        RECT 363.695 2288.375 364.025 2288.705 ;
        RECT 364.630 2285.985 364.930 2301.650 ;
        RECT 369.050 2296.850 369.350 2304.600 ;
        RECT 369.670 2303.650 369.970 2304.600 ;
        RECT 369.670 2303.350 371.370 2303.650 ;
        RECT 369.670 2300.000 369.970 2303.350 ;
        RECT 369.050 2296.550 369.530 2296.850 ;
        RECT 369.230 2290.745 369.530 2296.550 ;
        RECT 369.215 2290.415 369.545 2290.745 ;
        RECT 371.070 2287.345 371.370 2303.350 ;
        RECT 374.890 2296.850 375.190 2304.600 ;
        RECT 374.750 2296.550 375.190 2296.850 ;
        RECT 375.510 2296.850 375.810 2304.600 ;
        RECT 380.730 2303.650 381.030 2304.600 ;
        RECT 379.350 2303.350 381.030 2303.650 ;
        RECT 375.510 2296.550 375.970 2296.850 ;
        RECT 374.750 2290.745 375.050 2296.550 ;
        RECT 374.735 2290.415 375.065 2290.745 ;
        RECT 371.055 2287.015 371.385 2287.345 ;
        RECT 364.615 2285.655 364.945 2285.985 ;
        RECT 375.670 2285.305 375.970 2296.550 ;
        RECT 379.350 2288.025 379.650 2303.350 ;
        RECT 380.730 2300.000 381.030 2303.350 ;
        RECT 381.350 2296.850 381.650 2304.600 ;
        RECT 386.570 2297.545 386.870 2304.600 ;
        RECT 386.555 2297.215 386.885 2297.545 ;
        RECT 387.190 2296.850 387.490 2304.600 ;
        RECT 392.410 2296.850 392.710 2304.600 ;
        RECT 393.030 2301.950 393.330 2304.600 ;
        RECT 398.250 2303.650 398.550 2304.600 ;
        RECT 396.830 2303.350 398.550 2303.650 ;
        RECT 393.030 2300.000 393.450 2301.950 ;
        RECT 381.190 2296.550 381.650 2296.850 ;
        RECT 386.710 2296.550 387.490 2296.850 ;
        RECT 392.230 2296.550 392.710 2296.850 ;
        RECT 379.335 2287.695 379.665 2288.025 ;
        RECT 381.190 2287.345 381.490 2296.550 ;
        RECT 381.175 2287.015 381.505 2287.345 ;
        RECT 386.710 2285.985 387.010 2296.550 ;
        RECT 392.230 2289.385 392.530 2296.550 ;
        RECT 392.215 2289.055 392.545 2289.385 ;
        RECT 386.695 2285.655 387.025 2285.985 ;
        RECT 393.150 2285.305 393.450 2300.000 ;
        RECT 396.830 2290.745 397.130 2303.350 ;
        RECT 398.250 2300.000 398.550 2303.350 ;
        RECT 398.870 2296.850 399.170 2304.600 ;
        RECT 404.090 2301.950 404.390 2304.600 ;
        RECT 398.670 2296.550 399.170 2296.850 ;
        RECT 403.270 2301.650 404.390 2301.950 ;
        RECT 396.815 2290.415 397.145 2290.745 ;
        RECT 334.255 2284.295 334.585 2284.625 ;
        RECT 339.775 2284.295 340.105 2284.625 ;
        RECT 348.975 2284.295 349.305 2284.625 ;
        RECT 357.255 2284.295 357.585 2284.625 ;
        RECT 364.020 2215.000 367.020 2285.000 ;
        RECT 375.655 2284.975 375.985 2285.305 ;
        RECT 382.020 2215.000 385.020 2285.000 ;
        RECT 393.135 2284.975 393.465 2285.305 ;
        RECT 398.670 2284.625 398.970 2296.550 ;
        RECT 403.270 2290.065 403.570 2301.650 ;
        RECT 404.090 2300.000 404.390 2301.650 ;
        RECT 404.710 2296.850 405.010 2304.600 ;
        RECT 409.930 2296.850 410.230 2304.600 ;
        RECT 404.190 2296.550 405.010 2296.850 ;
        RECT 409.710 2296.550 410.230 2296.850 ;
        RECT 410.550 2296.850 410.850 2304.600 ;
        RECT 415.770 2303.650 416.070 2304.600 ;
        RECT 414.310 2303.350 416.070 2303.650 ;
        RECT 410.550 2296.550 410.930 2296.850 ;
        RECT 403.255 2289.735 403.585 2290.065 ;
        RECT 398.655 2284.295 398.985 2284.625 ;
        RECT 400.020 2215.000 403.020 2285.000 ;
        RECT 404.190 2284.625 404.490 2296.550 ;
        RECT 409.710 2290.745 410.010 2296.550 ;
        RECT 409.695 2290.415 410.025 2290.745 ;
        RECT 410.630 2284.625 410.930 2296.550 ;
        RECT 414.310 2290.745 414.610 2303.350 ;
        RECT 415.770 2300.000 416.070 2303.350 ;
        RECT 416.390 2296.850 416.690 2304.600 ;
        RECT 421.610 2301.950 421.910 2304.600 ;
        RECT 416.150 2296.550 416.690 2296.850 ;
        RECT 420.750 2301.650 421.910 2301.950 ;
        RECT 414.295 2290.415 414.625 2290.745 ;
        RECT 416.150 2284.625 416.450 2296.550 ;
        RECT 420.750 2290.745 421.050 2301.650 ;
        RECT 421.610 2300.000 421.910 2301.650 ;
        RECT 422.230 2296.850 422.530 2304.600 ;
        RECT 427.450 2296.850 427.750 2304.600 ;
        RECT 421.670 2296.550 422.530 2296.850 ;
        RECT 427.190 2296.550 427.750 2296.850 ;
        RECT 428.070 2296.850 428.370 2304.600 ;
        RECT 433.290 2303.650 433.590 2304.600 ;
        RECT 431.790 2303.350 433.590 2303.650 ;
        RECT 428.070 2296.550 428.410 2296.850 ;
        RECT 420.735 2290.415 421.065 2290.745 ;
        RECT 421.670 2284.625 421.970 2296.550 ;
        RECT 427.190 2290.745 427.490 2296.550 ;
        RECT 427.175 2290.415 427.505 2290.745 ;
        RECT 428.110 2284.625 428.410 2296.550 ;
        RECT 431.790 2290.745 432.090 2303.350 ;
        RECT 433.290 2300.000 433.590 2303.350 ;
        RECT 433.910 2296.850 434.210 2304.600 ;
        RECT 433.630 2296.550 434.210 2296.850 ;
        RECT 439.130 2296.850 439.430 2304.600 ;
        RECT 439.750 2296.850 440.050 2304.600 ;
        RECT 444.970 2296.850 445.270 2304.600 ;
        RECT 439.130 2296.550 439.450 2296.850 ;
        RECT 439.750 2296.550 440.370 2296.850 ;
        RECT 431.775 2290.415 432.105 2290.745 ;
        RECT 433.630 2284.625 433.930 2296.550 ;
        RECT 439.150 2290.745 439.450 2296.550 ;
        RECT 439.135 2290.415 439.465 2290.745 ;
        RECT 440.070 2284.625 440.370 2296.550 ;
        RECT 444.670 2296.550 445.270 2296.850 ;
        RECT 444.670 2290.745 444.970 2296.550 ;
        RECT 444.655 2290.415 444.985 2290.745 ;
        RECT 445.590 2284.625 445.890 2304.600 ;
        RECT 450.810 2296.850 451.110 2304.600 ;
        RECT 451.430 2301.950 451.730 2304.600 ;
        RECT 451.430 2301.650 453.250 2301.950 ;
        RECT 451.430 2300.000 451.730 2301.650 ;
        RECT 450.810 2296.550 451.410 2296.850 ;
        RECT 451.110 2290.745 451.410 2296.550 ;
        RECT 451.095 2290.415 451.425 2290.745 ;
        RECT 452.950 2284.625 453.250 2301.650 ;
        RECT 456.650 2296.850 456.950 2304.600 ;
        RECT 456.630 2296.550 456.950 2296.850 ;
        RECT 457.270 2296.850 457.570 2304.600 ;
        RECT 462.490 2296.850 462.790 2304.600 ;
        RECT 463.110 2301.950 463.410 2304.600 ;
        RECT 468.330 2301.950 468.630 2304.600 ;
        RECT 463.110 2301.650 466.130 2301.950 ;
        RECT 463.110 2300.000 463.410 2301.650 ;
        RECT 457.270 2296.550 457.850 2296.850 ;
        RECT 456.630 2290.745 456.930 2296.550 ;
        RECT 456.615 2290.415 456.945 2290.745 ;
        RECT 457.550 2284.625 457.850 2296.550 ;
        RECT 462.150 2296.550 462.790 2296.850 ;
        RECT 462.150 2290.745 462.450 2296.550 ;
        RECT 462.135 2290.415 462.465 2290.745 ;
        RECT 465.830 2285.305 466.130 2301.650 ;
        RECT 467.670 2301.650 468.630 2301.950 ;
        RECT 467.670 2290.745 467.970 2301.650 ;
        RECT 468.330 2300.000 468.630 2301.650 ;
        RECT 468.950 2296.850 469.250 2304.600 ;
        RECT 474.170 2296.850 474.470 2304.600 ;
        RECT 468.590 2296.550 469.250 2296.850 ;
        RECT 474.110 2296.550 474.470 2296.850 ;
        RECT 474.790 2296.850 475.090 2304.600 ;
        RECT 480.010 2303.650 480.310 2304.600 ;
        RECT 478.710 2303.350 480.310 2303.650 ;
        RECT 474.790 2296.550 475.330 2296.850 ;
        RECT 467.655 2290.415 467.985 2290.745 ;
        RECT 465.815 2284.975 466.145 2285.305 ;
        RECT 468.590 2284.625 468.890 2296.550 ;
        RECT 474.110 2290.745 474.410 2296.550 ;
        RECT 474.095 2290.415 474.425 2290.745 ;
        RECT 475.030 2285.985 475.330 2296.550 ;
        RECT 478.710 2290.745 479.010 2303.350 ;
        RECT 480.010 2300.000 480.310 2303.350 ;
        RECT 480.630 2296.850 480.930 2304.600 ;
        RECT 480.550 2296.550 480.930 2296.850 ;
        RECT 485.850 2296.850 486.150 2304.600 ;
        RECT 486.470 2301.950 486.770 2304.600 ;
        RECT 486.470 2301.650 489.130 2301.950 ;
        RECT 486.470 2300.000 486.770 2301.650 ;
        RECT 485.850 2296.550 486.370 2296.850 ;
        RECT 478.695 2290.415 479.025 2290.745 ;
        RECT 475.015 2285.655 475.345 2285.985 ;
        RECT 480.550 2284.625 480.850 2296.550 ;
        RECT 486.070 2290.745 486.370 2296.550 ;
        RECT 486.055 2290.415 486.385 2290.745 ;
        RECT 488.830 2284.625 489.130 2301.650 ;
        RECT 491.690 2296.850 491.990 2304.600 ;
        RECT 491.590 2296.550 491.990 2296.850 ;
        RECT 492.310 2296.850 492.610 2304.600 ;
        RECT 497.530 2296.850 497.830 2304.600 ;
        RECT 498.150 2301.950 498.450 2304.600 ;
        RECT 503.370 2301.950 503.670 2304.600 ;
        RECT 498.150 2301.650 501.090 2301.950 ;
        RECT 498.150 2300.000 498.450 2301.650 ;
        RECT 492.310 2296.550 492.810 2296.850 ;
        RECT 491.590 2290.745 491.890 2296.550 ;
        RECT 491.575 2290.415 491.905 2290.745 ;
        RECT 492.510 2285.985 492.810 2296.550 ;
        RECT 497.110 2296.550 497.830 2296.850 ;
        RECT 497.110 2290.745 497.410 2296.550 ;
        RECT 500.790 2290.745 501.090 2301.650 ;
        RECT 502.630 2301.650 503.670 2301.950 ;
        RECT 497.095 2290.415 497.425 2290.745 ;
        RECT 500.775 2290.415 501.105 2290.745 ;
        RECT 502.630 2290.065 502.930 2301.650 ;
        RECT 503.370 2300.000 503.670 2301.650 ;
        RECT 503.990 2301.950 504.290 2304.600 ;
        RECT 503.990 2301.650 507.530 2301.950 ;
        RECT 503.990 2300.000 504.290 2301.650 ;
        RECT 507.230 2290.065 507.530 2301.650 ;
        RECT 509.210 2296.850 509.510 2304.600 ;
        RECT 509.070 2296.550 509.510 2296.850 ;
        RECT 509.830 2296.850 510.130 2304.600 ;
        RECT 515.050 2303.650 515.350 2304.600 ;
        RECT 513.670 2303.350 515.350 2303.650 ;
        RECT 509.830 2296.550 510.290 2296.850 ;
        RECT 502.615 2289.735 502.945 2290.065 ;
        RECT 507.215 2289.735 507.545 2290.065 ;
        RECT 509.070 2289.385 509.370 2296.550 ;
        RECT 509.990 2290.745 510.290 2296.550 ;
        RECT 513.670 2290.745 513.970 2303.350 ;
        RECT 515.050 2300.000 515.350 2303.350 ;
        RECT 515.670 2296.850 515.970 2304.600 ;
        RECT 515.510 2296.550 515.970 2296.850 ;
        RECT 520.890 2296.850 521.190 2304.600 ;
        RECT 521.510 2301.950 521.810 2304.600 ;
        RECT 521.510 2301.650 524.090 2301.950 ;
        RECT 521.510 2300.000 521.810 2301.650 ;
        RECT 520.890 2296.550 521.330 2296.850 ;
        RECT 515.510 2290.745 515.810 2296.550 ;
        RECT 521.030 2290.745 521.330 2296.550 ;
        RECT 523.790 2290.745 524.090 2301.650 ;
        RECT 526.730 2296.850 527.030 2304.600 ;
        RECT 526.550 2296.550 527.030 2296.850 ;
        RECT 527.350 2296.850 527.650 2304.600 ;
        RECT 532.570 2296.850 532.870 2304.600 ;
        RECT 533.190 2301.950 533.490 2304.600 ;
        RECT 533.190 2301.650 536.050 2301.950 ;
        RECT 533.190 2300.000 533.490 2301.650 ;
        RECT 527.350 2296.550 527.770 2296.850 ;
        RECT 526.550 2290.745 526.850 2296.550 ;
        RECT 527.470 2290.745 527.770 2296.550 ;
        RECT 532.070 2296.550 532.870 2296.850 ;
        RECT 509.975 2290.415 510.305 2290.745 ;
        RECT 513.655 2290.415 513.985 2290.745 ;
        RECT 515.495 2290.415 515.825 2290.745 ;
        RECT 521.015 2290.415 521.345 2290.745 ;
        RECT 523.775 2290.415 524.105 2290.745 ;
        RECT 526.535 2290.415 526.865 2290.745 ;
        RECT 527.455 2290.415 527.785 2290.745 ;
        RECT 532.070 2290.065 532.370 2296.550 ;
        RECT 535.750 2290.745 536.050 2301.650 ;
        RECT 538.410 2296.850 538.710 2304.600 ;
        RECT 539.030 2301.950 539.330 2304.600 ;
        RECT 539.030 2301.650 542.490 2301.950 ;
        RECT 539.030 2300.000 539.330 2301.650 ;
        RECT 538.410 2296.550 538.810 2296.850 ;
        RECT 535.735 2290.415 536.065 2290.745 ;
        RECT 538.510 2290.065 538.810 2296.550 ;
        RECT 542.190 2290.065 542.490 2301.650 ;
        RECT 544.250 2296.850 544.550 2304.600 ;
        RECT 544.870 2301.950 545.170 2304.600 ;
        RECT 544.870 2300.000 545.250 2301.950 ;
        RECT 544.030 2296.550 544.550 2296.850 ;
        RECT 544.030 2290.745 544.330 2296.550 ;
        RECT 544.950 2290.745 545.250 2300.000 ;
        RECT 984.010 2296.850 984.310 2304.600 ;
        RECT 989.850 2301.950 990.150 2304.600 ;
        RECT 983.790 2296.550 984.310 2296.850 ;
        RECT 987.470 2301.650 990.150 2301.950 ;
        RECT 544.015 2290.415 544.345 2290.745 ;
        RECT 544.935 2290.415 545.265 2290.745 ;
        RECT 532.055 2289.735 532.385 2290.065 ;
        RECT 538.495 2289.735 538.825 2290.065 ;
        RECT 542.175 2289.735 542.505 2290.065 ;
        RECT 509.055 2289.055 509.385 2289.385 ;
        RECT 983.790 2288.025 984.090 2296.550 ;
        RECT 987.470 2290.065 987.770 2301.650 ;
        RECT 989.850 2300.000 990.150 2301.650 ;
        RECT 995.690 2296.850 995.990 2304.600 ;
        RECT 1001.530 2296.850 1001.830 2304.600 ;
        RECT 995.690 2296.550 996.050 2296.850 ;
        RECT 995.750 2290.065 996.050 2296.550 ;
        RECT 1001.270 2296.550 1001.830 2296.850 ;
        RECT 1007.370 2296.850 1007.670 2304.600 ;
        RECT 1013.210 2301.950 1013.510 2304.600 ;
        RECT 1012.310 2301.650 1013.510 2301.950 ;
        RECT 1007.370 2296.550 1008.010 2296.850 ;
        RECT 1001.270 2290.745 1001.570 2296.550 ;
        RECT 1001.255 2290.415 1001.585 2290.745 ;
        RECT 987.455 2289.735 987.785 2290.065 ;
        RECT 995.735 2289.735 996.065 2290.065 ;
        RECT 1007.710 2288.705 1008.010 2296.550 ;
        RECT 1007.695 2288.375 1008.025 2288.705 ;
        RECT 983.775 2287.695 984.105 2288.025 ;
        RECT 1012.310 2285.985 1012.610 2301.650 ;
        RECT 1013.210 2300.000 1013.510 2301.650 ;
        RECT 1013.830 2296.850 1014.130 2304.600 ;
        RECT 1019.050 2296.850 1019.350 2304.600 ;
        RECT 1013.230 2296.550 1014.130 2296.850 ;
        RECT 1018.750 2296.550 1019.350 2296.850 ;
        RECT 1013.230 2285.985 1013.530 2296.550 ;
        RECT 492.495 2285.655 492.825 2285.985 ;
        RECT 1012.295 2285.655 1012.625 2285.985 ;
        RECT 1013.215 2285.655 1013.545 2285.985 ;
        RECT 404.175 2284.295 404.505 2284.625 ;
        RECT 410.615 2284.295 410.945 2284.625 ;
        RECT 416.135 2284.295 416.465 2284.625 ;
        RECT 421.655 2284.295 421.985 2284.625 ;
        RECT 428.095 2284.295 428.425 2284.625 ;
        RECT 433.615 2284.295 433.945 2284.625 ;
        RECT 440.055 2284.295 440.385 2284.625 ;
        RECT 445.575 2284.295 445.905 2284.625 ;
        RECT 452.935 2284.295 453.265 2284.625 ;
        RECT 457.535 2284.295 457.865 2284.625 ;
        RECT 468.575 2284.295 468.905 2284.625 ;
        RECT 480.535 2284.295 480.865 2284.625 ;
        RECT 488.815 2284.295 489.145 2284.625 ;
        RECT 490.020 2215.000 493.020 2285.000 ;
        RECT 508.020 2215.000 511.020 2285.000 ;
        RECT 544.020 2215.000 547.020 2285.000 ;
        RECT 562.020 2215.000 565.020 2285.000 ;
        RECT 580.020 2215.000 583.020 2285.000 ;
        RECT 670.020 2215.000 673.020 2285.000 ;
        RECT 688.020 2215.000 691.020 2285.000 ;
        RECT 940.020 2215.000 943.020 2285.000 ;
        RECT 1018.750 2284.625 1019.050 2296.550 ;
        RECT 1019.670 2284.625 1019.970 2304.600 ;
        RECT 1024.890 2296.850 1025.190 2304.600 ;
        RECT 1025.510 2301.950 1025.810 2304.600 ;
        RECT 1025.510 2301.650 1027.330 2301.950 ;
        RECT 1025.510 2300.000 1025.810 2301.650 ;
        RECT 1024.890 2296.550 1025.490 2296.850 ;
        RECT 1025.190 2285.305 1025.490 2296.550 ;
        RECT 1025.175 2284.975 1025.505 2285.305 ;
        RECT 1027.030 2284.625 1027.330 2301.650 ;
        RECT 1030.730 2296.850 1031.030 2304.600 ;
        RECT 1030.710 2296.550 1031.030 2296.850 ;
        RECT 1031.350 2296.850 1031.650 2304.600 ;
        RECT 1036.570 2303.650 1036.870 2304.600 ;
        RECT 1035.310 2303.350 1036.870 2303.650 ;
        RECT 1031.350 2296.550 1031.930 2296.850 ;
        RECT 1030.710 2286.665 1031.010 2296.550 ;
        RECT 1030.695 2286.335 1031.025 2286.665 ;
        RECT 1031.630 2285.985 1031.930 2296.550 ;
        RECT 1035.310 2290.065 1035.610 2303.350 ;
        RECT 1036.570 2300.000 1036.870 2303.350 ;
        RECT 1037.190 2296.850 1037.490 2304.600 ;
        RECT 1037.150 2296.550 1037.490 2296.850 ;
        RECT 1042.410 2296.850 1042.710 2304.600 ;
        RECT 1043.030 2301.950 1043.330 2304.600 ;
        RECT 1043.030 2301.650 1046.650 2301.950 ;
        RECT 1043.030 2300.000 1043.330 2301.650 ;
        RECT 1042.410 2296.550 1042.970 2296.850 ;
        RECT 1035.295 2289.735 1035.625 2290.065 ;
        RECT 1031.615 2285.655 1031.945 2285.985 ;
        RECT 1018.735 2284.295 1019.065 2284.625 ;
        RECT 1019.655 2284.295 1019.985 2284.625 ;
        RECT 1027.015 2284.295 1027.345 2284.625 ;
        RECT 1030.020 2215.000 1033.020 2285.000 ;
        RECT 1037.150 2284.625 1037.450 2296.550 ;
        RECT 1042.670 2287.345 1042.970 2296.550 ;
        RECT 1042.655 2287.015 1042.985 2287.345 ;
        RECT 1046.350 2284.625 1046.650 2301.650 ;
        RECT 1048.250 2296.850 1048.550 2304.600 ;
        RECT 1048.190 2296.550 1048.550 2296.850 ;
        RECT 1048.870 2296.850 1049.170 2304.600 ;
        RECT 1054.090 2303.650 1054.390 2304.600 ;
        RECT 1052.790 2303.350 1054.390 2303.650 ;
        RECT 1048.870 2296.550 1049.410 2296.850 ;
        RECT 1048.190 2288.705 1048.490 2296.550 ;
        RECT 1048.175 2288.375 1048.505 2288.705 ;
        RECT 1049.110 2285.985 1049.410 2296.550 ;
        RECT 1052.790 2290.745 1053.090 2303.350 ;
        RECT 1054.090 2300.000 1054.390 2303.350 ;
        RECT 1054.710 2296.850 1055.010 2304.600 ;
        RECT 1054.630 2296.550 1055.010 2296.850 ;
        RECT 1059.930 2296.850 1060.230 2304.600 ;
        RECT 1060.550 2301.950 1060.850 2304.600 ;
        RECT 1060.550 2301.650 1062.290 2301.950 ;
        RECT 1060.550 2300.000 1060.850 2301.650 ;
        RECT 1059.930 2296.550 1060.450 2296.850 ;
        RECT 1052.775 2290.415 1053.105 2290.745 ;
        RECT 1049.095 2285.655 1049.425 2285.985 ;
        RECT 1037.135 2284.295 1037.465 2284.625 ;
        RECT 1046.335 2284.295 1046.665 2284.625 ;
        RECT 1048.020 2215.000 1051.020 2285.000 ;
        RECT 1054.630 2284.625 1054.930 2296.550 ;
        RECT 1060.150 2290.745 1060.450 2296.550 ;
        RECT 1060.135 2290.415 1060.465 2290.745 ;
        RECT 1061.990 2284.625 1062.290 2301.650 ;
        RECT 1065.770 2296.850 1066.070 2304.600 ;
        RECT 1065.670 2296.550 1066.070 2296.850 ;
        RECT 1066.390 2296.850 1066.690 2304.600 ;
        RECT 1071.610 2303.650 1071.910 2304.600 ;
        RECT 1070.270 2303.350 1071.910 2303.650 ;
        RECT 1066.390 2296.550 1066.890 2296.850 ;
        RECT 1065.670 2290.745 1065.970 2296.550 ;
        RECT 1065.655 2290.415 1065.985 2290.745 ;
        RECT 1066.590 2284.625 1066.890 2296.550 ;
        RECT 1070.270 2290.745 1070.570 2303.350 ;
        RECT 1071.610 2300.000 1071.910 2303.350 ;
        RECT 1072.230 2296.850 1072.530 2304.600 ;
        RECT 1077.450 2301.950 1077.750 2304.600 ;
        RECT 1072.110 2296.550 1072.530 2296.850 ;
        RECT 1076.710 2301.650 1077.750 2301.950 ;
        RECT 1070.255 2290.415 1070.585 2290.745 ;
        RECT 1072.110 2285.985 1072.410 2296.550 ;
        RECT 1076.710 2290.745 1077.010 2301.650 ;
        RECT 1077.450 2300.000 1077.750 2301.650 ;
        RECT 1078.070 2301.950 1078.370 2304.600 ;
        RECT 1078.070 2301.650 1081.610 2301.950 ;
        RECT 1078.070 2300.000 1078.370 2301.650 ;
        RECT 1076.695 2290.415 1077.025 2290.745 ;
        RECT 1081.310 2287.345 1081.610 2301.650 ;
        RECT 1083.290 2296.850 1083.590 2304.600 ;
        RECT 1083.150 2296.550 1083.590 2296.850 ;
        RECT 1083.910 2296.850 1084.210 2304.600 ;
        RECT 1089.130 2303.650 1089.430 2304.600 ;
        RECT 1087.750 2303.350 1089.430 2303.650 ;
        RECT 1083.910 2296.550 1084.370 2296.850 ;
        RECT 1083.150 2290.745 1083.450 2296.550 ;
        RECT 1083.135 2290.415 1083.465 2290.745 ;
        RECT 1081.295 2287.015 1081.625 2287.345 ;
        RECT 1084.070 2285.985 1084.370 2296.550 ;
        RECT 1087.750 2290.745 1088.050 2303.350 ;
        RECT 1089.130 2300.000 1089.430 2303.350 ;
        RECT 1089.750 2296.850 1090.050 2304.600 ;
        RECT 1094.970 2301.950 1095.270 2304.600 ;
        RECT 1089.590 2296.550 1090.050 2296.850 ;
        RECT 1094.190 2301.650 1095.270 2301.950 ;
        RECT 1087.735 2290.415 1088.065 2290.745 ;
        RECT 1072.095 2285.655 1072.425 2285.985 ;
        RECT 1084.055 2285.655 1084.385 2285.985 ;
        RECT 1054.615 2284.295 1054.945 2284.625 ;
        RECT 1061.975 2284.295 1062.305 2284.625 ;
        RECT 1066.575 2284.295 1066.905 2284.625 ;
        RECT 1084.020 2215.000 1087.020 2285.000 ;
        RECT 1089.590 2284.625 1089.890 2296.550 ;
        RECT 1094.190 2290.745 1094.490 2301.650 ;
        RECT 1094.970 2300.000 1095.270 2301.650 ;
        RECT 1095.590 2296.850 1095.890 2304.600 ;
        RECT 1100.810 2296.850 1101.110 2304.600 ;
        RECT 1095.590 2296.550 1096.330 2296.850 ;
        RECT 1094.175 2290.415 1094.505 2290.745 ;
        RECT 1096.030 2284.625 1096.330 2296.550 ;
        RECT 1100.630 2296.550 1101.110 2296.850 ;
        RECT 1101.430 2296.850 1101.730 2304.600 ;
        RECT 1106.650 2296.850 1106.950 2304.600 ;
        RECT 1107.270 2301.950 1107.570 2304.600 ;
        RECT 1107.270 2301.650 1110.130 2301.950 ;
        RECT 1107.270 2300.000 1107.570 2301.650 ;
        RECT 1101.430 2296.550 1101.850 2296.850 ;
        RECT 1106.650 2296.550 1107.370 2296.850 ;
        RECT 1100.630 2290.745 1100.930 2296.550 ;
        RECT 1100.615 2290.415 1100.945 2290.745 ;
        RECT 1101.550 2285.985 1101.850 2296.550 ;
        RECT 1107.070 2290.745 1107.370 2296.550 ;
        RECT 1107.055 2290.415 1107.385 2290.745 ;
        RECT 1101.535 2285.655 1101.865 2285.985 ;
        RECT 1089.575 2284.295 1089.905 2284.625 ;
        RECT 1096.015 2284.295 1096.345 2284.625 ;
        RECT 1102.020 2215.000 1105.020 2285.000 ;
        RECT 1109.830 2284.625 1110.130 2301.650 ;
        RECT 1112.490 2296.850 1112.790 2304.600 ;
        RECT 1113.110 2301.950 1113.410 2304.600 ;
        RECT 1113.110 2301.650 1116.570 2301.950 ;
        RECT 1113.110 2300.000 1113.410 2301.650 ;
        RECT 1112.490 2296.550 1112.890 2296.850 ;
        RECT 1112.590 2290.745 1112.890 2296.550 ;
        RECT 1112.575 2290.415 1112.905 2290.745 ;
        RECT 1116.270 2284.625 1116.570 2301.650 ;
        RECT 1118.330 2296.850 1118.630 2304.600 ;
        RECT 1118.110 2296.550 1118.630 2296.850 ;
        RECT 1118.950 2296.850 1119.250 2304.600 ;
        RECT 1124.170 2301.950 1124.470 2304.600 ;
        RECT 1121.790 2301.650 1124.470 2301.950 ;
        RECT 1118.950 2296.550 1119.330 2296.850 ;
        RECT 1118.110 2290.745 1118.410 2296.550 ;
        RECT 1118.095 2290.415 1118.425 2290.745 ;
        RECT 1119.030 2284.625 1119.330 2296.550 ;
        RECT 1121.790 2290.745 1122.090 2301.650 ;
        RECT 1124.170 2300.000 1124.470 2301.650 ;
        RECT 1124.790 2301.950 1125.090 2304.600 ;
        RECT 1130.010 2301.950 1130.310 2304.600 ;
        RECT 1124.790 2301.650 1128.530 2301.950 ;
        RECT 1124.790 2300.000 1125.090 2301.650 ;
        RECT 1121.775 2290.415 1122.105 2290.745 ;
        RECT 1128.230 2285.305 1128.530 2301.650 ;
        RECT 1129.150 2301.650 1130.310 2301.950 ;
        RECT 1129.150 2290.745 1129.450 2301.650 ;
        RECT 1130.010 2300.000 1130.310 2301.650 ;
        RECT 1130.630 2296.850 1130.930 2304.600 ;
        RECT 1135.850 2296.850 1136.150 2304.600 ;
        RECT 1130.630 2296.550 1131.290 2296.850 ;
        RECT 1129.135 2290.415 1129.465 2290.745 ;
        RECT 1109.815 2284.295 1110.145 2284.625 ;
        RECT 1116.255 2284.295 1116.585 2284.625 ;
        RECT 1119.015 2284.295 1119.345 2284.625 ;
        RECT 1120.020 2215.000 1123.020 2285.000 ;
        RECT 1128.215 2284.975 1128.545 2285.305 ;
        RECT 1130.990 2284.625 1131.290 2296.550 ;
        RECT 1135.590 2296.550 1136.150 2296.850 ;
        RECT 1136.470 2296.850 1136.770 2304.600 ;
        RECT 1141.690 2296.850 1141.990 2304.600 ;
        RECT 1142.310 2301.950 1142.610 2304.600 ;
        RECT 1142.310 2301.650 1145.090 2301.950 ;
        RECT 1142.310 2300.000 1142.610 2301.650 ;
        RECT 1136.470 2296.550 1136.810 2296.850 ;
        RECT 1141.690 2296.550 1142.330 2296.850 ;
        RECT 1135.590 2290.745 1135.890 2296.550 ;
        RECT 1135.575 2290.415 1135.905 2290.745 ;
        RECT 1136.510 2284.625 1136.810 2296.550 ;
        RECT 1142.030 2290.745 1142.330 2296.550 ;
        RECT 1142.015 2290.415 1142.345 2290.745 ;
        RECT 1144.790 2284.625 1145.090 2301.650 ;
        RECT 1147.530 2296.850 1147.830 2304.600 ;
        RECT 1148.150 2296.850 1148.450 2304.600 ;
        RECT 1153.370 2296.850 1153.670 2304.600 ;
        RECT 1147.530 2296.550 1147.850 2296.850 ;
        RECT 1148.150 2296.550 1148.770 2296.850 ;
        RECT 1147.550 2290.745 1147.850 2296.550 ;
        RECT 1147.535 2290.415 1147.865 2290.745 ;
        RECT 1148.470 2284.625 1148.770 2296.550 ;
        RECT 1153.070 2296.550 1153.670 2296.850 ;
        RECT 1153.070 2288.025 1153.370 2296.550 ;
        RECT 1153.055 2287.695 1153.385 2288.025 ;
        RECT 1153.990 2284.625 1154.290 2304.600 ;
        RECT 1159.210 2296.850 1159.510 2304.600 ;
        RECT 1159.830 2301.950 1160.130 2304.600 ;
        RECT 1165.050 2301.950 1165.350 2304.600 ;
        RECT 1159.830 2301.650 1163.490 2301.950 ;
        RECT 1159.830 2300.000 1160.130 2301.650 ;
        RECT 1159.210 2296.550 1159.810 2296.850 ;
        RECT 1159.510 2289.385 1159.810 2296.550 ;
        RECT 1159.495 2289.055 1159.825 2289.385 ;
        RECT 1163.190 2285.305 1163.490 2301.650 ;
        RECT 1164.110 2301.650 1165.350 2301.950 ;
        RECT 1164.110 2290.745 1164.410 2301.650 ;
        RECT 1165.050 2300.000 1165.350 2301.650 ;
        RECT 1165.670 2296.850 1165.970 2304.600 ;
        RECT 1170.890 2301.950 1171.190 2304.600 ;
        RECT 1165.030 2296.550 1165.970 2296.850 ;
        RECT 1167.790 2301.650 1171.190 2301.950 ;
        RECT 1164.095 2290.415 1164.425 2290.745 ;
        RECT 1163.175 2284.975 1163.505 2285.305 ;
        RECT 1165.030 2284.625 1165.330 2296.550 ;
        RECT 1167.790 2290.745 1168.090 2301.650 ;
        RECT 1170.890 2300.000 1171.190 2301.650 ;
        RECT 1171.510 2296.850 1171.810 2304.600 ;
        RECT 1176.730 2301.950 1177.030 2304.600 ;
        RECT 1171.470 2296.550 1171.810 2296.850 ;
        RECT 1173.310 2301.650 1177.030 2301.950 ;
        RECT 1167.775 2290.415 1168.105 2290.745 ;
        RECT 1171.470 2284.625 1171.770 2296.550 ;
        RECT 1173.310 2290.065 1173.610 2301.650 ;
        RECT 1176.730 2300.000 1177.030 2301.650 ;
        RECT 1177.350 2301.950 1177.650 2304.600 ;
        RECT 1177.350 2301.650 1179.130 2301.950 ;
        RECT 1177.350 2300.000 1177.650 2301.650 ;
        RECT 1173.295 2289.735 1173.625 2290.065 ;
        RECT 1178.830 2284.625 1179.130 2301.650 ;
        RECT 1182.570 2296.850 1182.870 2304.600 ;
        RECT 1182.510 2296.550 1182.870 2296.850 ;
        RECT 1183.190 2296.850 1183.490 2304.600 ;
        RECT 1188.410 2301.950 1188.710 2304.600 ;
        RECT 1187.110 2301.650 1188.710 2301.950 ;
        RECT 1183.190 2296.550 1183.730 2296.850 ;
        RECT 1182.510 2289.385 1182.810 2296.550 ;
        RECT 1182.495 2289.055 1182.825 2289.385 ;
        RECT 1183.430 2284.625 1183.730 2296.550 ;
        RECT 1187.110 2288.705 1187.410 2301.650 ;
        RECT 1188.410 2300.000 1188.710 2301.650 ;
        RECT 1189.030 2296.850 1189.330 2304.600 ;
        RECT 1188.950 2296.550 1189.330 2296.850 ;
        RECT 1194.250 2296.850 1194.550 2304.600 ;
        RECT 1194.870 2301.950 1195.170 2304.600 ;
        RECT 1584.010 2301.950 1584.310 2304.600 ;
        RECT 1589.850 2301.950 1590.150 2304.600 ;
        RECT 1194.870 2301.650 1198.450 2301.950 ;
        RECT 1194.870 2300.000 1195.170 2301.650 ;
        RECT 1194.250 2296.550 1194.770 2296.850 ;
        RECT 1187.095 2288.375 1187.425 2288.705 ;
        RECT 1188.950 2284.625 1189.250 2296.550 ;
        RECT 1194.470 2288.705 1194.770 2296.550 ;
        RECT 1194.455 2288.375 1194.785 2288.705 ;
        RECT 1198.150 2284.625 1198.450 2301.650 ;
        RECT 1580.870 2301.650 1584.310 2301.950 ;
        RECT 1130.975 2284.295 1131.305 2284.625 ;
        RECT 1136.495 2284.295 1136.825 2284.625 ;
        RECT 1144.775 2284.295 1145.105 2284.625 ;
        RECT 1148.455 2284.295 1148.785 2284.625 ;
        RECT 1153.975 2284.295 1154.305 2284.625 ;
        RECT 1165.015 2284.295 1165.345 2284.625 ;
        RECT 1171.455 2284.295 1171.785 2284.625 ;
        RECT 1178.815 2284.295 1179.145 2284.625 ;
        RECT 1183.415 2284.295 1183.745 2284.625 ;
        RECT 1188.935 2284.295 1189.265 2284.625 ;
        RECT 1198.135 2284.295 1198.465 2284.625 ;
        RECT 1210.020 2215.000 1213.020 2285.000 ;
        RECT 1228.020 2215.000 1231.020 2285.000 ;
        RECT 1264.020 2215.000 1267.020 2285.000 ;
        RECT 1282.020 2215.000 1285.020 2285.000 ;
        RECT 1300.020 2215.000 1303.020 2285.000 ;
        RECT 1580.870 2284.625 1581.170 2301.650 ;
        RECT 1584.010 2300.000 1584.310 2301.650 ;
        RECT 1587.310 2301.650 1590.150 2301.950 ;
        RECT 1587.310 2289.385 1587.610 2301.650 ;
        RECT 1589.850 2300.000 1590.150 2301.650 ;
        RECT 1595.690 2296.850 1595.990 2304.600 ;
        RECT 1601.530 2296.850 1601.830 2304.600 ;
        RECT 1607.370 2301.950 1607.670 2304.600 ;
        RECT 1595.590 2296.550 1595.990 2296.850 ;
        RECT 1601.110 2296.550 1601.830 2296.850 ;
        RECT 1604.790 2301.650 1607.670 2301.950 ;
        RECT 1587.295 2289.055 1587.625 2289.385 ;
        RECT 1595.590 2284.625 1595.890 2296.550 ;
        RECT 1601.110 2284.625 1601.410 2296.550 ;
        RECT 1604.790 2285.305 1605.090 2301.650 ;
        RECT 1607.370 2300.000 1607.670 2301.650 ;
        RECT 1613.210 2296.850 1613.510 2304.600 ;
        RECT 1613.070 2296.550 1613.510 2296.850 ;
        RECT 1613.830 2296.850 1614.130 2304.600 ;
        RECT 1619.050 2303.650 1619.350 2304.600 ;
        RECT 1617.670 2303.350 1619.350 2303.650 ;
        RECT 1613.830 2296.550 1614.290 2296.850 ;
        RECT 1613.070 2290.065 1613.370 2296.550 ;
        RECT 1613.990 2290.745 1614.290 2296.550 ;
        RECT 1613.975 2290.415 1614.305 2290.745 ;
        RECT 1617.670 2290.065 1617.970 2303.350 ;
        RECT 1619.050 2300.000 1619.350 2303.350 ;
        RECT 1619.670 2296.850 1619.970 2304.600 ;
        RECT 1624.890 2301.950 1625.190 2304.600 ;
        RECT 1619.510 2296.550 1619.970 2296.850 ;
        RECT 1624.110 2301.650 1625.190 2301.950 ;
        RECT 1619.510 2290.745 1619.810 2296.550 ;
        RECT 1619.495 2290.415 1619.825 2290.745 ;
        RECT 1613.055 2289.735 1613.385 2290.065 ;
        RECT 1617.655 2289.735 1617.985 2290.065 ;
        RECT 1624.110 2289.385 1624.410 2301.650 ;
        RECT 1624.890 2300.000 1625.190 2301.650 ;
        RECT 1625.510 2296.850 1625.810 2304.600 ;
        RECT 1630.730 2296.850 1631.030 2304.600 ;
        RECT 1625.030 2296.550 1625.810 2296.850 ;
        RECT 1630.550 2296.550 1631.030 2296.850 ;
        RECT 1631.350 2296.850 1631.650 2304.600 ;
        RECT 1636.570 2297.545 1636.870 2304.600 ;
        RECT 1636.555 2297.215 1636.885 2297.545 ;
        RECT 1637.190 2296.850 1637.490 2304.600 ;
        RECT 1642.410 2297.545 1642.710 2304.600 ;
        RECT 1642.395 2297.215 1642.725 2297.545 ;
        RECT 1643.030 2296.850 1643.330 2304.600 ;
        RECT 1644.335 2297.215 1644.665 2297.545 ;
        RECT 1631.350 2296.550 1631.770 2296.850 ;
        RECT 1624.095 2289.055 1624.425 2289.385 ;
        RECT 1625.030 2285.985 1625.330 2296.550 ;
        RECT 1630.550 2289.385 1630.850 2296.550 ;
        RECT 1631.470 2290.745 1631.770 2296.550 ;
        RECT 1636.990 2296.550 1637.490 2296.850 ;
        RECT 1642.510 2296.550 1643.330 2296.850 ;
        RECT 1636.990 2290.745 1637.290 2296.550 ;
        RECT 1631.455 2290.415 1631.785 2290.745 ;
        RECT 1636.975 2290.415 1637.305 2290.745 ;
        RECT 1630.535 2289.055 1630.865 2289.385 ;
        RECT 1642.510 2285.985 1642.810 2296.550 ;
        RECT 1644.350 2290.745 1644.650 2297.215 ;
        RECT 1648.250 2296.850 1648.550 2304.600 ;
        RECT 1648.870 2301.950 1649.170 2304.600 ;
        RECT 1654.090 2301.950 1654.390 2304.600 ;
        RECT 1648.870 2300.000 1649.250 2301.950 ;
        RECT 1648.030 2296.550 1648.550 2296.850 ;
        RECT 1644.335 2290.415 1644.665 2290.745 ;
        RECT 1648.030 2290.065 1648.330 2296.550 ;
        RECT 1648.015 2289.735 1648.345 2290.065 ;
        RECT 1648.950 2286.665 1649.250 2300.000 ;
        RECT 1652.630 2301.650 1654.390 2301.950 ;
        RECT 1652.630 2289.385 1652.930 2301.650 ;
        RECT 1654.090 2300.000 1654.390 2301.650 ;
        RECT 1654.710 2296.850 1655.010 2304.600 ;
        RECT 1659.930 2301.950 1660.230 2304.600 ;
        RECT 1654.470 2296.550 1655.010 2296.850 ;
        RECT 1659.070 2301.650 1660.230 2301.950 ;
        RECT 1654.470 2290.745 1654.770 2296.550 ;
        RECT 1659.070 2290.745 1659.370 2301.650 ;
        RECT 1659.930 2300.000 1660.230 2301.650 ;
        RECT 1660.550 2296.850 1660.850 2304.600 ;
        RECT 1665.770 2296.850 1666.070 2304.600 ;
        RECT 1659.990 2296.550 1660.850 2296.850 ;
        RECT 1665.510 2296.550 1666.070 2296.850 ;
        RECT 1666.390 2296.850 1666.690 2304.600 ;
        RECT 1671.610 2303.650 1671.910 2304.600 ;
        RECT 1670.110 2303.350 1671.910 2303.650 ;
        RECT 1666.390 2296.550 1666.730 2296.850 ;
        RECT 1654.455 2290.415 1654.785 2290.745 ;
        RECT 1659.055 2290.415 1659.385 2290.745 ;
        RECT 1652.615 2289.055 1652.945 2289.385 ;
        RECT 1659.990 2288.705 1660.290 2296.550 ;
        RECT 1665.510 2290.745 1665.810 2296.550 ;
        RECT 1665.495 2290.415 1665.825 2290.745 ;
        RECT 1659.975 2288.375 1660.305 2288.705 ;
        RECT 1648.935 2286.335 1649.265 2286.665 ;
        RECT 1625.015 2285.655 1625.345 2285.985 ;
        RECT 1642.495 2285.655 1642.825 2285.985 ;
        RECT 1604.775 2284.975 1605.105 2285.305 ;
        RECT 1666.430 2284.625 1666.730 2296.550 ;
        RECT 1670.110 2290.745 1670.410 2303.350 ;
        RECT 1671.610 2300.000 1671.910 2303.350 ;
        RECT 1672.230 2296.850 1672.530 2304.600 ;
        RECT 1677.450 2301.950 1677.750 2304.600 ;
        RECT 1671.950 2296.550 1672.530 2296.850 ;
        RECT 1676.550 2301.650 1677.750 2301.950 ;
        RECT 1670.095 2290.415 1670.425 2290.745 ;
        RECT 1671.950 2284.625 1672.250 2296.550 ;
        RECT 1676.550 2290.745 1676.850 2301.650 ;
        RECT 1677.450 2300.000 1677.750 2301.650 ;
        RECT 1678.070 2296.850 1678.370 2304.600 ;
        RECT 1683.290 2296.850 1683.590 2304.600 ;
        RECT 1677.470 2296.550 1678.370 2296.850 ;
        RECT 1682.990 2296.550 1683.590 2296.850 ;
        RECT 1676.535 2290.415 1676.865 2290.745 ;
        RECT 1677.470 2285.985 1677.770 2296.550 ;
        RECT 1682.990 2290.745 1683.290 2296.550 ;
        RECT 1682.975 2290.415 1683.305 2290.745 ;
        RECT 1677.455 2285.655 1677.785 2285.985 ;
        RECT 1683.910 2284.625 1684.210 2304.600 ;
        RECT 1689.130 2301.950 1689.430 2304.600 ;
        RECT 1688.510 2301.650 1689.430 2301.950 ;
        RECT 1688.510 2290.745 1688.810 2301.650 ;
        RECT 1689.130 2300.000 1689.430 2301.650 ;
        RECT 1689.750 2296.850 1690.050 2304.600 ;
        RECT 1694.970 2296.850 1695.270 2304.600 ;
        RECT 1689.430 2296.550 1690.050 2296.850 ;
        RECT 1694.950 2296.550 1695.270 2296.850 ;
        RECT 1695.590 2296.850 1695.890 2304.600 ;
        RECT 1700.810 2303.650 1701.110 2304.600 ;
        RECT 1699.550 2303.350 1701.110 2303.650 ;
        RECT 1695.590 2296.550 1696.170 2296.850 ;
        RECT 1688.495 2290.415 1688.825 2290.745 ;
        RECT 1689.430 2285.305 1689.730 2296.550 ;
        RECT 1694.950 2290.745 1695.250 2296.550 ;
        RECT 1694.935 2290.415 1695.265 2290.745 ;
        RECT 1689.415 2284.975 1689.745 2285.305 ;
        RECT 1695.870 2284.625 1696.170 2296.550 ;
        RECT 1699.550 2290.745 1699.850 2303.350 ;
        RECT 1700.810 2300.000 1701.110 2303.350 ;
        RECT 1701.430 2296.850 1701.730 2304.600 ;
        RECT 1706.650 2301.950 1706.950 2304.600 ;
        RECT 1701.390 2296.550 1701.730 2296.850 ;
        RECT 1705.990 2301.650 1706.950 2301.950 ;
        RECT 1699.535 2290.415 1699.865 2290.745 ;
        RECT 1701.390 2284.625 1701.690 2296.550 ;
        RECT 1705.990 2290.745 1706.290 2301.650 ;
        RECT 1706.650 2300.000 1706.950 2301.650 ;
        RECT 1707.270 2296.850 1707.570 2304.600 ;
        RECT 1712.490 2296.850 1712.790 2304.600 ;
        RECT 1706.910 2296.550 1707.570 2296.850 ;
        RECT 1712.430 2296.550 1712.790 2296.850 ;
        RECT 1713.110 2296.850 1713.410 2304.600 ;
        RECT 1718.330 2296.850 1718.630 2304.600 ;
        RECT 1718.950 2301.950 1719.250 2304.600 ;
        RECT 1724.170 2301.950 1724.470 2304.600 ;
        RECT 1718.950 2301.650 1720.090 2301.950 ;
        RECT 1718.950 2300.000 1719.250 2301.650 ;
        RECT 1713.110 2296.550 1713.650 2296.850 ;
        RECT 1705.975 2290.415 1706.305 2290.745 ;
        RECT 1706.910 2285.985 1707.210 2296.550 ;
        RECT 1712.430 2290.065 1712.730 2296.550 ;
        RECT 1713.350 2290.745 1713.650 2296.550 ;
        RECT 1717.950 2296.550 1718.630 2296.850 ;
        RECT 1713.335 2290.415 1713.665 2290.745 ;
        RECT 1717.950 2290.065 1718.250 2296.550 ;
        RECT 1719.790 2290.745 1720.090 2301.650 ;
        RECT 1723.470 2301.650 1724.470 2301.950 ;
        RECT 1723.470 2290.745 1723.770 2301.650 ;
        RECT 1724.170 2300.000 1724.470 2301.650 ;
        RECT 1724.790 2296.850 1725.090 2304.600 ;
        RECT 1730.010 2296.850 1730.310 2304.600 ;
        RECT 1724.390 2296.550 1725.090 2296.850 ;
        RECT 1729.910 2296.550 1730.310 2296.850 ;
        RECT 1730.630 2296.850 1730.930 2304.600 ;
        RECT 1735.850 2303.650 1736.150 2304.600 ;
        RECT 1734.510 2303.350 1736.150 2303.650 ;
        RECT 1730.630 2296.550 1731.130 2296.850 ;
        RECT 1719.775 2290.415 1720.105 2290.745 ;
        RECT 1723.455 2290.415 1723.785 2290.745 ;
        RECT 1712.415 2289.735 1712.745 2290.065 ;
        RECT 1717.935 2289.735 1718.265 2290.065 ;
        RECT 1724.390 2288.705 1724.690 2296.550 ;
        RECT 1729.910 2290.065 1730.210 2296.550 ;
        RECT 1730.830 2290.745 1731.130 2296.550 ;
        RECT 1730.815 2290.415 1731.145 2290.745 ;
        RECT 1734.510 2290.065 1734.810 2303.350 ;
        RECT 1735.850 2300.000 1736.150 2303.350 ;
        RECT 1736.470 2296.850 1736.770 2304.600 ;
        RECT 1741.690 2301.950 1741.990 2304.600 ;
        RECT 1736.350 2296.550 1736.770 2296.850 ;
        RECT 1740.950 2301.650 1741.990 2301.950 ;
        RECT 1736.350 2290.745 1736.650 2296.550 ;
        RECT 1736.335 2290.415 1736.665 2290.745 ;
        RECT 1740.950 2290.065 1741.250 2301.650 ;
        RECT 1741.690 2300.000 1741.990 2301.650 ;
        RECT 1742.310 2296.850 1742.610 2304.600 ;
        RECT 1747.530 2296.850 1747.830 2304.600 ;
        RECT 1741.870 2296.550 1742.610 2296.850 ;
        RECT 1747.390 2296.550 1747.830 2296.850 ;
        RECT 1748.150 2296.850 1748.450 2304.600 ;
        RECT 1753.370 2296.850 1753.670 2304.600 ;
        RECT 1753.990 2301.950 1754.290 2304.600 ;
        RECT 1753.990 2301.650 1755.050 2301.950 ;
        RECT 1753.990 2300.000 1754.290 2301.650 ;
        RECT 1748.150 2296.550 1748.610 2296.850 ;
        RECT 1741.870 2290.745 1742.170 2296.550 ;
        RECT 1741.855 2290.415 1742.185 2290.745 ;
        RECT 1747.390 2290.065 1747.690 2296.550 ;
        RECT 1748.310 2290.745 1748.610 2296.550 ;
        RECT 1752.910 2296.550 1753.670 2296.850 ;
        RECT 1748.295 2290.415 1748.625 2290.745 ;
        RECT 1752.910 2290.065 1753.210 2296.550 ;
        RECT 1729.895 2289.735 1730.225 2290.065 ;
        RECT 1734.495 2289.735 1734.825 2290.065 ;
        RECT 1740.935 2289.735 1741.265 2290.065 ;
        RECT 1747.375 2289.735 1747.705 2290.065 ;
        RECT 1752.895 2289.735 1753.225 2290.065 ;
        RECT 1724.375 2288.375 1724.705 2288.705 ;
        RECT 1706.895 2285.655 1707.225 2285.985 ;
        RECT 1754.750 2284.625 1755.050 2301.650 ;
        RECT 1759.210 2298.225 1759.510 2304.600 ;
        RECT 1759.195 2297.895 1759.525 2298.225 ;
        RECT 1759.830 2296.850 1760.130 2304.600 ;
        RECT 1765.050 2296.850 1765.350 2304.600 ;
        RECT 1759.350 2296.550 1760.130 2296.850 ;
        RECT 1764.870 2296.550 1765.350 2296.850 ;
        RECT 1765.670 2296.850 1765.970 2304.600 ;
        RECT 1770.890 2301.950 1771.190 2304.600 ;
        RECT 1767.630 2301.650 1771.190 2301.950 ;
        RECT 1765.670 2296.550 1766.090 2296.850 ;
        RECT 1759.350 2284.625 1759.650 2296.550 ;
        RECT 1764.870 2290.745 1765.170 2296.550 ;
        RECT 1764.855 2290.415 1765.185 2290.745 ;
        RECT 1765.790 2285.305 1766.090 2296.550 ;
        RECT 1767.630 2290.745 1767.930 2301.650 ;
        RECT 1770.890 2300.000 1771.190 2301.650 ;
        RECT 1771.510 2296.850 1771.810 2304.600 ;
        RECT 1776.730 2301.950 1777.030 2304.600 ;
        RECT 1771.310 2296.550 1771.810 2296.850 ;
        RECT 1775.910 2301.650 1777.030 2301.950 ;
        RECT 1767.615 2290.415 1767.945 2290.745 ;
        RECT 1771.310 2285.985 1771.610 2296.550 ;
        RECT 1775.910 2289.385 1776.210 2301.650 ;
        RECT 1776.730 2300.000 1777.030 2301.650 ;
        RECT 1777.350 2296.850 1777.650 2304.600 ;
        RECT 1782.570 2296.850 1782.870 2304.600 ;
        RECT 1776.830 2296.550 1777.650 2296.850 ;
        RECT 1782.350 2296.550 1782.870 2296.850 ;
        RECT 1783.190 2296.850 1783.490 2304.600 ;
        RECT 1788.410 2303.650 1788.710 2304.600 ;
        RECT 1786.950 2303.350 1788.710 2303.650 ;
        RECT 1783.190 2296.550 1783.570 2296.850 ;
        RECT 1775.895 2289.055 1776.225 2289.385 ;
        RECT 1771.295 2285.655 1771.625 2285.985 ;
        RECT 1765.775 2284.975 1766.105 2285.305 ;
        RECT 1776.830 2284.625 1777.130 2296.550 ;
        RECT 1782.350 2290.065 1782.650 2296.550 ;
        RECT 1782.335 2289.735 1782.665 2290.065 ;
        RECT 1783.270 2284.625 1783.570 2296.550 ;
        RECT 1786.950 2288.705 1787.250 2303.350 ;
        RECT 1788.410 2300.000 1788.710 2303.350 ;
        RECT 1789.030 2296.850 1789.330 2304.600 ;
        RECT 1794.250 2297.545 1794.550 2304.600 ;
        RECT 1794.235 2297.215 1794.565 2297.545 ;
        RECT 1794.870 2296.850 1795.170 2304.600 ;
        RECT 1788.790 2296.550 1789.330 2296.850 ;
        RECT 1794.310 2296.550 1795.170 2296.850 ;
        RECT 2234.010 2296.850 2234.310 2304.600 ;
        RECT 2239.850 2296.850 2240.150 2304.600 ;
        RECT 2245.690 2301.950 2245.990 2304.600 ;
        RECT 2234.010 2296.550 2234.370 2296.850 ;
        RECT 1786.935 2288.375 1787.265 2288.705 ;
        RECT 1788.790 2284.625 1789.090 2296.550 ;
        RECT 1794.310 2284.625 1794.610 2296.550 ;
        RECT 2234.070 2284.625 2234.370 2296.550 ;
        RECT 2239.590 2296.550 2240.150 2296.850 ;
        RECT 2242.350 2301.650 2245.990 2301.950 ;
        RECT 2239.590 2285.305 2239.890 2296.550 ;
        RECT 2239.575 2284.975 2239.905 2285.305 ;
        RECT 2242.350 2284.625 2242.650 2301.650 ;
        RECT 2245.690 2300.000 2245.990 2301.650 ;
        RECT 2251.530 2296.850 2251.830 2304.600 ;
        RECT 2257.370 2296.850 2257.670 2304.600 ;
        RECT 2263.210 2297.545 2263.510 2304.600 ;
        RECT 2263.195 2297.215 2263.525 2297.545 ;
        RECT 2263.830 2296.850 2264.130 2304.600 ;
        RECT 2269.050 2301.950 2269.350 2304.600 ;
        RECT 2268.110 2301.650 2269.350 2301.950 ;
        RECT 2265.335 2297.215 2265.665 2297.545 ;
        RECT 2251.530 2296.550 2251.850 2296.850 ;
        RECT 2251.550 2284.625 2251.850 2296.550 ;
        RECT 2257.070 2296.550 2257.670 2296.850 ;
        RECT 2263.510 2296.550 2264.130 2296.850 ;
        RECT 2257.070 2285.985 2257.370 2296.550 ;
        RECT 2257.055 2285.655 2257.385 2285.985 ;
        RECT 2263.510 2284.625 2263.810 2296.550 ;
        RECT 2265.350 2284.625 2265.650 2297.215 ;
        RECT 2268.110 2284.625 2268.410 2301.650 ;
        RECT 2269.050 2300.000 2269.350 2301.650 ;
        RECT 2269.670 2296.850 2269.970 2304.600 ;
        RECT 2274.890 2303.650 2275.190 2304.600 ;
        RECT 2269.030 2296.550 2269.970 2296.850 ;
        RECT 2273.630 2303.350 2275.190 2303.650 ;
        RECT 2269.030 2287.345 2269.330 2296.550 ;
        RECT 2269.015 2287.015 2269.345 2287.345 ;
        RECT 2273.630 2285.985 2273.930 2303.350 ;
        RECT 2274.890 2300.000 2275.190 2303.350 ;
        RECT 2275.510 2296.850 2275.810 2304.600 ;
        RECT 2280.730 2301.950 2281.030 2304.600 ;
        RECT 2275.470 2296.550 2275.810 2296.850 ;
        RECT 2280.070 2301.650 2281.030 2301.950 ;
        RECT 2275.470 2287.345 2275.770 2296.550 ;
        RECT 2275.455 2287.015 2275.785 2287.345 ;
        RECT 2273.615 2285.655 2273.945 2285.985 ;
        RECT 2280.070 2285.305 2280.370 2301.650 ;
        RECT 2280.730 2300.000 2281.030 2301.650 ;
        RECT 2281.350 2296.850 2281.650 2304.600 ;
        RECT 2286.570 2296.850 2286.870 2304.600 ;
        RECT 2280.990 2296.550 2281.650 2296.850 ;
        RECT 2286.510 2296.550 2286.870 2296.850 ;
        RECT 2287.190 2296.850 2287.490 2304.600 ;
        RECT 2292.410 2303.650 2292.710 2304.600 ;
        RECT 2291.110 2303.350 2292.710 2303.650 ;
        RECT 2287.190 2296.550 2287.730 2296.850 ;
        RECT 2280.055 2284.975 2280.385 2285.305 ;
        RECT 2280.990 2284.625 2281.290 2296.550 ;
        RECT 2286.510 2284.625 2286.810 2296.550 ;
        RECT 2287.430 2288.025 2287.730 2296.550 ;
        RECT 2287.415 2287.695 2287.745 2288.025 ;
        RECT 2291.110 2285.985 2291.410 2303.350 ;
        RECT 2292.410 2300.000 2292.710 2303.350 ;
        RECT 2293.030 2296.850 2293.330 2304.600 ;
        RECT 2298.250 2301.950 2298.550 2304.600 ;
        RECT 2292.950 2296.550 2293.330 2296.850 ;
        RECT 2297.550 2301.650 2298.550 2301.950 ;
        RECT 2292.950 2289.385 2293.250 2296.550 ;
        RECT 2297.550 2290.065 2297.850 2301.650 ;
        RECT 2298.250 2300.000 2298.550 2301.650 ;
        RECT 2298.870 2296.850 2299.170 2304.600 ;
        RECT 2304.090 2296.850 2304.390 2304.600 ;
        RECT 2298.470 2296.550 2299.170 2296.850 ;
        RECT 2303.990 2296.550 2304.390 2296.850 ;
        RECT 2304.710 2296.850 2305.010 2304.600 ;
        RECT 2309.930 2303.650 2310.230 2304.600 ;
        RECT 2308.590 2303.350 2310.230 2303.650 ;
        RECT 2304.710 2296.550 2305.210 2296.850 ;
        RECT 2297.535 2289.735 2297.865 2290.065 ;
        RECT 2292.935 2289.055 2293.265 2289.385 ;
        RECT 2298.470 2288.025 2298.770 2296.550 ;
        RECT 2303.990 2288.705 2304.290 2296.550 ;
        RECT 2303.975 2288.375 2304.305 2288.705 ;
        RECT 2298.455 2287.695 2298.785 2288.025 ;
        RECT 2291.095 2285.655 2291.425 2285.985 ;
        RECT 2304.910 2284.625 2305.210 2296.550 ;
        RECT 2308.590 2290.745 2308.890 2303.350 ;
        RECT 2309.930 2300.000 2310.230 2303.350 ;
        RECT 2310.550 2296.850 2310.850 2304.600 ;
        RECT 2315.770 2301.950 2316.070 2304.600 ;
        RECT 2310.430 2296.550 2310.850 2296.850 ;
        RECT 2315.030 2301.650 2316.070 2301.950 ;
        RECT 2308.575 2290.415 2308.905 2290.745 ;
        RECT 2310.430 2285.985 2310.730 2296.550 ;
        RECT 2315.030 2290.745 2315.330 2301.650 ;
        RECT 2315.770 2300.000 2316.070 2301.650 ;
        RECT 2316.390 2296.850 2316.690 2304.600 ;
        RECT 2321.610 2296.850 2321.910 2304.600 ;
        RECT 2315.950 2296.550 2316.690 2296.850 ;
        RECT 2321.470 2296.550 2321.910 2296.850 ;
        RECT 2322.230 2296.850 2322.530 2304.600 ;
        RECT 2327.450 2303.650 2327.750 2304.600 ;
        RECT 2326.070 2303.350 2327.750 2303.650 ;
        RECT 2322.230 2296.550 2322.690 2296.850 ;
        RECT 2315.015 2290.415 2315.345 2290.745 ;
        RECT 2310.415 2285.655 2310.745 2285.985 ;
        RECT 2315.950 2284.625 2316.250 2296.550 ;
        RECT 2321.470 2290.745 2321.770 2296.550 ;
        RECT 2321.455 2290.415 2321.785 2290.745 ;
        RECT 2322.390 2284.625 2322.690 2296.550 ;
        RECT 2326.070 2290.745 2326.370 2303.350 ;
        RECT 2327.450 2300.000 2327.750 2303.350 ;
        RECT 2328.070 2296.850 2328.370 2304.600 ;
        RECT 2333.290 2301.950 2333.590 2304.600 ;
        RECT 2327.910 2296.550 2328.370 2296.850 ;
        RECT 2332.510 2301.650 2333.590 2301.950 ;
        RECT 2326.055 2290.415 2326.385 2290.745 ;
        RECT 2327.910 2284.625 2328.210 2296.550 ;
        RECT 2332.510 2289.385 2332.810 2301.650 ;
        RECT 2333.290 2300.000 2333.590 2301.650 ;
        RECT 2333.910 2296.850 2334.210 2304.600 ;
        RECT 2339.130 2296.850 2339.430 2304.600 ;
        RECT 2333.430 2296.550 2334.210 2296.850 ;
        RECT 2338.950 2296.550 2339.430 2296.850 ;
        RECT 2339.750 2296.850 2340.050 2304.600 ;
        RECT 2344.970 2303.650 2345.270 2304.600 ;
        RECT 2343.550 2303.350 2345.270 2303.650 ;
        RECT 2339.750 2296.550 2340.170 2296.850 ;
        RECT 2332.495 2289.055 2332.825 2289.385 ;
        RECT 2333.430 2284.625 2333.730 2296.550 ;
        RECT 2338.950 2290.065 2339.250 2296.550 ;
        RECT 2338.935 2289.735 2339.265 2290.065 ;
        RECT 2339.870 2284.625 2340.170 2296.550 ;
        RECT 2343.550 2290.745 2343.850 2303.350 ;
        RECT 2344.970 2300.000 2345.270 2303.350 ;
        RECT 2345.590 2296.850 2345.890 2304.600 ;
        RECT 2350.810 2301.950 2351.110 2304.600 ;
        RECT 2345.390 2296.550 2345.890 2296.850 ;
        RECT 2349.990 2301.650 2351.110 2301.950 ;
        RECT 2343.535 2290.415 2343.865 2290.745 ;
        RECT 2345.390 2285.985 2345.690 2296.550 ;
        RECT 2349.990 2290.745 2350.290 2301.650 ;
        RECT 2350.810 2300.000 2351.110 2301.650 ;
        RECT 2351.430 2296.850 2351.730 2304.600 ;
        RECT 2356.650 2296.850 2356.950 2304.600 ;
        RECT 2350.910 2296.550 2351.730 2296.850 ;
        RECT 2356.430 2296.550 2356.950 2296.850 ;
        RECT 2357.270 2296.850 2357.570 2304.600 ;
        RECT 2362.490 2303.650 2362.790 2304.600 ;
        RECT 2361.030 2303.350 2362.790 2303.650 ;
        RECT 2357.270 2296.550 2357.650 2296.850 ;
        RECT 2349.975 2290.415 2350.305 2290.745 ;
        RECT 2345.375 2285.655 2345.705 2285.985 ;
        RECT 2350.910 2284.625 2351.210 2296.550 ;
        RECT 2356.430 2290.745 2356.730 2296.550 ;
        RECT 2356.415 2290.415 2356.745 2290.745 ;
        RECT 2357.350 2284.625 2357.650 2296.550 ;
        RECT 2361.030 2290.745 2361.330 2303.350 ;
        RECT 2362.490 2300.000 2362.790 2303.350 ;
        RECT 2363.110 2296.850 2363.410 2304.600 ;
        RECT 2368.330 2301.950 2368.630 2304.600 ;
        RECT 2362.870 2296.550 2363.410 2296.850 ;
        RECT 2367.470 2301.650 2368.630 2301.950 ;
        RECT 2361.015 2290.415 2361.345 2290.745 ;
        RECT 2362.870 2285.985 2363.170 2296.550 ;
        RECT 2367.470 2290.745 2367.770 2301.650 ;
        RECT 2368.330 2300.000 2368.630 2301.650 ;
        RECT 2368.950 2296.850 2369.250 2304.600 ;
        RECT 2374.170 2296.850 2374.470 2304.600 ;
        RECT 2368.390 2296.550 2369.250 2296.850 ;
        RECT 2373.910 2296.550 2374.470 2296.850 ;
        RECT 2374.790 2296.850 2375.090 2304.600 ;
        RECT 2380.010 2301.950 2380.310 2304.600 ;
        RECT 2377.590 2301.650 2380.310 2301.950 ;
        RECT 2374.790 2296.550 2375.130 2296.850 ;
        RECT 2367.455 2290.415 2367.785 2290.745 ;
        RECT 2362.855 2285.655 2363.185 2285.985 ;
        RECT 2368.390 2284.625 2368.690 2296.550 ;
        RECT 2373.910 2290.745 2374.210 2296.550 ;
        RECT 2373.895 2290.415 2374.225 2290.745 ;
        RECT 2374.830 2284.625 2375.130 2296.550 ;
        RECT 2377.590 2290.745 2377.890 2301.650 ;
        RECT 2380.010 2300.000 2380.310 2301.650 ;
        RECT 2380.630 2296.850 2380.930 2304.600 ;
        RECT 2385.850 2301.950 2386.150 2304.600 ;
        RECT 2380.350 2296.550 2380.930 2296.850 ;
        RECT 2384.950 2301.650 2386.150 2301.950 ;
        RECT 2377.575 2290.415 2377.905 2290.745 ;
        RECT 2380.350 2285.985 2380.650 2296.550 ;
        RECT 2384.950 2290.745 2385.250 2301.650 ;
        RECT 2385.850 2300.000 2386.150 2301.650 ;
        RECT 2386.470 2296.850 2386.770 2304.600 ;
        RECT 2391.690 2296.850 2391.990 2304.600 ;
        RECT 2385.870 2296.550 2386.770 2296.850 ;
        RECT 2391.390 2296.550 2391.990 2296.850 ;
        RECT 2384.935 2290.415 2385.265 2290.745 ;
        RECT 2385.870 2286.665 2386.170 2296.550 ;
        RECT 2391.390 2290.745 2391.690 2296.550 ;
        RECT 2391.375 2290.415 2391.705 2290.745 ;
        RECT 2392.310 2286.665 2392.610 2304.600 ;
        RECT 2397.530 2301.950 2397.830 2304.600 ;
        RECT 2396.910 2301.650 2397.830 2301.950 ;
        RECT 2396.910 2290.745 2397.210 2301.650 ;
        RECT 2397.530 2300.000 2397.830 2301.650 ;
        RECT 2398.150 2296.850 2398.450 2304.600 ;
        RECT 2403.370 2296.850 2403.670 2304.600 ;
        RECT 2397.830 2296.550 2398.450 2296.850 ;
        RECT 2403.350 2296.550 2403.670 2296.850 ;
        RECT 2403.990 2296.850 2404.290 2304.600 ;
        RECT 2409.210 2303.650 2409.510 2304.600 ;
        RECT 2407.950 2303.350 2409.510 2303.650 ;
        RECT 2403.990 2296.550 2404.570 2296.850 ;
        RECT 2396.895 2290.415 2397.225 2290.745 ;
        RECT 2397.830 2289.385 2398.130 2296.550 ;
        RECT 2403.350 2290.065 2403.650 2296.550 ;
        RECT 2403.335 2289.735 2403.665 2290.065 ;
        RECT 2404.270 2289.385 2404.570 2296.550 ;
        RECT 2397.815 2289.055 2398.145 2289.385 ;
        RECT 2404.255 2289.055 2404.585 2289.385 ;
        RECT 2407.950 2288.705 2408.250 2303.350 ;
        RECT 2409.210 2300.000 2409.510 2303.350 ;
        RECT 2409.830 2296.850 2410.130 2304.600 ;
        RECT 2415.050 2297.545 2415.350 2304.600 ;
        RECT 2415.035 2297.215 2415.365 2297.545 ;
        RECT 2415.670 2296.850 2415.970 2304.600 ;
        RECT 2420.890 2301.950 2421.190 2304.600 ;
        RECT 2409.790 2296.550 2410.130 2296.850 ;
        RECT 2415.310 2296.550 2415.970 2296.850 ;
        RECT 2418.070 2301.650 2421.190 2301.950 ;
        RECT 2407.935 2288.375 2408.265 2288.705 ;
        RECT 2385.855 2286.335 2386.185 2286.665 ;
        RECT 2392.295 2286.335 2392.625 2286.665 ;
        RECT 2409.790 2285.985 2410.090 2296.550 ;
        RECT 2415.310 2290.745 2415.610 2296.550 ;
        RECT 2415.295 2290.415 2415.625 2290.745 ;
        RECT 2418.070 2287.345 2418.370 2301.650 ;
        RECT 2420.890 2300.000 2421.190 2301.650 ;
        RECT 2421.510 2296.850 2421.810 2304.600 ;
        RECT 2426.730 2301.950 2427.030 2304.600 ;
        RECT 2420.830 2296.550 2421.810 2296.850 ;
        RECT 2423.590 2301.650 2427.030 2301.950 ;
        RECT 2420.830 2290.745 2421.130 2296.550 ;
        RECT 2420.815 2290.415 2421.145 2290.745 ;
        RECT 2423.590 2289.385 2423.890 2301.650 ;
        RECT 2426.730 2300.000 2427.030 2301.650 ;
        RECT 2427.350 2296.850 2427.650 2304.600 ;
        RECT 2432.570 2301.950 2432.870 2304.600 ;
        RECT 2427.270 2296.550 2427.650 2296.850 ;
        RECT 2430.030 2301.650 2432.870 2301.950 ;
        RECT 2427.270 2290.745 2427.570 2296.550 ;
        RECT 2427.255 2290.415 2427.585 2290.745 ;
        RECT 2423.575 2289.055 2423.905 2289.385 ;
        RECT 2430.030 2288.705 2430.330 2301.650 ;
        RECT 2432.570 2300.000 2432.870 2301.650 ;
        RECT 2433.190 2296.850 2433.490 2304.600 ;
        RECT 2438.410 2296.850 2438.710 2304.600 ;
        RECT 2432.790 2296.550 2433.490 2296.850 ;
        RECT 2438.310 2296.550 2438.710 2296.850 ;
        RECT 2439.030 2296.850 2439.330 2304.600 ;
        RECT 2444.250 2301.950 2444.550 2304.600 ;
        RECT 2442.910 2301.650 2444.550 2301.950 ;
        RECT 2439.030 2296.550 2439.530 2296.850 ;
        RECT 2430.015 2288.375 2430.345 2288.705 ;
        RECT 2432.790 2287.345 2433.090 2296.550 ;
        RECT 2438.310 2290.065 2438.610 2296.550 ;
        RECT 2438.295 2289.735 2438.625 2290.065 ;
        RECT 2439.230 2288.025 2439.530 2296.550 ;
        RECT 2442.910 2288.705 2443.210 2301.650 ;
        RECT 2444.250 2300.000 2444.550 2301.650 ;
        RECT 2444.870 2296.850 2445.170 2304.600 ;
        RECT 2444.750 2296.550 2445.170 2296.850 ;
        RECT 2442.895 2288.375 2443.225 2288.705 ;
        RECT 2439.215 2287.695 2439.545 2288.025 ;
        RECT 2444.750 2287.345 2445.050 2296.550 ;
        RECT 2418.055 2287.015 2418.385 2287.345 ;
        RECT 2432.775 2287.015 2433.105 2287.345 ;
        RECT 2444.735 2287.015 2445.065 2287.345 ;
        RECT 2380.335 2285.655 2380.665 2285.985 ;
        RECT 2409.775 2285.655 2410.105 2285.985 ;
        RECT 1580.855 2284.295 1581.185 2284.625 ;
        RECT 1595.575 2284.295 1595.905 2284.625 ;
        RECT 1601.095 2284.295 1601.425 2284.625 ;
        RECT 1666.415 2284.295 1666.745 2284.625 ;
        RECT 1671.935 2284.295 1672.265 2284.625 ;
        RECT 1683.895 2284.295 1684.225 2284.625 ;
        RECT 1695.855 2284.295 1696.185 2284.625 ;
        RECT 1701.375 2284.295 1701.705 2284.625 ;
        RECT 1754.735 2284.295 1755.065 2284.625 ;
        RECT 1759.335 2284.295 1759.665 2284.625 ;
        RECT 1776.815 2284.295 1777.145 2284.625 ;
        RECT 1783.255 2284.295 1783.585 2284.625 ;
        RECT 1788.775 2284.295 1789.105 2284.625 ;
        RECT 1794.295 2284.295 1794.625 2284.625 ;
        RECT 2234.055 2284.295 2234.385 2284.625 ;
        RECT 2242.335 2284.295 2242.665 2284.625 ;
        RECT 2251.535 2284.295 2251.865 2284.625 ;
        RECT 2263.495 2284.295 2263.825 2284.625 ;
        RECT 2265.335 2284.295 2265.665 2284.625 ;
        RECT 2268.095 2284.295 2268.425 2284.625 ;
        RECT 2280.975 2284.295 2281.305 2284.625 ;
        RECT 2286.495 2284.295 2286.825 2284.625 ;
        RECT 2304.895 2284.295 2305.225 2284.625 ;
        RECT 2315.935 2284.295 2316.265 2284.625 ;
        RECT 2322.375 2284.295 2322.705 2284.625 ;
        RECT 2327.895 2284.295 2328.225 2284.625 ;
        RECT 2333.415 2284.295 2333.745 2284.625 ;
        RECT 2339.855 2284.295 2340.185 2284.625 ;
        RECT 2350.895 2284.295 2351.225 2284.625 ;
        RECT 2357.335 2284.295 2357.665 2284.625 ;
        RECT 2368.375 2284.295 2368.705 2284.625 ;
        RECT 2374.815 2284.295 2375.145 2284.625 ;
      LAYER met4 ;
        RECT 306.735 1010.640 320.640 2188.880 ;
        RECT 323.040 1010.640 397.440 2188.880 ;
        RECT 399.840 1010.640 1486.505 2188.880 ;
  END
END user_project_wrapper
END LIBRARY

