VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 28.980 2924.800 30.180 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2374.980 2924.800 2376.180 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2609.580 2924.800 2610.780 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2844.180 2924.800 2845.380 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3078.780 2924.800 3079.980 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3313.380 2924.800 3314.580 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 263.580 2924.800 264.780 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3482.700 2.400 3483.900 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3195.060 2.400 3196.260 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2908.100 2.400 2909.300 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2620.460 2.400 2621.660 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2333.500 2.400 2334.700 ;
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2045.860 2.400 2047.060 ;
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 498.180 2924.800 499.380 ;
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1758.900 2.400 1760.100 ;
    END
  END analog_io[30]
  PIN analog_io[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 732.780 2924.800 733.980 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 967.380 2924.800 968.580 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1201.980 2924.800 1203.180 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1436.580 2924.800 1437.780 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1671.180 2924.800 1672.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1905.780 2924.800 1906.980 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2140.380 2924.800 2141.580 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 296.310 89.660 296.630 89.720 ;
        RECT 2898.990 89.660 2899.310 89.720 ;
        RECT 296.310 89.520 2899.310 89.660 ;
        RECT 296.310 89.460 296.630 89.520 ;
        RECT 2898.990 89.460 2899.310 89.520 ;
      LAYER via ;
        RECT 296.340 89.460 296.600 89.720 ;
        RECT 2899.020 89.460 2899.280 89.720 ;
      LAYER met2 ;
        RECT 296.330 1504.995 296.610 1505.365 ;
        RECT 296.400 89.750 296.540 1504.995 ;
        RECT 296.340 89.430 296.600 89.750 ;
        RECT 2899.020 89.430 2899.280 89.750 ;
        RECT 2899.080 88.245 2899.220 89.430 ;
        RECT 2899.010 87.875 2899.290 88.245 ;
      LAYER via2 ;
        RECT 296.330 1505.040 296.610 1505.320 ;
        RECT 2899.010 87.920 2899.290 88.200 ;
      LAYER met3 ;
        RECT 296.305 1505.330 296.635 1505.345 ;
        RECT 300.000 1505.330 304.000 1505.400 ;
        RECT 296.305 1505.030 304.000 1505.330 ;
        RECT 296.305 1505.015 296.635 1505.030 ;
        RECT 300.000 1504.800 304.000 1505.030 ;
        RECT 2898.985 88.210 2899.315 88.225 ;
        RECT 2917.600 88.210 2924.800 88.660 ;
        RECT 2898.985 87.910 2924.800 88.210 ;
        RECT 2898.985 87.895 2899.315 87.910 ;
        RECT 2917.600 87.460 2924.800 87.910 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 299.990 2691.680 300.310 2691.740 ;
        RECT 2818.490 2691.680 2818.810 2691.740 ;
        RECT 299.990 2691.540 2818.810 2691.680 ;
        RECT 299.990 2691.480 300.310 2691.540 ;
        RECT 2818.490 2691.480 2818.810 2691.540 ;
        RECT 2818.490 2650.200 2818.810 2650.260 ;
        RECT 2818.490 2650.060 2829.300 2650.200 ;
        RECT 2818.490 2650.000 2818.810 2650.060 ;
        RECT 2829.160 2649.520 2829.300 2650.060 ;
        RECT 2846.090 2649.520 2846.410 2649.580 ;
        RECT 2829.160 2649.380 2846.410 2649.520 ;
        RECT 2846.090 2649.320 2846.410 2649.380 ;
        RECT 2846.090 2608.040 2846.410 2608.100 ;
        RECT 2854.830 2608.040 2855.150 2608.100 ;
        RECT 2846.090 2607.900 2855.150 2608.040 ;
        RECT 2846.090 2607.840 2846.410 2607.900 ;
        RECT 2854.830 2607.840 2855.150 2607.900 ;
        RECT 2854.830 2587.640 2855.150 2587.700 ;
        RECT 2854.830 2587.500 2856.900 2587.640 ;
        RECT 2854.830 2587.440 2855.150 2587.500 ;
        RECT 2856.760 2587.300 2856.900 2587.500 ;
        RECT 2866.790 2587.300 2867.110 2587.360 ;
        RECT 2856.760 2587.160 2867.110 2587.300 ;
        RECT 2866.790 2587.100 2867.110 2587.160 ;
        RECT 2866.790 2497.880 2867.110 2497.940 ;
        RECT 2866.790 2497.740 2870.700 2497.880 ;
        RECT 2866.790 2497.680 2867.110 2497.740 ;
        RECT 2870.560 2497.540 2870.700 2497.740 ;
        RECT 2883.810 2497.540 2884.130 2497.600 ;
        RECT 2870.560 2497.400 2884.130 2497.540 ;
        RECT 2883.810 2497.340 2884.130 2497.400 ;
        RECT 2884.270 2469.320 2884.590 2469.380 ;
        RECT 2894.390 2469.320 2894.710 2469.380 ;
        RECT 2884.270 2469.180 2894.710 2469.320 ;
        RECT 2884.270 2469.120 2884.590 2469.180 ;
        RECT 2894.390 2469.120 2894.710 2469.180 ;
        RECT 293.550 2145.980 293.870 2146.040 ;
        RECT 299.990 2145.980 300.310 2146.040 ;
        RECT 293.550 2145.840 300.310 2145.980 ;
        RECT 293.550 2145.780 293.870 2145.840 ;
        RECT 299.990 2145.780 300.310 2145.840 ;
        RECT 288.490 2069.820 288.810 2069.880 ;
        RECT 293.550 2069.820 293.870 2069.880 ;
        RECT 288.490 2069.680 293.870 2069.820 ;
        RECT 288.490 2069.620 288.810 2069.680 ;
        RECT 293.550 2069.620 293.870 2069.680 ;
      LAYER via ;
        RECT 300.020 2691.480 300.280 2691.740 ;
        RECT 2818.520 2691.480 2818.780 2691.740 ;
        RECT 2818.520 2650.000 2818.780 2650.260 ;
        RECT 2846.120 2649.320 2846.380 2649.580 ;
        RECT 2846.120 2607.840 2846.380 2608.100 ;
        RECT 2854.860 2607.840 2855.120 2608.100 ;
        RECT 2854.860 2587.440 2855.120 2587.700 ;
        RECT 2866.820 2587.100 2867.080 2587.360 ;
        RECT 2866.820 2497.680 2867.080 2497.940 ;
        RECT 2883.840 2497.340 2884.100 2497.600 ;
        RECT 2884.300 2469.120 2884.560 2469.380 ;
        RECT 2894.420 2469.120 2894.680 2469.380 ;
        RECT 293.580 2145.780 293.840 2146.040 ;
        RECT 300.020 2145.780 300.280 2146.040 ;
        RECT 288.520 2069.620 288.780 2069.880 ;
        RECT 293.580 2069.620 293.840 2069.880 ;
      LAYER met2 ;
        RECT 300.020 2691.450 300.280 2691.770 ;
        RECT 2818.520 2691.450 2818.780 2691.770 ;
        RECT 300.080 2146.070 300.220 2691.450 ;
        RECT 2818.580 2650.290 2818.720 2691.450 ;
        RECT 2818.520 2649.970 2818.780 2650.290 ;
        RECT 2846.120 2649.290 2846.380 2649.610 ;
        RECT 2846.180 2608.130 2846.320 2649.290 ;
        RECT 2846.120 2607.810 2846.380 2608.130 ;
        RECT 2854.860 2607.810 2855.120 2608.130 ;
        RECT 2854.920 2587.730 2855.060 2607.810 ;
        RECT 2854.860 2587.410 2855.120 2587.730 ;
        RECT 2866.820 2587.070 2867.080 2587.390 ;
        RECT 2866.880 2497.970 2867.020 2587.070 ;
        RECT 2866.820 2497.650 2867.080 2497.970 ;
        RECT 2883.840 2497.310 2884.100 2497.630 ;
        RECT 2883.900 2483.770 2884.040 2497.310 ;
        RECT 2883.900 2483.630 2884.500 2483.770 ;
        RECT 2884.360 2469.410 2884.500 2483.630 ;
        RECT 2884.300 2469.090 2884.560 2469.410 ;
        RECT 2894.420 2469.090 2894.680 2469.410 ;
        RECT 2894.480 2434.245 2894.620 2469.090 ;
        RECT 2894.410 2433.875 2894.690 2434.245 ;
        RECT 293.580 2145.750 293.840 2146.070 ;
        RECT 300.020 2145.750 300.280 2146.070 ;
        RECT 293.640 2069.910 293.780 2145.750 ;
        RECT 288.520 2069.590 288.780 2069.910 ;
        RECT 293.580 2069.590 293.840 2069.910 ;
        RECT 288.580 1820.885 288.720 2069.590 ;
        RECT 288.510 1820.515 288.790 1820.885 ;
      LAYER via2 ;
        RECT 2894.410 2433.920 2894.690 2434.200 ;
        RECT 288.510 1820.560 288.790 1820.840 ;
      LAYER met3 ;
        RECT 2894.385 2434.210 2894.715 2434.225 ;
        RECT 2917.600 2434.210 2924.800 2434.660 ;
        RECT 2894.385 2433.910 2924.800 2434.210 ;
        RECT 2894.385 2433.895 2894.715 2433.910 ;
        RECT 2917.600 2433.460 2924.800 2433.910 ;
        RECT 288.485 1820.850 288.815 1820.865 ;
        RECT 300.000 1820.850 304.000 1820.920 ;
        RECT 288.485 1820.550 304.000 1820.850 ;
        RECT 288.485 1820.535 288.815 1820.550 ;
        RECT 300.000 1820.320 304.000 1820.550 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 290.790 2691.340 291.110 2691.400 ;
        RECT 2898.990 2691.340 2899.310 2691.400 ;
        RECT 290.790 2691.200 2899.310 2691.340 ;
        RECT 290.790 2691.140 291.110 2691.200 ;
        RECT 2898.990 2691.140 2899.310 2691.200 ;
      LAYER via ;
        RECT 290.820 2691.140 291.080 2691.400 ;
        RECT 2899.020 2691.140 2899.280 2691.400 ;
      LAYER met2 ;
        RECT 290.820 2691.110 291.080 2691.430 ;
        RECT 2899.020 2691.110 2899.280 2691.430 ;
        RECT 290.880 1852.165 291.020 2691.110 ;
        RECT 2899.080 2669.525 2899.220 2691.110 ;
        RECT 2899.010 2669.155 2899.290 2669.525 ;
        RECT 290.810 1851.795 291.090 1852.165 ;
      LAYER via2 ;
        RECT 2899.010 2669.200 2899.290 2669.480 ;
        RECT 290.810 1851.840 291.090 1852.120 ;
      LAYER met3 ;
        RECT 2898.985 2669.490 2899.315 2669.505 ;
        RECT 2917.600 2669.490 2924.800 2669.940 ;
        RECT 2898.985 2669.190 2924.800 2669.490 ;
        RECT 2898.985 2669.175 2899.315 2669.190 ;
        RECT 2917.600 2668.740 2924.800 2669.190 ;
        RECT 290.785 1852.130 291.115 1852.145 ;
        RECT 300.000 1852.130 304.000 1852.200 ;
        RECT 290.785 1851.830 304.000 1852.130 ;
        RECT 290.785 1851.815 291.115 1851.830 ;
        RECT 300.000 1851.600 304.000 1851.830 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 290.330 2694.740 290.650 2694.800 ;
        RECT 2903.130 2694.740 2903.450 2694.800 ;
        RECT 290.330 2694.600 2903.450 2694.740 ;
        RECT 290.330 2694.540 290.650 2694.600 ;
        RECT 2903.130 2694.540 2903.450 2694.600 ;
      LAYER via ;
        RECT 290.360 2694.540 290.620 2694.800 ;
        RECT 2903.160 2694.540 2903.420 2694.800 ;
      LAYER met2 ;
        RECT 2903.150 2903.755 2903.430 2904.125 ;
        RECT 2903.220 2694.830 2903.360 2903.755 ;
        RECT 290.360 2694.510 290.620 2694.830 ;
        RECT 2903.160 2694.510 2903.420 2694.830 ;
        RECT 290.420 1884.125 290.560 2694.510 ;
        RECT 290.350 1883.755 290.630 1884.125 ;
      LAYER via2 ;
        RECT 2903.150 2903.800 2903.430 2904.080 ;
        RECT 290.350 1883.800 290.630 1884.080 ;
      LAYER met3 ;
        RECT 2903.125 2904.090 2903.455 2904.105 ;
        RECT 2917.600 2904.090 2924.800 2904.540 ;
        RECT 2903.125 2903.790 2924.800 2904.090 ;
        RECT 2903.125 2903.775 2903.455 2903.790 ;
        RECT 2917.600 2903.340 2924.800 2903.790 ;
        RECT 290.325 1884.090 290.655 1884.105 ;
        RECT 300.000 1884.090 304.000 1884.160 ;
        RECT 290.325 1883.790 304.000 1884.090 ;
        RECT 290.325 1883.775 290.655 1883.790 ;
        RECT 300.000 1883.560 304.000 1883.790 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 289.870 2695.080 290.190 2695.140 ;
        RECT 2901.750 2695.080 2902.070 2695.140 ;
        RECT 289.870 2694.940 2902.070 2695.080 ;
        RECT 289.870 2694.880 290.190 2694.940 ;
        RECT 2901.750 2694.880 2902.070 2694.940 ;
      LAYER via ;
        RECT 289.900 2694.880 290.160 2695.140 ;
        RECT 2901.780 2694.880 2902.040 2695.140 ;
      LAYER met2 ;
        RECT 2901.770 3138.355 2902.050 3138.725 ;
        RECT 2901.840 2695.170 2901.980 3138.355 ;
        RECT 289.900 2694.850 290.160 2695.170 ;
        RECT 2901.780 2694.850 2902.040 2695.170 ;
        RECT 289.960 1915.405 290.100 2694.850 ;
        RECT 289.890 1915.035 290.170 1915.405 ;
      LAYER via2 ;
        RECT 2901.770 3138.400 2902.050 3138.680 ;
        RECT 289.890 1915.080 290.170 1915.360 ;
      LAYER met3 ;
        RECT 2901.745 3138.690 2902.075 3138.705 ;
        RECT 2917.600 3138.690 2924.800 3139.140 ;
        RECT 2901.745 3138.390 2924.800 3138.690 ;
        RECT 2901.745 3138.375 2902.075 3138.390 ;
        RECT 2917.600 3137.940 2924.800 3138.390 ;
        RECT 289.865 1915.370 290.195 1915.385 ;
        RECT 300.000 1915.370 304.000 1915.440 ;
        RECT 289.865 1915.070 304.000 1915.370 ;
        RECT 289.865 1915.055 290.195 1915.070 ;
        RECT 300.000 1914.840 304.000 1915.070 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 869.470 3369.640 869.790 3369.700 ;
        RECT 893.850 3369.640 894.170 3369.700 ;
        RECT 869.470 3369.500 894.170 3369.640 ;
        RECT 869.470 3369.440 869.790 3369.500 ;
        RECT 893.850 3369.440 894.170 3369.500 ;
        RECT 1835.470 3369.640 1835.790 3369.700 ;
        RECT 1859.850 3369.640 1860.170 3369.700 ;
        RECT 1835.470 3369.500 1860.170 3369.640 ;
        RECT 1835.470 3369.440 1835.790 3369.500 ;
        RECT 1859.850 3369.440 1860.170 3369.500 ;
        RECT 2801.470 3369.640 2801.790 3369.700 ;
        RECT 2825.850 3369.640 2826.170 3369.700 ;
        RECT 2801.470 3369.500 2826.170 3369.640 ;
        RECT 2801.470 3369.440 2801.790 3369.500 ;
        RECT 2825.850 3369.440 2826.170 3369.500 ;
        RECT 772.870 3368.960 773.190 3369.020 ;
        RECT 811.050 3368.960 811.370 3369.020 ;
        RECT 772.870 3368.820 811.370 3368.960 ;
        RECT 772.870 3368.760 773.190 3368.820 ;
        RECT 811.050 3368.760 811.370 3368.820 ;
        RECT 1449.070 3368.960 1449.390 3369.020 ;
        RECT 1463.330 3368.960 1463.650 3369.020 ;
        RECT 1449.070 3368.820 1463.650 3368.960 ;
        RECT 1449.070 3368.760 1449.390 3368.820 ;
        RECT 1463.330 3368.760 1463.650 3368.820 ;
        RECT 1738.870 3368.960 1739.190 3369.020 ;
        RECT 1777.050 3368.960 1777.370 3369.020 ;
        RECT 1738.870 3368.820 1777.370 3368.960 ;
        RECT 1738.870 3368.760 1739.190 3368.820 ;
        RECT 1777.050 3368.760 1777.370 3368.820 ;
        RECT 2704.870 3368.960 2705.190 3369.020 ;
        RECT 2743.050 3368.960 2743.370 3369.020 ;
        RECT 2704.870 3368.820 2743.370 3368.960 ;
        RECT 2704.870 3368.760 2705.190 3368.820 ;
        RECT 2743.050 3368.760 2743.370 3368.820 ;
      LAYER via ;
        RECT 869.500 3369.440 869.760 3369.700 ;
        RECT 893.880 3369.440 894.140 3369.700 ;
        RECT 1835.500 3369.440 1835.760 3369.700 ;
        RECT 1859.880 3369.440 1860.140 3369.700 ;
        RECT 2801.500 3369.440 2801.760 3369.700 ;
        RECT 2825.880 3369.440 2826.140 3369.700 ;
        RECT 772.900 3368.760 773.160 3369.020 ;
        RECT 811.080 3368.760 811.340 3369.020 ;
        RECT 1449.100 3368.760 1449.360 3369.020 ;
        RECT 1463.360 3368.760 1463.620 3369.020 ;
        RECT 1738.900 3368.760 1739.160 3369.020 ;
        RECT 1777.080 3368.760 1777.340 3369.020 ;
        RECT 2704.900 3368.760 2705.160 3369.020 ;
        RECT 2743.080 3368.760 2743.340 3369.020 ;
      LAYER met2 ;
        RECT 941.710 3370.235 941.990 3370.605 ;
        RECT 1897.590 3370.235 1897.870 3370.605 ;
        RECT 834.990 3369.555 835.270 3369.925 ;
        RECT 869.490 3369.555 869.770 3369.925 ;
        RECT 772.890 3368.875 773.170 3369.245 ;
        RECT 772.900 3368.730 773.160 3368.875 ;
        RECT 811.080 3368.730 811.340 3369.050 ;
        RECT 811.140 3367.885 811.280 3368.730 ;
        RECT 811.070 3367.515 811.350 3367.885 ;
        RECT 834.530 3367.770 834.810 3367.885 ;
        RECT 835.060 3367.770 835.200 3369.555 ;
        RECT 869.500 3369.410 869.760 3369.555 ;
        RECT 893.880 3369.410 894.140 3369.730 ;
        RECT 893.940 3369.245 894.080 3369.410 ;
        RECT 941.780 3369.245 941.920 3370.235 ;
        RECT 1800.530 3369.810 1800.810 3369.925 ;
        RECT 1801.450 3369.810 1801.730 3369.925 ;
        RECT 1800.530 3369.670 1801.730 3369.810 ;
        RECT 1800.530 3369.555 1800.810 3369.670 ;
        RECT 1801.450 3369.555 1801.730 3369.670 ;
        RECT 1835.490 3369.555 1835.770 3369.925 ;
        RECT 1835.500 3369.410 1835.760 3369.555 ;
        RECT 1859.880 3369.410 1860.140 3369.730 ;
        RECT 1859.940 3369.245 1860.080 3369.410 ;
        RECT 1897.660 3369.245 1897.800 3370.235 ;
        RECT 2766.990 3369.555 2767.270 3369.925 ;
        RECT 2801.490 3369.555 2801.770 3369.925 ;
        RECT 893.870 3368.875 894.150 3369.245 ;
        RECT 941.710 3368.875 941.990 3369.245 ;
        RECT 1449.090 3368.875 1449.370 3369.245 ;
        RECT 1449.100 3368.730 1449.360 3368.875 ;
        RECT 1463.360 3368.730 1463.620 3369.050 ;
        RECT 1738.890 3368.875 1739.170 3369.245 ;
        RECT 1738.900 3368.730 1739.160 3368.875 ;
        RECT 1777.080 3368.730 1777.340 3369.050 ;
        RECT 1859.870 3368.875 1860.150 3369.245 ;
        RECT 1897.590 3368.875 1897.870 3369.245 ;
        RECT 2704.890 3368.875 2705.170 3369.245 ;
        RECT 2704.900 3368.730 2705.160 3368.875 ;
        RECT 2743.080 3368.730 2743.340 3369.050 ;
        RECT 1463.420 3367.885 1463.560 3368.730 ;
        RECT 1777.140 3367.885 1777.280 3368.730 ;
        RECT 2743.140 3367.885 2743.280 3368.730 ;
        RECT 834.530 3367.630 835.200 3367.770 ;
        RECT 834.530 3367.515 834.810 3367.630 ;
        RECT 1463.350 3367.515 1463.630 3367.885 ;
        RECT 1777.070 3367.515 1777.350 3367.885 ;
        RECT 2743.070 3367.515 2743.350 3367.885 ;
        RECT 2766.530 3367.770 2766.810 3367.885 ;
        RECT 2767.060 3367.770 2767.200 3369.555 ;
        RECT 2801.500 3369.410 2801.760 3369.555 ;
        RECT 2825.880 3369.410 2826.140 3369.730 ;
        RECT 2825.940 3369.245 2826.080 3369.410 ;
        RECT 2825.870 3368.875 2826.150 3369.245 ;
        RECT 2863.590 3369.130 2863.870 3369.245 ;
        RECT 2863.200 3368.990 2863.870 3369.130 ;
        RECT 2863.200 3368.565 2863.340 3368.990 ;
        RECT 2863.590 3368.875 2863.870 3368.990 ;
        RECT 2863.130 3368.195 2863.410 3368.565 ;
        RECT 2766.530 3367.630 2767.200 3367.770 ;
        RECT 2766.530 3367.515 2766.810 3367.630 ;
      LAYER via2 ;
        RECT 941.710 3370.280 941.990 3370.560 ;
        RECT 1897.590 3370.280 1897.870 3370.560 ;
        RECT 834.990 3369.600 835.270 3369.880 ;
        RECT 869.490 3369.600 869.770 3369.880 ;
        RECT 772.890 3368.920 773.170 3369.200 ;
        RECT 811.070 3367.560 811.350 3367.840 ;
        RECT 834.530 3367.560 834.810 3367.840 ;
        RECT 1800.530 3369.600 1800.810 3369.880 ;
        RECT 1801.450 3369.600 1801.730 3369.880 ;
        RECT 1835.490 3369.600 1835.770 3369.880 ;
        RECT 2766.990 3369.600 2767.270 3369.880 ;
        RECT 2801.490 3369.600 2801.770 3369.880 ;
        RECT 893.870 3368.920 894.150 3369.200 ;
        RECT 941.710 3368.920 941.990 3369.200 ;
        RECT 1449.090 3368.920 1449.370 3369.200 ;
        RECT 1738.890 3368.920 1739.170 3369.200 ;
        RECT 1859.870 3368.920 1860.150 3369.200 ;
        RECT 1897.590 3368.920 1897.870 3369.200 ;
        RECT 2704.890 3368.920 2705.170 3369.200 ;
        RECT 1463.350 3367.560 1463.630 3367.840 ;
        RECT 1777.070 3367.560 1777.350 3367.840 ;
        RECT 2743.070 3367.560 2743.350 3367.840 ;
        RECT 2766.530 3367.560 2766.810 3367.840 ;
        RECT 2825.870 3368.920 2826.150 3369.200 ;
        RECT 2863.590 3368.920 2863.870 3369.200 ;
        RECT 2863.130 3368.240 2863.410 3368.520 ;
      LAYER met3 ;
        RECT 2917.600 3373.290 2924.800 3373.740 ;
        RECT 2916.710 3372.990 2924.800 3373.290 ;
        RECT 917.510 3370.570 917.890 3370.580 ;
        RECT 941.685 3370.570 942.015 3370.585 ;
        RECT 917.510 3370.270 942.015 3370.570 ;
        RECT 917.510 3370.260 917.890 3370.270 ;
        RECT 941.685 3370.255 942.015 3370.270 ;
        RECT 1883.510 3370.570 1883.890 3370.580 ;
        RECT 1897.565 3370.570 1897.895 3370.585 ;
        RECT 1883.510 3370.270 1897.895 3370.570 ;
        RECT 1883.510 3370.260 1883.890 3370.270 ;
        RECT 1897.565 3370.255 1897.895 3370.270 ;
        RECT 834.965 3369.890 835.295 3369.905 ;
        RECT 869.465 3369.890 869.795 3369.905 ;
        RECT 834.965 3369.590 869.795 3369.890 ;
        RECT 834.965 3369.575 835.295 3369.590 ;
        RECT 869.465 3369.575 869.795 3369.590 ;
        RECT 1786.910 3369.890 1787.290 3369.900 ;
        RECT 1800.505 3369.890 1800.835 3369.905 ;
        RECT 1786.910 3369.590 1800.835 3369.890 ;
        RECT 1786.910 3369.580 1787.290 3369.590 ;
        RECT 1800.505 3369.575 1800.835 3369.590 ;
        RECT 1801.425 3369.890 1801.755 3369.905 ;
        RECT 1835.465 3369.890 1835.795 3369.905 ;
        RECT 1801.425 3369.590 1835.795 3369.890 ;
        RECT 1801.425 3369.575 1801.755 3369.590 ;
        RECT 1835.465 3369.575 1835.795 3369.590 ;
        RECT 2766.965 3369.890 2767.295 3369.905 ;
        RECT 2801.465 3369.890 2801.795 3369.905 ;
        RECT 2766.965 3369.590 2801.795 3369.890 ;
        RECT 2766.965 3369.575 2767.295 3369.590 ;
        RECT 2801.465 3369.575 2801.795 3369.590 ;
        RECT 290.990 3369.210 291.370 3369.220 ;
        RECT 772.865 3369.210 773.195 3369.225 ;
        RECT 290.990 3368.910 324.450 3369.210 ;
        RECT 290.990 3368.900 291.370 3368.910 ;
        RECT 324.150 3368.530 324.450 3368.910 ;
        RECT 372.910 3368.910 421.050 3369.210 ;
        RECT 324.150 3368.230 372.290 3368.530 ;
        RECT 371.990 3367.850 372.290 3368.230 ;
        RECT 372.910 3367.850 373.210 3368.910 ;
        RECT 420.750 3368.530 421.050 3368.910 ;
        RECT 469.510 3368.910 517.650 3369.210 ;
        RECT 420.750 3368.230 468.890 3368.530 ;
        RECT 371.990 3367.550 373.210 3367.850 ;
        RECT 468.590 3367.850 468.890 3368.230 ;
        RECT 469.510 3367.850 469.810 3368.910 ;
        RECT 517.350 3368.530 517.650 3368.910 ;
        RECT 566.110 3368.910 614.250 3369.210 ;
        RECT 517.350 3368.230 565.490 3368.530 ;
        RECT 468.590 3367.550 469.810 3367.850 ;
        RECT 565.190 3367.850 565.490 3368.230 ;
        RECT 566.110 3367.850 566.410 3368.910 ;
        RECT 613.950 3368.530 614.250 3368.910 ;
        RECT 662.710 3368.910 710.850 3369.210 ;
        RECT 613.950 3368.230 662.090 3368.530 ;
        RECT 565.190 3367.550 566.410 3367.850 ;
        RECT 661.790 3367.850 662.090 3368.230 ;
        RECT 662.710 3367.850 663.010 3368.910 ;
        RECT 710.550 3368.530 710.850 3368.910 ;
        RECT 759.310 3368.910 773.195 3369.210 ;
        RECT 710.550 3368.230 758.690 3368.530 ;
        RECT 661.790 3367.550 663.010 3367.850 ;
        RECT 758.390 3367.850 758.690 3368.230 ;
        RECT 759.310 3367.850 759.610 3368.910 ;
        RECT 772.865 3368.895 773.195 3368.910 ;
        RECT 893.845 3369.210 894.175 3369.225 ;
        RECT 917.510 3369.210 917.890 3369.220 ;
        RECT 893.845 3368.910 917.890 3369.210 ;
        RECT 893.845 3368.895 894.175 3368.910 ;
        RECT 917.510 3368.900 917.890 3368.910 ;
        RECT 941.685 3369.210 942.015 3369.225 ;
        RECT 1449.065 3369.210 1449.395 3369.225 ;
        RECT 941.685 3368.910 1000.650 3369.210 ;
        RECT 941.685 3368.895 942.015 3368.910 ;
        RECT 1000.350 3368.530 1000.650 3368.910 ;
        RECT 1049.110 3368.910 1097.250 3369.210 ;
        RECT 1000.350 3368.230 1048.490 3368.530 ;
        RECT 758.390 3367.550 759.610 3367.850 ;
        RECT 811.045 3367.850 811.375 3367.865 ;
        RECT 834.505 3367.850 834.835 3367.865 ;
        RECT 811.045 3367.550 834.835 3367.850 ;
        RECT 1048.190 3367.850 1048.490 3368.230 ;
        RECT 1049.110 3367.850 1049.410 3368.910 ;
        RECT 1096.950 3368.530 1097.250 3368.910 ;
        RECT 1145.710 3368.910 1193.850 3369.210 ;
        RECT 1096.950 3368.230 1145.090 3368.530 ;
        RECT 1048.190 3367.550 1049.410 3367.850 ;
        RECT 1144.790 3367.850 1145.090 3368.230 ;
        RECT 1145.710 3367.850 1146.010 3368.910 ;
        RECT 1193.550 3368.530 1193.850 3368.910 ;
        RECT 1242.310 3368.910 1290.450 3369.210 ;
        RECT 1193.550 3368.230 1241.690 3368.530 ;
        RECT 1144.790 3367.550 1146.010 3367.850 ;
        RECT 1241.390 3367.850 1241.690 3368.230 ;
        RECT 1242.310 3367.850 1242.610 3368.910 ;
        RECT 1290.150 3368.530 1290.450 3368.910 ;
        RECT 1338.910 3368.910 1387.050 3369.210 ;
        RECT 1290.150 3368.230 1338.290 3368.530 ;
        RECT 1241.390 3367.550 1242.610 3367.850 ;
        RECT 1337.990 3367.850 1338.290 3368.230 ;
        RECT 1338.910 3367.850 1339.210 3368.910 ;
        RECT 1386.750 3368.530 1387.050 3368.910 ;
        RECT 1435.510 3368.910 1449.395 3369.210 ;
        RECT 1386.750 3368.230 1434.890 3368.530 ;
        RECT 1337.990 3367.550 1339.210 3367.850 ;
        RECT 1434.590 3367.850 1434.890 3368.230 ;
        RECT 1435.510 3367.850 1435.810 3368.910 ;
        RECT 1449.065 3368.895 1449.395 3368.910 ;
        RECT 1497.110 3369.210 1497.490 3369.220 ;
        RECT 1738.865 3369.210 1739.195 3369.225 ;
        RECT 1497.110 3368.910 1580.250 3369.210 ;
        RECT 1497.110 3368.900 1497.490 3368.910 ;
        RECT 1579.950 3368.530 1580.250 3368.910 ;
        RECT 1628.710 3368.910 1676.850 3369.210 ;
        RECT 1579.950 3368.230 1628.090 3368.530 ;
        RECT 1434.590 3367.550 1435.810 3367.850 ;
        RECT 1463.325 3367.850 1463.655 3367.865 ;
        RECT 1497.110 3367.850 1497.490 3367.860 ;
        RECT 1463.325 3367.550 1497.490 3367.850 ;
        RECT 1627.790 3367.850 1628.090 3368.230 ;
        RECT 1628.710 3367.850 1629.010 3368.910 ;
        RECT 1676.550 3368.530 1676.850 3368.910 ;
        RECT 1725.310 3368.910 1739.195 3369.210 ;
        RECT 1676.550 3368.230 1724.690 3368.530 ;
        RECT 1627.790 3367.550 1629.010 3367.850 ;
        RECT 1724.390 3367.850 1724.690 3368.230 ;
        RECT 1725.310 3367.850 1725.610 3368.910 ;
        RECT 1738.865 3368.895 1739.195 3368.910 ;
        RECT 1859.845 3369.210 1860.175 3369.225 ;
        RECT 1883.510 3369.210 1883.890 3369.220 ;
        RECT 1859.845 3368.910 1883.890 3369.210 ;
        RECT 1859.845 3368.895 1860.175 3368.910 ;
        RECT 1883.510 3368.900 1883.890 3368.910 ;
        RECT 1897.565 3369.210 1897.895 3369.225 ;
        RECT 2704.865 3369.210 2705.195 3369.225 ;
        RECT 1897.565 3368.910 1966.650 3369.210 ;
        RECT 1897.565 3368.895 1897.895 3368.910 ;
        RECT 1966.350 3368.530 1966.650 3368.910 ;
        RECT 2015.110 3368.910 2063.250 3369.210 ;
        RECT 1966.350 3368.230 2014.490 3368.530 ;
        RECT 1724.390 3367.550 1725.610 3367.850 ;
        RECT 1777.045 3367.850 1777.375 3367.865 ;
        RECT 1786.910 3367.850 1787.290 3367.860 ;
        RECT 1777.045 3367.550 1787.290 3367.850 ;
        RECT 2014.190 3367.850 2014.490 3368.230 ;
        RECT 2015.110 3367.850 2015.410 3368.910 ;
        RECT 2062.950 3368.530 2063.250 3368.910 ;
        RECT 2159.550 3368.910 2207.690 3369.210 ;
        RECT 2062.950 3368.230 2111.090 3368.530 ;
        RECT 2014.190 3367.550 2015.410 3367.850 ;
        RECT 2110.790 3367.850 2111.090 3368.230 ;
        RECT 2159.550 3367.850 2159.850 3368.910 ;
        RECT 2110.790 3367.550 2159.850 3367.850 ;
        RECT 2207.390 3367.850 2207.690 3368.910 ;
        RECT 2208.310 3368.910 2256.450 3369.210 ;
        RECT 2208.310 3367.850 2208.610 3368.910 ;
        RECT 2256.150 3368.530 2256.450 3368.910 ;
        RECT 2304.910 3368.910 2353.050 3369.210 ;
        RECT 2256.150 3368.230 2304.290 3368.530 ;
        RECT 2207.390 3367.550 2208.610 3367.850 ;
        RECT 2303.990 3367.850 2304.290 3368.230 ;
        RECT 2304.910 3367.850 2305.210 3368.910 ;
        RECT 2352.750 3368.530 2353.050 3368.910 ;
        RECT 2401.510 3368.910 2449.650 3369.210 ;
        RECT 2352.750 3368.230 2400.890 3368.530 ;
        RECT 2303.990 3367.550 2305.210 3367.850 ;
        RECT 2400.590 3367.850 2400.890 3368.230 ;
        RECT 2401.510 3367.850 2401.810 3368.910 ;
        RECT 2449.350 3368.530 2449.650 3368.910 ;
        RECT 2498.110 3368.910 2546.250 3369.210 ;
        RECT 2449.350 3368.230 2497.490 3368.530 ;
        RECT 2400.590 3367.550 2401.810 3367.850 ;
        RECT 2497.190 3367.850 2497.490 3368.230 ;
        RECT 2498.110 3367.850 2498.410 3368.910 ;
        RECT 2545.950 3368.530 2546.250 3368.910 ;
        RECT 2594.710 3368.910 2642.850 3369.210 ;
        RECT 2545.950 3368.230 2594.090 3368.530 ;
        RECT 2497.190 3367.550 2498.410 3367.850 ;
        RECT 2593.790 3367.850 2594.090 3368.230 ;
        RECT 2594.710 3367.850 2595.010 3368.910 ;
        RECT 2642.550 3368.530 2642.850 3368.910 ;
        RECT 2691.310 3368.910 2705.195 3369.210 ;
        RECT 2642.550 3368.230 2690.690 3368.530 ;
        RECT 2593.790 3367.550 2595.010 3367.850 ;
        RECT 2690.390 3367.850 2690.690 3368.230 ;
        RECT 2691.310 3367.850 2691.610 3368.910 ;
        RECT 2704.865 3368.895 2705.195 3368.910 ;
        RECT 2825.845 3369.210 2826.175 3369.225 ;
        RECT 2863.565 3369.210 2863.895 3369.225 ;
        RECT 2825.845 3368.910 2849.850 3369.210 ;
        RECT 2825.845 3368.895 2826.175 3368.910 ;
        RECT 2849.550 3368.530 2849.850 3368.910 ;
        RECT 2863.565 3368.910 2884.810 3369.210 ;
        RECT 2863.565 3368.895 2863.895 3368.910 ;
        RECT 2863.105 3368.530 2863.435 3368.545 ;
        RECT 2849.550 3368.230 2863.435 3368.530 ;
        RECT 2884.510 3368.530 2884.810 3368.910 ;
        RECT 2916.710 3368.530 2917.010 3372.990 ;
        RECT 2917.600 3372.540 2924.800 3372.990 ;
        RECT 2884.510 3368.230 2917.010 3368.530 ;
        RECT 2863.105 3368.215 2863.435 3368.230 ;
        RECT 2690.390 3367.550 2691.610 3367.850 ;
        RECT 2743.045 3367.850 2743.375 3367.865 ;
        RECT 2766.505 3367.850 2766.835 3367.865 ;
        RECT 2743.045 3367.550 2766.835 3367.850 ;
        RECT 811.045 3367.535 811.375 3367.550 ;
        RECT 834.505 3367.535 834.835 3367.550 ;
        RECT 1463.325 3367.535 1463.655 3367.550 ;
        RECT 1497.110 3367.540 1497.490 3367.550 ;
        RECT 1777.045 3367.535 1777.375 3367.550 ;
        RECT 1786.910 3367.540 1787.290 3367.550 ;
        RECT 2743.045 3367.535 2743.375 3367.550 ;
        RECT 2766.505 3367.535 2766.835 3367.550 ;
        RECT 290.990 1947.330 291.370 1947.340 ;
        RECT 300.000 1947.330 304.000 1947.400 ;
        RECT 290.990 1947.030 304.000 1947.330 ;
        RECT 290.990 1947.020 291.370 1947.030 ;
        RECT 300.000 1946.800 304.000 1947.030 ;
      LAYER via3 ;
        RECT 917.540 3370.260 917.860 3370.580 ;
        RECT 1883.540 3370.260 1883.860 3370.580 ;
        RECT 1786.940 3369.580 1787.260 3369.900 ;
        RECT 291.020 3368.900 291.340 3369.220 ;
        RECT 917.540 3368.900 917.860 3369.220 ;
        RECT 1497.140 3368.900 1497.460 3369.220 ;
        RECT 1497.140 3367.540 1497.460 3367.860 ;
        RECT 1883.540 3368.900 1883.860 3369.220 ;
        RECT 1786.940 3367.540 1787.260 3367.860 ;
        RECT 291.020 1947.020 291.340 1947.340 ;
      LAYER met4 ;
        RECT 917.535 3370.255 917.865 3370.585 ;
        RECT 1883.535 3370.255 1883.865 3370.585 ;
        RECT 917.550 3369.225 917.850 3370.255 ;
        RECT 1786.935 3369.575 1787.265 3369.905 ;
        RECT 291.015 3368.895 291.345 3369.225 ;
        RECT 917.535 3368.895 917.865 3369.225 ;
        RECT 1497.135 3368.895 1497.465 3369.225 ;
        RECT 291.030 1947.345 291.330 3368.895 ;
        RECT 1497.150 3367.865 1497.450 3368.895 ;
        RECT 1786.950 3367.865 1787.250 3369.575 ;
        RECT 1883.550 3369.225 1883.850 3370.255 ;
        RECT 1883.535 3368.895 1883.865 3369.225 ;
        RECT 1497.135 3367.535 1497.465 3367.865 ;
        RECT 1786.935 3367.535 1787.265 3367.865 ;
        RECT 291.015 1947.015 291.345 1947.345 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2795.030 3422.680 2795.350 3422.740 ;
        RECT 2798.250 3422.680 2798.570 3422.740 ;
        RECT 2795.030 3422.540 2798.570 3422.680 ;
        RECT 2795.030 3422.480 2795.350 3422.540 ;
        RECT 2798.250 3422.480 2798.570 3422.540 ;
        RECT 2795.030 3374.400 2795.350 3374.460 ;
        RECT 2796.870 3374.400 2797.190 3374.460 ;
        RECT 2795.030 3374.260 2797.190 3374.400 ;
        RECT 2795.030 3374.200 2795.350 3374.260 ;
        RECT 2796.870 3374.200 2797.190 3374.260 ;
        RECT 2795.490 3308.780 2795.810 3308.840 ;
        RECT 2796.870 3308.780 2797.190 3308.840 ;
        RECT 2795.490 3308.640 2797.190 3308.780 ;
        RECT 2795.490 3308.580 2795.810 3308.640 ;
        RECT 2796.870 3308.580 2797.190 3308.640 ;
        RECT 2795.490 3284.640 2795.810 3284.700 ;
        RECT 2795.950 3284.640 2796.270 3284.700 ;
        RECT 2795.490 3284.500 2796.270 3284.640 ;
        RECT 2795.490 3284.440 2795.810 3284.500 ;
        RECT 2795.950 3284.440 2796.270 3284.500 ;
        RECT 2795.490 3236.360 2795.810 3236.420 ;
        RECT 2795.950 3236.360 2796.270 3236.420 ;
        RECT 2795.490 3236.220 2796.270 3236.360 ;
        RECT 2795.490 3236.160 2795.810 3236.220 ;
        RECT 2795.950 3236.160 2796.270 3236.220 ;
        RECT 2795.490 3202.020 2795.810 3202.080 ;
        RECT 2795.950 3202.020 2796.270 3202.080 ;
        RECT 2795.490 3201.880 2796.270 3202.020 ;
        RECT 2795.490 3201.820 2795.810 3201.880 ;
        RECT 2795.950 3201.820 2796.270 3201.880 ;
        RECT 2795.030 3153.400 2795.350 3153.460 ;
        RECT 2795.950 3153.400 2796.270 3153.460 ;
        RECT 2795.030 3153.260 2796.270 3153.400 ;
        RECT 2795.030 3153.200 2795.350 3153.260 ;
        RECT 2795.950 3153.200 2796.270 3153.260 ;
        RECT 2795.030 3056.840 2795.350 3056.900 ;
        RECT 2795.950 3056.840 2796.270 3056.900 ;
        RECT 2795.030 3056.700 2796.270 3056.840 ;
        RECT 2795.030 3056.640 2795.350 3056.700 ;
        RECT 2795.950 3056.640 2796.270 3056.700 ;
        RECT 2795.030 3042.900 2795.350 3042.960 ;
        RECT 2795.490 3042.900 2795.810 3042.960 ;
        RECT 2795.030 3042.760 2795.810 3042.900 ;
        RECT 2795.030 3042.700 2795.350 3042.760 ;
        RECT 2795.490 3042.700 2795.810 3042.760 ;
        RECT 2795.030 3008.560 2795.350 3008.620 ;
        RECT 2796.410 3008.560 2796.730 3008.620 ;
        RECT 2795.030 3008.420 2796.730 3008.560 ;
        RECT 2795.030 3008.360 2795.350 3008.420 ;
        RECT 2796.410 3008.360 2796.730 3008.420 ;
        RECT 2795.490 2994.620 2795.810 2994.680 ;
        RECT 2796.410 2994.620 2796.730 2994.680 ;
        RECT 2795.490 2994.480 2796.730 2994.620 ;
        RECT 2795.490 2994.420 2795.810 2994.480 ;
        RECT 2796.410 2994.420 2796.730 2994.480 ;
        RECT 2795.490 2946.680 2795.810 2946.740 ;
        RECT 2796.870 2946.680 2797.190 2946.740 ;
        RECT 2795.490 2946.540 2797.190 2946.680 ;
        RECT 2795.490 2946.480 2795.810 2946.540 ;
        RECT 2796.870 2946.480 2797.190 2946.540 ;
        RECT 2796.870 2912.340 2797.190 2912.400 ;
        RECT 2796.500 2912.200 2797.190 2912.340 ;
        RECT 2796.500 2911.720 2796.640 2912.200 ;
        RECT 2796.870 2912.140 2797.190 2912.200 ;
        RECT 2796.410 2911.460 2796.730 2911.720 ;
        RECT 2795.030 2801.500 2795.350 2801.560 ;
        RECT 2795.490 2801.500 2795.810 2801.560 ;
        RECT 2795.030 2801.360 2795.810 2801.500 ;
        RECT 2795.030 2801.300 2795.350 2801.360 ;
        RECT 2795.490 2801.300 2795.810 2801.360 ;
        RECT 298.150 2695.420 298.470 2695.480 ;
        RECT 2795.950 2695.420 2796.270 2695.480 ;
        RECT 298.150 2695.280 2796.270 2695.420 ;
        RECT 298.150 2695.220 298.470 2695.280 ;
        RECT 2795.950 2695.220 2796.270 2695.280 ;
      LAYER via ;
        RECT 2795.060 3422.480 2795.320 3422.740 ;
        RECT 2798.280 3422.480 2798.540 3422.740 ;
        RECT 2795.060 3374.200 2795.320 3374.460 ;
        RECT 2796.900 3374.200 2797.160 3374.460 ;
        RECT 2795.520 3308.580 2795.780 3308.840 ;
        RECT 2796.900 3308.580 2797.160 3308.840 ;
        RECT 2795.520 3284.440 2795.780 3284.700 ;
        RECT 2795.980 3284.440 2796.240 3284.700 ;
        RECT 2795.520 3236.160 2795.780 3236.420 ;
        RECT 2795.980 3236.160 2796.240 3236.420 ;
        RECT 2795.520 3201.820 2795.780 3202.080 ;
        RECT 2795.980 3201.820 2796.240 3202.080 ;
        RECT 2795.060 3153.200 2795.320 3153.460 ;
        RECT 2795.980 3153.200 2796.240 3153.460 ;
        RECT 2795.060 3056.640 2795.320 3056.900 ;
        RECT 2795.980 3056.640 2796.240 3056.900 ;
        RECT 2795.060 3042.700 2795.320 3042.960 ;
        RECT 2795.520 3042.700 2795.780 3042.960 ;
        RECT 2795.060 3008.360 2795.320 3008.620 ;
        RECT 2796.440 3008.360 2796.700 3008.620 ;
        RECT 2795.520 2994.420 2795.780 2994.680 ;
        RECT 2796.440 2994.420 2796.700 2994.680 ;
        RECT 2795.520 2946.480 2795.780 2946.740 ;
        RECT 2796.900 2946.480 2797.160 2946.740 ;
        RECT 2796.900 2912.140 2797.160 2912.400 ;
        RECT 2796.440 2911.460 2796.700 2911.720 ;
        RECT 2795.060 2801.300 2795.320 2801.560 ;
        RECT 2795.520 2801.300 2795.780 2801.560 ;
        RECT 298.180 2695.220 298.440 2695.480 ;
        RECT 2795.980 2695.220 2796.240 2695.480 ;
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
        RECT 2798.340 3422.770 2798.480 3517.600 ;
        RECT 2795.060 3422.450 2795.320 3422.770 ;
        RECT 2798.280 3422.450 2798.540 3422.770 ;
        RECT 2795.120 3422.285 2795.260 3422.450 ;
        RECT 2795.050 3421.915 2795.330 3422.285 ;
        RECT 2795.050 3421.235 2795.330 3421.605 ;
        RECT 2795.120 3374.490 2795.260 3421.235 ;
        RECT 2795.060 3374.170 2795.320 3374.490 ;
        RECT 2796.900 3374.170 2797.160 3374.490 ;
        RECT 2796.960 3308.870 2797.100 3374.170 ;
        RECT 2795.520 3308.550 2795.780 3308.870 ;
        RECT 2796.900 3308.550 2797.160 3308.870 ;
        RECT 2795.580 3284.730 2795.720 3308.550 ;
        RECT 2795.520 3284.410 2795.780 3284.730 ;
        RECT 2795.980 3284.410 2796.240 3284.730 ;
        RECT 2796.040 3236.450 2796.180 3284.410 ;
        RECT 2795.520 3236.130 2795.780 3236.450 ;
        RECT 2795.980 3236.130 2796.240 3236.450 ;
        RECT 2795.580 3202.110 2795.720 3236.130 ;
        RECT 2795.520 3201.790 2795.780 3202.110 ;
        RECT 2795.980 3201.790 2796.240 3202.110 ;
        RECT 2796.040 3153.490 2796.180 3201.790 ;
        RECT 2795.060 3153.170 2795.320 3153.490 ;
        RECT 2795.980 3153.170 2796.240 3153.490 ;
        RECT 2795.120 3152.890 2795.260 3153.170 ;
        RECT 2795.120 3152.750 2795.720 3152.890 ;
        RECT 2795.580 3105.290 2795.720 3152.750 ;
        RECT 2795.580 3105.150 2796.180 3105.290 ;
        RECT 2796.040 3056.930 2796.180 3105.150 ;
        RECT 2795.060 3056.610 2795.320 3056.930 ;
        RECT 2795.980 3056.610 2796.240 3056.930 ;
        RECT 2795.120 3056.330 2795.260 3056.610 ;
        RECT 2795.120 3056.190 2795.720 3056.330 ;
        RECT 2795.580 3042.990 2795.720 3056.190 ;
        RECT 2795.060 3042.670 2795.320 3042.990 ;
        RECT 2795.520 3042.670 2795.780 3042.990 ;
        RECT 2795.120 3008.650 2795.260 3042.670 ;
        RECT 2795.060 3008.330 2795.320 3008.650 ;
        RECT 2796.440 3008.330 2796.700 3008.650 ;
        RECT 2796.500 2994.710 2796.640 3008.330 ;
        RECT 2795.520 2994.390 2795.780 2994.710 ;
        RECT 2796.440 2994.390 2796.700 2994.710 ;
        RECT 2795.580 2946.770 2795.720 2994.390 ;
        RECT 2795.520 2946.450 2795.780 2946.770 ;
        RECT 2796.900 2946.450 2797.160 2946.770 ;
        RECT 2796.960 2912.430 2797.100 2946.450 ;
        RECT 2796.900 2912.110 2797.160 2912.430 ;
        RECT 2796.440 2911.430 2796.700 2911.750 ;
        RECT 2796.500 2863.210 2796.640 2911.430 ;
        RECT 2795.580 2863.070 2796.640 2863.210 ;
        RECT 2795.580 2801.590 2795.720 2863.070 ;
        RECT 2795.060 2801.270 2795.320 2801.590 ;
        RECT 2795.520 2801.270 2795.780 2801.590 ;
        RECT 2795.120 2766.650 2795.260 2801.270 ;
        RECT 2795.120 2766.510 2795.720 2766.650 ;
        RECT 2795.580 2719.050 2795.720 2766.510 ;
        RECT 2795.580 2718.910 2796.180 2719.050 ;
        RECT 2796.040 2695.510 2796.180 2718.910 ;
        RECT 298.180 2695.190 298.440 2695.510 ;
        RECT 2795.980 2695.190 2796.240 2695.510 ;
        RECT 298.240 1978.645 298.380 2695.190 ;
        RECT 298.170 1978.275 298.450 1978.645 ;
      LAYER via2 ;
        RECT 2795.050 3421.960 2795.330 3422.240 ;
        RECT 2795.050 3421.280 2795.330 3421.560 ;
        RECT 298.170 1978.320 298.450 1978.600 ;
      LAYER met3 ;
        RECT 2795.025 3421.935 2795.355 3422.265 ;
        RECT 2795.040 3421.585 2795.340 3421.935 ;
        RECT 2795.025 3421.255 2795.355 3421.585 ;
        RECT 298.145 1978.610 298.475 1978.625 ;
        RECT 300.000 1978.610 304.000 1978.680 ;
        RECT 298.145 1978.310 304.000 1978.610 ;
        RECT 298.145 1978.295 298.475 1978.310 ;
        RECT 300.000 1978.080 304.000 1978.310 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2470.270 3464.160 2470.590 3464.220 ;
        RECT 2474.410 3464.160 2474.730 3464.220 ;
        RECT 2470.270 3464.020 2474.730 3464.160 ;
        RECT 2470.270 3463.960 2470.590 3464.020 ;
        RECT 2474.410 3463.960 2474.730 3464.020 ;
        RECT 2470.270 3367.600 2470.590 3367.660 ;
        RECT 2471.190 3367.600 2471.510 3367.660 ;
        RECT 2470.270 3367.460 2471.510 3367.600 ;
        RECT 2470.270 3367.400 2470.590 3367.460 ;
        RECT 2471.190 3367.400 2471.510 3367.460 ;
        RECT 2470.270 3270.700 2470.590 3270.760 ;
        RECT 2471.190 3270.700 2471.510 3270.760 ;
        RECT 2470.270 3270.560 2471.510 3270.700 ;
        RECT 2470.270 3270.500 2470.590 3270.560 ;
        RECT 2471.190 3270.500 2471.510 3270.560 ;
        RECT 297.230 3253.360 297.550 3253.420 ;
        RECT 2470.270 3253.360 2470.590 3253.420 ;
        RECT 297.230 3253.220 2470.590 3253.360 ;
        RECT 297.230 3253.160 297.550 3253.220 ;
        RECT 2470.270 3253.160 2470.590 3253.220 ;
      LAYER via ;
        RECT 2470.300 3463.960 2470.560 3464.220 ;
        RECT 2474.440 3463.960 2474.700 3464.220 ;
        RECT 2470.300 3367.400 2470.560 3367.660 ;
        RECT 2471.220 3367.400 2471.480 3367.660 ;
        RECT 2470.300 3270.500 2470.560 3270.760 ;
        RECT 2471.220 3270.500 2471.480 3270.760 ;
        RECT 297.260 3253.160 297.520 3253.420 ;
        RECT 2470.300 3253.160 2470.560 3253.420 ;
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
        RECT 2474.040 3517.370 2474.180 3517.600 ;
        RECT 2474.040 3517.230 2474.640 3517.370 ;
        RECT 2474.500 3464.250 2474.640 3517.230 ;
        RECT 2470.300 3463.930 2470.560 3464.250 ;
        RECT 2474.440 3463.930 2474.700 3464.250 ;
        RECT 2470.360 3415.370 2470.500 3463.930 ;
        RECT 2470.360 3415.230 2471.420 3415.370 ;
        RECT 2471.280 3367.690 2471.420 3415.230 ;
        RECT 2470.300 3367.370 2470.560 3367.690 ;
        RECT 2471.220 3367.370 2471.480 3367.690 ;
        RECT 2470.360 3318.810 2470.500 3367.370 ;
        RECT 2470.360 3318.670 2471.420 3318.810 ;
        RECT 2471.280 3270.790 2471.420 3318.670 ;
        RECT 2470.300 3270.470 2470.560 3270.790 ;
        RECT 2471.220 3270.470 2471.480 3270.790 ;
        RECT 2470.360 3253.450 2470.500 3270.470 ;
        RECT 297.260 3253.130 297.520 3253.450 ;
        RECT 2470.300 3253.130 2470.560 3253.450 ;
        RECT 297.320 2010.605 297.460 3253.130 ;
        RECT 297.250 2010.235 297.530 2010.605 ;
      LAYER via2 ;
        RECT 297.250 2010.280 297.530 2010.560 ;
      LAYER met3 ;
        RECT 297.225 2010.570 297.555 2010.585 ;
        RECT 300.000 2010.570 304.000 2010.640 ;
        RECT 297.225 2010.270 304.000 2010.570 ;
        RECT 297.225 2010.255 297.555 2010.270 ;
        RECT 300.000 2010.040 304.000 2010.270 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2145.970 3464.160 2146.290 3464.220 ;
        RECT 2149.650 3464.160 2149.970 3464.220 ;
        RECT 2145.970 3464.020 2149.970 3464.160 ;
        RECT 2145.970 3463.960 2146.290 3464.020 ;
        RECT 2149.650 3463.960 2149.970 3464.020 ;
        RECT 2145.970 3380.860 2146.290 3380.920 ;
        RECT 2146.430 3380.860 2146.750 3380.920 ;
        RECT 2145.970 3380.720 2146.750 3380.860 ;
        RECT 2145.970 3380.660 2146.290 3380.720 ;
        RECT 2146.430 3380.660 2146.750 3380.720 ;
        RECT 2146.430 3332.920 2146.750 3332.980 ;
        RECT 2146.890 3332.920 2147.210 3332.980 ;
        RECT 2146.430 3332.780 2147.210 3332.920 ;
        RECT 2146.430 3332.720 2146.750 3332.780 ;
        RECT 2146.890 3332.720 2147.210 3332.780 ;
        RECT 2146.890 3298.580 2147.210 3298.640 ;
        RECT 2146.520 3298.440 2147.210 3298.580 ;
        RECT 2146.520 3298.300 2146.660 3298.440 ;
        RECT 2146.890 3298.380 2147.210 3298.440 ;
        RECT 2146.430 3298.040 2146.750 3298.300 ;
        RECT 2146.430 3249.960 2146.750 3250.020 ;
        RECT 2147.350 3249.960 2147.670 3250.020 ;
        RECT 2146.430 3249.820 2147.670 3249.960 ;
        RECT 2146.430 3249.760 2146.750 3249.820 ;
        RECT 2147.350 3249.760 2147.670 3249.820 ;
        RECT 2145.970 3187.740 2146.290 3187.800 ;
        RECT 2146.890 3187.740 2147.210 3187.800 ;
        RECT 2145.970 3187.600 2147.210 3187.740 ;
        RECT 2145.970 3187.540 2146.290 3187.600 ;
        RECT 2146.890 3187.540 2147.210 3187.600 ;
        RECT 2145.970 3139.800 2146.290 3139.860 ;
        RECT 2147.810 3139.800 2148.130 3139.860 ;
        RECT 2145.970 3139.660 2148.130 3139.800 ;
        RECT 2145.970 3139.600 2146.290 3139.660 ;
        RECT 2147.810 3139.600 2148.130 3139.660 ;
        RECT 2147.810 3105.460 2148.130 3105.520 ;
        RECT 2147.440 3105.320 2148.130 3105.460 ;
        RECT 2147.440 3104.840 2147.580 3105.320 ;
        RECT 2147.810 3105.260 2148.130 3105.320 ;
        RECT 2147.350 3104.580 2147.670 3104.840 ;
        RECT 2146.430 3056.840 2146.750 3056.900 ;
        RECT 2147.350 3056.840 2147.670 3056.900 ;
        RECT 2146.430 3056.700 2147.670 3056.840 ;
        RECT 2146.430 3056.640 2146.750 3056.700 ;
        RECT 2147.350 3056.640 2147.670 3056.700 ;
        RECT 2146.430 3042.900 2146.750 3042.960 ;
        RECT 2146.890 3042.900 2147.210 3042.960 ;
        RECT 2146.430 3042.760 2147.210 3042.900 ;
        RECT 2146.430 3042.700 2146.750 3042.760 ;
        RECT 2146.890 3042.700 2147.210 3042.760 ;
        RECT 2146.430 3008.560 2146.750 3008.620 ;
        RECT 2147.810 3008.560 2148.130 3008.620 ;
        RECT 2146.430 3008.420 2148.130 3008.560 ;
        RECT 2146.430 3008.360 2146.750 3008.420 ;
        RECT 2147.810 3008.360 2148.130 3008.420 ;
        RECT 2146.890 2994.620 2147.210 2994.680 ;
        RECT 2147.810 2994.620 2148.130 2994.680 ;
        RECT 2146.890 2994.480 2148.130 2994.620 ;
        RECT 2146.890 2994.420 2147.210 2994.480 ;
        RECT 2147.810 2994.420 2148.130 2994.480 ;
        RECT 2146.890 2946.680 2147.210 2946.740 ;
        RECT 2148.270 2946.680 2148.590 2946.740 ;
        RECT 2146.890 2946.540 2148.590 2946.680 ;
        RECT 2146.890 2946.480 2147.210 2946.540 ;
        RECT 2148.270 2946.480 2148.590 2946.540 ;
        RECT 2148.270 2912.340 2148.590 2912.400 ;
        RECT 2147.900 2912.200 2148.590 2912.340 ;
        RECT 2147.900 2911.720 2148.040 2912.200 ;
        RECT 2148.270 2912.140 2148.590 2912.200 ;
        RECT 2147.810 2911.460 2148.130 2911.720 ;
        RECT 298.610 2695.760 298.930 2695.820 ;
        RECT 2147.350 2695.760 2147.670 2695.820 ;
        RECT 298.610 2695.620 2147.670 2695.760 ;
        RECT 298.610 2695.560 298.930 2695.620 ;
        RECT 2147.350 2695.560 2147.670 2695.620 ;
      LAYER via ;
        RECT 2146.000 3463.960 2146.260 3464.220 ;
        RECT 2149.680 3463.960 2149.940 3464.220 ;
        RECT 2146.000 3380.660 2146.260 3380.920 ;
        RECT 2146.460 3380.660 2146.720 3380.920 ;
        RECT 2146.460 3332.720 2146.720 3332.980 ;
        RECT 2146.920 3332.720 2147.180 3332.980 ;
        RECT 2146.920 3298.380 2147.180 3298.640 ;
        RECT 2146.460 3298.040 2146.720 3298.300 ;
        RECT 2146.460 3249.760 2146.720 3250.020 ;
        RECT 2147.380 3249.760 2147.640 3250.020 ;
        RECT 2146.000 3187.540 2146.260 3187.800 ;
        RECT 2146.920 3187.540 2147.180 3187.800 ;
        RECT 2146.000 3139.600 2146.260 3139.860 ;
        RECT 2147.840 3139.600 2148.100 3139.860 ;
        RECT 2147.840 3105.260 2148.100 3105.520 ;
        RECT 2147.380 3104.580 2147.640 3104.840 ;
        RECT 2146.460 3056.640 2146.720 3056.900 ;
        RECT 2147.380 3056.640 2147.640 3056.900 ;
        RECT 2146.460 3042.700 2146.720 3042.960 ;
        RECT 2146.920 3042.700 2147.180 3042.960 ;
        RECT 2146.460 3008.360 2146.720 3008.620 ;
        RECT 2147.840 3008.360 2148.100 3008.620 ;
        RECT 2146.920 2994.420 2147.180 2994.680 ;
        RECT 2147.840 2994.420 2148.100 2994.680 ;
        RECT 2146.920 2946.480 2147.180 2946.740 ;
        RECT 2148.300 2946.480 2148.560 2946.740 ;
        RECT 2148.300 2912.140 2148.560 2912.400 ;
        RECT 2147.840 2911.460 2148.100 2911.720 ;
        RECT 298.640 2695.560 298.900 2695.820 ;
        RECT 2147.380 2695.560 2147.640 2695.820 ;
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
        RECT 2149.280 3517.370 2149.420 3517.600 ;
        RECT 2149.280 3517.230 2149.880 3517.370 ;
        RECT 2149.740 3464.250 2149.880 3517.230 ;
        RECT 2146.000 3463.930 2146.260 3464.250 ;
        RECT 2149.680 3463.930 2149.940 3464.250 ;
        RECT 2146.060 3380.950 2146.200 3463.930 ;
        RECT 2146.000 3380.630 2146.260 3380.950 ;
        RECT 2146.460 3380.630 2146.720 3380.950 ;
        RECT 2146.520 3333.010 2146.660 3380.630 ;
        RECT 2146.460 3332.690 2146.720 3333.010 ;
        RECT 2146.920 3332.690 2147.180 3333.010 ;
        RECT 2146.980 3298.670 2147.120 3332.690 ;
        RECT 2146.920 3298.350 2147.180 3298.670 ;
        RECT 2146.460 3298.010 2146.720 3298.330 ;
        RECT 2146.520 3250.050 2146.660 3298.010 ;
        RECT 2146.460 3249.730 2146.720 3250.050 ;
        RECT 2147.380 3249.730 2147.640 3250.050 ;
        RECT 2147.440 3212.050 2147.580 3249.730 ;
        RECT 2146.520 3211.910 2147.580 3212.050 ;
        RECT 2146.520 3188.250 2146.660 3211.910 ;
        RECT 2146.520 3188.110 2147.120 3188.250 ;
        RECT 2146.980 3187.830 2147.120 3188.110 ;
        RECT 2146.000 3187.510 2146.260 3187.830 ;
        RECT 2146.920 3187.510 2147.180 3187.830 ;
        RECT 2146.060 3139.890 2146.200 3187.510 ;
        RECT 2146.000 3139.570 2146.260 3139.890 ;
        RECT 2147.840 3139.570 2148.100 3139.890 ;
        RECT 2147.900 3105.550 2148.040 3139.570 ;
        RECT 2147.840 3105.230 2148.100 3105.550 ;
        RECT 2147.380 3104.550 2147.640 3104.870 ;
        RECT 2147.440 3056.930 2147.580 3104.550 ;
        RECT 2146.460 3056.610 2146.720 3056.930 ;
        RECT 2147.380 3056.610 2147.640 3056.930 ;
        RECT 2146.520 3056.330 2146.660 3056.610 ;
        RECT 2146.520 3056.190 2147.120 3056.330 ;
        RECT 2146.980 3042.990 2147.120 3056.190 ;
        RECT 2146.460 3042.670 2146.720 3042.990 ;
        RECT 2146.920 3042.670 2147.180 3042.990 ;
        RECT 2146.520 3008.650 2146.660 3042.670 ;
        RECT 2146.460 3008.330 2146.720 3008.650 ;
        RECT 2147.840 3008.330 2148.100 3008.650 ;
        RECT 2147.900 2994.710 2148.040 3008.330 ;
        RECT 2146.920 2994.390 2147.180 2994.710 ;
        RECT 2147.840 2994.390 2148.100 2994.710 ;
        RECT 2146.980 2946.770 2147.120 2994.390 ;
        RECT 2146.920 2946.450 2147.180 2946.770 ;
        RECT 2148.300 2946.450 2148.560 2946.770 ;
        RECT 2148.360 2912.430 2148.500 2946.450 ;
        RECT 2148.300 2912.110 2148.560 2912.430 ;
        RECT 2147.840 2911.430 2148.100 2911.750 ;
        RECT 2147.900 2863.210 2148.040 2911.430 ;
        RECT 2146.980 2863.070 2148.040 2863.210 ;
        RECT 2146.980 2815.610 2147.120 2863.070 ;
        RECT 2146.520 2815.470 2147.120 2815.610 ;
        RECT 2146.520 2814.930 2146.660 2815.470 ;
        RECT 2146.520 2814.790 2147.120 2814.930 ;
        RECT 2146.980 2767.330 2147.120 2814.790 ;
        RECT 2146.980 2767.190 2147.580 2767.330 ;
        RECT 2147.440 2695.850 2147.580 2767.190 ;
        RECT 298.640 2695.530 298.900 2695.850 ;
        RECT 2147.380 2695.530 2147.640 2695.850 ;
        RECT 298.700 2041.885 298.840 2695.530 ;
        RECT 298.630 2041.515 298.910 2041.885 ;
      LAYER via2 ;
        RECT 298.630 2041.560 298.910 2041.840 ;
      LAYER met3 ;
        RECT 298.605 2041.850 298.935 2041.865 ;
        RECT 300.000 2041.850 304.000 2041.920 ;
        RECT 298.605 2041.550 304.000 2041.850 ;
        RECT 298.605 2041.535 298.935 2041.550 ;
        RECT 300.000 2041.320 304.000 2041.550 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1822.130 3491.360 1822.450 3491.420 ;
        RECT 1825.350 3491.360 1825.670 3491.420 ;
        RECT 1822.130 3491.220 1825.670 3491.360 ;
        RECT 1822.130 3491.160 1822.450 3491.220 ;
        RECT 1825.350 3491.160 1825.670 3491.220 ;
        RECT 1822.130 3347.000 1822.450 3347.260 ;
        RECT 1822.220 3346.580 1822.360 3347.000 ;
        RECT 1822.130 3346.320 1822.450 3346.580 ;
        RECT 1821.670 3270.700 1821.990 3270.760 ;
        RECT 1822.590 3270.700 1822.910 3270.760 ;
        RECT 1821.670 3270.560 1822.910 3270.700 ;
        RECT 1821.670 3270.500 1821.990 3270.560 ;
        RECT 1822.590 3270.500 1822.910 3270.560 ;
        RECT 297.690 3254.040 298.010 3254.100 ;
        RECT 1821.670 3254.040 1821.990 3254.100 ;
        RECT 297.690 3253.900 1821.990 3254.040 ;
        RECT 297.690 3253.840 298.010 3253.900 ;
        RECT 1821.670 3253.840 1821.990 3253.900 ;
      LAYER via ;
        RECT 1822.160 3491.160 1822.420 3491.420 ;
        RECT 1825.380 3491.160 1825.640 3491.420 ;
        RECT 1822.160 3347.000 1822.420 3347.260 ;
        RECT 1822.160 3346.320 1822.420 3346.580 ;
        RECT 1821.700 3270.500 1821.960 3270.760 ;
        RECT 1822.620 3270.500 1822.880 3270.760 ;
        RECT 297.720 3253.840 297.980 3254.100 ;
        RECT 1821.700 3253.840 1821.960 3254.100 ;
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
        RECT 1824.980 3517.370 1825.120 3517.600 ;
        RECT 1824.980 3517.230 1825.580 3517.370 ;
        RECT 1825.440 3491.450 1825.580 3517.230 ;
        RECT 1822.160 3491.130 1822.420 3491.450 ;
        RECT 1825.380 3491.130 1825.640 3491.450 ;
        RECT 1822.220 3443.250 1822.360 3491.130 ;
        RECT 1821.760 3443.110 1822.360 3443.250 ;
        RECT 1821.760 3442.570 1821.900 3443.110 ;
        RECT 1821.760 3442.430 1822.360 3442.570 ;
        RECT 1822.220 3347.290 1822.360 3442.430 ;
        RECT 1822.160 3346.970 1822.420 3347.290 ;
        RECT 1822.160 3346.290 1822.420 3346.610 ;
        RECT 1822.220 3298.410 1822.360 3346.290 ;
        RECT 1822.220 3298.270 1822.820 3298.410 ;
        RECT 1822.680 3270.790 1822.820 3298.270 ;
        RECT 1821.700 3270.470 1821.960 3270.790 ;
        RECT 1822.620 3270.470 1822.880 3270.790 ;
        RECT 1821.760 3254.130 1821.900 3270.470 ;
        RECT 297.720 3253.810 297.980 3254.130 ;
        RECT 1821.700 3253.810 1821.960 3254.130 ;
        RECT 297.780 2073.845 297.920 3253.810 ;
        RECT 297.710 2073.475 297.990 2073.845 ;
      LAYER via2 ;
        RECT 297.710 2073.520 297.990 2073.800 ;
      LAYER met3 ;
        RECT 297.685 2073.810 298.015 2073.825 ;
        RECT 300.000 2073.810 304.000 2073.880 ;
        RECT 297.685 2073.510 304.000 2073.810 ;
        RECT 297.685 2073.495 298.015 2073.510 ;
        RECT 300.000 2073.280 304.000 2073.510 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1497.830 3429.480 1498.150 3429.540 ;
        RECT 1500.590 3429.480 1500.910 3429.540 ;
        RECT 1497.830 3429.340 1500.910 3429.480 ;
        RECT 1497.830 3429.280 1498.150 3429.340 ;
        RECT 1500.590 3429.280 1500.910 3429.340 ;
        RECT 1497.830 3422.340 1498.150 3422.400 ;
        RECT 1498.290 3422.340 1498.610 3422.400 ;
        RECT 1497.830 3422.200 1498.610 3422.340 ;
        RECT 1497.830 3422.140 1498.150 3422.200 ;
        RECT 1498.290 3422.140 1498.610 3422.200 ;
        RECT 1498.290 3395.140 1498.610 3395.200 ;
        RECT 1497.920 3395.000 1498.610 3395.140 ;
        RECT 1497.920 3394.860 1498.060 3395.000 ;
        RECT 1498.290 3394.940 1498.610 3395.000 ;
        RECT 1497.830 3394.600 1498.150 3394.860 ;
        RECT 1497.830 3332.920 1498.150 3332.980 ;
        RECT 1498.750 3332.920 1499.070 3332.980 ;
        RECT 1497.830 3332.780 1499.070 3332.920 ;
        RECT 1497.830 3332.720 1498.150 3332.780 ;
        RECT 1498.750 3332.720 1499.070 3332.780 ;
        RECT 1498.750 3298.580 1499.070 3298.640 ;
        RECT 1497.920 3298.440 1499.070 3298.580 ;
        RECT 1497.920 3298.300 1498.060 3298.440 ;
        RECT 1498.750 3298.380 1499.070 3298.440 ;
        RECT 1497.830 3298.040 1498.150 3298.300 ;
        RECT 1497.830 3249.960 1498.150 3250.020 ;
        RECT 1498.750 3249.960 1499.070 3250.020 ;
        RECT 1497.830 3249.820 1499.070 3249.960 ;
        RECT 1497.830 3249.760 1498.150 3249.820 ;
        RECT 1498.750 3249.760 1499.070 3249.820 ;
        RECT 1497.370 3211.880 1497.690 3211.940 ;
        RECT 1498.750 3211.880 1499.070 3211.940 ;
        RECT 1497.370 3211.740 1499.070 3211.880 ;
        RECT 1497.370 3211.680 1497.690 3211.740 ;
        RECT 1498.750 3211.680 1499.070 3211.740 ;
        RECT 1497.370 3188.420 1497.690 3188.480 ;
        RECT 1497.370 3188.280 1498.520 3188.420 ;
        RECT 1497.370 3188.220 1497.690 3188.280 ;
        RECT 1498.380 3188.140 1498.520 3188.280 ;
        RECT 1498.290 3187.880 1498.610 3188.140 ;
        RECT 1499.210 3139.800 1499.530 3139.860 ;
        RECT 1500.130 3139.800 1500.450 3139.860 ;
        RECT 1499.210 3139.660 1500.450 3139.800 ;
        RECT 1499.210 3139.600 1499.530 3139.660 ;
        RECT 1500.130 3139.600 1500.450 3139.660 ;
        RECT 1499.210 3105.460 1499.530 3105.520 ;
        RECT 1498.840 3105.320 1499.530 3105.460 ;
        RECT 1498.840 3104.840 1498.980 3105.320 ;
        RECT 1499.210 3105.260 1499.530 3105.320 ;
        RECT 1498.750 3104.580 1499.070 3104.840 ;
        RECT 1497.830 3056.840 1498.150 3056.900 ;
        RECT 1498.750 3056.840 1499.070 3056.900 ;
        RECT 1497.830 3056.700 1499.070 3056.840 ;
        RECT 1497.830 3056.640 1498.150 3056.700 ;
        RECT 1498.750 3056.640 1499.070 3056.700 ;
        RECT 1497.830 3042.900 1498.150 3042.960 ;
        RECT 1498.290 3042.900 1498.610 3042.960 ;
        RECT 1497.830 3042.760 1498.610 3042.900 ;
        RECT 1497.830 3042.700 1498.150 3042.760 ;
        RECT 1498.290 3042.700 1498.610 3042.760 ;
        RECT 1497.830 3008.560 1498.150 3008.620 ;
        RECT 1499.210 3008.560 1499.530 3008.620 ;
        RECT 1497.830 3008.420 1499.530 3008.560 ;
        RECT 1497.830 3008.360 1498.150 3008.420 ;
        RECT 1499.210 3008.360 1499.530 3008.420 ;
        RECT 1498.290 2994.620 1498.610 2994.680 ;
        RECT 1499.210 2994.620 1499.530 2994.680 ;
        RECT 1498.290 2994.480 1499.530 2994.620 ;
        RECT 1498.290 2994.420 1498.610 2994.480 ;
        RECT 1499.210 2994.420 1499.530 2994.480 ;
        RECT 1498.290 2946.680 1498.610 2946.740 ;
        RECT 1499.670 2946.680 1499.990 2946.740 ;
        RECT 1498.290 2946.540 1499.990 2946.680 ;
        RECT 1498.290 2946.480 1498.610 2946.540 ;
        RECT 1499.670 2946.480 1499.990 2946.540 ;
        RECT 1499.670 2912.340 1499.990 2912.400 ;
        RECT 1499.300 2912.200 1499.990 2912.340 ;
        RECT 1499.300 2911.720 1499.440 2912.200 ;
        RECT 1499.670 2912.140 1499.990 2912.200 ;
        RECT 1499.210 2911.460 1499.530 2911.720 ;
        RECT 284.350 2696.100 284.670 2696.160 ;
        RECT 1498.750 2696.100 1499.070 2696.160 ;
        RECT 284.350 2695.960 1499.070 2696.100 ;
        RECT 284.350 2695.900 284.670 2695.960 ;
        RECT 1498.750 2695.900 1499.070 2695.960 ;
      LAYER via ;
        RECT 1497.860 3429.280 1498.120 3429.540 ;
        RECT 1500.620 3429.280 1500.880 3429.540 ;
        RECT 1497.860 3422.140 1498.120 3422.400 ;
        RECT 1498.320 3422.140 1498.580 3422.400 ;
        RECT 1498.320 3394.940 1498.580 3395.200 ;
        RECT 1497.860 3394.600 1498.120 3394.860 ;
        RECT 1497.860 3332.720 1498.120 3332.980 ;
        RECT 1498.780 3332.720 1499.040 3332.980 ;
        RECT 1498.780 3298.380 1499.040 3298.640 ;
        RECT 1497.860 3298.040 1498.120 3298.300 ;
        RECT 1497.860 3249.760 1498.120 3250.020 ;
        RECT 1498.780 3249.760 1499.040 3250.020 ;
        RECT 1497.400 3211.680 1497.660 3211.940 ;
        RECT 1498.780 3211.680 1499.040 3211.940 ;
        RECT 1497.400 3188.220 1497.660 3188.480 ;
        RECT 1498.320 3187.880 1498.580 3188.140 ;
        RECT 1499.240 3139.600 1499.500 3139.860 ;
        RECT 1500.160 3139.600 1500.420 3139.860 ;
        RECT 1499.240 3105.260 1499.500 3105.520 ;
        RECT 1498.780 3104.580 1499.040 3104.840 ;
        RECT 1497.860 3056.640 1498.120 3056.900 ;
        RECT 1498.780 3056.640 1499.040 3056.900 ;
        RECT 1497.860 3042.700 1498.120 3042.960 ;
        RECT 1498.320 3042.700 1498.580 3042.960 ;
        RECT 1497.860 3008.360 1498.120 3008.620 ;
        RECT 1499.240 3008.360 1499.500 3008.620 ;
        RECT 1498.320 2994.420 1498.580 2994.680 ;
        RECT 1499.240 2994.420 1499.500 2994.680 ;
        RECT 1498.320 2946.480 1498.580 2946.740 ;
        RECT 1499.700 2946.480 1499.960 2946.740 ;
        RECT 1499.700 2912.140 1499.960 2912.400 ;
        RECT 1499.240 2911.460 1499.500 2911.720 ;
        RECT 284.380 2695.900 284.640 2696.160 ;
        RECT 1498.780 2695.900 1499.040 2696.160 ;
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
        RECT 1500.680 3429.570 1500.820 3517.600 ;
        RECT 1497.860 3429.250 1498.120 3429.570 ;
        RECT 1500.620 3429.250 1500.880 3429.570 ;
        RECT 1497.920 3422.430 1498.060 3429.250 ;
        RECT 1497.860 3422.110 1498.120 3422.430 ;
        RECT 1498.320 3422.110 1498.580 3422.430 ;
        RECT 1498.380 3395.230 1498.520 3422.110 ;
        RECT 1498.320 3394.910 1498.580 3395.230 ;
        RECT 1497.860 3394.570 1498.120 3394.890 ;
        RECT 1497.920 3333.010 1498.060 3394.570 ;
        RECT 1497.860 3332.690 1498.120 3333.010 ;
        RECT 1498.780 3332.690 1499.040 3333.010 ;
        RECT 1498.840 3298.670 1498.980 3332.690 ;
        RECT 1498.780 3298.350 1499.040 3298.670 ;
        RECT 1497.860 3298.010 1498.120 3298.330 ;
        RECT 1497.920 3250.050 1498.060 3298.010 ;
        RECT 1497.860 3249.730 1498.120 3250.050 ;
        RECT 1498.780 3249.730 1499.040 3250.050 ;
        RECT 1498.840 3211.970 1498.980 3249.730 ;
        RECT 1497.400 3211.650 1497.660 3211.970 ;
        RECT 1498.780 3211.650 1499.040 3211.970 ;
        RECT 1497.460 3188.510 1497.600 3211.650 ;
        RECT 1497.400 3188.190 1497.660 3188.510 ;
        RECT 1498.320 3187.850 1498.580 3188.170 ;
        RECT 1498.380 3187.685 1498.520 3187.850 ;
        RECT 1498.310 3187.315 1498.590 3187.685 ;
        RECT 1500.150 3187.315 1500.430 3187.685 ;
        RECT 1500.220 3139.890 1500.360 3187.315 ;
        RECT 1499.240 3139.570 1499.500 3139.890 ;
        RECT 1500.160 3139.570 1500.420 3139.890 ;
        RECT 1499.300 3105.550 1499.440 3139.570 ;
        RECT 1499.240 3105.230 1499.500 3105.550 ;
        RECT 1498.780 3104.550 1499.040 3104.870 ;
        RECT 1498.840 3056.930 1498.980 3104.550 ;
        RECT 1497.860 3056.610 1498.120 3056.930 ;
        RECT 1498.780 3056.610 1499.040 3056.930 ;
        RECT 1497.920 3056.330 1498.060 3056.610 ;
        RECT 1497.920 3056.190 1498.520 3056.330 ;
        RECT 1498.380 3042.990 1498.520 3056.190 ;
        RECT 1497.860 3042.670 1498.120 3042.990 ;
        RECT 1498.320 3042.670 1498.580 3042.990 ;
        RECT 1497.920 3008.650 1498.060 3042.670 ;
        RECT 1497.860 3008.330 1498.120 3008.650 ;
        RECT 1499.240 3008.330 1499.500 3008.650 ;
        RECT 1499.300 2994.710 1499.440 3008.330 ;
        RECT 1498.320 2994.390 1498.580 2994.710 ;
        RECT 1499.240 2994.390 1499.500 2994.710 ;
        RECT 1498.380 2946.770 1498.520 2994.390 ;
        RECT 1498.320 2946.450 1498.580 2946.770 ;
        RECT 1499.700 2946.450 1499.960 2946.770 ;
        RECT 1499.760 2912.430 1499.900 2946.450 ;
        RECT 1499.700 2912.110 1499.960 2912.430 ;
        RECT 1499.240 2911.430 1499.500 2911.750 ;
        RECT 1499.300 2863.210 1499.440 2911.430 ;
        RECT 1498.380 2863.070 1499.440 2863.210 ;
        RECT 1498.380 2815.610 1498.520 2863.070 ;
        RECT 1497.920 2815.470 1498.520 2815.610 ;
        RECT 1497.920 2814.930 1498.060 2815.470 ;
        RECT 1497.920 2814.790 1498.520 2814.930 ;
        RECT 1498.380 2767.330 1498.520 2814.790 ;
        RECT 1498.380 2767.190 1498.980 2767.330 ;
        RECT 1498.840 2696.190 1498.980 2767.190 ;
        RECT 284.380 2695.870 284.640 2696.190 ;
        RECT 1498.780 2695.870 1499.040 2696.190 ;
        RECT 284.440 2105.125 284.580 2695.870 ;
        RECT 284.370 2104.755 284.650 2105.125 ;
      LAYER via2 ;
        RECT 1498.310 3187.360 1498.590 3187.640 ;
        RECT 1500.150 3187.360 1500.430 3187.640 ;
        RECT 284.370 2104.800 284.650 2105.080 ;
      LAYER met3 ;
        RECT 1498.285 3187.650 1498.615 3187.665 ;
        RECT 1500.125 3187.650 1500.455 3187.665 ;
        RECT 1498.285 3187.350 1500.455 3187.650 ;
        RECT 1498.285 3187.335 1498.615 3187.350 ;
        RECT 1500.125 3187.335 1500.455 3187.350 ;
        RECT 284.345 2105.090 284.675 2105.105 ;
        RECT 300.000 2105.090 304.000 2105.160 ;
        RECT 284.345 2104.790 304.000 2105.090 ;
        RECT 284.345 2104.775 284.675 2104.790 ;
        RECT 300.000 2104.560 304.000 2104.790 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 295.850 324.260 296.170 324.320 ;
        RECT 2898.990 324.260 2899.310 324.320 ;
        RECT 295.850 324.120 2899.310 324.260 ;
        RECT 295.850 324.060 296.170 324.120 ;
        RECT 2898.990 324.060 2899.310 324.120 ;
      LAYER via ;
        RECT 295.880 324.060 296.140 324.320 ;
        RECT 2899.020 324.060 2899.280 324.320 ;
      LAYER met2 ;
        RECT 295.870 1536.275 296.150 1536.645 ;
        RECT 295.940 324.350 296.080 1536.275 ;
        RECT 295.880 324.030 296.140 324.350 ;
        RECT 2899.020 324.030 2899.280 324.350 ;
        RECT 2899.080 322.845 2899.220 324.030 ;
        RECT 2899.010 322.475 2899.290 322.845 ;
      LAYER via2 ;
        RECT 295.870 1536.320 296.150 1536.600 ;
        RECT 2899.010 322.520 2899.290 322.800 ;
      LAYER met3 ;
        RECT 295.845 1536.610 296.175 1536.625 ;
        RECT 300.000 1536.610 304.000 1536.680 ;
        RECT 295.845 1536.310 304.000 1536.610 ;
        RECT 295.845 1536.295 296.175 1536.310 ;
        RECT 300.000 1536.080 304.000 1536.310 ;
        RECT 2898.985 322.810 2899.315 322.825 ;
        RECT 2917.600 322.810 2924.800 323.260 ;
        RECT 2898.985 322.510 2924.800 322.810 ;
        RECT 2898.985 322.495 2899.315 322.510 ;
        RECT 2917.600 322.060 2924.800 322.510 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 686.390 3501.220 686.710 3501.280 ;
        RECT 1175.830 3501.220 1176.150 3501.280 ;
        RECT 686.390 3501.080 1176.150 3501.220 ;
        RECT 686.390 3501.020 686.710 3501.080 ;
        RECT 1175.830 3501.020 1176.150 3501.080 ;
        RECT 283.890 2701.540 284.210 2701.600 ;
        RECT 686.390 2701.540 686.710 2701.600 ;
        RECT 283.890 2701.400 686.710 2701.540 ;
        RECT 283.890 2701.340 284.210 2701.400 ;
        RECT 686.390 2701.340 686.710 2701.400 ;
      LAYER via ;
        RECT 686.420 3501.020 686.680 3501.280 ;
        RECT 1175.860 3501.020 1176.120 3501.280 ;
        RECT 283.920 2701.340 284.180 2701.600 ;
        RECT 686.420 2701.340 686.680 2701.600 ;
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
        RECT 1175.920 3501.310 1176.060 3517.600 ;
        RECT 686.420 3500.990 686.680 3501.310 ;
        RECT 1175.860 3500.990 1176.120 3501.310 ;
        RECT 686.480 2701.630 686.620 3500.990 ;
        RECT 283.920 2701.310 284.180 2701.630 ;
        RECT 686.420 2701.310 686.680 2701.630 ;
        RECT 283.980 2136.405 284.120 2701.310 ;
        RECT 283.910 2136.035 284.190 2136.405 ;
      LAYER via2 ;
        RECT 283.910 2136.080 284.190 2136.360 ;
      LAYER met3 ;
        RECT 283.885 2136.370 284.215 2136.385 ;
        RECT 300.000 2136.370 304.000 2136.440 ;
        RECT 283.885 2136.070 304.000 2136.370 ;
        RECT 283.885 2136.055 284.215 2136.070 ;
        RECT 300.000 2135.840 304.000 2136.070 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 848.770 3477.420 849.090 3477.480 ;
        RECT 850.150 3477.420 850.470 3477.480 ;
        RECT 848.770 3477.280 850.470 3477.420 ;
        RECT 848.770 3477.220 849.090 3477.280 ;
        RECT 850.150 3477.220 850.470 3477.280 ;
        RECT 848.770 3429.480 849.090 3429.540 ;
        RECT 849.690 3429.480 850.010 3429.540 ;
        RECT 848.770 3429.340 850.010 3429.480 ;
        RECT 848.770 3429.280 849.090 3429.340 ;
        RECT 849.690 3429.280 850.010 3429.340 ;
        RECT 850.150 3298.580 850.470 3298.640 ;
        RECT 849.780 3298.440 850.470 3298.580 ;
        RECT 849.780 3298.300 849.920 3298.440 ;
        RECT 850.150 3298.380 850.470 3298.440 ;
        RECT 849.690 3298.040 850.010 3298.300 ;
        RECT 848.770 3277.500 849.090 3277.560 ;
        RECT 849.690 3277.500 850.010 3277.560 ;
        RECT 848.770 3277.360 850.010 3277.500 ;
        RECT 848.770 3277.300 849.090 3277.360 ;
        RECT 849.690 3277.300 850.010 3277.360 ;
        RECT 848.310 3181.280 848.630 3181.340 ;
        RECT 849.690 3181.280 850.010 3181.340 ;
        RECT 848.310 3181.140 850.010 3181.280 ;
        RECT 848.310 3181.080 848.630 3181.140 ;
        RECT 849.690 3181.080 850.010 3181.140 ;
        RECT 848.310 3139.800 848.630 3139.860 ;
        RECT 850.150 3139.800 850.470 3139.860 ;
        RECT 848.310 3139.660 850.470 3139.800 ;
        RECT 848.310 3139.600 848.630 3139.660 ;
        RECT 850.150 3139.600 850.470 3139.660 ;
        RECT 849.230 3091.520 849.550 3091.580 ;
        RECT 850.150 3091.520 850.470 3091.580 ;
        RECT 849.230 3091.380 850.470 3091.520 ;
        RECT 849.230 3091.320 849.550 3091.380 ;
        RECT 850.150 3091.320 850.470 3091.380 ;
        RECT 849.690 3057.180 850.010 3057.240 ;
        RECT 849.690 3057.040 850.380 3057.180 ;
        RECT 849.690 3056.980 850.010 3057.040 ;
        RECT 850.240 3056.220 850.380 3057.040 ;
        RECT 850.150 3055.960 850.470 3056.220 ;
        RECT 849.230 2994.960 849.550 2995.020 ;
        RECT 850.150 2994.960 850.470 2995.020 ;
        RECT 849.230 2994.820 850.470 2994.960 ;
        RECT 849.230 2994.760 849.550 2994.820 ;
        RECT 850.150 2994.760 850.470 2994.820 ;
        RECT 849.690 2960.620 850.010 2960.680 ;
        RECT 849.690 2960.480 850.380 2960.620 ;
        RECT 849.690 2960.420 850.010 2960.480 ;
        RECT 850.240 2959.660 850.380 2960.480 ;
        RECT 850.150 2959.400 850.470 2959.660 ;
        RECT 850.610 2891.260 850.930 2891.320 ;
        RECT 851.530 2891.260 851.850 2891.320 ;
        RECT 850.610 2891.120 851.850 2891.260 ;
        RECT 850.610 2891.060 850.930 2891.120 ;
        RECT 851.530 2891.060 851.850 2891.120 ;
        RECT 850.610 2863.520 850.930 2863.780 ;
        RECT 850.700 2863.100 850.840 2863.520 ;
        RECT 850.610 2862.840 850.930 2863.100 ;
        RECT 850.610 2815.780 850.930 2815.840 ;
        RECT 850.240 2815.640 850.930 2815.780 ;
        RECT 850.240 2815.160 850.380 2815.640 ;
        RECT 850.610 2815.580 850.930 2815.640 ;
        RECT 850.150 2814.900 850.470 2815.160 ;
        RECT 849.230 2767.160 849.550 2767.220 ;
        RECT 850.150 2767.160 850.470 2767.220 ;
        RECT 849.230 2767.020 850.470 2767.160 ;
        RECT 849.230 2766.960 849.550 2767.020 ;
        RECT 850.150 2766.960 850.470 2767.020 ;
        RECT 283.430 2701.200 283.750 2701.260 ;
        RECT 850.150 2701.200 850.470 2701.260 ;
        RECT 283.430 2701.060 850.470 2701.200 ;
        RECT 283.430 2701.000 283.750 2701.060 ;
        RECT 850.150 2701.000 850.470 2701.060 ;
      LAYER via ;
        RECT 848.800 3477.220 849.060 3477.480 ;
        RECT 850.180 3477.220 850.440 3477.480 ;
        RECT 848.800 3429.280 849.060 3429.540 ;
        RECT 849.720 3429.280 849.980 3429.540 ;
        RECT 850.180 3298.380 850.440 3298.640 ;
        RECT 849.720 3298.040 849.980 3298.300 ;
        RECT 848.800 3277.300 849.060 3277.560 ;
        RECT 849.720 3277.300 849.980 3277.560 ;
        RECT 848.340 3181.080 848.600 3181.340 ;
        RECT 849.720 3181.080 849.980 3181.340 ;
        RECT 848.340 3139.600 848.600 3139.860 ;
        RECT 850.180 3139.600 850.440 3139.860 ;
        RECT 849.260 3091.320 849.520 3091.580 ;
        RECT 850.180 3091.320 850.440 3091.580 ;
        RECT 849.720 3056.980 849.980 3057.240 ;
        RECT 850.180 3055.960 850.440 3056.220 ;
        RECT 849.260 2994.760 849.520 2995.020 ;
        RECT 850.180 2994.760 850.440 2995.020 ;
        RECT 849.720 2960.420 849.980 2960.680 ;
        RECT 850.180 2959.400 850.440 2959.660 ;
        RECT 850.640 2891.060 850.900 2891.320 ;
        RECT 851.560 2891.060 851.820 2891.320 ;
        RECT 850.640 2863.520 850.900 2863.780 ;
        RECT 850.640 2862.840 850.900 2863.100 ;
        RECT 850.640 2815.580 850.900 2815.840 ;
        RECT 850.180 2814.900 850.440 2815.160 ;
        RECT 849.260 2766.960 849.520 2767.220 ;
        RECT 850.180 2766.960 850.440 2767.220 ;
        RECT 283.460 2701.000 283.720 2701.260 ;
        RECT 850.180 2701.000 850.440 2701.260 ;
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
        RECT 851.620 3517.370 851.760 3517.600 ;
        RECT 850.700 3517.230 851.760 3517.370 ;
        RECT 850.700 3491.530 850.840 3517.230 ;
        RECT 850.240 3491.390 850.840 3491.530 ;
        RECT 850.240 3477.510 850.380 3491.390 ;
        RECT 848.800 3477.190 849.060 3477.510 ;
        RECT 850.180 3477.190 850.440 3477.510 ;
        RECT 848.860 3429.570 849.000 3477.190 ;
        RECT 848.800 3429.250 849.060 3429.570 ;
        RECT 849.720 3429.250 849.980 3429.570 ;
        RECT 849.780 3394.970 849.920 3429.250 ;
        RECT 849.320 3394.830 849.920 3394.970 ;
        RECT 849.320 3333.205 849.460 3394.830 ;
        RECT 849.250 3332.835 849.530 3333.205 ;
        RECT 850.170 3332.835 850.450 3333.205 ;
        RECT 850.240 3298.670 850.380 3332.835 ;
        RECT 850.180 3298.350 850.440 3298.670 ;
        RECT 849.720 3298.010 849.980 3298.330 ;
        RECT 849.780 3277.590 849.920 3298.010 ;
        RECT 848.800 3277.270 849.060 3277.590 ;
        RECT 849.720 3277.270 849.980 3277.590 ;
        RECT 848.860 3229.845 849.000 3277.270 ;
        RECT 848.790 3229.475 849.070 3229.845 ;
        RECT 850.170 3229.475 850.450 3229.845 ;
        RECT 850.240 3203.210 850.380 3229.475 ;
        RECT 849.780 3203.070 850.380 3203.210 ;
        RECT 849.780 3181.370 849.920 3203.070 ;
        RECT 848.340 3181.050 848.600 3181.370 ;
        RECT 849.720 3181.050 849.980 3181.370 ;
        RECT 848.400 3139.890 848.540 3181.050 ;
        RECT 848.340 3139.570 848.600 3139.890 ;
        RECT 850.180 3139.570 850.440 3139.890 ;
        RECT 850.240 3091.610 850.380 3139.570 ;
        RECT 849.260 3091.290 849.520 3091.610 ;
        RECT 850.180 3091.290 850.440 3091.610 ;
        RECT 849.320 3091.010 849.460 3091.290 ;
        RECT 849.320 3090.870 849.920 3091.010 ;
        RECT 849.780 3057.270 849.920 3090.870 ;
        RECT 849.720 3056.950 849.980 3057.270 ;
        RECT 850.180 3055.930 850.440 3056.250 ;
        RECT 850.240 2995.050 850.380 3055.930 ;
        RECT 849.260 2994.730 849.520 2995.050 ;
        RECT 850.180 2994.730 850.440 2995.050 ;
        RECT 849.320 2994.450 849.460 2994.730 ;
        RECT 849.320 2994.310 849.920 2994.450 ;
        RECT 849.780 2960.710 849.920 2994.310 ;
        RECT 849.720 2960.390 849.980 2960.710 ;
        RECT 850.180 2959.370 850.440 2959.690 ;
        RECT 850.240 2939.485 850.380 2959.370 ;
        RECT 850.170 2939.115 850.450 2939.485 ;
        RECT 851.550 2939.115 851.830 2939.485 ;
        RECT 851.620 2891.350 851.760 2939.115 ;
        RECT 850.640 2891.030 850.900 2891.350 ;
        RECT 851.560 2891.030 851.820 2891.350 ;
        RECT 850.700 2863.810 850.840 2891.030 ;
        RECT 850.640 2863.490 850.900 2863.810 ;
        RECT 850.640 2862.810 850.900 2863.130 ;
        RECT 850.700 2815.870 850.840 2862.810 ;
        RECT 850.640 2815.550 850.900 2815.870 ;
        RECT 850.180 2814.870 850.440 2815.190 ;
        RECT 850.240 2767.250 850.380 2814.870 ;
        RECT 849.260 2766.930 849.520 2767.250 ;
        RECT 850.180 2766.930 850.440 2767.250 ;
        RECT 849.320 2766.650 849.460 2766.930 ;
        RECT 849.320 2766.510 849.920 2766.650 ;
        RECT 849.780 2719.050 849.920 2766.510 ;
        RECT 849.780 2718.910 850.380 2719.050 ;
        RECT 850.240 2701.290 850.380 2718.910 ;
        RECT 283.460 2700.970 283.720 2701.290 ;
        RECT 850.180 2700.970 850.440 2701.290 ;
        RECT 283.520 2168.365 283.660 2700.970 ;
        RECT 283.450 2167.995 283.730 2168.365 ;
      LAYER via2 ;
        RECT 849.250 3332.880 849.530 3333.160 ;
        RECT 850.170 3332.880 850.450 3333.160 ;
        RECT 848.790 3229.520 849.070 3229.800 ;
        RECT 850.170 3229.520 850.450 3229.800 ;
        RECT 850.170 2939.160 850.450 2939.440 ;
        RECT 851.550 2939.160 851.830 2939.440 ;
        RECT 283.450 2168.040 283.730 2168.320 ;
      LAYER met3 ;
        RECT 849.225 3333.170 849.555 3333.185 ;
        RECT 850.145 3333.170 850.475 3333.185 ;
        RECT 849.225 3332.870 850.475 3333.170 ;
        RECT 849.225 3332.855 849.555 3332.870 ;
        RECT 850.145 3332.855 850.475 3332.870 ;
        RECT 848.765 3229.810 849.095 3229.825 ;
        RECT 850.145 3229.810 850.475 3229.825 ;
        RECT 848.765 3229.510 850.475 3229.810 ;
        RECT 848.765 3229.495 849.095 3229.510 ;
        RECT 850.145 3229.495 850.475 3229.510 ;
        RECT 850.145 2939.450 850.475 2939.465 ;
        RECT 851.525 2939.450 851.855 2939.465 ;
        RECT 850.145 2939.150 851.855 2939.450 ;
        RECT 850.145 2939.135 850.475 2939.150 ;
        RECT 851.525 2939.135 851.855 2939.150 ;
        RECT 283.425 2168.330 283.755 2168.345 ;
        RECT 300.000 2168.330 304.000 2168.400 ;
        RECT 283.425 2168.030 304.000 2168.330 ;
        RECT 283.425 2168.015 283.755 2168.030 ;
        RECT 300.000 2167.800 304.000 2168.030 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 524.930 3491.360 525.250 3491.420 ;
        RECT 527.690 3491.360 528.010 3491.420 ;
        RECT 524.930 3491.220 528.010 3491.360 ;
        RECT 524.930 3491.160 525.250 3491.220 ;
        RECT 527.690 3491.160 528.010 3491.220 ;
        RECT 524.470 3367.600 524.790 3367.660 ;
        RECT 525.390 3367.600 525.710 3367.660 ;
        RECT 524.470 3367.460 525.710 3367.600 ;
        RECT 524.470 3367.400 524.790 3367.460 ;
        RECT 525.390 3367.400 525.710 3367.460 ;
        RECT 524.470 3270.700 524.790 3270.760 ;
        RECT 525.390 3270.700 525.710 3270.760 ;
        RECT 524.470 3270.560 525.710 3270.700 ;
        RECT 524.470 3270.500 524.790 3270.560 ;
        RECT 525.390 3270.500 525.710 3270.560 ;
        RECT 287.110 3254.380 287.430 3254.440 ;
        RECT 524.470 3254.380 524.790 3254.440 ;
        RECT 287.110 3254.240 524.790 3254.380 ;
        RECT 287.110 3254.180 287.430 3254.240 ;
        RECT 524.470 3254.180 524.790 3254.240 ;
      LAYER via ;
        RECT 524.960 3491.160 525.220 3491.420 ;
        RECT 527.720 3491.160 527.980 3491.420 ;
        RECT 524.500 3367.400 524.760 3367.660 ;
        RECT 525.420 3367.400 525.680 3367.660 ;
        RECT 524.500 3270.500 524.760 3270.760 ;
        RECT 525.420 3270.500 525.680 3270.760 ;
        RECT 287.140 3254.180 287.400 3254.440 ;
        RECT 524.500 3254.180 524.760 3254.440 ;
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
        RECT 527.320 3517.370 527.460 3517.600 ;
        RECT 527.320 3517.230 527.920 3517.370 ;
        RECT 527.780 3491.450 527.920 3517.230 ;
        RECT 524.960 3491.130 525.220 3491.450 ;
        RECT 527.720 3491.130 527.980 3491.450 ;
        RECT 525.020 3443.250 525.160 3491.130 ;
        RECT 524.560 3443.110 525.160 3443.250 ;
        RECT 524.560 3415.370 524.700 3443.110 ;
        RECT 524.560 3415.230 525.620 3415.370 ;
        RECT 525.480 3367.690 525.620 3415.230 ;
        RECT 524.500 3367.370 524.760 3367.690 ;
        RECT 525.420 3367.370 525.680 3367.690 ;
        RECT 524.560 3318.810 524.700 3367.370 ;
        RECT 524.560 3318.670 525.620 3318.810 ;
        RECT 525.480 3270.790 525.620 3318.670 ;
        RECT 524.500 3270.470 524.760 3270.790 ;
        RECT 525.420 3270.470 525.680 3270.790 ;
        RECT 524.560 3254.470 524.700 3270.470 ;
        RECT 287.140 3254.150 287.400 3254.470 ;
        RECT 524.500 3254.150 524.760 3254.470 ;
        RECT 287.200 2199.645 287.340 3254.150 ;
        RECT 287.130 2199.275 287.410 2199.645 ;
      LAYER via2 ;
        RECT 287.130 2199.320 287.410 2199.600 ;
      LAYER met3 ;
        RECT 287.105 2199.610 287.435 2199.625 ;
        RECT 300.000 2199.610 304.000 2199.680 ;
        RECT 287.105 2199.310 304.000 2199.610 ;
        RECT 287.105 2199.295 287.435 2199.310 ;
        RECT 300.000 2199.080 304.000 2199.310 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 202.470 3499.860 202.790 3499.920 ;
        RECT 210.290 3499.860 210.610 3499.920 ;
        RECT 202.470 3499.720 210.610 3499.860 ;
        RECT 202.470 3499.660 202.790 3499.720 ;
        RECT 210.290 3499.660 210.610 3499.720 ;
        RECT 210.290 2235.400 210.610 2235.460 ;
        RECT 287.570 2235.400 287.890 2235.460 ;
        RECT 210.290 2235.260 287.890 2235.400 ;
        RECT 210.290 2235.200 210.610 2235.260 ;
        RECT 287.570 2235.200 287.890 2235.260 ;
      LAYER via ;
        RECT 202.500 3499.660 202.760 3499.920 ;
        RECT 210.320 3499.660 210.580 3499.920 ;
        RECT 210.320 2235.200 210.580 2235.460 ;
        RECT 287.600 2235.200 287.860 2235.460 ;
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
        RECT 202.560 3499.950 202.700 3517.600 ;
        RECT 202.500 3499.630 202.760 3499.950 ;
        RECT 210.320 3499.630 210.580 3499.950 ;
        RECT 210.380 2235.490 210.520 3499.630 ;
        RECT 210.320 2235.170 210.580 2235.490 ;
        RECT 287.600 2235.170 287.860 2235.490 ;
        RECT 287.660 2231.605 287.800 2235.170 ;
        RECT 287.590 2231.235 287.870 2231.605 ;
      LAYER via2 ;
        RECT 287.590 2231.280 287.870 2231.560 ;
      LAYER met3 ;
        RECT 287.565 2231.570 287.895 2231.585 ;
        RECT 300.000 2231.570 304.000 2231.640 ;
        RECT 287.565 2231.270 304.000 2231.570 ;
        RECT 287.565 2231.255 287.895 2231.270 ;
        RECT 300.000 2231.040 304.000 2231.270 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 13.870 3408.740 14.190 3408.800 ;
        RECT 25.370 3408.740 25.690 3408.800 ;
        RECT 13.870 3408.600 25.690 3408.740 ;
        RECT 13.870 3408.540 14.190 3408.600 ;
        RECT 25.370 3408.540 25.690 3408.600 ;
        RECT 25.370 2262.600 25.690 2262.660 ;
        RECT 282.970 2262.600 283.290 2262.660 ;
        RECT 25.370 2262.460 283.290 2262.600 ;
        RECT 25.370 2262.400 25.690 2262.460 ;
        RECT 282.970 2262.400 283.290 2262.460 ;
      LAYER via ;
        RECT 13.900 3408.540 14.160 3408.800 ;
        RECT 25.400 3408.540 25.660 3408.800 ;
        RECT 25.400 2262.400 25.660 2262.660 ;
        RECT 283.000 2262.400 283.260 2262.660 ;
      LAYER met2 ;
        RECT 13.890 3411.035 14.170 3411.405 ;
        RECT 13.960 3408.830 14.100 3411.035 ;
        RECT 13.900 3408.510 14.160 3408.830 ;
        RECT 25.400 3408.510 25.660 3408.830 ;
        RECT 25.460 2262.690 25.600 3408.510 ;
        RECT 25.400 2262.370 25.660 2262.690 ;
        RECT 282.990 2262.515 283.270 2262.885 ;
        RECT 283.000 2262.370 283.260 2262.515 ;
      LAYER via2 ;
        RECT 13.890 3411.080 14.170 3411.360 ;
        RECT 282.990 2262.560 283.270 2262.840 ;
      LAYER met3 ;
        RECT -4.800 3411.370 2.400 3411.820 ;
        RECT 13.865 3411.370 14.195 3411.385 ;
        RECT -4.800 3411.070 14.195 3411.370 ;
        RECT -4.800 3410.620 2.400 3411.070 ;
        RECT 13.865 3411.055 14.195 3411.070 ;
        RECT 282.965 2262.850 283.295 2262.865 ;
        RECT 300.000 2262.850 304.000 2262.920 ;
        RECT 282.965 2262.550 304.000 2262.850 ;
        RECT 282.965 2262.535 283.295 2262.550 ;
        RECT 300.000 2262.320 304.000 2262.550 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 19.390 3119.060 19.710 3119.120 ;
        RECT 25.830 3119.060 26.150 3119.120 ;
        RECT 19.390 3118.920 26.150 3119.060 ;
        RECT 19.390 3118.860 19.710 3118.920 ;
        RECT 25.830 3118.860 26.150 3118.920 ;
        RECT 25.830 2297.620 26.150 2297.680 ;
        RECT 282.970 2297.620 283.290 2297.680 ;
        RECT 25.830 2297.480 283.290 2297.620 ;
        RECT 25.830 2297.420 26.150 2297.480 ;
        RECT 282.970 2297.420 283.290 2297.480 ;
      LAYER via ;
        RECT 19.420 3118.860 19.680 3119.120 ;
        RECT 25.860 3118.860 26.120 3119.120 ;
        RECT 25.860 2297.420 26.120 2297.680 ;
        RECT 283.000 2297.420 283.260 2297.680 ;
      LAYER met2 ;
        RECT 19.410 3124.075 19.690 3124.445 ;
        RECT 19.480 3119.150 19.620 3124.075 ;
        RECT 19.420 3118.830 19.680 3119.150 ;
        RECT 25.860 3118.830 26.120 3119.150 ;
        RECT 25.920 2297.710 26.060 3118.830 ;
        RECT 25.860 2297.390 26.120 2297.710 ;
        RECT 283.000 2297.390 283.260 2297.710 ;
        RECT 283.060 2294.845 283.200 2297.390 ;
        RECT 282.990 2294.475 283.270 2294.845 ;
      LAYER via2 ;
        RECT 19.410 3124.120 19.690 3124.400 ;
        RECT 282.990 2294.520 283.270 2294.800 ;
      LAYER met3 ;
        RECT -4.800 3124.410 2.400 3124.860 ;
        RECT 19.385 3124.410 19.715 3124.425 ;
        RECT -4.800 3124.110 19.715 3124.410 ;
        RECT -4.800 3123.660 2.400 3124.110 ;
        RECT 19.385 3124.095 19.715 3124.110 ;
        RECT 282.965 2294.810 283.295 2294.825 ;
        RECT 300.000 2294.810 304.000 2294.880 ;
        RECT 282.965 2294.510 304.000 2294.810 ;
        RECT 282.965 2294.495 283.295 2294.510 ;
        RECT 300.000 2294.280 304.000 2294.510 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 19.850 2836.180 20.170 2836.240 ;
        RECT 26.290 2836.180 26.610 2836.240 ;
        RECT 19.850 2836.040 26.610 2836.180 ;
        RECT 19.850 2835.980 20.170 2836.040 ;
        RECT 26.290 2835.980 26.610 2836.040 ;
        RECT 26.290 2331.960 26.610 2332.020 ;
        RECT 282.510 2331.960 282.830 2332.020 ;
        RECT 26.290 2331.820 282.830 2331.960 ;
        RECT 26.290 2331.760 26.610 2331.820 ;
        RECT 282.510 2331.760 282.830 2331.820 ;
      LAYER via ;
        RECT 19.880 2835.980 20.140 2836.240 ;
        RECT 26.320 2835.980 26.580 2836.240 ;
        RECT 26.320 2331.760 26.580 2332.020 ;
        RECT 282.540 2331.760 282.800 2332.020 ;
      LAYER met2 ;
        RECT 19.870 2836.435 20.150 2836.805 ;
        RECT 19.940 2836.270 20.080 2836.435 ;
        RECT 19.880 2835.950 20.140 2836.270 ;
        RECT 26.320 2835.950 26.580 2836.270 ;
        RECT 26.380 2332.050 26.520 2835.950 ;
        RECT 26.320 2331.730 26.580 2332.050 ;
        RECT 282.540 2331.730 282.800 2332.050 ;
        RECT 282.600 2328.845 282.740 2331.730 ;
        RECT 282.530 2328.475 282.810 2328.845 ;
      LAYER via2 ;
        RECT 19.870 2836.480 20.150 2836.760 ;
        RECT 282.530 2328.520 282.810 2328.800 ;
      LAYER met3 ;
        RECT -4.800 2836.770 2.400 2837.220 ;
        RECT 19.845 2836.770 20.175 2836.785 ;
        RECT -4.800 2836.470 20.175 2836.770 ;
        RECT -4.800 2836.020 2.400 2836.470 ;
        RECT 19.845 2836.455 20.175 2836.470 ;
        RECT 282.505 2328.810 282.835 2328.825 ;
        RECT 282.505 2328.510 300.530 2328.810 ;
        RECT 282.505 2328.495 282.835 2328.510 ;
        RECT 300.230 2326.160 300.530 2328.510 ;
        RECT 300.000 2325.560 304.000 2326.160 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 13.870 2547.860 14.190 2547.920 ;
        RECT 27.210 2547.860 27.530 2547.920 ;
        RECT 13.870 2547.720 27.530 2547.860 ;
        RECT 13.870 2547.660 14.190 2547.720 ;
        RECT 27.210 2547.660 27.530 2547.720 ;
        RECT 27.210 2359.840 27.530 2359.900 ;
        RECT 282.970 2359.840 283.290 2359.900 ;
        RECT 27.210 2359.700 283.290 2359.840 ;
        RECT 27.210 2359.640 27.530 2359.700 ;
        RECT 282.970 2359.640 283.290 2359.700 ;
      LAYER via ;
        RECT 13.900 2547.660 14.160 2547.920 ;
        RECT 27.240 2547.660 27.500 2547.920 ;
        RECT 27.240 2359.640 27.500 2359.900 ;
        RECT 283.000 2359.640 283.260 2359.900 ;
      LAYER met2 ;
        RECT 13.890 2549.475 14.170 2549.845 ;
        RECT 13.960 2547.950 14.100 2549.475 ;
        RECT 13.900 2547.630 14.160 2547.950 ;
        RECT 27.240 2547.630 27.500 2547.950 ;
        RECT 27.300 2359.930 27.440 2547.630 ;
        RECT 27.240 2359.610 27.500 2359.930 ;
        RECT 283.000 2359.610 283.260 2359.930 ;
        RECT 283.060 2358.085 283.200 2359.610 ;
        RECT 282.990 2357.715 283.270 2358.085 ;
      LAYER via2 ;
        RECT 13.890 2549.520 14.170 2549.800 ;
        RECT 282.990 2357.760 283.270 2358.040 ;
      LAYER met3 ;
        RECT -4.800 2549.810 2.400 2550.260 ;
        RECT 13.865 2549.810 14.195 2549.825 ;
        RECT -4.800 2549.510 14.195 2549.810 ;
        RECT -4.800 2549.060 2.400 2549.510 ;
        RECT 13.865 2549.495 14.195 2549.510 ;
        RECT 282.965 2358.050 283.295 2358.065 ;
        RECT 300.000 2358.050 304.000 2358.120 ;
        RECT 282.965 2357.750 304.000 2358.050 ;
        RECT 282.965 2357.735 283.295 2357.750 ;
        RECT 300.000 2357.520 304.000 2357.750 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 16.630 2261.920 16.950 2261.980 ;
        RECT 282.510 2261.920 282.830 2261.980 ;
        RECT 16.630 2261.780 282.830 2261.920 ;
        RECT 16.630 2261.720 16.950 2261.780 ;
        RECT 282.510 2261.720 282.830 2261.780 ;
      LAYER via ;
        RECT 16.660 2261.720 16.920 2261.980 ;
        RECT 282.540 2261.720 282.800 2261.980 ;
      LAYER met2 ;
        RECT 282.990 2388.995 283.270 2389.365 ;
        RECT 283.060 2381.090 283.200 2388.995 ;
        RECT 282.600 2380.950 283.200 2381.090 ;
        RECT 282.600 2378.370 282.740 2380.950 ;
        RECT 282.600 2378.230 283.200 2378.370 ;
        RECT 283.060 2374.290 283.200 2378.230 ;
        RECT 282.600 2374.150 283.200 2374.290 ;
        RECT 282.600 2367.490 282.740 2374.150 ;
        RECT 282.600 2367.350 283.200 2367.490 ;
        RECT 283.060 2360.690 283.200 2367.350 ;
        RECT 282.600 2360.550 283.200 2360.690 ;
        RECT 282.600 2357.290 282.740 2360.550 ;
        RECT 282.600 2357.150 283.200 2357.290 ;
        RECT 283.060 2298.130 283.200 2357.150 ;
        RECT 282.600 2297.990 283.200 2298.130 ;
        RECT 282.600 2294.050 282.740 2297.990 ;
        RECT 282.600 2293.910 283.200 2294.050 ;
        RECT 283.060 2284.530 283.200 2293.910 ;
        RECT 282.600 2284.390 283.200 2284.530 ;
        RECT 282.600 2283.170 282.740 2284.390 ;
        RECT 282.600 2283.030 283.200 2283.170 ;
        RECT 283.060 2277.730 283.200 2283.030 ;
        RECT 282.600 2277.590 283.200 2277.730 ;
        RECT 282.600 2272.970 282.740 2277.590 ;
        RECT 282.600 2272.830 283.200 2272.970 ;
        RECT 283.060 2263.450 283.200 2272.830 ;
        RECT 282.600 2263.310 283.200 2263.450 ;
        RECT 16.650 2261.835 16.930 2262.205 ;
        RECT 282.600 2262.010 282.740 2263.310 ;
        RECT 16.660 2261.690 16.920 2261.835 ;
        RECT 282.540 2261.690 282.800 2262.010 ;
      LAYER via2 ;
        RECT 282.990 2389.040 283.270 2389.320 ;
        RECT 16.650 2261.880 16.930 2262.160 ;
      LAYER met3 ;
        RECT 282.965 2389.330 283.295 2389.345 ;
        RECT 300.000 2389.330 304.000 2389.400 ;
        RECT 282.965 2389.030 304.000 2389.330 ;
        RECT 282.965 2389.015 283.295 2389.030 ;
        RECT 300.000 2388.800 304.000 2389.030 ;
        RECT -4.800 2262.170 2.400 2262.620 ;
        RECT 16.625 2262.170 16.955 2262.185 ;
        RECT -4.800 2261.870 16.955 2262.170 ;
        RECT -4.800 2261.420 2.400 2261.870 ;
        RECT 16.625 2261.855 16.955 2261.870 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 18.930 2415.260 19.250 2415.320 ;
        RECT 282.970 2415.260 283.290 2415.320 ;
        RECT 18.930 2415.120 283.290 2415.260 ;
        RECT 18.930 2415.060 19.250 2415.120 ;
        RECT 282.970 2415.060 283.290 2415.120 ;
      LAYER via ;
        RECT 18.960 2415.060 19.220 2415.320 ;
        RECT 283.000 2415.060 283.260 2415.320 ;
      LAYER met2 ;
        RECT 282.990 2420.275 283.270 2420.645 ;
        RECT 283.060 2415.350 283.200 2420.275 ;
        RECT 18.960 2415.030 19.220 2415.350 ;
        RECT 283.000 2415.030 283.260 2415.350 ;
        RECT 19.020 1975.245 19.160 2415.030 ;
        RECT 18.950 1974.875 19.230 1975.245 ;
      LAYER via2 ;
        RECT 282.990 2420.320 283.270 2420.600 ;
        RECT 18.950 1974.920 19.230 1975.200 ;
      LAYER met3 ;
        RECT 282.965 2420.610 283.295 2420.625 ;
        RECT 300.000 2420.610 304.000 2420.680 ;
        RECT 282.965 2420.310 304.000 2420.610 ;
        RECT 282.965 2420.295 283.295 2420.310 ;
        RECT 300.000 2420.080 304.000 2420.310 ;
        RECT -4.800 1975.210 2.400 1975.660 ;
        RECT 18.925 1975.210 19.255 1975.225 ;
        RECT -4.800 1974.910 19.255 1975.210 ;
        RECT -4.800 1974.460 2.400 1974.910 ;
        RECT 18.925 1974.895 19.255 1974.910 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 295.390 558.860 295.710 558.920 ;
        RECT 2898.990 558.860 2899.310 558.920 ;
        RECT 295.390 558.720 2899.310 558.860 ;
        RECT 295.390 558.660 295.710 558.720 ;
        RECT 2898.990 558.660 2899.310 558.720 ;
      LAYER via ;
        RECT 295.420 558.660 295.680 558.920 ;
        RECT 2899.020 558.660 2899.280 558.920 ;
      LAYER met2 ;
        RECT 295.410 1567.555 295.690 1567.925 ;
        RECT 295.480 558.950 295.620 1567.555 ;
        RECT 295.420 558.630 295.680 558.950 ;
        RECT 2899.020 558.630 2899.280 558.950 ;
        RECT 2899.080 557.445 2899.220 558.630 ;
        RECT 2899.010 557.075 2899.290 557.445 ;
      LAYER via2 ;
        RECT 295.410 1567.600 295.690 1567.880 ;
        RECT 2899.010 557.120 2899.290 557.400 ;
      LAYER met3 ;
        RECT 295.385 1567.890 295.715 1567.905 ;
        RECT 300.000 1567.890 304.000 1567.960 ;
        RECT 295.385 1567.590 304.000 1567.890 ;
        RECT 295.385 1567.575 295.715 1567.590 ;
        RECT 300.000 1567.360 304.000 1567.590 ;
        RECT 2898.985 557.410 2899.315 557.425 ;
        RECT 2917.600 557.410 2924.800 557.860 ;
        RECT 2898.985 557.110 2924.800 557.410 ;
        RECT 2898.985 557.095 2899.315 557.110 ;
        RECT 2917.600 556.660 2924.800 557.110 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 16.630 1690.380 16.950 1690.440 ;
        RECT 284.810 1690.380 285.130 1690.440 ;
        RECT 16.630 1690.240 285.130 1690.380 ;
        RECT 16.630 1690.180 16.950 1690.240 ;
        RECT 284.810 1690.180 285.130 1690.240 ;
      LAYER via ;
        RECT 16.660 1690.180 16.920 1690.440 ;
        RECT 284.840 1690.180 285.100 1690.440 ;
      LAYER met2 ;
        RECT 284.830 2452.235 285.110 2452.605 ;
        RECT 284.900 1690.470 285.040 2452.235 ;
        RECT 16.660 1690.150 16.920 1690.470 ;
        RECT 284.840 1690.150 285.100 1690.470 ;
        RECT 16.720 1687.605 16.860 1690.150 ;
        RECT 16.650 1687.235 16.930 1687.605 ;
      LAYER via2 ;
        RECT 284.830 2452.280 285.110 2452.560 ;
        RECT 16.650 1687.280 16.930 1687.560 ;
      LAYER met3 ;
        RECT 284.805 2452.570 285.135 2452.585 ;
        RECT 300.000 2452.570 304.000 2452.640 ;
        RECT 284.805 2452.270 304.000 2452.570 ;
        RECT 284.805 2452.255 285.135 2452.270 ;
        RECT 300.000 2452.040 304.000 2452.270 ;
        RECT -4.800 1687.570 2.400 1688.020 ;
        RECT 16.625 1687.570 16.955 1687.585 ;
        RECT -4.800 1687.270 16.955 1687.570 ;
        RECT -4.800 1686.820 2.400 1687.270 ;
        RECT 16.625 1687.255 16.955 1687.270 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 284.810 2456.060 285.130 2456.120 ;
        RECT 286.190 2456.060 286.510 2456.120 ;
        RECT 284.810 2455.920 286.510 2456.060 ;
        RECT 284.810 2455.860 285.130 2455.920 ;
        RECT 286.190 2455.860 286.510 2455.920 ;
        RECT 14.790 1476.520 15.110 1476.580 ;
        RECT 286.190 1476.520 286.510 1476.580 ;
        RECT 14.790 1476.380 286.510 1476.520 ;
        RECT 14.790 1476.320 15.110 1476.380 ;
        RECT 286.190 1476.320 286.510 1476.380 ;
      LAYER via ;
        RECT 284.840 2455.860 285.100 2456.120 ;
        RECT 286.220 2455.860 286.480 2456.120 ;
        RECT 14.820 1476.320 15.080 1476.580 ;
        RECT 286.220 1476.320 286.480 1476.580 ;
      LAYER met2 ;
        RECT 284.830 2483.515 285.110 2483.885 ;
        RECT 284.900 2456.150 285.040 2483.515 ;
        RECT 284.840 2455.830 285.100 2456.150 ;
        RECT 286.220 2455.830 286.480 2456.150 ;
        RECT 286.280 1476.610 286.420 2455.830 ;
        RECT 14.820 1476.290 15.080 1476.610 ;
        RECT 286.220 1476.290 286.480 1476.610 ;
        RECT 14.880 1472.045 15.020 1476.290 ;
        RECT 14.810 1471.675 15.090 1472.045 ;
      LAYER via2 ;
        RECT 284.830 2483.560 285.110 2483.840 ;
        RECT 14.810 1471.720 15.090 1472.000 ;
      LAYER met3 ;
        RECT 284.805 2483.850 285.135 2483.865 ;
        RECT 300.000 2483.850 304.000 2483.920 ;
        RECT 284.805 2483.550 304.000 2483.850 ;
        RECT 284.805 2483.535 285.135 2483.550 ;
        RECT 300.000 2483.320 304.000 2483.550 ;
        RECT -4.800 1472.010 2.400 1472.460 ;
        RECT 14.785 1472.010 15.115 1472.025 ;
        RECT -4.800 1471.710 15.115 1472.010 ;
        RECT -4.800 1471.260 2.400 1471.710 ;
        RECT 14.785 1471.695 15.115 1471.710 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 18.010 2511.820 18.330 2511.880 ;
        RECT 286.190 2511.820 286.510 2511.880 ;
        RECT 18.010 2511.680 286.510 2511.820 ;
        RECT 18.010 2511.620 18.330 2511.680 ;
        RECT 286.190 2511.620 286.510 2511.680 ;
      LAYER via ;
        RECT 18.040 2511.620 18.300 2511.880 ;
        RECT 286.220 2511.620 286.480 2511.880 ;
      LAYER met2 ;
        RECT 286.210 2515.475 286.490 2515.845 ;
        RECT 286.280 2511.910 286.420 2515.475 ;
        RECT 18.040 2511.590 18.300 2511.910 ;
        RECT 286.220 2511.590 286.480 2511.910 ;
        RECT 18.100 1256.485 18.240 2511.590 ;
        RECT 18.030 1256.115 18.310 1256.485 ;
      LAYER via2 ;
        RECT 286.210 2515.520 286.490 2515.800 ;
        RECT 18.030 1256.160 18.310 1256.440 ;
      LAYER met3 ;
        RECT 286.185 2515.810 286.515 2515.825 ;
        RECT 300.000 2515.810 304.000 2515.880 ;
        RECT 286.185 2515.510 304.000 2515.810 ;
        RECT 286.185 2515.495 286.515 2515.510 ;
        RECT 300.000 2515.280 304.000 2515.510 ;
        RECT -4.800 1256.450 2.400 1256.900 ;
        RECT 18.005 1256.450 18.335 1256.465 ;
        RECT -4.800 1256.150 18.335 1256.450 ;
        RECT -4.800 1255.700 2.400 1256.150 ;
        RECT 18.005 1256.135 18.335 1256.150 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.550 2546.500 17.870 2546.560 ;
        RECT 286.190 2546.500 286.510 2546.560 ;
        RECT 17.550 2546.360 286.510 2546.500 ;
        RECT 17.550 2546.300 17.870 2546.360 ;
        RECT 286.190 2546.300 286.510 2546.360 ;
      LAYER via ;
        RECT 17.580 2546.300 17.840 2546.560 ;
        RECT 286.220 2546.300 286.480 2546.560 ;
      LAYER met2 ;
        RECT 286.210 2546.755 286.490 2547.125 ;
        RECT 286.280 2546.590 286.420 2546.755 ;
        RECT 17.580 2546.270 17.840 2546.590 ;
        RECT 286.220 2546.270 286.480 2546.590 ;
        RECT 17.640 1040.925 17.780 2546.270 ;
        RECT 17.570 1040.555 17.850 1040.925 ;
      LAYER via2 ;
        RECT 286.210 2546.800 286.490 2547.080 ;
        RECT 17.570 1040.600 17.850 1040.880 ;
      LAYER met3 ;
        RECT 286.185 2547.090 286.515 2547.105 ;
        RECT 300.000 2547.090 304.000 2547.160 ;
        RECT 286.185 2546.790 304.000 2547.090 ;
        RECT 286.185 2546.775 286.515 2546.790 ;
        RECT 300.000 2546.560 304.000 2546.790 ;
        RECT -4.800 1040.890 2.400 1041.340 ;
        RECT 17.545 1040.890 17.875 1040.905 ;
        RECT -4.800 1040.590 17.875 1040.890 ;
        RECT -4.800 1040.140 2.400 1040.590 ;
        RECT 17.545 1040.575 17.875 1040.590 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 2574.040 17.410 2574.100 ;
        RECT 286.190 2574.040 286.510 2574.100 ;
        RECT 17.090 2573.900 286.510 2574.040 ;
        RECT 17.090 2573.840 17.410 2573.900 ;
        RECT 286.190 2573.840 286.510 2573.900 ;
      LAYER via ;
        RECT 17.120 2573.840 17.380 2574.100 ;
        RECT 286.220 2573.840 286.480 2574.100 ;
      LAYER met2 ;
        RECT 286.210 2578.715 286.490 2579.085 ;
        RECT 286.280 2574.130 286.420 2578.715 ;
        RECT 17.120 2573.810 17.380 2574.130 ;
        RECT 286.220 2573.810 286.480 2574.130 ;
        RECT 17.180 825.365 17.320 2573.810 ;
        RECT 17.110 824.995 17.390 825.365 ;
      LAYER via2 ;
        RECT 286.210 2578.760 286.490 2579.040 ;
        RECT 17.110 825.040 17.390 825.320 ;
      LAYER met3 ;
        RECT 286.185 2579.050 286.515 2579.065 ;
        RECT 300.000 2579.050 304.000 2579.120 ;
        RECT 286.185 2578.750 304.000 2579.050 ;
        RECT 286.185 2578.735 286.515 2578.750 ;
        RECT 300.000 2578.520 304.000 2578.750 ;
        RECT -4.800 825.330 2.400 825.780 ;
        RECT 17.085 825.330 17.415 825.345 ;
        RECT -4.800 825.030 17.415 825.330 ;
        RECT -4.800 824.580 2.400 825.030 ;
        RECT 17.085 825.015 17.415 825.030 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 24.910 2608.380 25.230 2608.440 ;
        RECT 286.190 2608.380 286.510 2608.440 ;
        RECT 24.910 2608.240 286.510 2608.380 ;
        RECT 24.910 2608.180 25.230 2608.240 ;
        RECT 286.190 2608.180 286.510 2608.240 ;
        RECT 13.870 611.560 14.190 611.620 ;
        RECT 24.910 611.560 25.230 611.620 ;
        RECT 13.870 611.420 25.230 611.560 ;
        RECT 13.870 611.360 14.190 611.420 ;
        RECT 24.910 611.360 25.230 611.420 ;
      LAYER via ;
        RECT 24.940 2608.180 25.200 2608.440 ;
        RECT 286.220 2608.180 286.480 2608.440 ;
        RECT 13.900 611.360 14.160 611.620 ;
        RECT 24.940 611.360 25.200 611.620 ;
      LAYER met2 ;
        RECT 286.210 2609.995 286.490 2610.365 ;
        RECT 286.280 2608.470 286.420 2609.995 ;
        RECT 24.940 2608.150 25.200 2608.470 ;
        RECT 286.220 2608.150 286.480 2608.470 ;
        RECT 25.000 611.650 25.140 2608.150 ;
        RECT 13.900 611.330 14.160 611.650 ;
        RECT 24.940 611.330 25.200 611.650 ;
        RECT 13.960 610.485 14.100 611.330 ;
        RECT 13.890 610.115 14.170 610.485 ;
      LAYER via2 ;
        RECT 286.210 2610.040 286.490 2610.320 ;
        RECT 13.890 610.160 14.170 610.440 ;
      LAYER met3 ;
        RECT 286.185 2610.330 286.515 2610.345 ;
        RECT 300.000 2610.330 304.000 2610.400 ;
        RECT 286.185 2610.030 304.000 2610.330 ;
        RECT 286.185 2610.015 286.515 2610.030 ;
        RECT 300.000 2609.800 304.000 2610.030 ;
        RECT -4.800 610.450 2.400 610.900 ;
        RECT 13.865 610.450 14.195 610.465 ;
        RECT -4.800 610.150 14.195 610.450 ;
        RECT -4.800 609.700 2.400 610.150 ;
        RECT 13.865 610.135 14.195 610.150 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 24.450 2635.920 24.770 2635.980 ;
        RECT 286.190 2635.920 286.510 2635.980 ;
        RECT 24.450 2635.780 286.510 2635.920 ;
        RECT 24.450 2635.720 24.770 2635.780 ;
        RECT 286.190 2635.720 286.510 2635.780 ;
        RECT 13.870 399.060 14.190 399.120 ;
        RECT 24.450 399.060 24.770 399.120 ;
        RECT 13.870 398.920 24.770 399.060 ;
        RECT 13.870 398.860 14.190 398.920 ;
        RECT 24.450 398.860 24.770 398.920 ;
      LAYER via ;
        RECT 24.480 2635.720 24.740 2635.980 ;
        RECT 286.220 2635.720 286.480 2635.980 ;
        RECT 13.900 398.860 14.160 399.120 ;
        RECT 24.480 398.860 24.740 399.120 ;
      LAYER met2 ;
        RECT 286.210 2641.955 286.490 2642.325 ;
        RECT 286.280 2636.010 286.420 2641.955 ;
        RECT 24.480 2635.690 24.740 2636.010 ;
        RECT 286.220 2635.690 286.480 2636.010 ;
        RECT 24.540 399.150 24.680 2635.690 ;
        RECT 13.900 398.830 14.160 399.150 ;
        RECT 24.480 398.830 24.740 399.150 ;
        RECT 13.960 394.925 14.100 398.830 ;
        RECT 13.890 394.555 14.170 394.925 ;
      LAYER via2 ;
        RECT 286.210 2642.000 286.490 2642.280 ;
        RECT 13.890 394.600 14.170 394.880 ;
      LAYER met3 ;
        RECT 286.185 2642.290 286.515 2642.305 ;
        RECT 300.000 2642.290 304.000 2642.360 ;
        RECT 286.185 2641.990 304.000 2642.290 ;
        RECT 286.185 2641.975 286.515 2641.990 ;
        RECT 300.000 2641.760 304.000 2641.990 ;
        RECT -4.800 394.890 2.400 395.340 ;
        RECT 13.865 394.890 14.195 394.905 ;
        RECT -4.800 394.590 14.195 394.890 ;
        RECT -4.800 394.140 2.400 394.590 ;
        RECT 13.865 394.575 14.195 394.590 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 23.990 2670.600 24.310 2670.660 ;
        RECT 286.190 2670.600 286.510 2670.660 ;
        RECT 23.990 2670.460 286.510 2670.600 ;
        RECT 23.990 2670.400 24.310 2670.460 ;
        RECT 286.190 2670.400 286.510 2670.460 ;
        RECT 13.870 179.420 14.190 179.480 ;
        RECT 23.990 179.420 24.310 179.480 ;
        RECT 13.870 179.280 24.310 179.420 ;
        RECT 13.870 179.220 14.190 179.280 ;
        RECT 23.990 179.220 24.310 179.280 ;
      LAYER via ;
        RECT 24.020 2670.400 24.280 2670.660 ;
        RECT 286.220 2670.400 286.480 2670.660 ;
        RECT 13.900 179.220 14.160 179.480 ;
        RECT 24.020 179.220 24.280 179.480 ;
      LAYER met2 ;
        RECT 286.210 2673.235 286.490 2673.605 ;
        RECT 286.280 2670.690 286.420 2673.235 ;
        RECT 24.020 2670.370 24.280 2670.690 ;
        RECT 286.220 2670.370 286.480 2670.690 ;
        RECT 24.080 179.510 24.220 2670.370 ;
        RECT 13.900 179.365 14.160 179.510 ;
        RECT 13.890 178.995 14.170 179.365 ;
        RECT 24.020 179.190 24.280 179.510 ;
      LAYER via2 ;
        RECT 286.210 2673.280 286.490 2673.560 ;
        RECT 13.890 179.040 14.170 179.320 ;
      LAYER met3 ;
        RECT 286.185 2673.570 286.515 2673.585 ;
        RECT 300.000 2673.570 304.000 2673.640 ;
        RECT 286.185 2673.270 304.000 2673.570 ;
        RECT 286.185 2673.255 286.515 2673.270 ;
        RECT 300.000 2673.040 304.000 2673.270 ;
        RECT -4.800 179.330 2.400 179.780 ;
        RECT 13.865 179.330 14.195 179.345 ;
        RECT -4.800 179.030 14.195 179.330 ;
        RECT -4.800 178.580 2.400 179.030 ;
        RECT 13.865 179.015 14.195 179.030 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 296.770 793.460 297.090 793.520 ;
        RECT 2898.990 793.460 2899.310 793.520 ;
        RECT 296.770 793.320 2899.310 793.460 ;
        RECT 296.770 793.260 297.090 793.320 ;
        RECT 2898.990 793.260 2899.310 793.320 ;
      LAYER via ;
        RECT 296.800 793.260 297.060 793.520 ;
        RECT 2899.020 793.260 2899.280 793.520 ;
      LAYER met2 ;
        RECT 296.790 1599.515 297.070 1599.885 ;
        RECT 296.860 793.550 297.000 1599.515 ;
        RECT 296.800 793.230 297.060 793.550 ;
        RECT 2899.020 793.230 2899.280 793.550 ;
        RECT 2899.080 792.045 2899.220 793.230 ;
        RECT 2899.010 791.675 2899.290 792.045 ;
      LAYER via2 ;
        RECT 296.790 1599.560 297.070 1599.840 ;
        RECT 2899.010 791.720 2899.290 792.000 ;
      LAYER met3 ;
        RECT 296.765 1599.850 297.095 1599.865 ;
        RECT 300.000 1599.850 304.000 1599.920 ;
        RECT 296.765 1599.550 304.000 1599.850 ;
        RECT 296.765 1599.535 297.095 1599.550 ;
        RECT 300.000 1599.320 304.000 1599.550 ;
        RECT 2898.985 792.010 2899.315 792.025 ;
        RECT 2917.600 792.010 2924.800 792.460 ;
        RECT 2898.985 791.710 2924.800 792.010 ;
        RECT 2898.985 791.695 2899.315 791.710 ;
        RECT 2917.600 791.260 2924.800 791.710 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 287.110 1028.060 287.430 1028.120 ;
        RECT 2898.990 1028.060 2899.310 1028.120 ;
        RECT 287.110 1027.920 2899.310 1028.060 ;
        RECT 287.110 1027.860 287.430 1027.920 ;
        RECT 2898.990 1027.860 2899.310 1027.920 ;
      LAYER via ;
        RECT 287.140 1027.860 287.400 1028.120 ;
        RECT 2899.020 1027.860 2899.280 1028.120 ;
      LAYER met2 ;
        RECT 287.130 1630.795 287.410 1631.165 ;
        RECT 287.200 1028.150 287.340 1630.795 ;
        RECT 287.140 1027.830 287.400 1028.150 ;
        RECT 2899.020 1027.830 2899.280 1028.150 ;
        RECT 2899.080 1026.645 2899.220 1027.830 ;
        RECT 2899.010 1026.275 2899.290 1026.645 ;
      LAYER via2 ;
        RECT 287.130 1630.840 287.410 1631.120 ;
        RECT 2899.010 1026.320 2899.290 1026.600 ;
      LAYER met3 ;
        RECT 287.105 1631.130 287.435 1631.145 ;
        RECT 300.000 1631.130 304.000 1631.200 ;
        RECT 287.105 1630.830 304.000 1631.130 ;
        RECT 287.105 1630.815 287.435 1630.830 ;
        RECT 300.000 1630.600 304.000 1630.830 ;
        RECT 2898.985 1026.610 2899.315 1026.625 ;
        RECT 2917.600 1026.610 2924.800 1027.060 ;
        RECT 2898.985 1026.310 2924.800 1026.610 ;
        RECT 2898.985 1026.295 2899.315 1026.310 ;
        RECT 2917.600 1025.860 2924.800 1026.310 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 285.270 1262.660 285.590 1262.720 ;
        RECT 2898.990 1262.660 2899.310 1262.720 ;
        RECT 285.270 1262.520 2899.310 1262.660 ;
        RECT 285.270 1262.460 285.590 1262.520 ;
        RECT 2898.990 1262.460 2899.310 1262.520 ;
      LAYER via ;
        RECT 285.300 1262.460 285.560 1262.720 ;
        RECT 2899.020 1262.460 2899.280 1262.720 ;
      LAYER met2 ;
        RECT 285.290 1662.755 285.570 1663.125 ;
        RECT 285.360 1262.750 285.500 1662.755 ;
        RECT 285.300 1262.430 285.560 1262.750 ;
        RECT 2899.020 1262.430 2899.280 1262.750 ;
        RECT 2899.080 1261.245 2899.220 1262.430 ;
        RECT 2899.010 1260.875 2899.290 1261.245 ;
      LAYER via2 ;
        RECT 285.290 1662.800 285.570 1663.080 ;
        RECT 2899.010 1260.920 2899.290 1261.200 ;
      LAYER met3 ;
        RECT 285.265 1663.090 285.595 1663.105 ;
        RECT 300.000 1663.090 304.000 1663.160 ;
        RECT 285.265 1662.790 304.000 1663.090 ;
        RECT 285.265 1662.775 285.595 1662.790 ;
        RECT 300.000 1662.560 304.000 1662.790 ;
        RECT 2898.985 1261.210 2899.315 1261.225 ;
        RECT 2917.600 1261.210 2924.800 1261.660 ;
        RECT 2898.985 1260.910 2924.800 1261.210 ;
        RECT 2898.985 1260.895 2899.315 1260.910 ;
        RECT 2917.600 1260.460 2924.800 1260.910 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 283.890 1497.260 284.210 1497.320 ;
        RECT 2898.990 1497.260 2899.310 1497.320 ;
        RECT 283.890 1497.120 2899.310 1497.260 ;
        RECT 283.890 1497.060 284.210 1497.120 ;
        RECT 2898.990 1497.060 2899.310 1497.120 ;
      LAYER via ;
        RECT 283.920 1497.060 284.180 1497.320 ;
        RECT 2899.020 1497.060 2899.280 1497.320 ;
      LAYER met2 ;
        RECT 283.910 1694.035 284.190 1694.405 ;
        RECT 283.980 1497.350 284.120 1694.035 ;
        RECT 283.920 1497.030 284.180 1497.350 ;
        RECT 2899.020 1497.030 2899.280 1497.350 ;
        RECT 2899.080 1495.845 2899.220 1497.030 ;
        RECT 2899.010 1495.475 2899.290 1495.845 ;
      LAYER via2 ;
        RECT 283.910 1694.080 284.190 1694.360 ;
        RECT 2899.010 1495.520 2899.290 1495.800 ;
      LAYER met3 ;
        RECT 283.885 1694.370 284.215 1694.385 ;
        RECT 300.000 1694.370 304.000 1694.440 ;
        RECT 283.885 1694.070 304.000 1694.370 ;
        RECT 283.885 1694.055 284.215 1694.070 ;
        RECT 300.000 1693.840 304.000 1694.070 ;
        RECT 2898.985 1495.810 2899.315 1495.825 ;
        RECT 2917.600 1495.810 2924.800 1496.260 ;
        RECT 2898.985 1495.510 2924.800 1495.810 ;
        RECT 2898.985 1495.495 2899.315 1495.510 ;
        RECT 2917.600 1495.060 2924.800 1495.510 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2894.390 1700.920 2894.710 1700.980 ;
        RECT 2900.830 1700.920 2901.150 1700.980 ;
        RECT 2894.390 1700.780 2901.150 1700.920 ;
        RECT 2894.390 1700.720 2894.710 1700.780 ;
        RECT 2900.830 1700.720 2901.150 1700.780 ;
        RECT 2884.270 1642.100 2884.590 1642.160 ;
        RECT 2894.390 1642.100 2894.710 1642.160 ;
        RECT 2884.270 1641.960 2894.710 1642.100 ;
        RECT 2884.270 1641.900 2884.590 1641.960 ;
        RECT 2894.390 1641.900 2894.710 1641.960 ;
        RECT 288.030 1610.480 288.350 1610.540 ;
        RECT 296.310 1610.480 296.630 1610.540 ;
        RECT 288.030 1610.340 296.630 1610.480 ;
        RECT 288.030 1610.280 288.350 1610.340 ;
        RECT 296.310 1610.280 296.630 1610.340 ;
        RECT 2874.150 1594.160 2874.470 1594.220 ;
        RECT 2883.810 1594.160 2884.130 1594.220 ;
        RECT 2874.150 1594.020 2884.130 1594.160 ;
        RECT 2874.150 1593.960 2874.470 1594.020 ;
        RECT 2883.810 1593.960 2884.130 1594.020 ;
        RECT 2863.570 1585.320 2863.890 1585.380 ;
        RECT 2874.150 1585.320 2874.470 1585.380 ;
        RECT 2863.570 1585.180 2874.470 1585.320 ;
        RECT 2863.570 1585.120 2863.890 1585.180 ;
        RECT 2874.150 1585.120 2874.470 1585.180 ;
        RECT 2849.770 1545.880 2850.090 1545.940 ;
        RECT 2863.570 1545.880 2863.890 1545.940 ;
        RECT 2849.770 1545.740 2863.890 1545.880 ;
        RECT 2849.770 1545.680 2850.090 1545.740 ;
        RECT 2863.570 1545.680 2863.890 1545.740 ;
        RECT 2825.390 1542.140 2825.710 1542.200 ;
        RECT 2849.770 1542.140 2850.090 1542.200 ;
        RECT 2825.390 1542.000 2850.090 1542.140 ;
        RECT 2825.390 1541.940 2825.710 1542.000 ;
        RECT 2849.770 1541.940 2850.090 1542.000 ;
        RECT 296.310 1522.420 296.630 1522.480 ;
        RECT 297.230 1522.420 297.550 1522.480 ;
        RECT 296.310 1522.280 297.550 1522.420 ;
        RECT 296.310 1522.220 296.630 1522.280 ;
        RECT 297.230 1522.220 297.550 1522.280 ;
        RECT 297.230 1503.380 297.550 1503.440 ;
        RECT 2825.390 1503.380 2825.710 1503.440 ;
        RECT 297.230 1503.240 2825.710 1503.380 ;
        RECT 297.230 1503.180 297.550 1503.240 ;
        RECT 2825.390 1503.180 2825.710 1503.240 ;
      LAYER via ;
        RECT 2894.420 1700.720 2894.680 1700.980 ;
        RECT 2900.860 1700.720 2901.120 1700.980 ;
        RECT 2884.300 1641.900 2884.560 1642.160 ;
        RECT 2894.420 1641.900 2894.680 1642.160 ;
        RECT 288.060 1610.280 288.320 1610.540 ;
        RECT 296.340 1610.280 296.600 1610.540 ;
        RECT 2874.180 1593.960 2874.440 1594.220 ;
        RECT 2883.840 1593.960 2884.100 1594.220 ;
        RECT 2863.600 1585.120 2863.860 1585.380 ;
        RECT 2874.180 1585.120 2874.440 1585.380 ;
        RECT 2849.800 1545.680 2850.060 1545.940 ;
        RECT 2863.600 1545.680 2863.860 1545.940 ;
        RECT 2825.420 1541.940 2825.680 1542.200 ;
        RECT 2849.800 1541.940 2850.060 1542.200 ;
        RECT 296.340 1522.220 296.600 1522.480 ;
        RECT 297.260 1522.220 297.520 1522.480 ;
        RECT 297.260 1503.180 297.520 1503.440 ;
        RECT 2825.420 1503.180 2825.680 1503.440 ;
      LAYER met2 ;
        RECT 2900.850 1730.075 2901.130 1730.445 ;
        RECT 288.050 1725.995 288.330 1726.365 ;
        RECT 288.120 1610.570 288.260 1725.995 ;
        RECT 2900.920 1701.010 2901.060 1730.075 ;
        RECT 2894.420 1700.690 2894.680 1701.010 ;
        RECT 2900.860 1700.690 2901.120 1701.010 ;
        RECT 2894.480 1642.190 2894.620 1700.690 ;
        RECT 2884.300 1641.870 2884.560 1642.190 ;
        RECT 2894.420 1641.870 2894.680 1642.190 ;
        RECT 288.060 1610.250 288.320 1610.570 ;
        RECT 296.340 1610.250 296.600 1610.570 ;
        RECT 296.400 1522.510 296.540 1610.250 ;
        RECT 2884.360 1607.930 2884.500 1641.870 ;
        RECT 2883.900 1607.790 2884.500 1607.930 ;
        RECT 2883.900 1594.250 2884.040 1607.790 ;
        RECT 2874.180 1593.930 2874.440 1594.250 ;
        RECT 2883.840 1593.930 2884.100 1594.250 ;
        RECT 2874.240 1585.410 2874.380 1593.930 ;
        RECT 2863.600 1585.090 2863.860 1585.410 ;
        RECT 2874.180 1585.090 2874.440 1585.410 ;
        RECT 2863.660 1545.970 2863.800 1585.090 ;
        RECT 2849.800 1545.650 2850.060 1545.970 ;
        RECT 2863.600 1545.650 2863.860 1545.970 ;
        RECT 2849.860 1542.230 2850.000 1545.650 ;
        RECT 2825.420 1541.910 2825.680 1542.230 ;
        RECT 2849.800 1541.910 2850.060 1542.230 ;
        RECT 296.340 1522.190 296.600 1522.510 ;
        RECT 297.260 1522.190 297.520 1522.510 ;
        RECT 297.320 1503.470 297.460 1522.190 ;
        RECT 2825.480 1503.470 2825.620 1541.910 ;
        RECT 297.260 1503.150 297.520 1503.470 ;
        RECT 2825.420 1503.150 2825.680 1503.470 ;
      LAYER via2 ;
        RECT 2900.850 1730.120 2901.130 1730.400 ;
        RECT 288.050 1726.040 288.330 1726.320 ;
      LAYER met3 ;
        RECT 2900.825 1730.410 2901.155 1730.425 ;
        RECT 2917.600 1730.410 2924.800 1730.860 ;
        RECT 2900.825 1730.110 2924.800 1730.410 ;
        RECT 2900.825 1730.095 2901.155 1730.110 ;
        RECT 2917.600 1729.660 2924.800 1730.110 ;
        RECT 288.025 1726.330 288.355 1726.345 ;
        RECT 300.000 1726.330 304.000 1726.400 ;
        RECT 288.025 1726.030 304.000 1726.330 ;
        RECT 288.025 1726.015 288.355 1726.030 ;
        RECT 300.000 1725.800 304.000 1726.030 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2889.330 1960.000 2889.650 1960.060 ;
        RECT 2898.070 1960.000 2898.390 1960.060 ;
        RECT 2889.330 1959.860 2898.390 1960.000 ;
        RECT 2889.330 1959.800 2889.650 1959.860 ;
        RECT 2898.070 1959.800 2898.390 1959.860 ;
        RECT 2881.050 1925.320 2881.370 1925.380 ;
        RECT 2889.330 1925.320 2889.650 1925.380 ;
        RECT 2881.050 1925.180 2889.650 1925.320 ;
        RECT 2881.050 1925.120 2881.370 1925.180 ;
        RECT 2889.330 1925.120 2889.650 1925.180 ;
        RECT 2870.470 1911.380 2870.790 1911.440 ;
        RECT 2881.050 1911.380 2881.370 1911.440 ;
        RECT 2870.470 1911.240 2881.370 1911.380 ;
        RECT 2870.470 1911.180 2870.790 1911.240 ;
        RECT 2881.050 1911.180 2881.370 1911.240 ;
        RECT 2854.830 1881.800 2855.150 1881.860 ;
        RECT 2870.470 1881.800 2870.790 1881.860 ;
        RECT 2854.830 1881.660 2870.790 1881.800 ;
        RECT 2854.830 1881.600 2855.150 1881.660 ;
        RECT 2870.470 1881.600 2870.790 1881.660 ;
        RECT 2843.790 1858.000 2844.110 1858.060 ;
        RECT 2854.830 1858.000 2855.150 1858.060 ;
        RECT 2843.790 1857.860 2855.150 1858.000 ;
        RECT 2843.790 1857.800 2844.110 1857.860 ;
        RECT 2854.830 1857.800 2855.150 1857.860 ;
        RECT 2843.790 1849.500 2844.110 1849.560 ;
        RECT 2833.760 1849.360 2844.110 1849.500 ;
        RECT 2820.330 1849.160 2820.650 1849.220 ;
        RECT 2833.760 1849.160 2833.900 1849.360 ;
        RECT 2843.790 1849.300 2844.110 1849.360 ;
        RECT 2820.330 1849.020 2833.900 1849.160 ;
        RECT 2820.330 1848.960 2820.650 1849.020 ;
        RECT 2804.690 1835.560 2805.010 1835.620 ;
        RECT 2820.330 1835.560 2820.650 1835.620 ;
        RECT 2804.690 1835.420 2820.650 1835.560 ;
        RECT 2804.690 1835.360 2805.010 1835.420 ;
        RECT 2820.330 1835.360 2820.650 1835.420 ;
        RECT 2797.790 1742.060 2798.110 1742.120 ;
        RECT 2804.690 1742.060 2805.010 1742.120 ;
        RECT 2797.790 1741.920 2805.010 1742.060 ;
        RECT 2797.790 1741.860 2798.110 1741.920 ;
        RECT 2804.690 1741.860 2805.010 1741.920 ;
        RECT 2763.290 1626.800 2763.610 1626.860 ;
        RECT 2797.790 1626.800 2798.110 1626.860 ;
        RECT 2763.290 1626.660 2798.110 1626.800 ;
        RECT 2763.290 1626.600 2763.610 1626.660 ;
        RECT 2797.790 1626.600 2798.110 1626.660 ;
        RECT 2745.810 1614.900 2746.130 1614.960 ;
        RECT 2763.290 1614.900 2763.610 1614.960 ;
        RECT 2745.810 1614.760 2763.610 1614.900 ;
        RECT 2745.810 1614.700 2746.130 1614.760 ;
        RECT 2763.290 1614.700 2763.610 1614.760 ;
        RECT 2732.470 1598.920 2732.790 1598.980 ;
        RECT 2745.810 1598.920 2746.130 1598.980 ;
        RECT 2732.470 1598.780 2746.130 1598.920 ;
        RECT 2732.470 1598.720 2732.790 1598.780 ;
        RECT 2745.810 1598.720 2746.130 1598.780 ;
        RECT 287.570 1587.020 287.890 1587.080 ;
        RECT 292.170 1587.020 292.490 1587.080 ;
        RECT 287.570 1586.880 292.490 1587.020 ;
        RECT 287.570 1586.820 287.890 1586.880 ;
        RECT 292.170 1586.820 292.490 1586.880 ;
        RECT 2726.030 1583.280 2726.350 1583.340 ;
        RECT 2732.470 1583.280 2732.790 1583.340 ;
        RECT 2726.030 1583.140 2732.790 1583.280 ;
        RECT 2726.030 1583.080 2726.350 1583.140 ;
        RECT 2732.470 1583.080 2732.790 1583.140 ;
        RECT 2726.030 1559.480 2726.350 1559.540 ;
        RECT 2718.760 1559.340 2726.350 1559.480 ;
        RECT 2715.450 1559.140 2715.770 1559.200 ;
        RECT 2718.760 1559.140 2718.900 1559.340 ;
        RECT 2726.030 1559.280 2726.350 1559.340 ;
        RECT 2715.450 1559.000 2718.900 1559.140 ;
        RECT 2715.450 1558.940 2715.770 1559.000 ;
        RECT 2704.870 1525.140 2705.190 1525.200 ;
        RECT 2715.450 1525.140 2715.770 1525.200 ;
        RECT 2704.870 1525.000 2715.770 1525.140 ;
        RECT 2704.870 1524.940 2705.190 1525.000 ;
        RECT 2715.450 1524.940 2715.770 1525.000 ;
        RECT 292.170 1502.020 292.490 1502.080 ;
        RECT 2704.410 1502.020 2704.730 1502.080 ;
        RECT 292.170 1501.880 2704.730 1502.020 ;
        RECT 292.170 1501.820 292.490 1501.880 ;
        RECT 2704.410 1501.820 2704.730 1501.880 ;
      LAYER via ;
        RECT 2889.360 1959.800 2889.620 1960.060 ;
        RECT 2898.100 1959.800 2898.360 1960.060 ;
        RECT 2881.080 1925.120 2881.340 1925.380 ;
        RECT 2889.360 1925.120 2889.620 1925.380 ;
        RECT 2870.500 1911.180 2870.760 1911.440 ;
        RECT 2881.080 1911.180 2881.340 1911.440 ;
        RECT 2854.860 1881.600 2855.120 1881.860 ;
        RECT 2870.500 1881.600 2870.760 1881.860 ;
        RECT 2843.820 1857.800 2844.080 1858.060 ;
        RECT 2854.860 1857.800 2855.120 1858.060 ;
        RECT 2820.360 1848.960 2820.620 1849.220 ;
        RECT 2843.820 1849.300 2844.080 1849.560 ;
        RECT 2804.720 1835.360 2804.980 1835.620 ;
        RECT 2820.360 1835.360 2820.620 1835.620 ;
        RECT 2797.820 1741.860 2798.080 1742.120 ;
        RECT 2804.720 1741.860 2804.980 1742.120 ;
        RECT 2763.320 1626.600 2763.580 1626.860 ;
        RECT 2797.820 1626.600 2798.080 1626.860 ;
        RECT 2745.840 1614.700 2746.100 1614.960 ;
        RECT 2763.320 1614.700 2763.580 1614.960 ;
        RECT 2732.500 1598.720 2732.760 1598.980 ;
        RECT 2745.840 1598.720 2746.100 1598.980 ;
        RECT 287.600 1586.820 287.860 1587.080 ;
        RECT 292.200 1586.820 292.460 1587.080 ;
        RECT 2726.060 1583.080 2726.320 1583.340 ;
        RECT 2732.500 1583.080 2732.760 1583.340 ;
        RECT 2715.480 1558.940 2715.740 1559.200 ;
        RECT 2726.060 1559.280 2726.320 1559.540 ;
        RECT 2704.900 1524.940 2705.160 1525.200 ;
        RECT 2715.480 1524.940 2715.740 1525.200 ;
        RECT 292.200 1501.820 292.460 1502.080 ;
        RECT 2704.440 1501.820 2704.700 1502.080 ;
      LAYER met2 ;
        RECT 2898.090 1964.675 2898.370 1965.045 ;
        RECT 2898.160 1960.090 2898.300 1964.675 ;
        RECT 2889.360 1959.770 2889.620 1960.090 ;
        RECT 2898.100 1959.770 2898.360 1960.090 ;
        RECT 2889.420 1925.410 2889.560 1959.770 ;
        RECT 2881.080 1925.090 2881.340 1925.410 ;
        RECT 2889.360 1925.090 2889.620 1925.410 ;
        RECT 2881.140 1911.470 2881.280 1925.090 ;
        RECT 2870.500 1911.150 2870.760 1911.470 ;
        RECT 2881.080 1911.150 2881.340 1911.470 ;
        RECT 2870.560 1881.890 2870.700 1911.150 ;
        RECT 2854.860 1881.570 2855.120 1881.890 ;
        RECT 2870.500 1881.570 2870.760 1881.890 ;
        RECT 2854.920 1858.090 2855.060 1881.570 ;
        RECT 2843.820 1857.770 2844.080 1858.090 ;
        RECT 2854.860 1857.770 2855.120 1858.090 ;
        RECT 2843.880 1849.590 2844.020 1857.770 ;
        RECT 2843.820 1849.270 2844.080 1849.590 ;
        RECT 2820.360 1848.930 2820.620 1849.250 ;
        RECT 2820.420 1835.650 2820.560 1848.930 ;
        RECT 2804.720 1835.330 2804.980 1835.650 ;
        RECT 2820.360 1835.330 2820.620 1835.650 ;
        RECT 287.590 1757.275 287.870 1757.645 ;
        RECT 287.660 1587.110 287.800 1757.275 ;
        RECT 2804.780 1742.150 2804.920 1835.330 ;
        RECT 2797.820 1741.830 2798.080 1742.150 ;
        RECT 2804.720 1741.830 2804.980 1742.150 ;
        RECT 2797.880 1626.890 2798.020 1741.830 ;
        RECT 2763.320 1626.570 2763.580 1626.890 ;
        RECT 2797.820 1626.570 2798.080 1626.890 ;
        RECT 2763.380 1614.990 2763.520 1626.570 ;
        RECT 2745.840 1614.670 2746.100 1614.990 ;
        RECT 2763.320 1614.670 2763.580 1614.990 ;
        RECT 2745.900 1599.010 2746.040 1614.670 ;
        RECT 2732.500 1598.690 2732.760 1599.010 ;
        RECT 2745.840 1598.690 2746.100 1599.010 ;
        RECT 287.600 1586.790 287.860 1587.110 ;
        RECT 292.200 1586.790 292.460 1587.110 ;
        RECT 292.260 1502.110 292.400 1586.790 ;
        RECT 2732.560 1583.370 2732.700 1598.690 ;
        RECT 2726.060 1583.050 2726.320 1583.370 ;
        RECT 2732.500 1583.050 2732.760 1583.370 ;
        RECT 2726.120 1559.570 2726.260 1583.050 ;
        RECT 2726.060 1559.250 2726.320 1559.570 ;
        RECT 2715.480 1558.910 2715.740 1559.230 ;
        RECT 2715.540 1525.230 2715.680 1558.910 ;
        RECT 2704.900 1524.910 2705.160 1525.230 ;
        RECT 2715.480 1524.910 2715.740 1525.230 ;
        RECT 2704.960 1511.370 2705.100 1524.910 ;
        RECT 2704.500 1511.230 2705.100 1511.370 ;
        RECT 2704.500 1502.110 2704.640 1511.230 ;
        RECT 292.200 1501.790 292.460 1502.110 ;
        RECT 2704.440 1501.790 2704.700 1502.110 ;
      LAYER via2 ;
        RECT 2898.090 1964.720 2898.370 1965.000 ;
        RECT 287.590 1757.320 287.870 1757.600 ;
      LAYER met3 ;
        RECT 2898.065 1965.010 2898.395 1965.025 ;
        RECT 2917.600 1965.010 2924.800 1965.460 ;
        RECT 2898.065 1964.710 2924.800 1965.010 ;
        RECT 2898.065 1964.695 2898.395 1964.710 ;
        RECT 2917.600 1964.260 2924.800 1964.710 ;
        RECT 287.565 1757.610 287.895 1757.625 ;
        RECT 300.000 1757.610 304.000 1757.680 ;
        RECT 287.565 1757.310 304.000 1757.610 ;
        RECT 287.565 1757.295 287.895 1757.310 ;
        RECT 300.000 1757.080 304.000 1757.310 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2889.790 2188.140 2890.110 2188.200 ;
        RECT 2898.070 2188.140 2898.390 2188.200 ;
        RECT 2889.790 2188.000 2898.390 2188.140 ;
        RECT 2889.790 2187.940 2890.110 2188.000 ;
        RECT 2898.070 2187.940 2898.390 2188.000 ;
        RECT 2879.210 2177.600 2879.530 2177.660 ;
        RECT 2889.790 2177.600 2890.110 2177.660 ;
        RECT 2879.210 2177.460 2890.110 2177.600 ;
        RECT 2879.210 2177.400 2879.530 2177.460 ;
        RECT 2889.790 2177.400 2890.110 2177.460 ;
        RECT 2873.690 2162.640 2874.010 2162.700 ;
        RECT 2879.210 2162.640 2879.530 2162.700 ;
        RECT 2873.690 2162.500 2879.530 2162.640 ;
        RECT 2873.690 2162.440 2874.010 2162.500 ;
        RECT 2879.210 2162.440 2879.530 2162.500 ;
        RECT 2853.910 2113.680 2854.230 2113.740 ;
        RECT 2873.690 2113.680 2874.010 2113.740 ;
        RECT 2853.910 2113.540 2874.010 2113.680 ;
        RECT 2853.910 2113.480 2854.230 2113.540 ;
        RECT 2873.690 2113.480 2874.010 2113.540 ;
        RECT 2839.190 2097.700 2839.510 2097.760 ;
        RECT 2853.910 2097.700 2854.230 2097.760 ;
        RECT 2839.190 2097.560 2854.230 2097.700 ;
        RECT 2839.190 2097.500 2839.510 2097.560 ;
        RECT 2853.910 2097.500 2854.230 2097.560 ;
        RECT 2832.750 1960.000 2833.070 1960.060 ;
        RECT 2839.190 1960.000 2839.510 1960.060 ;
        RECT 2832.750 1959.860 2839.510 1960.000 ;
        RECT 2832.750 1959.800 2833.070 1959.860 ;
        RECT 2839.190 1959.800 2839.510 1959.860 ;
        RECT 2818.490 1842.360 2818.810 1842.420 ;
        RECT 2832.750 1842.360 2833.070 1842.420 ;
        RECT 2818.490 1842.220 2833.070 1842.360 ;
        RECT 2818.490 1842.160 2818.810 1842.220 ;
        RECT 2832.750 1842.160 2833.070 1842.220 ;
        RECT 2812.050 1785.240 2812.370 1785.300 ;
        RECT 2818.490 1785.240 2818.810 1785.300 ;
        RECT 2812.050 1785.100 2818.810 1785.240 ;
        RECT 2812.050 1785.040 2812.370 1785.100 ;
        RECT 2818.490 1785.040 2818.810 1785.100 ;
        RECT 2805.150 1752.940 2805.470 1753.000 ;
        RECT 2812.050 1752.940 2812.370 1753.000 ;
        RECT 2805.150 1752.800 2812.370 1752.940 ;
        RECT 2805.150 1752.740 2805.470 1752.800 ;
        RECT 2812.050 1752.740 2812.370 1752.800 ;
        RECT 2798.250 1718.260 2798.570 1718.320 ;
        RECT 2805.150 1718.260 2805.470 1718.320 ;
        RECT 2798.250 1718.120 2805.470 1718.260 ;
        RECT 2798.250 1718.060 2798.570 1718.120 ;
        RECT 2805.150 1718.060 2805.470 1718.120 ;
        RECT 287.110 1642.100 287.430 1642.160 ;
        RECT 294.470 1642.100 294.790 1642.160 ;
        RECT 287.110 1641.960 294.790 1642.100 ;
        RECT 287.110 1641.900 287.430 1641.960 ;
        RECT 294.470 1641.900 294.790 1641.960 ;
        RECT 2746.270 1638.700 2746.590 1638.760 ;
        RECT 2798.250 1638.700 2798.570 1638.760 ;
        RECT 2746.270 1638.560 2798.570 1638.700 ;
        RECT 2746.270 1638.500 2746.590 1638.560 ;
        RECT 2798.250 1638.500 2798.570 1638.560 ;
        RECT 2746.270 1608.100 2746.590 1608.160 ;
        RECT 2732.560 1607.960 2746.590 1608.100 ;
        RECT 2720.510 1607.420 2720.830 1607.480 ;
        RECT 2732.560 1607.420 2732.700 1607.960 ;
        RECT 2746.270 1607.900 2746.590 1607.960 ;
        RECT 2720.510 1607.280 2732.700 1607.420 ;
        RECT 2720.510 1607.220 2720.830 1607.280 ;
        RECT 2710.390 1584.980 2710.710 1585.040 ;
        RECT 2720.510 1584.980 2720.830 1585.040 ;
        RECT 2710.390 1584.840 2720.830 1584.980 ;
        RECT 2710.390 1584.780 2710.710 1584.840 ;
        RECT 2720.510 1584.780 2720.830 1584.840 ;
        RECT 2699.810 1559.820 2700.130 1559.880 ;
        RECT 2710.390 1559.820 2710.710 1559.880 ;
        RECT 2699.810 1559.680 2710.710 1559.820 ;
        RECT 2699.810 1559.620 2700.130 1559.680 ;
        RECT 2710.390 1559.620 2710.710 1559.680 ;
        RECT 2597.690 1548.940 2598.010 1549.000 ;
        RECT 2699.810 1548.940 2700.130 1549.000 ;
        RECT 2597.690 1548.800 2700.130 1548.940 ;
        RECT 2597.690 1548.740 2598.010 1548.800 ;
        RECT 2699.810 1548.740 2700.130 1548.800 ;
        RECT 2580.670 1525.140 2580.990 1525.200 ;
        RECT 2597.690 1525.140 2598.010 1525.200 ;
        RECT 2580.670 1525.000 2598.010 1525.140 ;
        RECT 2580.670 1524.940 2580.990 1525.000 ;
        RECT 2597.690 1524.940 2598.010 1525.000 ;
        RECT 294.470 1501.000 294.790 1501.060 ;
        RECT 2580.670 1501.000 2580.990 1501.060 ;
        RECT 294.470 1500.860 2580.990 1501.000 ;
        RECT 294.470 1500.800 294.790 1500.860 ;
        RECT 2580.670 1500.800 2580.990 1500.860 ;
      LAYER via ;
        RECT 2889.820 2187.940 2890.080 2188.200 ;
        RECT 2898.100 2187.940 2898.360 2188.200 ;
        RECT 2879.240 2177.400 2879.500 2177.660 ;
        RECT 2889.820 2177.400 2890.080 2177.660 ;
        RECT 2873.720 2162.440 2873.980 2162.700 ;
        RECT 2879.240 2162.440 2879.500 2162.700 ;
        RECT 2853.940 2113.480 2854.200 2113.740 ;
        RECT 2873.720 2113.480 2873.980 2113.740 ;
        RECT 2839.220 2097.500 2839.480 2097.760 ;
        RECT 2853.940 2097.500 2854.200 2097.760 ;
        RECT 2832.780 1959.800 2833.040 1960.060 ;
        RECT 2839.220 1959.800 2839.480 1960.060 ;
        RECT 2818.520 1842.160 2818.780 1842.420 ;
        RECT 2832.780 1842.160 2833.040 1842.420 ;
        RECT 2812.080 1785.040 2812.340 1785.300 ;
        RECT 2818.520 1785.040 2818.780 1785.300 ;
        RECT 2805.180 1752.740 2805.440 1753.000 ;
        RECT 2812.080 1752.740 2812.340 1753.000 ;
        RECT 2798.280 1718.060 2798.540 1718.320 ;
        RECT 2805.180 1718.060 2805.440 1718.320 ;
        RECT 287.140 1641.900 287.400 1642.160 ;
        RECT 294.500 1641.900 294.760 1642.160 ;
        RECT 2746.300 1638.500 2746.560 1638.760 ;
        RECT 2798.280 1638.500 2798.540 1638.760 ;
        RECT 2720.540 1607.220 2720.800 1607.480 ;
        RECT 2746.300 1607.900 2746.560 1608.160 ;
        RECT 2710.420 1584.780 2710.680 1585.040 ;
        RECT 2720.540 1584.780 2720.800 1585.040 ;
        RECT 2699.840 1559.620 2700.100 1559.880 ;
        RECT 2710.420 1559.620 2710.680 1559.880 ;
        RECT 2597.720 1548.740 2597.980 1549.000 ;
        RECT 2699.840 1548.740 2700.100 1549.000 ;
        RECT 2580.700 1524.940 2580.960 1525.200 ;
        RECT 2597.720 1524.940 2597.980 1525.200 ;
        RECT 294.500 1500.800 294.760 1501.060 ;
        RECT 2580.700 1500.800 2580.960 1501.060 ;
      LAYER met2 ;
        RECT 2898.090 2199.275 2898.370 2199.645 ;
        RECT 2898.160 2188.230 2898.300 2199.275 ;
        RECT 2889.820 2187.910 2890.080 2188.230 ;
        RECT 2898.100 2187.910 2898.360 2188.230 ;
        RECT 2889.880 2177.690 2890.020 2187.910 ;
        RECT 2879.240 2177.370 2879.500 2177.690 ;
        RECT 2889.820 2177.370 2890.080 2177.690 ;
        RECT 2879.300 2162.730 2879.440 2177.370 ;
        RECT 2873.720 2162.410 2873.980 2162.730 ;
        RECT 2879.240 2162.410 2879.500 2162.730 ;
        RECT 2873.780 2113.770 2873.920 2162.410 ;
        RECT 2853.940 2113.450 2854.200 2113.770 ;
        RECT 2873.720 2113.450 2873.980 2113.770 ;
        RECT 2854.000 2097.790 2854.140 2113.450 ;
        RECT 2839.220 2097.470 2839.480 2097.790 ;
        RECT 2853.940 2097.470 2854.200 2097.790 ;
        RECT 2839.280 1960.090 2839.420 2097.470 ;
        RECT 2832.780 1959.770 2833.040 1960.090 ;
        RECT 2839.220 1959.770 2839.480 1960.090 ;
        RECT 2832.840 1842.450 2832.980 1959.770 ;
        RECT 2818.520 1842.130 2818.780 1842.450 ;
        RECT 2832.780 1842.130 2833.040 1842.450 ;
        RECT 287.130 1789.235 287.410 1789.605 ;
        RECT 287.200 1642.190 287.340 1789.235 ;
        RECT 2818.580 1785.330 2818.720 1842.130 ;
        RECT 2812.080 1785.010 2812.340 1785.330 ;
        RECT 2818.520 1785.010 2818.780 1785.330 ;
        RECT 2812.140 1753.030 2812.280 1785.010 ;
        RECT 2805.180 1752.710 2805.440 1753.030 ;
        RECT 2812.080 1752.710 2812.340 1753.030 ;
        RECT 2805.240 1718.350 2805.380 1752.710 ;
        RECT 2798.280 1718.030 2798.540 1718.350 ;
        RECT 2805.180 1718.030 2805.440 1718.350 ;
        RECT 287.140 1641.870 287.400 1642.190 ;
        RECT 294.500 1641.870 294.760 1642.190 ;
        RECT 294.560 1501.090 294.700 1641.870 ;
        RECT 2798.340 1638.790 2798.480 1718.030 ;
        RECT 2746.300 1638.470 2746.560 1638.790 ;
        RECT 2798.280 1638.470 2798.540 1638.790 ;
        RECT 2746.360 1608.190 2746.500 1638.470 ;
        RECT 2746.300 1607.870 2746.560 1608.190 ;
        RECT 2720.540 1607.190 2720.800 1607.510 ;
        RECT 2720.600 1585.070 2720.740 1607.190 ;
        RECT 2710.420 1584.750 2710.680 1585.070 ;
        RECT 2720.540 1584.750 2720.800 1585.070 ;
        RECT 2710.480 1559.910 2710.620 1584.750 ;
        RECT 2699.840 1559.590 2700.100 1559.910 ;
        RECT 2710.420 1559.590 2710.680 1559.910 ;
        RECT 2699.900 1549.030 2700.040 1559.590 ;
        RECT 2597.720 1548.710 2597.980 1549.030 ;
        RECT 2699.840 1548.710 2700.100 1549.030 ;
        RECT 2597.780 1525.230 2597.920 1548.710 ;
        RECT 2580.700 1524.910 2580.960 1525.230 ;
        RECT 2597.720 1524.910 2597.980 1525.230 ;
        RECT 2580.760 1501.090 2580.900 1524.910 ;
        RECT 294.500 1500.770 294.760 1501.090 ;
        RECT 2580.700 1500.770 2580.960 1501.090 ;
      LAYER via2 ;
        RECT 2898.090 2199.320 2898.370 2199.600 ;
        RECT 287.130 1789.280 287.410 1789.560 ;
      LAYER met3 ;
        RECT 2898.065 2199.610 2898.395 2199.625 ;
        RECT 2917.600 2199.610 2924.800 2200.060 ;
        RECT 2898.065 2199.310 2924.800 2199.610 ;
        RECT 2898.065 2199.295 2898.395 2199.310 ;
        RECT 2917.600 2198.860 2924.800 2199.310 ;
        RECT 287.105 1789.570 287.435 1789.585 ;
        RECT 300.000 1789.570 304.000 1789.640 ;
        RECT 287.105 1789.270 304.000 1789.570 ;
        RECT 287.105 1789.255 287.435 1789.270 ;
        RECT 300.000 1789.040 304.000 1789.270 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 737.910 201.180 738.230 201.240 ;
        RECT 772.410 201.180 772.730 201.240 ;
        RECT 737.910 201.040 772.730 201.180 ;
        RECT 737.910 200.980 738.230 201.040 ;
        RECT 772.410 200.980 772.730 201.040 ;
        RECT 447.650 200.840 447.970 200.900 ;
        RECT 458.690 200.840 459.010 200.900 ;
        RECT 447.650 200.700 459.010 200.840 ;
        RECT 447.650 200.640 447.970 200.700 ;
        RECT 458.690 200.640 459.010 200.700 ;
        RECT 579.670 200.500 579.990 200.560 ;
        RECT 594.390 200.500 594.710 200.560 ;
        RECT 579.670 200.360 594.710 200.500 ;
        RECT 579.670 200.300 579.990 200.360 ;
        RECT 594.390 200.300 594.710 200.360 ;
      LAYER via ;
        RECT 737.940 200.980 738.200 201.240 ;
        RECT 772.440 200.980 772.700 201.240 ;
        RECT 447.680 200.640 447.940 200.900 ;
        RECT 458.720 200.640 458.980 200.900 ;
        RECT 579.700 200.300 579.960 200.560 ;
        RECT 594.420 200.300 594.680 200.560 ;
      LAYER met2 ;
        RECT 675.830 202.795 676.110 203.165 ;
        RECT 386.030 201.435 386.310 201.805 ;
        RECT 594.410 201.435 594.690 201.805 ;
        RECT 386.100 199.765 386.240 201.435 ;
        RECT 447.670 200.755 447.950 201.125 ;
        RECT 458.710 200.755 458.990 201.125 ;
        RECT 447.680 200.610 447.940 200.755 ;
        RECT 458.720 200.610 458.980 200.755 ;
        RECT 594.480 200.590 594.620 201.435 ;
        RECT 675.900 201.125 676.040 202.795 ;
        RECT 700.210 202.115 700.490 202.485 ;
        RECT 675.830 200.755 676.110 201.125 ;
        RECT 579.700 200.445 579.960 200.590 ;
        RECT 579.690 200.075 579.970 200.445 ;
        RECT 594.420 200.270 594.680 200.590 ;
        RECT 700.280 200.445 700.420 202.115 ;
        RECT 772.430 201.435 772.710 201.805 ;
        RECT 772.500 201.270 772.640 201.435 ;
        RECT 737.940 201.125 738.200 201.270 ;
        RECT 737.930 200.755 738.210 201.125 ;
        RECT 772.440 200.950 772.700 201.270 ;
        RECT 700.210 200.075 700.490 200.445 ;
        RECT 386.030 199.395 386.310 199.765 ;
      LAYER via2 ;
        RECT 675.830 202.840 676.110 203.120 ;
        RECT 386.030 201.480 386.310 201.760 ;
        RECT 594.410 201.480 594.690 201.760 ;
        RECT 447.670 200.800 447.950 201.080 ;
        RECT 458.710 200.800 458.990 201.080 ;
        RECT 700.210 202.160 700.490 202.440 ;
        RECT 675.830 200.800 676.110 201.080 ;
        RECT 579.690 200.120 579.970 200.400 ;
        RECT 772.430 201.480 772.710 201.760 ;
        RECT 737.930 200.800 738.210 201.080 ;
        RECT 700.210 200.120 700.490 200.400 ;
        RECT 386.030 199.440 386.310 199.720 ;
      LAYER met3 ;
        RECT 288.230 1515.530 288.610 1515.540 ;
        RECT 300.000 1515.530 304.000 1515.600 ;
        RECT 288.230 1515.230 304.000 1515.530 ;
        RECT 288.230 1515.220 288.610 1515.230 ;
        RECT 300.000 1515.000 304.000 1515.230 ;
        RECT 2917.600 205.170 2924.800 205.620 ;
        RECT 2916.710 204.870 2924.800 205.170 ;
        RECT 627.710 203.130 628.090 203.140 ;
        RECT 675.805 203.130 676.135 203.145 ;
        RECT 627.710 202.830 676.135 203.130 ;
        RECT 627.710 202.820 628.090 202.830 ;
        RECT 675.805 202.815 676.135 202.830 ;
        RECT 578.950 202.450 579.330 202.460 ;
        RECT 700.185 202.450 700.515 202.465 ;
        RECT 544.030 202.150 579.330 202.450 ;
        RECT 288.230 201.770 288.610 201.780 ;
        RECT 386.005 201.770 386.335 201.785 ;
        RECT 288.230 201.470 303.290 201.770 ;
        RECT 288.230 201.460 288.610 201.470 ;
        RECT 302.990 200.410 303.290 201.470 ;
        RECT 386.005 201.470 399.890 201.770 ;
        RECT 386.005 201.455 386.335 201.470 ;
        RECT 337.910 201.090 338.290 201.100 ;
        RECT 303.910 200.790 338.290 201.090 ;
        RECT 303.910 200.410 304.210 200.790 ;
        RECT 337.910 200.780 338.290 200.790 ;
        RECT 302.990 200.110 304.210 200.410 ;
        RECT 399.590 200.410 399.890 201.470 ;
        RECT 447.645 201.090 447.975 201.105 ;
        RECT 400.510 200.790 447.975 201.090 ;
        RECT 400.510 200.410 400.810 200.790 ;
        RECT 447.645 200.775 447.975 200.790 ;
        RECT 458.685 201.090 459.015 201.105 ;
        RECT 544.030 201.090 544.330 202.150 ;
        RECT 578.950 202.140 579.330 202.150 ;
        RECT 676.510 202.150 700.515 202.450 ;
        RECT 594.385 201.770 594.715 201.785 ;
        RECT 627.710 201.770 628.090 201.780 ;
        RECT 594.385 201.470 628.090 201.770 ;
        RECT 594.385 201.455 594.715 201.470 ;
        RECT 627.710 201.460 628.090 201.470 ;
        RECT 458.685 200.790 482.690 201.090 ;
        RECT 458.685 200.775 459.015 200.790 ;
        RECT 399.590 200.110 400.810 200.410 ;
        RECT 482.390 200.410 482.690 200.790 ;
        RECT 497.110 200.790 544.330 201.090 ;
        RECT 675.805 201.090 676.135 201.105 ;
        RECT 676.510 201.090 676.810 202.150 ;
        RECT 700.185 202.135 700.515 202.150 ;
        RECT 772.405 201.770 772.735 201.785 ;
        RECT 772.405 201.470 807.450 201.770 ;
        RECT 772.405 201.455 772.735 201.470 ;
        RECT 737.905 201.090 738.235 201.105 ;
        RECT 675.805 200.790 676.810 201.090 ;
        RECT 724.350 200.790 738.235 201.090 ;
        RECT 807.150 201.090 807.450 201.470 ;
        RECT 855.910 201.470 904.050 201.770 ;
        RECT 807.150 200.790 855.290 201.090 ;
        RECT 497.110 200.410 497.410 200.790 ;
        RECT 675.805 200.775 676.135 200.790 ;
        RECT 482.390 200.110 497.410 200.410 ;
        RECT 578.950 200.410 579.330 200.420 ;
        RECT 579.665 200.410 579.995 200.425 ;
        RECT 578.950 200.110 579.995 200.410 ;
        RECT 578.950 200.100 579.330 200.110 ;
        RECT 579.665 200.095 579.995 200.110 ;
        RECT 700.185 200.410 700.515 200.425 ;
        RECT 724.350 200.410 724.650 200.790 ;
        RECT 737.905 200.775 738.235 200.790 ;
        RECT 700.185 200.110 724.650 200.410 ;
        RECT 854.990 200.410 855.290 200.790 ;
        RECT 855.910 200.410 856.210 201.470 ;
        RECT 903.750 201.090 904.050 201.470 ;
        RECT 952.510 201.470 1000.650 201.770 ;
        RECT 903.750 200.790 951.890 201.090 ;
        RECT 854.990 200.110 856.210 200.410 ;
        RECT 951.590 200.410 951.890 200.790 ;
        RECT 952.510 200.410 952.810 201.470 ;
        RECT 1000.350 201.090 1000.650 201.470 ;
        RECT 1049.110 201.470 1097.250 201.770 ;
        RECT 1000.350 200.790 1048.490 201.090 ;
        RECT 951.590 200.110 952.810 200.410 ;
        RECT 1048.190 200.410 1048.490 200.790 ;
        RECT 1049.110 200.410 1049.410 201.470 ;
        RECT 1096.950 201.090 1097.250 201.470 ;
        RECT 1145.710 201.470 1193.850 201.770 ;
        RECT 1096.950 200.790 1145.090 201.090 ;
        RECT 1048.190 200.110 1049.410 200.410 ;
        RECT 1144.790 200.410 1145.090 200.790 ;
        RECT 1145.710 200.410 1146.010 201.470 ;
        RECT 1193.550 201.090 1193.850 201.470 ;
        RECT 1242.310 201.470 1290.450 201.770 ;
        RECT 1193.550 200.790 1241.690 201.090 ;
        RECT 1144.790 200.110 1146.010 200.410 ;
        RECT 1241.390 200.410 1241.690 200.790 ;
        RECT 1242.310 200.410 1242.610 201.470 ;
        RECT 1290.150 201.090 1290.450 201.470 ;
        RECT 1338.910 201.470 1387.050 201.770 ;
        RECT 1290.150 200.790 1338.290 201.090 ;
        RECT 1241.390 200.110 1242.610 200.410 ;
        RECT 1337.990 200.410 1338.290 200.790 ;
        RECT 1338.910 200.410 1339.210 201.470 ;
        RECT 1386.750 201.090 1387.050 201.470 ;
        RECT 1435.510 201.470 1483.650 201.770 ;
        RECT 1386.750 200.790 1434.890 201.090 ;
        RECT 1337.990 200.110 1339.210 200.410 ;
        RECT 1434.590 200.410 1434.890 200.790 ;
        RECT 1435.510 200.410 1435.810 201.470 ;
        RECT 1483.350 201.090 1483.650 201.470 ;
        RECT 1532.110 201.470 1580.250 201.770 ;
        RECT 1483.350 200.790 1531.490 201.090 ;
        RECT 1434.590 200.110 1435.810 200.410 ;
        RECT 1531.190 200.410 1531.490 200.790 ;
        RECT 1532.110 200.410 1532.410 201.470 ;
        RECT 1579.950 201.090 1580.250 201.470 ;
        RECT 1628.710 201.470 1676.850 201.770 ;
        RECT 1579.950 200.790 1628.090 201.090 ;
        RECT 1531.190 200.110 1532.410 200.410 ;
        RECT 1627.790 200.410 1628.090 200.790 ;
        RECT 1628.710 200.410 1629.010 201.470 ;
        RECT 1676.550 201.090 1676.850 201.470 ;
        RECT 1725.310 201.470 1773.450 201.770 ;
        RECT 1676.550 200.790 1724.690 201.090 ;
        RECT 1627.790 200.110 1629.010 200.410 ;
        RECT 1724.390 200.410 1724.690 200.790 ;
        RECT 1725.310 200.410 1725.610 201.470 ;
        RECT 1773.150 201.090 1773.450 201.470 ;
        RECT 1821.910 201.470 1870.050 201.770 ;
        RECT 1773.150 200.790 1821.290 201.090 ;
        RECT 1724.390 200.110 1725.610 200.410 ;
        RECT 1820.990 200.410 1821.290 200.790 ;
        RECT 1821.910 200.410 1822.210 201.470 ;
        RECT 1869.750 201.090 1870.050 201.470 ;
        RECT 1918.510 201.470 1966.650 201.770 ;
        RECT 1869.750 200.790 1917.890 201.090 ;
        RECT 1820.990 200.110 1822.210 200.410 ;
        RECT 1917.590 200.410 1917.890 200.790 ;
        RECT 1918.510 200.410 1918.810 201.470 ;
        RECT 1966.350 201.090 1966.650 201.470 ;
        RECT 2015.110 201.470 2063.250 201.770 ;
        RECT 1966.350 200.790 2014.490 201.090 ;
        RECT 1917.590 200.110 1918.810 200.410 ;
        RECT 2014.190 200.410 2014.490 200.790 ;
        RECT 2015.110 200.410 2015.410 201.470 ;
        RECT 2062.950 201.090 2063.250 201.470 ;
        RECT 2111.710 201.470 2159.850 201.770 ;
        RECT 2062.950 200.790 2111.090 201.090 ;
        RECT 2014.190 200.110 2015.410 200.410 ;
        RECT 2110.790 200.410 2111.090 200.790 ;
        RECT 2111.710 200.410 2112.010 201.470 ;
        RECT 2159.550 201.090 2159.850 201.470 ;
        RECT 2208.310 201.470 2256.450 201.770 ;
        RECT 2159.550 200.790 2207.690 201.090 ;
        RECT 2110.790 200.110 2112.010 200.410 ;
        RECT 2207.390 200.410 2207.690 200.790 ;
        RECT 2208.310 200.410 2208.610 201.470 ;
        RECT 2256.150 201.090 2256.450 201.470 ;
        RECT 2304.910 201.470 2353.050 201.770 ;
        RECT 2256.150 200.790 2304.290 201.090 ;
        RECT 2207.390 200.110 2208.610 200.410 ;
        RECT 2303.990 200.410 2304.290 200.790 ;
        RECT 2304.910 200.410 2305.210 201.470 ;
        RECT 2352.750 201.090 2353.050 201.470 ;
        RECT 2401.510 201.470 2449.650 201.770 ;
        RECT 2352.750 200.790 2400.890 201.090 ;
        RECT 2303.990 200.110 2305.210 200.410 ;
        RECT 2400.590 200.410 2400.890 200.790 ;
        RECT 2401.510 200.410 2401.810 201.470 ;
        RECT 2449.350 201.090 2449.650 201.470 ;
        RECT 2498.110 201.470 2546.250 201.770 ;
        RECT 2449.350 200.790 2497.490 201.090 ;
        RECT 2400.590 200.110 2401.810 200.410 ;
        RECT 2497.190 200.410 2497.490 200.790 ;
        RECT 2498.110 200.410 2498.410 201.470 ;
        RECT 2545.950 201.090 2546.250 201.470 ;
        RECT 2594.710 201.470 2642.850 201.770 ;
        RECT 2545.950 200.790 2594.090 201.090 ;
        RECT 2497.190 200.110 2498.410 200.410 ;
        RECT 2593.790 200.410 2594.090 200.790 ;
        RECT 2594.710 200.410 2595.010 201.470 ;
        RECT 2642.550 201.090 2642.850 201.470 ;
        RECT 2691.310 201.470 2739.450 201.770 ;
        RECT 2642.550 200.790 2690.690 201.090 ;
        RECT 2593.790 200.110 2595.010 200.410 ;
        RECT 2690.390 200.410 2690.690 200.790 ;
        RECT 2691.310 200.410 2691.610 201.470 ;
        RECT 2739.150 201.090 2739.450 201.470 ;
        RECT 2787.910 201.470 2836.050 201.770 ;
        RECT 2739.150 200.790 2787.290 201.090 ;
        RECT 2690.390 200.110 2691.610 200.410 ;
        RECT 2786.990 200.410 2787.290 200.790 ;
        RECT 2787.910 200.410 2788.210 201.470 ;
        RECT 2835.750 201.090 2836.050 201.470 ;
        RECT 2916.710 201.090 2917.010 204.870 ;
        RECT 2917.600 204.420 2924.800 204.870 ;
        RECT 2835.750 200.790 2883.890 201.090 ;
        RECT 2786.990 200.110 2788.210 200.410 ;
        RECT 2883.590 200.410 2883.890 200.790 ;
        RECT 2884.510 200.790 2917.010 201.090 ;
        RECT 2884.510 200.410 2884.810 200.790 ;
        RECT 2883.590 200.110 2884.810 200.410 ;
        RECT 700.185 200.095 700.515 200.110 ;
        RECT 337.910 199.730 338.290 199.740 ;
        RECT 386.005 199.730 386.335 199.745 ;
        RECT 337.910 199.430 386.335 199.730 ;
        RECT 337.910 199.420 338.290 199.430 ;
        RECT 386.005 199.415 386.335 199.430 ;
      LAYER via3 ;
        RECT 288.260 1515.220 288.580 1515.540 ;
        RECT 627.740 202.820 628.060 203.140 ;
        RECT 288.260 201.460 288.580 201.780 ;
        RECT 337.940 200.780 338.260 201.100 ;
        RECT 578.980 202.140 579.300 202.460 ;
        RECT 627.740 201.460 628.060 201.780 ;
        RECT 578.980 200.100 579.300 200.420 ;
        RECT 337.940 199.420 338.260 199.740 ;
      LAYER met4 ;
        RECT 288.255 1515.215 288.585 1515.545 ;
        RECT 288.270 201.785 288.570 1515.215 ;
        RECT 627.735 202.815 628.065 203.145 ;
        RECT 578.975 202.135 579.305 202.465 ;
        RECT 288.255 201.455 288.585 201.785 ;
        RECT 337.935 200.775 338.265 201.105 ;
        RECT 337.950 199.745 338.250 200.775 ;
        RECT 578.990 200.425 579.290 202.135 ;
        RECT 627.750 201.785 628.050 202.815 ;
        RECT 627.735 201.455 628.065 201.785 ;
        RECT 578.975 200.095 579.305 200.425 ;
        RECT 337.935 199.415 338.265 199.745 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 285.730 2689.640 286.050 2689.700 ;
        RECT 2901.290 2689.640 2901.610 2689.700 ;
        RECT 285.730 2689.500 2901.610 2689.640 ;
        RECT 285.730 2689.440 286.050 2689.500 ;
        RECT 2901.290 2689.440 2901.610 2689.500 ;
      LAYER via ;
        RECT 285.760 2689.440 286.020 2689.700 ;
        RECT 2901.320 2689.440 2901.580 2689.700 ;
      LAYER met2 ;
        RECT 285.760 2689.410 286.020 2689.730 ;
        RECT 2901.320 2689.410 2901.580 2689.730 ;
        RECT 285.820 1831.085 285.960 2689.410 ;
        RECT 2901.380 2551.885 2901.520 2689.410 ;
        RECT 2901.310 2551.515 2901.590 2551.885 ;
        RECT 285.750 1830.715 286.030 1831.085 ;
      LAYER via2 ;
        RECT 2901.310 2551.560 2901.590 2551.840 ;
        RECT 285.750 1830.760 286.030 1831.040 ;
      LAYER met3 ;
        RECT 2901.285 2551.850 2901.615 2551.865 ;
        RECT 2917.600 2551.850 2924.800 2552.300 ;
        RECT 2901.285 2551.550 2924.800 2551.850 ;
        RECT 2901.285 2551.535 2901.615 2551.550 ;
        RECT 2917.600 2551.100 2924.800 2551.550 ;
        RECT 285.725 1831.050 286.055 1831.065 ;
        RECT 300.000 1831.050 304.000 1831.120 ;
        RECT 285.725 1830.750 304.000 1831.050 ;
        RECT 285.725 1830.735 286.055 1830.750 ;
        RECT 300.000 1830.520 304.000 1830.750 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 291.250 2781.100 291.570 2781.160 ;
        RECT 2898.070 2781.100 2898.390 2781.160 ;
        RECT 291.250 2780.960 2898.390 2781.100 ;
        RECT 291.250 2780.900 291.570 2780.960 ;
        RECT 2898.070 2780.900 2898.390 2780.960 ;
      LAYER via ;
        RECT 291.280 2780.900 291.540 2781.160 ;
        RECT 2898.100 2780.900 2898.360 2781.160 ;
      LAYER met2 ;
        RECT 2898.090 2786.115 2898.370 2786.485 ;
        RECT 2898.160 2781.190 2898.300 2786.115 ;
        RECT 291.280 2780.870 291.540 2781.190 ;
        RECT 2898.100 2780.870 2898.360 2781.190 ;
        RECT 291.340 1863.045 291.480 2780.870 ;
        RECT 291.270 1862.675 291.550 1863.045 ;
      LAYER via2 ;
        RECT 2898.090 2786.160 2898.370 2786.440 ;
        RECT 291.270 1862.720 291.550 1863.000 ;
      LAYER met3 ;
        RECT 2898.065 2786.450 2898.395 2786.465 ;
        RECT 2917.600 2786.450 2924.800 2786.900 ;
        RECT 2898.065 2786.150 2924.800 2786.450 ;
        RECT 2898.065 2786.135 2898.395 2786.150 ;
        RECT 2917.600 2785.700 2924.800 2786.150 ;
        RECT 291.245 1863.010 291.575 1863.025 ;
        RECT 300.000 1863.010 304.000 1863.080 ;
        RECT 291.245 1862.710 304.000 1863.010 ;
        RECT 291.245 1862.695 291.575 1862.710 ;
        RECT 300.000 1862.480 304.000 1862.710 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2902.230 3020.715 2902.510 3021.085 ;
        RECT 2902.300 2695.365 2902.440 3020.715 ;
        RECT 2902.230 2694.995 2902.510 2695.365 ;
      LAYER via2 ;
        RECT 2902.230 3020.760 2902.510 3021.040 ;
        RECT 2902.230 2695.040 2902.510 2695.320 ;
      LAYER met3 ;
        RECT 2902.205 3021.050 2902.535 3021.065 ;
        RECT 2917.600 3021.050 2924.800 3021.500 ;
        RECT 2902.205 3020.750 2924.800 3021.050 ;
        RECT 2902.205 3020.735 2902.535 3020.750 ;
        RECT 2917.600 3020.300 2924.800 3020.750 ;
        RECT 288.230 2695.330 288.610 2695.340 ;
        RECT 2902.205 2695.330 2902.535 2695.345 ;
        RECT 288.230 2695.030 2902.535 2695.330 ;
        RECT 288.230 2695.020 288.610 2695.030 ;
        RECT 2902.205 2695.015 2902.535 2695.030 ;
        RECT 288.230 1894.290 288.610 1894.300 ;
        RECT 300.000 1894.290 304.000 1894.360 ;
        RECT 288.230 1893.990 304.000 1894.290 ;
        RECT 288.230 1893.980 288.610 1893.990 ;
        RECT 300.000 1893.760 304.000 1893.990 ;
      LAYER via3 ;
        RECT 288.260 2695.020 288.580 2695.340 ;
        RECT 288.260 1893.980 288.580 1894.300 ;
      LAYER met4 ;
        RECT 288.255 2695.015 288.585 2695.345 ;
        RECT 288.270 1894.305 288.570 2695.015 ;
        RECT 288.255 1893.975 288.585 1894.305 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 293.090 3251.660 293.410 3251.720 ;
        RECT 2900.830 3251.660 2901.150 3251.720 ;
        RECT 293.090 3251.520 2901.150 3251.660 ;
        RECT 293.090 3251.460 293.410 3251.520 ;
        RECT 2900.830 3251.460 2901.150 3251.520 ;
      LAYER via ;
        RECT 293.120 3251.460 293.380 3251.720 ;
        RECT 2900.860 3251.460 2901.120 3251.720 ;
      LAYER met2 ;
        RECT 2900.850 3255.315 2901.130 3255.685 ;
        RECT 2900.920 3251.750 2901.060 3255.315 ;
        RECT 293.120 3251.430 293.380 3251.750 ;
        RECT 2900.860 3251.430 2901.120 3251.750 ;
        RECT 293.180 1926.285 293.320 3251.430 ;
        RECT 293.110 1925.915 293.390 1926.285 ;
      LAYER via2 ;
        RECT 2900.850 3255.360 2901.130 3255.640 ;
        RECT 293.110 1925.960 293.390 1926.240 ;
      LAYER met3 ;
        RECT 2900.825 3255.650 2901.155 3255.665 ;
        RECT 2917.600 3255.650 2924.800 3256.100 ;
        RECT 2900.825 3255.350 2924.800 3255.650 ;
        RECT 2900.825 3255.335 2901.155 3255.350 ;
        RECT 2917.600 3254.900 2924.800 3255.350 ;
        RECT 293.085 1926.250 293.415 1926.265 ;
        RECT 300.000 1926.250 304.000 1926.320 ;
        RECT 293.085 1925.950 304.000 1926.250 ;
        RECT 293.085 1925.935 293.415 1925.950 ;
        RECT 300.000 1925.720 304.000 1925.950 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2801.470 3486.600 2801.790 3486.660 ;
        RECT 2825.850 3486.600 2826.170 3486.660 ;
        RECT 2801.470 3486.460 2826.170 3486.600 ;
        RECT 2801.470 3486.400 2801.790 3486.460 ;
        RECT 2825.850 3486.400 2826.170 3486.460 ;
        RECT 834.510 3485.920 834.830 3485.980 ;
        RECT 862.110 3485.920 862.430 3485.980 ;
        RECT 834.510 3485.780 862.430 3485.920 ;
        RECT 834.510 3485.720 834.830 3485.780 ;
        RECT 862.110 3485.720 862.430 3485.780 ;
        RECT 2704.870 3485.920 2705.190 3485.980 ;
        RECT 2743.050 3485.920 2743.370 3485.980 ;
        RECT 2704.870 3485.780 2743.370 3485.920 ;
        RECT 2704.870 3485.720 2705.190 3485.780 ;
        RECT 2743.050 3485.720 2743.370 3485.780 ;
        RECT 351.510 3485.580 351.830 3485.640 ;
        RECT 386.010 3485.580 386.330 3485.640 ;
        RECT 351.510 3485.440 386.330 3485.580 ;
        RECT 351.510 3485.380 351.830 3485.440 ;
        RECT 386.010 3485.380 386.330 3485.440 ;
        RECT 448.110 3485.580 448.430 3485.640 ;
        RECT 482.610 3485.580 482.930 3485.640 ;
        RECT 448.110 3485.440 482.930 3485.580 ;
        RECT 448.110 3485.380 448.430 3485.440 ;
        RECT 482.610 3485.380 482.930 3485.440 ;
        RECT 544.710 3485.580 545.030 3485.640 ;
        RECT 579.210 3485.580 579.530 3485.640 ;
        RECT 544.710 3485.440 579.530 3485.580 ;
        RECT 544.710 3485.380 545.030 3485.440 ;
        RECT 579.210 3485.380 579.530 3485.440 ;
        RECT 641.310 3485.580 641.630 3485.640 ;
        RECT 675.810 3485.580 676.130 3485.640 ;
        RECT 641.310 3485.440 676.130 3485.580 ;
        RECT 641.310 3485.380 641.630 3485.440 ;
        RECT 675.810 3485.380 676.130 3485.440 ;
        RECT 737.910 3485.580 738.230 3485.640 ;
        RECT 772.410 3485.580 772.730 3485.640 ;
        RECT 737.910 3485.440 772.730 3485.580 ;
        RECT 737.910 3485.380 738.230 3485.440 ;
        RECT 772.410 3485.380 772.730 3485.440 ;
        RECT 931.110 3485.580 931.430 3485.640 ;
        RECT 965.610 3485.580 965.930 3485.640 ;
        RECT 931.110 3485.440 965.930 3485.580 ;
        RECT 931.110 3485.380 931.430 3485.440 ;
        RECT 965.610 3485.380 965.930 3485.440 ;
        RECT 1027.710 3485.580 1028.030 3485.640 ;
        RECT 1062.210 3485.580 1062.530 3485.640 ;
        RECT 1027.710 3485.440 1062.530 3485.580 ;
        RECT 1027.710 3485.380 1028.030 3485.440 ;
        RECT 1062.210 3485.380 1062.530 3485.440 ;
        RECT 1124.310 3485.580 1124.630 3485.640 ;
        RECT 1158.810 3485.580 1159.130 3485.640 ;
        RECT 1124.310 3485.440 1159.130 3485.580 ;
        RECT 1124.310 3485.380 1124.630 3485.440 ;
        RECT 1158.810 3485.380 1159.130 3485.440 ;
        RECT 1220.910 3485.580 1221.230 3485.640 ;
        RECT 1255.410 3485.580 1255.730 3485.640 ;
        RECT 1220.910 3485.440 1255.730 3485.580 ;
        RECT 1220.910 3485.380 1221.230 3485.440 ;
        RECT 1255.410 3485.380 1255.730 3485.440 ;
        RECT 1317.510 3485.580 1317.830 3485.640 ;
        RECT 1352.010 3485.580 1352.330 3485.640 ;
        RECT 1317.510 3485.440 1352.330 3485.580 ;
        RECT 1317.510 3485.380 1317.830 3485.440 ;
        RECT 1352.010 3485.380 1352.330 3485.440 ;
        RECT 1414.110 3485.580 1414.430 3485.640 ;
        RECT 1448.610 3485.580 1448.930 3485.640 ;
        RECT 1414.110 3485.440 1448.930 3485.580 ;
        RECT 1414.110 3485.380 1414.430 3485.440 ;
        RECT 1448.610 3485.380 1448.930 3485.440 ;
        RECT 1510.710 3485.580 1511.030 3485.640 ;
        RECT 1545.210 3485.580 1545.530 3485.640 ;
        RECT 1510.710 3485.440 1545.530 3485.580 ;
        RECT 1510.710 3485.380 1511.030 3485.440 ;
        RECT 1545.210 3485.380 1545.530 3485.440 ;
        RECT 1607.310 3485.580 1607.630 3485.640 ;
        RECT 1641.810 3485.580 1642.130 3485.640 ;
        RECT 1607.310 3485.440 1642.130 3485.580 ;
        RECT 1607.310 3485.380 1607.630 3485.440 ;
        RECT 1641.810 3485.380 1642.130 3485.440 ;
      LAYER via ;
        RECT 2801.500 3486.400 2801.760 3486.660 ;
        RECT 2825.880 3486.400 2826.140 3486.660 ;
        RECT 834.540 3485.720 834.800 3485.980 ;
        RECT 862.140 3485.720 862.400 3485.980 ;
        RECT 2704.900 3485.720 2705.160 3485.980 ;
        RECT 2743.080 3485.720 2743.340 3485.980 ;
        RECT 351.540 3485.380 351.800 3485.640 ;
        RECT 386.040 3485.380 386.300 3485.640 ;
        RECT 448.140 3485.380 448.400 3485.640 ;
        RECT 482.640 3485.380 482.900 3485.640 ;
        RECT 544.740 3485.380 545.000 3485.640 ;
        RECT 579.240 3485.380 579.500 3485.640 ;
        RECT 641.340 3485.380 641.600 3485.640 ;
        RECT 675.840 3485.380 676.100 3485.640 ;
        RECT 737.940 3485.380 738.200 3485.640 ;
        RECT 772.440 3485.380 772.700 3485.640 ;
        RECT 931.140 3485.380 931.400 3485.640 ;
        RECT 965.640 3485.380 965.900 3485.640 ;
        RECT 1027.740 3485.380 1028.000 3485.640 ;
        RECT 1062.240 3485.380 1062.500 3485.640 ;
        RECT 1124.340 3485.380 1124.600 3485.640 ;
        RECT 1158.840 3485.380 1159.100 3485.640 ;
        RECT 1220.940 3485.380 1221.200 3485.640 ;
        RECT 1255.440 3485.380 1255.700 3485.640 ;
        RECT 1317.540 3485.380 1317.800 3485.640 ;
        RECT 1352.040 3485.380 1352.300 3485.640 ;
        RECT 1414.140 3485.380 1414.400 3485.640 ;
        RECT 1448.640 3485.380 1448.900 3485.640 ;
        RECT 1510.740 3485.380 1511.000 3485.640 ;
        RECT 1545.240 3485.380 1545.500 3485.640 ;
        RECT 1607.340 3485.380 1607.600 3485.640 ;
        RECT 1641.840 3485.380 1642.100 3485.640 ;
      LAYER met2 ;
        RECT 2766.530 3486.770 2766.810 3486.885 ;
        RECT 2767.450 3486.770 2767.730 3486.885 ;
        RECT 2766.530 3486.630 2767.730 3486.770 ;
        RECT 2766.530 3486.515 2766.810 3486.630 ;
        RECT 2767.450 3486.515 2767.730 3486.630 ;
        RECT 2801.490 3486.515 2801.770 3486.885 ;
        RECT 2801.500 3486.370 2801.760 3486.515 ;
        RECT 2825.880 3486.370 2826.140 3486.690 ;
        RECT 2825.940 3486.205 2826.080 3486.370 ;
        RECT 386.030 3485.835 386.310 3486.205 ;
        RECT 482.630 3485.835 482.910 3486.205 ;
        RECT 579.230 3485.835 579.510 3486.205 ;
        RECT 675.830 3485.835 676.110 3486.205 ;
        RECT 772.430 3485.835 772.710 3486.205 ;
        RECT 386.100 3485.670 386.240 3485.835 ;
        RECT 482.700 3485.670 482.840 3485.835 ;
        RECT 579.300 3485.670 579.440 3485.835 ;
        RECT 675.900 3485.670 676.040 3485.835 ;
        RECT 772.500 3485.670 772.640 3485.835 ;
        RECT 834.540 3485.690 834.800 3486.010 ;
        RECT 862.130 3485.835 862.410 3486.205 ;
        RECT 965.630 3485.835 965.910 3486.205 ;
        RECT 1062.230 3485.835 1062.510 3486.205 ;
        RECT 1158.830 3485.835 1159.110 3486.205 ;
        RECT 1255.430 3485.835 1255.710 3486.205 ;
        RECT 1352.030 3485.835 1352.310 3486.205 ;
        RECT 1448.630 3485.835 1448.910 3486.205 ;
        RECT 1545.230 3485.835 1545.510 3486.205 ;
        RECT 1641.830 3485.835 1642.110 3486.205 ;
        RECT 2704.890 3485.835 2705.170 3486.205 ;
        RECT 862.140 3485.690 862.400 3485.835 ;
        RECT 351.540 3485.525 351.800 3485.670 ;
        RECT 351.530 3485.155 351.810 3485.525 ;
        RECT 386.040 3485.350 386.300 3485.670 ;
        RECT 448.140 3485.525 448.400 3485.670 ;
        RECT 448.130 3485.155 448.410 3485.525 ;
        RECT 482.640 3485.350 482.900 3485.670 ;
        RECT 544.740 3485.525 545.000 3485.670 ;
        RECT 544.730 3485.155 545.010 3485.525 ;
        RECT 579.240 3485.350 579.500 3485.670 ;
        RECT 641.340 3485.525 641.600 3485.670 ;
        RECT 641.330 3485.155 641.610 3485.525 ;
        RECT 675.840 3485.350 676.100 3485.670 ;
        RECT 737.940 3485.525 738.200 3485.670 ;
        RECT 737.930 3485.155 738.210 3485.525 ;
        RECT 772.440 3485.350 772.700 3485.670 ;
        RECT 834.600 3485.525 834.740 3485.690 ;
        RECT 965.700 3485.670 965.840 3485.835 ;
        RECT 1062.300 3485.670 1062.440 3485.835 ;
        RECT 1158.900 3485.670 1159.040 3485.835 ;
        RECT 1255.500 3485.670 1255.640 3485.835 ;
        RECT 1352.100 3485.670 1352.240 3485.835 ;
        RECT 1448.700 3485.670 1448.840 3485.835 ;
        RECT 1545.300 3485.670 1545.440 3485.835 ;
        RECT 1641.900 3485.670 1642.040 3485.835 ;
        RECT 2704.900 3485.690 2705.160 3485.835 ;
        RECT 2743.080 3485.690 2743.340 3486.010 ;
        RECT 2825.870 3485.835 2826.150 3486.205 ;
        RECT 2863.590 3486.090 2863.870 3486.205 ;
        RECT 2863.200 3485.950 2863.870 3486.090 ;
        RECT 931.140 3485.525 931.400 3485.670 ;
        RECT 834.530 3485.155 834.810 3485.525 ;
        RECT 931.130 3485.155 931.410 3485.525 ;
        RECT 965.640 3485.350 965.900 3485.670 ;
        RECT 1027.740 3485.525 1028.000 3485.670 ;
        RECT 1027.730 3485.155 1028.010 3485.525 ;
        RECT 1062.240 3485.350 1062.500 3485.670 ;
        RECT 1124.340 3485.525 1124.600 3485.670 ;
        RECT 1124.330 3485.155 1124.610 3485.525 ;
        RECT 1158.840 3485.350 1159.100 3485.670 ;
        RECT 1220.940 3485.525 1221.200 3485.670 ;
        RECT 1220.930 3485.155 1221.210 3485.525 ;
        RECT 1255.440 3485.350 1255.700 3485.670 ;
        RECT 1317.540 3485.525 1317.800 3485.670 ;
        RECT 1317.530 3485.155 1317.810 3485.525 ;
        RECT 1352.040 3485.350 1352.300 3485.670 ;
        RECT 1414.140 3485.525 1414.400 3485.670 ;
        RECT 1414.130 3485.155 1414.410 3485.525 ;
        RECT 1448.640 3485.350 1448.900 3485.670 ;
        RECT 1510.740 3485.525 1511.000 3485.670 ;
        RECT 1510.730 3485.155 1511.010 3485.525 ;
        RECT 1545.240 3485.350 1545.500 3485.670 ;
        RECT 1607.340 3485.525 1607.600 3485.670 ;
        RECT 1607.330 3485.155 1607.610 3485.525 ;
        RECT 1641.840 3485.350 1642.100 3485.670 ;
        RECT 2743.140 3484.845 2743.280 3485.690 ;
        RECT 2863.200 3485.525 2863.340 3485.950 ;
        RECT 2863.590 3485.835 2863.870 3485.950 ;
        RECT 2863.130 3485.155 2863.410 3485.525 ;
        RECT 2743.070 3484.475 2743.350 3484.845 ;
      LAYER via2 ;
        RECT 2766.530 3486.560 2766.810 3486.840 ;
        RECT 2767.450 3486.560 2767.730 3486.840 ;
        RECT 2801.490 3486.560 2801.770 3486.840 ;
        RECT 386.030 3485.880 386.310 3486.160 ;
        RECT 482.630 3485.880 482.910 3486.160 ;
        RECT 579.230 3485.880 579.510 3486.160 ;
        RECT 675.830 3485.880 676.110 3486.160 ;
        RECT 772.430 3485.880 772.710 3486.160 ;
        RECT 862.130 3485.880 862.410 3486.160 ;
        RECT 965.630 3485.880 965.910 3486.160 ;
        RECT 1062.230 3485.880 1062.510 3486.160 ;
        RECT 1158.830 3485.880 1159.110 3486.160 ;
        RECT 1255.430 3485.880 1255.710 3486.160 ;
        RECT 1352.030 3485.880 1352.310 3486.160 ;
        RECT 1448.630 3485.880 1448.910 3486.160 ;
        RECT 1545.230 3485.880 1545.510 3486.160 ;
        RECT 1641.830 3485.880 1642.110 3486.160 ;
        RECT 2704.890 3485.880 2705.170 3486.160 ;
        RECT 351.530 3485.200 351.810 3485.480 ;
        RECT 448.130 3485.200 448.410 3485.480 ;
        RECT 544.730 3485.200 545.010 3485.480 ;
        RECT 641.330 3485.200 641.610 3485.480 ;
        RECT 737.930 3485.200 738.210 3485.480 ;
        RECT 2825.870 3485.880 2826.150 3486.160 ;
        RECT 834.530 3485.200 834.810 3485.480 ;
        RECT 931.130 3485.200 931.410 3485.480 ;
        RECT 1027.730 3485.200 1028.010 3485.480 ;
        RECT 1124.330 3485.200 1124.610 3485.480 ;
        RECT 1220.930 3485.200 1221.210 3485.480 ;
        RECT 1317.530 3485.200 1317.810 3485.480 ;
        RECT 1414.130 3485.200 1414.410 3485.480 ;
        RECT 1510.730 3485.200 1511.010 3485.480 ;
        RECT 1607.330 3485.200 1607.610 3485.480 ;
        RECT 2863.590 3485.880 2863.870 3486.160 ;
        RECT 2863.130 3485.200 2863.410 3485.480 ;
        RECT 2743.070 3484.520 2743.350 3484.800 ;
      LAYER met3 ;
        RECT 2917.600 3490.250 2924.800 3490.700 ;
        RECT 2916.710 3489.950 2924.800 3490.250 ;
        RECT 2752.910 3486.850 2753.290 3486.860 ;
        RECT 2766.505 3486.850 2766.835 3486.865 ;
        RECT 2752.910 3486.550 2766.835 3486.850 ;
        RECT 2752.910 3486.540 2753.290 3486.550 ;
        RECT 2766.505 3486.535 2766.835 3486.550 ;
        RECT 2767.425 3486.850 2767.755 3486.865 ;
        RECT 2801.465 3486.850 2801.795 3486.865 ;
        RECT 2767.425 3486.550 2801.795 3486.850 ;
        RECT 2767.425 3486.535 2767.755 3486.550 ;
        RECT 2801.465 3486.535 2801.795 3486.550 ;
        RECT 295.590 3486.170 295.970 3486.180 ;
        RECT 386.005 3486.170 386.335 3486.185 ;
        RECT 482.605 3486.170 482.935 3486.185 ;
        RECT 579.205 3486.170 579.535 3486.185 ;
        RECT 675.805 3486.170 676.135 3486.185 ;
        RECT 772.405 3486.170 772.735 3486.185 ;
        RECT 862.105 3486.170 862.435 3486.185 ;
        RECT 965.605 3486.170 965.935 3486.185 ;
        RECT 1062.205 3486.170 1062.535 3486.185 ;
        RECT 1158.805 3486.170 1159.135 3486.185 ;
        RECT 1255.405 3486.170 1255.735 3486.185 ;
        RECT 1352.005 3486.170 1352.335 3486.185 ;
        RECT 1448.605 3486.170 1448.935 3486.185 ;
        RECT 1545.205 3486.170 1545.535 3486.185 ;
        RECT 1641.805 3486.170 1642.135 3486.185 ;
        RECT 2704.865 3486.170 2705.195 3486.185 ;
        RECT 295.590 3485.870 304.210 3486.170 ;
        RECT 295.590 3485.860 295.970 3485.870 ;
        RECT 303.910 3485.490 304.210 3485.870 ;
        RECT 386.005 3485.870 400.810 3486.170 ;
        RECT 386.005 3485.855 386.335 3485.870 ;
        RECT 351.505 3485.490 351.835 3485.505 ;
        RECT 303.910 3485.190 351.835 3485.490 ;
        RECT 400.510 3485.490 400.810 3485.870 ;
        RECT 482.605 3485.870 497.410 3486.170 ;
        RECT 482.605 3485.855 482.935 3485.870 ;
        RECT 448.105 3485.490 448.435 3485.505 ;
        RECT 400.510 3485.190 448.435 3485.490 ;
        RECT 497.110 3485.490 497.410 3485.870 ;
        RECT 579.205 3485.870 594.010 3486.170 ;
        RECT 579.205 3485.855 579.535 3485.870 ;
        RECT 544.705 3485.490 545.035 3485.505 ;
        RECT 497.110 3485.190 545.035 3485.490 ;
        RECT 593.710 3485.490 594.010 3485.870 ;
        RECT 675.805 3485.870 690.610 3486.170 ;
        RECT 675.805 3485.855 676.135 3485.870 ;
        RECT 641.305 3485.490 641.635 3485.505 ;
        RECT 593.710 3485.190 641.635 3485.490 ;
        RECT 690.310 3485.490 690.610 3485.870 ;
        RECT 772.405 3485.870 787.210 3486.170 ;
        RECT 772.405 3485.855 772.735 3485.870 ;
        RECT 737.905 3485.490 738.235 3485.505 ;
        RECT 690.310 3485.190 738.235 3485.490 ;
        RECT 786.910 3485.490 787.210 3485.870 ;
        RECT 862.105 3485.870 883.810 3486.170 ;
        RECT 862.105 3485.855 862.435 3485.870 ;
        RECT 834.505 3485.490 834.835 3485.505 ;
        RECT 786.910 3485.190 834.835 3485.490 ;
        RECT 883.510 3485.490 883.810 3485.870 ;
        RECT 965.605 3485.870 980.410 3486.170 ;
        RECT 965.605 3485.855 965.935 3485.870 ;
        RECT 931.105 3485.490 931.435 3485.505 ;
        RECT 883.510 3485.190 931.435 3485.490 ;
        RECT 980.110 3485.490 980.410 3485.870 ;
        RECT 1062.205 3485.870 1077.010 3486.170 ;
        RECT 1062.205 3485.855 1062.535 3485.870 ;
        RECT 1027.705 3485.490 1028.035 3485.505 ;
        RECT 980.110 3485.190 1028.035 3485.490 ;
        RECT 1076.710 3485.490 1077.010 3485.870 ;
        RECT 1158.805 3485.870 1173.610 3486.170 ;
        RECT 1158.805 3485.855 1159.135 3485.870 ;
        RECT 1124.305 3485.490 1124.635 3485.505 ;
        RECT 1076.710 3485.190 1124.635 3485.490 ;
        RECT 1173.310 3485.490 1173.610 3485.870 ;
        RECT 1255.405 3485.870 1270.210 3486.170 ;
        RECT 1255.405 3485.855 1255.735 3485.870 ;
        RECT 1220.905 3485.490 1221.235 3485.505 ;
        RECT 1173.310 3485.190 1221.235 3485.490 ;
        RECT 1269.910 3485.490 1270.210 3485.870 ;
        RECT 1352.005 3485.870 1366.810 3486.170 ;
        RECT 1352.005 3485.855 1352.335 3485.870 ;
        RECT 1317.505 3485.490 1317.835 3485.505 ;
        RECT 1269.910 3485.190 1317.835 3485.490 ;
        RECT 1366.510 3485.490 1366.810 3485.870 ;
        RECT 1448.605 3485.870 1463.410 3486.170 ;
        RECT 1448.605 3485.855 1448.935 3485.870 ;
        RECT 1414.105 3485.490 1414.435 3485.505 ;
        RECT 1366.510 3485.190 1414.435 3485.490 ;
        RECT 1463.110 3485.490 1463.410 3485.870 ;
        RECT 1545.205 3485.870 1560.010 3486.170 ;
        RECT 1545.205 3485.855 1545.535 3485.870 ;
        RECT 1510.705 3485.490 1511.035 3485.505 ;
        RECT 1463.110 3485.190 1511.035 3485.490 ;
        RECT 1559.710 3485.490 1560.010 3485.870 ;
        RECT 1641.805 3485.870 1704.450 3486.170 ;
        RECT 1641.805 3485.855 1642.135 3485.870 ;
        RECT 1607.305 3485.490 1607.635 3485.505 ;
        RECT 1559.710 3485.190 1607.635 3485.490 ;
        RECT 1704.150 3485.490 1704.450 3485.870 ;
        RECT 1869.750 3485.870 1917.890 3486.170 ;
        RECT 1704.150 3485.190 1752.290 3485.490 ;
        RECT 351.505 3485.175 351.835 3485.190 ;
        RECT 448.105 3485.175 448.435 3485.190 ;
        RECT 544.705 3485.175 545.035 3485.190 ;
        RECT 641.305 3485.175 641.635 3485.190 ;
        RECT 737.905 3485.175 738.235 3485.190 ;
        RECT 834.505 3485.175 834.835 3485.190 ;
        RECT 931.105 3485.175 931.435 3485.190 ;
        RECT 1027.705 3485.175 1028.035 3485.190 ;
        RECT 1124.305 3485.175 1124.635 3485.190 ;
        RECT 1220.905 3485.175 1221.235 3485.190 ;
        RECT 1317.505 3485.175 1317.835 3485.190 ;
        RECT 1414.105 3485.175 1414.435 3485.190 ;
        RECT 1510.705 3485.175 1511.035 3485.190 ;
        RECT 1607.305 3485.175 1607.635 3485.190 ;
        RECT 1751.990 3484.810 1752.290 3485.190 ;
        RECT 1869.750 3484.810 1870.050 3485.870 ;
        RECT 1751.990 3484.510 1870.050 3484.810 ;
        RECT 1917.590 3484.810 1917.890 3485.870 ;
        RECT 1918.510 3485.870 1966.650 3486.170 ;
        RECT 1918.510 3484.810 1918.810 3485.870 ;
        RECT 1966.350 3485.490 1966.650 3485.870 ;
        RECT 2015.110 3485.870 2063.250 3486.170 ;
        RECT 1966.350 3485.190 2014.490 3485.490 ;
        RECT 1917.590 3484.510 1918.810 3484.810 ;
        RECT 2014.190 3484.810 2014.490 3485.190 ;
        RECT 2015.110 3484.810 2015.410 3485.870 ;
        RECT 2062.950 3485.490 2063.250 3485.870 ;
        RECT 2111.710 3485.870 2159.850 3486.170 ;
        RECT 2062.950 3485.190 2111.090 3485.490 ;
        RECT 2014.190 3484.510 2015.410 3484.810 ;
        RECT 2110.790 3484.810 2111.090 3485.190 ;
        RECT 2111.710 3484.810 2112.010 3485.870 ;
        RECT 2159.550 3485.490 2159.850 3485.870 ;
        RECT 2208.310 3485.870 2256.450 3486.170 ;
        RECT 2159.550 3485.190 2207.690 3485.490 ;
        RECT 2110.790 3484.510 2112.010 3484.810 ;
        RECT 2207.390 3484.810 2207.690 3485.190 ;
        RECT 2208.310 3484.810 2208.610 3485.870 ;
        RECT 2256.150 3485.490 2256.450 3485.870 ;
        RECT 2304.910 3485.870 2353.050 3486.170 ;
        RECT 2256.150 3485.190 2304.290 3485.490 ;
        RECT 2207.390 3484.510 2208.610 3484.810 ;
        RECT 2303.990 3484.810 2304.290 3485.190 ;
        RECT 2304.910 3484.810 2305.210 3485.870 ;
        RECT 2352.750 3485.490 2353.050 3485.870 ;
        RECT 2401.510 3485.870 2449.650 3486.170 ;
        RECT 2352.750 3485.190 2400.890 3485.490 ;
        RECT 2303.990 3484.510 2305.210 3484.810 ;
        RECT 2400.590 3484.810 2400.890 3485.190 ;
        RECT 2401.510 3484.810 2401.810 3485.870 ;
        RECT 2449.350 3485.490 2449.650 3485.870 ;
        RECT 2498.110 3485.870 2546.250 3486.170 ;
        RECT 2449.350 3485.190 2497.490 3485.490 ;
        RECT 2400.590 3484.510 2401.810 3484.810 ;
        RECT 2497.190 3484.810 2497.490 3485.190 ;
        RECT 2498.110 3484.810 2498.410 3485.870 ;
        RECT 2545.950 3485.490 2546.250 3485.870 ;
        RECT 2594.710 3485.870 2642.850 3486.170 ;
        RECT 2545.950 3485.190 2594.090 3485.490 ;
        RECT 2497.190 3484.510 2498.410 3484.810 ;
        RECT 2593.790 3484.810 2594.090 3485.190 ;
        RECT 2594.710 3484.810 2595.010 3485.870 ;
        RECT 2642.550 3485.490 2642.850 3485.870 ;
        RECT 2691.310 3485.870 2705.195 3486.170 ;
        RECT 2642.550 3485.190 2690.690 3485.490 ;
        RECT 2593.790 3484.510 2595.010 3484.810 ;
        RECT 2690.390 3484.810 2690.690 3485.190 ;
        RECT 2691.310 3484.810 2691.610 3485.870 ;
        RECT 2704.865 3485.855 2705.195 3485.870 ;
        RECT 2825.845 3486.170 2826.175 3486.185 ;
        RECT 2863.565 3486.170 2863.895 3486.185 ;
        RECT 2825.845 3485.870 2849.850 3486.170 ;
        RECT 2825.845 3485.855 2826.175 3485.870 ;
        RECT 2849.550 3485.490 2849.850 3485.870 ;
        RECT 2863.565 3485.870 2884.810 3486.170 ;
        RECT 2863.565 3485.855 2863.895 3485.870 ;
        RECT 2863.105 3485.490 2863.435 3485.505 ;
        RECT 2849.550 3485.190 2863.435 3485.490 ;
        RECT 2884.510 3485.490 2884.810 3485.870 ;
        RECT 2916.710 3485.490 2917.010 3489.950 ;
        RECT 2917.600 3489.500 2924.800 3489.950 ;
        RECT 2884.510 3485.190 2917.010 3485.490 ;
        RECT 2863.105 3485.175 2863.435 3485.190 ;
        RECT 2690.390 3484.510 2691.610 3484.810 ;
        RECT 2743.045 3484.810 2743.375 3484.825 ;
        RECT 2752.910 3484.810 2753.290 3484.820 ;
        RECT 2743.045 3484.510 2753.290 3484.810 ;
        RECT 2743.045 3484.495 2743.375 3484.510 ;
        RECT 2752.910 3484.500 2753.290 3484.510 ;
        RECT 295.590 1957.530 295.970 1957.540 ;
        RECT 300.000 1957.530 304.000 1957.600 ;
        RECT 295.590 1957.230 304.000 1957.530 ;
        RECT 295.590 1957.220 295.970 1957.230 ;
        RECT 300.000 1957.000 304.000 1957.230 ;
      LAYER via3 ;
        RECT 2752.940 3486.540 2753.260 3486.860 ;
        RECT 295.620 3485.860 295.940 3486.180 ;
        RECT 2752.940 3484.500 2753.260 3484.820 ;
        RECT 295.620 1957.220 295.940 1957.540 ;
      LAYER met4 ;
        RECT 2752.935 3486.535 2753.265 3486.865 ;
        RECT 295.615 3485.855 295.945 3486.185 ;
        RECT 295.630 1957.545 295.930 3485.855 ;
        RECT 2752.950 3484.825 2753.250 3486.535 ;
        RECT 2752.935 3484.495 2753.265 3484.825 ;
        RECT 295.615 1957.215 295.945 1957.545 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 296.310 3501.900 296.630 3501.960 ;
        RECT 2635.870 3501.900 2636.190 3501.960 ;
        RECT 296.310 3501.760 2636.190 3501.900 ;
        RECT 296.310 3501.700 296.630 3501.760 ;
        RECT 2635.870 3501.700 2636.190 3501.760 ;
      LAYER via ;
        RECT 296.340 3501.700 296.600 3501.960 ;
        RECT 2635.900 3501.700 2636.160 3501.960 ;
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
        RECT 2635.960 3501.990 2636.100 3517.600 ;
        RECT 296.340 3501.670 296.600 3501.990 ;
        RECT 2635.900 3501.670 2636.160 3501.990 ;
        RECT 296.400 1989.525 296.540 3501.670 ;
        RECT 296.330 1989.155 296.610 1989.525 ;
      LAYER via2 ;
        RECT 296.330 1989.200 296.610 1989.480 ;
      LAYER met3 ;
        RECT 296.305 1989.490 296.635 1989.505 ;
        RECT 300.000 1989.490 304.000 1989.560 ;
        RECT 296.305 1989.190 304.000 1989.490 ;
        RECT 296.305 1989.175 296.635 1989.190 ;
        RECT 300.000 1988.960 304.000 1989.190 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 291.710 3253.700 292.030 3253.760 ;
        RECT 2311.570 3253.700 2311.890 3253.760 ;
        RECT 291.710 3253.560 2311.890 3253.700 ;
        RECT 291.710 3253.500 292.030 3253.560 ;
        RECT 2311.570 3253.500 2311.890 3253.560 ;
      LAYER via ;
        RECT 291.740 3253.500 292.000 3253.760 ;
        RECT 2311.600 3253.500 2311.860 3253.760 ;
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
        RECT 2311.660 3253.790 2311.800 3517.600 ;
        RECT 291.740 3253.470 292.000 3253.790 ;
        RECT 2311.600 3253.470 2311.860 3253.790 ;
        RECT 291.800 2020.805 291.940 3253.470 ;
        RECT 291.730 2020.435 292.010 2020.805 ;
      LAYER via2 ;
        RECT 291.730 2020.480 292.010 2020.760 ;
      LAYER met3 ;
        RECT 291.705 2020.770 292.035 2020.785 ;
        RECT 300.000 2020.770 304.000 2020.840 ;
        RECT 291.705 2020.470 304.000 2020.770 ;
        RECT 291.705 2020.455 292.035 2020.470 ;
        RECT 300.000 2020.240 304.000 2020.470 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 295.850 3502.920 296.170 3502.980 ;
        RECT 1987.270 3502.920 1987.590 3502.980 ;
        RECT 295.850 3502.780 1987.590 3502.920 ;
        RECT 295.850 3502.720 296.170 3502.780 ;
        RECT 1987.270 3502.720 1987.590 3502.780 ;
      LAYER via ;
        RECT 295.880 3502.720 296.140 3502.980 ;
        RECT 1987.300 3502.720 1987.560 3502.980 ;
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
        RECT 1987.360 3503.010 1987.500 3517.600 ;
        RECT 295.880 3502.690 296.140 3503.010 ;
        RECT 1987.300 3502.690 1987.560 3503.010 ;
        RECT 295.940 2052.765 296.080 3502.690 ;
        RECT 295.870 2052.395 296.150 2052.765 ;
      LAYER via2 ;
        RECT 295.870 2052.440 296.150 2052.720 ;
      LAYER met3 ;
        RECT 295.845 2052.730 296.175 2052.745 ;
        RECT 300.000 2052.730 304.000 2052.800 ;
        RECT 295.845 2052.430 304.000 2052.730 ;
        RECT 295.845 2052.415 296.175 2052.430 ;
        RECT 300.000 2052.200 304.000 2052.430 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 295.390 3503.600 295.710 3503.660 ;
        RECT 1662.510 3503.600 1662.830 3503.660 ;
        RECT 295.390 3503.460 1662.830 3503.600 ;
        RECT 295.390 3503.400 295.710 3503.460 ;
        RECT 1662.510 3503.400 1662.830 3503.460 ;
      LAYER via ;
        RECT 295.420 3503.400 295.680 3503.660 ;
        RECT 1662.540 3503.400 1662.800 3503.660 ;
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
        RECT 1662.600 3503.690 1662.740 3517.600 ;
        RECT 295.420 3503.370 295.680 3503.690 ;
        RECT 1662.540 3503.370 1662.800 3503.690 ;
        RECT 295.480 2084.045 295.620 3503.370 ;
        RECT 295.410 2083.675 295.690 2084.045 ;
      LAYER via2 ;
        RECT 295.410 2083.720 295.690 2084.000 ;
      LAYER met3 ;
        RECT 295.385 2084.010 295.715 2084.025 ;
        RECT 300.000 2084.010 304.000 2084.080 ;
        RECT 295.385 2083.710 304.000 2084.010 ;
        RECT 295.385 2083.695 295.715 2083.710 ;
        RECT 300.000 2083.480 304.000 2083.710 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 294.930 3504.280 295.250 3504.340 ;
        RECT 1338.210 3504.280 1338.530 3504.340 ;
        RECT 294.930 3504.140 1338.530 3504.280 ;
        RECT 294.930 3504.080 295.250 3504.140 ;
        RECT 1338.210 3504.080 1338.530 3504.140 ;
      LAYER via ;
        RECT 294.960 3504.080 295.220 3504.340 ;
        RECT 1338.240 3504.080 1338.500 3504.340 ;
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
        RECT 1338.300 3504.370 1338.440 3517.600 ;
        RECT 294.960 3504.050 295.220 3504.370 ;
        RECT 1338.240 3504.050 1338.500 3504.370 ;
        RECT 295.020 2115.325 295.160 3504.050 ;
        RECT 294.950 2114.955 295.230 2115.325 ;
      LAYER via2 ;
        RECT 294.950 2115.000 295.230 2115.280 ;
      LAYER met3 ;
        RECT 294.925 2115.290 295.255 2115.305 ;
        RECT 300.000 2115.290 304.000 2115.360 ;
        RECT 294.925 2114.990 304.000 2115.290 ;
        RECT 294.925 2114.975 295.255 2114.990 ;
        RECT 300.000 2114.760 304.000 2114.990 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 282.970 441.560 283.290 441.620 ;
        RECT 2900.830 441.560 2901.150 441.620 ;
        RECT 282.970 441.420 2901.150 441.560 ;
        RECT 282.970 441.360 283.290 441.420 ;
        RECT 2900.830 441.360 2901.150 441.420 ;
      LAYER via ;
        RECT 283.000 441.360 283.260 441.620 ;
        RECT 2900.860 441.360 2901.120 441.620 ;
      LAYER met2 ;
        RECT 282.990 1546.475 283.270 1546.845 ;
        RECT 283.060 441.650 283.200 1546.475 ;
        RECT 283.000 441.330 283.260 441.650 ;
        RECT 2900.860 441.330 2901.120 441.650 ;
        RECT 2900.920 439.805 2901.060 441.330 ;
        RECT 2900.850 439.435 2901.130 439.805 ;
      LAYER via2 ;
        RECT 282.990 1546.520 283.270 1546.800 ;
        RECT 2900.850 439.480 2901.130 439.760 ;
      LAYER met3 ;
        RECT 282.965 1546.810 283.295 1546.825 ;
        RECT 300.000 1546.810 304.000 1546.880 ;
        RECT 282.965 1546.510 304.000 1546.810 ;
        RECT 282.965 1546.495 283.295 1546.510 ;
        RECT 300.000 1546.280 304.000 1546.510 ;
        RECT 2900.825 439.770 2901.155 439.785 ;
        RECT 2917.600 439.770 2924.800 440.220 ;
        RECT 2900.825 439.470 2924.800 439.770 ;
        RECT 2900.825 439.455 2901.155 439.470 ;
        RECT 2917.600 439.020 2924.800 439.470 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 294.010 3504.960 294.330 3505.020 ;
        RECT 1013.910 3504.960 1014.230 3505.020 ;
        RECT 294.010 3504.820 1014.230 3504.960 ;
        RECT 294.010 3504.760 294.330 3504.820 ;
        RECT 1013.910 3504.760 1014.230 3504.820 ;
      LAYER via ;
        RECT 294.040 3504.760 294.300 3505.020 ;
        RECT 1013.940 3504.760 1014.200 3505.020 ;
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
        RECT 1014.000 3505.050 1014.140 3517.600 ;
        RECT 294.040 3504.730 294.300 3505.050 ;
        RECT 1013.940 3504.730 1014.200 3505.050 ;
        RECT 294.100 2147.285 294.240 3504.730 ;
        RECT 294.030 2146.915 294.310 2147.285 ;
      LAYER via2 ;
        RECT 294.030 2146.960 294.310 2147.240 ;
      LAYER met3 ;
        RECT 294.005 2147.250 294.335 2147.265 ;
        RECT 300.000 2147.250 304.000 2147.320 ;
        RECT 294.005 2146.950 304.000 2147.250 ;
        RECT 294.005 2146.935 294.335 2146.950 ;
        RECT 300.000 2146.720 304.000 2146.950 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 292.630 3501.220 292.950 3501.280 ;
        RECT 683.170 3501.220 683.490 3501.280 ;
        RECT 292.630 3501.080 683.490 3501.220 ;
        RECT 292.630 3501.020 292.950 3501.080 ;
        RECT 683.170 3501.020 683.490 3501.080 ;
        RECT 683.170 3500.540 683.490 3500.600 ;
        RECT 689.150 3500.540 689.470 3500.600 ;
        RECT 683.170 3500.400 689.470 3500.540 ;
        RECT 683.170 3500.340 683.490 3500.400 ;
        RECT 689.150 3500.340 689.470 3500.400 ;
      LAYER via ;
        RECT 292.660 3501.020 292.920 3501.280 ;
        RECT 683.200 3501.020 683.460 3501.280 ;
        RECT 683.200 3500.340 683.460 3500.600 ;
        RECT 689.180 3500.340 689.440 3500.600 ;
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
        RECT 292.660 3500.990 292.920 3501.310 ;
        RECT 683.200 3500.990 683.460 3501.310 ;
        RECT 292.720 2178.565 292.860 3500.990 ;
        RECT 683.260 3500.630 683.400 3500.990 ;
        RECT 689.240 3500.630 689.380 3517.600 ;
        RECT 683.200 3500.310 683.460 3500.630 ;
        RECT 689.180 3500.310 689.440 3500.630 ;
        RECT 292.650 2178.195 292.930 2178.565 ;
      LAYER via2 ;
        RECT 292.650 2178.240 292.930 2178.520 ;
      LAYER met3 ;
        RECT 292.625 2178.530 292.955 2178.545 ;
        RECT 300.000 2178.530 304.000 2178.600 ;
        RECT 292.625 2178.230 304.000 2178.530 ;
        RECT 292.625 2178.215 292.955 2178.230 ;
        RECT 300.000 2178.000 304.000 2178.230 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 292.170 3500.200 292.490 3500.260 ;
        RECT 364.850 3500.200 365.170 3500.260 ;
        RECT 292.170 3500.060 365.170 3500.200 ;
        RECT 292.170 3500.000 292.490 3500.060 ;
        RECT 364.850 3500.000 365.170 3500.060 ;
      LAYER via ;
        RECT 292.200 3500.000 292.460 3500.260 ;
        RECT 364.880 3500.000 365.140 3500.260 ;
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
        RECT 364.940 3500.290 365.080 3517.600 ;
        RECT 292.200 3499.970 292.460 3500.290 ;
        RECT 364.880 3499.970 365.140 3500.290 ;
        RECT 292.260 2210.525 292.400 3499.970 ;
        RECT 292.190 2210.155 292.470 2210.525 ;
      LAYER via2 ;
        RECT 292.190 2210.200 292.470 2210.480 ;
      LAYER met3 ;
        RECT 292.165 2210.490 292.495 2210.505 ;
        RECT 300.000 2210.490 304.000 2210.560 ;
        RECT 292.165 2210.190 304.000 2210.490 ;
        RECT 292.165 2210.175 292.495 2210.190 ;
        RECT 300.000 2209.960 304.000 2210.190 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 40.550 3498.500 40.870 3498.560 ;
        RECT 51.590 3498.500 51.910 3498.560 ;
        RECT 40.550 3498.360 51.910 3498.500 ;
        RECT 40.550 3498.300 40.870 3498.360 ;
        RECT 51.590 3498.300 51.910 3498.360 ;
        RECT 51.590 2242.540 51.910 2242.600 ;
        RECT 287.570 2242.540 287.890 2242.600 ;
        RECT 51.590 2242.400 287.890 2242.540 ;
        RECT 51.590 2242.340 51.910 2242.400 ;
        RECT 287.570 2242.340 287.890 2242.400 ;
      LAYER via ;
        RECT 40.580 3498.300 40.840 3498.560 ;
        RECT 51.620 3498.300 51.880 3498.560 ;
        RECT 51.620 2242.340 51.880 2242.600 ;
        RECT 287.600 2242.340 287.860 2242.600 ;
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
        RECT 40.640 3498.590 40.780 3517.600 ;
        RECT 40.580 3498.270 40.840 3498.590 ;
        RECT 51.620 3498.270 51.880 3498.590 ;
        RECT 51.680 2242.630 51.820 3498.270 ;
        RECT 51.620 2242.310 51.880 2242.630 ;
        RECT 287.600 2242.310 287.860 2242.630 ;
        RECT 287.660 2241.805 287.800 2242.310 ;
        RECT 287.590 2241.435 287.870 2241.805 ;
      LAYER via2 ;
        RECT 287.590 2241.480 287.870 2241.760 ;
      LAYER met3 ;
        RECT 287.565 2241.770 287.895 2241.785 ;
        RECT 300.000 2241.770 304.000 2241.840 ;
        RECT 287.565 2241.470 304.000 2241.770 ;
        RECT 287.565 2241.455 287.895 2241.470 ;
        RECT 300.000 2241.240 304.000 2241.470 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.250 3263.900 15.570 3263.960 ;
        RECT 65.390 3263.900 65.710 3263.960 ;
        RECT 15.250 3263.760 65.710 3263.900 ;
        RECT 15.250 3263.700 15.570 3263.760 ;
        RECT 65.390 3263.700 65.710 3263.760 ;
        RECT 65.390 2276.880 65.710 2276.940 ;
        RECT 282.970 2276.880 283.290 2276.940 ;
        RECT 65.390 2276.740 283.290 2276.880 ;
        RECT 65.390 2276.680 65.710 2276.740 ;
        RECT 282.970 2276.680 283.290 2276.740 ;
      LAYER via ;
        RECT 15.280 3263.700 15.540 3263.960 ;
        RECT 65.420 3263.700 65.680 3263.960 ;
        RECT 65.420 2276.680 65.680 2276.940 ;
        RECT 283.000 2276.680 283.260 2276.940 ;
      LAYER met2 ;
        RECT 15.270 3267.555 15.550 3267.925 ;
        RECT 15.340 3263.990 15.480 3267.555 ;
        RECT 15.280 3263.670 15.540 3263.990 ;
        RECT 65.420 3263.670 65.680 3263.990 ;
        RECT 65.480 2276.970 65.620 3263.670 ;
        RECT 65.420 2276.650 65.680 2276.970 ;
        RECT 283.000 2276.650 283.260 2276.970 ;
        RECT 283.060 2273.765 283.200 2276.650 ;
        RECT 282.990 2273.395 283.270 2273.765 ;
      LAYER via2 ;
        RECT 15.270 3267.600 15.550 3267.880 ;
        RECT 282.990 2273.440 283.270 2273.720 ;
      LAYER met3 ;
        RECT -4.800 3267.890 2.400 3268.340 ;
        RECT 15.245 3267.890 15.575 3267.905 ;
        RECT -4.800 3267.590 15.575 3267.890 ;
        RECT -4.800 3267.140 2.400 3267.590 ;
        RECT 15.245 3267.575 15.575 3267.590 ;
        RECT 282.965 2273.730 283.295 2273.745 ;
        RECT 300.000 2273.730 304.000 2273.800 ;
        RECT 282.965 2273.430 304.000 2273.730 ;
        RECT 282.965 2273.415 283.295 2273.430 ;
        RECT 300.000 2273.200 304.000 2273.430 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.170 2974.220 16.490 2974.280 ;
        RECT 72.290 2974.220 72.610 2974.280 ;
        RECT 16.170 2974.080 72.610 2974.220 ;
        RECT 16.170 2974.020 16.490 2974.080 ;
        RECT 72.290 2974.020 72.610 2974.080 ;
        RECT 72.290 2311.560 72.610 2311.620 ;
        RECT 282.510 2311.560 282.830 2311.620 ;
        RECT 72.290 2311.420 282.830 2311.560 ;
        RECT 72.290 2311.360 72.610 2311.420 ;
        RECT 282.510 2311.360 282.830 2311.420 ;
      LAYER via ;
        RECT 16.200 2974.020 16.460 2974.280 ;
        RECT 72.320 2974.020 72.580 2974.280 ;
        RECT 72.320 2311.360 72.580 2311.620 ;
        RECT 282.540 2311.360 282.800 2311.620 ;
      LAYER met2 ;
        RECT 16.190 2979.915 16.470 2980.285 ;
        RECT 16.260 2974.310 16.400 2979.915 ;
        RECT 16.200 2973.990 16.460 2974.310 ;
        RECT 72.320 2973.990 72.580 2974.310 ;
        RECT 72.380 2311.650 72.520 2973.990 ;
        RECT 72.320 2311.330 72.580 2311.650 ;
        RECT 282.540 2311.330 282.800 2311.650 ;
        RECT 282.600 2307.765 282.740 2311.330 ;
        RECT 282.530 2307.395 282.810 2307.765 ;
      LAYER via2 ;
        RECT 16.190 2979.960 16.470 2980.240 ;
        RECT 282.530 2307.440 282.810 2307.720 ;
      LAYER met3 ;
        RECT -4.800 2980.250 2.400 2980.700 ;
        RECT 16.165 2980.250 16.495 2980.265 ;
        RECT -4.800 2979.950 16.495 2980.250 ;
        RECT -4.800 2979.500 2.400 2979.950 ;
        RECT 16.165 2979.935 16.495 2979.950 ;
        RECT 282.505 2307.730 282.835 2307.745 ;
        RECT 282.505 2307.430 300.530 2307.730 ;
        RECT 282.505 2307.415 282.835 2307.430 ;
        RECT 300.230 2305.080 300.530 2307.430 ;
        RECT 300.000 2304.480 304.000 2305.080 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 14.790 2692.020 15.110 2692.080 ;
        RECT 26.750 2692.020 27.070 2692.080 ;
        RECT 14.790 2691.880 27.070 2692.020 ;
        RECT 14.790 2691.820 15.110 2691.880 ;
        RECT 26.750 2691.820 27.070 2691.880 ;
        RECT 26.750 2339.100 27.070 2339.160 ;
        RECT 282.510 2339.100 282.830 2339.160 ;
        RECT 26.750 2338.960 282.830 2339.100 ;
        RECT 26.750 2338.900 27.070 2338.960 ;
        RECT 282.510 2338.900 282.830 2338.960 ;
      LAYER via ;
        RECT 14.820 2691.820 15.080 2692.080 ;
        RECT 26.780 2691.820 27.040 2692.080 ;
        RECT 26.780 2338.900 27.040 2339.160 ;
        RECT 282.540 2338.900 282.800 2339.160 ;
      LAYER met2 ;
        RECT 14.810 2692.955 15.090 2693.325 ;
        RECT 14.880 2692.110 15.020 2692.955 ;
        RECT 14.820 2691.790 15.080 2692.110 ;
        RECT 26.780 2691.790 27.040 2692.110 ;
        RECT 26.840 2339.190 26.980 2691.790 ;
        RECT 26.780 2338.870 27.040 2339.190 ;
        RECT 282.540 2339.045 282.800 2339.190 ;
        RECT 282.530 2338.675 282.810 2339.045 ;
      LAYER via2 ;
        RECT 14.810 2693.000 15.090 2693.280 ;
        RECT 282.530 2338.720 282.810 2339.000 ;
      LAYER met3 ;
        RECT -4.800 2693.290 2.400 2693.740 ;
        RECT 14.785 2693.290 15.115 2693.305 ;
        RECT -4.800 2692.990 15.115 2693.290 ;
        RECT -4.800 2692.540 2.400 2692.990 ;
        RECT 14.785 2692.975 15.115 2692.990 ;
        RECT 282.505 2339.010 282.835 2339.025 ;
        RECT 282.505 2338.710 300.530 2339.010 ;
        RECT 282.505 2338.695 282.835 2338.710 ;
        RECT 300.230 2337.040 300.530 2338.710 ;
        RECT 300.000 2336.440 304.000 2337.040 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.170 2403.360 16.490 2403.420 ;
        RECT 27.670 2403.360 27.990 2403.420 ;
        RECT 16.170 2403.220 27.990 2403.360 ;
        RECT 16.170 2403.160 16.490 2403.220 ;
        RECT 27.670 2403.160 27.990 2403.220 ;
        RECT 27.670 2373.440 27.990 2373.500 ;
        RECT 282.970 2373.440 283.290 2373.500 ;
        RECT 27.670 2373.300 283.290 2373.440 ;
        RECT 27.670 2373.240 27.990 2373.300 ;
        RECT 282.970 2373.240 283.290 2373.300 ;
      LAYER via ;
        RECT 16.200 2403.160 16.460 2403.420 ;
        RECT 27.700 2403.160 27.960 2403.420 ;
        RECT 27.700 2373.240 27.960 2373.500 ;
        RECT 283.000 2373.240 283.260 2373.500 ;
      LAYER met2 ;
        RECT 16.190 2405.315 16.470 2405.685 ;
        RECT 16.260 2403.450 16.400 2405.315 ;
        RECT 16.200 2403.130 16.460 2403.450 ;
        RECT 27.700 2403.130 27.960 2403.450 ;
        RECT 27.760 2373.530 27.900 2403.130 ;
        RECT 27.700 2373.210 27.960 2373.530 ;
        RECT 283.000 2373.210 283.260 2373.530 ;
        RECT 283.060 2368.285 283.200 2373.210 ;
        RECT 282.990 2367.915 283.270 2368.285 ;
      LAYER via2 ;
        RECT 16.190 2405.360 16.470 2405.640 ;
        RECT 282.990 2367.960 283.270 2368.240 ;
      LAYER met3 ;
        RECT -4.800 2405.650 2.400 2406.100 ;
        RECT 16.165 2405.650 16.495 2405.665 ;
        RECT -4.800 2405.350 16.495 2405.650 ;
        RECT -4.800 2404.900 2.400 2405.350 ;
        RECT 16.165 2405.335 16.495 2405.350 ;
        RECT 282.965 2368.250 283.295 2368.265 ;
        RECT 300.000 2368.250 304.000 2368.320 ;
        RECT 282.965 2367.950 304.000 2368.250 ;
        RECT 282.965 2367.935 283.295 2367.950 ;
        RECT 300.000 2367.720 304.000 2367.950 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 19.850 2394.520 20.170 2394.580 ;
        RECT 282.970 2394.520 283.290 2394.580 ;
        RECT 19.850 2394.380 283.290 2394.520 ;
        RECT 19.850 2394.320 20.170 2394.380 ;
        RECT 282.970 2394.320 283.290 2394.380 ;
      LAYER via ;
        RECT 19.880 2394.320 20.140 2394.580 ;
        RECT 283.000 2394.320 283.260 2394.580 ;
      LAYER met2 ;
        RECT 282.990 2399.875 283.270 2400.245 ;
        RECT 283.060 2394.610 283.200 2399.875 ;
        RECT 19.880 2394.290 20.140 2394.610 ;
        RECT 283.000 2394.290 283.260 2394.610 ;
        RECT 19.940 2118.725 20.080 2394.290 ;
        RECT 19.870 2118.355 20.150 2118.725 ;
      LAYER via2 ;
        RECT 282.990 2399.920 283.270 2400.200 ;
        RECT 19.870 2118.400 20.150 2118.680 ;
      LAYER met3 ;
        RECT 282.965 2400.210 283.295 2400.225 ;
        RECT 300.000 2400.210 304.000 2400.280 ;
        RECT 282.965 2399.910 304.000 2400.210 ;
        RECT 282.965 2399.895 283.295 2399.910 ;
        RECT 300.000 2399.680 304.000 2399.910 ;
        RECT -4.800 2118.690 2.400 2119.140 ;
        RECT 19.845 2118.690 20.175 2118.705 ;
        RECT -4.800 2118.390 20.175 2118.690 ;
        RECT -4.800 2117.940 2.400 2118.390 ;
        RECT 19.845 2118.375 20.175 2118.390 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 79.190 2429.200 79.510 2429.260 ;
        RECT 282.970 2429.200 283.290 2429.260 ;
        RECT 79.190 2429.060 283.290 2429.200 ;
        RECT 79.190 2429.000 79.510 2429.060 ;
        RECT 282.970 2429.000 283.290 2429.060 ;
        RECT 14.790 1835.220 15.110 1835.280 ;
        RECT 79.190 1835.220 79.510 1835.280 ;
        RECT 14.790 1835.080 79.510 1835.220 ;
        RECT 14.790 1835.020 15.110 1835.080 ;
        RECT 79.190 1835.020 79.510 1835.080 ;
      LAYER via ;
        RECT 79.220 2429.000 79.480 2429.260 ;
        RECT 283.000 2429.000 283.260 2429.260 ;
        RECT 14.820 1835.020 15.080 1835.280 ;
        RECT 79.220 1835.020 79.480 1835.280 ;
      LAYER met2 ;
        RECT 282.990 2431.155 283.270 2431.525 ;
        RECT 283.060 2429.290 283.200 2431.155 ;
        RECT 79.220 2428.970 79.480 2429.290 ;
        RECT 283.000 2428.970 283.260 2429.290 ;
        RECT 79.280 1835.310 79.420 2428.970 ;
        RECT 14.820 1834.990 15.080 1835.310 ;
        RECT 79.220 1834.990 79.480 1835.310 ;
        RECT 14.880 1831.085 15.020 1834.990 ;
        RECT 14.810 1830.715 15.090 1831.085 ;
      LAYER via2 ;
        RECT 282.990 2431.200 283.270 2431.480 ;
        RECT 14.810 1830.760 15.090 1831.040 ;
      LAYER met3 ;
        RECT 282.965 2431.490 283.295 2431.505 ;
        RECT 300.000 2431.490 304.000 2431.560 ;
        RECT 282.965 2431.190 304.000 2431.490 ;
        RECT 282.965 2431.175 283.295 2431.190 ;
        RECT 300.000 2430.960 304.000 2431.190 ;
        RECT -4.800 1831.050 2.400 1831.500 ;
        RECT 14.785 1831.050 15.115 1831.065 ;
        RECT -4.800 1830.750 15.115 1831.050 ;
        RECT -4.800 1830.300 2.400 1830.750 ;
        RECT 14.785 1830.735 15.115 1830.750 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 288.490 676.160 288.810 676.220 ;
        RECT 2900.830 676.160 2901.150 676.220 ;
        RECT 288.490 676.020 2901.150 676.160 ;
        RECT 288.490 675.960 288.810 676.020 ;
        RECT 2900.830 675.960 2901.150 676.020 ;
      LAYER via ;
        RECT 288.520 675.960 288.780 676.220 ;
        RECT 2900.860 675.960 2901.120 676.220 ;
      LAYER met2 ;
        RECT 288.510 1578.435 288.790 1578.805 ;
        RECT 288.580 676.250 288.720 1578.435 ;
        RECT 288.520 675.930 288.780 676.250 ;
        RECT 2900.860 675.930 2901.120 676.250 ;
        RECT 2900.920 674.405 2901.060 675.930 ;
        RECT 2900.850 674.035 2901.130 674.405 ;
      LAYER via2 ;
        RECT 288.510 1578.480 288.790 1578.760 ;
        RECT 2900.850 674.080 2901.130 674.360 ;
      LAYER met3 ;
        RECT 288.485 1578.770 288.815 1578.785 ;
        RECT 300.000 1578.770 304.000 1578.840 ;
        RECT 288.485 1578.470 304.000 1578.770 ;
        RECT 288.485 1578.455 288.815 1578.470 ;
        RECT 300.000 1578.240 304.000 1578.470 ;
        RECT 2900.825 674.370 2901.155 674.385 ;
        RECT 2917.600 674.370 2924.800 674.820 ;
        RECT 2900.825 674.070 2924.800 674.370 ;
        RECT 2900.825 674.055 2901.155 674.070 ;
        RECT 2917.600 673.620 2924.800 674.070 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 86.550 2456.740 86.870 2456.800 ;
        RECT 286.190 2456.740 286.510 2456.800 ;
        RECT 86.550 2456.600 286.510 2456.740 ;
        RECT 86.550 2456.540 86.870 2456.600 ;
        RECT 286.190 2456.540 286.510 2456.600 ;
        RECT 16.630 1545.540 16.950 1545.600 ;
        RECT 86.550 1545.540 86.870 1545.600 ;
        RECT 16.630 1545.400 86.870 1545.540 ;
        RECT 16.630 1545.340 16.950 1545.400 ;
        RECT 86.550 1545.340 86.870 1545.400 ;
      LAYER via ;
        RECT 86.580 2456.540 86.840 2456.800 ;
        RECT 286.220 2456.540 286.480 2456.800 ;
        RECT 16.660 1545.340 16.920 1545.600 ;
        RECT 86.580 1545.340 86.840 1545.600 ;
      LAYER met2 ;
        RECT 286.210 2462.435 286.490 2462.805 ;
        RECT 286.280 2456.830 286.420 2462.435 ;
        RECT 86.580 2456.510 86.840 2456.830 ;
        RECT 286.220 2456.510 286.480 2456.830 ;
        RECT 86.640 1545.630 86.780 2456.510 ;
        RECT 16.660 1545.310 16.920 1545.630 ;
        RECT 86.580 1545.310 86.840 1545.630 ;
        RECT 16.720 1544.125 16.860 1545.310 ;
        RECT 16.650 1543.755 16.930 1544.125 ;
      LAYER via2 ;
        RECT 286.210 2462.480 286.490 2462.760 ;
        RECT 16.650 1543.800 16.930 1544.080 ;
      LAYER met3 ;
        RECT 286.185 2462.770 286.515 2462.785 ;
        RECT 300.000 2462.770 304.000 2462.840 ;
        RECT 286.185 2462.470 304.000 2462.770 ;
        RECT 286.185 2462.455 286.515 2462.470 ;
        RECT 300.000 2462.240 304.000 2462.470 ;
        RECT -4.800 1544.090 2.400 1544.540 ;
        RECT 16.625 1544.090 16.955 1544.105 ;
        RECT -4.800 1543.790 16.955 1544.090 ;
        RECT -4.800 1543.340 2.400 1543.790 ;
        RECT 16.625 1543.775 16.955 1543.790 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 100.350 2491.080 100.670 2491.140 ;
        RECT 286.190 2491.080 286.510 2491.140 ;
        RECT 100.350 2490.940 286.510 2491.080 ;
        RECT 100.350 2490.880 100.670 2490.940 ;
        RECT 286.190 2490.880 286.510 2490.940 ;
        RECT 15.710 1331.680 16.030 1331.740 ;
        RECT 100.350 1331.680 100.670 1331.740 ;
        RECT 15.710 1331.540 100.670 1331.680 ;
        RECT 15.710 1331.480 16.030 1331.540 ;
        RECT 100.350 1331.480 100.670 1331.540 ;
      LAYER via ;
        RECT 100.380 2490.880 100.640 2491.140 ;
        RECT 286.220 2490.880 286.480 2491.140 ;
        RECT 15.740 1331.480 16.000 1331.740 ;
        RECT 100.380 1331.480 100.640 1331.740 ;
      LAYER met2 ;
        RECT 286.210 2494.395 286.490 2494.765 ;
        RECT 286.280 2491.170 286.420 2494.395 ;
        RECT 100.380 2490.850 100.640 2491.170 ;
        RECT 286.220 2490.850 286.480 2491.170 ;
        RECT 100.440 1331.770 100.580 2490.850 ;
        RECT 15.740 1331.450 16.000 1331.770 ;
        RECT 100.380 1331.450 100.640 1331.770 ;
        RECT 15.800 1328.565 15.940 1331.450 ;
        RECT 15.730 1328.195 16.010 1328.565 ;
      LAYER via2 ;
        RECT 286.210 2494.440 286.490 2494.720 ;
        RECT 15.730 1328.240 16.010 1328.520 ;
      LAYER met3 ;
        RECT 286.185 2494.730 286.515 2494.745 ;
        RECT 300.000 2494.730 304.000 2494.800 ;
        RECT 286.185 2494.430 304.000 2494.730 ;
        RECT 286.185 2494.415 286.515 2494.430 ;
        RECT 300.000 2494.200 304.000 2494.430 ;
        RECT -4.800 1328.530 2.400 1328.980 ;
        RECT 15.705 1328.530 16.035 1328.545 ;
        RECT -4.800 1328.230 16.035 1328.530 ;
        RECT -4.800 1327.780 2.400 1328.230 ;
        RECT 15.705 1328.215 16.035 1328.230 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 141.290 2525.760 141.610 2525.820 ;
        RECT 286.190 2525.760 286.510 2525.820 ;
        RECT 141.290 2525.620 286.510 2525.760 ;
        RECT 141.290 2525.560 141.610 2525.620 ;
        RECT 286.190 2525.560 286.510 2525.620 ;
        RECT 16.630 1117.820 16.950 1117.880 ;
        RECT 141.290 1117.820 141.610 1117.880 ;
        RECT 16.630 1117.680 141.610 1117.820 ;
        RECT 16.630 1117.620 16.950 1117.680 ;
        RECT 141.290 1117.620 141.610 1117.680 ;
      LAYER via ;
        RECT 141.320 2525.560 141.580 2525.820 ;
        RECT 286.220 2525.560 286.480 2525.820 ;
        RECT 16.660 1117.620 16.920 1117.880 ;
        RECT 141.320 1117.620 141.580 1117.880 ;
      LAYER met2 ;
        RECT 141.320 2525.530 141.580 2525.850 ;
        RECT 286.210 2525.675 286.490 2526.045 ;
        RECT 286.220 2525.530 286.480 2525.675 ;
        RECT 141.380 1117.910 141.520 2525.530 ;
        RECT 16.660 1117.590 16.920 1117.910 ;
        RECT 141.320 1117.590 141.580 1117.910 ;
        RECT 16.720 1113.005 16.860 1117.590 ;
        RECT 16.650 1112.635 16.930 1113.005 ;
      LAYER via2 ;
        RECT 286.210 2525.720 286.490 2526.000 ;
        RECT 16.650 1112.680 16.930 1112.960 ;
      LAYER met3 ;
        RECT 286.185 2526.010 286.515 2526.025 ;
        RECT 300.000 2526.010 304.000 2526.080 ;
        RECT 286.185 2525.710 304.000 2526.010 ;
        RECT 286.185 2525.695 286.515 2525.710 ;
        RECT 300.000 2525.480 304.000 2525.710 ;
        RECT -4.800 1112.970 2.400 1113.420 ;
        RECT 16.625 1112.970 16.955 1112.985 ;
        RECT -4.800 1112.670 16.955 1112.970 ;
        RECT -4.800 1112.220 2.400 1112.670 ;
        RECT 16.625 1112.655 16.955 1112.670 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 168.890 2553.300 169.210 2553.360 ;
        RECT 286.190 2553.300 286.510 2553.360 ;
        RECT 168.890 2553.160 286.510 2553.300 ;
        RECT 168.890 2553.100 169.210 2553.160 ;
        RECT 286.190 2553.100 286.510 2553.160 ;
        RECT 16.170 903.960 16.490 904.020 ;
        RECT 168.890 903.960 169.210 904.020 ;
        RECT 16.170 903.820 169.210 903.960 ;
        RECT 16.170 903.760 16.490 903.820 ;
        RECT 168.890 903.760 169.210 903.820 ;
      LAYER via ;
        RECT 168.920 2553.100 169.180 2553.360 ;
        RECT 286.220 2553.100 286.480 2553.360 ;
        RECT 16.200 903.760 16.460 904.020 ;
        RECT 168.920 903.760 169.180 904.020 ;
      LAYER met2 ;
        RECT 286.210 2557.635 286.490 2558.005 ;
        RECT 286.280 2553.390 286.420 2557.635 ;
        RECT 168.920 2553.070 169.180 2553.390 ;
        RECT 286.220 2553.070 286.480 2553.390 ;
        RECT 168.980 904.050 169.120 2553.070 ;
        RECT 16.200 903.730 16.460 904.050 ;
        RECT 168.920 903.730 169.180 904.050 ;
        RECT 16.260 897.445 16.400 903.730 ;
        RECT 16.190 897.075 16.470 897.445 ;
      LAYER via2 ;
        RECT 286.210 2557.680 286.490 2557.960 ;
        RECT 16.190 897.120 16.470 897.400 ;
      LAYER met3 ;
        RECT 286.185 2557.970 286.515 2557.985 ;
        RECT 300.000 2557.970 304.000 2558.040 ;
        RECT 286.185 2557.670 304.000 2557.970 ;
        RECT 286.185 2557.655 286.515 2557.670 ;
        RECT 300.000 2557.440 304.000 2557.670 ;
        RECT -4.800 897.410 2.400 897.860 ;
        RECT 16.165 897.410 16.495 897.425 ;
        RECT -4.800 897.110 16.495 897.410 ;
        RECT -4.800 896.660 2.400 897.110 ;
        RECT 16.165 897.095 16.495 897.110 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 175.790 2587.640 176.110 2587.700 ;
        RECT 286.190 2587.640 286.510 2587.700 ;
        RECT 175.790 2587.500 286.510 2587.640 ;
        RECT 175.790 2587.440 176.110 2587.500 ;
        RECT 286.190 2587.440 286.510 2587.500 ;
        RECT 16.170 682.960 16.490 683.020 ;
        RECT 175.790 682.960 176.110 683.020 ;
        RECT 16.170 682.820 176.110 682.960 ;
        RECT 16.170 682.760 16.490 682.820 ;
        RECT 175.790 682.760 176.110 682.820 ;
      LAYER via ;
        RECT 175.820 2587.440 176.080 2587.700 ;
        RECT 286.220 2587.440 286.480 2587.700 ;
        RECT 16.200 682.760 16.460 683.020 ;
        RECT 175.820 682.760 176.080 683.020 ;
      LAYER met2 ;
        RECT 286.210 2588.915 286.490 2589.285 ;
        RECT 286.280 2587.730 286.420 2588.915 ;
        RECT 175.820 2587.410 176.080 2587.730 ;
        RECT 286.220 2587.410 286.480 2587.730 ;
        RECT 175.880 683.050 176.020 2587.410 ;
        RECT 16.200 682.730 16.460 683.050 ;
        RECT 175.820 682.730 176.080 683.050 ;
        RECT 16.260 681.885 16.400 682.730 ;
        RECT 16.190 681.515 16.470 681.885 ;
      LAYER via2 ;
        RECT 286.210 2588.960 286.490 2589.240 ;
        RECT 16.190 681.560 16.470 681.840 ;
      LAYER met3 ;
        RECT 286.185 2589.250 286.515 2589.265 ;
        RECT 300.000 2589.250 304.000 2589.320 ;
        RECT 286.185 2588.950 304.000 2589.250 ;
        RECT 286.185 2588.935 286.515 2588.950 ;
        RECT 300.000 2588.720 304.000 2588.950 ;
        RECT -4.800 681.850 2.400 682.300 ;
        RECT 16.165 681.850 16.495 681.865 ;
        RECT -4.800 681.550 16.495 681.850 ;
        RECT -4.800 681.100 2.400 681.550 ;
        RECT 16.165 681.535 16.495 681.550 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 217.190 2615.180 217.510 2615.240 ;
        RECT 286.190 2615.180 286.510 2615.240 ;
        RECT 217.190 2615.040 286.510 2615.180 ;
        RECT 217.190 2614.980 217.510 2615.040 ;
        RECT 286.190 2614.980 286.510 2615.040 ;
        RECT 17.090 469.100 17.410 469.160 ;
        RECT 217.190 469.100 217.510 469.160 ;
        RECT 17.090 468.960 217.510 469.100 ;
        RECT 17.090 468.900 17.410 468.960 ;
        RECT 217.190 468.900 217.510 468.960 ;
      LAYER via ;
        RECT 217.220 2614.980 217.480 2615.240 ;
        RECT 286.220 2614.980 286.480 2615.240 ;
        RECT 17.120 468.900 17.380 469.160 ;
        RECT 217.220 468.900 217.480 469.160 ;
      LAYER met2 ;
        RECT 286.210 2620.875 286.490 2621.245 ;
        RECT 286.280 2615.270 286.420 2620.875 ;
        RECT 217.220 2614.950 217.480 2615.270 ;
        RECT 286.220 2614.950 286.480 2615.270 ;
        RECT 217.280 469.190 217.420 2614.950 ;
        RECT 17.120 468.870 17.380 469.190 ;
        RECT 217.220 468.870 217.480 469.190 ;
        RECT 17.180 466.325 17.320 468.870 ;
        RECT 17.110 465.955 17.390 466.325 ;
      LAYER via2 ;
        RECT 286.210 2620.920 286.490 2621.200 ;
        RECT 17.110 466.000 17.390 466.280 ;
      LAYER met3 ;
        RECT 286.185 2621.210 286.515 2621.225 ;
        RECT 300.000 2621.210 304.000 2621.280 ;
        RECT 286.185 2620.910 304.000 2621.210 ;
        RECT 286.185 2620.895 286.515 2620.910 ;
        RECT 300.000 2620.680 304.000 2620.910 ;
        RECT -4.800 466.290 2.400 466.740 ;
        RECT 17.085 466.290 17.415 466.305 ;
        RECT -4.800 465.990 17.415 466.290 ;
        RECT -4.800 465.540 2.400 465.990 ;
        RECT 17.085 465.975 17.415 465.990 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 230.990 2649.860 231.310 2649.920 ;
        RECT 286.190 2649.860 286.510 2649.920 ;
        RECT 230.990 2649.720 286.510 2649.860 ;
        RECT 230.990 2649.660 231.310 2649.720 ;
        RECT 286.190 2649.660 286.510 2649.720 ;
        RECT 17.090 255.240 17.410 255.300 ;
        RECT 230.990 255.240 231.310 255.300 ;
        RECT 17.090 255.100 231.310 255.240 ;
        RECT 17.090 255.040 17.410 255.100 ;
        RECT 230.990 255.040 231.310 255.100 ;
      LAYER via ;
        RECT 231.020 2649.660 231.280 2649.920 ;
        RECT 286.220 2649.660 286.480 2649.920 ;
        RECT 17.120 255.040 17.380 255.300 ;
        RECT 231.020 255.040 231.280 255.300 ;
      LAYER met2 ;
        RECT 286.210 2652.155 286.490 2652.525 ;
        RECT 286.280 2649.950 286.420 2652.155 ;
        RECT 231.020 2649.630 231.280 2649.950 ;
        RECT 286.220 2649.630 286.480 2649.950 ;
        RECT 231.080 255.330 231.220 2649.630 ;
        RECT 17.120 255.010 17.380 255.330 ;
        RECT 231.020 255.010 231.280 255.330 ;
        RECT 17.180 250.765 17.320 255.010 ;
        RECT 17.110 250.395 17.390 250.765 ;
      LAYER via2 ;
        RECT 286.210 2652.200 286.490 2652.480 ;
        RECT 17.110 250.440 17.390 250.720 ;
      LAYER met3 ;
        RECT 286.185 2652.490 286.515 2652.505 ;
        RECT 300.000 2652.490 304.000 2652.560 ;
        RECT 286.185 2652.190 304.000 2652.490 ;
        RECT 286.185 2652.175 286.515 2652.190 ;
        RECT 300.000 2651.960 304.000 2652.190 ;
        RECT -4.800 250.730 2.400 251.180 ;
        RECT 17.085 250.730 17.415 250.745 ;
        RECT -4.800 250.430 17.415 250.730 ;
        RECT -4.800 249.980 2.400 250.430 ;
        RECT 17.085 250.415 17.415 250.430 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 244.790 2684.200 245.110 2684.260 ;
        RECT 286.190 2684.200 286.510 2684.260 ;
        RECT 244.790 2684.060 286.510 2684.200 ;
        RECT 244.790 2684.000 245.110 2684.060 ;
        RECT 286.190 2684.000 286.510 2684.060 ;
        RECT 17.090 41.380 17.410 41.440 ;
        RECT 244.790 41.380 245.110 41.440 ;
        RECT 17.090 41.240 245.110 41.380 ;
        RECT 17.090 41.180 17.410 41.240 ;
        RECT 244.790 41.180 245.110 41.240 ;
      LAYER via ;
        RECT 244.820 2684.000 245.080 2684.260 ;
        RECT 286.220 2684.000 286.480 2684.260 ;
        RECT 17.120 41.180 17.380 41.440 ;
        RECT 244.820 41.180 245.080 41.440 ;
      LAYER met2 ;
        RECT 244.820 2683.970 245.080 2684.290 ;
        RECT 286.210 2684.115 286.490 2684.485 ;
        RECT 286.220 2683.970 286.480 2684.115 ;
        RECT 244.880 41.470 245.020 2683.970 ;
        RECT 17.120 41.150 17.380 41.470 ;
        RECT 244.820 41.150 245.080 41.470 ;
        RECT 17.180 35.885 17.320 41.150 ;
        RECT 17.110 35.515 17.390 35.885 ;
      LAYER via2 ;
        RECT 286.210 2684.160 286.490 2684.440 ;
        RECT 17.110 35.560 17.390 35.840 ;
      LAYER met3 ;
        RECT 286.185 2684.450 286.515 2684.465 ;
        RECT 300.000 2684.450 304.000 2684.520 ;
        RECT 286.185 2684.150 304.000 2684.450 ;
        RECT 286.185 2684.135 286.515 2684.150 ;
        RECT 300.000 2683.920 304.000 2684.150 ;
        RECT -4.800 35.850 2.400 36.300 ;
        RECT 17.085 35.850 17.415 35.865 ;
        RECT -4.800 35.550 17.415 35.850 ;
        RECT -4.800 35.100 2.400 35.550 ;
        RECT 17.085 35.535 17.415 35.550 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 288.950 1589.400 289.270 1589.460 ;
        RECT 287.200 1589.260 289.270 1589.400 ;
        RECT 287.200 1586.340 287.340 1589.260 ;
        RECT 288.950 1589.200 289.270 1589.260 ;
        RECT 287.570 1586.340 287.890 1586.400 ;
        RECT 287.200 1586.200 287.890 1586.340 ;
        RECT 287.570 1586.140 287.890 1586.200 ;
        RECT 282.970 1579.880 283.290 1579.940 ;
        RECT 287.570 1579.880 287.890 1579.940 ;
        RECT 282.970 1579.740 287.890 1579.880 ;
        RECT 282.970 1579.680 283.290 1579.740 ;
        RECT 287.570 1579.680 287.890 1579.740 ;
        RECT 282.510 1531.940 282.830 1532.000 ;
        RECT 287.570 1531.940 287.890 1532.000 ;
        RECT 282.510 1531.800 287.890 1531.940 ;
        RECT 282.510 1531.740 282.830 1531.800 ;
        RECT 287.570 1531.740 287.890 1531.800 ;
        RECT 287.570 1483.320 287.890 1483.380 ;
        RECT 289.410 1483.320 289.730 1483.380 ;
        RECT 287.570 1483.180 289.730 1483.320 ;
        RECT 287.570 1483.120 287.890 1483.180 ;
        RECT 289.410 1483.120 289.730 1483.180 ;
        RECT 287.570 1435.380 287.890 1435.440 ;
        RECT 289.410 1435.380 289.730 1435.440 ;
        RECT 287.570 1435.240 289.730 1435.380 ;
        RECT 287.570 1435.180 287.890 1435.240 ;
        RECT 289.410 1435.180 289.730 1435.240 ;
        RECT 286.190 1386.760 286.510 1386.820 ;
        RECT 287.570 1386.760 287.890 1386.820 ;
        RECT 286.190 1386.620 287.890 1386.760 ;
        RECT 286.190 1386.560 286.510 1386.620 ;
        RECT 287.570 1386.560 287.890 1386.620 ;
        RECT 286.190 1318.080 286.510 1318.140 ;
        RECT 287.570 1318.080 287.890 1318.140 ;
        RECT 286.190 1317.940 287.890 1318.080 ;
        RECT 286.190 1317.880 286.510 1317.940 ;
        RECT 287.570 1317.880 287.890 1317.940 ;
        RECT 287.570 910.760 287.890 910.820 ;
        RECT 2900.830 910.760 2901.150 910.820 ;
        RECT 287.570 910.620 2901.150 910.760 ;
        RECT 287.570 910.560 287.890 910.620 ;
        RECT 2900.830 910.560 2901.150 910.620 ;
      LAYER via ;
        RECT 288.980 1589.200 289.240 1589.460 ;
        RECT 287.600 1586.140 287.860 1586.400 ;
        RECT 283.000 1579.680 283.260 1579.940 ;
        RECT 287.600 1579.680 287.860 1579.940 ;
        RECT 282.540 1531.740 282.800 1532.000 ;
        RECT 287.600 1531.740 287.860 1532.000 ;
        RECT 287.600 1483.120 287.860 1483.380 ;
        RECT 289.440 1483.120 289.700 1483.380 ;
        RECT 287.600 1435.180 287.860 1435.440 ;
        RECT 289.440 1435.180 289.700 1435.440 ;
        RECT 286.220 1386.560 286.480 1386.820 ;
        RECT 287.600 1386.560 287.860 1386.820 ;
        RECT 286.220 1317.880 286.480 1318.140 ;
        RECT 287.600 1317.880 287.860 1318.140 ;
        RECT 287.600 910.560 287.860 910.820 ;
        RECT 2900.860 910.560 2901.120 910.820 ;
      LAYER met2 ;
        RECT 288.970 1609.715 289.250 1610.085 ;
        RECT 289.040 1589.490 289.180 1609.715 ;
        RECT 288.980 1589.170 289.240 1589.490 ;
        RECT 287.600 1586.110 287.860 1586.430 ;
        RECT 287.660 1579.970 287.800 1586.110 ;
        RECT 283.000 1579.650 283.260 1579.970 ;
        RECT 287.600 1579.650 287.860 1579.970 ;
        RECT 283.060 1547.410 283.200 1579.650 ;
        RECT 282.600 1547.270 283.200 1547.410 ;
        RECT 282.600 1532.030 282.740 1547.270 ;
        RECT 282.540 1531.710 282.800 1532.030 ;
        RECT 287.600 1531.710 287.860 1532.030 ;
        RECT 287.660 1483.410 287.800 1531.710 ;
        RECT 287.600 1483.090 287.860 1483.410 ;
        RECT 289.440 1483.090 289.700 1483.410 ;
        RECT 289.500 1435.470 289.640 1483.090 ;
        RECT 287.600 1435.150 287.860 1435.470 ;
        RECT 289.440 1435.150 289.700 1435.470 ;
        RECT 287.660 1386.850 287.800 1435.150 ;
        RECT 286.220 1386.530 286.480 1386.850 ;
        RECT 287.600 1386.530 287.860 1386.850 ;
        RECT 286.280 1318.170 286.420 1386.530 ;
        RECT 286.220 1317.850 286.480 1318.170 ;
        RECT 287.600 1317.850 287.860 1318.170 ;
        RECT 287.660 910.850 287.800 1317.850 ;
        RECT 287.600 910.530 287.860 910.850 ;
        RECT 2900.860 910.530 2901.120 910.850 ;
        RECT 2900.920 909.685 2901.060 910.530 ;
        RECT 2900.850 909.315 2901.130 909.685 ;
      LAYER via2 ;
        RECT 288.970 1609.760 289.250 1610.040 ;
        RECT 2900.850 909.360 2901.130 909.640 ;
      LAYER met3 ;
        RECT 288.945 1610.050 289.275 1610.065 ;
        RECT 300.000 1610.050 304.000 1610.120 ;
        RECT 288.945 1609.750 304.000 1610.050 ;
        RECT 288.945 1609.735 289.275 1609.750 ;
        RECT 300.000 1609.520 304.000 1609.750 ;
        RECT 2900.825 909.650 2901.155 909.665 ;
        RECT 2917.600 909.650 2924.800 910.100 ;
        RECT 2900.825 909.350 2924.800 909.650 ;
        RECT 2900.825 909.335 2901.155 909.350 ;
        RECT 2917.600 908.900 2924.800 909.350 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 285.730 1145.360 286.050 1145.420 ;
        RECT 2900.830 1145.360 2901.150 1145.420 ;
        RECT 285.730 1145.220 2901.150 1145.360 ;
        RECT 285.730 1145.160 286.050 1145.220 ;
        RECT 2900.830 1145.160 2901.150 1145.220 ;
      LAYER via ;
        RECT 285.760 1145.160 286.020 1145.420 ;
        RECT 2900.860 1145.160 2901.120 1145.420 ;
      LAYER met2 ;
        RECT 285.750 1641.675 286.030 1642.045 ;
        RECT 285.820 1145.450 285.960 1641.675 ;
        RECT 285.760 1145.130 286.020 1145.450 ;
        RECT 2900.860 1145.130 2901.120 1145.450 ;
        RECT 2900.920 1144.285 2901.060 1145.130 ;
        RECT 2900.850 1143.915 2901.130 1144.285 ;
      LAYER via2 ;
        RECT 285.750 1641.720 286.030 1642.000 ;
        RECT 2900.850 1143.960 2901.130 1144.240 ;
      LAYER met3 ;
        RECT 285.725 1642.010 286.055 1642.025 ;
        RECT 300.000 1642.010 304.000 1642.080 ;
        RECT 285.725 1641.710 304.000 1642.010 ;
        RECT 285.725 1641.695 286.055 1641.710 ;
        RECT 300.000 1641.480 304.000 1641.710 ;
        RECT 2900.825 1144.250 2901.155 1144.265 ;
        RECT 2917.600 1144.250 2924.800 1144.700 ;
        RECT 2900.825 1143.950 2924.800 1144.250 ;
        RECT 2900.825 1143.935 2901.155 1143.950 ;
        RECT 2917.600 1143.500 2924.800 1143.950 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 284.350 1379.960 284.670 1380.020 ;
        RECT 2900.830 1379.960 2901.150 1380.020 ;
        RECT 284.350 1379.820 2901.150 1379.960 ;
        RECT 284.350 1379.760 284.670 1379.820 ;
        RECT 2900.830 1379.760 2901.150 1379.820 ;
      LAYER via ;
        RECT 284.380 1379.760 284.640 1380.020 ;
        RECT 2900.860 1379.760 2901.120 1380.020 ;
      LAYER met2 ;
        RECT 284.370 1672.955 284.650 1673.325 ;
        RECT 284.440 1380.050 284.580 1672.955 ;
        RECT 284.380 1379.730 284.640 1380.050 ;
        RECT 2900.860 1379.730 2901.120 1380.050 ;
        RECT 2900.920 1378.885 2901.060 1379.730 ;
        RECT 2900.850 1378.515 2901.130 1378.885 ;
      LAYER via2 ;
        RECT 284.370 1673.000 284.650 1673.280 ;
        RECT 2900.850 1378.560 2901.130 1378.840 ;
      LAYER met3 ;
        RECT 284.345 1673.290 284.675 1673.305 ;
        RECT 300.000 1673.290 304.000 1673.360 ;
        RECT 284.345 1672.990 304.000 1673.290 ;
        RECT 284.345 1672.975 284.675 1672.990 ;
        RECT 300.000 1672.760 304.000 1672.990 ;
        RECT 2900.825 1378.850 2901.155 1378.865 ;
        RECT 2917.600 1378.850 2924.800 1379.300 ;
        RECT 2900.825 1378.550 2924.800 1378.850 ;
        RECT 2900.825 1378.535 2901.155 1378.550 ;
        RECT 2917.600 1378.100 2924.800 1378.550 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 289.410 1504.060 289.730 1504.120 ;
        RECT 2901.290 1504.060 2901.610 1504.120 ;
        RECT 289.410 1503.920 2901.610 1504.060 ;
        RECT 289.410 1503.860 289.730 1503.920 ;
        RECT 2901.290 1503.860 2901.610 1503.920 ;
      LAYER via ;
        RECT 289.440 1503.860 289.700 1504.120 ;
        RECT 2901.320 1503.860 2901.580 1504.120 ;
      LAYER met2 ;
        RECT 289.430 1704.915 289.710 1705.285 ;
        RECT 289.500 1504.150 289.640 1704.915 ;
        RECT 2901.310 1613.115 2901.590 1613.485 ;
        RECT 2901.380 1504.150 2901.520 1613.115 ;
        RECT 289.440 1503.830 289.700 1504.150 ;
        RECT 2901.320 1503.830 2901.580 1504.150 ;
      LAYER via2 ;
        RECT 289.430 1704.960 289.710 1705.240 ;
        RECT 2901.310 1613.160 2901.590 1613.440 ;
      LAYER met3 ;
        RECT 289.405 1705.250 289.735 1705.265 ;
        RECT 300.000 1705.250 304.000 1705.320 ;
        RECT 289.405 1704.950 304.000 1705.250 ;
        RECT 289.405 1704.935 289.735 1704.950 ;
        RECT 300.000 1704.720 304.000 1704.950 ;
        RECT 2901.285 1613.450 2901.615 1613.465 ;
        RECT 2917.600 1613.450 2924.800 1613.900 ;
        RECT 2901.285 1613.150 2924.800 1613.450 ;
        RECT 2901.285 1613.135 2901.615 1613.150 ;
        RECT 2917.600 1612.700 2924.800 1613.150 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2887.950 1835.560 2888.270 1835.620 ;
        RECT 2897.610 1835.560 2897.930 1835.620 ;
        RECT 2887.950 1835.420 2897.930 1835.560 ;
        RECT 2887.950 1835.360 2888.270 1835.420 ;
        RECT 2897.610 1835.360 2897.930 1835.420 ;
        RECT 2870.470 1725.400 2870.790 1725.460 ;
        RECT 2887.950 1725.400 2888.270 1725.460 ;
        RECT 2870.470 1725.260 2888.270 1725.400 ;
        RECT 2870.470 1725.200 2870.790 1725.260 ;
        RECT 2887.950 1725.200 2888.270 1725.260 ;
        RECT 2857.130 1704.660 2857.450 1704.720 ;
        RECT 2870.470 1704.660 2870.790 1704.720 ;
        RECT 2857.130 1704.520 2870.790 1704.660 ;
        RECT 2857.130 1704.460 2857.450 1704.520 ;
        RECT 2870.470 1704.460 2870.790 1704.520 ;
        RECT 2854.830 1681.880 2855.150 1681.940 ;
        RECT 2857.130 1681.880 2857.450 1681.940 ;
        RECT 2854.830 1681.740 2857.450 1681.880 ;
        RECT 2854.830 1681.680 2855.150 1681.740 ;
        RECT 2857.130 1681.680 2857.450 1681.740 ;
        RECT 2839.190 1656.720 2839.510 1656.780 ;
        RECT 2854.830 1656.720 2855.150 1656.780 ;
        RECT 2839.190 1656.580 2855.150 1656.720 ;
        RECT 2839.190 1656.520 2839.510 1656.580 ;
        RECT 2854.830 1656.520 2855.150 1656.580 ;
        RECT 2825.390 1650.600 2825.710 1650.660 ;
        RECT 2839.190 1650.600 2839.510 1650.660 ;
        RECT 2825.390 1650.460 2839.510 1650.600 ;
        RECT 2825.390 1650.400 2825.710 1650.460 ;
        RECT 2839.190 1650.400 2839.510 1650.460 ;
        RECT 288.950 1614.900 289.270 1614.960 ;
        RECT 295.390 1614.900 295.710 1614.960 ;
        RECT 288.950 1614.760 295.710 1614.900 ;
        RECT 288.950 1614.700 289.270 1614.760 ;
        RECT 295.390 1614.700 295.710 1614.760 ;
        RECT 295.390 1573.420 295.710 1573.480 ;
        RECT 299.990 1573.420 300.310 1573.480 ;
        RECT 295.390 1573.280 300.310 1573.420 ;
        RECT 295.390 1573.220 295.710 1573.280 ;
        RECT 299.990 1573.220 300.310 1573.280 ;
        RECT 2804.690 1573.420 2805.010 1573.480 ;
        RECT 2825.390 1573.420 2825.710 1573.480 ;
        RECT 2804.690 1573.280 2825.710 1573.420 ;
        RECT 2804.690 1573.220 2805.010 1573.280 ;
        RECT 2825.390 1573.220 2825.710 1573.280 ;
        RECT 2795.490 1511.880 2795.810 1511.940 ;
        RECT 2804.690 1511.880 2805.010 1511.940 ;
        RECT 2795.490 1511.740 2805.010 1511.880 ;
        RECT 2795.490 1511.680 2795.810 1511.740 ;
        RECT 2804.690 1511.680 2805.010 1511.740 ;
        RECT 299.990 1503.040 300.310 1503.100 ;
        RECT 2795.490 1503.040 2795.810 1503.100 ;
        RECT 299.990 1502.900 2795.810 1503.040 ;
        RECT 299.990 1502.840 300.310 1502.900 ;
        RECT 2795.490 1502.840 2795.810 1502.900 ;
      LAYER via ;
        RECT 2887.980 1835.360 2888.240 1835.620 ;
        RECT 2897.640 1835.360 2897.900 1835.620 ;
        RECT 2870.500 1725.200 2870.760 1725.460 ;
        RECT 2887.980 1725.200 2888.240 1725.460 ;
        RECT 2857.160 1704.460 2857.420 1704.720 ;
        RECT 2870.500 1704.460 2870.760 1704.720 ;
        RECT 2854.860 1681.680 2855.120 1681.940 ;
        RECT 2857.160 1681.680 2857.420 1681.940 ;
        RECT 2839.220 1656.520 2839.480 1656.780 ;
        RECT 2854.860 1656.520 2855.120 1656.780 ;
        RECT 2825.420 1650.400 2825.680 1650.660 ;
        RECT 2839.220 1650.400 2839.480 1650.660 ;
        RECT 288.980 1614.700 289.240 1614.960 ;
        RECT 295.420 1614.700 295.680 1614.960 ;
        RECT 295.420 1573.220 295.680 1573.480 ;
        RECT 300.020 1573.220 300.280 1573.480 ;
        RECT 2804.720 1573.220 2804.980 1573.480 ;
        RECT 2825.420 1573.220 2825.680 1573.480 ;
        RECT 2795.520 1511.680 2795.780 1511.940 ;
        RECT 2804.720 1511.680 2804.980 1511.940 ;
        RECT 300.020 1502.840 300.280 1503.100 ;
        RECT 2795.520 1502.840 2795.780 1503.100 ;
      LAYER met2 ;
        RECT 2897.630 1847.715 2897.910 1848.085 ;
        RECT 2897.700 1835.650 2897.840 1847.715 ;
        RECT 2887.980 1835.330 2888.240 1835.650 ;
        RECT 2897.640 1835.330 2897.900 1835.650 ;
        RECT 288.970 1736.195 289.250 1736.565 ;
        RECT 289.040 1614.990 289.180 1736.195 ;
        RECT 2888.040 1725.490 2888.180 1835.330 ;
        RECT 2870.500 1725.170 2870.760 1725.490 ;
        RECT 2887.980 1725.170 2888.240 1725.490 ;
        RECT 2870.560 1704.750 2870.700 1725.170 ;
        RECT 2857.160 1704.430 2857.420 1704.750 ;
        RECT 2870.500 1704.430 2870.760 1704.750 ;
        RECT 2857.220 1681.970 2857.360 1704.430 ;
        RECT 2854.860 1681.650 2855.120 1681.970 ;
        RECT 2857.160 1681.650 2857.420 1681.970 ;
        RECT 2854.920 1656.810 2855.060 1681.650 ;
        RECT 2839.220 1656.490 2839.480 1656.810 ;
        RECT 2854.860 1656.490 2855.120 1656.810 ;
        RECT 2839.280 1650.690 2839.420 1656.490 ;
        RECT 2825.420 1650.370 2825.680 1650.690 ;
        RECT 2839.220 1650.370 2839.480 1650.690 ;
        RECT 288.980 1614.670 289.240 1614.990 ;
        RECT 295.420 1614.670 295.680 1614.990 ;
        RECT 295.480 1573.510 295.620 1614.670 ;
        RECT 2825.480 1573.510 2825.620 1650.370 ;
        RECT 295.420 1573.190 295.680 1573.510 ;
        RECT 300.020 1573.190 300.280 1573.510 ;
        RECT 2804.720 1573.190 2804.980 1573.510 ;
        RECT 2825.420 1573.190 2825.680 1573.510 ;
        RECT 300.080 1503.130 300.220 1573.190 ;
        RECT 2804.780 1511.970 2804.920 1573.190 ;
        RECT 2795.520 1511.650 2795.780 1511.970 ;
        RECT 2804.720 1511.650 2804.980 1511.970 ;
        RECT 2795.580 1503.130 2795.720 1511.650 ;
        RECT 300.020 1502.810 300.280 1503.130 ;
        RECT 2795.520 1502.810 2795.780 1503.130 ;
      LAYER via2 ;
        RECT 2897.630 1847.760 2897.910 1848.040 ;
        RECT 288.970 1736.240 289.250 1736.520 ;
      LAYER met3 ;
        RECT 2897.605 1848.050 2897.935 1848.065 ;
        RECT 2917.600 1848.050 2924.800 1848.500 ;
        RECT 2897.605 1847.750 2924.800 1848.050 ;
        RECT 2897.605 1847.735 2897.935 1847.750 ;
        RECT 2917.600 1847.300 2924.800 1847.750 ;
        RECT 288.945 1736.530 289.275 1736.545 ;
        RECT 300.000 1736.530 304.000 1736.600 ;
        RECT 288.945 1736.230 304.000 1736.530 ;
        RECT 288.945 1736.215 289.275 1736.230 ;
        RECT 300.000 1736.000 304.000 1736.230 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2894.850 2028.680 2895.170 2028.740 ;
        RECT 2901.290 2028.680 2901.610 2028.740 ;
        RECT 2894.850 2028.540 2901.610 2028.680 ;
        RECT 2894.850 2028.480 2895.170 2028.540 ;
        RECT 2901.290 2028.480 2901.610 2028.540 ;
        RECT 2887.950 2017.800 2888.270 2017.860 ;
        RECT 2894.850 2017.800 2895.170 2017.860 ;
        RECT 2887.950 2017.660 2895.170 2017.800 ;
        RECT 2887.950 2017.600 2888.270 2017.660 ;
        RECT 2894.850 2017.600 2895.170 2017.660 ;
        RECT 2870.470 1953.200 2870.790 1953.260 ;
        RECT 2887.950 1953.200 2888.270 1953.260 ;
        RECT 2870.470 1953.060 2888.270 1953.200 ;
        RECT 2870.470 1953.000 2870.790 1953.060 ;
        RECT 2887.950 1953.000 2888.270 1953.060 ;
        RECT 2859.890 1935.860 2860.210 1935.920 ;
        RECT 2870.470 1935.860 2870.790 1935.920 ;
        RECT 2859.890 1935.720 2870.790 1935.860 ;
        RECT 2859.890 1935.660 2860.210 1935.720 ;
        RECT 2870.470 1935.660 2870.790 1935.720 ;
        RECT 2836.890 1911.380 2837.210 1911.440 ;
        RECT 2859.890 1911.380 2860.210 1911.440 ;
        RECT 2836.890 1911.240 2860.210 1911.380 ;
        RECT 2836.890 1911.180 2837.210 1911.240 ;
        RECT 2859.890 1911.180 2860.210 1911.240 ;
        RECT 2833.210 1888.600 2833.530 1888.660 ;
        RECT 2836.890 1888.600 2837.210 1888.660 ;
        RECT 2833.210 1888.460 2837.210 1888.600 ;
        RECT 2833.210 1888.400 2833.530 1888.460 ;
        RECT 2836.890 1888.400 2837.210 1888.460 ;
        RECT 2826.310 1849.500 2826.630 1849.560 ;
        RECT 2833.210 1849.500 2833.530 1849.560 ;
        RECT 2826.310 1849.360 2833.530 1849.500 ;
        RECT 2826.310 1849.300 2826.630 1849.360 ;
        RECT 2833.210 1849.300 2833.530 1849.360 ;
        RECT 2818.950 1840.320 2819.270 1840.380 ;
        RECT 2826.310 1840.320 2826.630 1840.380 ;
        RECT 2818.950 1840.180 2826.630 1840.320 ;
        RECT 2818.950 1840.120 2819.270 1840.180 ;
        RECT 2826.310 1840.120 2826.630 1840.180 ;
        RECT 2766.510 1804.280 2766.830 1804.340 ;
        RECT 2818.950 1804.280 2819.270 1804.340 ;
        RECT 2766.510 1804.140 2819.270 1804.280 ;
        RECT 2766.510 1804.080 2766.830 1804.140 ;
        RECT 2818.950 1804.080 2819.270 1804.140 ;
        RECT 2756.390 1783.200 2756.710 1783.260 ;
        RECT 2766.510 1783.200 2766.830 1783.260 ;
        RECT 2756.390 1783.060 2766.830 1783.200 ;
        RECT 2756.390 1783.000 2756.710 1783.060 ;
        RECT 2766.510 1783.000 2766.830 1783.060 ;
        RECT 2746.270 1759.740 2746.590 1759.800 ;
        RECT 2756.390 1759.740 2756.710 1759.800 ;
        RECT 2746.270 1759.600 2756.710 1759.740 ;
        RECT 2746.270 1759.540 2746.590 1759.600 ;
        RECT 2756.390 1759.540 2756.710 1759.600 ;
        RECT 2742.590 1729.480 2742.910 1729.540 ;
        RECT 2746.270 1729.480 2746.590 1729.540 ;
        RECT 2742.590 1729.340 2746.590 1729.480 ;
        RECT 2742.590 1729.280 2742.910 1729.340 ;
        RECT 2746.270 1729.280 2746.590 1729.340 ;
        RECT 2732.470 1656.040 2732.790 1656.100 ;
        RECT 2742.590 1656.040 2742.910 1656.100 ;
        RECT 2732.470 1655.900 2742.910 1656.040 ;
        RECT 2732.470 1655.840 2732.790 1655.900 ;
        RECT 2742.590 1655.840 2742.910 1655.900 ;
        RECT 2732.470 1628.500 2732.790 1628.560 ;
        RECT 2725.660 1628.360 2732.790 1628.500 ;
        RECT 2718.670 1628.160 2718.990 1628.220 ;
        RECT 2725.660 1628.160 2725.800 1628.360 ;
        RECT 2732.470 1628.300 2732.790 1628.360 ;
        RECT 2718.670 1628.020 2725.800 1628.160 ;
        RECT 2718.670 1627.960 2718.990 1628.020 ;
        RECT 2677.270 1617.960 2677.590 1618.020 ;
        RECT 2718.670 1617.960 2718.990 1618.020 ;
        RECT 2677.270 1617.820 2718.990 1617.960 ;
        RECT 2677.270 1617.760 2677.590 1617.820 ;
        RECT 2718.670 1617.760 2718.990 1617.820 ;
        RECT 2664.390 1608.100 2664.710 1608.160 ;
        RECT 2677.270 1608.100 2677.590 1608.160 ;
        RECT 2664.390 1607.960 2677.590 1608.100 ;
        RECT 2664.390 1607.900 2664.710 1607.960 ;
        RECT 2677.270 1607.900 2677.590 1607.960 ;
        RECT 282.970 1600.620 283.290 1600.680 ;
        RECT 292.630 1600.620 292.950 1600.680 ;
        RECT 282.970 1600.480 292.950 1600.620 ;
        RECT 282.970 1600.420 283.290 1600.480 ;
        RECT 292.630 1600.420 292.950 1600.480 ;
        RECT 2647.830 1596.200 2648.150 1596.260 ;
        RECT 2664.390 1596.200 2664.710 1596.260 ;
        RECT 2647.830 1596.060 2664.710 1596.200 ;
        RECT 2647.830 1596.000 2648.150 1596.060 ;
        RECT 2664.390 1596.000 2664.710 1596.060 ;
        RECT 2647.830 1580.220 2648.150 1580.280 ;
        RECT 2622.160 1580.080 2648.150 1580.220 ;
        RECT 2617.470 1579.880 2617.790 1579.940 ;
        RECT 2622.160 1579.880 2622.300 1580.080 ;
        RECT 2647.830 1580.020 2648.150 1580.080 ;
        RECT 2617.470 1579.740 2622.300 1579.880 ;
        RECT 2617.470 1579.680 2617.790 1579.740 ;
        RECT 2612.410 1535.680 2612.730 1535.740 ;
        RECT 2617.470 1535.680 2617.790 1535.740 ;
        RECT 2612.410 1535.540 2617.790 1535.680 ;
        RECT 2612.410 1535.480 2612.730 1535.540 ;
        RECT 2617.470 1535.480 2617.790 1535.540 ;
        RECT 2587.570 1528.200 2587.890 1528.260 ;
        RECT 2612.410 1528.200 2612.730 1528.260 ;
        RECT 2587.570 1528.060 2612.730 1528.200 ;
        RECT 2587.570 1528.000 2587.890 1528.060 ;
        RECT 2612.410 1528.000 2612.730 1528.060 ;
        RECT 2573.770 1504.400 2574.090 1504.460 ;
        RECT 2587.570 1504.400 2587.890 1504.460 ;
        RECT 2573.770 1504.260 2587.890 1504.400 ;
        RECT 2573.770 1504.200 2574.090 1504.260 ;
        RECT 2587.570 1504.200 2587.890 1504.260 ;
        RECT 292.630 1500.660 292.950 1500.720 ;
        RECT 2573.770 1500.660 2574.090 1500.720 ;
        RECT 292.630 1500.520 2574.090 1500.660 ;
        RECT 292.630 1500.460 292.950 1500.520 ;
        RECT 2573.770 1500.460 2574.090 1500.520 ;
      LAYER via ;
        RECT 2894.880 2028.480 2895.140 2028.740 ;
        RECT 2901.320 2028.480 2901.580 2028.740 ;
        RECT 2887.980 2017.600 2888.240 2017.860 ;
        RECT 2894.880 2017.600 2895.140 2017.860 ;
        RECT 2870.500 1953.000 2870.760 1953.260 ;
        RECT 2887.980 1953.000 2888.240 1953.260 ;
        RECT 2859.920 1935.660 2860.180 1935.920 ;
        RECT 2870.500 1935.660 2870.760 1935.920 ;
        RECT 2836.920 1911.180 2837.180 1911.440 ;
        RECT 2859.920 1911.180 2860.180 1911.440 ;
        RECT 2833.240 1888.400 2833.500 1888.660 ;
        RECT 2836.920 1888.400 2837.180 1888.660 ;
        RECT 2826.340 1849.300 2826.600 1849.560 ;
        RECT 2833.240 1849.300 2833.500 1849.560 ;
        RECT 2818.980 1840.120 2819.240 1840.380 ;
        RECT 2826.340 1840.120 2826.600 1840.380 ;
        RECT 2766.540 1804.080 2766.800 1804.340 ;
        RECT 2818.980 1804.080 2819.240 1804.340 ;
        RECT 2756.420 1783.000 2756.680 1783.260 ;
        RECT 2766.540 1783.000 2766.800 1783.260 ;
        RECT 2746.300 1759.540 2746.560 1759.800 ;
        RECT 2756.420 1759.540 2756.680 1759.800 ;
        RECT 2742.620 1729.280 2742.880 1729.540 ;
        RECT 2746.300 1729.280 2746.560 1729.540 ;
        RECT 2732.500 1655.840 2732.760 1656.100 ;
        RECT 2742.620 1655.840 2742.880 1656.100 ;
        RECT 2718.700 1627.960 2718.960 1628.220 ;
        RECT 2732.500 1628.300 2732.760 1628.560 ;
        RECT 2677.300 1617.760 2677.560 1618.020 ;
        RECT 2718.700 1617.760 2718.960 1618.020 ;
        RECT 2664.420 1607.900 2664.680 1608.160 ;
        RECT 2677.300 1607.900 2677.560 1608.160 ;
        RECT 283.000 1600.420 283.260 1600.680 ;
        RECT 292.660 1600.420 292.920 1600.680 ;
        RECT 2647.860 1596.000 2648.120 1596.260 ;
        RECT 2664.420 1596.000 2664.680 1596.260 ;
        RECT 2617.500 1579.680 2617.760 1579.940 ;
        RECT 2647.860 1580.020 2648.120 1580.280 ;
        RECT 2612.440 1535.480 2612.700 1535.740 ;
        RECT 2617.500 1535.480 2617.760 1535.740 ;
        RECT 2587.600 1528.000 2587.860 1528.260 ;
        RECT 2612.440 1528.000 2612.700 1528.260 ;
        RECT 2573.800 1504.200 2574.060 1504.460 ;
        RECT 2587.600 1504.200 2587.860 1504.460 ;
        RECT 292.660 1500.460 292.920 1500.720 ;
        RECT 2573.800 1500.460 2574.060 1500.720 ;
      LAYER met2 ;
        RECT 2901.310 2082.315 2901.590 2082.685 ;
        RECT 2901.380 2028.770 2901.520 2082.315 ;
        RECT 2894.880 2028.450 2895.140 2028.770 ;
        RECT 2901.320 2028.450 2901.580 2028.770 ;
        RECT 2894.940 2017.890 2895.080 2028.450 ;
        RECT 2887.980 2017.570 2888.240 2017.890 ;
        RECT 2894.880 2017.570 2895.140 2017.890 ;
        RECT 2888.040 1953.290 2888.180 2017.570 ;
        RECT 2870.500 1952.970 2870.760 1953.290 ;
        RECT 2887.980 1952.970 2888.240 1953.290 ;
        RECT 2870.560 1935.950 2870.700 1952.970 ;
        RECT 2859.920 1935.630 2860.180 1935.950 ;
        RECT 2870.500 1935.630 2870.760 1935.950 ;
        RECT 2859.980 1911.470 2860.120 1935.630 ;
        RECT 2836.920 1911.150 2837.180 1911.470 ;
        RECT 2859.920 1911.150 2860.180 1911.470 ;
        RECT 2836.980 1888.690 2837.120 1911.150 ;
        RECT 2833.240 1888.370 2833.500 1888.690 ;
        RECT 2836.920 1888.370 2837.180 1888.690 ;
        RECT 2833.300 1849.590 2833.440 1888.370 ;
        RECT 2826.340 1849.270 2826.600 1849.590 ;
        RECT 2833.240 1849.270 2833.500 1849.590 ;
        RECT 2826.400 1840.410 2826.540 1849.270 ;
        RECT 2818.980 1840.090 2819.240 1840.410 ;
        RECT 2826.340 1840.090 2826.600 1840.410 ;
        RECT 2819.040 1804.370 2819.180 1840.090 ;
        RECT 2766.540 1804.050 2766.800 1804.370 ;
        RECT 2818.980 1804.050 2819.240 1804.370 ;
        RECT 2766.600 1783.290 2766.740 1804.050 ;
        RECT 2756.420 1782.970 2756.680 1783.290 ;
        RECT 2766.540 1782.970 2766.800 1783.290 ;
        RECT 282.990 1768.155 283.270 1768.525 ;
        RECT 283.060 1600.710 283.200 1768.155 ;
        RECT 2756.480 1759.830 2756.620 1782.970 ;
        RECT 2746.300 1759.510 2746.560 1759.830 ;
        RECT 2756.420 1759.510 2756.680 1759.830 ;
        RECT 2746.360 1729.570 2746.500 1759.510 ;
        RECT 2742.620 1729.250 2742.880 1729.570 ;
        RECT 2746.300 1729.250 2746.560 1729.570 ;
        RECT 2742.680 1656.130 2742.820 1729.250 ;
        RECT 2732.500 1655.810 2732.760 1656.130 ;
        RECT 2742.620 1655.810 2742.880 1656.130 ;
        RECT 2732.560 1628.590 2732.700 1655.810 ;
        RECT 2732.500 1628.270 2732.760 1628.590 ;
        RECT 2718.700 1627.930 2718.960 1628.250 ;
        RECT 2718.760 1618.050 2718.900 1627.930 ;
        RECT 2677.300 1617.730 2677.560 1618.050 ;
        RECT 2718.700 1617.730 2718.960 1618.050 ;
        RECT 2677.360 1608.190 2677.500 1617.730 ;
        RECT 2664.420 1607.870 2664.680 1608.190 ;
        RECT 2677.300 1607.870 2677.560 1608.190 ;
        RECT 283.000 1600.390 283.260 1600.710 ;
        RECT 292.660 1600.390 292.920 1600.710 ;
        RECT 292.720 1500.750 292.860 1600.390 ;
        RECT 2664.480 1596.290 2664.620 1607.870 ;
        RECT 2647.860 1595.970 2648.120 1596.290 ;
        RECT 2664.420 1595.970 2664.680 1596.290 ;
        RECT 2647.920 1580.310 2648.060 1595.970 ;
        RECT 2647.860 1579.990 2648.120 1580.310 ;
        RECT 2617.500 1579.650 2617.760 1579.970 ;
        RECT 2617.560 1535.770 2617.700 1579.650 ;
        RECT 2612.440 1535.450 2612.700 1535.770 ;
        RECT 2617.500 1535.450 2617.760 1535.770 ;
        RECT 2612.500 1528.290 2612.640 1535.450 ;
        RECT 2587.600 1527.970 2587.860 1528.290 ;
        RECT 2612.440 1527.970 2612.700 1528.290 ;
        RECT 2587.660 1504.490 2587.800 1527.970 ;
        RECT 2573.800 1504.170 2574.060 1504.490 ;
        RECT 2587.600 1504.170 2587.860 1504.490 ;
        RECT 2573.860 1500.750 2574.000 1504.170 ;
        RECT 292.660 1500.430 292.920 1500.750 ;
        RECT 2573.800 1500.430 2574.060 1500.750 ;
      LAYER via2 ;
        RECT 2901.310 2082.360 2901.590 2082.640 ;
        RECT 282.990 1768.200 283.270 1768.480 ;
      LAYER met3 ;
        RECT 2901.285 2082.650 2901.615 2082.665 ;
        RECT 2917.600 2082.650 2924.800 2083.100 ;
        RECT 2901.285 2082.350 2924.800 2082.650 ;
        RECT 2901.285 2082.335 2901.615 2082.350 ;
        RECT 2917.600 2081.900 2924.800 2082.350 ;
        RECT 282.965 1768.490 283.295 1768.505 ;
        RECT 300.000 1768.490 304.000 1768.560 ;
        RECT 282.965 1768.190 304.000 1768.490 ;
        RECT 282.965 1768.175 283.295 1768.190 ;
        RECT 300.000 1767.960 304.000 1768.190 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2884.270 2310.200 2884.590 2310.260 ;
        RECT 2899.910 2310.200 2900.230 2310.260 ;
        RECT 2884.270 2310.060 2900.230 2310.200 ;
        RECT 2884.270 2310.000 2884.590 2310.060 ;
        RECT 2899.910 2310.000 2900.230 2310.060 ;
        RECT 2858.970 2297.960 2859.290 2298.020 ;
        RECT 2884.270 2297.960 2884.590 2298.020 ;
        RECT 2858.970 2297.820 2884.590 2297.960 ;
        RECT 2858.970 2297.760 2859.290 2297.820 ;
        RECT 2884.270 2297.760 2884.590 2297.820 ;
        RECT 2832.290 2280.280 2832.610 2280.340 ;
        RECT 2858.970 2280.280 2859.290 2280.340 ;
        RECT 2832.290 2280.140 2859.290 2280.280 ;
        RECT 2832.290 2280.080 2832.610 2280.140 ;
        RECT 2858.970 2280.080 2859.290 2280.140 ;
        RECT 2832.290 2228.940 2832.610 2229.000 ;
        RECT 2822.260 2228.800 2832.610 2228.940 ;
        RECT 2816.190 2228.600 2816.510 2228.660 ;
        RECT 2822.260 2228.600 2822.400 2228.800 ;
        RECT 2832.290 2228.740 2832.610 2228.800 ;
        RECT 2816.190 2228.460 2822.400 2228.600 ;
        RECT 2816.190 2228.400 2816.510 2228.460 ;
        RECT 2812.050 2210.920 2812.370 2210.980 ;
        RECT 2816.190 2210.920 2816.510 2210.980 ;
        RECT 2812.050 2210.780 2816.510 2210.920 ;
        RECT 2812.050 2210.720 2812.370 2210.780 ;
        RECT 2816.190 2210.720 2816.510 2210.780 ;
        RECT 2804.690 2194.600 2805.010 2194.660 ;
        RECT 2812.050 2194.600 2812.370 2194.660 ;
        RECT 2804.690 2194.460 2812.370 2194.600 ;
        RECT 2804.690 2194.400 2805.010 2194.460 ;
        RECT 2812.050 2194.400 2812.370 2194.460 ;
        RECT 2790.890 2090.900 2791.210 2090.960 ;
        RECT 2804.690 2090.900 2805.010 2090.960 ;
        RECT 2790.890 2090.760 2805.010 2090.900 ;
        RECT 2790.890 2090.700 2791.210 2090.760 ;
        RECT 2804.690 2090.700 2805.010 2090.760 ;
        RECT 2783.990 1998.420 2784.310 1998.480 ;
        RECT 2790.890 1998.420 2791.210 1998.480 ;
        RECT 2783.990 1998.280 2791.210 1998.420 ;
        RECT 2783.990 1998.220 2784.310 1998.280 ;
        RECT 2790.890 1998.220 2791.210 1998.280 ;
        RECT 2777.090 1938.920 2777.410 1938.980 ;
        RECT 2783.990 1938.920 2784.310 1938.980 ;
        RECT 2777.090 1938.780 2784.310 1938.920 ;
        RECT 2777.090 1938.720 2777.410 1938.780 ;
        RECT 2783.990 1938.720 2784.310 1938.780 ;
        RECT 2770.190 1759.740 2770.510 1759.800 ;
        RECT 2777.090 1759.740 2777.410 1759.800 ;
        RECT 2770.190 1759.600 2777.410 1759.740 ;
        RECT 2770.190 1759.540 2770.510 1759.600 ;
        RECT 2777.090 1759.540 2777.410 1759.600 ;
        RECT 2763.290 1711.460 2763.610 1711.520 ;
        RECT 2770.190 1711.460 2770.510 1711.520 ;
        RECT 2763.290 1711.320 2770.510 1711.460 ;
        RECT 2763.290 1711.260 2763.610 1711.320 ;
        RECT 2770.190 1711.260 2770.510 1711.320 ;
        RECT 288.490 1683.580 288.810 1683.640 ;
        RECT 293.090 1683.580 293.410 1683.640 ;
        RECT 288.490 1683.440 293.410 1683.580 ;
        RECT 288.490 1683.380 288.810 1683.440 ;
        RECT 293.090 1683.380 293.410 1683.440 ;
        RECT 2756.390 1669.980 2756.710 1670.040 ;
        RECT 2763.290 1669.980 2763.610 1670.040 ;
        RECT 2756.390 1669.840 2763.610 1669.980 ;
        RECT 2756.390 1669.780 2756.710 1669.840 ;
        RECT 2763.290 1669.780 2763.610 1669.840 ;
        RECT 2742.590 1603.680 2742.910 1603.740 ;
        RECT 2756.390 1603.680 2756.710 1603.740 ;
        RECT 2742.590 1603.540 2756.710 1603.680 ;
        RECT 2742.590 1603.480 2742.910 1603.540 ;
        RECT 2756.390 1603.480 2756.710 1603.540 ;
        RECT 2732.470 1525.140 2732.790 1525.200 ;
        RECT 2742.590 1525.140 2742.910 1525.200 ;
        RECT 2732.470 1525.000 2742.910 1525.140 ;
        RECT 2732.470 1524.940 2732.790 1525.000 ;
        RECT 2742.590 1524.940 2742.910 1525.000 ;
        RECT 293.090 1502.360 293.410 1502.420 ;
        RECT 2732.470 1502.360 2732.790 1502.420 ;
        RECT 293.090 1502.220 2732.790 1502.360 ;
        RECT 293.090 1502.160 293.410 1502.220 ;
        RECT 2732.470 1502.160 2732.790 1502.220 ;
      LAYER via ;
        RECT 2884.300 2310.000 2884.560 2310.260 ;
        RECT 2899.940 2310.000 2900.200 2310.260 ;
        RECT 2859.000 2297.760 2859.260 2298.020 ;
        RECT 2884.300 2297.760 2884.560 2298.020 ;
        RECT 2832.320 2280.080 2832.580 2280.340 ;
        RECT 2859.000 2280.080 2859.260 2280.340 ;
        RECT 2816.220 2228.400 2816.480 2228.660 ;
        RECT 2832.320 2228.740 2832.580 2229.000 ;
        RECT 2812.080 2210.720 2812.340 2210.980 ;
        RECT 2816.220 2210.720 2816.480 2210.980 ;
        RECT 2804.720 2194.400 2804.980 2194.660 ;
        RECT 2812.080 2194.400 2812.340 2194.660 ;
        RECT 2790.920 2090.700 2791.180 2090.960 ;
        RECT 2804.720 2090.700 2804.980 2090.960 ;
        RECT 2784.020 1998.220 2784.280 1998.480 ;
        RECT 2790.920 1998.220 2791.180 1998.480 ;
        RECT 2777.120 1938.720 2777.380 1938.980 ;
        RECT 2784.020 1938.720 2784.280 1938.980 ;
        RECT 2770.220 1759.540 2770.480 1759.800 ;
        RECT 2777.120 1759.540 2777.380 1759.800 ;
        RECT 2763.320 1711.260 2763.580 1711.520 ;
        RECT 2770.220 1711.260 2770.480 1711.520 ;
        RECT 288.520 1683.380 288.780 1683.640 ;
        RECT 293.120 1683.380 293.380 1683.640 ;
        RECT 2756.420 1669.780 2756.680 1670.040 ;
        RECT 2763.320 1669.780 2763.580 1670.040 ;
        RECT 2742.620 1603.480 2742.880 1603.740 ;
        RECT 2756.420 1603.480 2756.680 1603.740 ;
        RECT 2732.500 1524.940 2732.760 1525.200 ;
        RECT 2742.620 1524.940 2742.880 1525.200 ;
        RECT 293.120 1502.160 293.380 1502.420 ;
        RECT 2732.500 1502.160 2732.760 1502.420 ;
      LAYER met2 ;
        RECT 2899.930 2316.915 2900.210 2317.285 ;
        RECT 2900.000 2310.290 2900.140 2316.915 ;
        RECT 2884.300 2309.970 2884.560 2310.290 ;
        RECT 2899.940 2309.970 2900.200 2310.290 ;
        RECT 2884.360 2298.050 2884.500 2309.970 ;
        RECT 2859.000 2297.730 2859.260 2298.050 ;
        RECT 2884.300 2297.730 2884.560 2298.050 ;
        RECT 2859.060 2280.370 2859.200 2297.730 ;
        RECT 2832.320 2280.050 2832.580 2280.370 ;
        RECT 2859.000 2280.050 2859.260 2280.370 ;
        RECT 2832.380 2229.030 2832.520 2280.050 ;
        RECT 2832.320 2228.710 2832.580 2229.030 ;
        RECT 2816.220 2228.370 2816.480 2228.690 ;
        RECT 2816.280 2211.010 2816.420 2228.370 ;
        RECT 2812.080 2210.690 2812.340 2211.010 ;
        RECT 2816.220 2210.690 2816.480 2211.010 ;
        RECT 2812.140 2194.690 2812.280 2210.690 ;
        RECT 2804.720 2194.370 2804.980 2194.690 ;
        RECT 2812.080 2194.370 2812.340 2194.690 ;
        RECT 2804.780 2090.990 2804.920 2194.370 ;
        RECT 2790.920 2090.670 2791.180 2090.990 ;
        RECT 2804.720 2090.670 2804.980 2090.990 ;
        RECT 2790.980 1998.510 2791.120 2090.670 ;
        RECT 2784.020 1998.190 2784.280 1998.510 ;
        RECT 2790.920 1998.190 2791.180 1998.510 ;
        RECT 2784.080 1939.010 2784.220 1998.190 ;
        RECT 2777.120 1938.690 2777.380 1939.010 ;
        RECT 2784.020 1938.690 2784.280 1939.010 ;
        RECT 288.510 1799.435 288.790 1799.805 ;
        RECT 288.580 1683.670 288.720 1799.435 ;
        RECT 2777.180 1759.830 2777.320 1938.690 ;
        RECT 2770.220 1759.510 2770.480 1759.830 ;
        RECT 2777.120 1759.510 2777.380 1759.830 ;
        RECT 2770.280 1711.550 2770.420 1759.510 ;
        RECT 2763.320 1711.230 2763.580 1711.550 ;
        RECT 2770.220 1711.230 2770.480 1711.550 ;
        RECT 288.520 1683.350 288.780 1683.670 ;
        RECT 293.120 1683.350 293.380 1683.670 ;
        RECT 293.180 1502.450 293.320 1683.350 ;
        RECT 2763.380 1670.070 2763.520 1711.230 ;
        RECT 2756.420 1669.750 2756.680 1670.070 ;
        RECT 2763.320 1669.750 2763.580 1670.070 ;
        RECT 2756.480 1603.770 2756.620 1669.750 ;
        RECT 2742.620 1603.450 2742.880 1603.770 ;
        RECT 2756.420 1603.450 2756.680 1603.770 ;
        RECT 2742.680 1525.230 2742.820 1603.450 ;
        RECT 2732.500 1524.910 2732.760 1525.230 ;
        RECT 2742.620 1524.910 2742.880 1525.230 ;
        RECT 2732.560 1502.450 2732.700 1524.910 ;
        RECT 293.120 1502.130 293.380 1502.450 ;
        RECT 2732.500 1502.130 2732.760 1502.450 ;
      LAYER via2 ;
        RECT 2899.930 2316.960 2900.210 2317.240 ;
        RECT 288.510 1799.480 288.790 1799.760 ;
      LAYER met3 ;
        RECT 2899.905 2317.250 2900.235 2317.265 ;
        RECT 2917.600 2317.250 2924.800 2317.700 ;
        RECT 2899.905 2316.950 2924.800 2317.250 ;
        RECT 2899.905 2316.935 2900.235 2316.950 ;
        RECT 2917.600 2316.500 2924.800 2316.950 ;
        RECT 288.485 1799.770 288.815 1799.785 ;
        RECT 300.000 1799.770 304.000 1799.840 ;
        RECT 288.485 1799.470 304.000 1799.770 ;
        RECT 288.485 1799.455 288.815 1799.470 ;
        RECT 300.000 1799.240 304.000 1799.470 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 737.910 146.100 738.230 146.160 ;
        RECT 772.410 146.100 772.730 146.160 ;
        RECT 737.910 145.960 772.730 146.100 ;
        RECT 737.910 145.900 738.230 145.960 ;
        RECT 772.410 145.900 772.730 145.960 ;
        RECT 579.670 145.420 579.990 145.480 ;
        RECT 604.050 145.420 604.370 145.480 ;
        RECT 579.670 145.280 604.370 145.420 ;
        RECT 579.670 145.220 579.990 145.280 ;
        RECT 604.050 145.220 604.370 145.280 ;
      LAYER via ;
        RECT 737.940 145.900 738.200 146.160 ;
        RECT 772.440 145.900 772.700 146.160 ;
        RECT 579.700 145.220 579.960 145.480 ;
        RECT 604.080 145.220 604.340 145.480 ;
      LAYER met2 ;
        RECT 458.710 147.715 458.990 148.085 ;
        RECT 458.780 146.045 458.920 147.715 ;
        RECT 717.230 147.035 717.510 147.405 ;
        RECT 604.070 146.355 604.350 146.725 ;
        RECT 641.330 146.355 641.610 146.725 ;
        RECT 458.710 145.675 458.990 146.045 ;
        RECT 604.140 145.510 604.280 146.355 ;
        RECT 641.400 145.930 641.540 146.355 ;
        RECT 642.250 145.930 642.530 146.045 ;
        RECT 641.400 145.790 642.530 145.930 ;
        RECT 642.250 145.675 642.530 145.790 ;
        RECT 579.700 145.365 579.960 145.510 ;
        RECT 579.690 144.995 579.970 145.365 ;
        RECT 604.080 145.190 604.340 145.510 ;
        RECT 717.300 145.365 717.440 147.035 ;
        RECT 772.430 146.355 772.710 146.725 ;
        RECT 772.500 146.190 772.640 146.355 ;
        RECT 737.940 146.045 738.200 146.190 ;
        RECT 737.930 145.675 738.210 146.045 ;
        RECT 772.440 145.870 772.700 146.190 ;
        RECT 717.230 144.995 717.510 145.365 ;
      LAYER via2 ;
        RECT 458.710 147.760 458.990 148.040 ;
        RECT 717.230 147.080 717.510 147.360 ;
        RECT 604.070 146.400 604.350 146.680 ;
        RECT 641.330 146.400 641.610 146.680 ;
        RECT 458.710 145.720 458.990 146.000 ;
        RECT 642.250 145.720 642.530 146.000 ;
        RECT 579.690 145.040 579.970 145.320 ;
        RECT 772.430 146.400 772.710 146.680 ;
        RECT 737.930 145.720 738.210 146.000 ;
        RECT 717.230 145.040 717.510 145.320 ;
      LAYER met3 ;
        RECT 289.150 1525.730 289.530 1525.740 ;
        RECT 300.000 1525.730 304.000 1525.800 ;
        RECT 289.150 1525.430 304.000 1525.730 ;
        RECT 289.150 1525.420 289.530 1525.430 ;
        RECT 300.000 1525.200 304.000 1525.430 ;
        RECT 434.510 148.050 434.890 148.060 ;
        RECT 458.685 148.050 459.015 148.065 ;
        RECT 434.510 147.750 459.015 148.050 ;
        RECT 434.510 147.740 434.890 147.750 ;
        RECT 458.685 147.735 459.015 147.750 ;
        RECT 578.950 147.370 579.330 147.380 ;
        RECT 544.030 147.070 579.330 147.370 ;
        RECT 289.150 146.690 289.530 146.700 ;
        RECT 289.150 146.390 398.970 146.690 ;
        RECT 289.150 146.380 289.530 146.390 ;
        RECT 398.670 146.010 398.970 146.390 ;
        RECT 434.510 146.010 434.890 146.020 ;
        RECT 398.670 145.710 434.890 146.010 ;
        RECT 434.510 145.700 434.890 145.710 ;
        RECT 458.685 146.010 459.015 146.025 ;
        RECT 544.030 146.010 544.330 147.070 ;
        RECT 578.950 147.060 579.330 147.070 ;
        RECT 669.110 147.370 669.490 147.380 ;
        RECT 717.205 147.370 717.535 147.385 ;
        RECT 669.110 147.070 717.535 147.370 ;
        RECT 669.110 147.060 669.490 147.070 ;
        RECT 717.205 147.055 717.535 147.070 ;
        RECT 604.045 146.690 604.375 146.705 ;
        RECT 641.305 146.690 641.635 146.705 ;
        RECT 604.045 146.390 641.635 146.690 ;
        RECT 604.045 146.375 604.375 146.390 ;
        RECT 641.305 146.375 641.635 146.390 ;
        RECT 772.405 146.690 772.735 146.705 ;
        RECT 2917.600 146.690 2924.800 147.140 ;
        RECT 772.405 146.390 807.450 146.690 ;
        RECT 772.405 146.375 772.735 146.390 ;
        RECT 458.685 145.710 482.690 146.010 ;
        RECT 458.685 145.695 459.015 145.710 ;
        RECT 482.390 145.330 482.690 145.710 ;
        RECT 497.110 145.710 544.330 146.010 ;
        RECT 642.225 146.010 642.555 146.025 ;
        RECT 669.110 146.010 669.490 146.020 ;
        RECT 737.905 146.010 738.235 146.025 ;
        RECT 642.225 145.710 669.490 146.010 ;
        RECT 497.110 145.330 497.410 145.710 ;
        RECT 642.225 145.695 642.555 145.710 ;
        RECT 669.110 145.700 669.490 145.710 ;
        RECT 724.350 145.710 738.235 146.010 ;
        RECT 807.150 146.010 807.450 146.390 ;
        RECT 855.910 146.390 904.050 146.690 ;
        RECT 807.150 145.710 855.290 146.010 ;
        RECT 482.390 145.030 497.410 145.330 ;
        RECT 578.950 145.330 579.330 145.340 ;
        RECT 579.665 145.330 579.995 145.345 ;
        RECT 578.950 145.030 579.995 145.330 ;
        RECT 578.950 145.020 579.330 145.030 ;
        RECT 579.665 145.015 579.995 145.030 ;
        RECT 717.205 145.330 717.535 145.345 ;
        RECT 724.350 145.330 724.650 145.710 ;
        RECT 737.905 145.695 738.235 145.710 ;
        RECT 717.205 145.030 724.650 145.330 ;
        RECT 854.990 145.330 855.290 145.710 ;
        RECT 855.910 145.330 856.210 146.390 ;
        RECT 903.750 146.010 904.050 146.390 ;
        RECT 952.510 146.390 1000.650 146.690 ;
        RECT 903.750 145.710 951.890 146.010 ;
        RECT 854.990 145.030 856.210 145.330 ;
        RECT 951.590 145.330 951.890 145.710 ;
        RECT 952.510 145.330 952.810 146.390 ;
        RECT 1000.350 146.010 1000.650 146.390 ;
        RECT 1049.110 146.390 1097.250 146.690 ;
        RECT 1000.350 145.710 1048.490 146.010 ;
        RECT 951.590 145.030 952.810 145.330 ;
        RECT 1048.190 145.330 1048.490 145.710 ;
        RECT 1049.110 145.330 1049.410 146.390 ;
        RECT 1096.950 146.010 1097.250 146.390 ;
        RECT 1145.710 146.390 1193.850 146.690 ;
        RECT 1096.950 145.710 1145.090 146.010 ;
        RECT 1048.190 145.030 1049.410 145.330 ;
        RECT 1144.790 145.330 1145.090 145.710 ;
        RECT 1145.710 145.330 1146.010 146.390 ;
        RECT 1193.550 146.010 1193.850 146.390 ;
        RECT 1242.310 146.390 1290.450 146.690 ;
        RECT 1193.550 145.710 1241.690 146.010 ;
        RECT 1144.790 145.030 1146.010 145.330 ;
        RECT 1241.390 145.330 1241.690 145.710 ;
        RECT 1242.310 145.330 1242.610 146.390 ;
        RECT 1290.150 146.010 1290.450 146.390 ;
        RECT 1338.910 146.390 1387.050 146.690 ;
        RECT 1290.150 145.710 1338.290 146.010 ;
        RECT 1241.390 145.030 1242.610 145.330 ;
        RECT 1337.990 145.330 1338.290 145.710 ;
        RECT 1338.910 145.330 1339.210 146.390 ;
        RECT 1386.750 146.010 1387.050 146.390 ;
        RECT 1435.510 146.390 1483.650 146.690 ;
        RECT 1386.750 145.710 1434.890 146.010 ;
        RECT 1337.990 145.030 1339.210 145.330 ;
        RECT 1434.590 145.330 1434.890 145.710 ;
        RECT 1435.510 145.330 1435.810 146.390 ;
        RECT 1483.350 146.010 1483.650 146.390 ;
        RECT 1532.110 146.390 1580.250 146.690 ;
        RECT 1483.350 145.710 1531.490 146.010 ;
        RECT 1434.590 145.030 1435.810 145.330 ;
        RECT 1531.190 145.330 1531.490 145.710 ;
        RECT 1532.110 145.330 1532.410 146.390 ;
        RECT 1579.950 146.010 1580.250 146.390 ;
        RECT 1628.710 146.390 1676.850 146.690 ;
        RECT 1579.950 145.710 1628.090 146.010 ;
        RECT 1531.190 145.030 1532.410 145.330 ;
        RECT 1627.790 145.330 1628.090 145.710 ;
        RECT 1628.710 145.330 1629.010 146.390 ;
        RECT 1676.550 146.010 1676.850 146.390 ;
        RECT 1725.310 146.390 1773.450 146.690 ;
        RECT 1676.550 145.710 1724.690 146.010 ;
        RECT 1627.790 145.030 1629.010 145.330 ;
        RECT 1724.390 145.330 1724.690 145.710 ;
        RECT 1725.310 145.330 1725.610 146.390 ;
        RECT 1773.150 146.010 1773.450 146.390 ;
        RECT 1821.910 146.390 1870.050 146.690 ;
        RECT 1773.150 145.710 1821.290 146.010 ;
        RECT 1724.390 145.030 1725.610 145.330 ;
        RECT 1820.990 145.330 1821.290 145.710 ;
        RECT 1821.910 145.330 1822.210 146.390 ;
        RECT 1869.750 146.010 1870.050 146.390 ;
        RECT 1918.510 146.390 1966.650 146.690 ;
        RECT 1869.750 145.710 1917.890 146.010 ;
        RECT 1820.990 145.030 1822.210 145.330 ;
        RECT 1917.590 145.330 1917.890 145.710 ;
        RECT 1918.510 145.330 1918.810 146.390 ;
        RECT 1966.350 146.010 1966.650 146.390 ;
        RECT 2015.110 146.390 2063.250 146.690 ;
        RECT 1966.350 145.710 2014.490 146.010 ;
        RECT 1917.590 145.030 1918.810 145.330 ;
        RECT 2014.190 145.330 2014.490 145.710 ;
        RECT 2015.110 145.330 2015.410 146.390 ;
        RECT 2062.950 146.010 2063.250 146.390 ;
        RECT 2111.710 146.390 2159.850 146.690 ;
        RECT 2062.950 145.710 2111.090 146.010 ;
        RECT 2014.190 145.030 2015.410 145.330 ;
        RECT 2110.790 145.330 2111.090 145.710 ;
        RECT 2111.710 145.330 2112.010 146.390 ;
        RECT 2159.550 146.010 2159.850 146.390 ;
        RECT 2208.310 146.390 2256.450 146.690 ;
        RECT 2159.550 145.710 2207.690 146.010 ;
        RECT 2110.790 145.030 2112.010 145.330 ;
        RECT 2207.390 145.330 2207.690 145.710 ;
        RECT 2208.310 145.330 2208.610 146.390 ;
        RECT 2256.150 146.010 2256.450 146.390 ;
        RECT 2304.910 146.390 2353.050 146.690 ;
        RECT 2256.150 145.710 2304.290 146.010 ;
        RECT 2207.390 145.030 2208.610 145.330 ;
        RECT 2303.990 145.330 2304.290 145.710 ;
        RECT 2304.910 145.330 2305.210 146.390 ;
        RECT 2352.750 146.010 2353.050 146.390 ;
        RECT 2401.510 146.390 2449.650 146.690 ;
        RECT 2352.750 145.710 2400.890 146.010 ;
        RECT 2303.990 145.030 2305.210 145.330 ;
        RECT 2400.590 145.330 2400.890 145.710 ;
        RECT 2401.510 145.330 2401.810 146.390 ;
        RECT 2449.350 146.010 2449.650 146.390 ;
        RECT 2498.110 146.390 2546.250 146.690 ;
        RECT 2449.350 145.710 2497.490 146.010 ;
        RECT 2400.590 145.030 2401.810 145.330 ;
        RECT 2497.190 145.330 2497.490 145.710 ;
        RECT 2498.110 145.330 2498.410 146.390 ;
        RECT 2545.950 146.010 2546.250 146.390 ;
        RECT 2594.710 146.390 2642.850 146.690 ;
        RECT 2545.950 145.710 2594.090 146.010 ;
        RECT 2497.190 145.030 2498.410 145.330 ;
        RECT 2593.790 145.330 2594.090 145.710 ;
        RECT 2594.710 145.330 2595.010 146.390 ;
        RECT 2642.550 146.010 2642.850 146.390 ;
        RECT 2691.310 146.390 2739.450 146.690 ;
        RECT 2642.550 145.710 2690.690 146.010 ;
        RECT 2593.790 145.030 2595.010 145.330 ;
        RECT 2690.390 145.330 2690.690 145.710 ;
        RECT 2691.310 145.330 2691.610 146.390 ;
        RECT 2739.150 146.010 2739.450 146.390 ;
        RECT 2787.910 146.390 2836.050 146.690 ;
        RECT 2739.150 145.710 2787.290 146.010 ;
        RECT 2690.390 145.030 2691.610 145.330 ;
        RECT 2786.990 145.330 2787.290 145.710 ;
        RECT 2787.910 145.330 2788.210 146.390 ;
        RECT 2835.750 146.010 2836.050 146.390 ;
        RECT 2916.710 146.390 2924.800 146.690 ;
        RECT 2916.710 146.010 2917.010 146.390 ;
        RECT 2835.750 145.710 2883.890 146.010 ;
        RECT 2786.990 145.030 2788.210 145.330 ;
        RECT 2883.590 145.330 2883.890 145.710 ;
        RECT 2884.510 145.710 2917.010 146.010 ;
        RECT 2917.600 145.940 2924.800 146.390 ;
        RECT 2884.510 145.330 2884.810 145.710 ;
        RECT 2883.590 145.030 2884.810 145.330 ;
        RECT 717.205 145.015 717.535 145.030 ;
      LAYER via3 ;
        RECT 289.180 1525.420 289.500 1525.740 ;
        RECT 434.540 147.740 434.860 148.060 ;
        RECT 289.180 146.380 289.500 146.700 ;
        RECT 434.540 145.700 434.860 146.020 ;
        RECT 578.980 147.060 579.300 147.380 ;
        RECT 669.140 147.060 669.460 147.380 ;
        RECT 669.140 145.700 669.460 146.020 ;
        RECT 578.980 145.020 579.300 145.340 ;
      LAYER met4 ;
        RECT 289.175 1525.415 289.505 1525.745 ;
        RECT 289.190 146.705 289.490 1525.415 ;
        RECT 434.535 147.735 434.865 148.065 ;
        RECT 289.175 146.375 289.505 146.705 ;
        RECT 434.550 146.025 434.850 147.735 ;
        RECT 578.975 147.055 579.305 147.385 ;
        RECT 669.135 147.055 669.465 147.385 ;
        RECT 434.535 145.695 434.865 146.025 ;
        RECT 578.990 145.345 579.290 147.055 ;
        RECT 669.150 146.025 669.450 147.055 ;
        RECT 669.135 145.695 669.465 146.025 ;
        RECT 578.975 145.015 579.305 145.345 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 303.670 2692.020 303.990 2692.080 ;
        RECT 2708.090 2692.020 2708.410 2692.080 ;
        RECT 303.670 2691.880 2708.410 2692.020 ;
        RECT 303.670 2691.820 303.990 2691.880 ;
        RECT 2708.090 2691.820 2708.410 2691.880 ;
        RECT 300.450 2684.200 300.770 2684.260 ;
        RECT 303.670 2684.200 303.990 2684.260 ;
        RECT 300.450 2684.060 303.990 2684.200 ;
        RECT 300.450 2684.000 300.770 2684.060 ;
        RECT 303.670 2684.000 303.990 2684.060 ;
        RECT 2708.090 2652.920 2708.410 2652.980 ;
        RECT 2780.770 2652.920 2781.090 2652.980 ;
        RECT 2708.090 2652.780 2781.090 2652.920 ;
        RECT 2708.090 2652.720 2708.410 2652.780 ;
        RECT 2780.770 2652.720 2781.090 2652.780 ;
        RECT 2780.770 2646.120 2781.090 2646.180 ;
        RECT 2842.410 2646.120 2842.730 2646.180 ;
        RECT 2780.770 2645.980 2842.730 2646.120 ;
        RECT 2780.770 2645.920 2781.090 2645.980 ;
        RECT 2842.410 2645.920 2842.730 2645.980 ;
        RECT 2842.410 2629.120 2842.730 2629.180 ;
        RECT 2842.410 2628.980 2843.100 2629.120 ;
        RECT 2842.410 2628.920 2842.730 2628.980 ;
        RECT 2842.960 2628.780 2843.100 2628.980 ;
        RECT 2859.890 2628.780 2860.210 2628.840 ;
        RECT 2842.960 2628.640 2860.210 2628.780 ;
        RECT 2859.890 2628.580 2860.210 2628.640 ;
        RECT 2859.890 2566.560 2860.210 2566.620 ;
        RECT 2873.690 2566.560 2874.010 2566.620 ;
        RECT 2859.890 2566.420 2874.010 2566.560 ;
        RECT 2859.890 2566.360 2860.210 2566.420 ;
        RECT 2873.690 2566.360 2874.010 2566.420 ;
        RECT 2873.690 2539.020 2874.010 2539.080 ;
        RECT 2889.790 2539.020 2890.110 2539.080 ;
        RECT 2873.690 2538.880 2890.110 2539.020 ;
        RECT 2873.690 2538.820 2874.010 2538.880 ;
        RECT 2889.790 2538.820 2890.110 2538.880 ;
        RECT 2889.790 2531.540 2890.110 2531.600 ;
        RECT 2901.290 2531.540 2901.610 2531.600 ;
        RECT 2889.790 2531.400 2901.610 2531.540 ;
        RECT 2889.790 2531.340 2890.110 2531.400 ;
        RECT 2901.290 2531.340 2901.610 2531.400 ;
        RECT 288.030 2170.120 288.350 2170.180 ;
        RECT 300.450 2170.120 300.770 2170.180 ;
        RECT 288.030 2169.980 300.770 2170.120 ;
        RECT 288.030 2169.920 288.350 2169.980 ;
        RECT 300.450 2169.920 300.770 2169.980 ;
      LAYER via ;
        RECT 303.700 2691.820 303.960 2692.080 ;
        RECT 2708.120 2691.820 2708.380 2692.080 ;
        RECT 300.480 2684.000 300.740 2684.260 ;
        RECT 303.700 2684.000 303.960 2684.260 ;
        RECT 2708.120 2652.720 2708.380 2652.980 ;
        RECT 2780.800 2652.720 2781.060 2652.980 ;
        RECT 2780.800 2645.920 2781.060 2646.180 ;
        RECT 2842.440 2645.920 2842.700 2646.180 ;
        RECT 2842.440 2628.920 2842.700 2629.180 ;
        RECT 2859.920 2628.580 2860.180 2628.840 ;
        RECT 2859.920 2566.360 2860.180 2566.620 ;
        RECT 2873.720 2566.360 2873.980 2566.620 ;
        RECT 2873.720 2538.820 2873.980 2539.080 ;
        RECT 2889.820 2538.820 2890.080 2539.080 ;
        RECT 2889.820 2531.340 2890.080 2531.600 ;
        RECT 2901.320 2531.340 2901.580 2531.600 ;
        RECT 288.060 2169.920 288.320 2170.180 ;
        RECT 300.480 2169.920 300.740 2170.180 ;
      LAYER met2 ;
        RECT 303.700 2691.790 303.960 2692.110 ;
        RECT 2708.120 2691.790 2708.380 2692.110 ;
        RECT 303.760 2684.290 303.900 2691.790 ;
        RECT 300.480 2683.970 300.740 2684.290 ;
        RECT 303.700 2683.970 303.960 2684.290 ;
        RECT 300.540 2170.210 300.680 2683.970 ;
        RECT 2708.180 2653.010 2708.320 2691.790 ;
        RECT 2708.120 2652.690 2708.380 2653.010 ;
        RECT 2780.800 2652.690 2781.060 2653.010 ;
        RECT 2780.860 2646.210 2781.000 2652.690 ;
        RECT 2780.800 2645.890 2781.060 2646.210 ;
        RECT 2842.440 2645.890 2842.700 2646.210 ;
        RECT 2842.500 2629.210 2842.640 2645.890 ;
        RECT 2842.440 2628.890 2842.700 2629.210 ;
        RECT 2859.920 2628.550 2860.180 2628.870 ;
        RECT 2859.980 2566.650 2860.120 2628.550 ;
        RECT 2859.920 2566.330 2860.180 2566.650 ;
        RECT 2873.720 2566.330 2873.980 2566.650 ;
        RECT 2873.780 2539.110 2873.920 2566.330 ;
        RECT 2873.720 2538.790 2873.980 2539.110 ;
        RECT 2889.820 2538.790 2890.080 2539.110 ;
        RECT 2889.880 2531.630 2890.020 2538.790 ;
        RECT 2889.820 2531.310 2890.080 2531.630 ;
        RECT 2901.320 2531.310 2901.580 2531.630 ;
        RECT 2901.380 2493.405 2901.520 2531.310 ;
        RECT 2901.310 2493.035 2901.590 2493.405 ;
        RECT 288.060 2169.890 288.320 2170.210 ;
        RECT 300.480 2169.890 300.740 2170.210 ;
        RECT 288.120 1841.965 288.260 2169.890 ;
        RECT 288.050 1841.595 288.330 1841.965 ;
      LAYER via2 ;
        RECT 2901.310 2493.080 2901.590 2493.360 ;
        RECT 288.050 1841.640 288.330 1841.920 ;
      LAYER met3 ;
        RECT 2901.285 2493.370 2901.615 2493.385 ;
        RECT 2917.600 2493.370 2924.800 2493.820 ;
        RECT 2901.285 2493.070 2924.800 2493.370 ;
        RECT 2901.285 2493.055 2901.615 2493.070 ;
        RECT 2917.600 2492.620 2924.800 2493.070 ;
        RECT 288.025 1841.930 288.355 1841.945 ;
        RECT 300.000 1841.930 304.000 1842.000 ;
        RECT 288.025 1841.630 304.000 1841.930 ;
        RECT 288.025 1841.615 288.355 1841.630 ;
        RECT 300.000 1841.400 304.000 1841.630 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 286.650 2725.680 286.970 2725.740 ;
        RECT 2900.830 2725.680 2901.150 2725.740 ;
        RECT 286.650 2725.540 2901.150 2725.680 ;
        RECT 286.650 2725.480 286.970 2725.540 ;
        RECT 2900.830 2725.480 2901.150 2725.540 ;
      LAYER via ;
        RECT 286.680 2725.480 286.940 2725.740 ;
        RECT 2900.860 2725.480 2901.120 2725.740 ;
      LAYER met2 ;
        RECT 2900.850 2727.635 2901.130 2728.005 ;
        RECT 2900.920 2725.770 2901.060 2727.635 ;
        RECT 286.680 2725.450 286.940 2725.770 ;
        RECT 2900.860 2725.450 2901.120 2725.770 ;
        RECT 286.740 1873.245 286.880 2725.450 ;
        RECT 286.670 1872.875 286.950 1873.245 ;
      LAYER via2 ;
        RECT 2900.850 2727.680 2901.130 2727.960 ;
        RECT 286.670 1872.920 286.950 1873.200 ;
      LAYER met3 ;
        RECT 2900.825 2727.970 2901.155 2727.985 ;
        RECT 2917.600 2727.970 2924.800 2728.420 ;
        RECT 2900.825 2727.670 2924.800 2727.970 ;
        RECT 2900.825 2727.655 2901.155 2727.670 ;
        RECT 2917.600 2727.220 2924.800 2727.670 ;
        RECT 286.645 1873.210 286.975 1873.225 ;
        RECT 300.000 1873.210 304.000 1873.280 ;
        RECT 286.645 1872.910 304.000 1873.210 ;
        RECT 286.645 1872.895 286.975 1872.910 ;
        RECT 300.000 1872.680 304.000 1872.910 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 285.270 2694.400 285.590 2694.460 ;
        RECT 2902.670 2694.400 2902.990 2694.460 ;
        RECT 285.270 2694.260 2902.990 2694.400 ;
        RECT 285.270 2694.200 285.590 2694.260 ;
        RECT 2902.670 2694.200 2902.990 2694.260 ;
      LAYER via ;
        RECT 285.300 2694.200 285.560 2694.460 ;
        RECT 2902.700 2694.200 2902.960 2694.460 ;
      LAYER met2 ;
        RECT 2902.690 2962.235 2902.970 2962.605 ;
        RECT 2902.760 2694.490 2902.900 2962.235 ;
        RECT 285.300 2694.170 285.560 2694.490 ;
        RECT 2902.700 2694.170 2902.960 2694.490 ;
        RECT 285.360 1905.205 285.500 2694.170 ;
        RECT 285.290 1904.835 285.570 1905.205 ;
      LAYER via2 ;
        RECT 2902.690 2962.280 2902.970 2962.560 ;
        RECT 285.290 1904.880 285.570 1905.160 ;
      LAYER met3 ;
        RECT 2902.665 2962.570 2902.995 2962.585 ;
        RECT 2917.600 2962.570 2924.800 2963.020 ;
        RECT 2902.665 2962.270 2924.800 2962.570 ;
        RECT 2902.665 2962.255 2902.995 2962.270 ;
        RECT 2917.600 2961.820 2924.800 2962.270 ;
        RECT 285.265 1905.170 285.595 1905.185 ;
        RECT 300.000 1905.170 304.000 1905.240 ;
        RECT 285.265 1904.870 304.000 1905.170 ;
        RECT 285.265 1904.855 285.595 1904.870 ;
        RECT 300.000 1904.640 304.000 1904.870 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2901.310 3196.835 2901.590 3197.205 ;
        RECT 2901.380 2696.045 2901.520 3196.835 ;
        RECT 2901.310 2695.675 2901.590 2696.045 ;
      LAYER via2 ;
        RECT 2901.310 3196.880 2901.590 3197.160 ;
        RECT 2901.310 2695.720 2901.590 2696.000 ;
      LAYER met3 ;
        RECT 2901.285 3197.170 2901.615 3197.185 ;
        RECT 2917.600 3197.170 2924.800 3197.620 ;
        RECT 2901.285 3196.870 2924.800 3197.170 ;
        RECT 2901.285 3196.855 2901.615 3196.870 ;
        RECT 2917.600 3196.420 2924.800 3196.870 ;
        RECT 287.310 2696.010 287.690 2696.020 ;
        RECT 2901.285 2696.010 2901.615 2696.025 ;
        RECT 287.310 2695.710 2901.615 2696.010 ;
        RECT 287.310 2695.700 287.690 2695.710 ;
        RECT 2901.285 2695.695 2901.615 2695.710 ;
        RECT 287.310 1936.450 287.690 1936.460 ;
        RECT 300.000 1936.450 304.000 1936.520 ;
        RECT 287.310 1936.150 304.000 1936.450 ;
        RECT 287.310 1936.140 287.690 1936.150 ;
        RECT 300.000 1935.920 304.000 1936.150 ;
      LAYER via3 ;
        RECT 287.340 2695.700 287.660 2696.020 ;
        RECT 287.340 1936.140 287.660 1936.460 ;
      LAYER met4 ;
        RECT 287.335 2695.695 287.665 2696.025 ;
        RECT 287.350 1936.465 287.650 2695.695 ;
        RECT 287.335 1936.135 287.665 1936.465 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 869.470 3431.520 869.790 3431.580 ;
        RECT 893.850 3431.520 894.170 3431.580 ;
        RECT 869.470 3431.380 894.170 3431.520 ;
        RECT 869.470 3431.320 869.790 3431.380 ;
        RECT 893.850 3431.320 894.170 3431.380 ;
        RECT 1835.470 3431.520 1835.790 3431.580 ;
        RECT 1859.850 3431.520 1860.170 3431.580 ;
        RECT 1835.470 3431.380 1860.170 3431.520 ;
        RECT 1835.470 3431.320 1835.790 3431.380 ;
        RECT 1859.850 3431.320 1860.170 3431.380 ;
        RECT 2801.470 3431.520 2801.790 3431.580 ;
        RECT 2825.850 3431.520 2826.170 3431.580 ;
        RECT 2801.470 3431.380 2826.170 3431.520 ;
        RECT 2801.470 3431.320 2801.790 3431.380 ;
        RECT 2825.850 3431.320 2826.170 3431.380 ;
        RECT 772.870 3430.840 773.190 3430.900 ;
        RECT 811.050 3430.840 811.370 3430.900 ;
        RECT 772.870 3430.700 811.370 3430.840 ;
        RECT 772.870 3430.640 773.190 3430.700 ;
        RECT 811.050 3430.640 811.370 3430.700 ;
        RECT 1449.070 3430.840 1449.390 3430.900 ;
        RECT 1472.530 3430.840 1472.850 3430.900 ;
        RECT 1449.070 3430.700 1472.850 3430.840 ;
        RECT 1449.070 3430.640 1449.390 3430.700 ;
        RECT 1472.530 3430.640 1472.850 3430.700 ;
        RECT 1738.870 3430.840 1739.190 3430.900 ;
        RECT 1777.050 3430.840 1777.370 3430.900 ;
        RECT 1738.870 3430.700 1777.370 3430.840 ;
        RECT 1738.870 3430.640 1739.190 3430.700 ;
        RECT 1777.050 3430.640 1777.370 3430.700 ;
        RECT 2704.870 3430.840 2705.190 3430.900 ;
        RECT 2743.050 3430.840 2743.370 3430.900 ;
        RECT 2704.870 3430.700 2743.370 3430.840 ;
        RECT 2704.870 3430.640 2705.190 3430.700 ;
        RECT 2743.050 3430.640 2743.370 3430.700 ;
      LAYER via ;
        RECT 869.500 3431.320 869.760 3431.580 ;
        RECT 893.880 3431.320 894.140 3431.580 ;
        RECT 1835.500 3431.320 1835.760 3431.580 ;
        RECT 1859.880 3431.320 1860.140 3431.580 ;
        RECT 2801.500 3431.320 2801.760 3431.580 ;
        RECT 2825.880 3431.320 2826.140 3431.580 ;
        RECT 772.900 3430.640 773.160 3430.900 ;
        RECT 811.080 3430.640 811.340 3430.900 ;
        RECT 1449.100 3430.640 1449.360 3430.900 ;
        RECT 1472.560 3430.640 1472.820 3430.900 ;
        RECT 1738.900 3430.640 1739.160 3430.900 ;
        RECT 1777.080 3430.640 1777.340 3430.900 ;
        RECT 2704.900 3430.640 2705.160 3430.900 ;
        RECT 2743.080 3430.640 2743.340 3430.900 ;
      LAYER met2 ;
        RECT 941.710 3432.115 941.990 3432.485 ;
        RECT 1897.590 3432.115 1897.870 3432.485 ;
        RECT 2207.630 3432.115 2207.910 3432.485 ;
        RECT 834.530 3431.690 834.810 3431.805 ;
        RECT 835.450 3431.690 835.730 3431.805 ;
        RECT 834.530 3431.550 835.730 3431.690 ;
        RECT 834.530 3431.435 834.810 3431.550 ;
        RECT 835.450 3431.435 835.730 3431.550 ;
        RECT 869.490 3431.435 869.770 3431.805 ;
        RECT 869.500 3431.290 869.760 3431.435 ;
        RECT 893.880 3431.290 894.140 3431.610 ;
        RECT 893.940 3431.125 894.080 3431.290 ;
        RECT 941.780 3431.125 941.920 3432.115 ;
        RECT 1800.530 3431.690 1800.810 3431.805 ;
        RECT 1801.450 3431.690 1801.730 3431.805 ;
        RECT 1800.530 3431.550 1801.730 3431.690 ;
        RECT 1800.530 3431.435 1800.810 3431.550 ;
        RECT 1801.450 3431.435 1801.730 3431.550 ;
        RECT 1835.490 3431.435 1835.770 3431.805 ;
        RECT 1835.500 3431.290 1835.760 3431.435 ;
        RECT 1859.880 3431.290 1860.140 3431.610 ;
        RECT 1859.940 3431.125 1860.080 3431.290 ;
        RECT 1897.660 3431.125 1897.800 3432.115 ;
        RECT 2207.700 3431.125 2207.840 3432.115 ;
        RECT 2766.530 3431.690 2766.810 3431.805 ;
        RECT 2767.450 3431.690 2767.730 3431.805 ;
        RECT 2766.530 3431.550 2767.730 3431.690 ;
        RECT 2766.530 3431.435 2766.810 3431.550 ;
        RECT 2767.450 3431.435 2767.730 3431.550 ;
        RECT 2801.490 3431.435 2801.770 3431.805 ;
        RECT 2801.500 3431.290 2801.760 3431.435 ;
        RECT 2825.880 3431.290 2826.140 3431.610 ;
        RECT 2825.940 3431.125 2826.080 3431.290 ;
        RECT 772.890 3430.755 773.170 3431.125 ;
        RECT 772.900 3430.610 773.160 3430.755 ;
        RECT 811.080 3430.610 811.340 3430.930 ;
        RECT 893.870 3430.755 894.150 3431.125 ;
        RECT 941.710 3430.755 941.990 3431.125 ;
        RECT 1449.090 3430.755 1449.370 3431.125 ;
        RECT 1449.100 3430.610 1449.360 3430.755 ;
        RECT 1472.560 3430.610 1472.820 3430.930 ;
        RECT 1738.890 3430.755 1739.170 3431.125 ;
        RECT 1738.900 3430.610 1739.160 3430.755 ;
        RECT 1777.080 3430.610 1777.340 3430.930 ;
        RECT 1859.870 3430.755 1860.150 3431.125 ;
        RECT 1897.590 3430.755 1897.870 3431.125 ;
        RECT 2137.710 3431.010 2137.990 3431.125 ;
        RECT 2138.630 3431.010 2138.910 3431.125 ;
        RECT 2137.710 3430.870 2138.910 3431.010 ;
        RECT 2137.710 3430.755 2137.990 3430.870 ;
        RECT 2138.630 3430.755 2138.910 3430.870 ;
        RECT 2207.630 3430.755 2207.910 3431.125 ;
        RECT 2704.890 3430.755 2705.170 3431.125 ;
        RECT 2704.900 3430.610 2705.160 3430.755 ;
        RECT 2743.080 3430.610 2743.340 3430.930 ;
        RECT 2825.870 3430.755 2826.150 3431.125 ;
        RECT 2863.590 3431.010 2863.870 3431.125 ;
        RECT 2863.200 3430.870 2863.870 3431.010 ;
        RECT 811.140 3429.765 811.280 3430.610 ;
        RECT 1472.620 3429.765 1472.760 3430.610 ;
        RECT 1777.140 3429.765 1777.280 3430.610 ;
        RECT 2743.140 3429.765 2743.280 3430.610 ;
        RECT 2863.200 3430.445 2863.340 3430.870 ;
        RECT 2863.590 3430.755 2863.870 3430.870 ;
        RECT 2863.130 3430.075 2863.410 3430.445 ;
        RECT 811.070 3429.395 811.350 3429.765 ;
        RECT 1472.550 3429.395 1472.830 3429.765 ;
        RECT 1777.070 3429.395 1777.350 3429.765 ;
        RECT 2743.070 3429.395 2743.350 3429.765 ;
      LAYER via2 ;
        RECT 941.710 3432.160 941.990 3432.440 ;
        RECT 1897.590 3432.160 1897.870 3432.440 ;
        RECT 2207.630 3432.160 2207.910 3432.440 ;
        RECT 834.530 3431.480 834.810 3431.760 ;
        RECT 835.450 3431.480 835.730 3431.760 ;
        RECT 869.490 3431.480 869.770 3431.760 ;
        RECT 1800.530 3431.480 1800.810 3431.760 ;
        RECT 1801.450 3431.480 1801.730 3431.760 ;
        RECT 1835.490 3431.480 1835.770 3431.760 ;
        RECT 2766.530 3431.480 2766.810 3431.760 ;
        RECT 2767.450 3431.480 2767.730 3431.760 ;
        RECT 2801.490 3431.480 2801.770 3431.760 ;
        RECT 772.890 3430.800 773.170 3431.080 ;
        RECT 893.870 3430.800 894.150 3431.080 ;
        RECT 941.710 3430.800 941.990 3431.080 ;
        RECT 1449.090 3430.800 1449.370 3431.080 ;
        RECT 1738.890 3430.800 1739.170 3431.080 ;
        RECT 1859.870 3430.800 1860.150 3431.080 ;
        RECT 1897.590 3430.800 1897.870 3431.080 ;
        RECT 2137.710 3430.800 2137.990 3431.080 ;
        RECT 2138.630 3430.800 2138.910 3431.080 ;
        RECT 2207.630 3430.800 2207.910 3431.080 ;
        RECT 2704.890 3430.800 2705.170 3431.080 ;
        RECT 2825.870 3430.800 2826.150 3431.080 ;
        RECT 2863.590 3430.800 2863.870 3431.080 ;
        RECT 2863.130 3430.120 2863.410 3430.400 ;
        RECT 811.070 3429.440 811.350 3429.720 ;
        RECT 1472.550 3429.440 1472.830 3429.720 ;
        RECT 1777.070 3429.440 1777.350 3429.720 ;
        RECT 2743.070 3429.440 2743.350 3429.720 ;
      LAYER met3 ;
        RECT 917.510 3432.450 917.890 3432.460 ;
        RECT 941.685 3432.450 942.015 3432.465 ;
        RECT 917.510 3432.150 942.015 3432.450 ;
        RECT 917.510 3432.140 917.890 3432.150 ;
        RECT 941.685 3432.135 942.015 3432.150 ;
        RECT 1883.510 3432.450 1883.890 3432.460 ;
        RECT 1897.565 3432.450 1897.895 3432.465 ;
        RECT 1883.510 3432.150 1897.895 3432.450 ;
        RECT 1883.510 3432.140 1883.890 3432.150 ;
        RECT 1897.565 3432.135 1897.895 3432.150 ;
        RECT 2173.310 3432.450 2173.690 3432.460 ;
        RECT 2207.605 3432.450 2207.935 3432.465 ;
        RECT 2173.310 3432.150 2207.935 3432.450 ;
        RECT 2173.310 3432.140 2173.690 3432.150 ;
        RECT 2207.605 3432.135 2207.935 3432.150 ;
        RECT 820.910 3431.770 821.290 3431.780 ;
        RECT 834.505 3431.770 834.835 3431.785 ;
        RECT 820.910 3431.470 834.835 3431.770 ;
        RECT 820.910 3431.460 821.290 3431.470 ;
        RECT 834.505 3431.455 834.835 3431.470 ;
        RECT 835.425 3431.770 835.755 3431.785 ;
        RECT 869.465 3431.770 869.795 3431.785 ;
        RECT 835.425 3431.470 869.795 3431.770 ;
        RECT 835.425 3431.455 835.755 3431.470 ;
        RECT 869.465 3431.455 869.795 3431.470 ;
        RECT 1786.910 3431.770 1787.290 3431.780 ;
        RECT 1800.505 3431.770 1800.835 3431.785 ;
        RECT 1786.910 3431.470 1800.835 3431.770 ;
        RECT 1786.910 3431.460 1787.290 3431.470 ;
        RECT 1800.505 3431.455 1800.835 3431.470 ;
        RECT 1801.425 3431.770 1801.755 3431.785 ;
        RECT 1835.465 3431.770 1835.795 3431.785 ;
        RECT 1801.425 3431.470 1835.795 3431.770 ;
        RECT 1801.425 3431.455 1801.755 3431.470 ;
        RECT 1835.465 3431.455 1835.795 3431.470 ;
        RECT 2752.910 3431.770 2753.290 3431.780 ;
        RECT 2766.505 3431.770 2766.835 3431.785 ;
        RECT 2752.910 3431.470 2766.835 3431.770 ;
        RECT 2752.910 3431.460 2753.290 3431.470 ;
        RECT 2766.505 3431.455 2766.835 3431.470 ;
        RECT 2767.425 3431.770 2767.755 3431.785 ;
        RECT 2801.465 3431.770 2801.795 3431.785 ;
        RECT 2917.600 3431.770 2924.800 3432.220 ;
        RECT 2767.425 3431.470 2801.795 3431.770 ;
        RECT 2767.425 3431.455 2767.755 3431.470 ;
        RECT 2801.465 3431.455 2801.795 3431.470 ;
        RECT 2916.710 3431.470 2924.800 3431.770 ;
        RECT 289.150 3431.090 289.530 3431.100 ;
        RECT 772.865 3431.090 773.195 3431.105 ;
        RECT 289.150 3430.790 324.450 3431.090 ;
        RECT 289.150 3430.780 289.530 3430.790 ;
        RECT 324.150 3430.410 324.450 3430.790 ;
        RECT 372.910 3430.790 421.050 3431.090 ;
        RECT 324.150 3430.110 372.290 3430.410 ;
        RECT 371.990 3429.730 372.290 3430.110 ;
        RECT 372.910 3429.730 373.210 3430.790 ;
        RECT 420.750 3430.410 421.050 3430.790 ;
        RECT 469.510 3430.790 517.650 3431.090 ;
        RECT 420.750 3430.110 468.890 3430.410 ;
        RECT 371.990 3429.430 373.210 3429.730 ;
        RECT 468.590 3429.730 468.890 3430.110 ;
        RECT 469.510 3429.730 469.810 3430.790 ;
        RECT 517.350 3430.410 517.650 3430.790 ;
        RECT 566.110 3430.790 614.250 3431.090 ;
        RECT 517.350 3430.110 565.490 3430.410 ;
        RECT 468.590 3429.430 469.810 3429.730 ;
        RECT 565.190 3429.730 565.490 3430.110 ;
        RECT 566.110 3429.730 566.410 3430.790 ;
        RECT 613.950 3430.410 614.250 3430.790 ;
        RECT 662.710 3430.790 710.850 3431.090 ;
        RECT 613.950 3430.110 662.090 3430.410 ;
        RECT 565.190 3429.430 566.410 3429.730 ;
        RECT 661.790 3429.730 662.090 3430.110 ;
        RECT 662.710 3429.730 663.010 3430.790 ;
        RECT 710.550 3430.410 710.850 3430.790 ;
        RECT 759.310 3430.790 773.195 3431.090 ;
        RECT 710.550 3430.110 758.690 3430.410 ;
        RECT 661.790 3429.430 663.010 3429.730 ;
        RECT 758.390 3429.730 758.690 3430.110 ;
        RECT 759.310 3429.730 759.610 3430.790 ;
        RECT 772.865 3430.775 773.195 3430.790 ;
        RECT 893.845 3431.090 894.175 3431.105 ;
        RECT 917.510 3431.090 917.890 3431.100 ;
        RECT 893.845 3430.790 917.890 3431.090 ;
        RECT 893.845 3430.775 894.175 3430.790 ;
        RECT 917.510 3430.780 917.890 3430.790 ;
        RECT 941.685 3431.090 942.015 3431.105 ;
        RECT 1449.065 3431.090 1449.395 3431.105 ;
        RECT 941.685 3430.790 1000.650 3431.090 ;
        RECT 941.685 3430.775 942.015 3430.790 ;
        RECT 1000.350 3430.410 1000.650 3430.790 ;
        RECT 1049.110 3430.790 1097.250 3431.090 ;
        RECT 1000.350 3430.110 1048.490 3430.410 ;
        RECT 758.390 3429.430 759.610 3429.730 ;
        RECT 811.045 3429.730 811.375 3429.745 ;
        RECT 820.910 3429.730 821.290 3429.740 ;
        RECT 811.045 3429.430 821.290 3429.730 ;
        RECT 1048.190 3429.730 1048.490 3430.110 ;
        RECT 1049.110 3429.730 1049.410 3430.790 ;
        RECT 1096.950 3430.410 1097.250 3430.790 ;
        RECT 1145.710 3430.790 1193.850 3431.090 ;
        RECT 1096.950 3430.110 1145.090 3430.410 ;
        RECT 1048.190 3429.430 1049.410 3429.730 ;
        RECT 1144.790 3429.730 1145.090 3430.110 ;
        RECT 1145.710 3429.730 1146.010 3430.790 ;
        RECT 1193.550 3430.410 1193.850 3430.790 ;
        RECT 1242.310 3430.790 1290.450 3431.090 ;
        RECT 1193.550 3430.110 1241.690 3430.410 ;
        RECT 1144.790 3429.430 1146.010 3429.730 ;
        RECT 1241.390 3429.730 1241.690 3430.110 ;
        RECT 1242.310 3429.730 1242.610 3430.790 ;
        RECT 1290.150 3430.410 1290.450 3430.790 ;
        RECT 1338.910 3430.790 1387.050 3431.090 ;
        RECT 1290.150 3430.110 1338.290 3430.410 ;
        RECT 1241.390 3429.430 1242.610 3429.730 ;
        RECT 1337.990 3429.730 1338.290 3430.110 ;
        RECT 1338.910 3429.730 1339.210 3430.790 ;
        RECT 1386.750 3430.410 1387.050 3430.790 ;
        RECT 1435.510 3430.790 1449.395 3431.090 ;
        RECT 1386.750 3430.110 1434.890 3430.410 ;
        RECT 1337.990 3429.430 1339.210 3429.730 ;
        RECT 1434.590 3429.730 1434.890 3430.110 ;
        RECT 1435.510 3429.730 1435.810 3430.790 ;
        RECT 1449.065 3430.775 1449.395 3430.790 ;
        RECT 1497.110 3431.090 1497.490 3431.100 ;
        RECT 1738.865 3431.090 1739.195 3431.105 ;
        RECT 1497.110 3430.790 1580.250 3431.090 ;
        RECT 1497.110 3430.780 1497.490 3430.790 ;
        RECT 1579.950 3430.410 1580.250 3430.790 ;
        RECT 1628.710 3430.790 1676.850 3431.090 ;
        RECT 1579.950 3430.110 1628.090 3430.410 ;
        RECT 1434.590 3429.430 1435.810 3429.730 ;
        RECT 1472.525 3429.730 1472.855 3429.745 ;
        RECT 1497.110 3429.730 1497.490 3429.740 ;
        RECT 1472.525 3429.430 1497.490 3429.730 ;
        RECT 1627.790 3429.730 1628.090 3430.110 ;
        RECT 1628.710 3429.730 1629.010 3430.790 ;
        RECT 1676.550 3430.410 1676.850 3430.790 ;
        RECT 1725.310 3430.790 1739.195 3431.090 ;
        RECT 1676.550 3430.110 1724.690 3430.410 ;
        RECT 1627.790 3429.430 1629.010 3429.730 ;
        RECT 1724.390 3429.730 1724.690 3430.110 ;
        RECT 1725.310 3429.730 1725.610 3430.790 ;
        RECT 1738.865 3430.775 1739.195 3430.790 ;
        RECT 1859.845 3431.090 1860.175 3431.105 ;
        RECT 1883.510 3431.090 1883.890 3431.100 ;
        RECT 1859.845 3430.790 1883.890 3431.090 ;
        RECT 1859.845 3430.775 1860.175 3430.790 ;
        RECT 1883.510 3430.780 1883.890 3430.790 ;
        RECT 1897.565 3431.090 1897.895 3431.105 ;
        RECT 2137.685 3431.090 2138.015 3431.105 ;
        RECT 1897.565 3430.790 1966.650 3431.090 ;
        RECT 1897.565 3430.775 1897.895 3430.790 ;
        RECT 1966.350 3430.410 1966.650 3430.790 ;
        RECT 2015.110 3430.790 2138.015 3431.090 ;
        RECT 1966.350 3430.110 2014.490 3430.410 ;
        RECT 1724.390 3429.430 1725.610 3429.730 ;
        RECT 1777.045 3429.730 1777.375 3429.745 ;
        RECT 1786.910 3429.730 1787.290 3429.740 ;
        RECT 1777.045 3429.430 1787.290 3429.730 ;
        RECT 2014.190 3429.730 2014.490 3430.110 ;
        RECT 2015.110 3429.730 2015.410 3430.790 ;
        RECT 2137.685 3430.775 2138.015 3430.790 ;
        RECT 2138.605 3431.090 2138.935 3431.105 ;
        RECT 2207.605 3431.090 2207.935 3431.105 ;
        RECT 2704.865 3431.090 2705.195 3431.105 ;
        RECT 2138.605 3430.790 2148.810 3431.090 ;
        RECT 2138.605 3430.775 2138.935 3430.790 ;
        RECT 2148.510 3430.410 2148.810 3430.790 ;
        RECT 2207.605 3430.790 2256.450 3431.090 ;
        RECT 2207.605 3430.775 2207.935 3430.790 ;
        RECT 2173.310 3430.410 2173.690 3430.420 ;
        RECT 2148.510 3430.110 2173.690 3430.410 ;
        RECT 2256.150 3430.410 2256.450 3430.790 ;
        RECT 2304.910 3430.790 2353.050 3431.090 ;
        RECT 2256.150 3430.110 2304.290 3430.410 ;
        RECT 2173.310 3430.100 2173.690 3430.110 ;
        RECT 2014.190 3429.430 2015.410 3429.730 ;
        RECT 2303.990 3429.730 2304.290 3430.110 ;
        RECT 2304.910 3429.730 2305.210 3430.790 ;
        RECT 2352.750 3430.410 2353.050 3430.790 ;
        RECT 2401.510 3430.790 2449.650 3431.090 ;
        RECT 2352.750 3430.110 2400.890 3430.410 ;
        RECT 2303.990 3429.430 2305.210 3429.730 ;
        RECT 2400.590 3429.730 2400.890 3430.110 ;
        RECT 2401.510 3429.730 2401.810 3430.790 ;
        RECT 2449.350 3430.410 2449.650 3430.790 ;
        RECT 2498.110 3430.790 2546.250 3431.090 ;
        RECT 2449.350 3430.110 2497.490 3430.410 ;
        RECT 2400.590 3429.430 2401.810 3429.730 ;
        RECT 2497.190 3429.730 2497.490 3430.110 ;
        RECT 2498.110 3429.730 2498.410 3430.790 ;
        RECT 2545.950 3430.410 2546.250 3430.790 ;
        RECT 2594.710 3430.790 2642.850 3431.090 ;
        RECT 2545.950 3430.110 2594.090 3430.410 ;
        RECT 2497.190 3429.430 2498.410 3429.730 ;
        RECT 2593.790 3429.730 2594.090 3430.110 ;
        RECT 2594.710 3429.730 2595.010 3430.790 ;
        RECT 2642.550 3430.410 2642.850 3430.790 ;
        RECT 2691.310 3430.790 2705.195 3431.090 ;
        RECT 2642.550 3430.110 2690.690 3430.410 ;
        RECT 2593.790 3429.430 2595.010 3429.730 ;
        RECT 2690.390 3429.730 2690.690 3430.110 ;
        RECT 2691.310 3429.730 2691.610 3430.790 ;
        RECT 2704.865 3430.775 2705.195 3430.790 ;
        RECT 2825.845 3431.090 2826.175 3431.105 ;
        RECT 2863.565 3431.090 2863.895 3431.105 ;
        RECT 2825.845 3430.790 2849.850 3431.090 ;
        RECT 2825.845 3430.775 2826.175 3430.790 ;
        RECT 2849.550 3430.410 2849.850 3430.790 ;
        RECT 2863.565 3430.790 2884.810 3431.090 ;
        RECT 2863.565 3430.775 2863.895 3430.790 ;
        RECT 2863.105 3430.410 2863.435 3430.425 ;
        RECT 2849.550 3430.110 2863.435 3430.410 ;
        RECT 2884.510 3430.410 2884.810 3430.790 ;
        RECT 2916.710 3430.410 2917.010 3431.470 ;
        RECT 2917.600 3431.020 2924.800 3431.470 ;
        RECT 2884.510 3430.110 2917.010 3430.410 ;
        RECT 2863.105 3430.095 2863.435 3430.110 ;
        RECT 2690.390 3429.430 2691.610 3429.730 ;
        RECT 2743.045 3429.730 2743.375 3429.745 ;
        RECT 2752.910 3429.730 2753.290 3429.740 ;
        RECT 2743.045 3429.430 2753.290 3429.730 ;
        RECT 811.045 3429.415 811.375 3429.430 ;
        RECT 820.910 3429.420 821.290 3429.430 ;
        RECT 1472.525 3429.415 1472.855 3429.430 ;
        RECT 1497.110 3429.420 1497.490 3429.430 ;
        RECT 1777.045 3429.415 1777.375 3429.430 ;
        RECT 1786.910 3429.420 1787.290 3429.430 ;
        RECT 2743.045 3429.415 2743.375 3429.430 ;
        RECT 2752.910 3429.420 2753.290 3429.430 ;
        RECT 289.150 1968.410 289.530 1968.420 ;
        RECT 300.000 1968.410 304.000 1968.480 ;
        RECT 289.150 1968.110 304.000 1968.410 ;
        RECT 289.150 1968.100 289.530 1968.110 ;
        RECT 300.000 1967.880 304.000 1968.110 ;
      LAYER via3 ;
        RECT 917.540 3432.140 917.860 3432.460 ;
        RECT 1883.540 3432.140 1883.860 3432.460 ;
        RECT 2173.340 3432.140 2173.660 3432.460 ;
        RECT 820.940 3431.460 821.260 3431.780 ;
        RECT 1786.940 3431.460 1787.260 3431.780 ;
        RECT 2752.940 3431.460 2753.260 3431.780 ;
        RECT 289.180 3430.780 289.500 3431.100 ;
        RECT 917.540 3430.780 917.860 3431.100 ;
        RECT 820.940 3429.420 821.260 3429.740 ;
        RECT 1497.140 3430.780 1497.460 3431.100 ;
        RECT 1497.140 3429.420 1497.460 3429.740 ;
        RECT 1883.540 3430.780 1883.860 3431.100 ;
        RECT 1786.940 3429.420 1787.260 3429.740 ;
        RECT 2173.340 3430.100 2173.660 3430.420 ;
        RECT 2752.940 3429.420 2753.260 3429.740 ;
        RECT 289.180 1968.100 289.500 1968.420 ;
      LAYER met4 ;
        RECT 917.535 3432.135 917.865 3432.465 ;
        RECT 1883.535 3432.135 1883.865 3432.465 ;
        RECT 2173.335 3432.135 2173.665 3432.465 ;
        RECT 820.935 3431.455 821.265 3431.785 ;
        RECT 289.175 3430.775 289.505 3431.105 ;
        RECT 289.190 1968.425 289.490 3430.775 ;
        RECT 820.950 3429.745 821.250 3431.455 ;
        RECT 917.550 3431.105 917.850 3432.135 ;
        RECT 1786.935 3431.455 1787.265 3431.785 ;
        RECT 917.535 3430.775 917.865 3431.105 ;
        RECT 1497.135 3430.775 1497.465 3431.105 ;
        RECT 1497.150 3429.745 1497.450 3430.775 ;
        RECT 1786.950 3429.745 1787.250 3431.455 ;
        RECT 1883.550 3431.105 1883.850 3432.135 ;
        RECT 1883.535 3430.775 1883.865 3431.105 ;
        RECT 2173.350 3430.425 2173.650 3432.135 ;
        RECT 2752.935 3431.455 2753.265 3431.785 ;
        RECT 2173.335 3430.095 2173.665 3430.425 ;
        RECT 2752.950 3429.745 2753.250 3431.455 ;
        RECT 820.935 3429.415 821.265 3429.745 ;
        RECT 1497.135 3429.415 1497.465 3429.745 ;
        RECT 1786.935 3429.415 1787.265 3429.745 ;
        RECT 2752.935 3429.415 2753.265 3429.745 ;
        RECT 289.175 1968.095 289.505 1968.425 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 296.770 3501.560 297.090 3501.620 ;
        RECT 2717.290 3501.560 2717.610 3501.620 ;
        RECT 296.770 3501.420 2717.610 3501.560 ;
        RECT 296.770 3501.360 297.090 3501.420 ;
        RECT 2717.290 3501.360 2717.610 3501.420 ;
      LAYER via ;
        RECT 296.800 3501.360 297.060 3501.620 ;
        RECT 2717.320 3501.360 2717.580 3501.620 ;
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
        RECT 2717.380 3501.650 2717.520 3517.600 ;
        RECT 296.800 3501.330 297.060 3501.650 ;
        RECT 2717.320 3501.330 2717.580 3501.650 ;
        RECT 296.860 1999.725 297.000 3501.330 ;
        RECT 296.790 1999.355 297.070 1999.725 ;
      LAYER via2 ;
        RECT 296.790 1999.400 297.070 1999.680 ;
      LAYER met3 ;
        RECT 296.765 1999.690 297.095 1999.705 ;
        RECT 300.000 1999.690 304.000 1999.760 ;
        RECT 296.765 1999.390 304.000 1999.690 ;
        RECT 296.765 1999.375 297.095 1999.390 ;
        RECT 300.000 1999.160 304.000 1999.390 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 289.410 3502.240 289.730 3502.300 ;
        RECT 2392.530 3502.240 2392.850 3502.300 ;
        RECT 289.410 3502.100 2392.850 3502.240 ;
        RECT 289.410 3502.040 289.730 3502.100 ;
        RECT 2392.530 3502.040 2392.850 3502.100 ;
      LAYER via ;
        RECT 289.440 3502.040 289.700 3502.300 ;
        RECT 2392.560 3502.040 2392.820 3502.300 ;
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
        RECT 2392.620 3502.330 2392.760 3517.600 ;
        RECT 289.440 3502.010 289.700 3502.330 ;
        RECT 2392.560 3502.010 2392.820 3502.330 ;
        RECT 289.500 2031.685 289.640 3502.010 ;
        RECT 289.430 2031.315 289.710 2031.685 ;
      LAYER via2 ;
        RECT 289.430 2031.360 289.710 2031.640 ;
      LAYER met3 ;
        RECT 289.405 2031.650 289.735 2031.665 ;
        RECT 300.000 2031.650 304.000 2031.720 ;
        RECT 289.405 2031.350 304.000 2031.650 ;
        RECT 289.405 2031.335 289.735 2031.350 ;
        RECT 300.000 2031.120 304.000 2031.350 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 288.950 3502.580 289.270 3502.640 ;
        RECT 2068.230 3502.580 2068.550 3502.640 ;
        RECT 288.950 3502.440 2068.550 3502.580 ;
        RECT 288.950 3502.380 289.270 3502.440 ;
        RECT 2068.230 3502.380 2068.550 3502.440 ;
      LAYER via ;
        RECT 288.980 3502.380 289.240 3502.640 ;
        RECT 2068.260 3502.380 2068.520 3502.640 ;
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
        RECT 2068.320 3502.670 2068.460 3517.600 ;
        RECT 288.980 3502.350 289.240 3502.670 ;
        RECT 2068.260 3502.350 2068.520 3502.670 ;
        RECT 289.040 2062.965 289.180 3502.350 ;
        RECT 288.970 2062.595 289.250 2062.965 ;
      LAYER via2 ;
        RECT 288.970 2062.640 289.250 2062.920 ;
      LAYER met3 ;
        RECT 288.945 2062.930 289.275 2062.945 ;
        RECT 300.000 2062.930 304.000 2063.000 ;
        RECT 288.945 2062.630 304.000 2062.930 ;
        RECT 288.945 2062.615 289.275 2062.630 ;
        RECT 300.000 2062.400 304.000 2062.630 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 288.490 3503.260 288.810 3503.320 ;
        RECT 1743.930 3503.260 1744.250 3503.320 ;
        RECT 288.490 3503.120 1744.250 3503.260 ;
        RECT 288.490 3503.060 288.810 3503.120 ;
        RECT 1743.930 3503.060 1744.250 3503.120 ;
      LAYER via ;
        RECT 288.520 3503.060 288.780 3503.320 ;
        RECT 1743.960 3503.060 1744.220 3503.320 ;
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
        RECT 1744.020 3503.350 1744.160 3517.600 ;
        RECT 288.520 3503.030 288.780 3503.350 ;
        RECT 1743.960 3503.030 1744.220 3503.350 ;
        RECT 288.580 2094.925 288.720 3503.030 ;
        RECT 288.510 2094.555 288.790 2094.925 ;
      LAYER via2 ;
        RECT 288.510 2094.600 288.790 2094.880 ;
      LAYER met3 ;
        RECT 288.485 2094.890 288.815 2094.905 ;
        RECT 300.000 2094.890 304.000 2094.960 ;
        RECT 288.485 2094.590 304.000 2094.890 ;
        RECT 288.485 2094.575 288.815 2094.590 ;
        RECT 300.000 2094.360 304.000 2094.590 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 294.470 3503.940 294.790 3504.000 ;
        RECT 1419.170 3503.940 1419.490 3504.000 ;
        RECT 294.470 3503.800 1419.490 3503.940 ;
        RECT 294.470 3503.740 294.790 3503.800 ;
        RECT 1419.170 3503.740 1419.490 3503.800 ;
      LAYER via ;
        RECT 294.500 3503.740 294.760 3504.000 ;
        RECT 1419.200 3503.740 1419.460 3504.000 ;
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
        RECT 1419.260 3504.030 1419.400 3517.600 ;
        RECT 294.500 3503.710 294.760 3504.030 ;
        RECT 1419.200 3503.710 1419.460 3504.030 ;
        RECT 294.560 2126.205 294.700 3503.710 ;
        RECT 294.490 2125.835 294.770 2126.205 ;
      LAYER via2 ;
        RECT 294.490 2125.880 294.770 2126.160 ;
      LAYER met3 ;
        RECT 294.465 2126.170 294.795 2126.185 ;
        RECT 300.000 2126.170 304.000 2126.240 ;
        RECT 294.465 2125.870 304.000 2126.170 ;
        RECT 294.465 2125.855 294.795 2125.870 ;
        RECT 300.000 2125.640 304.000 2125.870 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 447.650 380.700 447.970 380.760 ;
        RECT 449.030 380.700 449.350 380.760 ;
        RECT 447.650 380.560 449.350 380.700 ;
        RECT 447.650 380.500 447.970 380.560 ;
        RECT 449.030 380.500 449.350 380.560 ;
        RECT 737.910 380.700 738.230 380.760 ;
        RECT 772.410 380.700 772.730 380.760 ;
        RECT 737.910 380.560 772.730 380.700 ;
        RECT 737.910 380.500 738.230 380.560 ;
        RECT 772.410 380.500 772.730 380.560 ;
        RECT 579.670 380.020 579.990 380.080 ;
        RECT 594.390 380.020 594.710 380.080 ;
        RECT 579.670 379.880 594.710 380.020 ;
        RECT 579.670 379.820 579.990 379.880 ;
        RECT 594.390 379.820 594.710 379.880 ;
      LAYER via ;
        RECT 447.680 380.500 447.940 380.760 ;
        RECT 449.060 380.500 449.320 380.760 ;
        RECT 737.940 380.500 738.200 380.760 ;
        RECT 772.440 380.500 772.700 380.760 ;
        RECT 579.700 379.820 579.960 380.080 ;
        RECT 594.420 379.820 594.680 380.080 ;
      LAYER met2 ;
        RECT 675.830 382.315 676.110 382.685 ;
        RECT 386.030 380.955 386.310 381.325 ;
        RECT 594.410 380.955 594.690 381.325 ;
        RECT 386.100 379.285 386.240 380.955 ;
        RECT 447.680 380.645 447.940 380.790 ;
        RECT 449.060 380.645 449.320 380.790 ;
        RECT 447.670 380.275 447.950 380.645 ;
        RECT 449.050 380.275 449.330 380.645 ;
        RECT 594.480 380.110 594.620 380.955 ;
        RECT 675.900 380.645 676.040 382.315 ;
        RECT 700.210 381.635 700.490 382.005 ;
        RECT 675.830 380.275 676.110 380.645 ;
        RECT 579.700 379.965 579.960 380.110 ;
        RECT 579.690 379.595 579.970 379.965 ;
        RECT 594.420 379.790 594.680 380.110 ;
        RECT 700.280 379.965 700.420 381.635 ;
        RECT 772.430 380.955 772.710 381.325 ;
        RECT 772.500 380.790 772.640 380.955 ;
        RECT 737.940 380.645 738.200 380.790 ;
        RECT 737.930 380.275 738.210 380.645 ;
        RECT 772.440 380.470 772.700 380.790 ;
        RECT 700.210 379.595 700.490 379.965 ;
        RECT 386.030 378.915 386.310 379.285 ;
      LAYER via2 ;
        RECT 675.830 382.360 676.110 382.640 ;
        RECT 386.030 381.000 386.310 381.280 ;
        RECT 594.410 381.000 594.690 381.280 ;
        RECT 447.670 380.320 447.950 380.600 ;
        RECT 449.050 380.320 449.330 380.600 ;
        RECT 700.210 381.680 700.490 381.960 ;
        RECT 675.830 380.320 676.110 380.600 ;
        RECT 579.690 379.640 579.970 379.920 ;
        RECT 772.430 381.000 772.710 381.280 ;
        RECT 737.930 380.320 738.210 380.600 ;
        RECT 700.210 379.640 700.490 379.920 ;
        RECT 386.030 378.960 386.310 379.240 ;
      LAYER met3 ;
        RECT 287.310 1557.690 287.690 1557.700 ;
        RECT 300.000 1557.690 304.000 1557.760 ;
        RECT 287.310 1557.390 304.000 1557.690 ;
        RECT 287.310 1557.380 287.690 1557.390 ;
        RECT 300.000 1557.160 304.000 1557.390 ;
        RECT 627.710 382.650 628.090 382.660 ;
        RECT 675.805 382.650 676.135 382.665 ;
        RECT 627.710 382.350 676.135 382.650 ;
        RECT 627.710 382.340 628.090 382.350 ;
        RECT 675.805 382.335 676.135 382.350 ;
        RECT 578.950 381.970 579.330 381.980 ;
        RECT 700.185 381.970 700.515 381.985 ;
        RECT 544.030 381.670 579.330 381.970 ;
        RECT 287.310 381.290 287.690 381.300 ;
        RECT 386.005 381.290 386.335 381.305 ;
        RECT 287.310 380.990 303.290 381.290 ;
        RECT 287.310 380.980 287.690 380.990 ;
        RECT 302.990 379.930 303.290 380.990 ;
        RECT 386.005 380.990 399.890 381.290 ;
        RECT 386.005 380.975 386.335 380.990 ;
        RECT 337.910 380.610 338.290 380.620 ;
        RECT 303.910 380.310 338.290 380.610 ;
        RECT 303.910 379.930 304.210 380.310 ;
        RECT 337.910 380.300 338.290 380.310 ;
        RECT 302.990 379.630 304.210 379.930 ;
        RECT 399.590 379.930 399.890 380.990 ;
        RECT 447.645 380.610 447.975 380.625 ;
        RECT 400.510 380.310 447.975 380.610 ;
        RECT 400.510 379.930 400.810 380.310 ;
        RECT 447.645 380.295 447.975 380.310 ;
        RECT 449.025 380.610 449.355 380.625 ;
        RECT 544.030 380.610 544.330 381.670 ;
        RECT 578.950 381.660 579.330 381.670 ;
        RECT 676.510 381.670 700.515 381.970 ;
        RECT 594.385 381.290 594.715 381.305 ;
        RECT 627.710 381.290 628.090 381.300 ;
        RECT 594.385 380.990 628.090 381.290 ;
        RECT 594.385 380.975 594.715 380.990 ;
        RECT 627.710 380.980 628.090 380.990 ;
        RECT 449.025 380.310 482.690 380.610 ;
        RECT 449.025 380.295 449.355 380.310 ;
        RECT 399.590 379.630 400.810 379.930 ;
        RECT 482.390 379.930 482.690 380.310 ;
        RECT 497.110 380.310 544.330 380.610 ;
        RECT 675.805 380.610 676.135 380.625 ;
        RECT 676.510 380.610 676.810 381.670 ;
        RECT 700.185 381.655 700.515 381.670 ;
        RECT 772.405 381.290 772.735 381.305 ;
        RECT 2917.600 381.290 2924.800 381.740 ;
        RECT 772.405 380.990 807.450 381.290 ;
        RECT 772.405 380.975 772.735 380.990 ;
        RECT 737.905 380.610 738.235 380.625 ;
        RECT 675.805 380.310 676.810 380.610 ;
        RECT 724.350 380.310 738.235 380.610 ;
        RECT 807.150 380.610 807.450 380.990 ;
        RECT 855.910 380.990 904.050 381.290 ;
        RECT 807.150 380.310 855.290 380.610 ;
        RECT 497.110 379.930 497.410 380.310 ;
        RECT 675.805 380.295 676.135 380.310 ;
        RECT 482.390 379.630 497.410 379.930 ;
        RECT 578.950 379.930 579.330 379.940 ;
        RECT 579.665 379.930 579.995 379.945 ;
        RECT 578.950 379.630 579.995 379.930 ;
        RECT 578.950 379.620 579.330 379.630 ;
        RECT 579.665 379.615 579.995 379.630 ;
        RECT 700.185 379.930 700.515 379.945 ;
        RECT 724.350 379.930 724.650 380.310 ;
        RECT 737.905 380.295 738.235 380.310 ;
        RECT 700.185 379.630 724.650 379.930 ;
        RECT 854.990 379.930 855.290 380.310 ;
        RECT 855.910 379.930 856.210 380.990 ;
        RECT 903.750 380.610 904.050 380.990 ;
        RECT 952.510 380.990 1000.650 381.290 ;
        RECT 903.750 380.310 951.890 380.610 ;
        RECT 854.990 379.630 856.210 379.930 ;
        RECT 951.590 379.930 951.890 380.310 ;
        RECT 952.510 379.930 952.810 380.990 ;
        RECT 1000.350 380.610 1000.650 380.990 ;
        RECT 1049.110 380.990 1097.250 381.290 ;
        RECT 1000.350 380.310 1048.490 380.610 ;
        RECT 951.590 379.630 952.810 379.930 ;
        RECT 1048.190 379.930 1048.490 380.310 ;
        RECT 1049.110 379.930 1049.410 380.990 ;
        RECT 1096.950 380.610 1097.250 380.990 ;
        RECT 1145.710 380.990 1193.850 381.290 ;
        RECT 1096.950 380.310 1145.090 380.610 ;
        RECT 1048.190 379.630 1049.410 379.930 ;
        RECT 1144.790 379.930 1145.090 380.310 ;
        RECT 1145.710 379.930 1146.010 380.990 ;
        RECT 1193.550 380.610 1193.850 380.990 ;
        RECT 1242.310 380.990 1290.450 381.290 ;
        RECT 1193.550 380.310 1241.690 380.610 ;
        RECT 1144.790 379.630 1146.010 379.930 ;
        RECT 1241.390 379.930 1241.690 380.310 ;
        RECT 1242.310 379.930 1242.610 380.990 ;
        RECT 1290.150 380.610 1290.450 380.990 ;
        RECT 1338.910 380.990 1387.050 381.290 ;
        RECT 1290.150 380.310 1338.290 380.610 ;
        RECT 1241.390 379.630 1242.610 379.930 ;
        RECT 1337.990 379.930 1338.290 380.310 ;
        RECT 1338.910 379.930 1339.210 380.990 ;
        RECT 1386.750 380.610 1387.050 380.990 ;
        RECT 1435.510 380.990 1483.650 381.290 ;
        RECT 1386.750 380.310 1434.890 380.610 ;
        RECT 1337.990 379.630 1339.210 379.930 ;
        RECT 1434.590 379.930 1434.890 380.310 ;
        RECT 1435.510 379.930 1435.810 380.990 ;
        RECT 1483.350 380.610 1483.650 380.990 ;
        RECT 1532.110 380.990 1580.250 381.290 ;
        RECT 1483.350 380.310 1531.490 380.610 ;
        RECT 1434.590 379.630 1435.810 379.930 ;
        RECT 1531.190 379.930 1531.490 380.310 ;
        RECT 1532.110 379.930 1532.410 380.990 ;
        RECT 1579.950 380.610 1580.250 380.990 ;
        RECT 1628.710 380.990 1676.850 381.290 ;
        RECT 1579.950 380.310 1628.090 380.610 ;
        RECT 1531.190 379.630 1532.410 379.930 ;
        RECT 1627.790 379.930 1628.090 380.310 ;
        RECT 1628.710 379.930 1629.010 380.990 ;
        RECT 1676.550 380.610 1676.850 380.990 ;
        RECT 1725.310 380.990 1773.450 381.290 ;
        RECT 1676.550 380.310 1724.690 380.610 ;
        RECT 1627.790 379.630 1629.010 379.930 ;
        RECT 1724.390 379.930 1724.690 380.310 ;
        RECT 1725.310 379.930 1725.610 380.990 ;
        RECT 1773.150 380.610 1773.450 380.990 ;
        RECT 1821.910 380.990 1870.050 381.290 ;
        RECT 1773.150 380.310 1821.290 380.610 ;
        RECT 1724.390 379.630 1725.610 379.930 ;
        RECT 1820.990 379.930 1821.290 380.310 ;
        RECT 1821.910 379.930 1822.210 380.990 ;
        RECT 1869.750 380.610 1870.050 380.990 ;
        RECT 1918.510 380.990 1966.650 381.290 ;
        RECT 1869.750 380.310 1917.890 380.610 ;
        RECT 1820.990 379.630 1822.210 379.930 ;
        RECT 1917.590 379.930 1917.890 380.310 ;
        RECT 1918.510 379.930 1918.810 380.990 ;
        RECT 1966.350 380.610 1966.650 380.990 ;
        RECT 2015.110 380.990 2063.250 381.290 ;
        RECT 1966.350 380.310 2014.490 380.610 ;
        RECT 1917.590 379.630 1918.810 379.930 ;
        RECT 2014.190 379.930 2014.490 380.310 ;
        RECT 2015.110 379.930 2015.410 380.990 ;
        RECT 2062.950 380.610 2063.250 380.990 ;
        RECT 2111.710 380.990 2159.850 381.290 ;
        RECT 2062.950 380.310 2111.090 380.610 ;
        RECT 2014.190 379.630 2015.410 379.930 ;
        RECT 2110.790 379.930 2111.090 380.310 ;
        RECT 2111.710 379.930 2112.010 380.990 ;
        RECT 2159.550 380.610 2159.850 380.990 ;
        RECT 2208.310 380.990 2256.450 381.290 ;
        RECT 2159.550 380.310 2207.690 380.610 ;
        RECT 2110.790 379.630 2112.010 379.930 ;
        RECT 2207.390 379.930 2207.690 380.310 ;
        RECT 2208.310 379.930 2208.610 380.990 ;
        RECT 2256.150 380.610 2256.450 380.990 ;
        RECT 2304.910 380.990 2353.050 381.290 ;
        RECT 2256.150 380.310 2304.290 380.610 ;
        RECT 2207.390 379.630 2208.610 379.930 ;
        RECT 2303.990 379.930 2304.290 380.310 ;
        RECT 2304.910 379.930 2305.210 380.990 ;
        RECT 2352.750 380.610 2353.050 380.990 ;
        RECT 2401.510 380.990 2449.650 381.290 ;
        RECT 2352.750 380.310 2400.890 380.610 ;
        RECT 2303.990 379.630 2305.210 379.930 ;
        RECT 2400.590 379.930 2400.890 380.310 ;
        RECT 2401.510 379.930 2401.810 380.990 ;
        RECT 2449.350 380.610 2449.650 380.990 ;
        RECT 2498.110 380.990 2546.250 381.290 ;
        RECT 2449.350 380.310 2497.490 380.610 ;
        RECT 2400.590 379.630 2401.810 379.930 ;
        RECT 2497.190 379.930 2497.490 380.310 ;
        RECT 2498.110 379.930 2498.410 380.990 ;
        RECT 2545.950 380.610 2546.250 380.990 ;
        RECT 2594.710 380.990 2642.850 381.290 ;
        RECT 2545.950 380.310 2594.090 380.610 ;
        RECT 2497.190 379.630 2498.410 379.930 ;
        RECT 2593.790 379.930 2594.090 380.310 ;
        RECT 2594.710 379.930 2595.010 380.990 ;
        RECT 2642.550 380.610 2642.850 380.990 ;
        RECT 2691.310 380.990 2739.450 381.290 ;
        RECT 2642.550 380.310 2690.690 380.610 ;
        RECT 2593.790 379.630 2595.010 379.930 ;
        RECT 2690.390 379.930 2690.690 380.310 ;
        RECT 2691.310 379.930 2691.610 380.990 ;
        RECT 2739.150 380.610 2739.450 380.990 ;
        RECT 2787.910 380.990 2836.050 381.290 ;
        RECT 2739.150 380.310 2787.290 380.610 ;
        RECT 2690.390 379.630 2691.610 379.930 ;
        RECT 2786.990 379.930 2787.290 380.310 ;
        RECT 2787.910 379.930 2788.210 380.990 ;
        RECT 2835.750 380.610 2836.050 380.990 ;
        RECT 2916.710 380.990 2924.800 381.290 ;
        RECT 2916.710 380.610 2917.010 380.990 ;
        RECT 2835.750 380.310 2883.890 380.610 ;
        RECT 2786.990 379.630 2788.210 379.930 ;
        RECT 2883.590 379.930 2883.890 380.310 ;
        RECT 2884.510 380.310 2917.010 380.610 ;
        RECT 2917.600 380.540 2924.800 380.990 ;
        RECT 2884.510 379.930 2884.810 380.310 ;
        RECT 2883.590 379.630 2884.810 379.930 ;
        RECT 700.185 379.615 700.515 379.630 ;
        RECT 337.910 379.250 338.290 379.260 ;
        RECT 386.005 379.250 386.335 379.265 ;
        RECT 337.910 378.950 386.335 379.250 ;
        RECT 337.910 378.940 338.290 378.950 ;
        RECT 386.005 378.935 386.335 378.950 ;
      LAYER via3 ;
        RECT 287.340 1557.380 287.660 1557.700 ;
        RECT 627.740 382.340 628.060 382.660 ;
        RECT 287.340 380.980 287.660 381.300 ;
        RECT 337.940 380.300 338.260 380.620 ;
        RECT 578.980 381.660 579.300 381.980 ;
        RECT 627.740 380.980 628.060 381.300 ;
        RECT 578.980 379.620 579.300 379.940 ;
        RECT 337.940 378.940 338.260 379.260 ;
      LAYER met4 ;
        RECT 287.335 1557.375 287.665 1557.705 ;
        RECT 287.350 381.305 287.650 1557.375 ;
        RECT 627.735 382.335 628.065 382.665 ;
        RECT 578.975 381.655 579.305 381.985 ;
        RECT 287.335 380.975 287.665 381.305 ;
        RECT 337.935 380.295 338.265 380.625 ;
        RECT 337.950 379.265 338.250 380.295 ;
        RECT 578.990 379.945 579.290 381.655 ;
        RECT 627.750 381.305 628.050 382.335 ;
        RECT 627.735 380.975 628.065 381.305 ;
        RECT 578.975 379.615 579.305 379.945 ;
        RECT 337.935 378.935 338.265 379.265 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 293.550 3504.620 293.870 3504.680 ;
        RECT 1094.870 3504.620 1095.190 3504.680 ;
        RECT 293.550 3504.480 1095.190 3504.620 ;
        RECT 293.550 3504.420 293.870 3504.480 ;
        RECT 1094.870 3504.420 1095.190 3504.480 ;
      LAYER via ;
        RECT 293.580 3504.420 293.840 3504.680 ;
        RECT 1094.900 3504.420 1095.160 3504.680 ;
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
        RECT 1094.960 3504.710 1095.100 3517.600 ;
        RECT 293.580 3504.390 293.840 3504.710 ;
        RECT 1094.900 3504.390 1095.160 3504.710 ;
        RECT 293.640 2157.485 293.780 3504.390 ;
        RECT 293.570 2157.115 293.850 2157.485 ;
      LAYER via2 ;
        RECT 293.570 2157.160 293.850 2157.440 ;
      LAYER met3 ;
        RECT 293.545 2157.450 293.875 2157.465 ;
        RECT 300.000 2157.450 304.000 2157.520 ;
        RECT 293.545 2157.150 304.000 2157.450 ;
        RECT 293.545 2157.135 293.875 2157.150 ;
        RECT 300.000 2156.920 304.000 2157.150 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 288.030 3500.880 288.350 3500.940 ;
        RECT 770.570 3500.880 770.890 3500.940 ;
        RECT 288.030 3500.740 770.890 3500.880 ;
        RECT 288.030 3500.680 288.350 3500.740 ;
        RECT 770.570 3500.680 770.890 3500.740 ;
      LAYER via ;
        RECT 288.060 3500.680 288.320 3500.940 ;
        RECT 770.600 3500.680 770.860 3500.940 ;
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
        RECT 770.660 3500.970 770.800 3517.600 ;
        RECT 288.060 3500.650 288.320 3500.970 ;
        RECT 770.600 3500.650 770.860 3500.970 ;
        RECT 288.120 2189.445 288.260 3500.650 ;
        RECT 288.050 2189.075 288.330 2189.445 ;
      LAYER via2 ;
        RECT 288.050 2189.120 288.330 2189.400 ;
      LAYER met3 ;
        RECT 288.025 2189.410 288.355 2189.425 ;
        RECT 300.000 2189.410 304.000 2189.480 ;
        RECT 288.025 2189.110 304.000 2189.410 ;
        RECT 288.025 2189.095 288.355 2189.110 ;
        RECT 300.000 2188.880 304.000 2189.110 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 287.570 3500.540 287.890 3500.600 ;
        RECT 445.810 3500.540 446.130 3500.600 ;
        RECT 287.570 3500.400 446.130 3500.540 ;
        RECT 287.570 3500.340 287.890 3500.400 ;
        RECT 445.810 3500.340 446.130 3500.400 ;
        RECT 282.970 2243.220 283.290 2243.280 ;
        RECT 287.570 2243.220 287.890 2243.280 ;
        RECT 282.970 2243.080 287.890 2243.220 ;
        RECT 282.970 2243.020 283.290 2243.080 ;
        RECT 287.570 2243.020 287.890 2243.080 ;
      LAYER via ;
        RECT 287.600 3500.340 287.860 3500.600 ;
        RECT 445.840 3500.340 446.100 3500.600 ;
        RECT 283.000 2243.020 283.260 2243.280 ;
        RECT 287.600 2243.020 287.860 2243.280 ;
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
        RECT 445.900 3500.630 446.040 3517.600 ;
        RECT 287.600 3500.310 287.860 3500.630 ;
        RECT 445.840 3500.310 446.100 3500.630 ;
        RECT 287.660 2243.310 287.800 3500.310 ;
        RECT 283.000 2242.990 283.260 2243.310 ;
        RECT 287.600 2242.990 287.860 2243.310 ;
        RECT 283.060 2220.725 283.200 2242.990 ;
        RECT 282.990 2220.355 283.270 2220.725 ;
      LAYER via2 ;
        RECT 282.990 2220.400 283.270 2220.680 ;
      LAYER met3 ;
        RECT 282.965 2220.690 283.295 2220.705 ;
        RECT 300.000 2220.690 304.000 2220.760 ;
        RECT 282.965 2220.390 304.000 2220.690 ;
        RECT 282.965 2220.375 283.295 2220.390 ;
        RECT 300.000 2220.160 304.000 2220.390 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 121.510 3498.500 121.830 3498.560 ;
        RECT 123.810 3498.500 124.130 3498.560 ;
        RECT 121.510 3498.360 124.130 3498.500 ;
        RECT 121.510 3498.300 121.830 3498.360 ;
        RECT 123.810 3498.300 124.130 3498.360 ;
        RECT 123.810 2256.140 124.130 2256.200 ;
        RECT 282.970 2256.140 283.290 2256.200 ;
        RECT 123.810 2256.000 283.290 2256.140 ;
        RECT 123.810 2255.940 124.130 2256.000 ;
        RECT 282.970 2255.940 283.290 2256.000 ;
      LAYER via ;
        RECT 121.540 3498.300 121.800 3498.560 ;
        RECT 123.840 3498.300 124.100 3498.560 ;
        RECT 123.840 2255.940 124.100 2256.200 ;
        RECT 283.000 2255.940 283.260 2256.200 ;
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
        RECT 121.600 3498.590 121.740 3517.600 ;
        RECT 121.540 3498.270 121.800 3498.590 ;
        RECT 123.840 3498.270 124.100 3498.590 ;
        RECT 123.900 2256.230 124.040 3498.270 ;
        RECT 123.840 2255.910 124.100 2256.230 ;
        RECT 283.000 2255.910 283.260 2256.230 ;
        RECT 283.060 2252.685 283.200 2255.910 ;
        RECT 282.990 2252.315 283.270 2252.685 ;
      LAYER via2 ;
        RECT 282.990 2252.360 283.270 2252.640 ;
      LAYER met3 ;
        RECT 282.965 2252.650 283.295 2252.665 ;
        RECT 300.000 2252.650 304.000 2252.720 ;
        RECT 282.965 2252.350 304.000 2252.650 ;
        RECT 282.965 2252.335 283.295 2252.350 ;
        RECT 300.000 2252.120 304.000 2252.350 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 3339.720 17.410 3339.780 ;
        RECT 106.790 3339.720 107.110 3339.780 ;
        RECT 17.090 3339.580 107.110 3339.720 ;
        RECT 17.090 3339.520 17.410 3339.580 ;
        RECT 106.790 3339.520 107.110 3339.580 ;
        RECT 106.790 2283.680 107.110 2283.740 ;
        RECT 282.970 2283.680 283.290 2283.740 ;
        RECT 106.790 2283.540 283.290 2283.680 ;
        RECT 106.790 2283.480 107.110 2283.540 ;
        RECT 282.970 2283.480 283.290 2283.540 ;
      LAYER via ;
        RECT 17.120 3339.520 17.380 3339.780 ;
        RECT 106.820 3339.520 107.080 3339.780 ;
        RECT 106.820 2283.480 107.080 2283.740 ;
        RECT 283.000 2283.480 283.260 2283.740 ;
      LAYER met2 ;
        RECT 17.110 3339.635 17.390 3340.005 ;
        RECT 17.120 3339.490 17.380 3339.635 ;
        RECT 106.820 3339.490 107.080 3339.810 ;
        RECT 106.880 2283.770 107.020 3339.490 ;
        RECT 106.820 2283.450 107.080 2283.770 ;
        RECT 282.990 2283.595 283.270 2283.965 ;
        RECT 283.000 2283.450 283.260 2283.595 ;
      LAYER via2 ;
        RECT 17.110 3339.680 17.390 3339.960 ;
        RECT 282.990 2283.640 283.270 2283.920 ;
      LAYER met3 ;
        RECT -4.800 3339.970 2.400 3340.420 ;
        RECT 17.085 3339.970 17.415 3339.985 ;
        RECT -4.800 3339.670 17.415 3339.970 ;
        RECT -4.800 3339.220 2.400 3339.670 ;
        RECT 17.085 3339.655 17.415 3339.670 ;
        RECT 282.965 2283.930 283.295 2283.945 ;
        RECT 300.000 2283.930 304.000 2284.000 ;
        RECT 282.965 2283.630 304.000 2283.930 ;
        RECT 282.965 2283.615 283.295 2283.630 ;
        RECT 300.000 2283.400 304.000 2283.630 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 3050.040 17.410 3050.100 ;
        RECT 155.090 3050.040 155.410 3050.100 ;
        RECT 17.090 3049.900 155.410 3050.040 ;
        RECT 17.090 3049.840 17.410 3049.900 ;
        RECT 155.090 3049.840 155.410 3049.900 ;
        RECT 155.090 2318.360 155.410 2318.420 ;
        RECT 282.510 2318.360 282.830 2318.420 ;
        RECT 155.090 2318.220 282.830 2318.360 ;
        RECT 155.090 2318.160 155.410 2318.220 ;
        RECT 282.510 2318.160 282.830 2318.220 ;
      LAYER via ;
        RECT 17.120 3049.840 17.380 3050.100 ;
        RECT 155.120 3049.840 155.380 3050.100 ;
        RECT 155.120 2318.160 155.380 2318.420 ;
        RECT 282.540 2318.160 282.800 2318.420 ;
      LAYER met2 ;
        RECT 17.110 3051.995 17.390 3052.365 ;
        RECT 17.180 3050.130 17.320 3051.995 ;
        RECT 17.120 3049.810 17.380 3050.130 ;
        RECT 155.120 3049.810 155.380 3050.130 ;
        RECT 155.180 2318.450 155.320 3049.810 ;
        RECT 155.120 2318.130 155.380 2318.450 ;
        RECT 282.540 2318.130 282.800 2318.450 ;
        RECT 282.600 2317.965 282.740 2318.130 ;
        RECT 282.530 2317.595 282.810 2317.965 ;
      LAYER via2 ;
        RECT 17.110 3052.040 17.390 3052.320 ;
        RECT 282.530 2317.640 282.810 2317.920 ;
      LAYER met3 ;
        RECT -4.800 3052.330 2.400 3052.780 ;
        RECT 17.085 3052.330 17.415 3052.345 ;
        RECT -4.800 3052.030 17.415 3052.330 ;
        RECT -4.800 3051.580 2.400 3052.030 ;
        RECT 17.085 3052.015 17.415 3052.030 ;
        RECT 282.505 2317.930 282.835 2317.945 ;
        RECT 282.505 2317.630 300.530 2317.930 ;
        RECT 282.505 2317.615 282.835 2317.630 ;
        RECT 300.230 2315.960 300.530 2317.630 ;
        RECT 300.000 2315.360 304.000 2315.960 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 19.390 2352.700 19.710 2352.760 ;
        RECT 282.510 2352.700 282.830 2352.760 ;
        RECT 19.390 2352.560 282.830 2352.700 ;
        RECT 19.390 2352.500 19.710 2352.560 ;
        RECT 282.510 2352.500 282.830 2352.560 ;
      LAYER via ;
        RECT 19.420 2352.500 19.680 2352.760 ;
        RECT 282.540 2352.500 282.800 2352.760 ;
      LAYER met2 ;
        RECT 19.410 2765.035 19.690 2765.405 ;
        RECT 19.480 2352.790 19.620 2765.035 ;
        RECT 19.420 2352.470 19.680 2352.790 ;
        RECT 282.540 2352.470 282.800 2352.790 ;
        RECT 282.600 2349.925 282.740 2352.470 ;
        RECT 282.530 2349.555 282.810 2349.925 ;
      LAYER via2 ;
        RECT 19.410 2765.080 19.690 2765.360 ;
        RECT 282.530 2349.600 282.810 2349.880 ;
      LAYER met3 ;
        RECT -4.800 2765.370 2.400 2765.820 ;
        RECT 19.385 2765.370 19.715 2765.385 ;
        RECT -4.800 2765.070 19.715 2765.370 ;
        RECT -4.800 2764.620 2.400 2765.070 ;
        RECT 19.385 2765.055 19.715 2765.070 ;
        RECT 282.505 2349.890 282.835 2349.905 ;
        RECT 282.505 2349.590 300.530 2349.890 ;
        RECT 282.505 2349.575 282.835 2349.590 ;
        RECT 300.230 2347.240 300.530 2349.590 ;
        RECT 300.000 2346.640 304.000 2347.240 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 2380.240 16.950 2380.300 ;
        RECT 282.970 2380.240 283.290 2380.300 ;
        RECT 16.630 2380.100 283.290 2380.240 ;
        RECT 16.630 2380.040 16.950 2380.100 ;
        RECT 282.970 2380.040 283.290 2380.100 ;
      LAYER via ;
        RECT 16.660 2380.040 16.920 2380.300 ;
        RECT 283.000 2380.040 283.260 2380.300 ;
      LAYER met2 ;
        RECT 16.650 2477.395 16.930 2477.765 ;
        RECT 16.720 2380.330 16.860 2477.395 ;
        RECT 16.660 2380.010 16.920 2380.330 ;
        RECT 283.000 2380.010 283.260 2380.330 ;
        RECT 283.060 2379.165 283.200 2380.010 ;
        RECT 282.990 2378.795 283.270 2379.165 ;
      LAYER via2 ;
        RECT 16.650 2477.440 16.930 2477.720 ;
        RECT 282.990 2378.840 283.270 2379.120 ;
      LAYER met3 ;
        RECT -4.800 2477.730 2.400 2478.180 ;
        RECT 16.625 2477.730 16.955 2477.745 ;
        RECT -4.800 2477.430 16.955 2477.730 ;
        RECT -4.800 2476.980 2.400 2477.430 ;
        RECT 16.625 2477.415 16.955 2477.430 ;
        RECT 282.965 2379.130 283.295 2379.145 ;
        RECT 300.000 2379.130 304.000 2379.200 ;
        RECT 282.965 2378.830 304.000 2379.130 ;
        RECT 282.965 2378.815 283.295 2378.830 ;
        RECT 300.000 2378.600 304.000 2378.830 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 20.310 2408.460 20.630 2408.520 ;
        RECT 282.970 2408.460 283.290 2408.520 ;
        RECT 20.310 2408.320 283.290 2408.460 ;
        RECT 20.310 2408.260 20.630 2408.320 ;
        RECT 282.970 2408.260 283.290 2408.320 ;
      LAYER via ;
        RECT 20.340 2408.260 20.600 2408.520 ;
        RECT 283.000 2408.260 283.260 2408.520 ;
      LAYER met2 ;
        RECT 282.990 2410.075 283.270 2410.445 ;
        RECT 283.060 2408.550 283.200 2410.075 ;
        RECT 20.340 2408.230 20.600 2408.550 ;
        RECT 283.000 2408.230 283.260 2408.550 ;
        RECT 20.400 2190.125 20.540 2408.230 ;
        RECT 20.330 2189.755 20.610 2190.125 ;
      LAYER via2 ;
        RECT 282.990 2410.120 283.270 2410.400 ;
        RECT 20.330 2189.800 20.610 2190.080 ;
      LAYER met3 ;
        RECT 282.965 2410.410 283.295 2410.425 ;
        RECT 300.000 2410.410 304.000 2410.480 ;
        RECT 282.965 2410.110 304.000 2410.410 ;
        RECT 282.965 2410.095 283.295 2410.110 ;
        RECT 300.000 2409.880 304.000 2410.110 ;
        RECT -4.800 2190.090 2.400 2190.540 ;
        RECT 20.305 2190.090 20.635 2190.105 ;
        RECT -4.800 2189.790 20.635 2190.090 ;
        RECT -4.800 2189.340 2.400 2189.790 ;
        RECT 20.305 2189.775 20.635 2189.790 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.470 2436.000 18.790 2436.060 ;
        RECT 282.970 2436.000 283.290 2436.060 ;
        RECT 18.470 2435.860 283.290 2436.000 ;
        RECT 18.470 2435.800 18.790 2435.860 ;
        RECT 282.970 2435.800 283.290 2435.860 ;
      LAYER via ;
        RECT 18.500 2435.800 18.760 2436.060 ;
        RECT 283.000 2435.800 283.260 2436.060 ;
      LAYER met2 ;
        RECT 282.990 2441.355 283.270 2441.725 ;
        RECT 283.060 2436.090 283.200 2441.355 ;
        RECT 18.500 2435.770 18.760 2436.090 ;
        RECT 283.000 2435.770 283.260 2436.090 ;
        RECT 18.560 1903.165 18.700 2435.770 ;
        RECT 18.490 1902.795 18.770 1903.165 ;
      LAYER via2 ;
        RECT 282.990 2441.400 283.270 2441.680 ;
        RECT 18.490 1902.840 18.770 1903.120 ;
      LAYER met3 ;
        RECT 282.965 2441.690 283.295 2441.705 ;
        RECT 300.000 2441.690 304.000 2441.760 ;
        RECT 282.965 2441.390 304.000 2441.690 ;
        RECT 282.965 2441.375 283.295 2441.390 ;
        RECT 300.000 2441.160 304.000 2441.390 ;
        RECT -4.800 1903.130 2.400 1903.580 ;
        RECT 18.465 1903.130 18.795 1903.145 ;
        RECT -4.800 1902.830 18.795 1903.130 ;
        RECT -4.800 1902.380 2.400 1902.830 ;
        RECT 18.465 1902.815 18.795 1902.830 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 288.950 620.740 289.270 620.800 ;
        RECT 2900.830 620.740 2901.150 620.800 ;
        RECT 288.950 620.600 2901.150 620.740 ;
        RECT 288.950 620.540 289.270 620.600 ;
        RECT 2900.830 620.540 2901.150 620.600 ;
      LAYER via ;
        RECT 288.980 620.540 289.240 620.800 ;
        RECT 2900.860 620.540 2901.120 620.800 ;
      LAYER met2 ;
        RECT 288.970 1588.635 289.250 1589.005 ;
        RECT 289.040 620.830 289.180 1588.635 ;
        RECT 288.980 620.510 289.240 620.830 ;
        RECT 2900.860 620.510 2901.120 620.830 ;
        RECT 2900.920 615.925 2901.060 620.510 ;
        RECT 2900.850 615.555 2901.130 615.925 ;
      LAYER via2 ;
        RECT 288.970 1588.680 289.250 1588.960 ;
        RECT 2900.850 615.600 2901.130 615.880 ;
      LAYER met3 ;
        RECT 288.945 1588.970 289.275 1588.985 ;
        RECT 300.000 1588.970 304.000 1589.040 ;
        RECT 288.945 1588.670 304.000 1588.970 ;
        RECT 288.945 1588.655 289.275 1588.670 ;
        RECT 300.000 1588.440 304.000 1588.670 ;
        RECT 2900.825 615.890 2901.155 615.905 ;
        RECT 2917.600 615.890 2924.800 616.340 ;
        RECT 2900.825 615.590 2924.800 615.890 ;
        RECT 2900.825 615.575 2901.155 615.590 ;
        RECT 2917.600 615.140 2924.800 615.590 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 161.990 2470.340 162.310 2470.400 ;
        RECT 286.190 2470.340 286.510 2470.400 ;
        RECT 161.990 2470.200 286.510 2470.340 ;
        RECT 161.990 2470.140 162.310 2470.200 ;
        RECT 286.190 2470.140 286.510 2470.200 ;
        RECT 15.250 1621.360 15.570 1621.420 ;
        RECT 161.990 1621.360 162.310 1621.420 ;
        RECT 15.250 1621.220 162.310 1621.360 ;
        RECT 15.250 1621.160 15.570 1621.220 ;
        RECT 161.990 1621.160 162.310 1621.220 ;
      LAYER via ;
        RECT 162.020 2470.140 162.280 2470.400 ;
        RECT 286.220 2470.140 286.480 2470.400 ;
        RECT 15.280 1621.160 15.540 1621.420 ;
        RECT 162.020 1621.160 162.280 1621.420 ;
      LAYER met2 ;
        RECT 286.210 2473.315 286.490 2473.685 ;
        RECT 286.280 2470.430 286.420 2473.315 ;
        RECT 162.020 2470.110 162.280 2470.430 ;
        RECT 286.220 2470.110 286.480 2470.430 ;
        RECT 162.080 1621.450 162.220 2470.110 ;
        RECT 15.280 1621.130 15.540 1621.450 ;
        RECT 162.020 1621.130 162.280 1621.450 ;
        RECT 15.340 1615.525 15.480 1621.130 ;
        RECT 15.270 1615.155 15.550 1615.525 ;
      LAYER via2 ;
        RECT 286.210 2473.360 286.490 2473.640 ;
        RECT 15.270 1615.200 15.550 1615.480 ;
      LAYER met3 ;
        RECT 286.185 2473.650 286.515 2473.665 ;
        RECT 300.000 2473.650 304.000 2473.720 ;
        RECT 286.185 2473.350 304.000 2473.650 ;
        RECT 286.185 2473.335 286.515 2473.350 ;
        RECT 300.000 2473.120 304.000 2473.350 ;
        RECT -4.800 1615.490 2.400 1615.940 ;
        RECT 15.245 1615.490 15.575 1615.505 ;
        RECT -4.800 1615.190 15.575 1615.490 ;
        RECT -4.800 1614.740 2.400 1615.190 ;
        RECT 15.245 1615.175 15.575 1615.190 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 189.590 2505.020 189.910 2505.080 ;
        RECT 286.190 2505.020 286.510 2505.080 ;
        RECT 189.590 2504.880 286.510 2505.020 ;
        RECT 189.590 2504.820 189.910 2504.880 ;
        RECT 286.190 2504.820 286.510 2504.880 ;
        RECT 16.630 1400.700 16.950 1400.760 ;
        RECT 189.590 1400.700 189.910 1400.760 ;
        RECT 16.630 1400.560 189.910 1400.700 ;
        RECT 16.630 1400.500 16.950 1400.560 ;
        RECT 189.590 1400.500 189.910 1400.560 ;
      LAYER via ;
        RECT 189.620 2504.820 189.880 2505.080 ;
        RECT 286.220 2504.820 286.480 2505.080 ;
        RECT 16.660 1400.500 16.920 1400.760 ;
        RECT 189.620 1400.500 189.880 1400.760 ;
      LAYER met2 ;
        RECT 189.620 2504.790 189.880 2505.110 ;
        RECT 286.220 2504.965 286.480 2505.110 ;
        RECT 189.680 1400.790 189.820 2504.790 ;
        RECT 286.210 2504.595 286.490 2504.965 ;
        RECT 16.660 1400.645 16.920 1400.790 ;
        RECT 16.650 1400.275 16.930 1400.645 ;
        RECT 189.620 1400.470 189.880 1400.790 ;
      LAYER via2 ;
        RECT 286.210 2504.640 286.490 2504.920 ;
        RECT 16.650 1400.320 16.930 1400.600 ;
      LAYER met3 ;
        RECT 286.185 2504.930 286.515 2504.945 ;
        RECT 300.000 2504.930 304.000 2505.000 ;
        RECT 286.185 2504.630 304.000 2504.930 ;
        RECT 286.185 2504.615 286.515 2504.630 ;
        RECT 300.000 2504.400 304.000 2504.630 ;
        RECT -4.800 1400.610 2.400 1401.060 ;
        RECT 16.625 1400.610 16.955 1400.625 ;
        RECT -4.800 1400.310 16.955 1400.610 ;
        RECT -4.800 1399.860 2.400 1400.310 ;
        RECT 16.625 1400.295 16.955 1400.310 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 196.950 2532.560 197.270 2532.620 ;
        RECT 286.190 2532.560 286.510 2532.620 ;
        RECT 196.950 2532.420 286.510 2532.560 ;
        RECT 196.950 2532.360 197.270 2532.420 ;
        RECT 286.190 2532.360 286.510 2532.420 ;
        RECT 16.170 1186.840 16.490 1186.900 ;
        RECT 196.950 1186.840 197.270 1186.900 ;
        RECT 16.170 1186.700 197.270 1186.840 ;
        RECT 16.170 1186.640 16.490 1186.700 ;
        RECT 196.950 1186.640 197.270 1186.700 ;
      LAYER via ;
        RECT 196.980 2532.360 197.240 2532.620 ;
        RECT 286.220 2532.360 286.480 2532.620 ;
        RECT 16.200 1186.640 16.460 1186.900 ;
        RECT 196.980 1186.640 197.240 1186.900 ;
      LAYER met2 ;
        RECT 286.210 2536.555 286.490 2536.925 ;
        RECT 286.280 2532.650 286.420 2536.555 ;
        RECT 196.980 2532.330 197.240 2532.650 ;
        RECT 286.220 2532.330 286.480 2532.650 ;
        RECT 197.040 1186.930 197.180 2532.330 ;
        RECT 16.200 1186.610 16.460 1186.930 ;
        RECT 196.980 1186.610 197.240 1186.930 ;
        RECT 16.260 1185.085 16.400 1186.610 ;
        RECT 16.190 1184.715 16.470 1185.085 ;
      LAYER via2 ;
        RECT 286.210 2536.600 286.490 2536.880 ;
        RECT 16.190 1184.760 16.470 1185.040 ;
      LAYER met3 ;
        RECT 286.185 2536.890 286.515 2536.905 ;
        RECT 300.000 2536.890 304.000 2536.960 ;
        RECT 286.185 2536.590 304.000 2536.890 ;
        RECT 286.185 2536.575 286.515 2536.590 ;
        RECT 300.000 2536.360 304.000 2536.590 ;
        RECT -4.800 1185.050 2.400 1185.500 ;
        RECT 16.165 1185.050 16.495 1185.065 ;
        RECT -4.800 1184.750 16.495 1185.050 ;
        RECT -4.800 1184.300 2.400 1184.750 ;
        RECT 16.165 1184.735 16.495 1184.750 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 251.690 2566.900 252.010 2566.960 ;
        RECT 286.190 2566.900 286.510 2566.960 ;
        RECT 251.690 2566.760 286.510 2566.900 ;
        RECT 251.690 2566.700 252.010 2566.760 ;
        RECT 286.190 2566.700 286.510 2566.760 ;
        RECT 17.550 972.640 17.870 972.700 ;
        RECT 251.690 972.640 252.010 972.700 ;
        RECT 17.550 972.500 252.010 972.640 ;
        RECT 17.550 972.440 17.870 972.500 ;
        RECT 251.690 972.440 252.010 972.500 ;
      LAYER via ;
        RECT 251.720 2566.700 251.980 2566.960 ;
        RECT 286.220 2566.700 286.480 2566.960 ;
        RECT 17.580 972.440 17.840 972.700 ;
        RECT 251.720 972.440 251.980 972.700 ;
      LAYER met2 ;
        RECT 286.210 2567.835 286.490 2568.205 ;
        RECT 286.280 2566.990 286.420 2567.835 ;
        RECT 251.720 2566.670 251.980 2566.990 ;
        RECT 286.220 2566.670 286.480 2566.990 ;
        RECT 251.780 972.730 251.920 2566.670 ;
        RECT 17.580 972.410 17.840 972.730 ;
        RECT 251.720 972.410 251.980 972.730 ;
        RECT 17.640 969.525 17.780 972.410 ;
        RECT 17.570 969.155 17.850 969.525 ;
      LAYER via2 ;
        RECT 286.210 2567.880 286.490 2568.160 ;
        RECT 17.570 969.200 17.850 969.480 ;
      LAYER met3 ;
        RECT 286.185 2568.170 286.515 2568.185 ;
        RECT 300.000 2568.170 304.000 2568.240 ;
        RECT 286.185 2567.870 304.000 2568.170 ;
        RECT 286.185 2567.855 286.515 2567.870 ;
        RECT 300.000 2567.640 304.000 2567.870 ;
        RECT -4.800 969.490 2.400 969.940 ;
        RECT 17.545 969.490 17.875 969.505 ;
        RECT -4.800 969.190 17.875 969.490 ;
        RECT -4.800 968.740 2.400 969.190 ;
        RECT 17.545 969.175 17.875 969.190 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 258.590 2594.780 258.910 2594.840 ;
        RECT 286.190 2594.780 286.510 2594.840 ;
        RECT 258.590 2594.640 286.510 2594.780 ;
        RECT 258.590 2594.580 258.910 2594.640 ;
        RECT 286.190 2594.580 286.510 2594.640 ;
        RECT 15.710 758.780 16.030 758.840 ;
        RECT 258.590 758.780 258.910 758.840 ;
        RECT 15.710 758.640 258.910 758.780 ;
        RECT 15.710 758.580 16.030 758.640 ;
        RECT 258.590 758.580 258.910 758.640 ;
      LAYER via ;
        RECT 258.620 2594.580 258.880 2594.840 ;
        RECT 286.220 2594.580 286.480 2594.840 ;
        RECT 15.740 758.580 16.000 758.840 ;
        RECT 258.620 758.580 258.880 758.840 ;
      LAYER met2 ;
        RECT 286.210 2599.795 286.490 2600.165 ;
        RECT 286.280 2594.870 286.420 2599.795 ;
        RECT 258.620 2594.550 258.880 2594.870 ;
        RECT 286.220 2594.550 286.480 2594.870 ;
        RECT 258.680 758.870 258.820 2594.550 ;
        RECT 15.740 758.550 16.000 758.870 ;
        RECT 258.620 758.550 258.880 758.870 ;
        RECT 15.800 753.965 15.940 758.550 ;
        RECT 15.730 753.595 16.010 753.965 ;
      LAYER via2 ;
        RECT 286.210 2599.840 286.490 2600.120 ;
        RECT 15.730 753.640 16.010 753.920 ;
      LAYER met3 ;
        RECT 286.185 2600.130 286.515 2600.145 ;
        RECT 300.000 2600.130 304.000 2600.200 ;
        RECT 286.185 2599.830 304.000 2600.130 ;
        RECT 286.185 2599.815 286.515 2599.830 ;
        RECT 300.000 2599.600 304.000 2599.830 ;
        RECT -4.800 753.930 2.400 754.380 ;
        RECT 15.705 753.930 16.035 753.945 ;
        RECT -4.800 753.630 16.035 753.930 ;
        RECT -4.800 753.180 2.400 753.630 ;
        RECT 15.705 753.615 16.035 753.630 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 86.090 2629.120 86.410 2629.180 ;
        RECT 286.190 2629.120 286.510 2629.180 ;
        RECT 86.090 2628.980 286.510 2629.120 ;
        RECT 86.090 2628.920 86.410 2628.980 ;
        RECT 286.190 2628.920 286.510 2628.980 ;
        RECT 16.170 544.920 16.490 544.980 ;
        RECT 86.090 544.920 86.410 544.980 ;
        RECT 16.170 544.780 86.410 544.920 ;
        RECT 16.170 544.720 16.490 544.780 ;
        RECT 86.090 544.720 86.410 544.780 ;
      LAYER via ;
        RECT 86.120 2628.920 86.380 2629.180 ;
        RECT 286.220 2628.920 286.480 2629.180 ;
        RECT 16.200 544.720 16.460 544.980 ;
        RECT 86.120 544.720 86.380 544.980 ;
      LAYER met2 ;
        RECT 286.210 2631.075 286.490 2631.445 ;
        RECT 286.280 2629.210 286.420 2631.075 ;
        RECT 86.120 2628.890 86.380 2629.210 ;
        RECT 286.220 2628.890 286.480 2629.210 ;
        RECT 86.180 545.010 86.320 2628.890 ;
        RECT 16.200 544.690 16.460 545.010 ;
        RECT 86.120 544.690 86.380 545.010 ;
        RECT 16.260 538.405 16.400 544.690 ;
        RECT 16.190 538.035 16.470 538.405 ;
      LAYER via2 ;
        RECT 286.210 2631.120 286.490 2631.400 ;
        RECT 16.190 538.080 16.470 538.360 ;
      LAYER met3 ;
        RECT 286.185 2631.410 286.515 2631.425 ;
        RECT 300.000 2631.410 304.000 2631.480 ;
        RECT 286.185 2631.110 304.000 2631.410 ;
        RECT 286.185 2631.095 286.515 2631.110 ;
        RECT 300.000 2630.880 304.000 2631.110 ;
        RECT -4.800 538.370 2.400 538.820 ;
        RECT 16.165 538.370 16.495 538.385 ;
        RECT -4.800 538.070 16.495 538.370 ;
        RECT -4.800 537.620 2.400 538.070 ;
        RECT 16.165 538.055 16.495 538.070 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 265.490 2657.000 265.810 2657.060 ;
        RECT 286.190 2657.000 286.510 2657.060 ;
        RECT 265.490 2656.860 286.510 2657.000 ;
        RECT 265.490 2656.800 265.810 2656.860 ;
        RECT 286.190 2656.800 286.510 2656.860 ;
        RECT 16.630 324.260 16.950 324.320 ;
        RECT 265.490 324.260 265.810 324.320 ;
        RECT 16.630 324.120 265.810 324.260 ;
        RECT 16.630 324.060 16.950 324.120 ;
        RECT 265.490 324.060 265.810 324.120 ;
      LAYER via ;
        RECT 265.520 2656.800 265.780 2657.060 ;
        RECT 286.220 2656.800 286.480 2657.060 ;
        RECT 16.660 324.060 16.920 324.320 ;
        RECT 265.520 324.060 265.780 324.320 ;
      LAYER met2 ;
        RECT 286.210 2663.035 286.490 2663.405 ;
        RECT 286.280 2657.090 286.420 2663.035 ;
        RECT 265.520 2656.770 265.780 2657.090 ;
        RECT 286.220 2656.770 286.480 2657.090 ;
        RECT 265.580 324.350 265.720 2656.770 ;
        RECT 16.660 324.030 16.920 324.350 ;
        RECT 265.520 324.030 265.780 324.350 ;
        RECT 16.720 322.845 16.860 324.030 ;
        RECT 16.650 322.475 16.930 322.845 ;
      LAYER via2 ;
        RECT 286.210 2663.080 286.490 2663.360 ;
        RECT 16.650 322.520 16.930 322.800 ;
      LAYER met3 ;
        RECT 286.185 2663.370 286.515 2663.385 ;
        RECT 300.000 2663.370 304.000 2663.440 ;
        RECT 286.185 2663.070 304.000 2663.370 ;
        RECT 286.185 2663.055 286.515 2663.070 ;
        RECT 300.000 2662.840 304.000 2663.070 ;
        RECT -4.800 322.810 2.400 323.260 ;
        RECT 16.625 322.810 16.955 322.825 ;
        RECT -4.800 322.510 16.955 322.810 ;
        RECT -4.800 322.060 2.400 322.510 ;
        RECT 16.625 322.495 16.955 322.510 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 99.890 2691.340 100.210 2691.400 ;
        RECT 286.190 2691.340 286.510 2691.400 ;
        RECT 99.890 2691.200 286.510 2691.340 ;
        RECT 99.890 2691.140 100.210 2691.200 ;
        RECT 286.190 2691.140 286.510 2691.200 ;
        RECT 14.330 110.400 14.650 110.460 ;
        RECT 99.890 110.400 100.210 110.460 ;
        RECT 14.330 110.260 100.210 110.400 ;
        RECT 14.330 110.200 14.650 110.260 ;
        RECT 99.890 110.200 100.210 110.260 ;
      LAYER via ;
        RECT 99.920 2691.140 100.180 2691.400 ;
        RECT 286.220 2691.140 286.480 2691.400 ;
        RECT 14.360 110.200 14.620 110.460 ;
        RECT 99.920 110.200 100.180 110.460 ;
      LAYER met2 ;
        RECT 286.210 2694.315 286.490 2694.685 ;
        RECT 286.280 2691.430 286.420 2694.315 ;
        RECT 99.920 2691.110 100.180 2691.430 ;
        RECT 286.220 2691.110 286.480 2691.430 ;
        RECT 99.980 110.490 100.120 2691.110 ;
        RECT 14.360 110.170 14.620 110.490 ;
        RECT 99.920 110.170 100.180 110.490 ;
        RECT 14.420 107.285 14.560 110.170 ;
        RECT 14.350 106.915 14.630 107.285 ;
      LAYER via2 ;
        RECT 286.210 2694.360 286.490 2694.640 ;
        RECT 14.350 106.960 14.630 107.240 ;
      LAYER met3 ;
        RECT 286.185 2694.650 286.515 2694.665 ;
        RECT 300.000 2694.650 304.000 2694.720 ;
        RECT 286.185 2694.350 304.000 2694.650 ;
        RECT 286.185 2694.335 286.515 2694.350 ;
        RECT 300.000 2694.120 304.000 2694.350 ;
        RECT -4.800 107.250 2.400 107.700 ;
        RECT 14.325 107.250 14.655 107.265 ;
        RECT -4.800 106.950 14.655 107.250 ;
        RECT -4.800 106.500 2.400 106.950 ;
        RECT 14.325 106.935 14.655 106.950 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 288.490 1579.200 288.810 1579.260 ;
        RECT 289.870 1579.200 290.190 1579.260 ;
        RECT 288.490 1579.060 290.190 1579.200 ;
        RECT 288.490 1579.000 288.810 1579.060 ;
        RECT 289.870 1579.000 290.190 1579.060 ;
        RECT 288.030 1531.940 288.350 1532.000 ;
        RECT 289.870 1531.940 290.190 1532.000 ;
        RECT 288.030 1531.800 290.190 1531.940 ;
        RECT 288.030 1531.740 288.350 1531.800 ;
        RECT 289.870 1531.740 290.190 1531.800 ;
        RECT 283.890 1435.720 284.210 1435.780 ;
        RECT 288.030 1435.720 288.350 1435.780 ;
        RECT 283.890 1435.580 288.350 1435.720 ;
        RECT 283.890 1435.520 284.210 1435.580 ;
        RECT 288.030 1435.520 288.350 1435.580 ;
        RECT 288.030 1386.760 288.350 1386.820 ;
        RECT 289.410 1386.760 289.730 1386.820 ;
        RECT 288.030 1386.620 289.730 1386.760 ;
        RECT 288.030 1386.560 288.350 1386.620 ;
        RECT 289.410 1386.560 289.730 1386.620 ;
        RECT 288.030 1342.220 288.350 1342.280 ;
        RECT 289.410 1342.220 289.730 1342.280 ;
        RECT 288.030 1342.080 289.730 1342.220 ;
        RECT 288.030 1342.020 288.350 1342.080 ;
        RECT 289.410 1342.020 289.730 1342.080 ;
        RECT 288.030 855.340 288.350 855.400 ;
        RECT 2900.830 855.340 2901.150 855.400 ;
        RECT 288.030 855.200 2901.150 855.340 ;
        RECT 288.030 855.140 288.350 855.200 ;
        RECT 2900.830 855.140 2901.150 855.200 ;
      LAYER via ;
        RECT 288.520 1579.000 288.780 1579.260 ;
        RECT 289.900 1579.000 290.160 1579.260 ;
        RECT 288.060 1531.740 288.320 1532.000 ;
        RECT 289.900 1531.740 290.160 1532.000 ;
        RECT 283.920 1435.520 284.180 1435.780 ;
        RECT 288.060 1435.520 288.320 1435.780 ;
        RECT 288.060 1386.560 288.320 1386.820 ;
        RECT 289.440 1386.560 289.700 1386.820 ;
        RECT 288.060 1342.020 288.320 1342.280 ;
        RECT 289.440 1342.020 289.700 1342.280 ;
        RECT 288.060 855.140 288.320 855.400 ;
        RECT 2900.860 855.140 2901.120 855.400 ;
      LAYER met2 ;
        RECT 288.510 1620.595 288.790 1620.965 ;
        RECT 288.580 1579.290 288.720 1620.595 ;
        RECT 288.520 1578.970 288.780 1579.290 ;
        RECT 289.900 1578.970 290.160 1579.290 ;
        RECT 289.960 1532.030 290.100 1578.970 ;
        RECT 288.060 1531.710 288.320 1532.030 ;
        RECT 289.900 1531.710 290.160 1532.030 ;
        RECT 288.120 1483.605 288.260 1531.710 ;
        RECT 283.910 1483.235 284.190 1483.605 ;
        RECT 288.050 1483.235 288.330 1483.605 ;
        RECT 283.980 1435.810 284.120 1483.235 ;
        RECT 283.920 1435.490 284.180 1435.810 ;
        RECT 288.060 1435.490 288.320 1435.810 ;
        RECT 288.120 1386.850 288.260 1435.490 ;
        RECT 288.060 1386.530 288.320 1386.850 ;
        RECT 289.440 1386.530 289.700 1386.850 ;
        RECT 289.500 1342.310 289.640 1386.530 ;
        RECT 288.060 1341.990 288.320 1342.310 ;
        RECT 289.440 1341.990 289.700 1342.310 ;
        RECT 288.120 855.430 288.260 1341.990 ;
        RECT 288.060 855.110 288.320 855.430 ;
        RECT 2900.860 855.110 2901.120 855.430 ;
        RECT 2900.920 850.525 2901.060 855.110 ;
        RECT 2900.850 850.155 2901.130 850.525 ;
      LAYER via2 ;
        RECT 288.510 1620.640 288.790 1620.920 ;
        RECT 283.910 1483.280 284.190 1483.560 ;
        RECT 288.050 1483.280 288.330 1483.560 ;
        RECT 2900.850 850.200 2901.130 850.480 ;
      LAYER met3 ;
        RECT 288.485 1620.930 288.815 1620.945 ;
        RECT 300.000 1620.930 304.000 1621.000 ;
        RECT 288.485 1620.630 304.000 1620.930 ;
        RECT 288.485 1620.615 288.815 1620.630 ;
        RECT 300.000 1620.400 304.000 1620.630 ;
        RECT 283.885 1483.570 284.215 1483.585 ;
        RECT 288.025 1483.570 288.355 1483.585 ;
        RECT 283.885 1483.270 288.355 1483.570 ;
        RECT 283.885 1483.255 284.215 1483.270 ;
        RECT 288.025 1483.255 288.355 1483.270 ;
        RECT 2900.825 850.490 2901.155 850.505 ;
        RECT 2917.600 850.490 2924.800 850.940 ;
        RECT 2900.825 850.190 2924.800 850.490 ;
        RECT 2900.825 850.175 2901.155 850.190 ;
        RECT 2917.600 849.740 2924.800 850.190 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 283.430 1483.320 283.750 1483.380 ;
        RECT 286.650 1483.320 286.970 1483.380 ;
        RECT 283.430 1483.180 286.970 1483.320 ;
        RECT 283.430 1483.120 283.750 1483.180 ;
        RECT 286.650 1483.120 286.970 1483.180 ;
        RECT 283.430 1435.380 283.750 1435.440 ;
        RECT 286.650 1435.380 286.970 1435.440 ;
        RECT 283.430 1435.240 286.970 1435.380 ;
        RECT 283.430 1435.180 283.750 1435.240 ;
        RECT 286.650 1435.180 286.970 1435.240 ;
        RECT 283.890 1342.220 284.210 1342.280 ;
        RECT 286.650 1342.220 286.970 1342.280 ;
        RECT 283.890 1342.080 286.970 1342.220 ;
        RECT 283.890 1342.020 284.210 1342.080 ;
        RECT 286.650 1342.020 286.970 1342.080 ;
        RECT 286.650 1089.940 286.970 1090.000 ;
        RECT 2900.830 1089.940 2901.150 1090.000 ;
        RECT 286.650 1089.800 2901.150 1089.940 ;
        RECT 286.650 1089.740 286.970 1089.800 ;
        RECT 2900.830 1089.740 2901.150 1089.800 ;
      LAYER via ;
        RECT 283.460 1483.120 283.720 1483.380 ;
        RECT 286.680 1483.120 286.940 1483.380 ;
        RECT 283.460 1435.180 283.720 1435.440 ;
        RECT 286.680 1435.180 286.940 1435.440 ;
        RECT 283.920 1342.020 284.180 1342.280 ;
        RECT 286.680 1342.020 286.940 1342.280 ;
        RECT 286.680 1089.740 286.940 1090.000 ;
        RECT 2900.860 1089.740 2901.120 1090.000 ;
      LAYER met2 ;
        RECT 286.670 1651.875 286.950 1652.245 ;
        RECT 286.740 1580.165 286.880 1651.875 ;
        RECT 286.670 1579.795 286.950 1580.165 ;
        RECT 286.670 1532.195 286.950 1532.565 ;
        RECT 286.740 1483.410 286.880 1532.195 ;
        RECT 283.460 1483.090 283.720 1483.410 ;
        RECT 286.680 1483.090 286.940 1483.410 ;
        RECT 283.520 1435.470 283.660 1483.090 ;
        RECT 283.460 1435.150 283.720 1435.470 ;
        RECT 286.680 1435.150 286.940 1435.470 ;
        RECT 286.740 1387.045 286.880 1435.150 ;
        RECT 283.910 1386.675 284.190 1387.045 ;
        RECT 286.670 1386.675 286.950 1387.045 ;
        RECT 283.980 1342.310 284.120 1386.675 ;
        RECT 283.920 1341.990 284.180 1342.310 ;
        RECT 286.680 1341.990 286.940 1342.310 ;
        RECT 286.740 1090.030 286.880 1341.990 ;
        RECT 286.680 1089.710 286.940 1090.030 ;
        RECT 2900.860 1089.710 2901.120 1090.030 ;
        RECT 2900.920 1085.125 2901.060 1089.710 ;
        RECT 2900.850 1084.755 2901.130 1085.125 ;
      LAYER via2 ;
        RECT 286.670 1651.920 286.950 1652.200 ;
        RECT 286.670 1579.840 286.950 1580.120 ;
        RECT 286.670 1532.240 286.950 1532.520 ;
        RECT 283.910 1386.720 284.190 1387.000 ;
        RECT 286.670 1386.720 286.950 1387.000 ;
        RECT 2900.850 1084.800 2901.130 1085.080 ;
      LAYER met3 ;
        RECT 286.645 1652.210 286.975 1652.225 ;
        RECT 300.000 1652.210 304.000 1652.280 ;
        RECT 286.645 1651.910 304.000 1652.210 ;
        RECT 286.645 1651.895 286.975 1651.910 ;
        RECT 300.000 1651.680 304.000 1651.910 ;
        RECT 286.645 1580.140 286.975 1580.145 ;
        RECT 286.390 1580.130 286.975 1580.140 ;
        RECT 286.190 1579.830 286.975 1580.130 ;
        RECT 286.390 1579.820 286.975 1579.830 ;
        RECT 286.645 1579.815 286.975 1579.820 ;
        RECT 286.645 1532.540 286.975 1532.545 ;
        RECT 286.390 1532.530 286.975 1532.540 ;
        RECT 286.390 1532.230 287.200 1532.530 ;
        RECT 286.390 1532.220 286.975 1532.230 ;
        RECT 286.645 1532.215 286.975 1532.220 ;
        RECT 283.885 1387.010 284.215 1387.025 ;
        RECT 286.645 1387.010 286.975 1387.025 ;
        RECT 283.885 1386.710 286.975 1387.010 ;
        RECT 283.885 1386.695 284.215 1386.710 ;
        RECT 286.645 1386.695 286.975 1386.710 ;
        RECT 2900.825 1085.090 2901.155 1085.105 ;
        RECT 2917.600 1085.090 2924.800 1085.540 ;
        RECT 2900.825 1084.790 2924.800 1085.090 ;
        RECT 2900.825 1084.775 2901.155 1084.790 ;
        RECT 2917.600 1084.340 2924.800 1084.790 ;
      LAYER via3 ;
        RECT 286.420 1579.820 286.740 1580.140 ;
        RECT 286.420 1532.220 286.740 1532.540 ;
      LAYER met4 ;
        RECT 286.415 1579.815 286.745 1580.145 ;
        RECT 286.430 1532.545 286.730 1579.815 ;
        RECT 286.415 1532.215 286.745 1532.545 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 284.810 1324.540 285.130 1324.600 ;
        RECT 2900.830 1324.540 2901.150 1324.600 ;
        RECT 284.810 1324.400 2901.150 1324.540 ;
        RECT 284.810 1324.340 285.130 1324.400 ;
        RECT 2900.830 1324.340 2901.150 1324.400 ;
      LAYER via ;
        RECT 284.840 1324.340 285.100 1324.600 ;
        RECT 2900.860 1324.340 2901.120 1324.600 ;
      LAYER met2 ;
        RECT 284.830 1683.835 285.110 1684.205 ;
        RECT 284.900 1324.630 285.040 1683.835 ;
        RECT 284.840 1324.310 285.100 1324.630 ;
        RECT 2900.860 1324.310 2901.120 1324.630 ;
        RECT 2900.920 1319.725 2901.060 1324.310 ;
        RECT 2900.850 1319.355 2901.130 1319.725 ;
      LAYER via2 ;
        RECT 284.830 1683.880 285.110 1684.160 ;
        RECT 2900.850 1319.400 2901.130 1319.680 ;
      LAYER met3 ;
        RECT 284.805 1684.170 285.135 1684.185 ;
        RECT 300.000 1684.170 304.000 1684.240 ;
        RECT 284.805 1683.870 304.000 1684.170 ;
        RECT 284.805 1683.855 285.135 1683.870 ;
        RECT 300.000 1683.640 304.000 1683.870 ;
        RECT 2900.825 1319.690 2901.155 1319.705 ;
        RECT 2917.600 1319.690 2924.800 1320.140 ;
        RECT 2900.825 1319.390 2924.800 1319.690 ;
        RECT 2900.825 1319.375 2901.155 1319.390 ;
        RECT 2917.600 1318.940 2924.800 1319.390 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 283.430 1503.720 283.750 1503.780 ;
        RECT 2901.750 1503.720 2902.070 1503.780 ;
        RECT 283.430 1503.580 2902.070 1503.720 ;
        RECT 283.430 1503.520 283.750 1503.580 ;
        RECT 2901.750 1503.520 2902.070 1503.580 ;
      LAYER via ;
        RECT 283.460 1503.520 283.720 1503.780 ;
        RECT 2901.780 1503.520 2902.040 1503.780 ;
      LAYER met2 ;
        RECT 283.450 1715.115 283.730 1715.485 ;
        RECT 283.520 1503.810 283.660 1715.115 ;
        RECT 2901.770 1553.955 2902.050 1554.325 ;
        RECT 2901.840 1503.810 2901.980 1553.955 ;
        RECT 283.460 1503.490 283.720 1503.810 ;
        RECT 2901.780 1503.490 2902.040 1503.810 ;
      LAYER via2 ;
        RECT 283.450 1715.160 283.730 1715.440 ;
        RECT 2901.770 1554.000 2902.050 1554.280 ;
      LAYER met3 ;
        RECT 283.425 1715.450 283.755 1715.465 ;
        RECT 300.000 1715.450 304.000 1715.520 ;
        RECT 283.425 1715.150 304.000 1715.450 ;
        RECT 283.425 1715.135 283.755 1715.150 ;
        RECT 300.000 1714.920 304.000 1715.150 ;
        RECT 2901.745 1554.290 2902.075 1554.305 ;
        RECT 2917.600 1554.290 2924.800 1554.740 ;
        RECT 2901.745 1553.990 2924.800 1554.290 ;
        RECT 2901.745 1553.975 2902.075 1553.990 ;
        RECT 2917.600 1553.540 2924.800 1553.990 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2884.270 1780.480 2884.590 1780.540 ;
        RECT 2897.610 1780.480 2897.930 1780.540 ;
        RECT 2884.270 1780.340 2897.930 1780.480 ;
        RECT 2884.270 1780.280 2884.590 1780.340 ;
        RECT 2897.610 1780.280 2897.930 1780.340 ;
        RECT 2859.890 1767.220 2860.210 1767.280 ;
        RECT 2884.270 1767.220 2884.590 1767.280 ;
        RECT 2859.890 1767.080 2884.590 1767.220 ;
        RECT 2859.890 1767.020 2860.210 1767.080 ;
        RECT 2884.270 1767.020 2884.590 1767.080 ;
        RECT 2822.170 1749.200 2822.490 1749.260 ;
        RECT 2859.890 1749.200 2860.210 1749.260 ;
        RECT 2822.170 1749.060 2860.210 1749.200 ;
        RECT 2822.170 1749.000 2822.490 1749.060 ;
        RECT 2859.890 1749.000 2860.210 1749.060 ;
        RECT 2808.370 1737.300 2808.690 1737.360 ;
        RECT 2822.170 1737.300 2822.490 1737.360 ;
        RECT 2808.370 1737.160 2822.490 1737.300 ;
        RECT 2808.370 1737.100 2808.690 1737.160 ;
        RECT 2822.170 1737.100 2822.490 1737.160 ;
        RECT 2808.370 1718.260 2808.690 1718.320 ;
        RECT 2805.700 1718.120 2808.690 1718.260 ;
        RECT 2792.270 1717.920 2792.590 1717.980 ;
        RECT 2805.700 1717.920 2805.840 1718.120 ;
        RECT 2808.370 1718.060 2808.690 1718.120 ;
        RECT 2792.270 1717.780 2805.840 1717.920 ;
        RECT 2792.270 1717.720 2792.590 1717.780 ;
        RECT 2766.970 1704.660 2767.290 1704.720 ;
        RECT 2792.270 1704.660 2792.590 1704.720 ;
        RECT 2766.970 1704.520 2792.590 1704.660 ;
        RECT 2766.970 1704.460 2767.290 1704.520 ;
        RECT 2792.270 1704.460 2792.590 1704.520 ;
        RECT 2756.850 1690.720 2757.170 1690.780 ;
        RECT 2766.970 1690.720 2767.290 1690.780 ;
        RECT 2756.850 1690.580 2767.290 1690.720 ;
        RECT 2756.850 1690.520 2757.170 1690.580 ;
        RECT 2766.970 1690.520 2767.290 1690.580 ;
        RECT 286.650 1652.640 286.970 1652.700 ;
        RECT 288.490 1652.640 288.810 1652.700 ;
        RECT 286.650 1652.500 288.810 1652.640 ;
        RECT 286.650 1652.440 286.970 1652.500 ;
        RECT 288.490 1652.440 288.810 1652.500 ;
        RECT 2746.730 1640.740 2747.050 1640.800 ;
        RECT 2756.850 1640.740 2757.170 1640.800 ;
        RECT 2746.730 1640.600 2757.170 1640.740 ;
        RECT 2746.730 1640.540 2747.050 1640.600 ;
        RECT 2756.850 1640.540 2757.170 1640.600 ;
        RECT 288.490 1635.300 288.810 1635.360 ;
        RECT 294.930 1635.300 295.250 1635.360 ;
        RECT 288.490 1635.160 295.250 1635.300 ;
        RECT 288.490 1635.100 288.810 1635.160 ;
        RECT 294.930 1635.100 295.250 1635.160 ;
        RECT 2725.570 1621.700 2725.890 1621.760 ;
        RECT 2746.730 1621.700 2747.050 1621.760 ;
        RECT 2725.570 1621.560 2747.050 1621.700 ;
        RECT 2725.570 1621.500 2725.890 1621.560 ;
        RECT 2746.730 1621.500 2747.050 1621.560 ;
        RECT 2714.990 1600.960 2715.310 1601.020 ;
        RECT 2725.570 1600.960 2725.890 1601.020 ;
        RECT 2714.990 1600.820 2725.890 1600.960 ;
        RECT 2714.990 1600.760 2715.310 1600.820 ;
        RECT 2725.570 1600.760 2725.890 1600.820 ;
        RECT 2677.270 1555.740 2677.590 1555.800 ;
        RECT 2714.990 1555.740 2715.310 1555.800 ;
        RECT 2677.270 1555.600 2715.310 1555.740 ;
        RECT 2677.270 1555.540 2677.590 1555.600 ;
        RECT 2714.990 1555.540 2715.310 1555.600 ;
        RECT 2677.270 1545.880 2677.590 1545.940 ;
        RECT 2663.560 1545.740 2677.590 1545.880 ;
        RECT 2661.630 1545.540 2661.950 1545.600 ;
        RECT 2663.560 1545.540 2663.700 1545.740 ;
        RECT 2677.270 1545.680 2677.590 1545.740 ;
        RECT 2661.630 1545.400 2663.700 1545.540 ;
        RECT 2661.630 1545.340 2661.950 1545.400 ;
        RECT 294.930 1501.340 295.250 1501.400 ;
        RECT 2661.630 1501.340 2661.950 1501.400 ;
        RECT 294.930 1501.200 2661.950 1501.340 ;
        RECT 294.930 1501.140 295.250 1501.200 ;
        RECT 2661.630 1501.140 2661.950 1501.200 ;
      LAYER via ;
        RECT 2884.300 1780.280 2884.560 1780.540 ;
        RECT 2897.640 1780.280 2897.900 1780.540 ;
        RECT 2859.920 1767.020 2860.180 1767.280 ;
        RECT 2884.300 1767.020 2884.560 1767.280 ;
        RECT 2822.200 1749.000 2822.460 1749.260 ;
        RECT 2859.920 1749.000 2860.180 1749.260 ;
        RECT 2808.400 1737.100 2808.660 1737.360 ;
        RECT 2822.200 1737.100 2822.460 1737.360 ;
        RECT 2792.300 1717.720 2792.560 1717.980 ;
        RECT 2808.400 1718.060 2808.660 1718.320 ;
        RECT 2767.000 1704.460 2767.260 1704.720 ;
        RECT 2792.300 1704.460 2792.560 1704.720 ;
        RECT 2756.880 1690.520 2757.140 1690.780 ;
        RECT 2767.000 1690.520 2767.260 1690.780 ;
        RECT 286.680 1652.440 286.940 1652.700 ;
        RECT 288.520 1652.440 288.780 1652.700 ;
        RECT 2746.760 1640.540 2747.020 1640.800 ;
        RECT 2756.880 1640.540 2757.140 1640.800 ;
        RECT 288.520 1635.100 288.780 1635.360 ;
        RECT 294.960 1635.100 295.220 1635.360 ;
        RECT 2725.600 1621.500 2725.860 1621.760 ;
        RECT 2746.760 1621.500 2747.020 1621.760 ;
        RECT 2715.020 1600.760 2715.280 1601.020 ;
        RECT 2725.600 1600.760 2725.860 1601.020 ;
        RECT 2677.300 1555.540 2677.560 1555.800 ;
        RECT 2715.020 1555.540 2715.280 1555.800 ;
        RECT 2661.660 1545.340 2661.920 1545.600 ;
        RECT 2677.300 1545.680 2677.560 1545.940 ;
        RECT 294.960 1501.140 295.220 1501.400 ;
        RECT 2661.660 1501.140 2661.920 1501.400 ;
      LAYER met2 ;
        RECT 2897.630 1789.235 2897.910 1789.605 ;
        RECT 2897.700 1780.570 2897.840 1789.235 ;
        RECT 2884.300 1780.250 2884.560 1780.570 ;
        RECT 2897.640 1780.250 2897.900 1780.570 ;
        RECT 2884.360 1767.310 2884.500 1780.250 ;
        RECT 2859.920 1766.990 2860.180 1767.310 ;
        RECT 2884.300 1766.990 2884.560 1767.310 ;
        RECT 2859.980 1749.290 2860.120 1766.990 ;
        RECT 2822.200 1748.970 2822.460 1749.290 ;
        RECT 2859.920 1748.970 2860.180 1749.290 ;
        RECT 286.670 1747.075 286.950 1747.445 ;
        RECT 286.740 1652.730 286.880 1747.075 ;
        RECT 2822.260 1737.390 2822.400 1748.970 ;
        RECT 2808.400 1737.070 2808.660 1737.390 ;
        RECT 2822.200 1737.070 2822.460 1737.390 ;
        RECT 2808.460 1718.350 2808.600 1737.070 ;
        RECT 2808.400 1718.030 2808.660 1718.350 ;
        RECT 2792.300 1717.690 2792.560 1718.010 ;
        RECT 2792.360 1704.750 2792.500 1717.690 ;
        RECT 2767.000 1704.430 2767.260 1704.750 ;
        RECT 2792.300 1704.430 2792.560 1704.750 ;
        RECT 2767.060 1690.810 2767.200 1704.430 ;
        RECT 2756.880 1690.490 2757.140 1690.810 ;
        RECT 2767.000 1690.490 2767.260 1690.810 ;
        RECT 286.680 1652.410 286.940 1652.730 ;
        RECT 288.520 1652.410 288.780 1652.730 ;
        RECT 288.580 1635.390 288.720 1652.410 ;
        RECT 2756.940 1640.830 2757.080 1690.490 ;
        RECT 2746.760 1640.510 2747.020 1640.830 ;
        RECT 2756.880 1640.510 2757.140 1640.830 ;
        RECT 288.520 1635.070 288.780 1635.390 ;
        RECT 294.960 1635.070 295.220 1635.390 ;
        RECT 295.020 1501.430 295.160 1635.070 ;
        RECT 2746.820 1621.790 2746.960 1640.510 ;
        RECT 2725.600 1621.470 2725.860 1621.790 ;
        RECT 2746.760 1621.470 2747.020 1621.790 ;
        RECT 2725.660 1601.050 2725.800 1621.470 ;
        RECT 2715.020 1600.730 2715.280 1601.050 ;
        RECT 2725.600 1600.730 2725.860 1601.050 ;
        RECT 2715.080 1555.830 2715.220 1600.730 ;
        RECT 2677.300 1555.510 2677.560 1555.830 ;
        RECT 2715.020 1555.510 2715.280 1555.830 ;
        RECT 2677.360 1545.970 2677.500 1555.510 ;
        RECT 2677.300 1545.650 2677.560 1545.970 ;
        RECT 2661.660 1545.310 2661.920 1545.630 ;
        RECT 2661.720 1501.430 2661.860 1545.310 ;
        RECT 294.960 1501.110 295.220 1501.430 ;
        RECT 2661.660 1501.110 2661.920 1501.430 ;
      LAYER via2 ;
        RECT 2897.630 1789.280 2897.910 1789.560 ;
        RECT 286.670 1747.120 286.950 1747.400 ;
      LAYER met3 ;
        RECT 2897.605 1789.570 2897.935 1789.585 ;
        RECT 2917.600 1789.570 2924.800 1790.020 ;
        RECT 2897.605 1789.270 2924.800 1789.570 ;
        RECT 2897.605 1789.255 2897.935 1789.270 ;
        RECT 2917.600 1788.820 2924.800 1789.270 ;
        RECT 286.645 1747.410 286.975 1747.425 ;
        RECT 300.000 1747.410 304.000 1747.480 ;
        RECT 286.645 1747.110 304.000 1747.410 ;
        RECT 286.645 1747.095 286.975 1747.110 ;
        RECT 300.000 1746.880 304.000 1747.110 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2887.490 2001.140 2887.810 2001.200 ;
        RECT 2904.510 2001.140 2904.830 2001.200 ;
        RECT 2887.490 2001.000 2904.830 2001.140 ;
        RECT 2887.490 2000.940 2887.810 2001.000 ;
        RECT 2904.510 2000.940 2904.830 2001.000 ;
        RECT 2873.690 1773.680 2874.010 1773.740 ;
        RECT 2887.490 1773.680 2887.810 1773.740 ;
        RECT 2873.690 1773.540 2887.810 1773.680 ;
        RECT 2873.690 1773.480 2874.010 1773.540 ;
        RECT 2887.490 1773.480 2887.810 1773.540 ;
        RECT 2866.790 1737.300 2867.110 1737.360 ;
        RECT 2873.690 1737.300 2874.010 1737.360 ;
        RECT 2866.790 1737.160 2874.010 1737.300 ;
        RECT 2866.790 1737.100 2867.110 1737.160 ;
        RECT 2873.690 1737.100 2874.010 1737.160 ;
        RECT 285.730 1658.080 286.050 1658.140 ;
        RECT 294.010 1658.080 294.330 1658.140 ;
        RECT 285.730 1657.940 294.330 1658.080 ;
        RECT 285.730 1657.880 286.050 1657.940 ;
        RECT 294.010 1657.880 294.330 1657.940 ;
        RECT 2866.790 1559.480 2867.110 1559.540 ;
        RECT 2849.860 1559.340 2867.110 1559.480 ;
        RECT 2839.650 1559.140 2839.970 1559.200 ;
        RECT 2849.860 1559.140 2850.000 1559.340 ;
        RECT 2866.790 1559.280 2867.110 1559.340 ;
        RECT 2839.650 1559.000 2850.000 1559.140 ;
        RECT 2839.650 1558.940 2839.970 1559.000 ;
        RECT 2815.270 1549.960 2815.590 1550.020 ;
        RECT 2839.650 1549.960 2839.970 1550.020 ;
        RECT 2815.270 1549.820 2839.970 1549.960 ;
        RECT 2815.270 1549.760 2815.590 1549.820 ;
        RECT 2839.650 1549.760 2839.970 1549.820 ;
        RECT 2815.270 1539.080 2815.590 1539.140 ;
        RECT 2808.460 1538.940 2815.590 1539.080 ;
        RECT 2787.670 1538.740 2787.990 1538.800 ;
        RECT 2808.460 1538.740 2808.600 1538.940 ;
        RECT 2815.270 1538.880 2815.590 1538.940 ;
        RECT 2787.670 1538.600 2808.600 1538.740 ;
        RECT 2787.670 1538.540 2787.990 1538.600 ;
        RECT 294.010 1517.320 294.330 1517.380 ;
        RECT 303.210 1517.320 303.530 1517.380 ;
        RECT 294.010 1517.180 303.530 1517.320 ;
        RECT 294.010 1517.120 294.330 1517.180 ;
        RECT 303.210 1517.120 303.530 1517.180 ;
        RECT 2766.970 1513.920 2767.290 1513.980 ;
        RECT 2787.670 1513.920 2787.990 1513.980 ;
        RECT 2766.970 1513.780 2787.990 1513.920 ;
        RECT 2766.970 1513.720 2767.290 1513.780 ;
        RECT 2787.670 1513.720 2787.990 1513.780 ;
        RECT 303.210 1502.700 303.530 1502.760 ;
        RECT 2766.970 1502.700 2767.290 1502.760 ;
        RECT 303.210 1502.560 2767.290 1502.700 ;
        RECT 303.210 1502.500 303.530 1502.560 ;
        RECT 2766.970 1502.500 2767.290 1502.560 ;
      LAYER via ;
        RECT 2887.520 2000.940 2887.780 2001.200 ;
        RECT 2904.540 2000.940 2904.800 2001.200 ;
        RECT 2873.720 1773.480 2873.980 1773.740 ;
        RECT 2887.520 1773.480 2887.780 1773.740 ;
        RECT 2866.820 1737.100 2867.080 1737.360 ;
        RECT 2873.720 1737.100 2873.980 1737.360 ;
        RECT 285.760 1657.880 286.020 1658.140 ;
        RECT 294.040 1657.880 294.300 1658.140 ;
        RECT 2839.680 1558.940 2839.940 1559.200 ;
        RECT 2866.820 1559.280 2867.080 1559.540 ;
        RECT 2815.300 1549.760 2815.560 1550.020 ;
        RECT 2839.680 1549.760 2839.940 1550.020 ;
        RECT 2787.700 1538.540 2787.960 1538.800 ;
        RECT 2815.300 1538.880 2815.560 1539.140 ;
        RECT 294.040 1517.120 294.300 1517.380 ;
        RECT 303.240 1517.120 303.500 1517.380 ;
        RECT 2767.000 1513.720 2767.260 1513.980 ;
        RECT 2787.700 1513.720 2787.960 1513.980 ;
        RECT 303.240 1502.500 303.500 1502.760 ;
        RECT 2767.000 1502.500 2767.260 1502.760 ;
      LAYER met2 ;
        RECT 2904.530 2023.835 2904.810 2024.205 ;
        RECT 2904.600 2001.230 2904.740 2023.835 ;
        RECT 2887.520 2000.910 2887.780 2001.230 ;
        RECT 2904.540 2000.910 2904.800 2001.230 ;
        RECT 285.750 1778.355 286.030 1778.725 ;
        RECT 285.820 1658.170 285.960 1778.355 ;
        RECT 2887.580 1773.770 2887.720 2000.910 ;
        RECT 2873.720 1773.450 2873.980 1773.770 ;
        RECT 2887.520 1773.450 2887.780 1773.770 ;
        RECT 2873.780 1737.390 2873.920 1773.450 ;
        RECT 2866.820 1737.070 2867.080 1737.390 ;
        RECT 2873.720 1737.070 2873.980 1737.390 ;
        RECT 285.760 1657.850 286.020 1658.170 ;
        RECT 294.040 1657.850 294.300 1658.170 ;
        RECT 294.100 1517.410 294.240 1657.850 ;
        RECT 2866.880 1559.570 2867.020 1737.070 ;
        RECT 2866.820 1559.250 2867.080 1559.570 ;
        RECT 2839.680 1558.910 2839.940 1559.230 ;
        RECT 2839.740 1550.050 2839.880 1558.910 ;
        RECT 2815.300 1549.730 2815.560 1550.050 ;
        RECT 2839.680 1549.730 2839.940 1550.050 ;
        RECT 2815.360 1539.170 2815.500 1549.730 ;
        RECT 2815.300 1538.850 2815.560 1539.170 ;
        RECT 2787.700 1538.510 2787.960 1538.830 ;
        RECT 294.040 1517.090 294.300 1517.410 ;
        RECT 303.240 1517.090 303.500 1517.410 ;
        RECT 303.300 1502.790 303.440 1517.090 ;
        RECT 2787.760 1514.010 2787.900 1538.510 ;
        RECT 2767.000 1513.690 2767.260 1514.010 ;
        RECT 2787.700 1513.690 2787.960 1514.010 ;
        RECT 2767.060 1502.790 2767.200 1513.690 ;
        RECT 303.240 1502.470 303.500 1502.790 ;
        RECT 2767.000 1502.470 2767.260 1502.790 ;
      LAYER via2 ;
        RECT 2904.530 2023.880 2904.810 2024.160 ;
        RECT 285.750 1778.400 286.030 1778.680 ;
      LAYER met3 ;
        RECT 2904.505 2024.170 2904.835 2024.185 ;
        RECT 2917.600 2024.170 2924.800 2024.620 ;
        RECT 2904.505 2023.870 2924.800 2024.170 ;
        RECT 2904.505 2023.855 2904.835 2023.870 ;
        RECT 2917.600 2023.420 2924.800 2023.870 ;
        RECT 285.725 1778.690 286.055 1778.705 ;
        RECT 300.000 1778.690 304.000 1778.760 ;
        RECT 285.725 1778.390 304.000 1778.690 ;
        RECT 285.725 1778.375 286.055 1778.390 ;
        RECT 300.000 1778.160 304.000 1778.390 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2893.010 2201.400 2893.330 2201.460 ;
        RECT 2901.290 2201.400 2901.610 2201.460 ;
        RECT 2893.010 2201.260 2901.610 2201.400 ;
        RECT 2893.010 2201.200 2893.330 2201.260 ;
        RECT 2901.290 2201.200 2901.610 2201.260 ;
        RECT 2880.590 2194.600 2880.910 2194.660 ;
        RECT 2893.010 2194.600 2893.330 2194.660 ;
        RECT 2880.590 2194.460 2893.330 2194.600 ;
        RECT 2880.590 2194.400 2880.910 2194.460 ;
        RECT 2893.010 2194.400 2893.330 2194.460 ;
        RECT 2852.990 2134.080 2853.310 2134.140 ;
        RECT 2880.590 2134.080 2880.910 2134.140 ;
        RECT 2852.990 2133.940 2880.910 2134.080 ;
        RECT 2852.990 2133.880 2853.310 2133.940 ;
        RECT 2880.590 2133.880 2880.910 2133.940 ;
        RECT 2846.090 1973.260 2846.410 1973.320 ;
        RECT 2852.990 1973.260 2853.310 1973.320 ;
        RECT 2846.090 1973.120 2853.310 1973.260 ;
        RECT 2846.090 1973.060 2846.410 1973.120 ;
        RECT 2852.990 1973.060 2853.310 1973.120 ;
        RECT 2832.290 1858.680 2832.610 1858.740 ;
        RECT 2846.090 1858.680 2846.410 1858.740 ;
        RECT 2832.290 1858.540 2846.410 1858.680 ;
        RECT 2832.290 1858.480 2832.610 1858.540 ;
        RECT 2846.090 1858.480 2846.410 1858.540 ;
        RECT 285.270 1697.180 285.590 1697.240 ;
        RECT 293.550 1697.180 293.870 1697.240 ;
        RECT 285.270 1697.040 293.870 1697.180 ;
        RECT 285.270 1696.980 285.590 1697.040 ;
        RECT 293.550 1696.980 293.870 1697.040 ;
        RECT 2817.110 1693.440 2817.430 1693.500 ;
        RECT 2832.290 1693.440 2832.610 1693.500 ;
        RECT 2817.110 1693.300 2832.610 1693.440 ;
        RECT 2817.110 1693.240 2817.430 1693.300 ;
        RECT 2832.290 1693.240 2832.610 1693.300 ;
        RECT 2808.830 1683.240 2809.150 1683.300 ;
        RECT 2817.110 1683.240 2817.430 1683.300 ;
        RECT 2808.830 1683.100 2817.430 1683.240 ;
        RECT 2808.830 1683.040 2809.150 1683.100 ;
        RECT 2817.110 1683.040 2817.430 1683.100 ;
        RECT 2794.110 1669.980 2794.430 1670.040 ;
        RECT 2808.830 1669.980 2809.150 1670.040 ;
        RECT 2794.110 1669.840 2809.150 1669.980 ;
        RECT 2794.110 1669.780 2794.430 1669.840 ;
        RECT 2808.830 1669.780 2809.150 1669.840 ;
        RECT 2783.990 1657.400 2784.310 1657.460 ;
        RECT 2794.110 1657.400 2794.430 1657.460 ;
        RECT 2783.990 1657.260 2794.430 1657.400 ;
        RECT 2783.990 1657.200 2784.310 1657.260 ;
        RECT 2794.110 1657.200 2794.430 1657.260 ;
        RECT 2766.970 1621.700 2767.290 1621.760 ;
        RECT 2783.990 1621.700 2784.310 1621.760 ;
        RECT 2766.970 1621.560 2784.310 1621.700 ;
        RECT 2766.970 1621.500 2767.290 1621.560 ;
        RECT 2783.990 1621.500 2784.310 1621.560 ;
        RECT 2749.490 1597.560 2749.810 1597.620 ;
        RECT 2766.970 1597.560 2767.290 1597.620 ;
        RECT 2749.490 1597.420 2767.290 1597.560 ;
        RECT 2749.490 1597.360 2749.810 1597.420 ;
        RECT 2766.970 1597.360 2767.290 1597.420 ;
        RECT 2725.570 1555.060 2725.890 1555.120 ;
        RECT 2749.490 1555.060 2749.810 1555.120 ;
        RECT 2725.570 1554.920 2749.810 1555.060 ;
        RECT 2725.570 1554.860 2725.890 1554.920 ;
        RECT 2749.490 1554.860 2749.810 1554.920 ;
        RECT 2698.430 1543.500 2698.750 1543.560 ;
        RECT 2725.570 1543.500 2725.890 1543.560 ;
        RECT 2698.430 1543.360 2725.890 1543.500 ;
        RECT 2698.430 1543.300 2698.750 1543.360 ;
        RECT 2725.570 1543.300 2725.890 1543.360 ;
        RECT 293.550 1521.740 293.870 1521.800 ;
        RECT 297.690 1521.740 298.010 1521.800 ;
        RECT 293.550 1521.600 298.010 1521.740 ;
        RECT 293.550 1521.540 293.870 1521.600 ;
        RECT 297.690 1521.540 298.010 1521.600 ;
        RECT 2684.170 1505.080 2684.490 1505.140 ;
        RECT 2698.430 1505.080 2698.750 1505.140 ;
        RECT 2684.170 1504.940 2698.750 1505.080 ;
        RECT 2684.170 1504.880 2684.490 1504.940 ;
        RECT 2698.430 1504.880 2698.750 1504.940 ;
        RECT 297.690 1501.680 298.010 1501.740 ;
        RECT 2684.170 1501.680 2684.490 1501.740 ;
        RECT 297.690 1501.540 2684.490 1501.680 ;
        RECT 297.690 1501.480 298.010 1501.540 ;
        RECT 2684.170 1501.480 2684.490 1501.540 ;
      LAYER via ;
        RECT 2893.040 2201.200 2893.300 2201.460 ;
        RECT 2901.320 2201.200 2901.580 2201.460 ;
        RECT 2880.620 2194.400 2880.880 2194.660 ;
        RECT 2893.040 2194.400 2893.300 2194.660 ;
        RECT 2853.020 2133.880 2853.280 2134.140 ;
        RECT 2880.620 2133.880 2880.880 2134.140 ;
        RECT 2846.120 1973.060 2846.380 1973.320 ;
        RECT 2853.020 1973.060 2853.280 1973.320 ;
        RECT 2832.320 1858.480 2832.580 1858.740 ;
        RECT 2846.120 1858.480 2846.380 1858.740 ;
        RECT 285.300 1696.980 285.560 1697.240 ;
        RECT 293.580 1696.980 293.840 1697.240 ;
        RECT 2817.140 1693.240 2817.400 1693.500 ;
        RECT 2832.320 1693.240 2832.580 1693.500 ;
        RECT 2808.860 1683.040 2809.120 1683.300 ;
        RECT 2817.140 1683.040 2817.400 1683.300 ;
        RECT 2794.140 1669.780 2794.400 1670.040 ;
        RECT 2808.860 1669.780 2809.120 1670.040 ;
        RECT 2784.020 1657.200 2784.280 1657.460 ;
        RECT 2794.140 1657.200 2794.400 1657.460 ;
        RECT 2767.000 1621.500 2767.260 1621.760 ;
        RECT 2784.020 1621.500 2784.280 1621.760 ;
        RECT 2749.520 1597.360 2749.780 1597.620 ;
        RECT 2767.000 1597.360 2767.260 1597.620 ;
        RECT 2725.600 1554.860 2725.860 1555.120 ;
        RECT 2749.520 1554.860 2749.780 1555.120 ;
        RECT 2698.460 1543.300 2698.720 1543.560 ;
        RECT 2725.600 1543.300 2725.860 1543.560 ;
        RECT 293.580 1521.540 293.840 1521.800 ;
        RECT 297.720 1521.540 297.980 1521.800 ;
        RECT 2684.200 1504.880 2684.460 1505.140 ;
        RECT 2698.460 1504.880 2698.720 1505.140 ;
        RECT 297.720 1501.480 297.980 1501.740 ;
        RECT 2684.200 1501.480 2684.460 1501.740 ;
      LAYER met2 ;
        RECT 2901.310 2258.435 2901.590 2258.805 ;
        RECT 2901.380 2201.490 2901.520 2258.435 ;
        RECT 2893.040 2201.170 2893.300 2201.490 ;
        RECT 2901.320 2201.170 2901.580 2201.490 ;
        RECT 2893.100 2194.690 2893.240 2201.170 ;
        RECT 2880.620 2194.370 2880.880 2194.690 ;
        RECT 2893.040 2194.370 2893.300 2194.690 ;
        RECT 2880.680 2134.170 2880.820 2194.370 ;
        RECT 2853.020 2133.850 2853.280 2134.170 ;
        RECT 2880.620 2133.850 2880.880 2134.170 ;
        RECT 2853.080 1973.350 2853.220 2133.850 ;
        RECT 2846.120 1973.030 2846.380 1973.350 ;
        RECT 2853.020 1973.030 2853.280 1973.350 ;
        RECT 2846.180 1858.770 2846.320 1973.030 ;
        RECT 2832.320 1858.450 2832.580 1858.770 ;
        RECT 2846.120 1858.450 2846.380 1858.770 ;
        RECT 285.290 1809.635 285.570 1810.005 ;
        RECT 285.360 1697.270 285.500 1809.635 ;
        RECT 285.300 1696.950 285.560 1697.270 ;
        RECT 293.580 1696.950 293.840 1697.270 ;
        RECT 293.640 1521.830 293.780 1696.950 ;
        RECT 2832.380 1693.530 2832.520 1858.450 ;
        RECT 2817.140 1693.210 2817.400 1693.530 ;
        RECT 2832.320 1693.210 2832.580 1693.530 ;
        RECT 2817.200 1683.330 2817.340 1693.210 ;
        RECT 2808.860 1683.010 2809.120 1683.330 ;
        RECT 2817.140 1683.010 2817.400 1683.330 ;
        RECT 2808.920 1670.070 2809.060 1683.010 ;
        RECT 2794.140 1669.750 2794.400 1670.070 ;
        RECT 2808.860 1669.750 2809.120 1670.070 ;
        RECT 2794.200 1657.490 2794.340 1669.750 ;
        RECT 2784.020 1657.170 2784.280 1657.490 ;
        RECT 2794.140 1657.170 2794.400 1657.490 ;
        RECT 2784.080 1621.790 2784.220 1657.170 ;
        RECT 2767.000 1621.470 2767.260 1621.790 ;
        RECT 2784.020 1621.470 2784.280 1621.790 ;
        RECT 2767.060 1597.650 2767.200 1621.470 ;
        RECT 2749.520 1597.330 2749.780 1597.650 ;
        RECT 2767.000 1597.330 2767.260 1597.650 ;
        RECT 2749.580 1555.150 2749.720 1597.330 ;
        RECT 2725.600 1554.830 2725.860 1555.150 ;
        RECT 2749.520 1554.830 2749.780 1555.150 ;
        RECT 2725.660 1543.590 2725.800 1554.830 ;
        RECT 2698.460 1543.270 2698.720 1543.590 ;
        RECT 2725.600 1543.270 2725.860 1543.590 ;
        RECT 293.580 1521.510 293.840 1521.830 ;
        RECT 297.720 1521.510 297.980 1521.830 ;
        RECT 297.780 1501.770 297.920 1521.510 ;
        RECT 2698.520 1505.170 2698.660 1543.270 ;
        RECT 2684.200 1504.850 2684.460 1505.170 ;
        RECT 2698.460 1504.850 2698.720 1505.170 ;
        RECT 2684.260 1501.770 2684.400 1504.850 ;
        RECT 297.720 1501.450 297.980 1501.770 ;
        RECT 2684.200 1501.450 2684.460 1501.770 ;
      LAYER via2 ;
        RECT 2901.310 2258.480 2901.590 2258.760 ;
        RECT 285.290 1809.680 285.570 1809.960 ;
      LAYER met3 ;
        RECT 2901.285 2258.770 2901.615 2258.785 ;
        RECT 2917.600 2258.770 2924.800 2259.220 ;
        RECT 2901.285 2258.470 2924.800 2258.770 ;
        RECT 2901.285 2258.455 2901.615 2258.470 ;
        RECT 2917.600 2258.020 2924.800 2258.470 ;
        RECT 285.265 1809.970 285.595 1809.985 ;
        RECT 300.000 1809.970 304.000 1810.040 ;
        RECT 285.265 1809.670 304.000 1809.970 ;
        RECT 285.265 1809.655 285.595 1809.670 ;
        RECT 300.000 1809.440 304.000 1809.670 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 688.230 25.740 688.550 25.800 ;
        RECT 1331.770 25.740 1332.090 25.800 ;
        RECT 688.230 25.600 1332.090 25.740 ;
        RECT 688.230 25.540 688.550 25.600 ;
        RECT 1331.770 25.540 1332.090 25.600 ;
        RECT 633.030 24.720 633.350 24.780 ;
        RECT 633.030 24.580 637.400 24.720 ;
        RECT 633.030 24.520 633.350 24.580 ;
        RECT 637.260 24.380 637.400 24.580 ;
        RECT 687.310 24.380 687.630 24.440 ;
        RECT 637.260 24.240 687.630 24.380 ;
        RECT 687.310 24.180 687.630 24.240 ;
      LAYER via ;
        RECT 688.260 25.540 688.520 25.800 ;
        RECT 1331.800 25.540 1332.060 25.800 ;
        RECT 633.060 24.520 633.320 24.780 ;
        RECT 687.340 24.180 687.600 24.440 ;
      LAYER met2 ;
        RECT 1336.010 1500.490 1336.290 1504.000 ;
        RECT 1331.860 1500.350 1336.290 1500.490 ;
        RECT 1331.860 25.830 1332.000 1500.350 ;
        RECT 1336.010 1500.000 1336.290 1500.350 ;
        RECT 688.260 25.510 688.520 25.830 ;
        RECT 1331.800 25.510 1332.060 25.830 ;
        RECT 633.060 24.490 633.320 24.810 ;
        RECT 633.120 2.400 633.260 24.490 ;
        RECT 687.340 24.150 687.600 24.470 ;
        RECT 687.400 23.530 687.540 24.150 ;
        RECT 688.320 23.530 688.460 25.510 ;
        RECT 687.400 23.390 688.460 23.530 ;
        RECT 632.910 -4.800 633.470 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2417.250 -4.800 2417.810 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2434.730 -4.800 2435.290 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2452.670 -4.800 2453.230 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2470.610 -4.800 2471.170 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2488.550 -4.800 2489.110 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2506.030 -4.800 2506.590 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2523.970 -4.800 2524.530 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2541.910 -4.800 2542.470 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2559.850 -4.800 2560.410 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2577.790 -4.800 2578.350 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 811.390 -4.800 811.950 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2595.270 -4.800 2595.830 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2613.210 -4.800 2613.770 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2631.150 -4.800 2631.710 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2649.090 -4.800 2649.650 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2667.030 -4.800 2667.590 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2684.510 -4.800 2685.070 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2702.450 -4.800 2703.010 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2720.390 -4.800 2720.950 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2738.330 -4.800 2738.890 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2755.810 -4.800 2756.370 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 829.330 -4.800 829.890 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2773.750 -4.800 2774.310 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2791.690 -4.800 2792.250 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2809.630 -4.800 2810.190 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2827.570 -4.800 2828.130 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2845.050 -4.800 2845.610 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2862.990 -4.800 2863.550 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2880.930 -4.800 2881.490 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 846.810 -4.800 847.370 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 864.750 -4.800 865.310 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 882.690 -4.800 883.250 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 900.630 -4.800 901.190 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 918.570 -4.800 919.130 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 936.050 -4.800 936.610 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1359.370 25.400 1359.690 25.460 ;
        RECT 686.480 25.260 1359.690 25.400 ;
        RECT 650.970 25.060 651.290 25.120 ;
        RECT 686.480 25.060 686.620 25.260 ;
        RECT 1359.370 25.200 1359.690 25.260 ;
        RECT 650.970 24.920 686.620 25.060 ;
        RECT 650.970 24.860 651.290 24.920 ;
      LAYER via ;
        RECT 651.000 24.860 651.260 25.120 ;
        RECT 1359.400 25.200 1359.660 25.460 ;
      LAYER met2 ;
        RECT 1365.450 1500.490 1365.730 1504.000 ;
        RECT 1359.460 1500.350 1365.730 1500.490 ;
        RECT 1359.460 25.490 1359.600 1500.350 ;
        RECT 1365.450 1500.000 1365.730 1500.350 ;
        RECT 1359.400 25.170 1359.660 25.490 ;
        RECT 651.000 24.830 651.260 25.150 ;
        RECT 651.060 2.400 651.200 24.830 ;
        RECT 650.850 -4.800 651.410 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 989.870 -4.800 990.430 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1043.230 -4.800 1043.790 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1061.170 -4.800 1061.730 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1079.110 -4.800 1079.670 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1096.590 -4.800 1097.150 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1114.530 -4.800 1115.090 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1132.470 -4.800 1133.030 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1150.410 -4.800 1150.970 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 668.790 -4.800 669.350 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1168.350 -4.800 1168.910 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1185.830 -4.800 1186.390 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1203.770 -4.800 1204.330 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1221.710 -4.800 1222.270 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1239.650 -4.800 1240.210 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 -4.800 1257.690 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1275.070 -4.800 1275.630 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1293.010 -4.800 1293.570 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1310.950 -4.800 1311.510 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1328.890 -4.800 1329.450 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 686.270 -4.800 686.830 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1346.370 -4.800 1346.930 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1364.310 -4.800 1364.870 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1382.250 -4.800 1382.810 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1400.190 -4.800 1400.750 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1418.130 -4.800 1418.690 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1435.610 -4.800 1436.170 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1453.550 -4.800 1454.110 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1471.490 -4.800 1472.050 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1489.430 -4.800 1489.990 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1506.910 -4.800 1507.470 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 704.210 -4.800 704.770 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1524.850 -4.800 1525.410 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1542.790 -4.800 1543.350 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1560.730 -4.800 1561.290 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1578.670 -4.800 1579.230 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1596.150 -4.800 1596.710 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1614.090 -4.800 1614.650 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1632.030 -4.800 1632.590 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1649.970 -4.800 1650.530 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1667.910 -4.800 1668.470 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1685.390 -4.800 1685.950 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 722.150 -4.800 722.710 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1703.330 -4.800 1703.890 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1721.270 -4.800 1721.830 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1739.210 -4.800 1739.770 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1756.690 -4.800 1757.250 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1774.630 -4.800 1775.190 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1792.570 -4.800 1793.130 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1810.510 -4.800 1811.070 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1828.450 -4.800 1829.010 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1845.930 -4.800 1846.490 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1863.870 -4.800 1864.430 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 740.090 -4.800 740.650 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1881.810 -4.800 1882.370 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1935.170 -4.800 1935.730 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1988.990 -4.800 1989.550 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2024.410 -4.800 2024.970 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2042.350 -4.800 2042.910 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 757.570 -4.800 758.130 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2060.290 -4.800 2060.850 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2078.230 -4.800 2078.790 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2095.710 -4.800 2096.270 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2113.650 -4.800 2114.210 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2131.590 -4.800 2132.150 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2149.530 -4.800 2150.090 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2167.470 -4.800 2168.030 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2184.950 -4.800 2185.510 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2202.890 -4.800 2203.450 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2220.830 -4.800 2221.390 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 775.510 -4.800 776.070 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2238.770 -4.800 2239.330 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2256.250 -4.800 2256.810 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2274.190 -4.800 2274.750 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2292.130 -4.800 2292.690 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2310.070 -4.800 2310.630 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2328.010 -4.800 2328.570 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2345.490 -4.800 2346.050 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2363.430 -4.800 2363.990 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2381.370 -4.800 2381.930 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2399.310 -4.800 2399.870 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 793.450 -4.800 794.010 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 639.010 25.740 639.330 25.800 ;
        RECT 686.850 25.740 687.170 25.800 ;
        RECT 639.010 25.600 687.170 25.740 ;
        RECT 639.010 25.540 639.330 25.600 ;
        RECT 686.850 25.540 687.170 25.600 ;
        RECT 687.310 25.060 687.630 25.120 ;
        RECT 1345.570 25.060 1345.890 25.120 ;
        RECT 687.310 24.920 1345.890 25.060 ;
        RECT 687.310 24.860 687.630 24.920 ;
        RECT 1345.570 24.860 1345.890 24.920 ;
      LAYER via ;
        RECT 639.040 25.540 639.300 25.800 ;
        RECT 686.880 25.540 687.140 25.800 ;
        RECT 687.340 24.860 687.600 25.120 ;
        RECT 1345.600 24.860 1345.860 25.120 ;
      LAYER met2 ;
        RECT 1346.130 1500.490 1346.410 1504.000 ;
        RECT 1345.660 1500.350 1346.410 1500.490 ;
        RECT 639.040 25.510 639.300 25.830 ;
        RECT 686.880 25.570 687.140 25.830 ;
        RECT 686.880 25.510 687.540 25.570 ;
        RECT 639.100 2.400 639.240 25.510 ;
        RECT 686.940 25.430 687.540 25.510 ;
        RECT 687.400 25.150 687.540 25.430 ;
        RECT 1345.660 25.150 1345.800 1500.350 ;
        RECT 1346.130 1500.000 1346.410 1500.350 ;
        RECT 687.340 24.830 687.600 25.150 ;
        RECT 1345.600 24.830 1345.860 25.150 ;
        RECT 638.890 -4.800 639.450 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2422.770 -4.800 2423.330 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2440.710 -4.800 2441.270 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2458.650 -4.800 2459.210 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2476.590 -4.800 2477.150 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2494.530 -4.800 2495.090 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2512.010 -4.800 2512.570 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2529.950 -4.800 2530.510 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2547.890 -4.800 2548.450 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2565.830 -4.800 2566.390 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2583.770 -4.800 2584.330 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 817.370 -4.800 817.930 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2601.250 -4.800 2601.810 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2619.190 -4.800 2619.750 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2637.130 -4.800 2637.690 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2655.070 -4.800 2655.630 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2672.550 -4.800 2673.110 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2690.490 -4.800 2691.050 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2708.430 -4.800 2708.990 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2726.370 -4.800 2726.930 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2744.310 -4.800 2744.870 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2761.790 -4.800 2762.350 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 835.310 -4.800 835.870 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2779.730 -4.800 2780.290 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2797.670 -4.800 2798.230 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2815.610 -4.800 2816.170 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2833.550 -4.800 2834.110 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2851.030 -4.800 2851.590 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2868.970 -4.800 2869.530 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 852.790 -4.800 853.350 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 870.730 -4.800 871.290 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 888.670 -4.800 889.230 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 906.610 -4.800 907.170 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 924.090 -4.800 924.650 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 942.030 -4.800 942.590 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 977.910 -4.800 978.470 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1375.110 1500.490 1375.390 1504.000 ;
        RECT 1373.260 1500.350 1375.390 1500.490 ;
        RECT 1373.260 24.325 1373.400 1500.350 ;
        RECT 1375.110 1500.000 1375.390 1500.350 ;
        RECT 656.970 23.955 657.250 24.325 ;
        RECT 1373.190 23.955 1373.470 24.325 ;
        RECT 657.040 2.400 657.180 23.955 ;
        RECT 656.830 -4.800 657.390 2.400 ;
      LAYER via2 ;
        RECT 656.970 24.000 657.250 24.280 ;
        RECT 1373.190 24.000 1373.470 24.280 ;
      LAYER met3 ;
        RECT 656.945 24.290 657.275 24.305 ;
        RECT 1373.165 24.290 1373.495 24.305 ;
        RECT 656.945 23.990 1373.495 24.290 ;
        RECT 656.945 23.975 657.275 23.990 ;
        RECT 1373.165 23.975 1373.495 23.990 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 995.850 -4.800 996.410 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1031.270 -4.800 1031.830 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1049.210 -4.800 1049.770 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1067.150 -4.800 1067.710 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1085.090 -4.800 1085.650 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1102.570 -4.800 1103.130 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1120.510 -4.800 1121.070 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1138.450 -4.800 1139.010 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1156.390 -4.800 1156.950 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 674.430 24.040 674.750 24.100 ;
        RECT 1393.870 24.040 1394.190 24.100 ;
        RECT 674.430 23.900 1394.190 24.040 ;
        RECT 674.430 23.840 674.750 23.900 ;
        RECT 1393.870 23.840 1394.190 23.900 ;
      LAYER via ;
        RECT 674.460 23.840 674.720 24.100 ;
        RECT 1393.900 23.840 1394.160 24.100 ;
      LAYER met2 ;
        RECT 1394.430 1500.490 1394.710 1504.000 ;
        RECT 1393.960 1500.350 1394.710 1500.490 ;
        RECT 1393.960 24.130 1394.100 1500.350 ;
        RECT 1394.430 1500.000 1394.710 1500.350 ;
        RECT 674.460 23.810 674.720 24.130 ;
        RECT 1393.900 23.810 1394.160 24.130 ;
        RECT 674.520 2.400 674.660 23.810 ;
        RECT 674.310 -4.800 674.870 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1173.870 -4.800 1174.430 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1191.810 -4.800 1192.370 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1209.750 -4.800 1210.310 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1227.690 -4.800 1228.250 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1245.630 -4.800 1246.190 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1263.110 -4.800 1263.670 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1281.050 -4.800 1281.610 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1298.990 -4.800 1299.550 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1316.930 -4.800 1317.490 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1334.870 -4.800 1335.430 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 692.250 -4.800 692.810 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1352.350 -4.800 1352.910 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1370.290 -4.800 1370.850 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1388.230 -4.800 1388.790 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1406.170 -4.800 1406.730 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1423.650 -4.800 1424.210 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1441.590 -4.800 1442.150 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1459.530 -4.800 1460.090 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1477.470 -4.800 1478.030 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1495.410 -4.800 1495.970 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1512.890 -4.800 1513.450 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 710.190 -4.800 710.750 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1530.830 -4.800 1531.390 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1548.770 -4.800 1549.330 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1566.710 -4.800 1567.270 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1584.650 -4.800 1585.210 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1602.130 -4.800 1602.690 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1620.070 -4.800 1620.630 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1638.010 -4.800 1638.570 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1655.950 -4.800 1656.510 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1673.430 -4.800 1673.990 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1691.370 -4.800 1691.930 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 728.130 -4.800 728.690 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1709.310 -4.800 1709.870 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1727.250 -4.800 1727.810 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1745.190 -4.800 1745.750 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1762.670 -4.800 1763.230 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1780.610 -4.800 1781.170 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1798.550 -4.800 1799.110 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1816.490 -4.800 1817.050 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1834.430 -4.800 1834.990 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1851.910 -4.800 1852.470 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1869.850 -4.800 1870.410 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 746.070 -4.800 746.630 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1887.790 -4.800 1888.350 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1923.210 -4.800 1923.770 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1977.030 -4.800 1977.590 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1994.970 -4.800 1995.530 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2030.390 -4.800 2030.950 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2048.330 -4.800 2048.890 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 763.550 -4.800 764.110 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2066.270 -4.800 2066.830 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2084.210 -4.800 2084.770 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2101.690 -4.800 2102.250 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2119.630 -4.800 2120.190 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2137.570 -4.800 2138.130 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2155.510 -4.800 2156.070 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2172.990 -4.800 2173.550 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2190.930 -4.800 2191.490 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2208.870 -4.800 2209.430 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2226.810 -4.800 2227.370 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 781.490 -4.800 782.050 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2244.750 -4.800 2245.310 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2262.230 -4.800 2262.790 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2280.170 -4.800 2280.730 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2298.110 -4.800 2298.670 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2316.050 -4.800 2316.610 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2333.990 -4.800 2334.550 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2351.470 -4.800 2352.030 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2369.410 -4.800 2369.970 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2387.350 -4.800 2387.910 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2405.290 -4.800 2405.850 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 799.430 -4.800 799.990 2.400 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 644.990 24.720 645.310 24.780 ;
        RECT 1352.470 24.720 1352.790 24.780 ;
        RECT 644.990 24.580 1352.790 24.720 ;
        RECT 644.990 24.520 645.310 24.580 ;
        RECT 1352.470 24.520 1352.790 24.580 ;
      LAYER via ;
        RECT 645.020 24.520 645.280 24.780 ;
        RECT 1352.500 24.520 1352.760 24.780 ;
      LAYER met2 ;
        RECT 1355.790 1500.490 1356.070 1504.000 ;
        RECT 1352.560 1500.350 1356.070 1500.490 ;
        RECT 1352.560 24.810 1352.700 1500.350 ;
        RECT 1355.790 1500.000 1356.070 1500.350 ;
        RECT 645.020 24.490 645.280 24.810 ;
        RECT 1352.500 24.490 1352.760 24.810 ;
        RECT 645.080 2.400 645.220 24.490 ;
        RECT 644.870 -4.800 645.430 2.400 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2428.750 -4.800 2429.310 2.400 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2446.690 -4.800 2447.250 2.400 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2464.630 -4.800 2465.190 2.400 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2482.570 -4.800 2483.130 2.400 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2500.510 -4.800 2501.070 2.400 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2517.990 -4.800 2518.550 2.400 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2535.930 -4.800 2536.490 2.400 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2553.870 -4.800 2554.430 2.400 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2571.810 -4.800 2572.370 2.400 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2589.290 -4.800 2589.850 2.400 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 823.350 -4.800 823.910 2.400 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2607.230 -4.800 2607.790 2.400 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2625.170 -4.800 2625.730 2.400 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2643.110 -4.800 2643.670 2.400 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2661.050 -4.800 2661.610 2.400 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2678.530 -4.800 2679.090 2.400 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2696.470 -4.800 2697.030 2.400 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2714.410 -4.800 2714.970 2.400 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2732.350 -4.800 2732.910 2.400 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2750.290 -4.800 2750.850 2.400 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2767.770 -4.800 2768.330 2.400 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 840.830 -4.800 841.390 2.400 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2785.710 -4.800 2786.270 2.400 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2803.650 -4.800 2804.210 2.400 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2821.590 -4.800 2822.150 2.400 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2839.070 -4.800 2839.630 2.400 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2857.010 -4.800 2857.570 2.400 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2874.950 -4.800 2875.510 2.400 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 858.770 -4.800 859.330 2.400 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 876.710 -4.800 877.270 2.400 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 894.650 -4.800 895.210 2.400 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 912.590 -4.800 913.150 2.400 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 930.070 -4.800 930.630 2.400 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 948.010 -4.800 948.570 2.400 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 983.890 -4.800 984.450 2.400 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 673.050 25.400 673.370 25.460 ;
        RECT 685.930 25.400 686.250 25.460 ;
        RECT 673.050 25.260 686.250 25.400 ;
        RECT 673.050 25.200 673.370 25.260 ;
        RECT 685.930 25.200 686.250 25.260 ;
        RECT 687.770 24.380 688.090 24.440 ;
        RECT 1380.070 24.380 1380.390 24.440 ;
        RECT 687.770 24.240 1380.390 24.380 ;
        RECT 687.770 24.180 688.090 24.240 ;
        RECT 1380.070 24.180 1380.390 24.240 ;
        RECT 662.930 24.040 663.250 24.100 ;
        RECT 673.050 24.040 673.370 24.100 ;
        RECT 662.930 23.900 673.370 24.040 ;
        RECT 662.930 23.840 663.250 23.900 ;
        RECT 673.050 23.840 673.370 23.900 ;
      LAYER via ;
        RECT 673.080 25.200 673.340 25.460 ;
        RECT 685.960 25.200 686.220 25.460 ;
        RECT 687.800 24.180 688.060 24.440 ;
        RECT 1380.100 24.180 1380.360 24.440 ;
        RECT 662.960 23.840 663.220 24.100 ;
        RECT 673.080 23.840 673.340 24.100 ;
      LAYER met2 ;
        RECT 1384.770 1500.490 1385.050 1504.000 ;
        RECT 1380.160 1500.350 1385.050 1500.490 ;
        RECT 686.020 26.110 688.000 26.250 ;
        RECT 686.020 25.490 686.160 26.110 ;
        RECT 673.080 25.170 673.340 25.490 ;
        RECT 685.960 25.170 686.220 25.490 ;
        RECT 673.140 24.130 673.280 25.170 ;
        RECT 687.860 24.470 688.000 26.110 ;
        RECT 1380.160 24.470 1380.300 1500.350 ;
        RECT 1384.770 1500.000 1385.050 1500.350 ;
        RECT 687.800 24.150 688.060 24.470 ;
        RECT 1380.100 24.150 1380.360 24.470 ;
        RECT 662.960 23.810 663.220 24.130 ;
        RECT 673.080 23.810 673.340 24.130 ;
        RECT 663.020 2.400 663.160 23.810 ;
        RECT 662.810 -4.800 663.370 2.400 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1001.830 -4.800 1002.390 2.400 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1037.250 -4.800 1037.810 2.400 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1055.190 -4.800 1055.750 2.400 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1073.130 -4.800 1073.690 2.400 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1090.610 -4.800 1091.170 2.400 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1108.550 -4.800 1109.110 2.400 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1126.490 -4.800 1127.050 2.400 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1144.430 -4.800 1144.990 2.400 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1162.370 -4.800 1162.930 2.400 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 680.290 -4.800 680.850 2.400 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1179.850 -4.800 1180.410 2.400 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1197.790 -4.800 1198.350 2.400 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1215.730 -4.800 1216.290 2.400 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1233.670 -4.800 1234.230 2.400 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1251.610 -4.800 1252.170 2.400 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1269.090 -4.800 1269.650 2.400 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1287.030 -4.800 1287.590 2.400 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1304.970 -4.800 1305.530 2.400 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1322.910 -4.800 1323.470 2.400 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1340.390 -4.800 1340.950 2.400 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 698.230 -4.800 698.790 2.400 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1358.330 -4.800 1358.890 2.400 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1376.270 -4.800 1376.830 2.400 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1394.210 -4.800 1394.770 2.400 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1412.150 -4.800 1412.710 2.400 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1429.630 -4.800 1430.190 2.400 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1447.570 -4.800 1448.130 2.400 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1465.510 -4.800 1466.070 2.400 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1483.450 -4.800 1484.010 2.400 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1501.390 -4.800 1501.950 2.400 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1518.870 -4.800 1519.430 2.400 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 716.170 -4.800 716.730 2.400 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1536.810 -4.800 1537.370 2.400 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1554.750 -4.800 1555.310 2.400 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1572.690 -4.800 1573.250 2.400 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1590.170 -4.800 1590.730 2.400 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1608.110 -4.800 1608.670 2.400 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1626.050 -4.800 1626.610 2.400 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1643.990 -4.800 1644.550 2.400 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1661.930 -4.800 1662.490 2.400 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1679.410 -4.800 1679.970 2.400 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1697.350 -4.800 1697.910 2.400 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 734.110 -4.800 734.670 2.400 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1715.290 -4.800 1715.850 2.400 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1733.230 -4.800 1733.790 2.400 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1751.170 -4.800 1751.730 2.400 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1768.650 -4.800 1769.210 2.400 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1786.590 -4.800 1787.150 2.400 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1804.530 -4.800 1805.090 2.400 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1822.470 -4.800 1823.030 2.400 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1839.950 -4.800 1840.510 2.400 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1857.890 -4.800 1858.450 2.400 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1875.830 -4.800 1876.390 2.400 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 752.050 -4.800 752.610 2.400 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1893.770 -4.800 1894.330 2.400 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1929.190 -4.800 1929.750 2.400 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1983.010 -4.800 1983.570 2.400 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2000.950 -4.800 2001.510 2.400 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2018.430 -4.800 2018.990 2.400 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2036.370 -4.800 2036.930 2.400 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2054.310 -4.800 2054.870 2.400 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 769.530 -4.800 770.090 2.400 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2072.250 -4.800 2072.810 2.400 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2089.730 -4.800 2090.290 2.400 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2107.670 -4.800 2108.230 2.400 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2125.610 -4.800 2126.170 2.400 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2143.550 -4.800 2144.110 2.400 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2161.490 -4.800 2162.050 2.400 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2178.970 -4.800 2179.530 2.400 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2196.910 -4.800 2197.470 2.400 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2214.850 -4.800 2215.410 2.400 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2232.790 -4.800 2233.350 2.400 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 787.470 -4.800 788.030 2.400 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2250.730 -4.800 2251.290 2.400 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2268.210 -4.800 2268.770 2.400 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2286.150 -4.800 2286.710 2.400 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2304.090 -4.800 2304.650 2.400 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2322.030 -4.800 2322.590 2.400 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2339.510 -4.800 2340.070 2.400 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2357.450 -4.800 2358.010 2.400 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2375.390 -4.800 2375.950 2.400 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2393.330 -4.800 2393.890 2.400 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2411.270 -4.800 2411.830 2.400 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 805.410 -4.800 805.970 2.400 ;
    END
  END la_oen[9]
  PIN user_clock2
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 321.610 2790.960 321.930 2791.020 ;
        RECT 968.830 2790.960 969.150 2791.020 ;
        RECT 1568.670 2790.960 1568.990 2791.020 ;
        RECT 2215.430 2790.960 2215.750 2791.020 ;
        RECT 321.610 2790.820 2215.750 2790.960 ;
        RECT 321.610 2790.760 321.930 2790.820 ;
        RECT 968.830 2790.760 969.150 2790.820 ;
        RECT 1568.670 2790.760 1568.990 2790.820 ;
        RECT 2215.430 2790.760 2215.750 2790.820 ;
        RECT 305.050 1462.720 305.370 1462.980 ;
        RECT 305.140 1462.580 305.280 1462.720 ;
        RECT 305.510 1462.580 305.830 1462.640 ;
        RECT 305.140 1462.440 305.830 1462.580 ;
        RECT 305.510 1462.380 305.830 1462.440 ;
        RECT 305.050 1442.180 305.370 1442.240 ;
        RECT 305.510 1442.180 305.830 1442.240 ;
        RECT 305.050 1442.040 305.830 1442.180 ;
        RECT 305.050 1441.980 305.370 1442.040 ;
        RECT 305.510 1441.980 305.830 1442.040 ;
        RECT 303.670 1366.360 303.990 1366.420 ;
        RECT 305.510 1366.360 305.830 1366.420 ;
        RECT 303.670 1366.220 305.830 1366.360 ;
        RECT 303.670 1366.160 303.990 1366.220 ;
        RECT 305.510 1366.160 305.830 1366.220 ;
        RECT 304.590 1317.740 304.910 1317.800 ;
        RECT 305.510 1317.740 305.830 1317.800 ;
        RECT 304.590 1317.600 305.830 1317.740 ;
        RECT 304.590 1317.540 304.910 1317.600 ;
        RECT 305.510 1317.540 305.830 1317.600 ;
        RECT 304.130 1304.140 304.450 1304.200 ;
        RECT 305.510 1304.140 305.830 1304.200 ;
        RECT 304.130 1304.000 305.830 1304.140 ;
        RECT 304.130 1303.940 304.450 1304.000 ;
        RECT 305.510 1303.940 305.830 1304.000 ;
        RECT 304.130 1256.200 304.450 1256.260 ;
        RECT 305.050 1256.200 305.370 1256.260 ;
        RECT 304.130 1256.060 305.370 1256.200 ;
        RECT 304.130 1256.000 304.450 1256.060 ;
        RECT 305.050 1256.000 305.370 1256.060 ;
        RECT 303.670 1124.760 303.990 1125.020 ;
        RECT 303.760 1124.280 303.900 1124.760 ;
        RECT 304.590 1124.280 304.910 1124.340 ;
        RECT 303.760 1124.140 304.910 1124.280 ;
        RECT 304.590 1124.080 304.910 1124.140 ;
        RECT 303.670 1076.680 303.990 1076.740 ;
        RECT 304.590 1076.680 304.910 1076.740 ;
        RECT 303.670 1076.540 304.910 1076.680 ;
        RECT 303.670 1076.480 303.990 1076.540 ;
        RECT 304.590 1076.480 304.910 1076.540 ;
        RECT 303.210 1027.720 303.530 1027.780 ;
        RECT 304.590 1027.720 304.910 1027.780 ;
        RECT 303.210 1027.580 304.910 1027.720 ;
        RECT 303.210 1027.520 303.530 1027.580 ;
        RECT 304.590 1027.520 304.910 1027.580 ;
        RECT 304.590 979.920 304.910 980.180 ;
        RECT 304.680 979.780 304.820 979.920 ;
        RECT 305.050 979.780 305.370 979.840 ;
        RECT 304.680 979.640 305.370 979.780 ;
        RECT 305.050 979.580 305.370 979.640 ;
        RECT 304.590 907.700 304.910 907.760 ;
        RECT 305.510 907.700 305.830 907.760 ;
        RECT 304.590 907.560 305.830 907.700 ;
        RECT 304.590 907.500 304.910 907.560 ;
        RECT 305.510 907.500 305.830 907.560 ;
        RECT 304.590 834.940 304.910 835.000 ;
        RECT 305.510 834.940 305.830 835.000 ;
        RECT 304.590 834.800 305.830 834.940 ;
        RECT 304.590 834.740 304.910 834.800 ;
        RECT 305.510 834.740 305.830 834.800 ;
        RECT 305.970 787.340 306.290 787.400 ;
        RECT 305.140 787.200 306.290 787.340 ;
        RECT 305.140 786.380 305.280 787.200 ;
        RECT 305.970 787.140 306.290 787.200 ;
        RECT 305.050 786.120 305.370 786.380 ;
        RECT 305.050 765.920 305.370 765.980 ;
        RECT 305.970 765.920 306.290 765.980 ;
        RECT 305.050 765.780 306.290 765.920 ;
        RECT 305.050 765.720 305.370 765.780 ;
        RECT 305.970 765.720 306.290 765.780 ;
        RECT 304.590 689.900 304.910 690.160 ;
        RECT 304.680 689.760 304.820 689.900 ;
        RECT 305.050 689.760 305.370 689.820 ;
        RECT 304.680 689.620 305.370 689.760 ;
        RECT 305.050 689.560 305.370 689.620 ;
        RECT 304.590 593.340 304.910 593.600 ;
        RECT 304.680 593.200 304.820 593.340 ;
        RECT 305.050 593.200 305.370 593.260 ;
        RECT 304.680 593.060 305.370 593.200 ;
        RECT 305.050 593.000 305.370 593.060 ;
        RECT 303.670 496.780 303.990 497.040 ;
        RECT 303.760 496.300 303.900 496.780 ;
        RECT 305.510 496.300 305.830 496.360 ;
        RECT 303.760 496.160 305.830 496.300 ;
        RECT 305.510 496.100 305.830 496.160 ;
        RECT 303.670 434.760 303.990 434.820 ;
        RECT 305.050 434.760 305.370 434.820 ;
        RECT 303.670 434.620 305.370 434.760 ;
        RECT 303.670 434.560 303.990 434.620 ;
        RECT 305.050 434.560 305.370 434.620 ;
        RECT 303.670 386.480 303.990 386.540 ;
        RECT 304.590 386.480 304.910 386.540 ;
        RECT 303.670 386.340 304.910 386.480 ;
        RECT 303.670 386.280 303.990 386.340 ;
        RECT 304.590 386.280 304.910 386.340 ;
        RECT 303.210 379.340 303.530 379.400 ;
        RECT 304.590 379.340 304.910 379.400 ;
        RECT 303.210 379.200 304.910 379.340 ;
        RECT 303.210 379.140 303.530 379.200 ;
        RECT 304.590 379.140 304.910 379.200 ;
        RECT 304.590 303.520 304.910 303.580 ;
        RECT 305.510 303.520 305.830 303.580 ;
        RECT 304.590 303.380 305.830 303.520 ;
        RECT 304.590 303.320 304.910 303.380 ;
        RECT 305.510 303.320 305.830 303.380 ;
        RECT 304.130 289.580 304.450 289.640 ;
        RECT 305.510 289.580 305.830 289.640 ;
        RECT 304.130 289.440 305.830 289.580 ;
        RECT 304.130 289.380 304.450 289.440 ;
        RECT 305.510 289.380 305.830 289.440 ;
        RECT 304.130 241.640 304.450 241.700 ;
        RECT 305.050 241.640 305.370 241.700 ;
        RECT 304.130 241.500 305.370 241.640 ;
        RECT 304.130 241.440 304.450 241.500 ;
        RECT 305.050 241.440 305.370 241.500 ;
        RECT 304.590 159.160 304.910 159.420 ;
        RECT 304.680 158.740 304.820 159.160 ;
        RECT 304.590 158.480 304.910 158.740 ;
        RECT 303.670 62.260 303.990 62.520 ;
        RECT 303.760 61.780 303.900 62.260 ;
        RECT 304.130 61.780 304.450 61.840 ;
        RECT 303.760 61.640 304.450 61.780 ;
        RECT 304.130 61.580 304.450 61.640 ;
        RECT 295.850 48.180 296.170 48.240 ;
        RECT 304.130 48.180 304.450 48.240 ;
        RECT 295.850 48.040 304.450 48.180 ;
        RECT 295.850 47.980 296.170 48.040 ;
        RECT 304.130 47.980 304.450 48.040 ;
        RECT 2.830 16.900 3.150 16.960 ;
        RECT 295.850 16.900 296.170 16.960 ;
        RECT 2.830 16.760 296.170 16.900 ;
        RECT 2.830 16.700 3.150 16.760 ;
        RECT 295.850 16.700 296.170 16.760 ;
      LAYER via ;
        RECT 321.640 2790.760 321.900 2791.020 ;
        RECT 968.860 2790.760 969.120 2791.020 ;
        RECT 1568.700 2790.760 1568.960 2791.020 ;
        RECT 2215.460 2790.760 2215.720 2791.020 ;
        RECT 305.080 1462.720 305.340 1462.980 ;
        RECT 305.540 1462.380 305.800 1462.640 ;
        RECT 305.080 1441.980 305.340 1442.240 ;
        RECT 305.540 1441.980 305.800 1442.240 ;
        RECT 303.700 1366.160 303.960 1366.420 ;
        RECT 305.540 1366.160 305.800 1366.420 ;
        RECT 304.620 1317.540 304.880 1317.800 ;
        RECT 305.540 1317.540 305.800 1317.800 ;
        RECT 304.160 1303.940 304.420 1304.200 ;
        RECT 305.540 1303.940 305.800 1304.200 ;
        RECT 304.160 1256.000 304.420 1256.260 ;
        RECT 305.080 1256.000 305.340 1256.260 ;
        RECT 303.700 1124.760 303.960 1125.020 ;
        RECT 304.620 1124.080 304.880 1124.340 ;
        RECT 303.700 1076.480 303.960 1076.740 ;
        RECT 304.620 1076.480 304.880 1076.740 ;
        RECT 303.240 1027.520 303.500 1027.780 ;
        RECT 304.620 1027.520 304.880 1027.780 ;
        RECT 304.620 979.920 304.880 980.180 ;
        RECT 305.080 979.580 305.340 979.840 ;
        RECT 304.620 907.500 304.880 907.760 ;
        RECT 305.540 907.500 305.800 907.760 ;
        RECT 304.620 834.740 304.880 835.000 ;
        RECT 305.540 834.740 305.800 835.000 ;
        RECT 306.000 787.140 306.260 787.400 ;
        RECT 305.080 786.120 305.340 786.380 ;
        RECT 305.080 765.720 305.340 765.980 ;
        RECT 306.000 765.720 306.260 765.980 ;
        RECT 304.620 689.900 304.880 690.160 ;
        RECT 305.080 689.560 305.340 689.820 ;
        RECT 304.620 593.340 304.880 593.600 ;
        RECT 305.080 593.000 305.340 593.260 ;
        RECT 303.700 496.780 303.960 497.040 ;
        RECT 305.540 496.100 305.800 496.360 ;
        RECT 303.700 434.560 303.960 434.820 ;
        RECT 305.080 434.560 305.340 434.820 ;
        RECT 303.700 386.280 303.960 386.540 ;
        RECT 304.620 386.280 304.880 386.540 ;
        RECT 303.240 379.140 303.500 379.400 ;
        RECT 304.620 379.140 304.880 379.400 ;
        RECT 304.620 303.320 304.880 303.580 ;
        RECT 305.540 303.320 305.800 303.580 ;
        RECT 304.160 289.380 304.420 289.640 ;
        RECT 305.540 289.380 305.800 289.640 ;
        RECT 304.160 241.440 304.420 241.700 ;
        RECT 305.080 241.440 305.340 241.700 ;
        RECT 304.620 159.160 304.880 159.420 ;
        RECT 304.620 158.480 304.880 158.740 ;
        RECT 303.700 62.260 303.960 62.520 ;
        RECT 304.160 61.580 304.420 61.840 ;
        RECT 295.880 47.980 296.140 48.240 ;
        RECT 304.160 47.980 304.420 48.240 ;
        RECT 2.860 16.700 3.120 16.960 ;
        RECT 295.880 16.700 296.140 16.960 ;
      LAYER met2 ;
        RECT 968.850 2794.275 969.130 2794.645 ;
        RECT 1568.690 2794.275 1568.970 2794.645 ;
        RECT 2215.450 2794.275 2215.730 2794.645 ;
        RECT 321.630 2793.595 321.910 2793.965 ;
        RECT 321.700 2791.050 321.840 2793.595 ;
        RECT 968.920 2791.050 969.060 2794.275 ;
        RECT 1568.760 2791.050 1568.900 2794.275 ;
        RECT 2215.520 2791.050 2215.660 2794.275 ;
        RECT 321.640 2790.730 321.900 2791.050 ;
        RECT 968.860 2790.730 969.120 2791.050 ;
        RECT 1568.700 2790.730 1568.960 2791.050 ;
        RECT 2215.460 2790.730 2215.720 2791.050 ;
        RECT 304.690 1503.890 304.970 1504.000 ;
        RECT 304.220 1503.750 304.970 1503.890 ;
        RECT 304.220 1503.325 304.360 1503.750 ;
        RECT 304.150 1502.955 304.430 1503.325 ;
        RECT 304.690 1500.000 304.970 1503.750 ;
        RECT 305.530 1497.515 305.810 1497.885 ;
        RECT 305.600 1490.290 305.740 1497.515 ;
        RECT 305.140 1490.150 305.740 1490.290 ;
        RECT 305.140 1463.010 305.280 1490.150 ;
        RECT 305.080 1462.690 305.340 1463.010 ;
        RECT 305.540 1462.350 305.800 1462.670 ;
        RECT 305.600 1442.270 305.740 1462.350 ;
        RECT 305.080 1441.950 305.340 1442.270 ;
        RECT 305.540 1441.950 305.800 1442.270 ;
        RECT 305.140 1425.010 305.280 1441.950 ;
        RECT 305.140 1424.870 305.740 1425.010 ;
        RECT 305.600 1366.450 305.740 1424.870 ;
        RECT 303.700 1366.130 303.960 1366.450 ;
        RECT 305.540 1366.130 305.800 1366.450 ;
        RECT 303.760 1365.850 303.900 1366.130 ;
        RECT 303.760 1365.710 304.360 1365.850 ;
        RECT 304.220 1318.250 304.360 1365.710 ;
        RECT 304.220 1318.110 304.820 1318.250 ;
        RECT 304.680 1317.830 304.820 1318.110 ;
        RECT 304.620 1317.510 304.880 1317.830 ;
        RECT 305.540 1317.510 305.800 1317.830 ;
        RECT 305.600 1304.230 305.740 1317.510 ;
        RECT 304.160 1303.910 304.420 1304.230 ;
        RECT 305.540 1303.910 305.800 1304.230 ;
        RECT 304.220 1256.290 304.360 1303.910 ;
        RECT 304.160 1255.970 304.420 1256.290 ;
        RECT 305.080 1255.970 305.340 1256.290 ;
        RECT 305.140 1221.010 305.280 1255.970 ;
        RECT 304.220 1220.870 305.280 1221.010 ;
        RECT 304.220 1173.410 304.360 1220.870 ;
        RECT 303.760 1173.270 304.360 1173.410 ;
        RECT 303.760 1125.050 303.900 1173.270 ;
        RECT 303.700 1124.730 303.960 1125.050 ;
        RECT 304.620 1124.050 304.880 1124.370 ;
        RECT 304.680 1076.770 304.820 1124.050 ;
        RECT 303.700 1076.450 303.960 1076.770 ;
        RECT 304.620 1076.450 304.880 1076.770 ;
        RECT 303.760 1038.770 303.900 1076.450 ;
        RECT 303.300 1038.630 303.900 1038.770 ;
        RECT 303.300 1027.810 303.440 1038.630 ;
        RECT 303.240 1027.490 303.500 1027.810 ;
        RECT 304.620 1027.490 304.880 1027.810 ;
        RECT 304.680 980.210 304.820 1027.490 ;
        RECT 304.620 979.890 304.880 980.210 ;
        RECT 305.080 979.550 305.340 979.870 ;
        RECT 305.140 931.330 305.280 979.550 ;
        RECT 304.680 931.190 305.280 931.330 ;
        RECT 304.680 907.790 304.820 931.190 ;
        RECT 304.620 907.470 304.880 907.790 ;
        RECT 305.540 907.470 305.800 907.790 ;
        RECT 305.600 869.565 305.740 907.470 ;
        RECT 304.610 869.195 304.890 869.565 ;
        RECT 305.530 869.195 305.810 869.565 ;
        RECT 304.680 835.030 304.820 869.195 ;
        RECT 304.620 834.710 304.880 835.030 ;
        RECT 305.540 834.710 305.800 835.030 ;
        RECT 305.600 821.170 305.740 834.710 ;
        RECT 305.600 821.030 306.200 821.170 ;
        RECT 306.060 787.430 306.200 821.030 ;
        RECT 306.000 787.110 306.260 787.430 ;
        RECT 305.080 786.090 305.340 786.410 ;
        RECT 305.140 766.010 305.280 786.090 ;
        RECT 305.080 765.690 305.340 766.010 ;
        RECT 306.000 765.690 306.260 766.010 ;
        RECT 306.060 717.925 306.200 765.690 ;
        RECT 304.610 717.555 304.890 717.925 ;
        RECT 305.990 717.555 306.270 717.925 ;
        RECT 304.680 690.190 304.820 717.555 ;
        RECT 304.620 689.870 304.880 690.190 ;
        RECT 305.080 689.530 305.340 689.850 ;
        RECT 305.140 676.160 305.280 689.530 ;
        RECT 304.220 676.020 305.280 676.160 ;
        RECT 304.220 628.050 304.360 676.020 ;
        RECT 304.220 627.910 304.820 628.050 ;
        RECT 304.680 593.630 304.820 627.910 ;
        RECT 304.620 593.310 304.880 593.630 ;
        RECT 305.080 592.970 305.340 593.290 ;
        RECT 305.140 531.605 305.280 592.970 ;
        RECT 303.690 531.235 303.970 531.605 ;
        RECT 305.070 531.235 305.350 531.605 ;
        RECT 303.760 497.070 303.900 531.235 ;
        RECT 303.700 496.750 303.960 497.070 ;
        RECT 305.540 496.070 305.800 496.390 ;
        RECT 305.600 448.530 305.740 496.070 ;
        RECT 305.140 448.390 305.740 448.530 ;
        RECT 305.140 434.850 305.280 448.390 ;
        RECT 303.700 434.530 303.960 434.850 ;
        RECT 305.080 434.530 305.340 434.850 ;
        RECT 303.760 386.570 303.900 434.530 ;
        RECT 303.700 386.250 303.960 386.570 ;
        RECT 304.620 386.250 304.880 386.570 ;
        RECT 304.680 379.430 304.820 386.250 ;
        RECT 303.240 379.110 303.500 379.430 ;
        RECT 304.620 379.110 304.880 379.430 ;
        RECT 303.300 351.290 303.440 379.110 ;
        RECT 303.300 351.150 304.360 351.290 ;
        RECT 304.220 303.690 304.360 351.150 ;
        RECT 304.220 303.610 304.820 303.690 ;
        RECT 304.220 303.550 304.880 303.610 ;
        RECT 304.620 303.290 304.880 303.550 ;
        RECT 305.540 303.290 305.800 303.610 ;
        RECT 305.600 289.670 305.740 303.290 ;
        RECT 304.160 289.350 304.420 289.670 ;
        RECT 305.540 289.350 305.800 289.670 ;
        RECT 304.220 241.730 304.360 289.350 ;
        RECT 304.160 241.410 304.420 241.730 ;
        RECT 305.080 241.410 305.340 241.730 ;
        RECT 305.140 207.130 305.280 241.410 ;
        RECT 304.680 206.990 305.280 207.130 ;
        RECT 304.680 159.450 304.820 206.990 ;
        RECT 304.620 159.130 304.880 159.450 ;
        RECT 304.620 158.450 304.880 158.770 ;
        RECT 304.680 110.570 304.820 158.450 ;
        RECT 303.760 110.430 304.820 110.570 ;
        RECT 303.760 62.550 303.900 110.430 ;
        RECT 303.700 62.230 303.960 62.550 ;
        RECT 304.160 61.550 304.420 61.870 ;
        RECT 304.220 48.270 304.360 61.550 ;
        RECT 295.880 47.950 296.140 48.270 ;
        RECT 304.160 47.950 304.420 48.270 ;
        RECT 295.940 16.990 296.080 47.950 ;
        RECT 2.860 16.670 3.120 16.990 ;
        RECT 295.880 16.670 296.140 16.990 ;
        RECT 2.920 2.400 3.060 16.670 ;
        RECT 2.710 -4.800 3.270 2.400 ;
      LAYER via2 ;
        RECT 968.850 2794.320 969.130 2794.600 ;
        RECT 1568.690 2794.320 1568.970 2794.600 ;
        RECT 2215.450 2794.320 2215.730 2794.600 ;
        RECT 321.630 2793.640 321.910 2793.920 ;
        RECT 304.150 1503.000 304.430 1503.280 ;
        RECT 305.530 1497.560 305.810 1497.840 ;
        RECT 304.610 869.240 304.890 869.520 ;
        RECT 305.530 869.240 305.810 869.520 ;
        RECT 304.610 717.600 304.890 717.880 ;
        RECT 305.990 717.600 306.270 717.880 ;
        RECT 303.690 531.280 303.970 531.560 ;
        RECT 305.070 531.280 305.350 531.560 ;
      LAYER met3 ;
        RECT 968.825 2794.620 969.155 2794.625 ;
        RECT 1568.665 2794.620 1568.995 2794.625 ;
        RECT 2215.425 2794.620 2215.755 2794.625 ;
        RECT 968.825 2794.610 969.410 2794.620 ;
        RECT 1568.665 2794.610 1569.250 2794.620 ;
        RECT 2215.425 2794.610 2216.010 2794.620 ;
        RECT 968.825 2794.310 969.610 2794.610 ;
        RECT 1568.665 2794.310 1569.450 2794.610 ;
        RECT 2215.425 2794.310 2216.210 2794.610 ;
        RECT 968.825 2794.300 969.410 2794.310 ;
        RECT 1568.665 2794.300 1569.250 2794.310 ;
        RECT 2215.425 2794.300 2216.010 2794.310 ;
        RECT 968.825 2794.295 969.155 2794.300 ;
        RECT 1568.665 2794.295 1568.995 2794.300 ;
        RECT 2215.425 2794.295 2215.755 2794.300 ;
        RECT 308.470 2793.930 308.850 2793.940 ;
        RECT 317.670 2793.930 318.050 2793.940 ;
        RECT 321.605 2793.930 321.935 2793.945 ;
        RECT 308.470 2793.630 321.935 2793.930 ;
        RECT 308.470 2793.620 308.850 2793.630 ;
        RECT 317.670 2793.620 318.050 2793.630 ;
        RECT 321.605 2793.615 321.935 2793.630 ;
        RECT 304.125 1503.290 304.455 1503.305 ;
        RECT 305.710 1503.290 306.090 1503.300 ;
        RECT 308.470 1503.290 308.850 1503.300 ;
        RECT 304.125 1502.990 308.850 1503.290 ;
        RECT 304.125 1502.975 304.455 1502.990 ;
        RECT 305.710 1502.980 306.090 1502.990 ;
        RECT 308.470 1502.980 308.850 1502.990 ;
        RECT 305.505 1497.860 305.835 1497.865 ;
        RECT 305.505 1497.850 306.090 1497.860 ;
        RECT 305.505 1497.550 306.290 1497.850 ;
        RECT 305.505 1497.540 306.090 1497.550 ;
        RECT 305.505 1497.535 305.835 1497.540 ;
        RECT 304.585 869.530 304.915 869.545 ;
        RECT 305.505 869.530 305.835 869.545 ;
        RECT 304.585 869.230 305.835 869.530 ;
        RECT 304.585 869.215 304.915 869.230 ;
        RECT 305.505 869.215 305.835 869.230 ;
        RECT 304.585 717.890 304.915 717.905 ;
        RECT 305.965 717.890 306.295 717.905 ;
        RECT 304.585 717.590 306.295 717.890 ;
        RECT 304.585 717.575 304.915 717.590 ;
        RECT 305.965 717.575 306.295 717.590 ;
        RECT 303.665 531.570 303.995 531.585 ;
        RECT 305.045 531.570 305.375 531.585 ;
        RECT 303.665 531.270 305.375 531.570 ;
        RECT 303.665 531.255 303.995 531.270 ;
        RECT 305.045 531.255 305.375 531.270 ;
      LAYER via3 ;
        RECT 969.060 2794.300 969.380 2794.620 ;
        RECT 1568.900 2794.300 1569.220 2794.620 ;
        RECT 2215.660 2794.300 2215.980 2794.620 ;
        RECT 308.500 2793.620 308.820 2793.940 ;
        RECT 317.700 2793.620 318.020 2793.940 ;
        RECT 305.740 1502.980 306.060 1503.300 ;
        RECT 308.500 1502.980 308.820 1503.300 ;
        RECT 305.740 1497.540 306.060 1497.860 ;
      LAYER met4 ;
        RECT 319.015 2801.750 319.315 2804.600 ;
        RECT 317.710 2801.450 319.315 2801.750 ;
        RECT 317.710 2793.945 318.010 2801.450 ;
        RECT 319.015 2800.000 319.315 2801.450 ;
        RECT 969.015 2801.750 969.315 2804.600 ;
        RECT 1569.015 2801.750 1569.315 2804.600 ;
        RECT 2219.015 2801.750 2219.315 2804.600 ;
        RECT 969.015 2800.000 969.370 2801.750 ;
        RECT 969.070 2794.625 969.370 2800.000 ;
        RECT 1568.910 2800.000 1569.315 2801.750 ;
        RECT 2215.670 2801.450 2219.315 2801.750 ;
        RECT 1568.910 2794.625 1569.210 2800.000 ;
        RECT 2215.670 2794.625 2215.970 2801.450 ;
        RECT 2219.015 2800.000 2219.315 2801.450 ;
        RECT 969.055 2794.295 969.385 2794.625 ;
        RECT 1568.895 2794.295 1569.225 2794.625 ;
        RECT 2215.655 2794.295 2215.985 2794.625 ;
        RECT 308.495 2793.615 308.825 2793.945 ;
        RECT 317.695 2793.615 318.025 2793.945 ;
        RECT 308.510 1503.305 308.810 2793.615 ;
        RECT 305.735 1502.975 306.065 1503.305 ;
        RECT 308.495 1502.975 308.825 1503.305 ;
        RECT 305.750 1497.865 306.050 1502.975 ;
        RECT 305.735 1497.535 306.065 1497.865 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 8.350 16.560 8.670 16.620 ;
        RECT 311.030 16.560 311.350 16.620 ;
        RECT 8.350 16.420 311.350 16.560 ;
        RECT 8.350 16.360 8.670 16.420 ;
        RECT 311.030 16.360 311.350 16.420 ;
      LAYER via ;
        RECT 8.380 16.360 8.640 16.620 ;
        RECT 311.060 16.360 311.320 16.620 ;
      LAYER met2 ;
        RECT 314.350 1500.490 314.630 1504.000 ;
        RECT 311.120 1500.350 314.630 1500.490 ;
        RECT 311.120 16.650 311.260 1500.350 ;
        RECT 314.350 1500.000 314.630 1500.350 ;
        RECT 8.380 16.330 8.640 16.650 ;
        RECT 311.060 16.330 311.320 16.650 ;
        RECT 8.440 2.400 8.580 16.330 ;
        RECT 8.230 -4.800 8.790 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 20.310 1489.780 20.630 1489.840 ;
        RECT 323.910 1489.780 324.230 1489.840 ;
        RECT 20.310 1489.640 324.230 1489.780 ;
        RECT 20.310 1489.580 20.630 1489.640 ;
        RECT 323.910 1489.580 324.230 1489.640 ;
        RECT 14.330 17.580 14.650 17.640 ;
        RECT 20.310 17.580 20.630 17.640 ;
        RECT 14.330 17.440 20.630 17.580 ;
        RECT 14.330 17.380 14.650 17.440 ;
        RECT 20.310 17.380 20.630 17.440 ;
      LAYER via ;
        RECT 20.340 1489.580 20.600 1489.840 ;
        RECT 323.940 1489.580 324.200 1489.840 ;
        RECT 14.360 17.380 14.620 17.640 ;
        RECT 20.340 17.380 20.600 17.640 ;
      LAYER met2 ;
        RECT 324.010 1500.420 324.290 1504.000 ;
        RECT 324.000 1500.000 324.290 1500.420 ;
        RECT 324.000 1489.870 324.140 1500.000 ;
        RECT 20.340 1489.550 20.600 1489.870 ;
        RECT 323.940 1489.550 324.200 1489.870 ;
        RECT 20.400 17.670 20.540 1489.550 ;
        RECT 14.360 17.350 14.620 17.670 ;
        RECT 20.340 17.350 20.600 17.670 ;
        RECT 14.420 2.400 14.560 17.350 ;
        RECT 14.210 -4.800 14.770 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 38.250 27.440 38.570 27.500 ;
        RECT 358.870 27.440 359.190 27.500 ;
        RECT 38.250 27.300 359.190 27.440 ;
        RECT 38.250 27.240 38.570 27.300 ;
        RECT 358.870 27.240 359.190 27.300 ;
      LAYER via ;
        RECT 38.280 27.240 38.540 27.500 ;
        RECT 358.900 27.240 359.160 27.500 ;
      LAYER met2 ;
        RECT 362.650 1500.490 362.930 1504.000 ;
        RECT 358.960 1500.350 362.930 1500.490 ;
        RECT 358.960 27.530 359.100 1500.350 ;
        RECT 362.650 1500.000 362.930 1500.350 ;
        RECT 38.280 27.210 38.540 27.530 ;
        RECT 358.900 27.210 359.160 27.530 ;
        RECT 38.340 2.400 38.480 27.210 ;
        RECT 38.130 -4.800 38.690 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 241.110 20.980 241.430 21.040 ;
        RECT 690.070 20.980 690.390 21.040 ;
        RECT 241.110 20.840 690.390 20.980 ;
        RECT 241.110 20.780 241.430 20.840 ;
        RECT 690.070 20.780 690.390 20.840 ;
      LAYER via ;
        RECT 241.140 20.780 241.400 21.040 ;
        RECT 690.100 20.780 690.360 21.040 ;
      LAYER met2 ;
        RECT 693.850 1500.490 694.130 1504.000 ;
        RECT 690.160 1500.350 694.130 1500.490 ;
        RECT 690.160 21.070 690.300 1500.350 ;
        RECT 693.850 1500.000 694.130 1500.350 ;
        RECT 241.140 20.750 241.400 21.070 ;
        RECT 690.100 20.750 690.360 21.070 ;
        RECT 241.200 10.610 241.340 20.750 ;
        RECT 240.740 10.470 241.340 10.610 ;
        RECT 240.740 2.400 240.880 10.470 ;
        RECT 240.530 -4.800 241.090 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 258.130 21.320 258.450 21.380 ;
        RECT 717.670 21.320 717.990 21.380 ;
        RECT 258.130 21.180 717.990 21.320 ;
        RECT 258.130 21.120 258.450 21.180 ;
        RECT 717.670 21.120 717.990 21.180 ;
      LAYER via ;
        RECT 258.160 21.120 258.420 21.380 ;
        RECT 717.700 21.120 717.960 21.380 ;
      LAYER met2 ;
        RECT 722.830 1500.490 723.110 1504.000 ;
        RECT 717.760 1500.350 723.110 1500.490 ;
        RECT 717.760 21.410 717.900 1500.350 ;
        RECT 722.830 1500.000 723.110 1500.350 ;
        RECT 258.160 21.090 258.420 21.410 ;
        RECT 717.700 21.090 717.960 21.410 ;
        RECT 258.220 2.400 258.360 21.090 ;
        RECT 258.010 -4.800 258.570 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 276.070 21.660 276.390 21.720 ;
        RECT 752.170 21.660 752.490 21.720 ;
        RECT 276.070 21.520 752.490 21.660 ;
        RECT 276.070 21.460 276.390 21.520 ;
        RECT 752.170 21.460 752.490 21.520 ;
      LAYER via ;
        RECT 276.100 21.460 276.360 21.720 ;
        RECT 752.200 21.460 752.460 21.720 ;
      LAYER met2 ;
        RECT 752.270 1500.420 752.550 1504.000 ;
        RECT 752.260 1500.000 752.550 1500.420 ;
        RECT 752.260 21.750 752.400 1500.000 ;
        RECT 276.100 21.430 276.360 21.750 ;
        RECT 752.200 21.430 752.460 21.750 ;
        RECT 276.160 2.400 276.300 21.430 ;
        RECT 275.950 -4.800 276.510 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 294.010 22.000 294.330 22.060 ;
        RECT 779.770 22.000 780.090 22.060 ;
        RECT 294.010 21.860 780.090 22.000 ;
        RECT 294.010 21.800 294.330 21.860 ;
        RECT 779.770 21.800 780.090 21.860 ;
      LAYER via ;
        RECT 294.040 21.800 294.300 22.060 ;
        RECT 779.800 21.800 780.060 22.060 ;
      LAYER met2 ;
        RECT 781.250 1500.490 781.530 1504.000 ;
        RECT 779.860 1500.350 781.530 1500.490 ;
        RECT 779.860 22.090 780.000 1500.350 ;
        RECT 781.250 1500.000 781.530 1500.350 ;
        RECT 294.040 21.770 294.300 22.090 ;
        RECT 779.800 21.770 780.060 22.090 ;
        RECT 294.100 2.400 294.240 21.770 ;
        RECT 293.890 -4.800 294.450 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 311.950 22.340 312.270 22.400 ;
        RECT 807.370 22.340 807.690 22.400 ;
        RECT 311.950 22.200 807.690 22.340 ;
        RECT 311.950 22.140 312.270 22.200 ;
        RECT 807.370 22.140 807.690 22.200 ;
      LAYER via ;
        RECT 311.980 22.140 312.240 22.400 ;
        RECT 807.400 22.140 807.660 22.400 ;
      LAYER met2 ;
        RECT 810.690 1500.490 810.970 1504.000 ;
        RECT 807.460 1500.350 810.970 1500.490 ;
        RECT 807.460 22.430 807.600 1500.350 ;
        RECT 810.690 1500.000 810.970 1500.350 ;
        RECT 311.980 22.110 312.240 22.430 ;
        RECT 807.400 22.110 807.660 22.430 ;
        RECT 312.040 2.400 312.180 22.110 ;
        RECT 311.830 -4.800 312.390 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 329.890 22.680 330.210 22.740 ;
        RECT 834.970 22.680 835.290 22.740 ;
        RECT 329.890 22.540 835.290 22.680 ;
        RECT 329.890 22.480 330.210 22.540 ;
        RECT 834.970 22.480 835.290 22.540 ;
      LAYER via ;
        RECT 329.920 22.480 330.180 22.740 ;
        RECT 835.000 22.480 835.260 22.740 ;
      LAYER met2 ;
        RECT 839.670 1500.490 839.950 1504.000 ;
        RECT 835.060 1500.350 839.950 1500.490 ;
        RECT 835.060 22.770 835.200 1500.350 ;
        RECT 839.670 1500.000 839.950 1500.350 ;
        RECT 329.920 22.450 330.180 22.770 ;
        RECT 835.000 22.450 835.260 22.770 ;
        RECT 329.980 2.400 330.120 22.450 ;
        RECT 329.770 -4.800 330.330 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 347.370 23.020 347.690 23.080 ;
        RECT 862.570 23.020 862.890 23.080 ;
        RECT 347.370 22.880 862.890 23.020 ;
        RECT 347.370 22.820 347.690 22.880 ;
        RECT 862.570 22.820 862.890 22.880 ;
      LAYER via ;
        RECT 347.400 22.820 347.660 23.080 ;
        RECT 862.600 22.820 862.860 23.080 ;
      LAYER met2 ;
        RECT 869.110 1500.490 869.390 1504.000 ;
        RECT 862.660 1500.350 869.390 1500.490 ;
        RECT 862.660 23.110 862.800 1500.350 ;
        RECT 869.110 1500.000 869.390 1500.350 ;
        RECT 347.400 22.790 347.660 23.110 ;
        RECT 862.600 22.790 862.860 23.110 ;
        RECT 347.460 2.400 347.600 22.790 ;
        RECT 347.250 -4.800 347.810 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 365.310 23.360 365.630 23.420 ;
        RECT 897.070 23.360 897.390 23.420 ;
        RECT 365.310 23.220 897.390 23.360 ;
        RECT 365.310 23.160 365.630 23.220 ;
        RECT 897.070 23.160 897.390 23.220 ;
      LAYER via ;
        RECT 365.340 23.160 365.600 23.420 ;
        RECT 897.100 23.160 897.360 23.420 ;
      LAYER met2 ;
        RECT 898.090 1500.490 898.370 1504.000 ;
        RECT 897.160 1500.350 898.370 1500.490 ;
        RECT 897.160 23.450 897.300 1500.350 ;
        RECT 898.090 1500.000 898.370 1500.350 ;
        RECT 365.340 23.130 365.600 23.450 ;
        RECT 897.100 23.130 897.360 23.450 ;
        RECT 365.400 2.400 365.540 23.130 ;
        RECT 365.190 -4.800 365.750 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 383.250 23.700 383.570 23.760 ;
        RECT 924.670 23.700 924.990 23.760 ;
        RECT 383.250 23.560 924.990 23.700 ;
        RECT 383.250 23.500 383.570 23.560 ;
        RECT 924.670 23.500 924.990 23.560 ;
      LAYER via ;
        RECT 383.280 23.500 383.540 23.760 ;
        RECT 924.700 23.500 924.960 23.760 ;
      LAYER met2 ;
        RECT 927.530 1500.490 927.810 1504.000 ;
        RECT 924.760 1500.350 927.810 1500.490 ;
        RECT 924.760 23.790 924.900 1500.350 ;
        RECT 927.530 1500.000 927.810 1500.350 ;
        RECT 383.280 23.470 383.540 23.790 ;
        RECT 924.700 23.470 924.960 23.790 ;
        RECT 383.340 2.400 383.480 23.470 ;
        RECT 383.130 -4.800 383.690 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 401.190 27.440 401.510 27.500 ;
        RECT 952.270 27.440 952.590 27.500 ;
        RECT 401.190 27.300 952.590 27.440 ;
        RECT 401.190 27.240 401.510 27.300 ;
        RECT 952.270 27.240 952.590 27.300 ;
      LAYER via ;
        RECT 401.220 27.240 401.480 27.500 ;
        RECT 952.300 27.240 952.560 27.500 ;
      LAYER met2 ;
        RECT 956.510 1500.490 956.790 1504.000 ;
        RECT 952.360 1500.350 956.790 1500.490 ;
        RECT 952.360 27.530 952.500 1500.350 ;
        RECT 956.510 1500.000 956.790 1500.350 ;
        RECT 401.220 27.210 401.480 27.530 ;
        RECT 952.300 27.210 952.560 27.530 ;
        RECT 401.280 2.400 401.420 27.210 ;
        RECT 401.070 -4.800 401.630 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 62.170 27.100 62.490 27.160 ;
        RECT 400.270 27.100 400.590 27.160 ;
        RECT 62.170 26.960 400.590 27.100 ;
        RECT 62.170 26.900 62.490 26.960 ;
        RECT 400.270 26.900 400.590 26.960 ;
      LAYER via ;
        RECT 62.200 26.900 62.460 27.160 ;
        RECT 400.300 26.900 400.560 27.160 ;
      LAYER met2 ;
        RECT 401.750 1500.490 402.030 1504.000 ;
        RECT 400.360 1500.350 402.030 1500.490 ;
        RECT 400.360 27.190 400.500 1500.350 ;
        RECT 401.750 1500.000 402.030 1500.350 ;
        RECT 62.200 26.870 62.460 27.190 ;
        RECT 400.300 26.870 400.560 27.190 ;
        RECT 62.260 2.400 62.400 26.870 ;
        RECT 62.050 -4.800 62.610 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 419.130 27.100 419.450 27.160 ;
        RECT 979.870 27.100 980.190 27.160 ;
        RECT 419.130 26.960 980.190 27.100 ;
        RECT 419.130 26.900 419.450 26.960 ;
        RECT 979.870 26.900 980.190 26.960 ;
      LAYER via ;
        RECT 419.160 26.900 419.420 27.160 ;
        RECT 979.900 26.900 980.160 27.160 ;
      LAYER met2 ;
        RECT 985.950 1500.490 986.230 1504.000 ;
        RECT 979.960 1500.350 986.230 1500.490 ;
        RECT 979.960 27.190 980.100 1500.350 ;
        RECT 985.950 1500.000 986.230 1500.350 ;
        RECT 419.160 26.870 419.420 27.190 ;
        RECT 979.900 26.870 980.160 27.190 ;
        RECT 419.220 2.400 419.360 26.870 ;
        RECT 419.010 -4.800 419.570 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 436.610 26.760 436.930 26.820 ;
        RECT 1014.370 26.760 1014.690 26.820 ;
        RECT 436.610 26.620 1014.690 26.760 ;
        RECT 436.610 26.560 436.930 26.620 ;
        RECT 1014.370 26.560 1014.690 26.620 ;
      LAYER via ;
        RECT 436.640 26.560 436.900 26.820 ;
        RECT 1014.400 26.560 1014.660 26.820 ;
      LAYER met2 ;
        RECT 1014.930 1500.490 1015.210 1504.000 ;
        RECT 1014.460 1500.350 1015.210 1500.490 ;
        RECT 1014.460 26.850 1014.600 1500.350 ;
        RECT 1014.930 1500.000 1015.210 1500.350 ;
        RECT 436.640 26.530 436.900 26.850 ;
        RECT 1014.400 26.530 1014.660 26.850 ;
        RECT 436.700 2.400 436.840 26.530 ;
        RECT 436.490 -4.800 437.050 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1044.370 1500.490 1044.650 1504.000 ;
        RECT 1042.060 1500.350 1044.650 1500.490 ;
        RECT 1042.060 26.365 1042.200 1500.350 ;
        RECT 1044.370 1500.000 1044.650 1500.350 ;
        RECT 454.570 25.995 454.850 26.365 ;
        RECT 1041.990 25.995 1042.270 26.365 ;
        RECT 454.640 2.400 454.780 25.995 ;
        RECT 454.430 -4.800 454.990 2.400 ;
      LAYER via2 ;
        RECT 454.570 26.040 454.850 26.320 ;
        RECT 1041.990 26.040 1042.270 26.320 ;
      LAYER met3 ;
        RECT 454.545 26.330 454.875 26.345 ;
        RECT 1041.965 26.330 1042.295 26.345 ;
        RECT 454.545 26.030 1042.295 26.330 ;
        RECT 454.545 26.015 454.875 26.030 ;
        RECT 1041.965 26.015 1042.295 26.030 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1073.350 1500.490 1073.630 1504.000 ;
        RECT 1069.660 1500.350 1073.630 1500.490 ;
        RECT 1069.660 25.685 1069.800 1500.350 ;
        RECT 1073.350 1500.000 1073.630 1500.350 ;
        RECT 472.510 25.315 472.790 25.685 ;
        RECT 1069.590 25.315 1069.870 25.685 ;
        RECT 472.580 2.400 472.720 25.315 ;
        RECT 472.370 -4.800 472.930 2.400 ;
      LAYER via2 ;
        RECT 472.510 25.360 472.790 25.640 ;
        RECT 1069.590 25.360 1069.870 25.640 ;
      LAYER met3 ;
        RECT 472.485 25.650 472.815 25.665 ;
        RECT 1069.565 25.650 1069.895 25.665 ;
        RECT 472.485 25.350 1069.895 25.650 ;
        RECT 472.485 25.335 472.815 25.350 ;
        RECT 1069.565 25.335 1069.895 25.350 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 544.710 27.780 545.030 27.840 ;
        RECT 545.170 27.780 545.490 27.840 ;
        RECT 544.710 27.640 545.490 27.780 ;
        RECT 544.710 27.580 545.030 27.640 ;
        RECT 545.170 27.580 545.490 27.640 ;
        RECT 544.710 26.420 545.030 26.480 ;
        RECT 496.960 26.280 545.030 26.420 ;
        RECT 490.430 26.080 490.750 26.140 ;
        RECT 496.960 26.080 497.100 26.280 ;
        RECT 544.710 26.220 545.030 26.280 ;
        RECT 545.170 26.420 545.490 26.480 ;
        RECT 1097.170 26.420 1097.490 26.480 ;
        RECT 545.170 26.280 1097.490 26.420 ;
        RECT 545.170 26.220 545.490 26.280 ;
        RECT 1097.170 26.220 1097.490 26.280 ;
        RECT 490.430 25.940 497.100 26.080 ;
        RECT 490.430 25.880 490.750 25.940 ;
      LAYER via ;
        RECT 544.740 27.580 545.000 27.840 ;
        RECT 545.200 27.580 545.460 27.840 ;
        RECT 490.460 25.880 490.720 26.140 ;
        RECT 544.740 26.220 545.000 26.480 ;
        RECT 545.200 26.220 545.460 26.480 ;
        RECT 1097.200 26.220 1097.460 26.480 ;
      LAYER met2 ;
        RECT 1102.790 1500.490 1103.070 1504.000 ;
        RECT 1097.260 1500.350 1103.070 1500.490 ;
        RECT 544.740 27.550 545.000 27.870 ;
        RECT 545.200 27.550 545.460 27.870 ;
        RECT 544.800 26.510 544.940 27.550 ;
        RECT 545.260 26.510 545.400 27.550 ;
        RECT 1097.260 26.510 1097.400 1500.350 ;
        RECT 1102.790 1500.000 1103.070 1500.350 ;
        RECT 544.740 26.190 545.000 26.510 ;
        RECT 545.200 26.190 545.460 26.510 ;
        RECT 1097.200 26.190 1097.460 26.510 ;
        RECT 490.460 25.850 490.720 26.170 ;
        RECT 490.520 2.400 490.660 25.850 ;
        RECT 490.310 -4.800 490.870 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1131.770 1500.420 1132.050 1504.000 ;
        RECT 1131.760 1500.000 1132.050 1500.420 ;
        RECT 1131.760 25.005 1131.900 1500.000 ;
        RECT 507.930 24.635 508.210 25.005 ;
        RECT 1131.690 24.635 1131.970 25.005 ;
        RECT 508.000 2.400 508.140 24.635 ;
        RECT 507.790 -4.800 508.350 2.400 ;
      LAYER via2 ;
        RECT 507.930 24.680 508.210 24.960 ;
        RECT 1131.690 24.680 1131.970 24.960 ;
      LAYER met3 ;
        RECT 507.905 24.970 508.235 24.985 ;
        RECT 1131.665 24.970 1131.995 24.985 ;
        RECT 507.905 24.670 1131.995 24.970 ;
        RECT 507.905 24.655 508.235 24.670 ;
        RECT 1131.665 24.655 1131.995 24.670 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 525.850 26.080 526.170 26.140 ;
        RECT 1159.270 26.080 1159.590 26.140 ;
        RECT 525.850 25.940 1159.590 26.080 ;
        RECT 525.850 25.880 526.170 25.940 ;
        RECT 1159.270 25.880 1159.590 25.940 ;
      LAYER via ;
        RECT 525.880 25.880 526.140 26.140 ;
        RECT 1159.300 25.880 1159.560 26.140 ;
      LAYER met2 ;
        RECT 1161.210 1500.490 1161.490 1504.000 ;
        RECT 1159.360 1500.350 1161.490 1500.490 ;
        RECT 1159.360 26.170 1159.500 1500.350 ;
        RECT 1161.210 1500.000 1161.490 1500.350 ;
        RECT 525.880 25.850 526.140 26.170 ;
        RECT 1159.300 25.850 1159.560 26.170 ;
        RECT 525.940 2.400 526.080 25.850 ;
        RECT 525.730 -4.800 526.290 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 543.790 31.860 544.110 31.920 ;
        RECT 1186.870 31.860 1187.190 31.920 ;
        RECT 543.790 31.720 1187.190 31.860 ;
        RECT 543.790 31.660 544.110 31.720 ;
        RECT 1186.870 31.660 1187.190 31.720 ;
      LAYER via ;
        RECT 543.820 31.660 544.080 31.920 ;
        RECT 1186.900 31.660 1187.160 31.920 ;
      LAYER met2 ;
        RECT 1190.190 1500.490 1190.470 1504.000 ;
        RECT 1186.960 1500.350 1190.470 1500.490 ;
        RECT 1186.960 31.950 1187.100 1500.350 ;
        RECT 1190.190 1500.000 1190.470 1500.350 ;
        RECT 543.820 31.630 544.080 31.950 ;
        RECT 1186.900 31.630 1187.160 31.950 ;
        RECT 543.880 2.400 544.020 31.630 ;
        RECT 543.670 -4.800 544.230 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 561.730 31.520 562.050 31.580 ;
        RECT 1214.470 31.520 1214.790 31.580 ;
        RECT 561.730 31.380 1214.790 31.520 ;
        RECT 561.730 31.320 562.050 31.380 ;
        RECT 1214.470 31.320 1214.790 31.380 ;
      LAYER via ;
        RECT 561.760 31.320 562.020 31.580 ;
        RECT 1214.500 31.320 1214.760 31.580 ;
      LAYER met2 ;
        RECT 1219.170 1500.490 1219.450 1504.000 ;
        RECT 1214.560 1500.350 1219.450 1500.490 ;
        RECT 1214.560 31.610 1214.700 1500.350 ;
        RECT 1219.170 1500.000 1219.450 1500.350 ;
        RECT 561.760 31.290 562.020 31.610 ;
        RECT 1214.500 31.290 1214.760 31.610 ;
        RECT 561.820 2.400 561.960 31.290 ;
        RECT 561.610 -4.800 562.170 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 579.670 31.180 579.990 31.240 ;
        RECT 1242.070 31.180 1242.390 31.240 ;
        RECT 579.670 31.040 1242.390 31.180 ;
        RECT 579.670 30.980 579.990 31.040 ;
        RECT 1242.070 30.980 1242.390 31.040 ;
      LAYER via ;
        RECT 579.700 30.980 579.960 31.240 ;
        RECT 1242.100 30.980 1242.360 31.240 ;
      LAYER met2 ;
        RECT 1248.610 1500.490 1248.890 1504.000 ;
        RECT 1242.160 1500.350 1248.890 1500.490 ;
        RECT 1242.160 31.270 1242.300 1500.350 ;
        RECT 1248.610 1500.000 1248.890 1500.350 ;
        RECT 579.700 30.950 579.960 31.270 ;
        RECT 1242.100 30.950 1242.360 31.270 ;
        RECT 579.760 2.400 579.900 30.950 ;
        RECT 579.550 -4.800 580.110 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 86.090 26.760 86.410 26.820 ;
        RECT 434.770 26.760 435.090 26.820 ;
        RECT 86.090 26.620 435.090 26.760 ;
        RECT 86.090 26.560 86.410 26.620 ;
        RECT 434.770 26.560 435.090 26.620 ;
      LAYER via ;
        RECT 86.120 26.560 86.380 26.820 ;
        RECT 434.800 26.560 435.060 26.820 ;
      LAYER met2 ;
        RECT 440.850 1500.490 441.130 1504.000 ;
        RECT 434.860 1500.350 441.130 1500.490 ;
        RECT 434.860 26.850 435.000 1500.350 ;
        RECT 440.850 1500.000 441.130 1500.350 ;
        RECT 86.120 26.530 86.380 26.850 ;
        RECT 434.800 26.530 435.060 26.850 ;
        RECT 86.180 2.400 86.320 26.530 ;
        RECT 85.970 -4.800 86.530 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 672.590 1488.760 672.910 1488.820 ;
        RECT 1277.490 1488.760 1277.810 1488.820 ;
        RECT 672.590 1488.620 1277.810 1488.760 ;
        RECT 672.590 1488.560 672.910 1488.620 ;
        RECT 1277.490 1488.560 1277.810 1488.620 ;
        RECT 597.150 25.400 597.470 25.460 ;
        RECT 672.590 25.400 672.910 25.460 ;
        RECT 597.150 25.260 672.910 25.400 ;
        RECT 597.150 25.200 597.470 25.260 ;
        RECT 672.590 25.200 672.910 25.260 ;
      LAYER via ;
        RECT 672.620 1488.560 672.880 1488.820 ;
        RECT 1277.520 1488.560 1277.780 1488.820 ;
        RECT 597.180 25.200 597.440 25.460 ;
        RECT 672.620 25.200 672.880 25.460 ;
      LAYER met2 ;
        RECT 1277.590 1500.420 1277.870 1504.000 ;
        RECT 1277.580 1500.000 1277.870 1500.420 ;
        RECT 1277.580 1488.850 1277.720 1500.000 ;
        RECT 672.620 1488.530 672.880 1488.850 ;
        RECT 1277.520 1488.530 1277.780 1488.850 ;
        RECT 672.680 25.490 672.820 1488.530 ;
        RECT 597.180 25.170 597.440 25.490 ;
        RECT 672.620 25.170 672.880 25.490 ;
        RECT 597.240 2.400 597.380 25.170 ;
        RECT 597.030 -4.800 597.590 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 615.090 30.840 615.410 30.900 ;
        RECT 1304.170 30.840 1304.490 30.900 ;
        RECT 615.090 30.700 1304.490 30.840 ;
        RECT 615.090 30.640 615.410 30.700 ;
        RECT 1304.170 30.640 1304.490 30.700 ;
      LAYER via ;
        RECT 615.120 30.640 615.380 30.900 ;
        RECT 1304.200 30.640 1304.460 30.900 ;
      LAYER met2 ;
        RECT 1307.030 1500.490 1307.310 1504.000 ;
        RECT 1304.260 1500.350 1307.310 1500.490 ;
        RECT 1304.260 30.930 1304.400 1500.350 ;
        RECT 1307.030 1500.000 1307.310 1500.350 ;
        RECT 615.120 30.610 615.380 30.930 ;
        RECT 1304.200 30.610 1304.460 30.930 ;
        RECT 615.180 2.400 615.320 30.610 ;
        RECT 614.970 -4.800 615.530 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 110.010 26.080 110.330 26.140 ;
        RECT 476.170 26.080 476.490 26.140 ;
        RECT 110.010 25.940 476.490 26.080 ;
        RECT 110.010 25.880 110.330 25.940 ;
        RECT 476.170 25.880 476.490 25.940 ;
      LAYER via ;
        RECT 110.040 25.880 110.300 26.140 ;
        RECT 476.200 25.880 476.460 26.140 ;
      LAYER met2 ;
        RECT 479.490 1500.490 479.770 1504.000 ;
        RECT 476.260 1500.350 479.770 1500.490 ;
        RECT 476.260 26.170 476.400 1500.350 ;
        RECT 479.490 1500.000 479.770 1500.350 ;
        RECT 110.040 25.850 110.300 26.170 ;
        RECT 476.200 25.850 476.460 26.170 ;
        RECT 110.100 13.330 110.240 25.850 ;
        RECT 109.640 13.190 110.240 13.330 ;
        RECT 109.640 2.400 109.780 13.190 ;
        RECT 109.430 -4.800 109.990 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 133.470 25.740 133.790 25.800 ;
        RECT 517.570 25.740 517.890 25.800 ;
        RECT 133.470 25.600 517.890 25.740 ;
        RECT 133.470 25.540 133.790 25.600 ;
        RECT 517.570 25.540 517.890 25.600 ;
      LAYER via ;
        RECT 133.500 25.540 133.760 25.800 ;
        RECT 517.600 25.540 517.860 25.800 ;
      LAYER met2 ;
        RECT 518.590 1500.490 518.870 1504.000 ;
        RECT 517.660 1500.350 518.870 1500.490 ;
        RECT 517.660 25.830 517.800 1500.350 ;
        RECT 518.590 1500.000 518.870 1500.350 ;
        RECT 133.500 25.510 133.760 25.830 ;
        RECT 517.600 25.510 517.860 25.830 ;
        RECT 133.560 2.400 133.700 25.510 ;
        RECT 133.350 -4.800 133.910 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 151.410 25.400 151.730 25.460 ;
        RECT 545.630 25.400 545.950 25.460 ;
        RECT 151.410 25.260 545.950 25.400 ;
        RECT 151.410 25.200 151.730 25.260 ;
        RECT 545.630 25.200 545.950 25.260 ;
      LAYER via ;
        RECT 151.440 25.200 151.700 25.460 ;
        RECT 545.660 25.200 545.920 25.460 ;
      LAYER met2 ;
        RECT 547.570 1500.490 547.850 1504.000 ;
        RECT 545.260 1500.350 547.850 1500.490 ;
        RECT 545.260 28.290 545.400 1500.350 ;
        RECT 547.570 1500.000 547.850 1500.350 ;
        RECT 545.260 28.150 545.860 28.290 ;
        RECT 545.720 25.490 545.860 28.150 ;
        RECT 151.440 25.170 151.700 25.490 ;
        RECT 545.660 25.170 545.920 25.490 ;
        RECT 151.500 2.400 151.640 25.170 ;
        RECT 151.290 -4.800 151.850 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 169.350 25.060 169.670 25.120 ;
        RECT 572.770 25.060 573.090 25.120 ;
        RECT 169.350 24.920 573.090 25.060 ;
        RECT 169.350 24.860 169.670 24.920 ;
        RECT 572.770 24.860 573.090 24.920 ;
      LAYER via ;
        RECT 169.380 24.860 169.640 25.120 ;
        RECT 572.800 24.860 573.060 25.120 ;
      LAYER met2 ;
        RECT 577.010 1500.490 577.290 1504.000 ;
        RECT 572.860 1500.350 577.290 1500.490 ;
        RECT 572.860 25.150 573.000 1500.350 ;
        RECT 577.010 1500.000 577.290 1500.350 ;
        RECT 169.380 24.830 169.640 25.150 ;
        RECT 572.800 24.830 573.060 25.150 ;
        RECT 169.440 2.400 169.580 24.830 ;
        RECT 169.230 -4.800 169.790 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 186.830 24.720 187.150 24.780 ;
        RECT 600.370 24.720 600.690 24.780 ;
        RECT 186.830 24.580 600.690 24.720 ;
        RECT 186.830 24.520 187.150 24.580 ;
        RECT 600.370 24.520 600.690 24.580 ;
      LAYER via ;
        RECT 186.860 24.520 187.120 24.780 ;
        RECT 600.400 24.520 600.660 24.780 ;
      LAYER met2 ;
        RECT 605.990 1500.490 606.270 1504.000 ;
        RECT 600.460 1500.350 606.270 1500.490 ;
        RECT 600.460 24.810 600.600 1500.350 ;
        RECT 605.990 1500.000 606.270 1500.350 ;
        RECT 186.860 24.490 187.120 24.810 ;
        RECT 600.400 24.490 600.660 24.810 ;
        RECT 186.920 2.400 187.060 24.490 ;
        RECT 186.710 -4.800 187.270 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 204.770 24.380 205.090 24.440 ;
        RECT 634.870 24.380 635.190 24.440 ;
        RECT 204.770 24.240 635.190 24.380 ;
        RECT 204.770 24.180 205.090 24.240 ;
        RECT 634.870 24.180 635.190 24.240 ;
      LAYER via ;
        RECT 204.800 24.180 205.060 24.440 ;
        RECT 634.900 24.180 635.160 24.440 ;
      LAYER met2 ;
        RECT 635.430 1500.490 635.710 1504.000 ;
        RECT 634.960 1500.350 635.710 1500.490 ;
        RECT 634.960 24.470 635.100 1500.350 ;
        RECT 635.430 1500.000 635.710 1500.350 ;
        RECT 204.800 24.150 205.060 24.470 ;
        RECT 634.900 24.150 635.160 24.470 ;
        RECT 204.860 2.400 205.000 24.150 ;
        RECT 204.650 -4.800 205.210 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 222.710 24.040 223.030 24.100 ;
        RECT 662.470 24.040 662.790 24.100 ;
        RECT 222.710 23.900 662.790 24.040 ;
        RECT 222.710 23.840 223.030 23.900 ;
        RECT 662.470 23.840 662.790 23.900 ;
      LAYER via ;
        RECT 222.740 23.840 223.000 24.100 ;
        RECT 662.500 23.840 662.760 24.100 ;
      LAYER met2 ;
        RECT 664.410 1500.490 664.690 1504.000 ;
        RECT 662.560 1500.350 664.690 1500.490 ;
        RECT 662.560 24.130 662.700 1500.350 ;
        RECT 664.410 1500.000 664.690 1500.350 ;
        RECT 222.740 23.810 223.000 24.130 ;
        RECT 662.500 23.810 662.760 24.130 ;
        RECT 222.800 2.400 222.940 23.810 ;
        RECT 222.590 -4.800 223.150 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 19.850 20.640 20.170 20.700 ;
        RECT 305.510 20.640 305.830 20.700 ;
        RECT 19.850 20.500 305.830 20.640 ;
        RECT 19.850 20.440 20.170 20.500 ;
        RECT 305.510 20.440 305.830 20.500 ;
        RECT 305.510 17.240 305.830 17.300 ;
        RECT 331.270 17.240 331.590 17.300 ;
        RECT 305.510 17.100 331.590 17.240 ;
        RECT 305.510 17.040 305.830 17.100 ;
        RECT 331.270 17.040 331.590 17.100 ;
      LAYER via ;
        RECT 19.880 20.440 20.140 20.700 ;
        RECT 305.540 20.440 305.800 20.700 ;
        RECT 305.540 17.040 305.800 17.300 ;
        RECT 331.300 17.040 331.560 17.300 ;
      LAYER met2 ;
        RECT 333.670 1500.490 333.950 1504.000 ;
        RECT 331.360 1500.350 333.950 1500.490 ;
        RECT 19.880 20.410 20.140 20.730 ;
        RECT 305.540 20.410 305.800 20.730 ;
        RECT 19.940 10.610 20.080 20.410 ;
        RECT 305.600 17.330 305.740 20.410 ;
        RECT 331.360 17.330 331.500 1500.350 ;
        RECT 333.670 1500.000 333.950 1500.350 ;
        RECT 305.540 17.010 305.800 17.330 ;
        RECT 331.300 17.010 331.560 17.330 ;
        RECT 19.940 10.470 20.540 10.610 ;
        RECT 20.400 2.400 20.540 10.470 ;
        RECT 20.190 -4.800 20.750 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 44.230 20.300 44.550 20.360 ;
        RECT 372.670 20.300 372.990 20.360 ;
        RECT 44.230 20.160 372.990 20.300 ;
        RECT 44.230 20.100 44.550 20.160 ;
        RECT 372.670 20.100 372.990 20.160 ;
      LAYER via ;
        RECT 44.260 20.100 44.520 20.360 ;
        RECT 372.700 20.100 372.960 20.360 ;
      LAYER met2 ;
        RECT 372.770 1500.420 373.050 1504.000 ;
        RECT 372.760 1500.000 373.050 1500.420 ;
        RECT 372.760 20.390 372.900 1500.000 ;
        RECT 44.260 20.070 44.520 20.390 ;
        RECT 372.700 20.070 372.960 20.390 ;
        RECT 44.320 2.400 44.460 20.070 ;
        RECT 44.110 -4.800 44.670 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 246.630 14.860 246.950 14.920 ;
        RECT 696.970 14.860 697.290 14.920 ;
        RECT 246.630 14.720 697.290 14.860 ;
        RECT 246.630 14.660 246.950 14.720 ;
        RECT 696.970 14.660 697.290 14.720 ;
      LAYER via ;
        RECT 246.660 14.660 246.920 14.920 ;
        RECT 697.000 14.660 697.260 14.920 ;
      LAYER met2 ;
        RECT 703.510 1500.490 703.790 1504.000 ;
        RECT 697.060 1500.350 703.790 1500.490 ;
        RECT 697.060 14.950 697.200 1500.350 ;
        RECT 703.510 1500.000 703.790 1500.350 ;
        RECT 246.660 14.630 246.920 14.950 ;
        RECT 697.000 14.630 697.260 14.950 ;
        RECT 246.720 2.400 246.860 14.630 ;
        RECT 246.510 -4.800 247.070 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 624.290 1484.000 624.610 1484.060 ;
        RECT 732.850 1484.000 733.170 1484.060 ;
        RECT 624.290 1483.860 733.170 1484.000 ;
        RECT 624.290 1483.800 624.610 1483.860 ;
        RECT 732.850 1483.800 733.170 1483.860 ;
        RECT 469.270 27.780 469.590 27.840 ;
        RECT 497.330 27.780 497.650 27.840 ;
        RECT 469.270 27.640 497.650 27.780 ;
        RECT 469.270 27.580 469.590 27.640 ;
        RECT 497.330 27.580 497.650 27.640 ;
        RECT 359.330 27.440 359.650 27.500 ;
        RECT 359.330 27.300 400.960 27.440 ;
        RECT 359.330 27.240 359.650 27.300 ;
        RECT 400.820 27.100 400.960 27.300 ;
        RECT 418.670 27.100 418.990 27.160 ;
        RECT 400.820 26.960 418.990 27.100 ;
        RECT 418.670 26.900 418.990 26.960 ;
        RECT 327.590 26.420 327.910 26.480 ;
        RECT 359.330 26.420 359.650 26.480 ;
        RECT 327.590 26.280 359.650 26.420 ;
        RECT 327.590 26.220 327.910 26.280 ;
        RECT 359.330 26.220 359.650 26.280 ;
        RECT 420.510 26.420 420.830 26.480 ;
        RECT 469.270 26.420 469.590 26.480 ;
        RECT 420.510 26.280 469.590 26.420 ;
        RECT 420.510 26.220 420.830 26.280 ;
        RECT 469.270 26.220 469.590 26.280 ;
        RECT 497.330 26.080 497.650 26.140 ;
        RECT 497.330 25.940 520.560 26.080 ;
        RECT 497.330 25.880 497.650 25.940 ;
        RECT 520.420 25.740 520.560 25.940 ;
        RECT 624.290 25.740 624.610 25.800 ;
        RECT 520.420 25.600 624.610 25.740 ;
        RECT 624.290 25.540 624.610 25.600 ;
        RECT 264.110 23.700 264.430 23.760 ;
        RECT 327.590 23.700 327.910 23.760 ;
        RECT 264.110 23.560 327.910 23.700 ;
        RECT 264.110 23.500 264.430 23.560 ;
        RECT 327.590 23.500 327.910 23.560 ;
      LAYER via ;
        RECT 624.320 1483.800 624.580 1484.060 ;
        RECT 732.880 1483.800 733.140 1484.060 ;
        RECT 469.300 27.580 469.560 27.840 ;
        RECT 497.360 27.580 497.620 27.840 ;
        RECT 359.360 27.240 359.620 27.500 ;
        RECT 418.700 26.900 418.960 27.160 ;
        RECT 327.620 26.220 327.880 26.480 ;
        RECT 359.360 26.220 359.620 26.480 ;
        RECT 420.540 26.220 420.800 26.480 ;
        RECT 469.300 26.220 469.560 26.480 ;
        RECT 497.360 25.880 497.620 26.140 ;
        RECT 624.320 25.540 624.580 25.800 ;
        RECT 264.140 23.500 264.400 23.760 ;
        RECT 327.620 23.500 327.880 23.760 ;
      LAYER met2 ;
        RECT 732.950 1500.420 733.230 1504.000 ;
        RECT 732.940 1500.000 733.230 1500.420 ;
        RECT 732.940 1484.090 733.080 1500.000 ;
        RECT 624.320 1483.770 624.580 1484.090 ;
        RECT 732.880 1483.770 733.140 1484.090 ;
        RECT 359.360 27.210 359.620 27.530 ;
        RECT 418.760 27.470 419.820 27.610 ;
        RECT 469.300 27.550 469.560 27.870 ;
        RECT 497.360 27.550 497.620 27.870 ;
        RECT 359.420 26.510 359.560 27.210 ;
        RECT 418.760 27.190 418.900 27.470 ;
        RECT 418.700 26.870 418.960 27.190 ;
        RECT 419.680 26.930 419.820 27.470 ;
        RECT 419.680 26.790 420.740 26.930 ;
        RECT 420.600 26.510 420.740 26.790 ;
        RECT 469.360 26.510 469.500 27.550 ;
        RECT 327.620 26.190 327.880 26.510 ;
        RECT 359.360 26.190 359.620 26.510 ;
        RECT 420.540 26.190 420.800 26.510 ;
        RECT 469.300 26.190 469.560 26.510 ;
        RECT 327.680 23.790 327.820 26.190 ;
        RECT 497.420 26.170 497.560 27.550 ;
        RECT 497.360 25.850 497.620 26.170 ;
        RECT 624.380 25.830 624.520 1483.770 ;
        RECT 624.320 25.510 624.580 25.830 ;
        RECT 264.140 23.470 264.400 23.790 ;
        RECT 327.620 23.470 327.880 23.790 ;
        RECT 264.200 2.400 264.340 23.470 ;
        RECT 263.990 -4.800 264.550 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 282.050 15.540 282.370 15.600 ;
        RECT 759.070 15.540 759.390 15.600 ;
        RECT 282.050 15.400 759.390 15.540 ;
        RECT 282.050 15.340 282.370 15.400 ;
        RECT 759.070 15.340 759.390 15.400 ;
      LAYER via ;
        RECT 282.080 15.340 282.340 15.600 ;
        RECT 759.100 15.340 759.360 15.600 ;
      LAYER met2 ;
        RECT 761.930 1500.490 762.210 1504.000 ;
        RECT 759.160 1500.350 762.210 1500.490 ;
        RECT 759.160 15.630 759.300 1500.350 ;
        RECT 761.930 1500.000 762.210 1500.350 ;
        RECT 282.080 15.310 282.340 15.630 ;
        RECT 759.100 15.310 759.360 15.630 ;
        RECT 282.140 2.400 282.280 15.310 ;
        RECT 281.930 -4.800 282.490 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 299.990 32.200 300.310 32.260 ;
        RECT 786.670 32.200 786.990 32.260 ;
        RECT 299.990 32.060 786.990 32.200 ;
        RECT 299.990 32.000 300.310 32.060 ;
        RECT 786.670 32.000 786.990 32.060 ;
      LAYER via ;
        RECT 300.020 32.000 300.280 32.260 ;
        RECT 786.700 32.000 786.960 32.260 ;
      LAYER met2 ;
        RECT 790.910 1500.490 791.190 1504.000 ;
        RECT 786.760 1500.350 791.190 1500.490 ;
        RECT 786.760 32.290 786.900 1500.350 ;
        RECT 790.910 1500.000 791.190 1500.350 ;
        RECT 300.020 31.970 300.280 32.290 ;
        RECT 786.700 31.970 786.960 32.290 ;
        RECT 300.080 2.400 300.220 31.970 ;
        RECT 299.870 -4.800 300.430 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 317.930 16.900 318.250 16.960 ;
        RECT 320.690 16.900 321.010 16.960 ;
        RECT 317.930 16.760 321.010 16.900 ;
        RECT 317.930 16.700 318.250 16.760 ;
        RECT 320.690 16.700 321.010 16.760 ;
        RECT 320.690 16.220 321.010 16.280 ;
        RECT 814.270 16.220 814.590 16.280 ;
        RECT 320.690 16.080 814.590 16.220 ;
        RECT 320.690 16.020 321.010 16.080 ;
        RECT 814.270 16.020 814.590 16.080 ;
      LAYER via ;
        RECT 317.960 16.700 318.220 16.960 ;
        RECT 320.720 16.700 320.980 16.960 ;
        RECT 320.720 16.020 320.980 16.280 ;
        RECT 814.300 16.020 814.560 16.280 ;
      LAYER met2 ;
        RECT 820.350 1500.490 820.630 1504.000 ;
        RECT 814.360 1500.350 820.630 1500.490 ;
        RECT 317.960 16.670 318.220 16.990 ;
        RECT 320.720 16.670 320.980 16.990 ;
        RECT 318.020 2.400 318.160 16.670 ;
        RECT 320.780 16.310 320.920 16.670 ;
        RECT 814.360 16.310 814.500 1500.350 ;
        RECT 820.350 1500.000 820.630 1500.350 ;
        RECT 320.720 15.990 320.980 16.310 ;
        RECT 814.300 15.990 814.560 16.310 ;
        RECT 317.810 -4.800 318.370 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 337.710 1485.700 338.030 1485.760 ;
        RECT 849.230 1485.700 849.550 1485.760 ;
        RECT 337.710 1485.560 849.550 1485.700 ;
        RECT 337.710 1485.500 338.030 1485.560 ;
        RECT 849.230 1485.500 849.550 1485.560 ;
        RECT 337.710 1401.860 338.030 1402.120 ;
        RECT 337.800 1401.440 337.940 1401.860 ;
        RECT 337.710 1401.180 338.030 1401.440 ;
        RECT 336.790 1159.100 337.110 1159.360 ;
        RECT 336.880 1158.680 337.020 1159.100 ;
        RECT 336.790 1158.420 337.110 1158.680 ;
        RECT 336.330 1152.160 336.650 1152.220 ;
        RECT 336.790 1152.160 337.110 1152.220 ;
        RECT 336.330 1152.020 337.110 1152.160 ;
        RECT 336.330 1151.960 336.650 1152.020 ;
        RECT 336.790 1151.960 337.110 1152.020 ;
        RECT 336.330 1104.220 336.650 1104.280 ;
        RECT 337.710 1104.220 338.030 1104.280 ;
        RECT 336.330 1104.080 338.030 1104.220 ;
        RECT 336.330 1104.020 336.650 1104.080 ;
        RECT 337.710 1104.020 338.030 1104.080 ;
        RECT 337.710 1062.740 338.030 1062.800 ;
        RECT 337.340 1062.600 338.030 1062.740 ;
        RECT 337.340 1062.460 337.480 1062.600 ;
        RECT 337.710 1062.540 338.030 1062.600 ;
        RECT 337.250 1062.200 337.570 1062.460 ;
        RECT 337.250 1055.600 337.570 1055.660 ;
        RECT 337.710 1055.600 338.030 1055.660 ;
        RECT 337.250 1055.460 338.030 1055.600 ;
        RECT 337.250 1055.400 337.570 1055.460 ;
        RECT 337.710 1055.400 338.030 1055.460 ;
        RECT 337.710 1014.260 338.030 1014.520 ;
        RECT 337.250 1014.120 337.570 1014.180 ;
        RECT 337.800 1014.120 337.940 1014.260 ;
        RECT 337.250 1013.980 337.940 1014.120 ;
        RECT 337.250 1013.920 337.570 1013.980 ;
        RECT 337.250 579.600 337.570 579.660 ;
        RECT 337.710 579.600 338.030 579.660 ;
        RECT 337.250 579.460 338.030 579.600 ;
        RECT 337.250 579.400 337.570 579.460 ;
        RECT 337.710 579.400 338.030 579.460 ;
        RECT 336.330 572.460 336.650 572.520 ;
        RECT 337.250 572.460 337.570 572.520 ;
        RECT 336.330 572.320 337.570 572.460 ;
        RECT 336.330 572.260 336.650 572.320 ;
        RECT 337.250 572.260 337.570 572.320 ;
        RECT 336.330 524.520 336.650 524.580 ;
        RECT 337.710 524.520 338.030 524.580 ;
        RECT 336.330 524.380 338.030 524.520 ;
        RECT 336.330 524.320 336.650 524.380 ;
        RECT 337.710 524.320 338.030 524.380 ;
        RECT 337.250 289.580 337.570 289.640 ;
        RECT 337.710 289.580 338.030 289.640 ;
        RECT 337.250 289.440 338.030 289.580 ;
        RECT 337.250 289.380 337.570 289.440 ;
        RECT 337.710 289.380 338.030 289.440 ;
        RECT 336.330 282.780 336.650 282.840 ;
        RECT 337.250 282.780 337.570 282.840 ;
        RECT 336.330 282.640 337.570 282.780 ;
        RECT 336.330 282.580 336.650 282.640 ;
        RECT 337.250 282.580 337.570 282.640 ;
        RECT 336.330 234.840 336.650 234.900 ;
        RECT 337.710 234.840 338.030 234.900 ;
        RECT 336.330 234.700 338.030 234.840 ;
        RECT 336.330 234.640 336.650 234.700 ;
        RECT 337.710 234.640 338.030 234.700 ;
        RECT 337.250 186.560 337.570 186.620 ;
        RECT 337.710 186.560 338.030 186.620 ;
        RECT 337.250 186.420 338.030 186.560 ;
        RECT 337.250 186.360 337.570 186.420 ;
        RECT 337.710 186.360 338.030 186.420 ;
        RECT 337.710 138.280 338.030 138.340 ;
        RECT 338.630 138.280 338.950 138.340 ;
        RECT 337.710 138.140 338.950 138.280 ;
        RECT 337.710 138.080 338.030 138.140 ;
        RECT 338.630 138.080 338.950 138.140 ;
        RECT 337.710 96.260 338.030 96.520 ;
        RECT 334.950 96.120 335.270 96.180 ;
        RECT 337.800 96.120 337.940 96.260 ;
        RECT 334.950 95.980 337.940 96.120 ;
        RECT 334.950 95.920 335.270 95.980 ;
      LAYER via ;
        RECT 337.740 1485.500 338.000 1485.760 ;
        RECT 849.260 1485.500 849.520 1485.760 ;
        RECT 337.740 1401.860 338.000 1402.120 ;
        RECT 337.740 1401.180 338.000 1401.440 ;
        RECT 336.820 1159.100 337.080 1159.360 ;
        RECT 336.820 1158.420 337.080 1158.680 ;
        RECT 336.360 1151.960 336.620 1152.220 ;
        RECT 336.820 1151.960 337.080 1152.220 ;
        RECT 336.360 1104.020 336.620 1104.280 ;
        RECT 337.740 1104.020 338.000 1104.280 ;
        RECT 337.740 1062.540 338.000 1062.800 ;
        RECT 337.280 1062.200 337.540 1062.460 ;
        RECT 337.280 1055.400 337.540 1055.660 ;
        RECT 337.740 1055.400 338.000 1055.660 ;
        RECT 337.740 1014.260 338.000 1014.520 ;
        RECT 337.280 1013.920 337.540 1014.180 ;
        RECT 337.280 579.400 337.540 579.660 ;
        RECT 337.740 579.400 338.000 579.660 ;
        RECT 336.360 572.260 336.620 572.520 ;
        RECT 337.280 572.260 337.540 572.520 ;
        RECT 336.360 524.320 336.620 524.580 ;
        RECT 337.740 524.320 338.000 524.580 ;
        RECT 337.280 289.380 337.540 289.640 ;
        RECT 337.740 289.380 338.000 289.640 ;
        RECT 336.360 282.580 336.620 282.840 ;
        RECT 337.280 282.580 337.540 282.840 ;
        RECT 336.360 234.640 336.620 234.900 ;
        RECT 337.740 234.640 338.000 234.900 ;
        RECT 337.280 186.360 337.540 186.620 ;
        RECT 337.740 186.360 338.000 186.620 ;
        RECT 337.740 138.080 338.000 138.340 ;
        RECT 338.660 138.080 338.920 138.340 ;
        RECT 337.740 96.260 338.000 96.520 ;
        RECT 334.980 95.920 335.240 96.180 ;
      LAYER met2 ;
        RECT 849.330 1500.420 849.610 1504.000 ;
        RECT 849.320 1500.000 849.610 1500.420 ;
        RECT 849.320 1485.790 849.460 1500.000 ;
        RECT 337.740 1485.470 338.000 1485.790 ;
        RECT 849.260 1485.470 849.520 1485.790 ;
        RECT 337.800 1402.150 337.940 1485.470 ;
        RECT 337.740 1401.830 338.000 1402.150 ;
        RECT 337.740 1401.150 338.000 1401.470 ;
        RECT 337.800 1200.725 337.940 1401.150 ;
        RECT 336.810 1200.355 337.090 1200.725 ;
        RECT 337.730 1200.355 338.010 1200.725 ;
        RECT 336.880 1159.390 337.020 1200.355 ;
        RECT 336.820 1159.070 337.080 1159.390 ;
        RECT 336.820 1158.390 337.080 1158.710 ;
        RECT 336.880 1152.250 337.020 1158.390 ;
        RECT 336.360 1151.930 336.620 1152.250 ;
        RECT 336.820 1151.930 337.080 1152.250 ;
        RECT 336.420 1104.310 336.560 1151.930 ;
        RECT 336.360 1103.990 336.620 1104.310 ;
        RECT 337.740 1103.990 338.000 1104.310 ;
        RECT 337.800 1062.830 337.940 1103.990 ;
        RECT 337.740 1062.510 338.000 1062.830 ;
        RECT 337.280 1062.170 337.540 1062.490 ;
        RECT 337.340 1055.690 337.480 1062.170 ;
        RECT 337.280 1055.370 337.540 1055.690 ;
        RECT 337.740 1055.370 338.000 1055.690 ;
        RECT 337.800 1014.550 337.940 1055.370 ;
        RECT 337.740 1014.230 338.000 1014.550 ;
        RECT 337.280 1013.890 337.540 1014.210 ;
        RECT 337.340 1007.490 337.480 1013.890 ;
        RECT 337.340 1007.350 337.940 1007.490 ;
        RECT 337.800 886.565 337.940 1007.350 ;
        RECT 337.730 886.195 338.010 886.565 ;
        RECT 337.730 820.915 338.010 821.285 ;
        RECT 337.800 630.205 337.940 820.915 ;
        RECT 337.730 629.835 338.010 630.205 ;
        RECT 337.730 627.795 338.010 628.165 ;
        RECT 337.800 579.690 337.940 627.795 ;
        RECT 337.280 579.370 337.540 579.690 ;
        RECT 337.740 579.370 338.000 579.690 ;
        RECT 337.340 572.550 337.480 579.370 ;
        RECT 336.360 572.230 336.620 572.550 ;
        RECT 337.280 572.230 337.540 572.550 ;
        RECT 336.420 524.610 336.560 572.230 ;
        RECT 336.360 524.290 336.620 524.610 ;
        RECT 337.740 524.290 338.000 524.610 ;
        RECT 337.800 289.670 337.940 524.290 ;
        RECT 337.280 289.350 337.540 289.670 ;
        RECT 337.740 289.350 338.000 289.670 ;
        RECT 337.340 282.870 337.480 289.350 ;
        RECT 336.360 282.550 336.620 282.870 ;
        RECT 337.280 282.550 337.540 282.870 ;
        RECT 336.420 234.930 336.560 282.550 ;
        RECT 336.360 234.610 336.620 234.930 ;
        RECT 337.740 234.610 338.000 234.930 ;
        RECT 337.800 186.650 337.940 234.610 ;
        RECT 337.280 186.330 337.540 186.650 ;
        RECT 337.740 186.330 338.000 186.650 ;
        RECT 337.340 186.165 337.480 186.330 ;
        RECT 337.270 185.795 337.550 186.165 ;
        RECT 338.650 185.795 338.930 186.165 ;
        RECT 338.720 138.370 338.860 185.795 ;
        RECT 337.740 138.050 338.000 138.370 ;
        RECT 338.660 138.050 338.920 138.370 ;
        RECT 337.800 96.550 337.940 138.050 ;
        RECT 337.740 96.230 338.000 96.550 ;
        RECT 334.980 95.890 335.240 96.210 ;
        RECT 335.040 24.210 335.180 95.890 ;
        RECT 335.040 24.070 336.100 24.210 ;
        RECT 335.960 2.400 336.100 24.070 ;
        RECT 335.750 -4.800 336.310 2.400 ;
      LAYER via2 ;
        RECT 336.810 1200.400 337.090 1200.680 ;
        RECT 337.730 1200.400 338.010 1200.680 ;
        RECT 337.730 886.240 338.010 886.520 ;
        RECT 337.730 820.960 338.010 821.240 ;
        RECT 337.730 629.880 338.010 630.160 ;
        RECT 337.730 627.840 338.010 628.120 ;
        RECT 337.270 185.840 337.550 186.120 ;
        RECT 338.650 185.840 338.930 186.120 ;
      LAYER met3 ;
        RECT 336.785 1200.690 337.115 1200.705 ;
        RECT 337.705 1200.690 338.035 1200.705 ;
        RECT 336.785 1200.390 338.035 1200.690 ;
        RECT 336.785 1200.375 337.115 1200.390 ;
        RECT 337.705 1200.375 338.035 1200.390 ;
        RECT 336.990 886.530 337.370 886.540 ;
        RECT 337.705 886.530 338.035 886.545 ;
        RECT 336.990 886.230 338.035 886.530 ;
        RECT 336.990 886.220 337.370 886.230 ;
        RECT 337.705 886.215 338.035 886.230 ;
        RECT 336.990 821.250 337.370 821.260 ;
        RECT 337.705 821.250 338.035 821.265 ;
        RECT 336.990 820.950 338.035 821.250 ;
        RECT 336.990 820.940 337.370 820.950 ;
        RECT 337.705 820.935 338.035 820.950 ;
        RECT 336.990 630.170 337.370 630.180 ;
        RECT 337.705 630.170 338.035 630.185 ;
        RECT 336.990 629.870 338.035 630.170 ;
        RECT 336.990 629.860 337.370 629.870 ;
        RECT 337.705 629.855 338.035 629.870 ;
        RECT 336.990 628.130 337.370 628.140 ;
        RECT 337.705 628.130 338.035 628.145 ;
        RECT 336.990 627.830 338.035 628.130 ;
        RECT 336.990 627.820 337.370 627.830 ;
        RECT 337.705 627.815 338.035 627.830 ;
        RECT 337.245 186.130 337.575 186.145 ;
        RECT 338.625 186.130 338.955 186.145 ;
        RECT 337.245 185.830 338.955 186.130 ;
        RECT 337.245 185.815 337.575 185.830 ;
        RECT 338.625 185.815 338.955 185.830 ;
      LAYER via3 ;
        RECT 337.020 886.220 337.340 886.540 ;
        RECT 337.020 820.940 337.340 821.260 ;
        RECT 337.020 629.860 337.340 630.180 ;
        RECT 337.020 627.820 337.340 628.140 ;
      LAYER met4 ;
        RECT 337.015 886.215 337.345 886.545 ;
        RECT 337.030 821.265 337.330 886.215 ;
        RECT 337.015 820.935 337.345 821.265 ;
        RECT 337.015 629.855 337.345 630.185 ;
        RECT 337.030 628.145 337.330 629.855 ;
        RECT 337.015 627.815 337.345 628.145 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 366.230 16.900 366.550 16.960 ;
        RECT 876.370 16.900 876.690 16.960 ;
        RECT 366.230 16.760 876.690 16.900 ;
        RECT 366.230 16.700 366.550 16.760 ;
        RECT 876.370 16.700 876.690 16.760 ;
        RECT 353.350 5.680 353.670 5.740 ;
        RECT 366.230 5.680 366.550 5.740 ;
        RECT 353.350 5.540 366.550 5.680 ;
        RECT 353.350 5.480 353.670 5.540 ;
        RECT 366.230 5.480 366.550 5.540 ;
      LAYER via ;
        RECT 366.260 16.700 366.520 16.960 ;
        RECT 876.400 16.700 876.660 16.960 ;
        RECT 353.380 5.480 353.640 5.740 ;
        RECT 366.260 5.480 366.520 5.740 ;
      LAYER met2 ;
        RECT 878.770 1500.490 879.050 1504.000 ;
        RECT 876.460 1500.350 879.050 1500.490 ;
        RECT 876.460 16.990 876.600 1500.350 ;
        RECT 878.770 1500.000 879.050 1500.350 ;
        RECT 366.260 16.670 366.520 16.990 ;
        RECT 876.400 16.670 876.660 16.990 ;
        RECT 366.320 5.770 366.460 16.670 ;
        RECT 353.380 5.450 353.640 5.770 ;
        RECT 366.260 5.450 366.520 5.770 ;
        RECT 353.440 2.400 353.580 5.450 ;
        RECT 353.230 -4.800 353.790 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 372.210 1486.380 372.530 1486.440 ;
        RECT 907.650 1486.380 907.970 1486.440 ;
        RECT 372.210 1486.240 907.970 1486.380 ;
        RECT 372.210 1486.180 372.530 1486.240 ;
        RECT 907.650 1486.180 907.970 1486.240 ;
      LAYER via ;
        RECT 372.240 1486.180 372.500 1486.440 ;
        RECT 907.680 1486.180 907.940 1486.440 ;
      LAYER met2 ;
        RECT 907.750 1500.420 908.030 1504.000 ;
        RECT 907.740 1500.000 908.030 1500.420 ;
        RECT 907.740 1486.470 907.880 1500.000 ;
        RECT 372.240 1486.150 372.500 1486.470 ;
        RECT 907.680 1486.150 907.940 1486.470 ;
        RECT 372.300 17.240 372.440 1486.150 ;
        RECT 371.380 17.100 372.440 17.240 ;
        RECT 371.380 2.400 371.520 17.100 ;
        RECT 371.170 -4.800 371.730 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 407.720 20.500 414.760 20.640 ;
        RECT 389.230 20.300 389.550 20.360 ;
        RECT 407.720 20.300 407.860 20.500 ;
        RECT 389.230 20.160 407.860 20.300 ;
        RECT 414.620 20.300 414.760 20.500 ;
        RECT 931.570 20.300 931.890 20.360 ;
        RECT 414.620 20.160 931.890 20.300 ;
        RECT 389.230 20.100 389.550 20.160 ;
        RECT 931.570 20.100 931.890 20.160 ;
      LAYER via ;
        RECT 389.260 20.100 389.520 20.360 ;
        RECT 931.600 20.100 931.860 20.360 ;
      LAYER met2 ;
        RECT 937.190 1500.490 937.470 1504.000 ;
        RECT 931.660 1500.350 937.470 1500.490 ;
        RECT 931.660 20.390 931.800 1500.350 ;
        RECT 937.190 1500.000 937.470 1500.350 ;
        RECT 389.260 20.070 389.520 20.390 ;
        RECT 931.600 20.070 931.860 20.390 ;
        RECT 389.320 2.400 389.460 20.070 ;
        RECT 389.110 -4.800 389.670 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 413.610 1490.460 413.930 1490.520 ;
        RECT 966.070 1490.460 966.390 1490.520 ;
        RECT 413.610 1490.320 966.390 1490.460 ;
        RECT 413.610 1490.260 413.930 1490.320 ;
        RECT 966.070 1490.260 966.390 1490.320 ;
        RECT 407.170 19.960 407.490 20.020 ;
        RECT 413.610 19.960 413.930 20.020 ;
        RECT 407.170 19.820 413.930 19.960 ;
        RECT 407.170 19.760 407.490 19.820 ;
        RECT 413.610 19.760 413.930 19.820 ;
      LAYER via ;
        RECT 413.640 1490.260 413.900 1490.520 ;
        RECT 966.100 1490.260 966.360 1490.520 ;
        RECT 407.200 19.760 407.460 20.020 ;
        RECT 413.640 19.760 413.900 20.020 ;
      LAYER met2 ;
        RECT 966.170 1500.420 966.450 1504.000 ;
        RECT 966.160 1500.000 966.450 1500.420 ;
        RECT 966.160 1490.550 966.300 1500.000 ;
        RECT 413.640 1490.230 413.900 1490.550 ;
        RECT 966.100 1490.230 966.360 1490.550 ;
        RECT 413.700 20.050 413.840 1490.230 ;
        RECT 407.200 19.730 407.460 20.050 ;
        RECT 413.640 19.730 413.900 20.050 ;
        RECT 407.260 2.400 407.400 19.730 ;
        RECT 407.050 -4.800 407.610 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 407.170 20.640 407.490 20.700 ;
        RECT 373.220 20.500 407.490 20.640 ;
        RECT 68.150 19.960 68.470 20.020 ;
        RECT 373.220 19.960 373.360 20.500 ;
        RECT 407.170 20.440 407.490 20.500 ;
        RECT 68.150 19.820 373.360 19.960 ;
        RECT 68.150 19.760 68.470 19.820 ;
      LAYER via ;
        RECT 68.180 19.760 68.440 20.020 ;
        RECT 407.200 20.440 407.460 20.700 ;
      LAYER met2 ;
        RECT 411.410 1500.490 411.690 1504.000 ;
        RECT 407.260 1500.350 411.690 1500.490 ;
        RECT 407.260 20.730 407.400 1500.350 ;
        RECT 411.410 1500.000 411.690 1500.350 ;
        RECT 407.200 20.410 407.460 20.730 ;
        RECT 68.180 19.730 68.440 20.050 ;
        RECT 68.240 2.400 68.380 19.730 ;
        RECT 68.030 -4.800 68.590 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 995.610 1500.490 995.890 1504.000 ;
        RECT 993.760 1500.350 995.890 1500.490 ;
        RECT 993.760 18.885 993.900 1500.350 ;
        RECT 995.610 1500.000 995.890 1500.350 ;
        RECT 424.670 18.515 424.950 18.885 ;
        RECT 993.690 18.515 993.970 18.885 ;
        RECT 424.740 2.400 424.880 18.515 ;
        RECT 424.530 -4.800 425.090 2.400 ;
      LAYER via2 ;
        RECT 424.670 18.560 424.950 18.840 ;
        RECT 993.690 18.560 993.970 18.840 ;
      LAYER met3 ;
        RECT 424.645 18.850 424.975 18.865 ;
        RECT 993.665 18.850 993.995 18.865 ;
        RECT 424.645 18.550 993.995 18.850 ;
        RECT 424.645 18.535 424.975 18.550 ;
        RECT 993.665 18.535 993.995 18.550 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 448.110 1489.780 448.430 1489.840 ;
        RECT 1024.490 1489.780 1024.810 1489.840 ;
        RECT 448.110 1489.640 1024.810 1489.780 ;
        RECT 448.110 1489.580 448.430 1489.640 ;
        RECT 1024.490 1489.580 1024.810 1489.640 ;
        RECT 442.590 19.620 442.910 19.680 ;
        RECT 448.110 19.620 448.430 19.680 ;
        RECT 442.590 19.480 448.430 19.620 ;
        RECT 442.590 19.420 442.910 19.480 ;
        RECT 448.110 19.420 448.430 19.480 ;
      LAYER via ;
        RECT 448.140 1489.580 448.400 1489.840 ;
        RECT 1024.520 1489.580 1024.780 1489.840 ;
        RECT 442.620 19.420 442.880 19.680 ;
        RECT 448.140 19.420 448.400 19.680 ;
      LAYER met2 ;
        RECT 1024.590 1500.420 1024.870 1504.000 ;
        RECT 1024.580 1500.000 1024.870 1500.420 ;
        RECT 1024.580 1489.870 1024.720 1500.000 ;
        RECT 448.140 1489.550 448.400 1489.870 ;
        RECT 1024.520 1489.550 1024.780 1489.870 ;
        RECT 448.200 19.710 448.340 1489.550 ;
        RECT 442.620 19.390 442.880 19.710 ;
        RECT 448.140 19.390 448.400 19.710 ;
        RECT 442.680 2.400 442.820 19.390 ;
        RECT 442.470 -4.800 443.030 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1054.030 1500.490 1054.310 1504.000 ;
        RECT 1048.960 1500.350 1054.310 1500.490 ;
        RECT 1048.960 18.205 1049.100 1500.350 ;
        RECT 1054.030 1500.000 1054.310 1500.350 ;
        RECT 460.550 17.835 460.830 18.205 ;
        RECT 1048.890 17.835 1049.170 18.205 ;
        RECT 460.620 2.400 460.760 17.835 ;
        RECT 460.410 -4.800 460.970 2.400 ;
      LAYER via2 ;
        RECT 460.550 17.880 460.830 18.160 ;
        RECT 1048.890 17.880 1049.170 18.160 ;
      LAYER met3 ;
        RECT 460.525 18.170 460.855 18.185 ;
        RECT 1048.865 18.170 1049.195 18.185 ;
        RECT 460.525 17.870 1049.195 18.170 ;
        RECT 460.525 17.855 460.855 17.870 ;
        RECT 1048.865 17.855 1049.195 17.870 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 482.610 1489.440 482.930 1489.500 ;
        RECT 1082.910 1489.440 1083.230 1489.500 ;
        RECT 482.610 1489.300 1083.230 1489.440 ;
        RECT 482.610 1489.240 482.930 1489.300 ;
        RECT 1082.910 1489.240 1083.230 1489.300 ;
        RECT 478.470 18.940 478.790 19.000 ;
        RECT 482.610 18.940 482.930 19.000 ;
        RECT 478.470 18.800 482.930 18.940 ;
        RECT 478.470 18.740 478.790 18.800 ;
        RECT 482.610 18.740 482.930 18.800 ;
      LAYER via ;
        RECT 482.640 1489.240 482.900 1489.500 ;
        RECT 1082.940 1489.240 1083.200 1489.500 ;
        RECT 478.500 18.740 478.760 19.000 ;
        RECT 482.640 18.740 482.900 19.000 ;
      LAYER met2 ;
        RECT 1083.010 1500.420 1083.290 1504.000 ;
        RECT 1083.000 1500.000 1083.290 1500.420 ;
        RECT 1083.000 1489.530 1083.140 1500.000 ;
        RECT 482.640 1489.210 482.900 1489.530 ;
        RECT 1082.940 1489.210 1083.200 1489.530 ;
        RECT 482.700 19.030 482.840 1489.210 ;
        RECT 478.500 18.710 478.760 19.030 ;
        RECT 482.640 18.710 482.900 19.030 ;
        RECT 478.560 2.400 478.700 18.710 ;
        RECT 478.350 -4.800 478.910 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1112.450 1500.490 1112.730 1504.000 ;
        RECT 1111.060 1500.350 1112.730 1500.490 ;
        RECT 1111.060 17.525 1111.200 1500.350 ;
        RECT 1112.450 1500.000 1112.730 1500.350 ;
        RECT 496.430 17.155 496.710 17.525 ;
        RECT 1110.990 17.155 1111.270 17.525 ;
        RECT 496.500 2.400 496.640 17.155 ;
        RECT 496.290 -4.800 496.850 2.400 ;
      LAYER via2 ;
        RECT 496.430 17.200 496.710 17.480 ;
        RECT 1110.990 17.200 1111.270 17.480 ;
      LAYER met3 ;
        RECT 496.405 17.490 496.735 17.505 ;
        RECT 1110.965 17.490 1111.295 17.505 ;
        RECT 496.405 17.190 1111.295 17.490 ;
        RECT 496.405 17.175 496.735 17.190 ;
        RECT 1110.965 17.175 1111.295 17.190 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 517.110 1488.080 517.430 1488.140 ;
        RECT 1141.330 1488.080 1141.650 1488.140 ;
        RECT 517.110 1487.940 1141.650 1488.080 ;
        RECT 517.110 1487.880 517.430 1487.940 ;
        RECT 1141.330 1487.880 1141.650 1487.940 ;
        RECT 513.890 18.940 514.210 19.000 ;
        RECT 517.110 18.940 517.430 19.000 ;
        RECT 513.890 18.800 517.430 18.940 ;
        RECT 513.890 18.740 514.210 18.800 ;
        RECT 517.110 18.740 517.430 18.800 ;
      LAYER via ;
        RECT 517.140 1487.880 517.400 1488.140 ;
        RECT 1141.360 1487.880 1141.620 1488.140 ;
        RECT 513.920 18.740 514.180 19.000 ;
        RECT 517.140 18.740 517.400 19.000 ;
      LAYER met2 ;
        RECT 1141.430 1500.420 1141.710 1504.000 ;
        RECT 1141.420 1500.000 1141.710 1500.420 ;
        RECT 1141.420 1488.170 1141.560 1500.000 ;
        RECT 517.140 1487.850 517.400 1488.170 ;
        RECT 1141.360 1487.850 1141.620 1488.170 ;
        RECT 517.200 19.030 517.340 1487.850 ;
        RECT 513.920 18.710 514.180 19.030 ;
        RECT 517.140 18.710 517.400 19.030 ;
        RECT 513.980 2.400 514.120 18.710 ;
        RECT 513.770 -4.800 514.330 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 537.810 1487.740 538.130 1487.800 ;
        RECT 1170.770 1487.740 1171.090 1487.800 ;
        RECT 537.810 1487.600 1171.090 1487.740 ;
        RECT 537.810 1487.540 538.130 1487.600 ;
        RECT 1170.770 1487.540 1171.090 1487.600 ;
        RECT 531.830 18.940 532.150 19.000 ;
        RECT 537.810 18.940 538.130 19.000 ;
        RECT 531.830 18.800 538.130 18.940 ;
        RECT 531.830 18.740 532.150 18.800 ;
        RECT 537.810 18.740 538.130 18.800 ;
      LAYER via ;
        RECT 537.840 1487.540 538.100 1487.800 ;
        RECT 1170.800 1487.540 1171.060 1487.800 ;
        RECT 531.860 18.740 532.120 19.000 ;
        RECT 537.840 18.740 538.100 19.000 ;
      LAYER met2 ;
        RECT 1170.870 1500.420 1171.150 1504.000 ;
        RECT 1170.860 1500.000 1171.150 1500.420 ;
        RECT 1170.860 1487.830 1171.000 1500.000 ;
        RECT 537.840 1487.510 538.100 1487.830 ;
        RECT 1170.800 1487.510 1171.060 1487.830 ;
        RECT 537.900 19.030 538.040 1487.510 ;
        RECT 531.860 18.710 532.120 19.030 ;
        RECT 537.840 18.710 538.100 19.030 ;
        RECT 531.920 2.400 532.060 18.710 ;
        RECT 531.710 -4.800 532.270 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1193.770 18.940 1194.090 19.000 ;
        RECT 579.760 18.800 1194.090 18.940 ;
        RECT 549.770 18.260 550.090 18.320 ;
        RECT 579.760 18.260 579.900 18.800 ;
        RECT 1193.770 18.740 1194.090 18.800 ;
        RECT 549.770 18.120 579.900 18.260 ;
        RECT 549.770 18.060 550.090 18.120 ;
      LAYER via ;
        RECT 549.800 18.060 550.060 18.320 ;
        RECT 1193.800 18.740 1194.060 19.000 ;
      LAYER met2 ;
        RECT 1199.850 1500.490 1200.130 1504.000 ;
        RECT 1193.860 1500.350 1200.130 1500.490 ;
        RECT 1193.860 19.030 1194.000 1500.350 ;
        RECT 1199.850 1500.000 1200.130 1500.350 ;
        RECT 1193.800 18.710 1194.060 19.030 ;
        RECT 549.800 18.030 550.060 18.350 ;
        RECT 549.860 2.400 550.000 18.030 ;
        RECT 549.650 -4.800 550.210 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 572.310 1487.060 572.630 1487.120 ;
        RECT 1229.190 1487.060 1229.510 1487.120 ;
        RECT 572.310 1486.920 1229.510 1487.060 ;
        RECT 572.310 1486.860 572.630 1486.920 ;
        RECT 1229.190 1486.860 1229.510 1486.920 ;
        RECT 567.710 18.940 568.030 19.000 ;
        RECT 572.310 18.940 572.630 19.000 ;
        RECT 567.710 18.800 572.630 18.940 ;
        RECT 567.710 18.740 568.030 18.800 ;
        RECT 572.310 18.740 572.630 18.800 ;
      LAYER via ;
        RECT 572.340 1486.860 572.600 1487.120 ;
        RECT 1229.220 1486.860 1229.480 1487.120 ;
        RECT 567.740 18.740 568.000 19.000 ;
        RECT 572.340 18.740 572.600 19.000 ;
      LAYER met2 ;
        RECT 1229.290 1500.420 1229.570 1504.000 ;
        RECT 1229.280 1500.000 1229.570 1500.420 ;
        RECT 1229.280 1487.150 1229.420 1500.000 ;
        RECT 572.340 1486.830 572.600 1487.150 ;
        RECT 1229.220 1486.830 1229.480 1487.150 ;
        RECT 572.400 19.030 572.540 1486.830 ;
        RECT 567.740 18.710 568.000 19.030 ;
        RECT 572.340 18.710 572.600 19.030 ;
        RECT 567.800 2.400 567.940 18.710 ;
        RECT 567.590 -4.800 568.150 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 585.650 18.260 585.970 18.320 ;
        RECT 585.650 18.120 602.900 18.260 ;
        RECT 585.650 18.060 585.970 18.120 ;
        RECT 602.760 17.920 602.900 18.120 ;
        RECT 1255.870 17.920 1256.190 17.980 ;
        RECT 602.760 17.780 613.940 17.920 ;
        RECT 613.800 17.580 613.940 17.780 ;
        RECT 615.180 17.780 1256.190 17.920 ;
        RECT 615.180 17.580 615.320 17.780 ;
        RECT 1255.870 17.720 1256.190 17.780 ;
        RECT 613.800 17.440 615.320 17.580 ;
      LAYER via ;
        RECT 585.680 18.060 585.940 18.320 ;
        RECT 1255.900 17.720 1256.160 17.980 ;
      LAYER met2 ;
        RECT 1258.270 1500.490 1258.550 1504.000 ;
        RECT 1255.960 1500.350 1258.550 1500.490 ;
        RECT 585.680 18.030 585.940 18.350 ;
        RECT 585.740 2.400 585.880 18.030 ;
        RECT 1255.960 18.010 1256.100 1500.350 ;
        RECT 1258.270 1500.000 1258.550 1500.350 ;
        RECT 1255.900 17.690 1256.160 18.010 ;
        RECT 585.530 -4.800 586.090 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 91.610 19.620 91.930 19.680 ;
        RECT 430.170 19.620 430.490 19.680 ;
        RECT 91.610 19.480 430.490 19.620 ;
        RECT 91.610 19.420 91.930 19.480 ;
        RECT 430.170 19.420 430.490 19.480 ;
      LAYER via ;
        RECT 91.640 19.420 91.900 19.680 ;
        RECT 430.200 19.420 430.460 19.680 ;
      LAYER met2 ;
        RECT 450.510 1500.490 450.790 1504.000 ;
        RECT 448.660 1500.350 450.790 1500.490 ;
        RECT 448.660 20.245 448.800 1500.350 ;
        RECT 450.510 1500.000 450.790 1500.350 ;
        RECT 430.190 19.875 430.470 20.245 ;
        RECT 448.590 19.875 448.870 20.245 ;
        RECT 430.260 19.710 430.400 19.875 ;
        RECT 91.640 19.390 91.900 19.710 ;
        RECT 430.200 19.390 430.460 19.710 ;
        RECT 91.700 2.400 91.840 19.390 ;
        RECT 91.490 -4.800 92.050 2.400 ;
      LAYER via2 ;
        RECT 430.190 19.920 430.470 20.200 ;
        RECT 448.590 19.920 448.870 20.200 ;
      LAYER met3 ;
        RECT 430.165 20.210 430.495 20.225 ;
        RECT 448.565 20.210 448.895 20.225 ;
        RECT 430.165 19.910 448.895 20.210 ;
        RECT 430.165 19.895 430.495 19.910 ;
        RECT 448.565 19.895 448.895 19.910 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 603.130 18.260 603.450 18.320 ;
        RECT 606.810 18.260 607.130 18.320 ;
        RECT 603.130 18.120 607.130 18.260 ;
        RECT 603.130 18.060 603.450 18.120 ;
        RECT 606.810 18.060 607.130 18.120 ;
      LAYER via ;
        RECT 603.160 18.060 603.420 18.320 ;
        RECT 606.840 18.060 607.100 18.320 ;
      LAYER met2 ;
        RECT 1287.710 1500.420 1287.990 1504.000 ;
        RECT 1287.700 1500.000 1287.990 1500.420 ;
        RECT 1287.700 1487.685 1287.840 1500.000 ;
        RECT 606.830 1487.315 607.110 1487.685 ;
        RECT 1287.630 1487.315 1287.910 1487.685 ;
        RECT 606.900 18.350 607.040 1487.315 ;
        RECT 603.160 18.030 603.420 18.350 ;
        RECT 606.840 18.030 607.100 18.350 ;
        RECT 603.220 2.400 603.360 18.030 ;
        RECT 603.010 -4.800 603.570 2.400 ;
      LAYER via2 ;
        RECT 606.830 1487.360 607.110 1487.640 ;
        RECT 1287.630 1487.360 1287.910 1487.640 ;
      LAYER met3 ;
        RECT 606.805 1487.650 607.135 1487.665 ;
        RECT 1287.605 1487.650 1287.935 1487.665 ;
        RECT 606.805 1487.350 1287.935 1487.650 ;
        RECT 606.805 1487.335 607.135 1487.350 ;
        RECT 1287.605 1487.335 1287.935 1487.350 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 621.070 17.580 621.390 17.640 ;
        RECT 1311.070 17.580 1311.390 17.640 ;
        RECT 621.070 17.440 1311.390 17.580 ;
        RECT 621.070 17.380 621.390 17.440 ;
        RECT 1311.070 17.380 1311.390 17.440 ;
      LAYER via ;
        RECT 621.100 17.380 621.360 17.640 ;
        RECT 1311.100 17.380 1311.360 17.640 ;
      LAYER met2 ;
        RECT 1316.690 1500.490 1316.970 1504.000 ;
        RECT 1311.160 1500.350 1316.970 1500.490 ;
        RECT 1311.160 17.670 1311.300 1500.350 ;
        RECT 1316.690 1500.000 1316.970 1500.350 ;
        RECT 621.100 17.350 621.360 17.670 ;
        RECT 1311.100 17.350 1311.360 17.670 ;
        RECT 621.160 2.400 621.300 17.350 ;
        RECT 620.950 -4.800 621.510 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 477.550 19.280 477.870 19.340 ;
        RECT 131.260 19.140 477.870 19.280 ;
        RECT 115.530 18.940 115.850 19.000 ;
        RECT 131.260 18.940 131.400 19.140 ;
        RECT 477.550 19.080 477.870 19.140 ;
        RECT 115.530 18.800 131.400 18.940 ;
        RECT 115.530 18.740 115.850 18.800 ;
      LAYER via ;
        RECT 115.560 18.740 115.820 19.000 ;
        RECT 477.580 19.080 477.840 19.340 ;
      LAYER met2 ;
        RECT 489.610 1500.490 489.890 1504.000 ;
        RECT 483.160 1500.350 489.890 1500.490 ;
        RECT 483.160 19.565 483.300 1500.350 ;
        RECT 489.610 1500.000 489.890 1500.350 ;
        RECT 477.570 19.195 477.850 19.565 ;
        RECT 483.090 19.195 483.370 19.565 ;
        RECT 477.580 19.050 477.840 19.195 ;
        RECT 115.560 18.710 115.820 19.030 ;
        RECT 115.620 2.400 115.760 18.710 ;
        RECT 115.410 -4.800 115.970 2.400 ;
      LAYER via2 ;
        RECT 477.570 19.240 477.850 19.520 ;
        RECT 483.090 19.240 483.370 19.520 ;
      LAYER met3 ;
        RECT 477.545 19.530 477.875 19.545 ;
        RECT 483.065 19.530 483.395 19.545 ;
        RECT 477.545 19.230 483.395 19.530 ;
        RECT 477.545 19.215 477.875 19.230 ;
        RECT 483.065 19.215 483.395 19.230 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 478.100 19.140 483.300 19.280 ;
        RECT 139.450 18.940 139.770 19.000 ;
        RECT 478.100 18.940 478.240 19.140 ;
        RECT 139.450 18.800 478.240 18.940 ;
        RECT 483.160 18.940 483.300 19.140 ;
        RECT 513.430 18.940 513.750 19.000 ;
        RECT 483.160 18.800 513.750 18.940 ;
        RECT 139.450 18.740 139.770 18.800 ;
        RECT 513.430 18.740 513.750 18.800 ;
      LAYER via ;
        RECT 139.480 18.740 139.740 19.000 ;
        RECT 513.460 18.740 513.720 19.000 ;
      LAYER met2 ;
        RECT 528.250 1500.490 528.530 1504.000 ;
        RECT 524.560 1500.350 528.530 1500.490 ;
        RECT 524.560 19.565 524.700 1500.350 ;
        RECT 528.250 1500.000 528.530 1500.350 ;
        RECT 513.450 19.195 513.730 19.565 ;
        RECT 524.490 19.195 524.770 19.565 ;
        RECT 513.520 19.030 513.660 19.195 ;
        RECT 139.480 18.710 139.740 19.030 ;
        RECT 513.460 18.710 513.720 19.030 ;
        RECT 139.540 2.400 139.680 18.710 ;
        RECT 139.330 -4.800 139.890 2.400 ;
      LAYER via2 ;
        RECT 513.450 19.240 513.730 19.520 ;
        RECT 524.490 19.240 524.770 19.520 ;
      LAYER met3 ;
        RECT 513.425 19.530 513.755 19.545 ;
        RECT 524.465 19.530 524.795 19.545 ;
        RECT 513.425 19.230 524.795 19.530 ;
        RECT 513.425 19.215 513.755 19.230 ;
        RECT 524.465 19.215 524.795 19.230 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 157.390 18.600 157.710 18.660 ;
        RECT 552.070 18.600 552.390 18.660 ;
        RECT 157.390 18.460 552.390 18.600 ;
        RECT 157.390 18.400 157.710 18.460 ;
        RECT 552.070 18.400 552.390 18.460 ;
      LAYER via ;
        RECT 157.420 18.400 157.680 18.660 ;
        RECT 552.100 18.400 552.360 18.660 ;
      LAYER met2 ;
        RECT 557.690 1500.490 557.970 1504.000 ;
        RECT 552.160 1500.350 557.970 1500.490 ;
        RECT 552.160 18.690 552.300 1500.350 ;
        RECT 557.690 1500.000 557.970 1500.350 ;
        RECT 157.420 18.370 157.680 18.690 ;
        RECT 552.100 18.370 552.360 18.690 ;
        RECT 157.480 2.400 157.620 18.370 ;
        RECT 157.270 -4.800 157.830 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 174.870 18.260 175.190 18.320 ;
        RECT 549.310 18.260 549.630 18.320 ;
        RECT 174.870 18.120 549.630 18.260 ;
        RECT 174.870 18.060 175.190 18.120 ;
        RECT 549.310 18.060 549.630 18.120 ;
      LAYER via ;
        RECT 174.900 18.060 175.160 18.320 ;
        RECT 549.340 18.060 549.600 18.320 ;
      LAYER met2 ;
        RECT 586.670 1500.420 586.950 1504.000 ;
        RECT 586.660 1500.000 586.950 1500.420 ;
        RECT 586.660 19.565 586.800 1500.000 ;
        RECT 549.330 19.195 549.610 19.565 ;
        RECT 586.590 19.195 586.870 19.565 ;
        RECT 549.400 18.350 549.540 19.195 ;
        RECT 174.900 18.030 175.160 18.350 ;
        RECT 549.340 18.030 549.600 18.350 ;
        RECT 174.960 2.400 175.100 18.030 ;
        RECT 174.750 -4.800 175.310 2.400 ;
      LAYER via2 ;
        RECT 549.330 19.240 549.610 19.520 ;
        RECT 586.590 19.240 586.870 19.520 ;
      LAYER met3 ;
        RECT 549.305 19.530 549.635 19.545 ;
        RECT 586.565 19.530 586.895 19.545 ;
        RECT 549.305 19.230 586.895 19.530 ;
        RECT 549.305 19.215 549.635 19.230 ;
        RECT 586.565 19.215 586.895 19.230 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 227.310 17.240 227.630 17.300 ;
        RECT 234.210 17.240 234.530 17.300 ;
        RECT 227.310 17.100 234.530 17.240 ;
        RECT 227.310 17.040 227.630 17.100 ;
        RECT 234.210 17.040 234.530 17.100 ;
        RECT 420.510 17.240 420.830 17.300 ;
        RECT 469.270 17.240 469.590 17.300 ;
        RECT 420.510 17.100 469.590 17.240 ;
        RECT 420.510 17.040 420.830 17.100 ;
        RECT 469.270 17.040 469.590 17.100 ;
        RECT 496.870 17.240 497.190 17.300 ;
        RECT 614.630 17.240 614.950 17.300 ;
        RECT 496.870 17.100 614.950 17.240 ;
        RECT 496.870 17.040 497.190 17.100 ;
        RECT 614.630 17.040 614.950 17.100 ;
        RECT 343.230 16.560 343.550 16.620 ;
        RECT 320.320 16.420 343.550 16.560 ;
        RECT 234.210 16.220 234.530 16.280 ;
        RECT 320.320 16.220 320.460 16.420 ;
        RECT 343.230 16.360 343.550 16.420 ;
        RECT 234.210 16.080 320.460 16.220 ;
        RECT 234.210 16.020 234.530 16.080 ;
        RECT 192.810 14.520 193.130 14.580 ;
        RECT 227.310 14.520 227.630 14.580 ;
        RECT 192.810 14.380 227.630 14.520 ;
        RECT 192.810 14.320 193.130 14.380 ;
        RECT 227.310 14.320 227.630 14.380 ;
      LAYER via ;
        RECT 227.340 17.040 227.600 17.300 ;
        RECT 234.240 17.040 234.500 17.300 ;
        RECT 420.540 17.040 420.800 17.300 ;
        RECT 469.300 17.040 469.560 17.300 ;
        RECT 496.900 17.040 497.160 17.300 ;
        RECT 614.660 17.040 614.920 17.300 ;
        RECT 234.240 16.020 234.500 16.280 ;
        RECT 343.260 16.360 343.520 16.620 ;
        RECT 192.840 14.320 193.100 14.580 ;
        RECT 227.340 14.320 227.600 14.580 ;
      LAYER met2 ;
        RECT 616.110 1500.490 616.390 1504.000 ;
        RECT 614.720 1500.350 616.390 1500.490 ;
        RECT 227.340 17.010 227.600 17.330 ;
        RECT 234.240 17.010 234.500 17.330 ;
        RECT 343.250 17.155 343.530 17.525 ;
        RECT 420.530 17.155 420.810 17.525 ;
        RECT 614.720 17.330 614.860 1500.350 ;
        RECT 616.110 1500.000 616.390 1500.350 ;
        RECT 227.400 14.610 227.540 17.010 ;
        RECT 234.300 16.310 234.440 17.010 ;
        RECT 343.320 16.650 343.460 17.155 ;
        RECT 420.540 17.010 420.800 17.155 ;
        RECT 469.300 17.010 469.560 17.330 ;
        RECT 496.900 17.010 497.160 17.330 ;
        RECT 614.660 17.010 614.920 17.330 ;
        RECT 469.360 16.845 469.500 17.010 ;
        RECT 496.960 16.845 497.100 17.010 ;
        RECT 343.260 16.330 343.520 16.650 ;
        RECT 469.290 16.475 469.570 16.845 ;
        RECT 496.890 16.475 497.170 16.845 ;
        RECT 234.240 15.990 234.500 16.310 ;
        RECT 192.840 14.290 193.100 14.610 ;
        RECT 227.340 14.290 227.600 14.610 ;
        RECT 192.900 2.400 193.040 14.290 ;
        RECT 192.690 -4.800 193.250 2.400 ;
      LAYER via2 ;
        RECT 343.250 17.200 343.530 17.480 ;
        RECT 420.530 17.200 420.810 17.480 ;
        RECT 469.290 16.520 469.570 16.800 ;
        RECT 496.890 16.520 497.170 16.800 ;
      LAYER met3 ;
        RECT 343.225 17.490 343.555 17.505 ;
        RECT 420.505 17.490 420.835 17.505 ;
        RECT 343.225 17.190 420.835 17.490 ;
        RECT 343.225 17.175 343.555 17.190 ;
        RECT 420.505 17.175 420.835 17.190 ;
        RECT 469.265 16.810 469.595 16.825 ;
        RECT 496.865 16.810 497.195 16.825 ;
        RECT 469.265 16.510 497.195 16.810 ;
        RECT 469.265 16.495 469.595 16.510 ;
        RECT 496.865 16.495 497.195 16.510 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 213.510 1488.760 213.830 1488.820 ;
        RECT 644.990 1488.760 645.310 1488.820 ;
        RECT 213.510 1488.620 645.310 1488.760 ;
        RECT 213.510 1488.560 213.830 1488.620 ;
        RECT 644.990 1488.560 645.310 1488.620 ;
        RECT 210.750 17.580 211.070 17.640 ;
        RECT 213.510 17.580 213.830 17.640 ;
        RECT 210.750 17.440 213.830 17.580 ;
        RECT 210.750 17.380 211.070 17.440 ;
        RECT 213.510 17.380 213.830 17.440 ;
      LAYER via ;
        RECT 213.540 1488.560 213.800 1488.820 ;
        RECT 645.020 1488.560 645.280 1488.820 ;
        RECT 210.780 17.380 211.040 17.640 ;
        RECT 213.540 17.380 213.800 17.640 ;
      LAYER met2 ;
        RECT 645.090 1500.420 645.370 1504.000 ;
        RECT 645.080 1500.000 645.370 1500.420 ;
        RECT 645.080 1488.850 645.220 1500.000 ;
        RECT 213.540 1488.530 213.800 1488.850 ;
        RECT 645.020 1488.530 645.280 1488.850 ;
        RECT 213.600 17.670 213.740 1488.530 ;
        RECT 210.780 17.350 211.040 17.670 ;
        RECT 213.540 17.350 213.800 17.670 ;
        RECT 210.840 2.400 210.980 17.350 ;
        RECT 210.630 -4.800 211.190 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 228.690 14.520 229.010 14.580 ;
        RECT 669.830 14.520 670.150 14.580 ;
        RECT 228.690 14.380 670.150 14.520 ;
        RECT 228.690 14.320 229.010 14.380 ;
        RECT 669.830 14.320 670.150 14.380 ;
      LAYER via ;
        RECT 228.720 14.320 228.980 14.580 ;
        RECT 669.860 14.320 670.120 14.580 ;
      LAYER met2 ;
        RECT 674.530 1500.490 674.810 1504.000 ;
        RECT 669.920 1500.350 674.810 1500.490 ;
        RECT 669.920 14.610 670.060 1500.350 ;
        RECT 674.530 1500.000 674.810 1500.350 ;
        RECT 228.720 14.290 228.980 14.610 ;
        RECT 669.860 14.290 670.120 14.610 ;
        RECT 228.780 2.400 228.920 14.290 ;
        RECT 228.570 -4.800 229.130 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 54.810 1489.440 55.130 1489.500 ;
        RECT 382.330 1489.440 382.650 1489.500 ;
        RECT 54.810 1489.300 382.650 1489.440 ;
        RECT 54.810 1489.240 55.130 1489.300 ;
        RECT 382.330 1489.240 382.650 1489.300 ;
        RECT 50.210 17.580 50.530 17.640 ;
        RECT 54.810 17.580 55.130 17.640 ;
        RECT 50.210 17.440 55.130 17.580 ;
        RECT 50.210 17.380 50.530 17.440 ;
        RECT 54.810 17.380 55.130 17.440 ;
      LAYER via ;
        RECT 54.840 1489.240 55.100 1489.500 ;
        RECT 382.360 1489.240 382.620 1489.500 ;
        RECT 50.240 17.380 50.500 17.640 ;
        RECT 54.840 17.380 55.100 17.640 ;
      LAYER met2 ;
        RECT 382.430 1500.420 382.710 1504.000 ;
        RECT 382.420 1500.000 382.710 1500.420 ;
        RECT 382.420 1489.530 382.560 1500.000 ;
        RECT 54.840 1489.210 55.100 1489.530 ;
        RECT 382.360 1489.210 382.620 1489.530 ;
        RECT 54.900 17.670 55.040 1489.210 ;
        RECT 50.240 17.350 50.500 17.670 ;
        RECT 54.840 17.350 55.100 17.670 ;
        RECT 50.300 2.400 50.440 17.350 ;
        RECT 50.090 -4.800 50.650 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 254.910 1484.680 255.230 1484.740 ;
        RECT 713.070 1484.680 713.390 1484.740 ;
        RECT 254.910 1484.540 713.390 1484.680 ;
        RECT 254.910 1484.480 255.230 1484.540 ;
        RECT 713.070 1484.480 713.390 1484.540 ;
        RECT 252.610 17.240 252.930 17.300 ;
        RECT 254.910 17.240 255.230 17.300 ;
        RECT 252.610 17.100 255.230 17.240 ;
        RECT 252.610 17.040 252.930 17.100 ;
        RECT 254.910 17.040 255.230 17.100 ;
      LAYER via ;
        RECT 254.940 1484.480 255.200 1484.740 ;
        RECT 713.100 1484.480 713.360 1484.740 ;
        RECT 252.640 17.040 252.900 17.300 ;
        RECT 254.940 17.040 255.200 17.300 ;
      LAYER met2 ;
        RECT 713.170 1500.420 713.450 1504.000 ;
        RECT 713.160 1500.000 713.450 1500.420 ;
        RECT 713.160 1484.770 713.300 1500.000 ;
        RECT 254.940 1484.450 255.200 1484.770 ;
        RECT 713.100 1484.450 713.360 1484.770 ;
        RECT 255.000 17.330 255.140 1484.450 ;
        RECT 252.640 17.010 252.900 17.330 ;
        RECT 254.940 17.010 255.200 17.330 ;
        RECT 252.700 2.400 252.840 17.010 ;
        RECT 252.490 -4.800 253.050 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 270.090 15.200 270.410 15.260 ;
        RECT 738.370 15.200 738.690 15.260 ;
        RECT 270.090 15.060 738.690 15.200 ;
        RECT 270.090 15.000 270.410 15.060 ;
        RECT 738.370 15.000 738.690 15.060 ;
      LAYER via ;
        RECT 270.120 15.000 270.380 15.260 ;
        RECT 738.400 15.000 738.660 15.260 ;
      LAYER met2 ;
        RECT 742.610 1500.490 742.890 1504.000 ;
        RECT 738.460 1500.350 742.890 1500.490 ;
        RECT 738.460 15.290 738.600 1500.350 ;
        RECT 742.610 1500.000 742.890 1500.350 ;
        RECT 270.120 14.970 270.380 15.290 ;
        RECT 738.400 14.970 738.660 15.290 ;
        RECT 270.180 2.400 270.320 14.970 ;
        RECT 269.970 -4.800 270.530 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 288.030 15.880 288.350 15.940 ;
        RECT 765.970 15.880 766.290 15.940 ;
        RECT 288.030 15.740 766.290 15.880 ;
        RECT 288.030 15.680 288.350 15.740 ;
        RECT 765.970 15.680 766.290 15.740 ;
      LAYER via ;
        RECT 288.060 15.680 288.320 15.940 ;
        RECT 766.000 15.680 766.260 15.940 ;
      LAYER met2 ;
        RECT 771.590 1500.490 771.870 1504.000 ;
        RECT 766.060 1500.350 771.870 1500.490 ;
        RECT 766.060 15.970 766.200 1500.350 ;
        RECT 771.590 1500.000 771.870 1500.350 ;
        RECT 288.060 15.650 288.320 15.970 ;
        RECT 766.000 15.650 766.260 15.970 ;
        RECT 288.120 2.400 288.260 15.650 ;
        RECT 287.910 -4.800 288.470 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 310.110 1485.020 310.430 1485.080 ;
        RECT 800.930 1485.020 801.250 1485.080 ;
        RECT 310.110 1484.880 801.250 1485.020 ;
        RECT 310.110 1484.820 310.430 1484.880 ;
        RECT 800.930 1484.820 801.250 1484.880 ;
        RECT 305.970 20.640 306.290 20.700 ;
        RECT 310.110 20.640 310.430 20.700 ;
        RECT 305.970 20.500 310.430 20.640 ;
        RECT 305.970 20.440 306.290 20.500 ;
        RECT 310.110 20.440 310.430 20.500 ;
      LAYER via ;
        RECT 310.140 1484.820 310.400 1485.080 ;
        RECT 800.960 1484.820 801.220 1485.080 ;
        RECT 306.000 20.440 306.260 20.700 ;
        RECT 310.140 20.440 310.400 20.700 ;
      LAYER met2 ;
        RECT 801.030 1500.420 801.310 1504.000 ;
        RECT 801.020 1500.000 801.310 1500.420 ;
        RECT 801.020 1485.110 801.160 1500.000 ;
        RECT 310.140 1484.790 310.400 1485.110 ;
        RECT 800.960 1484.790 801.220 1485.110 ;
        RECT 310.200 20.730 310.340 1484.790 ;
        RECT 306.000 20.410 306.260 20.730 ;
        RECT 310.140 20.410 310.400 20.730 ;
        RECT 306.060 2.400 306.200 20.410 ;
        RECT 305.850 -4.800 306.410 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 323.910 1485.360 324.230 1485.420 ;
        RECT 829.910 1485.360 830.230 1485.420 ;
        RECT 323.910 1485.220 830.230 1485.360 ;
        RECT 323.910 1485.160 324.230 1485.220 ;
        RECT 829.910 1485.160 830.230 1485.220 ;
      LAYER via ;
        RECT 323.940 1485.160 324.200 1485.420 ;
        RECT 829.940 1485.160 830.200 1485.420 ;
      LAYER met2 ;
        RECT 830.010 1500.420 830.290 1504.000 ;
        RECT 830.000 1500.000 830.290 1500.420 ;
        RECT 830.000 1485.450 830.140 1500.000 ;
        RECT 323.940 1485.130 324.200 1485.450 ;
        RECT 829.940 1485.130 830.200 1485.450 ;
        RECT 324.000 2.400 324.140 1485.130 ;
        RECT 323.790 -4.800 324.350 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 341.390 20.640 341.710 20.700 ;
        RECT 366.690 20.640 367.010 20.700 ;
        RECT 341.390 20.500 367.010 20.640 ;
        RECT 341.390 20.440 341.710 20.500 ;
        RECT 366.690 20.440 367.010 20.500 ;
        RECT 366.690 16.560 367.010 16.620 ;
        RECT 855.670 16.560 855.990 16.620 ;
        RECT 366.690 16.420 855.990 16.560 ;
        RECT 366.690 16.360 367.010 16.420 ;
        RECT 855.670 16.360 855.990 16.420 ;
      LAYER via ;
        RECT 341.420 20.440 341.680 20.700 ;
        RECT 366.720 20.440 366.980 20.700 ;
        RECT 366.720 16.360 366.980 16.620 ;
        RECT 855.700 16.360 855.960 16.620 ;
      LAYER met2 ;
        RECT 859.450 1500.490 859.730 1504.000 ;
        RECT 855.760 1500.350 859.730 1500.490 ;
        RECT 341.420 20.410 341.680 20.730 ;
        RECT 366.720 20.410 366.980 20.730 ;
        RECT 341.480 2.400 341.620 20.410 ;
        RECT 366.780 16.650 366.920 20.410 ;
        RECT 855.760 16.650 855.900 1500.350 ;
        RECT 859.450 1500.000 859.730 1500.350 ;
        RECT 366.720 16.330 366.980 16.650 ;
        RECT 855.700 16.330 855.960 16.650 ;
        RECT 341.270 -4.800 341.830 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 364.850 1486.040 365.170 1486.100 ;
        RECT 888.330 1486.040 888.650 1486.100 ;
        RECT 364.850 1485.900 888.650 1486.040 ;
        RECT 364.850 1485.840 365.170 1485.900 ;
        RECT 888.330 1485.840 888.650 1485.900 ;
        RECT 359.330 17.240 359.650 17.300 ;
        RECT 364.850 17.240 365.170 17.300 ;
        RECT 359.330 17.100 365.170 17.240 ;
        RECT 359.330 17.040 359.650 17.100 ;
        RECT 364.850 17.040 365.170 17.100 ;
      LAYER via ;
        RECT 364.880 1485.840 365.140 1486.100 ;
        RECT 888.360 1485.840 888.620 1486.100 ;
        RECT 359.360 17.040 359.620 17.300 ;
        RECT 364.880 17.040 365.140 17.300 ;
      LAYER met2 ;
        RECT 888.430 1500.420 888.710 1504.000 ;
        RECT 888.420 1500.000 888.710 1500.420 ;
        RECT 888.420 1486.130 888.560 1500.000 ;
        RECT 364.880 1485.810 365.140 1486.130 ;
        RECT 888.360 1485.810 888.620 1486.130 ;
        RECT 364.940 17.330 365.080 1485.810 ;
        RECT 359.360 17.010 359.620 17.330 ;
        RECT 364.880 17.010 365.140 17.330 ;
        RECT 359.420 2.400 359.560 17.010 ;
        RECT 359.210 -4.800 359.770 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 414.990 20.640 415.310 20.700 ;
        RECT 917.770 20.640 918.090 20.700 ;
        RECT 414.990 20.500 918.090 20.640 ;
        RECT 414.990 20.440 415.310 20.500 ;
        RECT 917.770 20.440 918.090 20.500 ;
        RECT 377.270 19.960 377.590 20.020 ;
        RECT 394.750 19.960 395.070 20.020 ;
        RECT 377.270 19.820 395.070 19.960 ;
        RECT 377.270 19.760 377.590 19.820 ;
        RECT 394.750 19.760 395.070 19.820 ;
      LAYER via ;
        RECT 415.020 20.440 415.280 20.700 ;
        RECT 917.800 20.440 918.060 20.700 ;
        RECT 377.300 19.760 377.560 20.020 ;
        RECT 394.780 19.760 395.040 20.020 ;
      LAYER met2 ;
        RECT 917.870 1500.420 918.150 1504.000 ;
        RECT 917.860 1500.000 918.150 1500.420 ;
        RECT 917.860 20.730 918.000 1500.000 ;
        RECT 415.020 20.410 415.280 20.730 ;
        RECT 917.800 20.410 918.060 20.730 ;
        RECT 415.080 20.245 415.220 20.410 ;
        RECT 377.300 19.730 377.560 20.050 ;
        RECT 394.770 19.875 395.050 20.245 ;
        RECT 415.010 19.875 415.290 20.245 ;
        RECT 394.780 19.730 395.040 19.875 ;
        RECT 377.360 2.400 377.500 19.730 ;
        RECT 377.150 -4.800 377.710 2.400 ;
      LAYER via2 ;
        RECT 394.770 19.920 395.050 20.200 ;
        RECT 415.010 19.920 415.290 20.200 ;
      LAYER met3 ;
        RECT 394.745 20.210 395.075 20.225 ;
        RECT 414.985 20.210 415.315 20.225 ;
        RECT 394.745 19.910 415.315 20.210 ;
        RECT 394.745 19.895 395.075 19.910 ;
        RECT 414.985 19.895 415.315 19.910 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 399.810 1486.720 400.130 1486.780 ;
        RECT 946.750 1486.720 947.070 1486.780 ;
        RECT 399.810 1486.580 947.070 1486.720 ;
        RECT 399.810 1486.520 400.130 1486.580 ;
        RECT 946.750 1486.520 947.070 1486.580 ;
        RECT 395.210 19.960 395.530 20.020 ;
        RECT 399.810 19.960 400.130 20.020 ;
        RECT 395.210 19.820 400.130 19.960 ;
        RECT 395.210 19.760 395.530 19.820 ;
        RECT 399.810 19.760 400.130 19.820 ;
      LAYER via ;
        RECT 399.840 1486.520 400.100 1486.780 ;
        RECT 946.780 1486.520 947.040 1486.780 ;
        RECT 395.240 19.760 395.500 20.020 ;
        RECT 399.840 19.760 400.100 20.020 ;
      LAYER met2 ;
        RECT 946.850 1500.420 947.130 1504.000 ;
        RECT 946.840 1500.000 947.130 1500.420 ;
        RECT 946.840 1486.810 946.980 1500.000 ;
        RECT 399.840 1486.490 400.100 1486.810 ;
        RECT 946.780 1486.490 947.040 1486.810 ;
        RECT 399.900 20.050 400.040 1486.490 ;
        RECT 395.240 19.730 395.500 20.050 ;
        RECT 399.840 19.730 400.100 20.050 ;
        RECT 395.300 2.400 395.440 19.730 ;
        RECT 395.090 -4.800 395.650 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 413.150 20.300 413.470 20.360 ;
        RECT 413.150 20.160 414.300 20.300 ;
        RECT 413.150 20.100 413.470 20.160 ;
        RECT 414.160 19.960 414.300 20.160 ;
        RECT 972.970 19.960 973.290 20.020 ;
        RECT 414.160 19.820 973.290 19.960 ;
        RECT 972.970 19.760 973.290 19.820 ;
      LAYER via ;
        RECT 413.180 20.100 413.440 20.360 ;
        RECT 973.000 19.760 973.260 20.020 ;
      LAYER met2 ;
        RECT 975.830 1500.490 976.110 1504.000 ;
        RECT 973.060 1500.350 976.110 1500.490 ;
        RECT 413.180 20.070 413.440 20.390 ;
        RECT 413.240 2.400 413.380 20.070 ;
        RECT 973.060 20.050 973.200 1500.350 ;
        RECT 975.830 1500.000 976.110 1500.350 ;
        RECT 973.000 19.730 973.260 20.050 ;
        RECT 413.030 -4.800 413.590 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 75.510 1488.420 75.830 1488.480 ;
        RECT 420.970 1488.420 421.290 1488.480 ;
        RECT 75.510 1488.280 421.290 1488.420 ;
        RECT 75.510 1488.220 75.830 1488.280 ;
        RECT 420.970 1488.220 421.290 1488.280 ;
      LAYER via ;
        RECT 75.540 1488.220 75.800 1488.480 ;
        RECT 421.000 1488.220 421.260 1488.480 ;
      LAYER met2 ;
        RECT 421.070 1500.420 421.350 1504.000 ;
        RECT 421.060 1500.000 421.350 1500.420 ;
        RECT 421.060 1488.510 421.200 1500.000 ;
        RECT 75.540 1488.190 75.800 1488.510 ;
        RECT 421.000 1488.190 421.260 1488.510 ;
        RECT 75.600 17.410 75.740 1488.190 ;
        RECT 74.220 17.270 75.740 17.410 ;
        RECT 74.220 2.400 74.360 17.270 ;
        RECT 74.010 -4.800 74.570 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 434.310 1490.120 434.630 1490.180 ;
        RECT 1005.170 1490.120 1005.490 1490.180 ;
        RECT 434.310 1489.980 1005.490 1490.120 ;
        RECT 434.310 1489.920 434.630 1489.980 ;
        RECT 1005.170 1489.920 1005.490 1489.980 ;
        RECT 434.310 146.240 434.630 146.500 ;
        RECT 434.400 145.820 434.540 146.240 ;
        RECT 434.310 145.560 434.630 145.820 ;
        RECT 430.630 19.620 430.950 19.680 ;
        RECT 434.310 19.620 434.630 19.680 ;
        RECT 430.630 19.480 434.630 19.620 ;
        RECT 430.630 19.420 430.950 19.480 ;
        RECT 434.310 19.420 434.630 19.480 ;
      LAYER via ;
        RECT 434.340 1489.920 434.600 1490.180 ;
        RECT 1005.200 1489.920 1005.460 1490.180 ;
        RECT 434.340 146.240 434.600 146.500 ;
        RECT 434.340 145.560 434.600 145.820 ;
        RECT 430.660 19.420 430.920 19.680 ;
        RECT 434.340 19.420 434.600 19.680 ;
      LAYER met2 ;
        RECT 1005.270 1500.420 1005.550 1504.000 ;
        RECT 1005.260 1500.000 1005.550 1500.420 ;
        RECT 1005.260 1490.210 1005.400 1500.000 ;
        RECT 434.340 1489.890 434.600 1490.210 ;
        RECT 1005.200 1489.890 1005.460 1490.210 ;
        RECT 434.400 146.530 434.540 1489.890 ;
        RECT 434.340 146.210 434.600 146.530 ;
        RECT 434.340 145.530 434.600 145.850 ;
        RECT 434.400 19.710 434.540 145.530 ;
        RECT 430.660 19.390 430.920 19.710 ;
        RECT 434.340 19.390 434.600 19.710 ;
        RECT 430.720 2.400 430.860 19.390 ;
        RECT 430.510 -4.800 431.070 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 448.570 19.620 448.890 19.680 ;
        RECT 466.050 19.620 466.370 19.680 ;
        RECT 448.570 19.480 466.370 19.620 ;
        RECT 448.570 19.420 448.890 19.480 ;
        RECT 466.050 19.420 466.370 19.480 ;
        RECT 469.270 19.620 469.590 19.680 ;
        RECT 1028.170 19.620 1028.490 19.680 ;
        RECT 469.270 19.480 1028.490 19.620 ;
        RECT 469.270 19.420 469.590 19.480 ;
        RECT 1028.170 19.420 1028.490 19.480 ;
      LAYER via ;
        RECT 448.600 19.420 448.860 19.680 ;
        RECT 466.080 19.420 466.340 19.680 ;
        RECT 469.300 19.420 469.560 19.680 ;
        RECT 1028.200 19.420 1028.460 19.680 ;
      LAYER met2 ;
        RECT 1034.250 1500.490 1034.530 1504.000 ;
        RECT 1028.260 1500.350 1034.530 1500.490 ;
        RECT 1028.260 19.710 1028.400 1500.350 ;
        RECT 1034.250 1500.000 1034.530 1500.350 ;
        RECT 448.600 19.390 448.860 19.710 ;
        RECT 466.080 19.565 466.340 19.710 ;
        RECT 469.300 19.565 469.560 19.710 ;
        RECT 448.660 2.400 448.800 19.390 ;
        RECT 466.070 19.195 466.350 19.565 ;
        RECT 469.290 19.195 469.570 19.565 ;
        RECT 1028.200 19.390 1028.460 19.710 ;
        RECT 448.450 -4.800 449.010 2.400 ;
      LAYER via2 ;
        RECT 466.070 19.240 466.350 19.520 ;
        RECT 469.290 19.240 469.570 19.520 ;
      LAYER met3 ;
        RECT 466.045 19.530 466.375 19.545 ;
        RECT 469.265 19.530 469.595 19.545 ;
        RECT 466.045 19.230 469.595 19.530 ;
        RECT 466.045 19.215 466.375 19.230 ;
        RECT 469.265 19.215 469.595 19.230 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 468.810 1489.100 469.130 1489.160 ;
        RECT 1063.590 1489.100 1063.910 1489.160 ;
        RECT 468.810 1488.960 1063.910 1489.100 ;
        RECT 468.810 1488.900 469.130 1488.960 ;
        RECT 1063.590 1488.900 1063.910 1488.960 ;
        RECT 466.510 19.620 466.830 19.680 ;
        RECT 468.810 19.620 469.130 19.680 ;
        RECT 466.510 19.480 469.130 19.620 ;
        RECT 466.510 19.420 466.830 19.480 ;
        RECT 468.810 19.420 469.130 19.480 ;
      LAYER via ;
        RECT 468.840 1488.900 469.100 1489.160 ;
        RECT 1063.620 1488.900 1063.880 1489.160 ;
        RECT 466.540 19.420 466.800 19.680 ;
        RECT 468.840 19.420 469.100 19.680 ;
      LAYER met2 ;
        RECT 1063.690 1500.420 1063.970 1504.000 ;
        RECT 1063.680 1500.000 1063.970 1500.420 ;
        RECT 1063.680 1489.190 1063.820 1500.000 ;
        RECT 468.840 1488.870 469.100 1489.190 ;
        RECT 1063.620 1488.870 1063.880 1489.190 ;
        RECT 468.900 19.710 469.040 1488.870 ;
        RECT 466.540 19.390 466.800 19.710 ;
        RECT 468.840 19.390 469.100 19.710 ;
        RECT 466.600 2.400 466.740 19.390 ;
        RECT 466.390 -4.800 466.950 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 484.450 19.280 484.770 19.340 ;
        RECT 1090.270 19.280 1090.590 19.340 ;
        RECT 484.450 19.140 1090.590 19.280 ;
        RECT 484.450 19.080 484.770 19.140 ;
        RECT 1090.270 19.080 1090.590 19.140 ;
      LAYER via ;
        RECT 484.480 19.080 484.740 19.340 ;
        RECT 1090.300 19.080 1090.560 19.340 ;
      LAYER met2 ;
        RECT 1092.670 1500.490 1092.950 1504.000 ;
        RECT 1090.360 1500.350 1092.950 1500.490 ;
        RECT 1090.360 19.370 1090.500 1500.350 ;
        RECT 1092.670 1500.000 1092.950 1500.350 ;
        RECT 484.480 19.050 484.740 19.370 ;
        RECT 1090.300 19.050 1090.560 19.370 ;
        RECT 484.540 2.400 484.680 19.050 ;
        RECT 484.330 -4.800 484.890 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 503.310 1488.420 503.630 1488.480 ;
        RECT 1122.010 1488.420 1122.330 1488.480 ;
        RECT 503.310 1488.280 1122.330 1488.420 ;
        RECT 503.310 1488.220 503.630 1488.280 ;
        RECT 1122.010 1488.220 1122.330 1488.280 ;
      LAYER via ;
        RECT 503.340 1488.220 503.600 1488.480 ;
        RECT 1122.040 1488.220 1122.300 1488.480 ;
      LAYER met2 ;
        RECT 1122.110 1500.420 1122.390 1504.000 ;
        RECT 1122.100 1500.000 1122.390 1500.420 ;
        RECT 1122.100 1488.510 1122.240 1500.000 ;
        RECT 503.340 1488.190 503.600 1488.510 ;
        RECT 1122.040 1488.190 1122.300 1488.510 ;
        RECT 503.400 3.130 503.540 1488.190 ;
        RECT 502.480 2.990 503.540 3.130 ;
        RECT 502.480 2.400 502.620 2.990 ;
        RECT 502.270 -4.800 502.830 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1151.090 1500.490 1151.370 1504.000 ;
        RECT 1145.560 1500.350 1151.370 1500.490 ;
        RECT 1145.560 16.845 1145.700 1500.350 ;
        RECT 1151.090 1500.000 1151.370 1500.350 ;
        RECT 519.890 16.475 520.170 16.845 ;
        RECT 1145.490 16.475 1145.770 16.845 ;
        RECT 519.960 2.400 520.100 16.475 ;
        RECT 519.750 -4.800 520.310 2.400 ;
      LAYER via2 ;
        RECT 519.890 16.520 520.170 16.800 ;
        RECT 1145.490 16.520 1145.770 16.800 ;
      LAYER met3 ;
        RECT 519.865 16.810 520.195 16.825 ;
        RECT 1145.465 16.810 1145.795 16.825 ;
        RECT 519.865 16.510 1145.795 16.810 ;
        RECT 519.865 16.495 520.195 16.510 ;
        RECT 1145.465 16.495 1145.795 16.510 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 537.350 1487.400 537.670 1487.460 ;
        RECT 1180.430 1487.400 1180.750 1487.460 ;
        RECT 537.350 1487.260 1180.750 1487.400 ;
        RECT 537.350 1487.200 537.670 1487.260 ;
        RECT 1180.430 1487.200 1180.750 1487.260 ;
      LAYER via ;
        RECT 537.380 1487.200 537.640 1487.460 ;
        RECT 1180.460 1487.200 1180.720 1487.460 ;
      LAYER met2 ;
        RECT 1180.530 1500.420 1180.810 1504.000 ;
        RECT 1180.520 1500.000 1180.810 1500.420 ;
        RECT 1180.520 1487.490 1180.660 1500.000 ;
        RECT 537.380 1487.170 537.640 1487.490 ;
        RECT 1180.460 1487.170 1180.720 1487.490 ;
        RECT 537.440 18.090 537.580 1487.170 ;
        RECT 537.440 17.950 538.040 18.090 ;
        RECT 537.900 2.400 538.040 17.950 ;
        RECT 537.690 -4.800 538.250 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1207.570 18.600 1207.890 18.660 ;
        RECT 580.680 18.460 1207.890 18.600 ;
        RECT 555.750 17.920 556.070 17.980 ;
        RECT 580.680 17.920 580.820 18.460 ;
        RECT 1207.570 18.400 1207.890 18.460 ;
        RECT 555.750 17.780 580.820 17.920 ;
        RECT 555.750 17.720 556.070 17.780 ;
      LAYER via ;
        RECT 555.780 17.720 556.040 17.980 ;
        RECT 1207.600 18.400 1207.860 18.660 ;
      LAYER met2 ;
        RECT 1209.510 1500.490 1209.790 1504.000 ;
        RECT 1207.660 1500.350 1209.790 1500.490 ;
        RECT 1207.660 18.690 1207.800 1500.350 ;
        RECT 1209.510 1500.000 1209.790 1500.350 ;
        RECT 1207.600 18.370 1207.860 18.690 ;
        RECT 555.780 17.690 556.040 18.010 ;
        RECT 555.840 2.400 555.980 17.690 ;
        RECT 555.630 -4.800 556.190 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 573.690 18.940 574.010 19.000 ;
        RECT 579.210 18.940 579.530 19.000 ;
        RECT 573.690 18.800 579.530 18.940 ;
        RECT 573.690 18.740 574.010 18.800 ;
        RECT 579.210 18.740 579.530 18.800 ;
      LAYER via ;
        RECT 573.720 18.740 573.980 19.000 ;
        RECT 579.240 18.740 579.500 19.000 ;
      LAYER met2 ;
        RECT 1238.950 1500.420 1239.230 1504.000 ;
        RECT 1238.940 1500.000 1239.230 1500.420 ;
        RECT 1238.940 1488.365 1239.080 1500.000 ;
        RECT 579.230 1487.995 579.510 1488.365 ;
        RECT 1238.870 1487.995 1239.150 1488.365 ;
        RECT 579.300 19.030 579.440 1487.995 ;
        RECT 573.720 18.710 573.980 19.030 ;
        RECT 579.240 18.710 579.500 19.030 ;
        RECT 573.780 2.400 573.920 18.710 ;
        RECT 573.570 -4.800 574.130 2.400 ;
      LAYER via2 ;
        RECT 579.230 1488.040 579.510 1488.320 ;
        RECT 1238.870 1488.040 1239.150 1488.320 ;
      LAYER met3 ;
        RECT 579.205 1488.330 579.535 1488.345 ;
        RECT 1238.845 1488.330 1239.175 1488.345 ;
        RECT 579.205 1488.030 1239.175 1488.330 ;
        RECT 579.205 1488.015 579.535 1488.030 ;
        RECT 1238.845 1488.015 1239.175 1488.030 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 614.170 18.260 614.490 18.320 ;
        RECT 1262.770 18.260 1263.090 18.320 ;
        RECT 614.170 18.120 1263.090 18.260 ;
        RECT 614.170 18.060 614.490 18.120 ;
        RECT 1262.770 18.060 1263.090 18.120 ;
        RECT 591.170 17.920 591.490 17.980 ;
        RECT 591.170 17.780 602.440 17.920 ;
        RECT 591.170 17.720 591.490 17.780 ;
        RECT 602.300 17.580 602.440 17.780 ;
        RECT 613.250 17.580 613.570 17.640 ;
        RECT 602.300 17.440 613.570 17.580 ;
        RECT 613.250 17.380 613.570 17.440 ;
      LAYER via ;
        RECT 614.200 18.060 614.460 18.320 ;
        RECT 1262.800 18.060 1263.060 18.320 ;
        RECT 591.200 17.720 591.460 17.980 ;
        RECT 613.280 17.380 613.540 17.640 ;
      LAYER met2 ;
        RECT 1267.930 1500.490 1268.210 1504.000 ;
        RECT 1262.860 1500.350 1268.210 1500.490 ;
        RECT 1262.860 18.350 1263.000 1500.350 ;
        RECT 1267.930 1500.000 1268.210 1500.350 ;
        RECT 614.200 18.030 614.460 18.350 ;
        RECT 1262.800 18.030 1263.060 18.350 ;
        RECT 591.200 17.690 591.460 18.010 ;
        RECT 591.260 2.400 591.400 17.690 ;
        RECT 613.280 17.410 613.540 17.670 ;
        RECT 614.260 17.410 614.400 18.030 ;
        RECT 613.280 17.350 614.400 17.410 ;
        RECT 613.340 17.270 614.400 17.350 ;
        RECT 591.050 -4.800 591.610 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 103.110 1488.080 103.430 1488.140 ;
        RECT 460.070 1488.080 460.390 1488.140 ;
        RECT 103.110 1487.940 460.390 1488.080 ;
        RECT 103.110 1487.880 103.430 1487.940 ;
        RECT 460.070 1487.880 460.390 1487.940 ;
        RECT 97.590 17.580 97.910 17.640 ;
        RECT 103.110 17.580 103.430 17.640 ;
        RECT 97.590 17.440 103.430 17.580 ;
        RECT 97.590 17.380 97.910 17.440 ;
        RECT 103.110 17.380 103.430 17.440 ;
      LAYER via ;
        RECT 103.140 1487.880 103.400 1488.140 ;
        RECT 460.100 1487.880 460.360 1488.140 ;
        RECT 97.620 17.380 97.880 17.640 ;
        RECT 103.140 17.380 103.400 17.640 ;
      LAYER met2 ;
        RECT 460.170 1500.420 460.450 1504.000 ;
        RECT 460.160 1500.000 460.450 1500.420 ;
        RECT 460.160 1488.170 460.300 1500.000 ;
        RECT 103.140 1487.850 103.400 1488.170 ;
        RECT 460.100 1487.850 460.360 1488.170 ;
        RECT 103.200 17.670 103.340 1487.850 ;
        RECT 97.620 17.350 97.880 17.670 ;
        RECT 103.140 17.350 103.400 17.670 ;
        RECT 97.680 2.400 97.820 17.350 ;
        RECT 97.470 -4.800 98.030 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 609.110 18.260 609.430 18.320 ;
        RECT 613.710 18.260 614.030 18.320 ;
        RECT 609.110 18.120 614.030 18.260 ;
        RECT 609.110 18.060 609.430 18.120 ;
        RECT 613.710 18.060 614.030 18.120 ;
      LAYER via ;
        RECT 609.140 18.060 609.400 18.320 ;
        RECT 613.740 18.060 614.000 18.320 ;
      LAYER met2 ;
        RECT 1297.370 1500.420 1297.650 1504.000 ;
        RECT 1297.360 1500.000 1297.650 1500.420 ;
        RECT 1297.360 1487.005 1297.500 1500.000 ;
        RECT 613.730 1486.635 614.010 1487.005 ;
        RECT 1297.290 1486.635 1297.570 1487.005 ;
        RECT 613.800 18.350 613.940 1486.635 ;
        RECT 609.140 18.030 609.400 18.350 ;
        RECT 613.740 18.030 614.000 18.350 ;
        RECT 609.200 2.400 609.340 18.030 ;
        RECT 608.990 -4.800 609.550 2.400 ;
      LAYER via2 ;
        RECT 613.730 1486.680 614.010 1486.960 ;
        RECT 1297.290 1486.680 1297.570 1486.960 ;
      LAYER met3 ;
        RECT 613.705 1486.970 614.035 1486.985 ;
        RECT 1297.265 1486.970 1297.595 1486.985 ;
        RECT 613.705 1486.670 1297.595 1486.970 ;
        RECT 613.705 1486.655 614.035 1486.670 ;
        RECT 1297.265 1486.655 1297.595 1486.670 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 627.050 17.240 627.370 17.300 ;
        RECT 1324.870 17.240 1325.190 17.300 ;
        RECT 627.050 17.100 1325.190 17.240 ;
        RECT 627.050 17.040 627.370 17.100 ;
        RECT 1324.870 17.040 1325.190 17.100 ;
      LAYER via ;
        RECT 627.080 17.040 627.340 17.300 ;
        RECT 1324.900 17.040 1325.160 17.300 ;
      LAYER met2 ;
        RECT 1326.350 1500.490 1326.630 1504.000 ;
        RECT 1324.960 1500.350 1326.630 1500.490 ;
        RECT 1324.960 17.330 1325.100 1500.350 ;
        RECT 1326.350 1500.000 1326.630 1500.350 ;
        RECT 627.080 17.010 627.340 17.330 ;
        RECT 1324.900 17.010 1325.160 17.330 ;
        RECT 627.140 2.400 627.280 17.010 ;
        RECT 626.930 -4.800 627.490 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 123.810 1487.400 124.130 1487.460 ;
        RECT 499.170 1487.400 499.490 1487.460 ;
        RECT 123.810 1487.260 499.490 1487.400 ;
        RECT 123.810 1487.200 124.130 1487.260 ;
        RECT 499.170 1487.200 499.490 1487.260 ;
        RECT 121.510 19.280 121.830 19.340 ;
        RECT 123.810 19.280 124.130 19.340 ;
        RECT 121.510 19.140 124.130 19.280 ;
        RECT 121.510 19.080 121.830 19.140 ;
        RECT 123.810 19.080 124.130 19.140 ;
      LAYER via ;
        RECT 123.840 1487.200 124.100 1487.460 ;
        RECT 499.200 1487.200 499.460 1487.460 ;
        RECT 121.540 19.080 121.800 19.340 ;
        RECT 123.840 19.080 124.100 19.340 ;
      LAYER met2 ;
        RECT 499.270 1500.420 499.550 1504.000 ;
        RECT 499.260 1500.000 499.550 1500.420 ;
        RECT 499.260 1487.490 499.400 1500.000 ;
        RECT 123.840 1487.170 124.100 1487.490 ;
        RECT 499.200 1487.170 499.460 1487.490 ;
        RECT 123.900 19.370 124.040 1487.170 ;
        RECT 121.540 19.050 121.800 19.370 ;
        RECT 123.840 19.050 124.100 19.370 ;
        RECT 121.600 2.400 121.740 19.050 ;
        RECT 121.390 -4.800 121.950 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 210.290 1483.660 210.610 1483.720 ;
        RECT 536.430 1483.660 536.750 1483.720 ;
        RECT 210.290 1483.520 536.750 1483.660 ;
        RECT 210.290 1483.460 210.610 1483.520 ;
        RECT 536.430 1483.460 536.750 1483.520 ;
        RECT 145.430 15.540 145.750 15.600 ;
        RECT 145.430 15.400 179.700 15.540 ;
        RECT 145.430 15.340 145.750 15.400 ;
        RECT 179.560 14.860 179.700 15.400 ;
        RECT 210.290 14.860 210.610 14.920 ;
        RECT 179.560 14.720 210.610 14.860 ;
        RECT 210.290 14.660 210.610 14.720 ;
      LAYER via ;
        RECT 210.320 1483.460 210.580 1483.720 ;
        RECT 536.460 1483.460 536.720 1483.720 ;
        RECT 145.460 15.340 145.720 15.600 ;
        RECT 210.320 14.660 210.580 14.920 ;
      LAYER met2 ;
        RECT 537.910 1500.490 538.190 1504.000 ;
        RECT 536.520 1500.350 538.190 1500.490 ;
        RECT 536.520 1483.750 536.660 1500.350 ;
        RECT 537.910 1500.000 538.190 1500.350 ;
        RECT 210.320 1483.430 210.580 1483.750 ;
        RECT 536.460 1483.430 536.720 1483.750 ;
        RECT 145.460 15.310 145.720 15.630 ;
        RECT 145.520 2.400 145.660 15.310 ;
        RECT 210.380 14.950 210.520 1483.430 ;
        RECT 210.320 14.630 210.580 14.950 ;
        RECT 145.310 -4.800 145.870 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 538.270 18.940 538.590 19.000 ;
        RECT 565.870 18.940 566.190 19.000 ;
        RECT 538.270 18.800 566.190 18.940 ;
        RECT 538.270 18.740 538.590 18.800 ;
        RECT 565.870 18.740 566.190 18.800 ;
        RECT 163.370 17.920 163.690 17.980 ;
        RECT 538.270 17.920 538.590 17.980 ;
        RECT 163.370 17.780 538.590 17.920 ;
        RECT 163.370 17.720 163.690 17.780 ;
        RECT 538.270 17.720 538.590 17.780 ;
      LAYER via ;
        RECT 538.300 18.740 538.560 19.000 ;
        RECT 565.900 18.740 566.160 19.000 ;
        RECT 163.400 17.720 163.660 17.980 ;
        RECT 538.300 17.720 538.560 17.980 ;
      LAYER met2 ;
        RECT 567.350 1500.490 567.630 1504.000 ;
        RECT 565.960 1500.350 567.630 1500.490 ;
        RECT 565.960 19.030 566.100 1500.350 ;
        RECT 567.350 1500.000 567.630 1500.350 ;
        RECT 538.300 18.710 538.560 19.030 ;
        RECT 565.900 18.710 566.160 19.030 ;
        RECT 538.360 18.010 538.500 18.710 ;
        RECT 163.400 17.690 163.660 18.010 ;
        RECT 538.300 17.690 538.560 18.010 ;
        RECT 163.460 2.400 163.600 17.690 ;
        RECT 163.250 -4.800 163.810 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 226.850 17.580 227.170 17.640 ;
        RECT 373.130 17.580 373.450 17.640 ;
        RECT 226.850 17.440 373.450 17.580 ;
        RECT 226.850 17.380 227.170 17.440 ;
        RECT 373.130 17.380 373.450 17.440 ;
        RECT 420.050 17.580 420.370 17.640 ;
        RECT 469.730 17.580 470.050 17.640 ;
        RECT 420.050 17.440 470.050 17.580 ;
        RECT 420.050 17.380 420.370 17.440 ;
        RECT 469.730 17.380 470.050 17.440 ;
        RECT 497.330 17.580 497.650 17.640 ;
        RECT 593.930 17.580 594.250 17.640 ;
        RECT 497.330 17.440 594.250 17.580 ;
        RECT 497.330 17.380 497.650 17.440 ;
        RECT 593.930 17.380 594.250 17.440 ;
        RECT 180.850 16.220 181.170 16.280 ;
        RECT 226.850 16.220 227.170 16.280 ;
        RECT 180.850 16.080 227.170 16.220 ;
        RECT 180.850 16.020 181.170 16.080 ;
        RECT 226.850 16.020 227.170 16.080 ;
      LAYER via ;
        RECT 226.880 17.380 227.140 17.640 ;
        RECT 373.160 17.380 373.420 17.640 ;
        RECT 420.080 17.380 420.340 17.640 ;
        RECT 469.760 17.380 470.020 17.640 ;
        RECT 497.360 17.380 497.620 17.640 ;
        RECT 593.960 17.380 594.220 17.640 ;
        RECT 180.880 16.020 181.140 16.280 ;
        RECT 226.880 16.020 227.140 16.280 ;
      LAYER met2 ;
        RECT 596.330 1500.490 596.610 1504.000 ;
        RECT 594.020 1500.350 596.610 1500.490 ;
        RECT 373.150 17.835 373.430 18.205 ;
        RECT 420.070 17.835 420.350 18.205 ;
        RECT 373.220 17.670 373.360 17.835 ;
        RECT 420.140 17.670 420.280 17.835 ;
        RECT 594.020 17.670 594.160 1500.350 ;
        RECT 596.330 1500.000 596.610 1500.350 ;
        RECT 226.880 17.350 227.140 17.670 ;
        RECT 373.160 17.350 373.420 17.670 ;
        RECT 420.080 17.350 420.340 17.670 ;
        RECT 469.760 17.350 470.020 17.670 ;
        RECT 497.360 17.350 497.620 17.670 ;
        RECT 593.960 17.350 594.220 17.670 ;
        RECT 226.940 16.310 227.080 17.350 ;
        RECT 180.880 15.990 181.140 16.310 ;
        RECT 226.880 15.990 227.140 16.310 ;
        RECT 469.820 16.165 469.960 17.350 ;
        RECT 497.420 16.165 497.560 17.350 ;
        RECT 180.940 2.400 181.080 15.990 ;
        RECT 469.750 15.795 470.030 16.165 ;
        RECT 497.350 15.795 497.630 16.165 ;
        RECT 180.730 -4.800 181.290 2.400 ;
      LAYER via2 ;
        RECT 373.150 17.880 373.430 18.160 ;
        RECT 420.070 17.880 420.350 18.160 ;
        RECT 469.750 15.840 470.030 16.120 ;
        RECT 497.350 15.840 497.630 16.120 ;
      LAYER met3 ;
        RECT 373.125 18.170 373.455 18.185 ;
        RECT 420.045 18.170 420.375 18.185 ;
        RECT 373.125 17.870 420.375 18.170 ;
        RECT 373.125 17.855 373.455 17.870 ;
        RECT 420.045 17.855 420.375 17.870 ;
        RECT 469.725 16.130 470.055 16.145 ;
        RECT 497.325 16.130 497.655 16.145 ;
        RECT 469.725 15.830 497.655 16.130 ;
        RECT 469.725 15.815 470.055 15.830 ;
        RECT 497.325 15.815 497.655 15.830 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 199.710 1484.000 200.030 1484.060 ;
        RECT 623.830 1484.000 624.150 1484.060 ;
        RECT 199.710 1483.860 624.150 1484.000 ;
        RECT 199.710 1483.800 200.030 1483.860 ;
        RECT 623.830 1483.800 624.150 1483.860 ;
      LAYER via ;
        RECT 199.740 1483.800 200.000 1484.060 ;
        RECT 623.860 1483.800 624.120 1484.060 ;
      LAYER met2 ;
        RECT 625.770 1500.490 626.050 1504.000 ;
        RECT 623.920 1500.350 626.050 1500.490 ;
        RECT 623.920 1484.090 624.060 1500.350 ;
        RECT 625.770 1500.000 626.050 1500.350 ;
        RECT 199.740 1483.770 200.000 1484.090 ;
        RECT 623.860 1483.770 624.120 1484.090 ;
        RECT 199.800 16.730 199.940 1483.770 ;
        RECT 198.880 16.590 199.940 16.730 ;
        RECT 198.880 2.400 199.020 16.590 ;
        RECT 198.670 -4.800 199.230 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 216.730 14.180 217.050 14.240 ;
        RECT 649.130 14.180 649.450 14.240 ;
        RECT 216.730 14.040 620.840 14.180 ;
        RECT 216.730 13.980 217.050 14.040 ;
        RECT 620.700 13.840 620.840 14.040 ;
        RECT 639.100 14.040 649.450 14.180 ;
        RECT 639.100 13.840 639.240 14.040 ;
        RECT 649.130 13.980 649.450 14.040 ;
        RECT 620.700 13.700 639.240 13.840 ;
      LAYER via ;
        RECT 216.760 13.980 217.020 14.240 ;
        RECT 649.160 13.980 649.420 14.240 ;
      LAYER met2 ;
        RECT 654.750 1500.490 655.030 1504.000 ;
        RECT 649.220 1500.350 655.030 1500.490 ;
        RECT 649.220 14.270 649.360 1500.350 ;
        RECT 654.750 1500.000 655.030 1500.350 ;
        RECT 216.760 13.950 217.020 14.270 ;
        RECT 649.160 13.950 649.420 14.270 ;
        RECT 216.820 2.400 216.960 13.950 ;
        RECT 216.610 -4.800 217.170 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 240.650 1484.340 240.970 1484.400 ;
        RECT 684.090 1484.340 684.410 1484.400 ;
        RECT 240.650 1484.200 684.410 1484.340 ;
        RECT 240.650 1484.140 240.970 1484.200 ;
        RECT 684.090 1484.140 684.410 1484.200 ;
        RECT 234.670 17.240 234.990 17.300 ;
        RECT 240.650 17.240 240.970 17.300 ;
        RECT 234.670 17.100 240.970 17.240 ;
        RECT 234.670 17.040 234.990 17.100 ;
        RECT 240.650 17.040 240.970 17.100 ;
      LAYER via ;
        RECT 240.680 1484.140 240.940 1484.400 ;
        RECT 684.120 1484.140 684.380 1484.400 ;
        RECT 234.700 17.040 234.960 17.300 ;
        RECT 240.680 17.040 240.940 17.300 ;
      LAYER met2 ;
        RECT 684.190 1500.420 684.470 1504.000 ;
        RECT 684.180 1500.000 684.470 1500.420 ;
        RECT 684.180 1484.430 684.320 1500.000 ;
        RECT 240.680 1484.110 240.940 1484.430 ;
        RECT 684.120 1484.110 684.380 1484.430 ;
        RECT 240.740 17.330 240.880 1484.110 ;
        RECT 234.700 17.010 234.960 17.330 ;
        RECT 240.680 17.010 240.940 17.330 ;
        RECT 234.760 2.400 234.900 17.010 ;
        RECT 234.550 -4.800 235.110 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 161.990 1490.120 162.310 1490.180 ;
        RECT 391.990 1490.120 392.310 1490.180 ;
        RECT 161.990 1489.980 392.310 1490.120 ;
        RECT 161.990 1489.920 162.310 1489.980 ;
        RECT 391.990 1489.920 392.310 1489.980 ;
        RECT 56.190 17.240 56.510 17.300 ;
        RECT 161.990 17.240 162.310 17.300 ;
        RECT 56.190 17.100 162.310 17.240 ;
        RECT 56.190 17.040 56.510 17.100 ;
        RECT 161.990 17.040 162.310 17.100 ;
      LAYER via ;
        RECT 162.020 1489.920 162.280 1490.180 ;
        RECT 392.020 1489.920 392.280 1490.180 ;
        RECT 56.220 17.040 56.480 17.300 ;
        RECT 162.020 17.040 162.280 17.300 ;
      LAYER met2 ;
        RECT 392.090 1500.420 392.370 1504.000 ;
        RECT 392.080 1500.000 392.370 1500.420 ;
        RECT 392.080 1490.210 392.220 1500.000 ;
        RECT 162.020 1489.890 162.280 1490.210 ;
        RECT 392.020 1489.890 392.280 1490.210 ;
        RECT 162.080 17.330 162.220 1489.890 ;
        RECT 56.220 17.010 56.480 17.330 ;
        RECT 162.020 17.010 162.280 17.330 ;
        RECT 56.280 2.400 56.420 17.010 ;
        RECT 56.070 -4.800 56.630 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 82.410 1489.100 82.730 1489.160 ;
        RECT 431.090 1489.100 431.410 1489.160 ;
        RECT 82.410 1488.960 431.410 1489.100 ;
        RECT 82.410 1488.900 82.730 1488.960 ;
        RECT 431.090 1488.900 431.410 1488.960 ;
        RECT 80.110 17.580 80.430 17.640 ;
        RECT 82.410 17.580 82.730 17.640 ;
        RECT 80.110 17.440 82.730 17.580 ;
        RECT 80.110 17.380 80.430 17.440 ;
        RECT 82.410 17.380 82.730 17.440 ;
      LAYER via ;
        RECT 82.440 1488.900 82.700 1489.160 ;
        RECT 431.120 1488.900 431.380 1489.160 ;
        RECT 80.140 17.380 80.400 17.640 ;
        RECT 82.440 17.380 82.700 17.640 ;
      LAYER met2 ;
        RECT 431.190 1500.420 431.470 1504.000 ;
        RECT 431.180 1500.000 431.470 1500.420 ;
        RECT 431.180 1489.190 431.320 1500.000 ;
        RECT 82.440 1488.870 82.700 1489.190 ;
        RECT 431.120 1488.870 431.380 1489.190 ;
        RECT 82.500 17.670 82.640 1488.870 ;
        RECT 80.140 17.350 80.400 17.670 ;
        RECT 82.440 17.350 82.700 17.670 ;
        RECT 80.200 2.400 80.340 17.350 ;
        RECT 79.990 -4.800 80.550 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 109.550 1487.740 109.870 1487.800 ;
        RECT 469.730 1487.740 470.050 1487.800 ;
        RECT 109.550 1487.600 470.050 1487.740 ;
        RECT 109.550 1487.540 109.870 1487.600 ;
        RECT 469.730 1487.540 470.050 1487.600 ;
        RECT 103.570 17.580 103.890 17.640 ;
        RECT 109.550 17.580 109.870 17.640 ;
        RECT 103.570 17.440 109.870 17.580 ;
        RECT 103.570 17.380 103.890 17.440 ;
        RECT 109.550 17.380 109.870 17.440 ;
      LAYER via ;
        RECT 109.580 1487.540 109.840 1487.800 ;
        RECT 469.760 1487.540 470.020 1487.800 ;
        RECT 103.600 17.380 103.860 17.640 ;
        RECT 109.580 17.380 109.840 17.640 ;
      LAYER met2 ;
        RECT 469.830 1500.420 470.110 1504.000 ;
        RECT 469.820 1500.000 470.110 1500.420 ;
        RECT 469.820 1487.830 469.960 1500.000 ;
        RECT 109.580 1487.510 109.840 1487.830 ;
        RECT 469.760 1487.510 470.020 1487.830 ;
        RECT 109.640 17.670 109.780 1487.510 ;
        RECT 103.600 17.350 103.860 17.670 ;
        RECT 109.580 17.350 109.840 17.670 ;
        RECT 103.660 2.400 103.800 17.350 ;
        RECT 103.450 -4.800 104.010 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 130.710 1487.060 131.030 1487.120 ;
        RECT 508.830 1487.060 509.150 1487.120 ;
        RECT 130.710 1486.920 509.150 1487.060 ;
        RECT 130.710 1486.860 131.030 1486.920 ;
        RECT 508.830 1486.860 509.150 1486.920 ;
        RECT 127.490 19.280 127.810 19.340 ;
        RECT 130.710 19.280 131.030 19.340 ;
        RECT 127.490 19.140 131.030 19.280 ;
        RECT 127.490 19.080 127.810 19.140 ;
        RECT 130.710 19.080 131.030 19.140 ;
      LAYER via ;
        RECT 130.740 1486.860 131.000 1487.120 ;
        RECT 508.860 1486.860 509.120 1487.120 ;
        RECT 127.520 19.080 127.780 19.340 ;
        RECT 130.740 19.080 131.000 19.340 ;
      LAYER met2 ;
        RECT 508.930 1500.420 509.210 1504.000 ;
        RECT 508.920 1500.000 509.210 1500.420 ;
        RECT 508.920 1487.150 509.060 1500.000 ;
        RECT 130.740 1486.830 131.000 1487.150 ;
        RECT 508.860 1486.830 509.120 1487.150 ;
        RECT 130.800 19.370 130.940 1486.830 ;
        RECT 127.520 19.050 127.780 19.370 ;
        RECT 130.740 19.050 131.000 19.370 ;
        RECT 127.580 2.400 127.720 19.050 ;
        RECT 127.370 -4.800 127.930 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 196.490 1490.460 196.810 1490.520 ;
        RECT 343.230 1490.460 343.550 1490.520 ;
        RECT 196.490 1490.320 343.550 1490.460 ;
        RECT 196.490 1490.260 196.810 1490.320 ;
        RECT 343.230 1490.260 343.550 1490.320 ;
        RECT 26.290 15.880 26.610 15.940 ;
        RECT 26.290 15.740 121.740 15.880 ;
        RECT 26.290 15.680 26.610 15.740 ;
        RECT 121.600 15.540 121.740 15.740 ;
        RECT 134.020 15.740 180.620 15.880 ;
        RECT 134.020 15.540 134.160 15.740 ;
        RECT 121.600 15.400 134.160 15.540 ;
        RECT 180.480 15.540 180.620 15.740 ;
        RECT 196.490 15.540 196.810 15.600 ;
        RECT 180.480 15.400 196.810 15.540 ;
        RECT 196.490 15.340 196.810 15.400 ;
      LAYER via ;
        RECT 196.520 1490.260 196.780 1490.520 ;
        RECT 343.260 1490.260 343.520 1490.520 ;
        RECT 26.320 15.680 26.580 15.940 ;
        RECT 196.520 15.340 196.780 15.600 ;
      LAYER met2 ;
        RECT 343.330 1500.420 343.610 1504.000 ;
        RECT 343.320 1500.000 343.610 1500.420 ;
        RECT 343.320 1490.550 343.460 1500.000 ;
        RECT 196.520 1490.230 196.780 1490.550 ;
        RECT 343.260 1490.230 343.520 1490.550 ;
        RECT 26.320 15.650 26.580 15.970 ;
        RECT 26.380 2.400 26.520 15.650 ;
        RECT 196.580 15.630 196.720 1490.230 ;
        RECT 196.520 15.310 196.780 15.630 ;
        RECT 26.170 -4.800 26.730 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 259.050 1486.720 259.370 1486.780 ;
        RECT 352.890 1486.720 353.210 1486.780 ;
        RECT 259.050 1486.580 353.210 1486.720 ;
        RECT 259.050 1486.520 259.370 1486.580 ;
        RECT 352.890 1486.520 353.210 1486.580 ;
        RECT 32.270 16.220 32.590 16.280 ;
        RECT 34.570 16.220 34.890 16.280 ;
        RECT 32.270 16.080 34.890 16.220 ;
        RECT 32.270 16.020 32.590 16.080 ;
        RECT 34.570 16.020 34.890 16.080 ;
        RECT 106.790 16.220 107.110 16.280 ;
        RECT 179.470 16.220 179.790 16.280 ;
        RECT 106.790 16.080 179.790 16.220 ;
        RECT 106.790 16.020 107.110 16.080 ;
        RECT 179.470 16.020 179.790 16.080 ;
        RECT 34.570 15.540 34.890 15.600 ;
        RECT 106.790 15.540 107.110 15.600 ;
        RECT 34.570 15.400 107.110 15.540 ;
        RECT 34.570 15.340 34.890 15.400 ;
        RECT 106.790 15.340 107.110 15.400 ;
        RECT 179.930 15.200 180.250 15.260 ;
        RECT 259.050 15.200 259.370 15.260 ;
        RECT 179.930 15.060 259.370 15.200 ;
        RECT 179.930 15.000 180.250 15.060 ;
        RECT 259.050 15.000 259.370 15.060 ;
      LAYER via ;
        RECT 259.080 1486.520 259.340 1486.780 ;
        RECT 352.920 1486.520 353.180 1486.780 ;
        RECT 32.300 16.020 32.560 16.280 ;
        RECT 34.600 16.020 34.860 16.280 ;
        RECT 106.820 16.020 107.080 16.280 ;
        RECT 179.500 16.020 179.760 16.280 ;
        RECT 34.600 15.340 34.860 15.600 ;
        RECT 106.820 15.340 107.080 15.600 ;
        RECT 179.960 15.000 180.220 15.260 ;
        RECT 259.080 15.000 259.340 15.260 ;
      LAYER met2 ;
        RECT 352.990 1500.420 353.270 1504.000 ;
        RECT 352.980 1500.000 353.270 1500.420 ;
        RECT 352.980 1486.810 353.120 1500.000 ;
        RECT 259.080 1486.490 259.340 1486.810 ;
        RECT 352.920 1486.490 353.180 1486.810 ;
        RECT 32.300 15.990 32.560 16.310 ;
        RECT 34.600 15.990 34.860 16.310 ;
        RECT 106.820 15.990 107.080 16.310 ;
        RECT 179.500 16.050 179.760 16.310 ;
        RECT 179.500 15.990 180.160 16.050 ;
        RECT 32.360 2.400 32.500 15.990 ;
        RECT 34.660 15.630 34.800 15.990 ;
        RECT 106.880 15.630 107.020 15.990 ;
        RECT 179.560 15.910 180.160 15.990 ;
        RECT 34.600 15.310 34.860 15.630 ;
        RECT 106.820 15.310 107.080 15.630 ;
        RECT 180.020 15.290 180.160 15.910 ;
        RECT 259.140 15.290 259.280 1486.490 ;
        RECT 179.960 14.970 180.220 15.290 ;
        RECT 259.080 14.970 259.340 15.290 ;
        RECT 32.150 -4.800 32.710 2.400 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 681.480 3243.600 684.050 3244.660 ;
        RECT 1331.480 3243.600 1334.050 3244.660 ;
        RECT 1931.480 3243.600 1934.050 3244.660 ;
        RECT 2581.480 3243.600 2584.050 3244.660 ;
      LAYER via3 ;
        RECT 682.500 3243.620 684.020 3244.630 ;
        RECT 1332.500 3243.620 1334.020 3244.630 ;
        RECT 1932.500 3243.620 1934.020 3244.630 ;
        RECT 2582.500 3243.620 2584.020 3244.630 ;
      LAYER met4 ;
        RECT -38.180 -32.820 -35.180 3552.500 ;
        RECT -28.780 -23.420 -25.780 3543.100 ;
        RECT -19.380 -14.020 -16.380 3533.700 ;
        RECT -9.980 -4.620 -6.980 3524.300 ;
        RECT 4.020 -9.320 7.020 3529.000 ;
        RECT 22.020 -18.720 25.020 3538.400 ;
        RECT 40.020 -28.120 43.020 3547.800 ;
        RECT 58.020 -37.520 61.020 3557.200 ;
        RECT 184.020 -9.320 187.020 3529.000 ;
        RECT 202.020 -18.720 205.020 3538.400 ;
        RECT 220.020 -28.120 223.020 3547.800 ;
        RECT 238.020 -37.520 241.020 3557.200 ;
        RECT 364.020 3271.235 367.020 3529.000 ;
        RECT 382.020 3271.235 385.020 3538.400 ;
        RECT 400.020 3271.235 403.020 3547.800 ;
        RECT 418.020 3271.235 421.020 3557.200 ;
        RECT 544.020 3271.235 547.020 3529.000 ;
        RECT 562.020 3271.235 565.020 3538.400 ;
        RECT 580.020 3271.235 583.020 3547.800 ;
        RECT 598.020 3271.235 601.020 3557.200 ;
        RECT 682.470 2803.670 684.070 3244.680 ;
        RECT 382.020 2715.000 385.020 2785.000 ;
        RECT 400.020 2715.000 403.020 2785.000 ;
        RECT 418.020 2715.000 421.020 2785.000 ;
        RECT 562.020 2715.000 565.020 2785.000 ;
        RECT 580.020 2715.000 583.020 2785.000 ;
        RECT 598.020 2715.000 601.020 2785.000 ;
        RECT 724.020 2715.000 727.020 3529.000 ;
        RECT 742.020 2715.000 745.020 3538.400 ;
        RECT 760.020 2715.000 763.020 3547.800 ;
        RECT 778.020 2715.000 781.020 3557.200 ;
        RECT 904.020 2715.000 907.020 3529.000 ;
        RECT 922.020 2715.000 925.020 3538.400 ;
        RECT 940.020 3271.235 943.020 3547.800 ;
        RECT 958.020 3271.235 961.020 3557.200 ;
        RECT 1084.020 3271.235 1087.020 3529.000 ;
        RECT 1102.020 3271.235 1105.020 3538.400 ;
        RECT 1120.020 3271.235 1123.020 3547.800 ;
        RECT 1138.020 3271.235 1141.020 3557.200 ;
        RECT 1264.020 3271.235 1267.020 3529.000 ;
        RECT 1282.020 3271.235 1285.020 3538.400 ;
        RECT 1300.020 3271.235 1303.020 3547.800 ;
        RECT 1318.020 3271.235 1321.020 3557.200 ;
        RECT 1332.470 2803.670 1334.070 3244.680 ;
        RECT 940.020 2715.000 943.020 2785.000 ;
        RECT 958.020 2715.000 961.020 2785.000 ;
        RECT 1102.020 2715.000 1105.020 2785.000 ;
        RECT 1120.020 2715.000 1123.020 2785.000 ;
        RECT 1138.020 2715.000 1141.020 2785.000 ;
        RECT 1282.020 2715.000 1285.020 2785.000 ;
        RECT 1300.020 2715.000 1303.020 2785.000 ;
        RECT 1318.020 2715.000 1321.020 2785.000 ;
        RECT 321.040 1510.640 322.640 2688.880 ;
        RECT 364.020 -9.320 367.020 1485.000 ;
        RECT 382.020 -18.720 385.020 1485.000 ;
        RECT 400.020 -28.120 403.020 1485.000 ;
        RECT 418.020 -37.520 421.020 1485.000 ;
        RECT 544.020 -9.320 547.020 1485.000 ;
        RECT 562.020 -18.720 565.020 1485.000 ;
        RECT 580.020 -28.120 583.020 1485.000 ;
        RECT 598.020 -37.520 601.020 1485.000 ;
        RECT 724.020 -9.320 727.020 1485.000 ;
        RECT 742.020 -18.720 745.020 1485.000 ;
        RECT 760.020 -28.120 763.020 1485.000 ;
        RECT 778.020 -37.520 781.020 1485.000 ;
        RECT 904.020 -9.320 907.020 1485.000 ;
        RECT 922.020 -18.720 925.020 1485.000 ;
        RECT 940.020 -28.120 943.020 1485.000 ;
        RECT 958.020 -37.520 961.020 1485.000 ;
        RECT 1084.020 -9.320 1087.020 1485.000 ;
        RECT 1102.020 -18.720 1105.020 1485.000 ;
        RECT 1120.020 -28.120 1123.020 1485.000 ;
        RECT 1138.020 -37.520 1141.020 1485.000 ;
        RECT 1264.020 -9.320 1267.020 1485.000 ;
        RECT 1282.020 -18.720 1285.020 1485.000 ;
        RECT 1300.020 -28.120 1303.020 1485.000 ;
        RECT 1318.020 -37.520 1321.020 1485.000 ;
        RECT 1444.020 -9.320 1447.020 3529.000 ;
        RECT 1462.020 -18.720 1465.020 3538.400 ;
        RECT 1480.020 -28.120 1483.020 3547.800 ;
        RECT 1498.020 -37.520 1501.020 3557.200 ;
        RECT 1624.020 3271.235 1627.020 3529.000 ;
        RECT 1642.020 3271.235 1645.020 3538.400 ;
        RECT 1660.020 3271.235 1663.020 3547.800 ;
        RECT 1678.020 3271.235 1681.020 3557.200 ;
        RECT 1804.020 3271.235 1807.020 3529.000 ;
        RECT 1822.020 3271.235 1825.020 3538.400 ;
        RECT 1840.020 3271.235 1843.020 3547.800 ;
        RECT 1858.020 3271.235 1861.020 3557.200 ;
        RECT 1932.470 2803.670 1934.070 3244.680 ;
        RECT 1624.020 -9.320 1627.020 2785.000 ;
        RECT 1642.020 -18.720 1645.020 2785.000 ;
        RECT 1660.020 -28.120 1663.020 2785.000 ;
        RECT 1678.020 -37.520 1681.020 2785.000 ;
        RECT 1804.020 -9.320 1807.020 2785.000 ;
        RECT 1822.020 -18.720 1825.020 2785.000 ;
        RECT 1840.020 -28.120 1843.020 2785.000 ;
        RECT 1858.020 -37.520 1861.020 2785.000 ;
        RECT 1984.020 -9.320 1987.020 3529.000 ;
        RECT 2002.020 -18.720 2005.020 3538.400 ;
        RECT 2020.020 -28.120 2023.020 3547.800 ;
        RECT 2038.020 -37.520 2041.020 3557.200 ;
        RECT 2164.020 -9.320 2167.020 3529.000 ;
        RECT 2182.020 3271.235 2185.020 3538.400 ;
        RECT 2200.020 3271.235 2203.020 3547.800 ;
        RECT 2218.020 3271.235 2221.020 3557.200 ;
        RECT 2344.020 3271.235 2347.020 3529.000 ;
        RECT 2362.020 3271.235 2365.020 3538.400 ;
        RECT 2380.020 3271.235 2383.020 3547.800 ;
        RECT 2398.020 3271.235 2401.020 3557.200 ;
        RECT 2524.020 3271.235 2527.020 3529.000 ;
        RECT 2542.020 3271.235 2545.020 3538.400 ;
        RECT 2560.020 3271.235 2563.020 3547.800 ;
        RECT 2578.020 3271.235 2581.020 3557.200 ;
        RECT 2582.470 2803.670 2584.070 3244.680 ;
        RECT 2182.020 -18.720 2185.020 2785.000 ;
        RECT 2200.020 -28.120 2203.020 2785.000 ;
        RECT 2218.020 -37.520 2221.020 2785.000 ;
        RECT 2344.020 -9.320 2347.020 2785.000 ;
        RECT 2362.020 -18.720 2365.020 2785.000 ;
        RECT 2380.020 -28.120 2383.020 2785.000 ;
        RECT 2398.020 -37.520 2401.020 2785.000 ;
        RECT 2524.020 -9.320 2527.020 2785.000 ;
        RECT 2542.020 -18.720 2545.020 2785.000 ;
        RECT 2560.020 -28.120 2563.020 2785.000 ;
        RECT 2578.020 -37.520 2581.020 2785.000 ;
        RECT 2704.020 -9.320 2707.020 3529.000 ;
        RECT 2722.020 -18.720 2725.020 3538.400 ;
        RECT 2740.020 -28.120 2743.020 3547.800 ;
        RECT 2758.020 -37.520 2761.020 3557.200 ;
        RECT 2884.020 -9.320 2887.020 3529.000 ;
        RECT 2902.020 -18.720 2905.020 3538.400 ;
        RECT 2926.600 -4.620 2929.600 3524.300 ;
        RECT 2936.000 -14.020 2939.000 3533.700 ;
        RECT 2945.400 -23.420 2948.400 3543.100 ;
        RECT 2954.800 -32.820 2957.800 3552.500 ;
      LAYER via4 ;
        RECT -37.270 3551.210 -36.090 3552.390 ;
        RECT -37.270 3549.610 -36.090 3550.790 ;
        RECT 58.930 3551.210 60.110 3552.390 ;
        RECT 58.930 3549.610 60.110 3550.790 ;
        RECT -37.270 3485.090 -36.090 3486.270 ;
        RECT -37.270 3483.490 -36.090 3484.670 ;
        RECT -37.270 3305.090 -36.090 3306.270 ;
        RECT -37.270 3303.490 -36.090 3304.670 ;
        RECT -37.270 3125.090 -36.090 3126.270 ;
        RECT -37.270 3123.490 -36.090 3124.670 ;
        RECT -37.270 2945.090 -36.090 2946.270 ;
        RECT -37.270 2943.490 -36.090 2944.670 ;
        RECT -37.270 2765.090 -36.090 2766.270 ;
        RECT -37.270 2763.490 -36.090 2764.670 ;
        RECT -37.270 2585.090 -36.090 2586.270 ;
        RECT -37.270 2583.490 -36.090 2584.670 ;
        RECT -37.270 2405.090 -36.090 2406.270 ;
        RECT -37.270 2403.490 -36.090 2404.670 ;
        RECT -37.270 2225.090 -36.090 2226.270 ;
        RECT -37.270 2223.490 -36.090 2224.670 ;
        RECT -37.270 2045.090 -36.090 2046.270 ;
        RECT -37.270 2043.490 -36.090 2044.670 ;
        RECT -37.270 1865.090 -36.090 1866.270 ;
        RECT -37.270 1863.490 -36.090 1864.670 ;
        RECT -37.270 1685.090 -36.090 1686.270 ;
        RECT -37.270 1683.490 -36.090 1684.670 ;
        RECT -37.270 1505.090 -36.090 1506.270 ;
        RECT -37.270 1503.490 -36.090 1504.670 ;
        RECT -37.270 1325.090 -36.090 1326.270 ;
        RECT -37.270 1323.490 -36.090 1324.670 ;
        RECT -37.270 1145.090 -36.090 1146.270 ;
        RECT -37.270 1143.490 -36.090 1144.670 ;
        RECT -37.270 965.090 -36.090 966.270 ;
        RECT -37.270 963.490 -36.090 964.670 ;
        RECT -37.270 785.090 -36.090 786.270 ;
        RECT -37.270 783.490 -36.090 784.670 ;
        RECT -37.270 605.090 -36.090 606.270 ;
        RECT -37.270 603.490 -36.090 604.670 ;
        RECT -37.270 425.090 -36.090 426.270 ;
        RECT -37.270 423.490 -36.090 424.670 ;
        RECT -37.270 245.090 -36.090 246.270 ;
        RECT -37.270 243.490 -36.090 244.670 ;
        RECT -37.270 65.090 -36.090 66.270 ;
        RECT -37.270 63.490 -36.090 64.670 ;
        RECT -27.870 3541.810 -26.690 3542.990 ;
        RECT -27.870 3540.210 -26.690 3541.390 ;
        RECT 40.930 3541.810 42.110 3542.990 ;
        RECT 40.930 3540.210 42.110 3541.390 ;
        RECT -27.870 3467.090 -26.690 3468.270 ;
        RECT -27.870 3465.490 -26.690 3466.670 ;
        RECT -27.870 3287.090 -26.690 3288.270 ;
        RECT -27.870 3285.490 -26.690 3286.670 ;
        RECT -27.870 3107.090 -26.690 3108.270 ;
        RECT -27.870 3105.490 -26.690 3106.670 ;
        RECT -27.870 2927.090 -26.690 2928.270 ;
        RECT -27.870 2925.490 -26.690 2926.670 ;
        RECT -27.870 2747.090 -26.690 2748.270 ;
        RECT -27.870 2745.490 -26.690 2746.670 ;
        RECT -27.870 2567.090 -26.690 2568.270 ;
        RECT -27.870 2565.490 -26.690 2566.670 ;
        RECT -27.870 2387.090 -26.690 2388.270 ;
        RECT -27.870 2385.490 -26.690 2386.670 ;
        RECT -27.870 2207.090 -26.690 2208.270 ;
        RECT -27.870 2205.490 -26.690 2206.670 ;
        RECT -27.870 2027.090 -26.690 2028.270 ;
        RECT -27.870 2025.490 -26.690 2026.670 ;
        RECT -27.870 1847.090 -26.690 1848.270 ;
        RECT -27.870 1845.490 -26.690 1846.670 ;
        RECT -27.870 1667.090 -26.690 1668.270 ;
        RECT -27.870 1665.490 -26.690 1666.670 ;
        RECT -27.870 1487.090 -26.690 1488.270 ;
        RECT -27.870 1485.490 -26.690 1486.670 ;
        RECT -27.870 1307.090 -26.690 1308.270 ;
        RECT -27.870 1305.490 -26.690 1306.670 ;
        RECT -27.870 1127.090 -26.690 1128.270 ;
        RECT -27.870 1125.490 -26.690 1126.670 ;
        RECT -27.870 947.090 -26.690 948.270 ;
        RECT -27.870 945.490 -26.690 946.670 ;
        RECT -27.870 767.090 -26.690 768.270 ;
        RECT -27.870 765.490 -26.690 766.670 ;
        RECT -27.870 587.090 -26.690 588.270 ;
        RECT -27.870 585.490 -26.690 586.670 ;
        RECT -27.870 407.090 -26.690 408.270 ;
        RECT -27.870 405.490 -26.690 406.670 ;
        RECT -27.870 227.090 -26.690 228.270 ;
        RECT -27.870 225.490 -26.690 226.670 ;
        RECT -27.870 47.090 -26.690 48.270 ;
        RECT -27.870 45.490 -26.690 46.670 ;
        RECT -18.470 3532.410 -17.290 3533.590 ;
        RECT -18.470 3530.810 -17.290 3531.990 ;
        RECT 22.930 3532.410 24.110 3533.590 ;
        RECT 22.930 3530.810 24.110 3531.990 ;
        RECT -18.470 3449.090 -17.290 3450.270 ;
        RECT -18.470 3447.490 -17.290 3448.670 ;
        RECT -18.470 3269.090 -17.290 3270.270 ;
        RECT -18.470 3267.490 -17.290 3268.670 ;
        RECT -18.470 3089.090 -17.290 3090.270 ;
        RECT -18.470 3087.490 -17.290 3088.670 ;
        RECT -18.470 2909.090 -17.290 2910.270 ;
        RECT -18.470 2907.490 -17.290 2908.670 ;
        RECT -18.470 2729.090 -17.290 2730.270 ;
        RECT -18.470 2727.490 -17.290 2728.670 ;
        RECT -18.470 2549.090 -17.290 2550.270 ;
        RECT -18.470 2547.490 -17.290 2548.670 ;
        RECT -18.470 2369.090 -17.290 2370.270 ;
        RECT -18.470 2367.490 -17.290 2368.670 ;
        RECT -18.470 2189.090 -17.290 2190.270 ;
        RECT -18.470 2187.490 -17.290 2188.670 ;
        RECT -18.470 2009.090 -17.290 2010.270 ;
        RECT -18.470 2007.490 -17.290 2008.670 ;
        RECT -18.470 1829.090 -17.290 1830.270 ;
        RECT -18.470 1827.490 -17.290 1828.670 ;
        RECT -18.470 1649.090 -17.290 1650.270 ;
        RECT -18.470 1647.490 -17.290 1648.670 ;
        RECT -18.470 1469.090 -17.290 1470.270 ;
        RECT -18.470 1467.490 -17.290 1468.670 ;
        RECT -18.470 1289.090 -17.290 1290.270 ;
        RECT -18.470 1287.490 -17.290 1288.670 ;
        RECT -18.470 1109.090 -17.290 1110.270 ;
        RECT -18.470 1107.490 -17.290 1108.670 ;
        RECT -18.470 929.090 -17.290 930.270 ;
        RECT -18.470 927.490 -17.290 928.670 ;
        RECT -18.470 749.090 -17.290 750.270 ;
        RECT -18.470 747.490 -17.290 748.670 ;
        RECT -18.470 569.090 -17.290 570.270 ;
        RECT -18.470 567.490 -17.290 568.670 ;
        RECT -18.470 389.090 -17.290 390.270 ;
        RECT -18.470 387.490 -17.290 388.670 ;
        RECT -18.470 209.090 -17.290 210.270 ;
        RECT -18.470 207.490 -17.290 208.670 ;
        RECT -18.470 29.090 -17.290 30.270 ;
        RECT -18.470 27.490 -17.290 28.670 ;
        RECT -9.070 3523.010 -7.890 3524.190 ;
        RECT -9.070 3521.410 -7.890 3522.590 ;
        RECT -9.070 3431.090 -7.890 3432.270 ;
        RECT -9.070 3429.490 -7.890 3430.670 ;
        RECT -9.070 3251.090 -7.890 3252.270 ;
        RECT -9.070 3249.490 -7.890 3250.670 ;
        RECT -9.070 3071.090 -7.890 3072.270 ;
        RECT -9.070 3069.490 -7.890 3070.670 ;
        RECT -9.070 2891.090 -7.890 2892.270 ;
        RECT -9.070 2889.490 -7.890 2890.670 ;
        RECT -9.070 2711.090 -7.890 2712.270 ;
        RECT -9.070 2709.490 -7.890 2710.670 ;
        RECT -9.070 2531.090 -7.890 2532.270 ;
        RECT -9.070 2529.490 -7.890 2530.670 ;
        RECT -9.070 2351.090 -7.890 2352.270 ;
        RECT -9.070 2349.490 -7.890 2350.670 ;
        RECT -9.070 2171.090 -7.890 2172.270 ;
        RECT -9.070 2169.490 -7.890 2170.670 ;
        RECT -9.070 1991.090 -7.890 1992.270 ;
        RECT -9.070 1989.490 -7.890 1990.670 ;
        RECT -9.070 1811.090 -7.890 1812.270 ;
        RECT -9.070 1809.490 -7.890 1810.670 ;
        RECT -9.070 1631.090 -7.890 1632.270 ;
        RECT -9.070 1629.490 -7.890 1630.670 ;
        RECT -9.070 1451.090 -7.890 1452.270 ;
        RECT -9.070 1449.490 -7.890 1450.670 ;
        RECT -9.070 1271.090 -7.890 1272.270 ;
        RECT -9.070 1269.490 -7.890 1270.670 ;
        RECT -9.070 1091.090 -7.890 1092.270 ;
        RECT -9.070 1089.490 -7.890 1090.670 ;
        RECT -9.070 911.090 -7.890 912.270 ;
        RECT -9.070 909.490 -7.890 910.670 ;
        RECT -9.070 731.090 -7.890 732.270 ;
        RECT -9.070 729.490 -7.890 730.670 ;
        RECT -9.070 551.090 -7.890 552.270 ;
        RECT -9.070 549.490 -7.890 550.670 ;
        RECT -9.070 371.090 -7.890 372.270 ;
        RECT -9.070 369.490 -7.890 370.670 ;
        RECT -9.070 191.090 -7.890 192.270 ;
        RECT -9.070 189.490 -7.890 190.670 ;
        RECT -9.070 11.090 -7.890 12.270 ;
        RECT -9.070 9.490 -7.890 10.670 ;
        RECT -9.070 -2.910 -7.890 -1.730 ;
        RECT -9.070 -4.510 -7.890 -3.330 ;
        RECT 4.930 3523.010 6.110 3524.190 ;
        RECT 4.930 3521.410 6.110 3522.590 ;
        RECT 4.930 3431.090 6.110 3432.270 ;
        RECT 4.930 3429.490 6.110 3430.670 ;
        RECT 4.930 3251.090 6.110 3252.270 ;
        RECT 4.930 3249.490 6.110 3250.670 ;
        RECT 4.930 3071.090 6.110 3072.270 ;
        RECT 4.930 3069.490 6.110 3070.670 ;
        RECT 4.930 2891.090 6.110 2892.270 ;
        RECT 4.930 2889.490 6.110 2890.670 ;
        RECT 4.930 2711.090 6.110 2712.270 ;
        RECT 4.930 2709.490 6.110 2710.670 ;
        RECT 4.930 2531.090 6.110 2532.270 ;
        RECT 4.930 2529.490 6.110 2530.670 ;
        RECT 4.930 2351.090 6.110 2352.270 ;
        RECT 4.930 2349.490 6.110 2350.670 ;
        RECT 4.930 2171.090 6.110 2172.270 ;
        RECT 4.930 2169.490 6.110 2170.670 ;
        RECT 4.930 1991.090 6.110 1992.270 ;
        RECT 4.930 1989.490 6.110 1990.670 ;
        RECT 4.930 1811.090 6.110 1812.270 ;
        RECT 4.930 1809.490 6.110 1810.670 ;
        RECT 4.930 1631.090 6.110 1632.270 ;
        RECT 4.930 1629.490 6.110 1630.670 ;
        RECT 4.930 1451.090 6.110 1452.270 ;
        RECT 4.930 1449.490 6.110 1450.670 ;
        RECT 4.930 1271.090 6.110 1272.270 ;
        RECT 4.930 1269.490 6.110 1270.670 ;
        RECT 4.930 1091.090 6.110 1092.270 ;
        RECT 4.930 1089.490 6.110 1090.670 ;
        RECT 4.930 911.090 6.110 912.270 ;
        RECT 4.930 909.490 6.110 910.670 ;
        RECT 4.930 731.090 6.110 732.270 ;
        RECT 4.930 729.490 6.110 730.670 ;
        RECT 4.930 551.090 6.110 552.270 ;
        RECT 4.930 549.490 6.110 550.670 ;
        RECT 4.930 371.090 6.110 372.270 ;
        RECT 4.930 369.490 6.110 370.670 ;
        RECT 4.930 191.090 6.110 192.270 ;
        RECT 4.930 189.490 6.110 190.670 ;
        RECT 4.930 11.090 6.110 12.270 ;
        RECT 4.930 9.490 6.110 10.670 ;
        RECT 4.930 -2.910 6.110 -1.730 ;
        RECT 4.930 -4.510 6.110 -3.330 ;
        RECT 22.930 3449.090 24.110 3450.270 ;
        RECT 22.930 3447.490 24.110 3448.670 ;
        RECT 22.930 3269.090 24.110 3270.270 ;
        RECT 22.930 3267.490 24.110 3268.670 ;
        RECT 22.930 3089.090 24.110 3090.270 ;
        RECT 22.930 3087.490 24.110 3088.670 ;
        RECT 22.930 2909.090 24.110 2910.270 ;
        RECT 22.930 2907.490 24.110 2908.670 ;
        RECT 22.930 2729.090 24.110 2730.270 ;
        RECT 22.930 2727.490 24.110 2728.670 ;
        RECT 22.930 2549.090 24.110 2550.270 ;
        RECT 22.930 2547.490 24.110 2548.670 ;
        RECT 22.930 2369.090 24.110 2370.270 ;
        RECT 22.930 2367.490 24.110 2368.670 ;
        RECT 22.930 2189.090 24.110 2190.270 ;
        RECT 22.930 2187.490 24.110 2188.670 ;
        RECT 22.930 2009.090 24.110 2010.270 ;
        RECT 22.930 2007.490 24.110 2008.670 ;
        RECT 22.930 1829.090 24.110 1830.270 ;
        RECT 22.930 1827.490 24.110 1828.670 ;
        RECT 22.930 1649.090 24.110 1650.270 ;
        RECT 22.930 1647.490 24.110 1648.670 ;
        RECT 22.930 1469.090 24.110 1470.270 ;
        RECT 22.930 1467.490 24.110 1468.670 ;
        RECT 22.930 1289.090 24.110 1290.270 ;
        RECT 22.930 1287.490 24.110 1288.670 ;
        RECT 22.930 1109.090 24.110 1110.270 ;
        RECT 22.930 1107.490 24.110 1108.670 ;
        RECT 22.930 929.090 24.110 930.270 ;
        RECT 22.930 927.490 24.110 928.670 ;
        RECT 22.930 749.090 24.110 750.270 ;
        RECT 22.930 747.490 24.110 748.670 ;
        RECT 22.930 569.090 24.110 570.270 ;
        RECT 22.930 567.490 24.110 568.670 ;
        RECT 22.930 389.090 24.110 390.270 ;
        RECT 22.930 387.490 24.110 388.670 ;
        RECT 22.930 209.090 24.110 210.270 ;
        RECT 22.930 207.490 24.110 208.670 ;
        RECT 22.930 29.090 24.110 30.270 ;
        RECT 22.930 27.490 24.110 28.670 ;
        RECT -18.470 -12.310 -17.290 -11.130 ;
        RECT -18.470 -13.910 -17.290 -12.730 ;
        RECT 22.930 -12.310 24.110 -11.130 ;
        RECT 22.930 -13.910 24.110 -12.730 ;
        RECT 40.930 3467.090 42.110 3468.270 ;
        RECT 40.930 3465.490 42.110 3466.670 ;
        RECT 40.930 3287.090 42.110 3288.270 ;
        RECT 40.930 3285.490 42.110 3286.670 ;
        RECT 40.930 3107.090 42.110 3108.270 ;
        RECT 40.930 3105.490 42.110 3106.670 ;
        RECT 40.930 2927.090 42.110 2928.270 ;
        RECT 40.930 2925.490 42.110 2926.670 ;
        RECT 40.930 2747.090 42.110 2748.270 ;
        RECT 40.930 2745.490 42.110 2746.670 ;
        RECT 40.930 2567.090 42.110 2568.270 ;
        RECT 40.930 2565.490 42.110 2566.670 ;
        RECT 40.930 2387.090 42.110 2388.270 ;
        RECT 40.930 2385.490 42.110 2386.670 ;
        RECT 40.930 2207.090 42.110 2208.270 ;
        RECT 40.930 2205.490 42.110 2206.670 ;
        RECT 40.930 2027.090 42.110 2028.270 ;
        RECT 40.930 2025.490 42.110 2026.670 ;
        RECT 40.930 1847.090 42.110 1848.270 ;
        RECT 40.930 1845.490 42.110 1846.670 ;
        RECT 40.930 1667.090 42.110 1668.270 ;
        RECT 40.930 1665.490 42.110 1666.670 ;
        RECT 40.930 1487.090 42.110 1488.270 ;
        RECT 40.930 1485.490 42.110 1486.670 ;
        RECT 40.930 1307.090 42.110 1308.270 ;
        RECT 40.930 1305.490 42.110 1306.670 ;
        RECT 40.930 1127.090 42.110 1128.270 ;
        RECT 40.930 1125.490 42.110 1126.670 ;
        RECT 40.930 947.090 42.110 948.270 ;
        RECT 40.930 945.490 42.110 946.670 ;
        RECT 40.930 767.090 42.110 768.270 ;
        RECT 40.930 765.490 42.110 766.670 ;
        RECT 40.930 587.090 42.110 588.270 ;
        RECT 40.930 585.490 42.110 586.670 ;
        RECT 40.930 407.090 42.110 408.270 ;
        RECT 40.930 405.490 42.110 406.670 ;
        RECT 40.930 227.090 42.110 228.270 ;
        RECT 40.930 225.490 42.110 226.670 ;
        RECT 40.930 47.090 42.110 48.270 ;
        RECT 40.930 45.490 42.110 46.670 ;
        RECT -27.870 -21.710 -26.690 -20.530 ;
        RECT -27.870 -23.310 -26.690 -22.130 ;
        RECT 40.930 -21.710 42.110 -20.530 ;
        RECT 40.930 -23.310 42.110 -22.130 ;
        RECT 238.930 3551.210 240.110 3552.390 ;
        RECT 238.930 3549.610 240.110 3550.790 ;
        RECT 220.930 3541.810 222.110 3542.990 ;
        RECT 220.930 3540.210 222.110 3541.390 ;
        RECT 202.930 3532.410 204.110 3533.590 ;
        RECT 202.930 3530.810 204.110 3531.990 ;
        RECT 58.930 3485.090 60.110 3486.270 ;
        RECT 58.930 3483.490 60.110 3484.670 ;
        RECT 58.930 3305.090 60.110 3306.270 ;
        RECT 58.930 3303.490 60.110 3304.670 ;
        RECT 58.930 3125.090 60.110 3126.270 ;
        RECT 58.930 3123.490 60.110 3124.670 ;
        RECT 58.930 2945.090 60.110 2946.270 ;
        RECT 58.930 2943.490 60.110 2944.670 ;
        RECT 58.930 2765.090 60.110 2766.270 ;
        RECT 58.930 2763.490 60.110 2764.670 ;
        RECT 58.930 2585.090 60.110 2586.270 ;
        RECT 58.930 2583.490 60.110 2584.670 ;
        RECT 58.930 2405.090 60.110 2406.270 ;
        RECT 58.930 2403.490 60.110 2404.670 ;
        RECT 58.930 2225.090 60.110 2226.270 ;
        RECT 58.930 2223.490 60.110 2224.670 ;
        RECT 58.930 2045.090 60.110 2046.270 ;
        RECT 58.930 2043.490 60.110 2044.670 ;
        RECT 58.930 1865.090 60.110 1866.270 ;
        RECT 58.930 1863.490 60.110 1864.670 ;
        RECT 58.930 1685.090 60.110 1686.270 ;
        RECT 58.930 1683.490 60.110 1684.670 ;
        RECT 58.930 1505.090 60.110 1506.270 ;
        RECT 58.930 1503.490 60.110 1504.670 ;
        RECT 58.930 1325.090 60.110 1326.270 ;
        RECT 58.930 1323.490 60.110 1324.670 ;
        RECT 58.930 1145.090 60.110 1146.270 ;
        RECT 58.930 1143.490 60.110 1144.670 ;
        RECT 58.930 965.090 60.110 966.270 ;
        RECT 58.930 963.490 60.110 964.670 ;
        RECT 58.930 785.090 60.110 786.270 ;
        RECT 58.930 783.490 60.110 784.670 ;
        RECT 58.930 605.090 60.110 606.270 ;
        RECT 58.930 603.490 60.110 604.670 ;
        RECT 58.930 425.090 60.110 426.270 ;
        RECT 58.930 423.490 60.110 424.670 ;
        RECT 58.930 245.090 60.110 246.270 ;
        RECT 58.930 243.490 60.110 244.670 ;
        RECT 58.930 65.090 60.110 66.270 ;
        RECT 58.930 63.490 60.110 64.670 ;
        RECT -37.270 -31.110 -36.090 -29.930 ;
        RECT -37.270 -32.710 -36.090 -31.530 ;
        RECT 184.930 3523.010 186.110 3524.190 ;
        RECT 184.930 3521.410 186.110 3522.590 ;
        RECT 184.930 3431.090 186.110 3432.270 ;
        RECT 184.930 3429.490 186.110 3430.670 ;
        RECT 184.930 3251.090 186.110 3252.270 ;
        RECT 184.930 3249.490 186.110 3250.670 ;
        RECT 184.930 3071.090 186.110 3072.270 ;
        RECT 184.930 3069.490 186.110 3070.670 ;
        RECT 184.930 2891.090 186.110 2892.270 ;
        RECT 184.930 2889.490 186.110 2890.670 ;
        RECT 184.930 2711.090 186.110 2712.270 ;
        RECT 184.930 2709.490 186.110 2710.670 ;
        RECT 184.930 2531.090 186.110 2532.270 ;
        RECT 184.930 2529.490 186.110 2530.670 ;
        RECT 184.930 2351.090 186.110 2352.270 ;
        RECT 184.930 2349.490 186.110 2350.670 ;
        RECT 184.930 2171.090 186.110 2172.270 ;
        RECT 184.930 2169.490 186.110 2170.670 ;
        RECT 184.930 1991.090 186.110 1992.270 ;
        RECT 184.930 1989.490 186.110 1990.670 ;
        RECT 184.930 1811.090 186.110 1812.270 ;
        RECT 184.930 1809.490 186.110 1810.670 ;
        RECT 184.930 1631.090 186.110 1632.270 ;
        RECT 184.930 1629.490 186.110 1630.670 ;
        RECT 184.930 1451.090 186.110 1452.270 ;
        RECT 184.930 1449.490 186.110 1450.670 ;
        RECT 184.930 1271.090 186.110 1272.270 ;
        RECT 184.930 1269.490 186.110 1270.670 ;
        RECT 184.930 1091.090 186.110 1092.270 ;
        RECT 184.930 1089.490 186.110 1090.670 ;
        RECT 184.930 911.090 186.110 912.270 ;
        RECT 184.930 909.490 186.110 910.670 ;
        RECT 184.930 731.090 186.110 732.270 ;
        RECT 184.930 729.490 186.110 730.670 ;
        RECT 184.930 551.090 186.110 552.270 ;
        RECT 184.930 549.490 186.110 550.670 ;
        RECT 184.930 371.090 186.110 372.270 ;
        RECT 184.930 369.490 186.110 370.670 ;
        RECT 184.930 191.090 186.110 192.270 ;
        RECT 184.930 189.490 186.110 190.670 ;
        RECT 184.930 11.090 186.110 12.270 ;
        RECT 184.930 9.490 186.110 10.670 ;
        RECT 184.930 -2.910 186.110 -1.730 ;
        RECT 184.930 -4.510 186.110 -3.330 ;
        RECT 202.930 3449.090 204.110 3450.270 ;
        RECT 202.930 3447.490 204.110 3448.670 ;
        RECT 202.930 3269.090 204.110 3270.270 ;
        RECT 202.930 3267.490 204.110 3268.670 ;
        RECT 202.930 3089.090 204.110 3090.270 ;
        RECT 202.930 3087.490 204.110 3088.670 ;
        RECT 202.930 2909.090 204.110 2910.270 ;
        RECT 202.930 2907.490 204.110 2908.670 ;
        RECT 202.930 2729.090 204.110 2730.270 ;
        RECT 202.930 2727.490 204.110 2728.670 ;
        RECT 202.930 2549.090 204.110 2550.270 ;
        RECT 202.930 2547.490 204.110 2548.670 ;
        RECT 202.930 2369.090 204.110 2370.270 ;
        RECT 202.930 2367.490 204.110 2368.670 ;
        RECT 202.930 2189.090 204.110 2190.270 ;
        RECT 202.930 2187.490 204.110 2188.670 ;
        RECT 202.930 2009.090 204.110 2010.270 ;
        RECT 202.930 2007.490 204.110 2008.670 ;
        RECT 202.930 1829.090 204.110 1830.270 ;
        RECT 202.930 1827.490 204.110 1828.670 ;
        RECT 202.930 1649.090 204.110 1650.270 ;
        RECT 202.930 1647.490 204.110 1648.670 ;
        RECT 202.930 1469.090 204.110 1470.270 ;
        RECT 202.930 1467.490 204.110 1468.670 ;
        RECT 202.930 1289.090 204.110 1290.270 ;
        RECT 202.930 1287.490 204.110 1288.670 ;
        RECT 202.930 1109.090 204.110 1110.270 ;
        RECT 202.930 1107.490 204.110 1108.670 ;
        RECT 202.930 929.090 204.110 930.270 ;
        RECT 202.930 927.490 204.110 928.670 ;
        RECT 202.930 749.090 204.110 750.270 ;
        RECT 202.930 747.490 204.110 748.670 ;
        RECT 202.930 569.090 204.110 570.270 ;
        RECT 202.930 567.490 204.110 568.670 ;
        RECT 202.930 389.090 204.110 390.270 ;
        RECT 202.930 387.490 204.110 388.670 ;
        RECT 202.930 209.090 204.110 210.270 ;
        RECT 202.930 207.490 204.110 208.670 ;
        RECT 202.930 29.090 204.110 30.270 ;
        RECT 202.930 27.490 204.110 28.670 ;
        RECT 202.930 -12.310 204.110 -11.130 ;
        RECT 202.930 -13.910 204.110 -12.730 ;
        RECT 220.930 3467.090 222.110 3468.270 ;
        RECT 220.930 3465.490 222.110 3466.670 ;
        RECT 220.930 3287.090 222.110 3288.270 ;
        RECT 220.930 3285.490 222.110 3286.670 ;
        RECT 220.930 3107.090 222.110 3108.270 ;
        RECT 220.930 3105.490 222.110 3106.670 ;
        RECT 220.930 2927.090 222.110 2928.270 ;
        RECT 220.930 2925.490 222.110 2926.670 ;
        RECT 220.930 2747.090 222.110 2748.270 ;
        RECT 220.930 2745.490 222.110 2746.670 ;
        RECT 220.930 2567.090 222.110 2568.270 ;
        RECT 220.930 2565.490 222.110 2566.670 ;
        RECT 220.930 2387.090 222.110 2388.270 ;
        RECT 220.930 2385.490 222.110 2386.670 ;
        RECT 220.930 2207.090 222.110 2208.270 ;
        RECT 220.930 2205.490 222.110 2206.670 ;
        RECT 220.930 2027.090 222.110 2028.270 ;
        RECT 220.930 2025.490 222.110 2026.670 ;
        RECT 220.930 1847.090 222.110 1848.270 ;
        RECT 220.930 1845.490 222.110 1846.670 ;
        RECT 220.930 1667.090 222.110 1668.270 ;
        RECT 220.930 1665.490 222.110 1666.670 ;
        RECT 220.930 1487.090 222.110 1488.270 ;
        RECT 220.930 1485.490 222.110 1486.670 ;
        RECT 220.930 1307.090 222.110 1308.270 ;
        RECT 220.930 1305.490 222.110 1306.670 ;
        RECT 220.930 1127.090 222.110 1128.270 ;
        RECT 220.930 1125.490 222.110 1126.670 ;
        RECT 220.930 947.090 222.110 948.270 ;
        RECT 220.930 945.490 222.110 946.670 ;
        RECT 220.930 767.090 222.110 768.270 ;
        RECT 220.930 765.490 222.110 766.670 ;
        RECT 220.930 587.090 222.110 588.270 ;
        RECT 220.930 585.490 222.110 586.670 ;
        RECT 220.930 407.090 222.110 408.270 ;
        RECT 220.930 405.490 222.110 406.670 ;
        RECT 220.930 227.090 222.110 228.270 ;
        RECT 220.930 225.490 222.110 226.670 ;
        RECT 220.930 47.090 222.110 48.270 ;
        RECT 220.930 45.490 222.110 46.670 ;
        RECT 220.930 -21.710 222.110 -20.530 ;
        RECT 220.930 -23.310 222.110 -22.130 ;
        RECT 418.930 3551.210 420.110 3552.390 ;
        RECT 418.930 3549.610 420.110 3550.790 ;
        RECT 400.930 3541.810 402.110 3542.990 ;
        RECT 400.930 3540.210 402.110 3541.390 ;
        RECT 382.930 3532.410 384.110 3533.590 ;
        RECT 382.930 3530.810 384.110 3531.990 ;
        RECT 238.930 3485.090 240.110 3486.270 ;
        RECT 238.930 3483.490 240.110 3484.670 ;
        RECT 238.930 3305.090 240.110 3306.270 ;
        RECT 238.930 3303.490 240.110 3304.670 ;
        RECT 364.930 3523.010 366.110 3524.190 ;
        RECT 364.930 3521.410 366.110 3522.590 ;
        RECT 364.930 3431.090 366.110 3432.270 ;
        RECT 364.930 3429.490 366.110 3430.670 ;
        RECT 382.930 3449.090 384.110 3450.270 ;
        RECT 382.930 3447.490 384.110 3448.670 ;
        RECT 400.930 3467.090 402.110 3468.270 ;
        RECT 400.930 3465.490 402.110 3466.670 ;
        RECT 400.930 3287.090 402.110 3288.270 ;
        RECT 400.930 3285.490 402.110 3286.670 ;
        RECT 598.930 3551.210 600.110 3552.390 ;
        RECT 598.930 3549.610 600.110 3550.790 ;
        RECT 580.930 3541.810 582.110 3542.990 ;
        RECT 580.930 3540.210 582.110 3541.390 ;
        RECT 562.930 3532.410 564.110 3533.590 ;
        RECT 562.930 3530.810 564.110 3531.990 ;
        RECT 418.930 3485.090 420.110 3486.270 ;
        RECT 418.930 3483.490 420.110 3484.670 ;
        RECT 418.930 3305.090 420.110 3306.270 ;
        RECT 418.930 3303.490 420.110 3304.670 ;
        RECT 544.930 3523.010 546.110 3524.190 ;
        RECT 544.930 3521.410 546.110 3522.590 ;
        RECT 544.930 3431.090 546.110 3432.270 ;
        RECT 544.930 3429.490 546.110 3430.670 ;
        RECT 562.930 3449.090 564.110 3450.270 ;
        RECT 562.930 3447.490 564.110 3448.670 ;
        RECT 580.930 3467.090 582.110 3468.270 ;
        RECT 580.930 3465.490 582.110 3466.670 ;
        RECT 580.930 3287.090 582.110 3288.270 ;
        RECT 580.930 3285.490 582.110 3286.670 ;
        RECT 778.930 3551.210 780.110 3552.390 ;
        RECT 778.930 3549.610 780.110 3550.790 ;
        RECT 760.930 3541.810 762.110 3542.990 ;
        RECT 760.930 3540.210 762.110 3541.390 ;
        RECT 742.930 3532.410 744.110 3533.590 ;
        RECT 742.930 3530.810 744.110 3531.990 ;
        RECT 598.930 3485.090 600.110 3486.270 ;
        RECT 598.930 3483.490 600.110 3484.670 ;
        RECT 598.930 3305.090 600.110 3306.270 ;
        RECT 598.930 3303.490 600.110 3304.670 ;
        RECT 724.930 3523.010 726.110 3524.190 ;
        RECT 724.930 3521.410 726.110 3522.590 ;
        RECT 724.930 3431.090 726.110 3432.270 ;
        RECT 724.930 3429.490 726.110 3430.670 ;
        RECT 724.930 3251.090 726.110 3252.270 ;
        RECT 724.930 3249.490 726.110 3250.670 ;
        RECT 238.930 3125.090 240.110 3126.270 ;
        RECT 238.930 3123.490 240.110 3124.670 ;
        RECT 238.930 2945.090 240.110 2946.270 ;
        RECT 238.930 2943.490 240.110 2944.670 ;
        RECT 682.680 3125.090 683.860 3126.270 ;
        RECT 682.680 3123.490 683.860 3124.670 ;
        RECT 682.680 3107.090 683.860 3108.270 ;
        RECT 682.680 3105.490 683.860 3106.670 ;
        RECT 682.680 3089.090 683.860 3090.270 ;
        RECT 682.680 3087.490 683.860 3088.670 ;
        RECT 682.680 3071.090 683.860 3072.270 ;
        RECT 682.680 3069.490 683.860 3070.670 ;
        RECT 682.680 2945.090 683.860 2946.270 ;
        RECT 682.680 2943.490 683.860 2944.670 ;
        RECT 682.680 2927.090 683.860 2928.270 ;
        RECT 682.680 2925.490 683.860 2926.670 ;
        RECT 682.680 2909.090 683.860 2910.270 ;
        RECT 682.680 2907.490 683.860 2908.670 ;
        RECT 682.680 2891.090 683.860 2892.270 ;
        RECT 682.680 2889.490 683.860 2890.670 ;
        RECT 724.930 3071.090 726.110 3072.270 ;
        RECT 724.930 3069.490 726.110 3070.670 ;
        RECT 724.930 2891.090 726.110 2892.270 ;
        RECT 724.930 2889.490 726.110 2890.670 ;
        RECT 238.930 2765.090 240.110 2766.270 ;
        RECT 238.930 2763.490 240.110 2764.670 ;
        RECT 382.930 2729.090 384.110 2730.270 ;
        RECT 382.930 2727.490 384.110 2728.670 ;
        RECT 400.930 2747.090 402.110 2748.270 ;
        RECT 400.930 2745.490 402.110 2746.670 ;
        RECT 418.930 2765.090 420.110 2766.270 ;
        RECT 418.930 2763.490 420.110 2764.670 ;
        RECT 562.930 2729.090 564.110 2730.270 ;
        RECT 562.930 2727.490 564.110 2728.670 ;
        RECT 580.930 2747.090 582.110 2748.270 ;
        RECT 580.930 2745.490 582.110 2746.670 ;
        RECT 598.930 2765.090 600.110 2766.270 ;
        RECT 598.930 2763.490 600.110 2764.670 ;
        RECT 742.930 3449.090 744.110 3450.270 ;
        RECT 742.930 3447.490 744.110 3448.670 ;
        RECT 742.930 3269.090 744.110 3270.270 ;
        RECT 742.930 3267.490 744.110 3268.670 ;
        RECT 742.930 3089.090 744.110 3090.270 ;
        RECT 742.930 3087.490 744.110 3088.670 ;
        RECT 742.930 2909.090 744.110 2910.270 ;
        RECT 742.930 2907.490 744.110 2908.670 ;
        RECT 742.930 2729.090 744.110 2730.270 ;
        RECT 742.930 2727.490 744.110 2728.670 ;
        RECT 760.930 3467.090 762.110 3468.270 ;
        RECT 760.930 3465.490 762.110 3466.670 ;
        RECT 760.930 3287.090 762.110 3288.270 ;
        RECT 760.930 3285.490 762.110 3286.670 ;
        RECT 760.930 3107.090 762.110 3108.270 ;
        RECT 760.930 3105.490 762.110 3106.670 ;
        RECT 760.930 2927.090 762.110 2928.270 ;
        RECT 760.930 2925.490 762.110 2926.670 ;
        RECT 760.930 2747.090 762.110 2748.270 ;
        RECT 760.930 2745.490 762.110 2746.670 ;
        RECT 958.930 3551.210 960.110 3552.390 ;
        RECT 958.930 3549.610 960.110 3550.790 ;
        RECT 940.930 3541.810 942.110 3542.990 ;
        RECT 940.930 3540.210 942.110 3541.390 ;
        RECT 922.930 3532.410 924.110 3533.590 ;
        RECT 922.930 3530.810 924.110 3531.990 ;
        RECT 778.930 3485.090 780.110 3486.270 ;
        RECT 778.930 3483.490 780.110 3484.670 ;
        RECT 778.930 3305.090 780.110 3306.270 ;
        RECT 778.930 3303.490 780.110 3304.670 ;
        RECT 778.930 3125.090 780.110 3126.270 ;
        RECT 778.930 3123.490 780.110 3124.670 ;
        RECT 778.930 2945.090 780.110 2946.270 ;
        RECT 778.930 2943.490 780.110 2944.670 ;
        RECT 778.930 2765.090 780.110 2766.270 ;
        RECT 778.930 2763.490 780.110 2764.670 ;
        RECT 904.930 3523.010 906.110 3524.190 ;
        RECT 904.930 3521.410 906.110 3522.590 ;
        RECT 904.930 3431.090 906.110 3432.270 ;
        RECT 904.930 3429.490 906.110 3430.670 ;
        RECT 904.930 3251.090 906.110 3252.270 ;
        RECT 904.930 3249.490 906.110 3250.670 ;
        RECT 904.930 3071.090 906.110 3072.270 ;
        RECT 904.930 3069.490 906.110 3070.670 ;
        RECT 904.930 2891.090 906.110 2892.270 ;
        RECT 904.930 2889.490 906.110 2890.670 ;
        RECT 922.930 3449.090 924.110 3450.270 ;
        RECT 922.930 3447.490 924.110 3448.670 ;
        RECT 940.930 3467.090 942.110 3468.270 ;
        RECT 940.930 3465.490 942.110 3466.670 ;
        RECT 940.930 3287.090 942.110 3288.270 ;
        RECT 940.930 3285.490 942.110 3286.670 ;
        RECT 1138.930 3551.210 1140.110 3552.390 ;
        RECT 1138.930 3549.610 1140.110 3550.790 ;
        RECT 1120.930 3541.810 1122.110 3542.990 ;
        RECT 1120.930 3540.210 1122.110 3541.390 ;
        RECT 1102.930 3532.410 1104.110 3533.590 ;
        RECT 1102.930 3530.810 1104.110 3531.990 ;
        RECT 958.930 3485.090 960.110 3486.270 ;
        RECT 958.930 3483.490 960.110 3484.670 ;
        RECT 958.930 3305.090 960.110 3306.270 ;
        RECT 958.930 3303.490 960.110 3304.670 ;
        RECT 1084.930 3523.010 1086.110 3524.190 ;
        RECT 1084.930 3521.410 1086.110 3522.590 ;
        RECT 1084.930 3431.090 1086.110 3432.270 ;
        RECT 1084.930 3429.490 1086.110 3430.670 ;
        RECT 1102.930 3449.090 1104.110 3450.270 ;
        RECT 1102.930 3447.490 1104.110 3448.670 ;
        RECT 1120.930 3467.090 1122.110 3468.270 ;
        RECT 1120.930 3465.490 1122.110 3466.670 ;
        RECT 1120.930 3287.090 1122.110 3288.270 ;
        RECT 1120.930 3285.490 1122.110 3286.670 ;
        RECT 1318.930 3551.210 1320.110 3552.390 ;
        RECT 1318.930 3549.610 1320.110 3550.790 ;
        RECT 1300.930 3541.810 1302.110 3542.990 ;
        RECT 1300.930 3540.210 1302.110 3541.390 ;
        RECT 1282.930 3532.410 1284.110 3533.590 ;
        RECT 1282.930 3530.810 1284.110 3531.990 ;
        RECT 1138.930 3485.090 1140.110 3486.270 ;
        RECT 1138.930 3483.490 1140.110 3484.670 ;
        RECT 1138.930 3305.090 1140.110 3306.270 ;
        RECT 1138.930 3303.490 1140.110 3304.670 ;
        RECT 1264.930 3523.010 1266.110 3524.190 ;
        RECT 1264.930 3521.410 1266.110 3522.590 ;
        RECT 1264.930 3431.090 1266.110 3432.270 ;
        RECT 1264.930 3429.490 1266.110 3430.670 ;
        RECT 1282.930 3449.090 1284.110 3450.270 ;
        RECT 1282.930 3447.490 1284.110 3448.670 ;
        RECT 1300.930 3467.090 1302.110 3468.270 ;
        RECT 1300.930 3465.490 1302.110 3466.670 ;
        RECT 1300.930 3287.090 1302.110 3288.270 ;
        RECT 1300.930 3285.490 1302.110 3286.670 ;
        RECT 1498.930 3551.210 1500.110 3552.390 ;
        RECT 1498.930 3549.610 1500.110 3550.790 ;
        RECT 1480.930 3541.810 1482.110 3542.990 ;
        RECT 1480.930 3540.210 1482.110 3541.390 ;
        RECT 1462.930 3532.410 1464.110 3533.590 ;
        RECT 1462.930 3530.810 1464.110 3531.990 ;
        RECT 1318.930 3485.090 1320.110 3486.270 ;
        RECT 1318.930 3483.490 1320.110 3484.670 ;
        RECT 1318.930 3305.090 1320.110 3306.270 ;
        RECT 1318.930 3303.490 1320.110 3304.670 ;
        RECT 1444.930 3523.010 1446.110 3524.190 ;
        RECT 1444.930 3521.410 1446.110 3522.590 ;
        RECT 1444.930 3431.090 1446.110 3432.270 ;
        RECT 1444.930 3429.490 1446.110 3430.670 ;
        RECT 922.930 3269.090 924.110 3270.270 ;
        RECT 922.930 3267.490 924.110 3268.670 ;
        RECT 1444.930 3251.090 1446.110 3252.270 ;
        RECT 1444.930 3249.490 1446.110 3250.670 ;
        RECT 922.930 3089.090 924.110 3090.270 ;
        RECT 922.930 3087.490 924.110 3088.670 ;
        RECT 922.930 2909.090 924.110 2910.270 ;
        RECT 922.930 2907.490 924.110 2908.670 ;
        RECT 1332.680 3125.090 1333.860 3126.270 ;
        RECT 1332.680 3123.490 1333.860 3124.670 ;
        RECT 1332.680 3107.090 1333.860 3108.270 ;
        RECT 1332.680 3105.490 1333.860 3106.670 ;
        RECT 1332.680 3089.090 1333.860 3090.270 ;
        RECT 1332.680 3087.490 1333.860 3088.670 ;
        RECT 1332.680 3071.090 1333.860 3072.270 ;
        RECT 1332.680 3069.490 1333.860 3070.670 ;
        RECT 1332.680 2945.090 1333.860 2946.270 ;
        RECT 1332.680 2943.490 1333.860 2944.670 ;
        RECT 1332.680 2927.090 1333.860 2928.270 ;
        RECT 1332.680 2925.490 1333.860 2926.670 ;
        RECT 1332.680 2909.090 1333.860 2910.270 ;
        RECT 1332.680 2907.490 1333.860 2908.670 ;
        RECT 1332.680 2891.090 1333.860 2892.270 ;
        RECT 1332.680 2889.490 1333.860 2890.670 ;
        RECT 1444.930 3071.090 1446.110 3072.270 ;
        RECT 1444.930 3069.490 1446.110 3070.670 ;
        RECT 1444.930 2891.090 1446.110 2892.270 ;
        RECT 1444.930 2889.490 1446.110 2890.670 ;
        RECT 922.930 2729.090 924.110 2730.270 ;
        RECT 922.930 2727.490 924.110 2728.670 ;
        RECT 940.930 2747.090 942.110 2748.270 ;
        RECT 940.930 2745.490 942.110 2746.670 ;
        RECT 958.930 2765.090 960.110 2766.270 ;
        RECT 958.930 2763.490 960.110 2764.670 ;
        RECT 1102.930 2729.090 1104.110 2730.270 ;
        RECT 1102.930 2727.490 1104.110 2728.670 ;
        RECT 1120.930 2747.090 1122.110 2748.270 ;
        RECT 1120.930 2745.490 1122.110 2746.670 ;
        RECT 1138.930 2765.090 1140.110 2766.270 ;
        RECT 1138.930 2763.490 1140.110 2764.670 ;
        RECT 1282.930 2729.090 1284.110 2730.270 ;
        RECT 1282.930 2727.490 1284.110 2728.670 ;
        RECT 1300.930 2747.090 1302.110 2748.270 ;
        RECT 1300.930 2745.490 1302.110 2746.670 ;
        RECT 1318.930 2765.090 1320.110 2766.270 ;
        RECT 1318.930 2763.490 1320.110 2764.670 ;
        RECT 1444.930 2711.090 1446.110 2712.270 ;
        RECT 1444.930 2709.490 1446.110 2710.670 ;
        RECT 238.930 2585.090 240.110 2586.270 ;
        RECT 238.930 2583.490 240.110 2584.670 ;
        RECT 238.930 2405.090 240.110 2406.270 ;
        RECT 238.930 2403.490 240.110 2404.670 ;
        RECT 238.930 2225.090 240.110 2226.270 ;
        RECT 238.930 2223.490 240.110 2224.670 ;
        RECT 238.930 2045.090 240.110 2046.270 ;
        RECT 238.930 2043.490 240.110 2044.670 ;
        RECT 238.930 1865.090 240.110 1866.270 ;
        RECT 238.930 1863.490 240.110 1864.670 ;
        RECT 238.930 1685.090 240.110 1686.270 ;
        RECT 238.930 1683.490 240.110 1684.670 ;
        RECT 321.250 2585.090 322.430 2586.270 ;
        RECT 321.250 2583.490 322.430 2584.670 ;
        RECT 321.250 2567.090 322.430 2568.270 ;
        RECT 321.250 2565.490 322.430 2566.670 ;
        RECT 321.250 2549.090 322.430 2550.270 ;
        RECT 321.250 2547.490 322.430 2548.670 ;
        RECT 321.250 2531.090 322.430 2532.270 ;
        RECT 321.250 2529.490 322.430 2530.670 ;
        RECT 321.250 2405.090 322.430 2406.270 ;
        RECT 321.250 2403.490 322.430 2404.670 ;
        RECT 321.250 2387.090 322.430 2388.270 ;
        RECT 321.250 2385.490 322.430 2386.670 ;
        RECT 321.250 2369.090 322.430 2370.270 ;
        RECT 321.250 2367.490 322.430 2368.670 ;
        RECT 321.250 2351.090 322.430 2352.270 ;
        RECT 321.250 2349.490 322.430 2350.670 ;
        RECT 321.250 2225.090 322.430 2226.270 ;
        RECT 321.250 2223.490 322.430 2224.670 ;
        RECT 321.250 2207.090 322.430 2208.270 ;
        RECT 321.250 2205.490 322.430 2206.670 ;
        RECT 321.250 2189.090 322.430 2190.270 ;
        RECT 321.250 2187.490 322.430 2188.670 ;
        RECT 321.250 2171.090 322.430 2172.270 ;
        RECT 321.250 2169.490 322.430 2170.670 ;
        RECT 321.250 2045.090 322.430 2046.270 ;
        RECT 321.250 2043.490 322.430 2044.670 ;
        RECT 321.250 2027.090 322.430 2028.270 ;
        RECT 321.250 2025.490 322.430 2026.670 ;
        RECT 321.250 2009.090 322.430 2010.270 ;
        RECT 321.250 2007.490 322.430 2008.670 ;
        RECT 321.250 1991.090 322.430 1992.270 ;
        RECT 321.250 1989.490 322.430 1990.670 ;
        RECT 321.250 1865.090 322.430 1866.270 ;
        RECT 321.250 1863.490 322.430 1864.670 ;
        RECT 321.250 1847.090 322.430 1848.270 ;
        RECT 321.250 1845.490 322.430 1846.670 ;
        RECT 321.250 1829.090 322.430 1830.270 ;
        RECT 321.250 1827.490 322.430 1828.670 ;
        RECT 321.250 1811.090 322.430 1812.270 ;
        RECT 321.250 1809.490 322.430 1810.670 ;
        RECT 321.250 1685.090 322.430 1686.270 ;
        RECT 321.250 1683.490 322.430 1684.670 ;
        RECT 321.250 1667.090 322.430 1668.270 ;
        RECT 321.250 1665.490 322.430 1666.670 ;
        RECT 321.250 1649.090 322.430 1650.270 ;
        RECT 321.250 1647.490 322.430 1648.670 ;
        RECT 321.250 1631.090 322.430 1632.270 ;
        RECT 321.250 1629.490 322.430 1630.670 ;
        RECT 1444.930 2531.090 1446.110 2532.270 ;
        RECT 1444.930 2529.490 1446.110 2530.670 ;
        RECT 1444.930 2351.090 1446.110 2352.270 ;
        RECT 1444.930 2349.490 1446.110 2350.670 ;
        RECT 1444.930 2171.090 1446.110 2172.270 ;
        RECT 1444.930 2169.490 1446.110 2170.670 ;
        RECT 1444.930 1991.090 1446.110 1992.270 ;
        RECT 1444.930 1989.490 1446.110 1990.670 ;
        RECT 1444.930 1811.090 1446.110 1812.270 ;
        RECT 1444.930 1809.490 1446.110 1810.670 ;
        RECT 1444.930 1631.090 1446.110 1632.270 ;
        RECT 1444.930 1629.490 1446.110 1630.670 ;
        RECT 238.930 1505.090 240.110 1506.270 ;
        RECT 238.930 1503.490 240.110 1504.670 ;
        RECT 238.930 1325.090 240.110 1326.270 ;
        RECT 238.930 1323.490 240.110 1324.670 ;
        RECT 238.930 1145.090 240.110 1146.270 ;
        RECT 238.930 1143.490 240.110 1144.670 ;
        RECT 238.930 965.090 240.110 966.270 ;
        RECT 238.930 963.490 240.110 964.670 ;
        RECT 238.930 785.090 240.110 786.270 ;
        RECT 238.930 783.490 240.110 784.670 ;
        RECT 238.930 605.090 240.110 606.270 ;
        RECT 238.930 603.490 240.110 604.670 ;
        RECT 238.930 425.090 240.110 426.270 ;
        RECT 238.930 423.490 240.110 424.670 ;
        RECT 238.930 245.090 240.110 246.270 ;
        RECT 238.930 243.490 240.110 244.670 ;
        RECT 238.930 65.090 240.110 66.270 ;
        RECT 238.930 63.490 240.110 64.670 ;
        RECT 58.930 -31.110 60.110 -29.930 ;
        RECT 58.930 -32.710 60.110 -31.530 ;
        RECT 364.930 1451.090 366.110 1452.270 ;
        RECT 364.930 1449.490 366.110 1450.670 ;
        RECT 364.930 1271.090 366.110 1272.270 ;
        RECT 364.930 1269.490 366.110 1270.670 ;
        RECT 364.930 1091.090 366.110 1092.270 ;
        RECT 364.930 1089.490 366.110 1090.670 ;
        RECT 364.930 911.090 366.110 912.270 ;
        RECT 364.930 909.490 366.110 910.670 ;
        RECT 364.930 731.090 366.110 732.270 ;
        RECT 364.930 729.490 366.110 730.670 ;
        RECT 364.930 551.090 366.110 552.270 ;
        RECT 364.930 549.490 366.110 550.670 ;
        RECT 364.930 371.090 366.110 372.270 ;
        RECT 364.930 369.490 366.110 370.670 ;
        RECT 364.930 191.090 366.110 192.270 ;
        RECT 364.930 189.490 366.110 190.670 ;
        RECT 364.930 11.090 366.110 12.270 ;
        RECT 364.930 9.490 366.110 10.670 ;
        RECT 364.930 -2.910 366.110 -1.730 ;
        RECT 364.930 -4.510 366.110 -3.330 ;
        RECT 382.930 1469.090 384.110 1470.270 ;
        RECT 382.930 1467.490 384.110 1468.670 ;
        RECT 382.930 1289.090 384.110 1290.270 ;
        RECT 382.930 1287.490 384.110 1288.670 ;
        RECT 382.930 1109.090 384.110 1110.270 ;
        RECT 382.930 1107.490 384.110 1108.670 ;
        RECT 382.930 929.090 384.110 930.270 ;
        RECT 382.930 927.490 384.110 928.670 ;
        RECT 382.930 749.090 384.110 750.270 ;
        RECT 382.930 747.490 384.110 748.670 ;
        RECT 382.930 569.090 384.110 570.270 ;
        RECT 382.930 567.490 384.110 568.670 ;
        RECT 382.930 389.090 384.110 390.270 ;
        RECT 382.930 387.490 384.110 388.670 ;
        RECT 382.930 209.090 384.110 210.270 ;
        RECT 382.930 207.490 384.110 208.670 ;
        RECT 382.930 29.090 384.110 30.270 ;
        RECT 382.930 27.490 384.110 28.670 ;
        RECT 382.930 -12.310 384.110 -11.130 ;
        RECT 382.930 -13.910 384.110 -12.730 ;
        RECT 400.930 1307.090 402.110 1308.270 ;
        RECT 400.930 1305.490 402.110 1306.670 ;
        RECT 400.930 1127.090 402.110 1128.270 ;
        RECT 400.930 1125.490 402.110 1126.670 ;
        RECT 400.930 947.090 402.110 948.270 ;
        RECT 400.930 945.490 402.110 946.670 ;
        RECT 400.930 767.090 402.110 768.270 ;
        RECT 400.930 765.490 402.110 766.670 ;
        RECT 400.930 587.090 402.110 588.270 ;
        RECT 400.930 585.490 402.110 586.670 ;
        RECT 400.930 407.090 402.110 408.270 ;
        RECT 400.930 405.490 402.110 406.670 ;
        RECT 400.930 227.090 402.110 228.270 ;
        RECT 400.930 225.490 402.110 226.670 ;
        RECT 400.930 47.090 402.110 48.270 ;
        RECT 400.930 45.490 402.110 46.670 ;
        RECT 400.930 -21.710 402.110 -20.530 ;
        RECT 400.930 -23.310 402.110 -22.130 ;
        RECT 418.930 1325.090 420.110 1326.270 ;
        RECT 418.930 1323.490 420.110 1324.670 ;
        RECT 418.930 1145.090 420.110 1146.270 ;
        RECT 418.930 1143.490 420.110 1144.670 ;
        RECT 418.930 965.090 420.110 966.270 ;
        RECT 418.930 963.490 420.110 964.670 ;
        RECT 418.930 785.090 420.110 786.270 ;
        RECT 418.930 783.490 420.110 784.670 ;
        RECT 418.930 605.090 420.110 606.270 ;
        RECT 418.930 603.490 420.110 604.670 ;
        RECT 418.930 425.090 420.110 426.270 ;
        RECT 418.930 423.490 420.110 424.670 ;
        RECT 418.930 245.090 420.110 246.270 ;
        RECT 418.930 243.490 420.110 244.670 ;
        RECT 418.930 65.090 420.110 66.270 ;
        RECT 418.930 63.490 420.110 64.670 ;
        RECT 238.930 -31.110 240.110 -29.930 ;
        RECT 238.930 -32.710 240.110 -31.530 ;
        RECT 544.930 1451.090 546.110 1452.270 ;
        RECT 544.930 1449.490 546.110 1450.670 ;
        RECT 544.930 1271.090 546.110 1272.270 ;
        RECT 544.930 1269.490 546.110 1270.670 ;
        RECT 544.930 1091.090 546.110 1092.270 ;
        RECT 544.930 1089.490 546.110 1090.670 ;
        RECT 544.930 911.090 546.110 912.270 ;
        RECT 544.930 909.490 546.110 910.670 ;
        RECT 544.930 731.090 546.110 732.270 ;
        RECT 544.930 729.490 546.110 730.670 ;
        RECT 544.930 551.090 546.110 552.270 ;
        RECT 544.930 549.490 546.110 550.670 ;
        RECT 544.930 371.090 546.110 372.270 ;
        RECT 544.930 369.490 546.110 370.670 ;
        RECT 544.930 191.090 546.110 192.270 ;
        RECT 544.930 189.490 546.110 190.670 ;
        RECT 544.930 11.090 546.110 12.270 ;
        RECT 544.930 9.490 546.110 10.670 ;
        RECT 544.930 -2.910 546.110 -1.730 ;
        RECT 544.930 -4.510 546.110 -3.330 ;
        RECT 562.930 1469.090 564.110 1470.270 ;
        RECT 562.930 1467.490 564.110 1468.670 ;
        RECT 562.930 1289.090 564.110 1290.270 ;
        RECT 562.930 1287.490 564.110 1288.670 ;
        RECT 562.930 1109.090 564.110 1110.270 ;
        RECT 562.930 1107.490 564.110 1108.670 ;
        RECT 562.930 929.090 564.110 930.270 ;
        RECT 562.930 927.490 564.110 928.670 ;
        RECT 562.930 749.090 564.110 750.270 ;
        RECT 562.930 747.490 564.110 748.670 ;
        RECT 562.930 569.090 564.110 570.270 ;
        RECT 562.930 567.490 564.110 568.670 ;
        RECT 562.930 389.090 564.110 390.270 ;
        RECT 562.930 387.490 564.110 388.670 ;
        RECT 562.930 209.090 564.110 210.270 ;
        RECT 562.930 207.490 564.110 208.670 ;
        RECT 562.930 29.090 564.110 30.270 ;
        RECT 562.930 27.490 564.110 28.670 ;
        RECT 562.930 -12.310 564.110 -11.130 ;
        RECT 562.930 -13.910 564.110 -12.730 ;
        RECT 580.930 1307.090 582.110 1308.270 ;
        RECT 580.930 1305.490 582.110 1306.670 ;
        RECT 580.930 1127.090 582.110 1128.270 ;
        RECT 580.930 1125.490 582.110 1126.670 ;
        RECT 580.930 947.090 582.110 948.270 ;
        RECT 580.930 945.490 582.110 946.670 ;
        RECT 580.930 767.090 582.110 768.270 ;
        RECT 580.930 765.490 582.110 766.670 ;
        RECT 580.930 587.090 582.110 588.270 ;
        RECT 580.930 585.490 582.110 586.670 ;
        RECT 580.930 407.090 582.110 408.270 ;
        RECT 580.930 405.490 582.110 406.670 ;
        RECT 580.930 227.090 582.110 228.270 ;
        RECT 580.930 225.490 582.110 226.670 ;
        RECT 580.930 47.090 582.110 48.270 ;
        RECT 580.930 45.490 582.110 46.670 ;
        RECT 580.930 -21.710 582.110 -20.530 ;
        RECT 580.930 -23.310 582.110 -22.130 ;
        RECT 598.930 1325.090 600.110 1326.270 ;
        RECT 598.930 1323.490 600.110 1324.670 ;
        RECT 598.930 1145.090 600.110 1146.270 ;
        RECT 598.930 1143.490 600.110 1144.670 ;
        RECT 598.930 965.090 600.110 966.270 ;
        RECT 598.930 963.490 600.110 964.670 ;
        RECT 598.930 785.090 600.110 786.270 ;
        RECT 598.930 783.490 600.110 784.670 ;
        RECT 598.930 605.090 600.110 606.270 ;
        RECT 598.930 603.490 600.110 604.670 ;
        RECT 598.930 425.090 600.110 426.270 ;
        RECT 598.930 423.490 600.110 424.670 ;
        RECT 598.930 245.090 600.110 246.270 ;
        RECT 598.930 243.490 600.110 244.670 ;
        RECT 598.930 65.090 600.110 66.270 ;
        RECT 598.930 63.490 600.110 64.670 ;
        RECT 418.930 -31.110 420.110 -29.930 ;
        RECT 418.930 -32.710 420.110 -31.530 ;
        RECT 724.930 1451.090 726.110 1452.270 ;
        RECT 724.930 1449.490 726.110 1450.670 ;
        RECT 724.930 1271.090 726.110 1272.270 ;
        RECT 724.930 1269.490 726.110 1270.670 ;
        RECT 724.930 1091.090 726.110 1092.270 ;
        RECT 724.930 1089.490 726.110 1090.670 ;
        RECT 724.930 911.090 726.110 912.270 ;
        RECT 724.930 909.490 726.110 910.670 ;
        RECT 724.930 731.090 726.110 732.270 ;
        RECT 724.930 729.490 726.110 730.670 ;
        RECT 724.930 551.090 726.110 552.270 ;
        RECT 724.930 549.490 726.110 550.670 ;
        RECT 724.930 371.090 726.110 372.270 ;
        RECT 724.930 369.490 726.110 370.670 ;
        RECT 724.930 191.090 726.110 192.270 ;
        RECT 724.930 189.490 726.110 190.670 ;
        RECT 724.930 11.090 726.110 12.270 ;
        RECT 724.930 9.490 726.110 10.670 ;
        RECT 724.930 -2.910 726.110 -1.730 ;
        RECT 724.930 -4.510 726.110 -3.330 ;
        RECT 742.930 1469.090 744.110 1470.270 ;
        RECT 742.930 1467.490 744.110 1468.670 ;
        RECT 742.930 1289.090 744.110 1290.270 ;
        RECT 742.930 1287.490 744.110 1288.670 ;
        RECT 742.930 1109.090 744.110 1110.270 ;
        RECT 742.930 1107.490 744.110 1108.670 ;
        RECT 742.930 929.090 744.110 930.270 ;
        RECT 742.930 927.490 744.110 928.670 ;
        RECT 742.930 749.090 744.110 750.270 ;
        RECT 742.930 747.490 744.110 748.670 ;
        RECT 742.930 569.090 744.110 570.270 ;
        RECT 742.930 567.490 744.110 568.670 ;
        RECT 742.930 389.090 744.110 390.270 ;
        RECT 742.930 387.490 744.110 388.670 ;
        RECT 742.930 209.090 744.110 210.270 ;
        RECT 742.930 207.490 744.110 208.670 ;
        RECT 742.930 29.090 744.110 30.270 ;
        RECT 742.930 27.490 744.110 28.670 ;
        RECT 742.930 -12.310 744.110 -11.130 ;
        RECT 742.930 -13.910 744.110 -12.730 ;
        RECT 760.930 1307.090 762.110 1308.270 ;
        RECT 760.930 1305.490 762.110 1306.670 ;
        RECT 760.930 1127.090 762.110 1128.270 ;
        RECT 760.930 1125.490 762.110 1126.670 ;
        RECT 760.930 947.090 762.110 948.270 ;
        RECT 760.930 945.490 762.110 946.670 ;
        RECT 760.930 767.090 762.110 768.270 ;
        RECT 760.930 765.490 762.110 766.670 ;
        RECT 760.930 587.090 762.110 588.270 ;
        RECT 760.930 585.490 762.110 586.670 ;
        RECT 760.930 407.090 762.110 408.270 ;
        RECT 760.930 405.490 762.110 406.670 ;
        RECT 760.930 227.090 762.110 228.270 ;
        RECT 760.930 225.490 762.110 226.670 ;
        RECT 760.930 47.090 762.110 48.270 ;
        RECT 760.930 45.490 762.110 46.670 ;
        RECT 760.930 -21.710 762.110 -20.530 ;
        RECT 760.930 -23.310 762.110 -22.130 ;
        RECT 778.930 1325.090 780.110 1326.270 ;
        RECT 778.930 1323.490 780.110 1324.670 ;
        RECT 778.930 1145.090 780.110 1146.270 ;
        RECT 778.930 1143.490 780.110 1144.670 ;
        RECT 778.930 965.090 780.110 966.270 ;
        RECT 778.930 963.490 780.110 964.670 ;
        RECT 778.930 785.090 780.110 786.270 ;
        RECT 778.930 783.490 780.110 784.670 ;
        RECT 778.930 605.090 780.110 606.270 ;
        RECT 778.930 603.490 780.110 604.670 ;
        RECT 778.930 425.090 780.110 426.270 ;
        RECT 778.930 423.490 780.110 424.670 ;
        RECT 778.930 245.090 780.110 246.270 ;
        RECT 778.930 243.490 780.110 244.670 ;
        RECT 778.930 65.090 780.110 66.270 ;
        RECT 778.930 63.490 780.110 64.670 ;
        RECT 598.930 -31.110 600.110 -29.930 ;
        RECT 598.930 -32.710 600.110 -31.530 ;
        RECT 904.930 1451.090 906.110 1452.270 ;
        RECT 904.930 1449.490 906.110 1450.670 ;
        RECT 904.930 1271.090 906.110 1272.270 ;
        RECT 904.930 1269.490 906.110 1270.670 ;
        RECT 904.930 1091.090 906.110 1092.270 ;
        RECT 904.930 1089.490 906.110 1090.670 ;
        RECT 904.930 911.090 906.110 912.270 ;
        RECT 904.930 909.490 906.110 910.670 ;
        RECT 904.930 731.090 906.110 732.270 ;
        RECT 904.930 729.490 906.110 730.670 ;
        RECT 904.930 551.090 906.110 552.270 ;
        RECT 904.930 549.490 906.110 550.670 ;
        RECT 904.930 371.090 906.110 372.270 ;
        RECT 904.930 369.490 906.110 370.670 ;
        RECT 904.930 191.090 906.110 192.270 ;
        RECT 904.930 189.490 906.110 190.670 ;
        RECT 904.930 11.090 906.110 12.270 ;
        RECT 904.930 9.490 906.110 10.670 ;
        RECT 904.930 -2.910 906.110 -1.730 ;
        RECT 904.930 -4.510 906.110 -3.330 ;
        RECT 922.930 1469.090 924.110 1470.270 ;
        RECT 922.930 1467.490 924.110 1468.670 ;
        RECT 922.930 1289.090 924.110 1290.270 ;
        RECT 922.930 1287.490 924.110 1288.670 ;
        RECT 922.930 1109.090 924.110 1110.270 ;
        RECT 922.930 1107.490 924.110 1108.670 ;
        RECT 922.930 929.090 924.110 930.270 ;
        RECT 922.930 927.490 924.110 928.670 ;
        RECT 922.930 749.090 924.110 750.270 ;
        RECT 922.930 747.490 924.110 748.670 ;
        RECT 922.930 569.090 924.110 570.270 ;
        RECT 922.930 567.490 924.110 568.670 ;
        RECT 922.930 389.090 924.110 390.270 ;
        RECT 922.930 387.490 924.110 388.670 ;
        RECT 922.930 209.090 924.110 210.270 ;
        RECT 922.930 207.490 924.110 208.670 ;
        RECT 922.930 29.090 924.110 30.270 ;
        RECT 922.930 27.490 924.110 28.670 ;
        RECT 922.930 -12.310 924.110 -11.130 ;
        RECT 922.930 -13.910 924.110 -12.730 ;
        RECT 940.930 1307.090 942.110 1308.270 ;
        RECT 940.930 1305.490 942.110 1306.670 ;
        RECT 940.930 1127.090 942.110 1128.270 ;
        RECT 940.930 1125.490 942.110 1126.670 ;
        RECT 940.930 947.090 942.110 948.270 ;
        RECT 940.930 945.490 942.110 946.670 ;
        RECT 940.930 767.090 942.110 768.270 ;
        RECT 940.930 765.490 942.110 766.670 ;
        RECT 940.930 587.090 942.110 588.270 ;
        RECT 940.930 585.490 942.110 586.670 ;
        RECT 940.930 407.090 942.110 408.270 ;
        RECT 940.930 405.490 942.110 406.670 ;
        RECT 940.930 227.090 942.110 228.270 ;
        RECT 940.930 225.490 942.110 226.670 ;
        RECT 940.930 47.090 942.110 48.270 ;
        RECT 940.930 45.490 942.110 46.670 ;
        RECT 940.930 -21.710 942.110 -20.530 ;
        RECT 940.930 -23.310 942.110 -22.130 ;
        RECT 958.930 1325.090 960.110 1326.270 ;
        RECT 958.930 1323.490 960.110 1324.670 ;
        RECT 958.930 1145.090 960.110 1146.270 ;
        RECT 958.930 1143.490 960.110 1144.670 ;
        RECT 958.930 965.090 960.110 966.270 ;
        RECT 958.930 963.490 960.110 964.670 ;
        RECT 958.930 785.090 960.110 786.270 ;
        RECT 958.930 783.490 960.110 784.670 ;
        RECT 958.930 605.090 960.110 606.270 ;
        RECT 958.930 603.490 960.110 604.670 ;
        RECT 958.930 425.090 960.110 426.270 ;
        RECT 958.930 423.490 960.110 424.670 ;
        RECT 958.930 245.090 960.110 246.270 ;
        RECT 958.930 243.490 960.110 244.670 ;
        RECT 958.930 65.090 960.110 66.270 ;
        RECT 958.930 63.490 960.110 64.670 ;
        RECT 778.930 -31.110 780.110 -29.930 ;
        RECT 778.930 -32.710 780.110 -31.530 ;
        RECT 1084.930 1451.090 1086.110 1452.270 ;
        RECT 1084.930 1449.490 1086.110 1450.670 ;
        RECT 1084.930 1271.090 1086.110 1272.270 ;
        RECT 1084.930 1269.490 1086.110 1270.670 ;
        RECT 1084.930 1091.090 1086.110 1092.270 ;
        RECT 1084.930 1089.490 1086.110 1090.670 ;
        RECT 1084.930 911.090 1086.110 912.270 ;
        RECT 1084.930 909.490 1086.110 910.670 ;
        RECT 1084.930 731.090 1086.110 732.270 ;
        RECT 1084.930 729.490 1086.110 730.670 ;
        RECT 1084.930 551.090 1086.110 552.270 ;
        RECT 1084.930 549.490 1086.110 550.670 ;
        RECT 1084.930 371.090 1086.110 372.270 ;
        RECT 1084.930 369.490 1086.110 370.670 ;
        RECT 1084.930 191.090 1086.110 192.270 ;
        RECT 1084.930 189.490 1086.110 190.670 ;
        RECT 1084.930 11.090 1086.110 12.270 ;
        RECT 1084.930 9.490 1086.110 10.670 ;
        RECT 1084.930 -2.910 1086.110 -1.730 ;
        RECT 1084.930 -4.510 1086.110 -3.330 ;
        RECT 1102.930 1469.090 1104.110 1470.270 ;
        RECT 1102.930 1467.490 1104.110 1468.670 ;
        RECT 1102.930 1289.090 1104.110 1290.270 ;
        RECT 1102.930 1287.490 1104.110 1288.670 ;
        RECT 1102.930 1109.090 1104.110 1110.270 ;
        RECT 1102.930 1107.490 1104.110 1108.670 ;
        RECT 1102.930 929.090 1104.110 930.270 ;
        RECT 1102.930 927.490 1104.110 928.670 ;
        RECT 1102.930 749.090 1104.110 750.270 ;
        RECT 1102.930 747.490 1104.110 748.670 ;
        RECT 1102.930 569.090 1104.110 570.270 ;
        RECT 1102.930 567.490 1104.110 568.670 ;
        RECT 1102.930 389.090 1104.110 390.270 ;
        RECT 1102.930 387.490 1104.110 388.670 ;
        RECT 1102.930 209.090 1104.110 210.270 ;
        RECT 1102.930 207.490 1104.110 208.670 ;
        RECT 1102.930 29.090 1104.110 30.270 ;
        RECT 1102.930 27.490 1104.110 28.670 ;
        RECT 1102.930 -12.310 1104.110 -11.130 ;
        RECT 1102.930 -13.910 1104.110 -12.730 ;
        RECT 1120.930 1307.090 1122.110 1308.270 ;
        RECT 1120.930 1305.490 1122.110 1306.670 ;
        RECT 1120.930 1127.090 1122.110 1128.270 ;
        RECT 1120.930 1125.490 1122.110 1126.670 ;
        RECT 1120.930 947.090 1122.110 948.270 ;
        RECT 1120.930 945.490 1122.110 946.670 ;
        RECT 1120.930 767.090 1122.110 768.270 ;
        RECT 1120.930 765.490 1122.110 766.670 ;
        RECT 1120.930 587.090 1122.110 588.270 ;
        RECT 1120.930 585.490 1122.110 586.670 ;
        RECT 1120.930 407.090 1122.110 408.270 ;
        RECT 1120.930 405.490 1122.110 406.670 ;
        RECT 1120.930 227.090 1122.110 228.270 ;
        RECT 1120.930 225.490 1122.110 226.670 ;
        RECT 1120.930 47.090 1122.110 48.270 ;
        RECT 1120.930 45.490 1122.110 46.670 ;
        RECT 1120.930 -21.710 1122.110 -20.530 ;
        RECT 1120.930 -23.310 1122.110 -22.130 ;
        RECT 1138.930 1325.090 1140.110 1326.270 ;
        RECT 1138.930 1323.490 1140.110 1324.670 ;
        RECT 1138.930 1145.090 1140.110 1146.270 ;
        RECT 1138.930 1143.490 1140.110 1144.670 ;
        RECT 1138.930 965.090 1140.110 966.270 ;
        RECT 1138.930 963.490 1140.110 964.670 ;
        RECT 1138.930 785.090 1140.110 786.270 ;
        RECT 1138.930 783.490 1140.110 784.670 ;
        RECT 1138.930 605.090 1140.110 606.270 ;
        RECT 1138.930 603.490 1140.110 604.670 ;
        RECT 1138.930 425.090 1140.110 426.270 ;
        RECT 1138.930 423.490 1140.110 424.670 ;
        RECT 1138.930 245.090 1140.110 246.270 ;
        RECT 1138.930 243.490 1140.110 244.670 ;
        RECT 1138.930 65.090 1140.110 66.270 ;
        RECT 1138.930 63.490 1140.110 64.670 ;
        RECT 958.930 -31.110 960.110 -29.930 ;
        RECT 958.930 -32.710 960.110 -31.530 ;
        RECT 1264.930 1451.090 1266.110 1452.270 ;
        RECT 1264.930 1449.490 1266.110 1450.670 ;
        RECT 1264.930 1271.090 1266.110 1272.270 ;
        RECT 1264.930 1269.490 1266.110 1270.670 ;
        RECT 1264.930 1091.090 1266.110 1092.270 ;
        RECT 1264.930 1089.490 1266.110 1090.670 ;
        RECT 1264.930 911.090 1266.110 912.270 ;
        RECT 1264.930 909.490 1266.110 910.670 ;
        RECT 1264.930 731.090 1266.110 732.270 ;
        RECT 1264.930 729.490 1266.110 730.670 ;
        RECT 1264.930 551.090 1266.110 552.270 ;
        RECT 1264.930 549.490 1266.110 550.670 ;
        RECT 1264.930 371.090 1266.110 372.270 ;
        RECT 1264.930 369.490 1266.110 370.670 ;
        RECT 1264.930 191.090 1266.110 192.270 ;
        RECT 1264.930 189.490 1266.110 190.670 ;
        RECT 1264.930 11.090 1266.110 12.270 ;
        RECT 1264.930 9.490 1266.110 10.670 ;
        RECT 1264.930 -2.910 1266.110 -1.730 ;
        RECT 1264.930 -4.510 1266.110 -3.330 ;
        RECT 1282.930 1469.090 1284.110 1470.270 ;
        RECT 1282.930 1467.490 1284.110 1468.670 ;
        RECT 1282.930 1289.090 1284.110 1290.270 ;
        RECT 1282.930 1287.490 1284.110 1288.670 ;
        RECT 1282.930 1109.090 1284.110 1110.270 ;
        RECT 1282.930 1107.490 1284.110 1108.670 ;
        RECT 1282.930 929.090 1284.110 930.270 ;
        RECT 1282.930 927.490 1284.110 928.670 ;
        RECT 1282.930 749.090 1284.110 750.270 ;
        RECT 1282.930 747.490 1284.110 748.670 ;
        RECT 1282.930 569.090 1284.110 570.270 ;
        RECT 1282.930 567.490 1284.110 568.670 ;
        RECT 1282.930 389.090 1284.110 390.270 ;
        RECT 1282.930 387.490 1284.110 388.670 ;
        RECT 1282.930 209.090 1284.110 210.270 ;
        RECT 1282.930 207.490 1284.110 208.670 ;
        RECT 1282.930 29.090 1284.110 30.270 ;
        RECT 1282.930 27.490 1284.110 28.670 ;
        RECT 1282.930 -12.310 1284.110 -11.130 ;
        RECT 1282.930 -13.910 1284.110 -12.730 ;
        RECT 1300.930 1307.090 1302.110 1308.270 ;
        RECT 1300.930 1305.490 1302.110 1306.670 ;
        RECT 1300.930 1127.090 1302.110 1128.270 ;
        RECT 1300.930 1125.490 1302.110 1126.670 ;
        RECT 1300.930 947.090 1302.110 948.270 ;
        RECT 1300.930 945.490 1302.110 946.670 ;
        RECT 1300.930 767.090 1302.110 768.270 ;
        RECT 1300.930 765.490 1302.110 766.670 ;
        RECT 1300.930 587.090 1302.110 588.270 ;
        RECT 1300.930 585.490 1302.110 586.670 ;
        RECT 1300.930 407.090 1302.110 408.270 ;
        RECT 1300.930 405.490 1302.110 406.670 ;
        RECT 1300.930 227.090 1302.110 228.270 ;
        RECT 1300.930 225.490 1302.110 226.670 ;
        RECT 1300.930 47.090 1302.110 48.270 ;
        RECT 1300.930 45.490 1302.110 46.670 ;
        RECT 1300.930 -21.710 1302.110 -20.530 ;
        RECT 1300.930 -23.310 1302.110 -22.130 ;
        RECT 1318.930 1325.090 1320.110 1326.270 ;
        RECT 1318.930 1323.490 1320.110 1324.670 ;
        RECT 1318.930 1145.090 1320.110 1146.270 ;
        RECT 1318.930 1143.490 1320.110 1144.670 ;
        RECT 1318.930 965.090 1320.110 966.270 ;
        RECT 1318.930 963.490 1320.110 964.670 ;
        RECT 1318.930 785.090 1320.110 786.270 ;
        RECT 1318.930 783.490 1320.110 784.670 ;
        RECT 1318.930 605.090 1320.110 606.270 ;
        RECT 1318.930 603.490 1320.110 604.670 ;
        RECT 1318.930 425.090 1320.110 426.270 ;
        RECT 1318.930 423.490 1320.110 424.670 ;
        RECT 1318.930 245.090 1320.110 246.270 ;
        RECT 1318.930 243.490 1320.110 244.670 ;
        RECT 1318.930 65.090 1320.110 66.270 ;
        RECT 1318.930 63.490 1320.110 64.670 ;
        RECT 1138.930 -31.110 1140.110 -29.930 ;
        RECT 1138.930 -32.710 1140.110 -31.530 ;
        RECT 1444.930 1451.090 1446.110 1452.270 ;
        RECT 1444.930 1449.490 1446.110 1450.670 ;
        RECT 1444.930 1271.090 1446.110 1272.270 ;
        RECT 1444.930 1269.490 1446.110 1270.670 ;
        RECT 1444.930 1091.090 1446.110 1092.270 ;
        RECT 1444.930 1089.490 1446.110 1090.670 ;
        RECT 1444.930 911.090 1446.110 912.270 ;
        RECT 1444.930 909.490 1446.110 910.670 ;
        RECT 1444.930 731.090 1446.110 732.270 ;
        RECT 1444.930 729.490 1446.110 730.670 ;
        RECT 1444.930 551.090 1446.110 552.270 ;
        RECT 1444.930 549.490 1446.110 550.670 ;
        RECT 1444.930 371.090 1446.110 372.270 ;
        RECT 1444.930 369.490 1446.110 370.670 ;
        RECT 1444.930 191.090 1446.110 192.270 ;
        RECT 1444.930 189.490 1446.110 190.670 ;
        RECT 1444.930 11.090 1446.110 12.270 ;
        RECT 1444.930 9.490 1446.110 10.670 ;
        RECT 1444.930 -2.910 1446.110 -1.730 ;
        RECT 1444.930 -4.510 1446.110 -3.330 ;
        RECT 1462.930 3449.090 1464.110 3450.270 ;
        RECT 1462.930 3447.490 1464.110 3448.670 ;
        RECT 1462.930 3269.090 1464.110 3270.270 ;
        RECT 1462.930 3267.490 1464.110 3268.670 ;
        RECT 1462.930 3089.090 1464.110 3090.270 ;
        RECT 1462.930 3087.490 1464.110 3088.670 ;
        RECT 1462.930 2909.090 1464.110 2910.270 ;
        RECT 1462.930 2907.490 1464.110 2908.670 ;
        RECT 1462.930 2729.090 1464.110 2730.270 ;
        RECT 1462.930 2727.490 1464.110 2728.670 ;
        RECT 1462.930 2549.090 1464.110 2550.270 ;
        RECT 1462.930 2547.490 1464.110 2548.670 ;
        RECT 1462.930 2369.090 1464.110 2370.270 ;
        RECT 1462.930 2367.490 1464.110 2368.670 ;
        RECT 1462.930 2189.090 1464.110 2190.270 ;
        RECT 1462.930 2187.490 1464.110 2188.670 ;
        RECT 1462.930 2009.090 1464.110 2010.270 ;
        RECT 1462.930 2007.490 1464.110 2008.670 ;
        RECT 1462.930 1829.090 1464.110 1830.270 ;
        RECT 1462.930 1827.490 1464.110 1828.670 ;
        RECT 1462.930 1649.090 1464.110 1650.270 ;
        RECT 1462.930 1647.490 1464.110 1648.670 ;
        RECT 1462.930 1469.090 1464.110 1470.270 ;
        RECT 1462.930 1467.490 1464.110 1468.670 ;
        RECT 1462.930 1289.090 1464.110 1290.270 ;
        RECT 1462.930 1287.490 1464.110 1288.670 ;
        RECT 1462.930 1109.090 1464.110 1110.270 ;
        RECT 1462.930 1107.490 1464.110 1108.670 ;
        RECT 1462.930 929.090 1464.110 930.270 ;
        RECT 1462.930 927.490 1464.110 928.670 ;
        RECT 1462.930 749.090 1464.110 750.270 ;
        RECT 1462.930 747.490 1464.110 748.670 ;
        RECT 1462.930 569.090 1464.110 570.270 ;
        RECT 1462.930 567.490 1464.110 568.670 ;
        RECT 1462.930 389.090 1464.110 390.270 ;
        RECT 1462.930 387.490 1464.110 388.670 ;
        RECT 1462.930 209.090 1464.110 210.270 ;
        RECT 1462.930 207.490 1464.110 208.670 ;
        RECT 1462.930 29.090 1464.110 30.270 ;
        RECT 1462.930 27.490 1464.110 28.670 ;
        RECT 1462.930 -12.310 1464.110 -11.130 ;
        RECT 1462.930 -13.910 1464.110 -12.730 ;
        RECT 1480.930 3467.090 1482.110 3468.270 ;
        RECT 1480.930 3465.490 1482.110 3466.670 ;
        RECT 1480.930 3287.090 1482.110 3288.270 ;
        RECT 1480.930 3285.490 1482.110 3286.670 ;
        RECT 1480.930 3107.090 1482.110 3108.270 ;
        RECT 1480.930 3105.490 1482.110 3106.670 ;
        RECT 1480.930 2927.090 1482.110 2928.270 ;
        RECT 1480.930 2925.490 1482.110 2926.670 ;
        RECT 1480.930 2747.090 1482.110 2748.270 ;
        RECT 1480.930 2745.490 1482.110 2746.670 ;
        RECT 1480.930 2567.090 1482.110 2568.270 ;
        RECT 1480.930 2565.490 1482.110 2566.670 ;
        RECT 1480.930 2387.090 1482.110 2388.270 ;
        RECT 1480.930 2385.490 1482.110 2386.670 ;
        RECT 1480.930 2207.090 1482.110 2208.270 ;
        RECT 1480.930 2205.490 1482.110 2206.670 ;
        RECT 1480.930 2027.090 1482.110 2028.270 ;
        RECT 1480.930 2025.490 1482.110 2026.670 ;
        RECT 1480.930 1847.090 1482.110 1848.270 ;
        RECT 1480.930 1845.490 1482.110 1846.670 ;
        RECT 1480.930 1667.090 1482.110 1668.270 ;
        RECT 1480.930 1665.490 1482.110 1666.670 ;
        RECT 1480.930 1487.090 1482.110 1488.270 ;
        RECT 1480.930 1485.490 1482.110 1486.670 ;
        RECT 1480.930 1307.090 1482.110 1308.270 ;
        RECT 1480.930 1305.490 1482.110 1306.670 ;
        RECT 1480.930 1127.090 1482.110 1128.270 ;
        RECT 1480.930 1125.490 1482.110 1126.670 ;
        RECT 1480.930 947.090 1482.110 948.270 ;
        RECT 1480.930 945.490 1482.110 946.670 ;
        RECT 1480.930 767.090 1482.110 768.270 ;
        RECT 1480.930 765.490 1482.110 766.670 ;
        RECT 1480.930 587.090 1482.110 588.270 ;
        RECT 1480.930 585.490 1482.110 586.670 ;
        RECT 1480.930 407.090 1482.110 408.270 ;
        RECT 1480.930 405.490 1482.110 406.670 ;
        RECT 1480.930 227.090 1482.110 228.270 ;
        RECT 1480.930 225.490 1482.110 226.670 ;
        RECT 1480.930 47.090 1482.110 48.270 ;
        RECT 1480.930 45.490 1482.110 46.670 ;
        RECT 1480.930 -21.710 1482.110 -20.530 ;
        RECT 1480.930 -23.310 1482.110 -22.130 ;
        RECT 1678.930 3551.210 1680.110 3552.390 ;
        RECT 1678.930 3549.610 1680.110 3550.790 ;
        RECT 1660.930 3541.810 1662.110 3542.990 ;
        RECT 1660.930 3540.210 1662.110 3541.390 ;
        RECT 1642.930 3532.410 1644.110 3533.590 ;
        RECT 1642.930 3530.810 1644.110 3531.990 ;
        RECT 1498.930 3485.090 1500.110 3486.270 ;
        RECT 1498.930 3483.490 1500.110 3484.670 ;
        RECT 1498.930 3305.090 1500.110 3306.270 ;
        RECT 1498.930 3303.490 1500.110 3304.670 ;
        RECT 1624.930 3523.010 1626.110 3524.190 ;
        RECT 1624.930 3521.410 1626.110 3522.590 ;
        RECT 1624.930 3431.090 1626.110 3432.270 ;
        RECT 1624.930 3429.490 1626.110 3430.670 ;
        RECT 1642.930 3449.090 1644.110 3450.270 ;
        RECT 1642.930 3447.490 1644.110 3448.670 ;
        RECT 1660.930 3467.090 1662.110 3468.270 ;
        RECT 1660.930 3465.490 1662.110 3466.670 ;
        RECT 1660.930 3287.090 1662.110 3288.270 ;
        RECT 1660.930 3285.490 1662.110 3286.670 ;
        RECT 1858.930 3551.210 1860.110 3552.390 ;
        RECT 1858.930 3549.610 1860.110 3550.790 ;
        RECT 1840.930 3541.810 1842.110 3542.990 ;
        RECT 1840.930 3540.210 1842.110 3541.390 ;
        RECT 1822.930 3532.410 1824.110 3533.590 ;
        RECT 1822.930 3530.810 1824.110 3531.990 ;
        RECT 1678.930 3485.090 1680.110 3486.270 ;
        RECT 1678.930 3483.490 1680.110 3484.670 ;
        RECT 1678.930 3305.090 1680.110 3306.270 ;
        RECT 1678.930 3303.490 1680.110 3304.670 ;
        RECT 1804.930 3523.010 1806.110 3524.190 ;
        RECT 1804.930 3521.410 1806.110 3522.590 ;
        RECT 1804.930 3431.090 1806.110 3432.270 ;
        RECT 1804.930 3429.490 1806.110 3430.670 ;
        RECT 1822.930 3449.090 1824.110 3450.270 ;
        RECT 1822.930 3447.490 1824.110 3448.670 ;
        RECT 1840.930 3467.090 1842.110 3468.270 ;
        RECT 1840.930 3465.490 1842.110 3466.670 ;
        RECT 1840.930 3287.090 1842.110 3288.270 ;
        RECT 1840.930 3285.490 1842.110 3286.670 ;
        RECT 2038.930 3551.210 2040.110 3552.390 ;
        RECT 2038.930 3549.610 2040.110 3550.790 ;
        RECT 2020.930 3541.810 2022.110 3542.990 ;
        RECT 2020.930 3540.210 2022.110 3541.390 ;
        RECT 2002.930 3532.410 2004.110 3533.590 ;
        RECT 2002.930 3530.810 2004.110 3531.990 ;
        RECT 1858.930 3485.090 1860.110 3486.270 ;
        RECT 1858.930 3483.490 1860.110 3484.670 ;
        RECT 1858.930 3305.090 1860.110 3306.270 ;
        RECT 1858.930 3303.490 1860.110 3304.670 ;
        RECT 1984.930 3523.010 1986.110 3524.190 ;
        RECT 1984.930 3521.410 1986.110 3522.590 ;
        RECT 1984.930 3431.090 1986.110 3432.270 ;
        RECT 1984.930 3429.490 1986.110 3430.670 ;
        RECT 1984.930 3251.090 1986.110 3252.270 ;
        RECT 1984.930 3249.490 1986.110 3250.670 ;
        RECT 1498.930 3125.090 1500.110 3126.270 ;
        RECT 1498.930 3123.490 1500.110 3124.670 ;
        RECT 1498.930 2945.090 1500.110 2946.270 ;
        RECT 1498.930 2943.490 1500.110 2944.670 ;
        RECT 1932.680 3125.090 1933.860 3126.270 ;
        RECT 1932.680 3123.490 1933.860 3124.670 ;
        RECT 1932.680 3107.090 1933.860 3108.270 ;
        RECT 1932.680 3105.490 1933.860 3106.670 ;
        RECT 1932.680 3089.090 1933.860 3090.270 ;
        RECT 1932.680 3087.490 1933.860 3088.670 ;
        RECT 1932.680 3071.090 1933.860 3072.270 ;
        RECT 1932.680 3069.490 1933.860 3070.670 ;
        RECT 1932.680 2945.090 1933.860 2946.270 ;
        RECT 1932.680 2943.490 1933.860 2944.670 ;
        RECT 1932.680 2927.090 1933.860 2928.270 ;
        RECT 1932.680 2925.490 1933.860 2926.670 ;
        RECT 1932.680 2909.090 1933.860 2910.270 ;
        RECT 1932.680 2907.490 1933.860 2908.670 ;
        RECT 1932.680 2891.090 1933.860 2892.270 ;
        RECT 1932.680 2889.490 1933.860 2890.670 ;
        RECT 1984.930 3071.090 1986.110 3072.270 ;
        RECT 1984.930 3069.490 1986.110 3070.670 ;
        RECT 1984.930 2891.090 1986.110 2892.270 ;
        RECT 1984.930 2889.490 1986.110 2890.670 ;
        RECT 1498.930 2765.090 1500.110 2766.270 ;
        RECT 1498.930 2763.490 1500.110 2764.670 ;
        RECT 1498.930 2585.090 1500.110 2586.270 ;
        RECT 1498.930 2583.490 1500.110 2584.670 ;
        RECT 1498.930 2405.090 1500.110 2406.270 ;
        RECT 1498.930 2403.490 1500.110 2404.670 ;
        RECT 1498.930 2225.090 1500.110 2226.270 ;
        RECT 1498.930 2223.490 1500.110 2224.670 ;
        RECT 1498.930 2045.090 1500.110 2046.270 ;
        RECT 1498.930 2043.490 1500.110 2044.670 ;
        RECT 1498.930 1865.090 1500.110 1866.270 ;
        RECT 1498.930 1863.490 1500.110 1864.670 ;
        RECT 1498.930 1685.090 1500.110 1686.270 ;
        RECT 1498.930 1683.490 1500.110 1684.670 ;
        RECT 1498.930 1505.090 1500.110 1506.270 ;
        RECT 1498.930 1503.490 1500.110 1504.670 ;
        RECT 1498.930 1325.090 1500.110 1326.270 ;
        RECT 1498.930 1323.490 1500.110 1324.670 ;
        RECT 1498.930 1145.090 1500.110 1146.270 ;
        RECT 1498.930 1143.490 1500.110 1144.670 ;
        RECT 1498.930 965.090 1500.110 966.270 ;
        RECT 1498.930 963.490 1500.110 964.670 ;
        RECT 1498.930 785.090 1500.110 786.270 ;
        RECT 1498.930 783.490 1500.110 784.670 ;
        RECT 1498.930 605.090 1500.110 606.270 ;
        RECT 1498.930 603.490 1500.110 604.670 ;
        RECT 1498.930 425.090 1500.110 426.270 ;
        RECT 1498.930 423.490 1500.110 424.670 ;
        RECT 1498.930 245.090 1500.110 246.270 ;
        RECT 1498.930 243.490 1500.110 244.670 ;
        RECT 1498.930 65.090 1500.110 66.270 ;
        RECT 1498.930 63.490 1500.110 64.670 ;
        RECT 1318.930 -31.110 1320.110 -29.930 ;
        RECT 1318.930 -32.710 1320.110 -31.530 ;
        RECT 1624.930 2711.090 1626.110 2712.270 ;
        RECT 1624.930 2709.490 1626.110 2710.670 ;
        RECT 1624.930 2531.090 1626.110 2532.270 ;
        RECT 1624.930 2529.490 1626.110 2530.670 ;
        RECT 1624.930 2351.090 1626.110 2352.270 ;
        RECT 1624.930 2349.490 1626.110 2350.670 ;
        RECT 1624.930 2171.090 1626.110 2172.270 ;
        RECT 1624.930 2169.490 1626.110 2170.670 ;
        RECT 1624.930 1991.090 1626.110 1992.270 ;
        RECT 1624.930 1989.490 1626.110 1990.670 ;
        RECT 1624.930 1811.090 1626.110 1812.270 ;
        RECT 1624.930 1809.490 1626.110 1810.670 ;
        RECT 1624.930 1631.090 1626.110 1632.270 ;
        RECT 1624.930 1629.490 1626.110 1630.670 ;
        RECT 1624.930 1451.090 1626.110 1452.270 ;
        RECT 1624.930 1449.490 1626.110 1450.670 ;
        RECT 1624.930 1271.090 1626.110 1272.270 ;
        RECT 1624.930 1269.490 1626.110 1270.670 ;
        RECT 1624.930 1091.090 1626.110 1092.270 ;
        RECT 1624.930 1089.490 1626.110 1090.670 ;
        RECT 1624.930 911.090 1626.110 912.270 ;
        RECT 1624.930 909.490 1626.110 910.670 ;
        RECT 1624.930 731.090 1626.110 732.270 ;
        RECT 1624.930 729.490 1626.110 730.670 ;
        RECT 1624.930 551.090 1626.110 552.270 ;
        RECT 1624.930 549.490 1626.110 550.670 ;
        RECT 1624.930 371.090 1626.110 372.270 ;
        RECT 1624.930 369.490 1626.110 370.670 ;
        RECT 1624.930 191.090 1626.110 192.270 ;
        RECT 1624.930 189.490 1626.110 190.670 ;
        RECT 1624.930 11.090 1626.110 12.270 ;
        RECT 1624.930 9.490 1626.110 10.670 ;
        RECT 1624.930 -2.910 1626.110 -1.730 ;
        RECT 1624.930 -4.510 1626.110 -3.330 ;
        RECT 1642.930 2729.090 1644.110 2730.270 ;
        RECT 1642.930 2727.490 1644.110 2728.670 ;
        RECT 1642.930 2549.090 1644.110 2550.270 ;
        RECT 1642.930 2547.490 1644.110 2548.670 ;
        RECT 1642.930 2369.090 1644.110 2370.270 ;
        RECT 1642.930 2367.490 1644.110 2368.670 ;
        RECT 1642.930 2189.090 1644.110 2190.270 ;
        RECT 1642.930 2187.490 1644.110 2188.670 ;
        RECT 1642.930 2009.090 1644.110 2010.270 ;
        RECT 1642.930 2007.490 1644.110 2008.670 ;
        RECT 1642.930 1829.090 1644.110 1830.270 ;
        RECT 1642.930 1827.490 1644.110 1828.670 ;
        RECT 1642.930 1649.090 1644.110 1650.270 ;
        RECT 1642.930 1647.490 1644.110 1648.670 ;
        RECT 1642.930 1469.090 1644.110 1470.270 ;
        RECT 1642.930 1467.490 1644.110 1468.670 ;
        RECT 1642.930 1289.090 1644.110 1290.270 ;
        RECT 1642.930 1287.490 1644.110 1288.670 ;
        RECT 1642.930 1109.090 1644.110 1110.270 ;
        RECT 1642.930 1107.490 1644.110 1108.670 ;
        RECT 1642.930 929.090 1644.110 930.270 ;
        RECT 1642.930 927.490 1644.110 928.670 ;
        RECT 1642.930 749.090 1644.110 750.270 ;
        RECT 1642.930 747.490 1644.110 748.670 ;
        RECT 1642.930 569.090 1644.110 570.270 ;
        RECT 1642.930 567.490 1644.110 568.670 ;
        RECT 1642.930 389.090 1644.110 390.270 ;
        RECT 1642.930 387.490 1644.110 388.670 ;
        RECT 1642.930 209.090 1644.110 210.270 ;
        RECT 1642.930 207.490 1644.110 208.670 ;
        RECT 1642.930 29.090 1644.110 30.270 ;
        RECT 1642.930 27.490 1644.110 28.670 ;
        RECT 1642.930 -12.310 1644.110 -11.130 ;
        RECT 1642.930 -13.910 1644.110 -12.730 ;
        RECT 1660.930 2747.090 1662.110 2748.270 ;
        RECT 1660.930 2745.490 1662.110 2746.670 ;
        RECT 1660.930 2567.090 1662.110 2568.270 ;
        RECT 1660.930 2565.490 1662.110 2566.670 ;
        RECT 1660.930 2387.090 1662.110 2388.270 ;
        RECT 1660.930 2385.490 1662.110 2386.670 ;
        RECT 1660.930 2207.090 1662.110 2208.270 ;
        RECT 1660.930 2205.490 1662.110 2206.670 ;
        RECT 1660.930 2027.090 1662.110 2028.270 ;
        RECT 1660.930 2025.490 1662.110 2026.670 ;
        RECT 1660.930 1847.090 1662.110 1848.270 ;
        RECT 1660.930 1845.490 1662.110 1846.670 ;
        RECT 1660.930 1667.090 1662.110 1668.270 ;
        RECT 1660.930 1665.490 1662.110 1666.670 ;
        RECT 1660.930 1487.090 1662.110 1488.270 ;
        RECT 1660.930 1485.490 1662.110 1486.670 ;
        RECT 1660.930 1307.090 1662.110 1308.270 ;
        RECT 1660.930 1305.490 1662.110 1306.670 ;
        RECT 1660.930 1127.090 1662.110 1128.270 ;
        RECT 1660.930 1125.490 1662.110 1126.670 ;
        RECT 1660.930 947.090 1662.110 948.270 ;
        RECT 1660.930 945.490 1662.110 946.670 ;
        RECT 1660.930 767.090 1662.110 768.270 ;
        RECT 1660.930 765.490 1662.110 766.670 ;
        RECT 1660.930 587.090 1662.110 588.270 ;
        RECT 1660.930 585.490 1662.110 586.670 ;
        RECT 1660.930 407.090 1662.110 408.270 ;
        RECT 1660.930 405.490 1662.110 406.670 ;
        RECT 1660.930 227.090 1662.110 228.270 ;
        RECT 1660.930 225.490 1662.110 226.670 ;
        RECT 1660.930 47.090 1662.110 48.270 ;
        RECT 1660.930 45.490 1662.110 46.670 ;
        RECT 1660.930 -21.710 1662.110 -20.530 ;
        RECT 1660.930 -23.310 1662.110 -22.130 ;
        RECT 1678.930 2765.090 1680.110 2766.270 ;
        RECT 1678.930 2763.490 1680.110 2764.670 ;
        RECT 1678.930 2585.090 1680.110 2586.270 ;
        RECT 1678.930 2583.490 1680.110 2584.670 ;
        RECT 1678.930 2405.090 1680.110 2406.270 ;
        RECT 1678.930 2403.490 1680.110 2404.670 ;
        RECT 1678.930 2225.090 1680.110 2226.270 ;
        RECT 1678.930 2223.490 1680.110 2224.670 ;
        RECT 1678.930 2045.090 1680.110 2046.270 ;
        RECT 1678.930 2043.490 1680.110 2044.670 ;
        RECT 1678.930 1865.090 1680.110 1866.270 ;
        RECT 1678.930 1863.490 1680.110 1864.670 ;
        RECT 1678.930 1685.090 1680.110 1686.270 ;
        RECT 1678.930 1683.490 1680.110 1684.670 ;
        RECT 1678.930 1505.090 1680.110 1506.270 ;
        RECT 1678.930 1503.490 1680.110 1504.670 ;
        RECT 1678.930 1325.090 1680.110 1326.270 ;
        RECT 1678.930 1323.490 1680.110 1324.670 ;
        RECT 1678.930 1145.090 1680.110 1146.270 ;
        RECT 1678.930 1143.490 1680.110 1144.670 ;
        RECT 1678.930 965.090 1680.110 966.270 ;
        RECT 1678.930 963.490 1680.110 964.670 ;
        RECT 1678.930 785.090 1680.110 786.270 ;
        RECT 1678.930 783.490 1680.110 784.670 ;
        RECT 1678.930 605.090 1680.110 606.270 ;
        RECT 1678.930 603.490 1680.110 604.670 ;
        RECT 1678.930 425.090 1680.110 426.270 ;
        RECT 1678.930 423.490 1680.110 424.670 ;
        RECT 1678.930 245.090 1680.110 246.270 ;
        RECT 1678.930 243.490 1680.110 244.670 ;
        RECT 1678.930 65.090 1680.110 66.270 ;
        RECT 1678.930 63.490 1680.110 64.670 ;
        RECT 1498.930 -31.110 1500.110 -29.930 ;
        RECT 1498.930 -32.710 1500.110 -31.530 ;
        RECT 1804.930 2711.090 1806.110 2712.270 ;
        RECT 1804.930 2709.490 1806.110 2710.670 ;
        RECT 1804.930 2531.090 1806.110 2532.270 ;
        RECT 1804.930 2529.490 1806.110 2530.670 ;
        RECT 1804.930 2351.090 1806.110 2352.270 ;
        RECT 1804.930 2349.490 1806.110 2350.670 ;
        RECT 1804.930 2171.090 1806.110 2172.270 ;
        RECT 1804.930 2169.490 1806.110 2170.670 ;
        RECT 1804.930 1991.090 1806.110 1992.270 ;
        RECT 1804.930 1989.490 1806.110 1990.670 ;
        RECT 1804.930 1811.090 1806.110 1812.270 ;
        RECT 1804.930 1809.490 1806.110 1810.670 ;
        RECT 1804.930 1631.090 1806.110 1632.270 ;
        RECT 1804.930 1629.490 1806.110 1630.670 ;
        RECT 1804.930 1451.090 1806.110 1452.270 ;
        RECT 1804.930 1449.490 1806.110 1450.670 ;
        RECT 1804.930 1271.090 1806.110 1272.270 ;
        RECT 1804.930 1269.490 1806.110 1270.670 ;
        RECT 1804.930 1091.090 1806.110 1092.270 ;
        RECT 1804.930 1089.490 1806.110 1090.670 ;
        RECT 1804.930 911.090 1806.110 912.270 ;
        RECT 1804.930 909.490 1806.110 910.670 ;
        RECT 1804.930 731.090 1806.110 732.270 ;
        RECT 1804.930 729.490 1806.110 730.670 ;
        RECT 1804.930 551.090 1806.110 552.270 ;
        RECT 1804.930 549.490 1806.110 550.670 ;
        RECT 1804.930 371.090 1806.110 372.270 ;
        RECT 1804.930 369.490 1806.110 370.670 ;
        RECT 1804.930 191.090 1806.110 192.270 ;
        RECT 1804.930 189.490 1806.110 190.670 ;
        RECT 1804.930 11.090 1806.110 12.270 ;
        RECT 1804.930 9.490 1806.110 10.670 ;
        RECT 1804.930 -2.910 1806.110 -1.730 ;
        RECT 1804.930 -4.510 1806.110 -3.330 ;
        RECT 1822.930 2729.090 1824.110 2730.270 ;
        RECT 1822.930 2727.490 1824.110 2728.670 ;
        RECT 1822.930 2549.090 1824.110 2550.270 ;
        RECT 1822.930 2547.490 1824.110 2548.670 ;
        RECT 1822.930 2369.090 1824.110 2370.270 ;
        RECT 1822.930 2367.490 1824.110 2368.670 ;
        RECT 1822.930 2189.090 1824.110 2190.270 ;
        RECT 1822.930 2187.490 1824.110 2188.670 ;
        RECT 1822.930 2009.090 1824.110 2010.270 ;
        RECT 1822.930 2007.490 1824.110 2008.670 ;
        RECT 1822.930 1829.090 1824.110 1830.270 ;
        RECT 1822.930 1827.490 1824.110 1828.670 ;
        RECT 1822.930 1649.090 1824.110 1650.270 ;
        RECT 1822.930 1647.490 1824.110 1648.670 ;
        RECT 1822.930 1469.090 1824.110 1470.270 ;
        RECT 1822.930 1467.490 1824.110 1468.670 ;
        RECT 1822.930 1289.090 1824.110 1290.270 ;
        RECT 1822.930 1287.490 1824.110 1288.670 ;
        RECT 1822.930 1109.090 1824.110 1110.270 ;
        RECT 1822.930 1107.490 1824.110 1108.670 ;
        RECT 1822.930 929.090 1824.110 930.270 ;
        RECT 1822.930 927.490 1824.110 928.670 ;
        RECT 1822.930 749.090 1824.110 750.270 ;
        RECT 1822.930 747.490 1824.110 748.670 ;
        RECT 1822.930 569.090 1824.110 570.270 ;
        RECT 1822.930 567.490 1824.110 568.670 ;
        RECT 1822.930 389.090 1824.110 390.270 ;
        RECT 1822.930 387.490 1824.110 388.670 ;
        RECT 1822.930 209.090 1824.110 210.270 ;
        RECT 1822.930 207.490 1824.110 208.670 ;
        RECT 1822.930 29.090 1824.110 30.270 ;
        RECT 1822.930 27.490 1824.110 28.670 ;
        RECT 1822.930 -12.310 1824.110 -11.130 ;
        RECT 1822.930 -13.910 1824.110 -12.730 ;
        RECT 1840.930 2747.090 1842.110 2748.270 ;
        RECT 1840.930 2745.490 1842.110 2746.670 ;
        RECT 1840.930 2567.090 1842.110 2568.270 ;
        RECT 1840.930 2565.490 1842.110 2566.670 ;
        RECT 1840.930 2387.090 1842.110 2388.270 ;
        RECT 1840.930 2385.490 1842.110 2386.670 ;
        RECT 1840.930 2207.090 1842.110 2208.270 ;
        RECT 1840.930 2205.490 1842.110 2206.670 ;
        RECT 1840.930 2027.090 1842.110 2028.270 ;
        RECT 1840.930 2025.490 1842.110 2026.670 ;
        RECT 1840.930 1847.090 1842.110 1848.270 ;
        RECT 1840.930 1845.490 1842.110 1846.670 ;
        RECT 1840.930 1667.090 1842.110 1668.270 ;
        RECT 1840.930 1665.490 1842.110 1666.670 ;
        RECT 1840.930 1487.090 1842.110 1488.270 ;
        RECT 1840.930 1485.490 1842.110 1486.670 ;
        RECT 1840.930 1307.090 1842.110 1308.270 ;
        RECT 1840.930 1305.490 1842.110 1306.670 ;
        RECT 1840.930 1127.090 1842.110 1128.270 ;
        RECT 1840.930 1125.490 1842.110 1126.670 ;
        RECT 1840.930 947.090 1842.110 948.270 ;
        RECT 1840.930 945.490 1842.110 946.670 ;
        RECT 1840.930 767.090 1842.110 768.270 ;
        RECT 1840.930 765.490 1842.110 766.670 ;
        RECT 1840.930 587.090 1842.110 588.270 ;
        RECT 1840.930 585.490 1842.110 586.670 ;
        RECT 1840.930 407.090 1842.110 408.270 ;
        RECT 1840.930 405.490 1842.110 406.670 ;
        RECT 1840.930 227.090 1842.110 228.270 ;
        RECT 1840.930 225.490 1842.110 226.670 ;
        RECT 1840.930 47.090 1842.110 48.270 ;
        RECT 1840.930 45.490 1842.110 46.670 ;
        RECT 1840.930 -21.710 1842.110 -20.530 ;
        RECT 1840.930 -23.310 1842.110 -22.130 ;
        RECT 1858.930 2765.090 1860.110 2766.270 ;
        RECT 1858.930 2763.490 1860.110 2764.670 ;
        RECT 1858.930 2585.090 1860.110 2586.270 ;
        RECT 1858.930 2583.490 1860.110 2584.670 ;
        RECT 1858.930 2405.090 1860.110 2406.270 ;
        RECT 1858.930 2403.490 1860.110 2404.670 ;
        RECT 1858.930 2225.090 1860.110 2226.270 ;
        RECT 1858.930 2223.490 1860.110 2224.670 ;
        RECT 1858.930 2045.090 1860.110 2046.270 ;
        RECT 1858.930 2043.490 1860.110 2044.670 ;
        RECT 1858.930 1865.090 1860.110 1866.270 ;
        RECT 1858.930 1863.490 1860.110 1864.670 ;
        RECT 1858.930 1685.090 1860.110 1686.270 ;
        RECT 1858.930 1683.490 1860.110 1684.670 ;
        RECT 1858.930 1505.090 1860.110 1506.270 ;
        RECT 1858.930 1503.490 1860.110 1504.670 ;
        RECT 1858.930 1325.090 1860.110 1326.270 ;
        RECT 1858.930 1323.490 1860.110 1324.670 ;
        RECT 1858.930 1145.090 1860.110 1146.270 ;
        RECT 1858.930 1143.490 1860.110 1144.670 ;
        RECT 1858.930 965.090 1860.110 966.270 ;
        RECT 1858.930 963.490 1860.110 964.670 ;
        RECT 1858.930 785.090 1860.110 786.270 ;
        RECT 1858.930 783.490 1860.110 784.670 ;
        RECT 1858.930 605.090 1860.110 606.270 ;
        RECT 1858.930 603.490 1860.110 604.670 ;
        RECT 1858.930 425.090 1860.110 426.270 ;
        RECT 1858.930 423.490 1860.110 424.670 ;
        RECT 1858.930 245.090 1860.110 246.270 ;
        RECT 1858.930 243.490 1860.110 244.670 ;
        RECT 1858.930 65.090 1860.110 66.270 ;
        RECT 1858.930 63.490 1860.110 64.670 ;
        RECT 1678.930 -31.110 1680.110 -29.930 ;
        RECT 1678.930 -32.710 1680.110 -31.530 ;
        RECT 1984.930 2711.090 1986.110 2712.270 ;
        RECT 1984.930 2709.490 1986.110 2710.670 ;
        RECT 1984.930 2531.090 1986.110 2532.270 ;
        RECT 1984.930 2529.490 1986.110 2530.670 ;
        RECT 1984.930 2351.090 1986.110 2352.270 ;
        RECT 1984.930 2349.490 1986.110 2350.670 ;
        RECT 1984.930 2171.090 1986.110 2172.270 ;
        RECT 1984.930 2169.490 1986.110 2170.670 ;
        RECT 1984.930 1991.090 1986.110 1992.270 ;
        RECT 1984.930 1989.490 1986.110 1990.670 ;
        RECT 1984.930 1811.090 1986.110 1812.270 ;
        RECT 1984.930 1809.490 1986.110 1810.670 ;
        RECT 1984.930 1631.090 1986.110 1632.270 ;
        RECT 1984.930 1629.490 1986.110 1630.670 ;
        RECT 1984.930 1451.090 1986.110 1452.270 ;
        RECT 1984.930 1449.490 1986.110 1450.670 ;
        RECT 1984.930 1271.090 1986.110 1272.270 ;
        RECT 1984.930 1269.490 1986.110 1270.670 ;
        RECT 1984.930 1091.090 1986.110 1092.270 ;
        RECT 1984.930 1089.490 1986.110 1090.670 ;
        RECT 1984.930 911.090 1986.110 912.270 ;
        RECT 1984.930 909.490 1986.110 910.670 ;
        RECT 1984.930 731.090 1986.110 732.270 ;
        RECT 1984.930 729.490 1986.110 730.670 ;
        RECT 1984.930 551.090 1986.110 552.270 ;
        RECT 1984.930 549.490 1986.110 550.670 ;
        RECT 1984.930 371.090 1986.110 372.270 ;
        RECT 1984.930 369.490 1986.110 370.670 ;
        RECT 1984.930 191.090 1986.110 192.270 ;
        RECT 1984.930 189.490 1986.110 190.670 ;
        RECT 1984.930 11.090 1986.110 12.270 ;
        RECT 1984.930 9.490 1986.110 10.670 ;
        RECT 1984.930 -2.910 1986.110 -1.730 ;
        RECT 1984.930 -4.510 1986.110 -3.330 ;
        RECT 2002.930 3449.090 2004.110 3450.270 ;
        RECT 2002.930 3447.490 2004.110 3448.670 ;
        RECT 2002.930 3269.090 2004.110 3270.270 ;
        RECT 2002.930 3267.490 2004.110 3268.670 ;
        RECT 2002.930 3089.090 2004.110 3090.270 ;
        RECT 2002.930 3087.490 2004.110 3088.670 ;
        RECT 2002.930 2909.090 2004.110 2910.270 ;
        RECT 2002.930 2907.490 2004.110 2908.670 ;
        RECT 2002.930 2729.090 2004.110 2730.270 ;
        RECT 2002.930 2727.490 2004.110 2728.670 ;
        RECT 2002.930 2549.090 2004.110 2550.270 ;
        RECT 2002.930 2547.490 2004.110 2548.670 ;
        RECT 2002.930 2369.090 2004.110 2370.270 ;
        RECT 2002.930 2367.490 2004.110 2368.670 ;
        RECT 2002.930 2189.090 2004.110 2190.270 ;
        RECT 2002.930 2187.490 2004.110 2188.670 ;
        RECT 2002.930 2009.090 2004.110 2010.270 ;
        RECT 2002.930 2007.490 2004.110 2008.670 ;
        RECT 2002.930 1829.090 2004.110 1830.270 ;
        RECT 2002.930 1827.490 2004.110 1828.670 ;
        RECT 2002.930 1649.090 2004.110 1650.270 ;
        RECT 2002.930 1647.490 2004.110 1648.670 ;
        RECT 2002.930 1469.090 2004.110 1470.270 ;
        RECT 2002.930 1467.490 2004.110 1468.670 ;
        RECT 2002.930 1289.090 2004.110 1290.270 ;
        RECT 2002.930 1287.490 2004.110 1288.670 ;
        RECT 2002.930 1109.090 2004.110 1110.270 ;
        RECT 2002.930 1107.490 2004.110 1108.670 ;
        RECT 2002.930 929.090 2004.110 930.270 ;
        RECT 2002.930 927.490 2004.110 928.670 ;
        RECT 2002.930 749.090 2004.110 750.270 ;
        RECT 2002.930 747.490 2004.110 748.670 ;
        RECT 2002.930 569.090 2004.110 570.270 ;
        RECT 2002.930 567.490 2004.110 568.670 ;
        RECT 2002.930 389.090 2004.110 390.270 ;
        RECT 2002.930 387.490 2004.110 388.670 ;
        RECT 2002.930 209.090 2004.110 210.270 ;
        RECT 2002.930 207.490 2004.110 208.670 ;
        RECT 2002.930 29.090 2004.110 30.270 ;
        RECT 2002.930 27.490 2004.110 28.670 ;
        RECT 2002.930 -12.310 2004.110 -11.130 ;
        RECT 2002.930 -13.910 2004.110 -12.730 ;
        RECT 2020.930 3467.090 2022.110 3468.270 ;
        RECT 2020.930 3465.490 2022.110 3466.670 ;
        RECT 2020.930 3287.090 2022.110 3288.270 ;
        RECT 2020.930 3285.490 2022.110 3286.670 ;
        RECT 2020.930 3107.090 2022.110 3108.270 ;
        RECT 2020.930 3105.490 2022.110 3106.670 ;
        RECT 2020.930 2927.090 2022.110 2928.270 ;
        RECT 2020.930 2925.490 2022.110 2926.670 ;
        RECT 2020.930 2747.090 2022.110 2748.270 ;
        RECT 2020.930 2745.490 2022.110 2746.670 ;
        RECT 2020.930 2567.090 2022.110 2568.270 ;
        RECT 2020.930 2565.490 2022.110 2566.670 ;
        RECT 2020.930 2387.090 2022.110 2388.270 ;
        RECT 2020.930 2385.490 2022.110 2386.670 ;
        RECT 2020.930 2207.090 2022.110 2208.270 ;
        RECT 2020.930 2205.490 2022.110 2206.670 ;
        RECT 2020.930 2027.090 2022.110 2028.270 ;
        RECT 2020.930 2025.490 2022.110 2026.670 ;
        RECT 2020.930 1847.090 2022.110 1848.270 ;
        RECT 2020.930 1845.490 2022.110 1846.670 ;
        RECT 2020.930 1667.090 2022.110 1668.270 ;
        RECT 2020.930 1665.490 2022.110 1666.670 ;
        RECT 2020.930 1487.090 2022.110 1488.270 ;
        RECT 2020.930 1485.490 2022.110 1486.670 ;
        RECT 2020.930 1307.090 2022.110 1308.270 ;
        RECT 2020.930 1305.490 2022.110 1306.670 ;
        RECT 2020.930 1127.090 2022.110 1128.270 ;
        RECT 2020.930 1125.490 2022.110 1126.670 ;
        RECT 2020.930 947.090 2022.110 948.270 ;
        RECT 2020.930 945.490 2022.110 946.670 ;
        RECT 2020.930 767.090 2022.110 768.270 ;
        RECT 2020.930 765.490 2022.110 766.670 ;
        RECT 2020.930 587.090 2022.110 588.270 ;
        RECT 2020.930 585.490 2022.110 586.670 ;
        RECT 2020.930 407.090 2022.110 408.270 ;
        RECT 2020.930 405.490 2022.110 406.670 ;
        RECT 2020.930 227.090 2022.110 228.270 ;
        RECT 2020.930 225.490 2022.110 226.670 ;
        RECT 2020.930 47.090 2022.110 48.270 ;
        RECT 2020.930 45.490 2022.110 46.670 ;
        RECT 2020.930 -21.710 2022.110 -20.530 ;
        RECT 2020.930 -23.310 2022.110 -22.130 ;
        RECT 2218.930 3551.210 2220.110 3552.390 ;
        RECT 2218.930 3549.610 2220.110 3550.790 ;
        RECT 2200.930 3541.810 2202.110 3542.990 ;
        RECT 2200.930 3540.210 2202.110 3541.390 ;
        RECT 2182.930 3532.410 2184.110 3533.590 ;
        RECT 2182.930 3530.810 2184.110 3531.990 ;
        RECT 2038.930 3485.090 2040.110 3486.270 ;
        RECT 2038.930 3483.490 2040.110 3484.670 ;
        RECT 2038.930 3305.090 2040.110 3306.270 ;
        RECT 2038.930 3303.490 2040.110 3304.670 ;
        RECT 2038.930 3125.090 2040.110 3126.270 ;
        RECT 2038.930 3123.490 2040.110 3124.670 ;
        RECT 2038.930 2945.090 2040.110 2946.270 ;
        RECT 2038.930 2943.490 2040.110 2944.670 ;
        RECT 2038.930 2765.090 2040.110 2766.270 ;
        RECT 2038.930 2763.490 2040.110 2764.670 ;
        RECT 2038.930 2585.090 2040.110 2586.270 ;
        RECT 2038.930 2583.490 2040.110 2584.670 ;
        RECT 2038.930 2405.090 2040.110 2406.270 ;
        RECT 2038.930 2403.490 2040.110 2404.670 ;
        RECT 2038.930 2225.090 2040.110 2226.270 ;
        RECT 2038.930 2223.490 2040.110 2224.670 ;
        RECT 2038.930 2045.090 2040.110 2046.270 ;
        RECT 2038.930 2043.490 2040.110 2044.670 ;
        RECT 2038.930 1865.090 2040.110 1866.270 ;
        RECT 2038.930 1863.490 2040.110 1864.670 ;
        RECT 2038.930 1685.090 2040.110 1686.270 ;
        RECT 2038.930 1683.490 2040.110 1684.670 ;
        RECT 2038.930 1505.090 2040.110 1506.270 ;
        RECT 2038.930 1503.490 2040.110 1504.670 ;
        RECT 2038.930 1325.090 2040.110 1326.270 ;
        RECT 2038.930 1323.490 2040.110 1324.670 ;
        RECT 2038.930 1145.090 2040.110 1146.270 ;
        RECT 2038.930 1143.490 2040.110 1144.670 ;
        RECT 2038.930 965.090 2040.110 966.270 ;
        RECT 2038.930 963.490 2040.110 964.670 ;
        RECT 2038.930 785.090 2040.110 786.270 ;
        RECT 2038.930 783.490 2040.110 784.670 ;
        RECT 2038.930 605.090 2040.110 606.270 ;
        RECT 2038.930 603.490 2040.110 604.670 ;
        RECT 2038.930 425.090 2040.110 426.270 ;
        RECT 2038.930 423.490 2040.110 424.670 ;
        RECT 2038.930 245.090 2040.110 246.270 ;
        RECT 2038.930 243.490 2040.110 244.670 ;
        RECT 2038.930 65.090 2040.110 66.270 ;
        RECT 2038.930 63.490 2040.110 64.670 ;
        RECT 1858.930 -31.110 1860.110 -29.930 ;
        RECT 1858.930 -32.710 1860.110 -31.530 ;
        RECT 2164.930 3523.010 2166.110 3524.190 ;
        RECT 2164.930 3521.410 2166.110 3522.590 ;
        RECT 2164.930 3431.090 2166.110 3432.270 ;
        RECT 2164.930 3429.490 2166.110 3430.670 ;
        RECT 2182.930 3449.090 2184.110 3450.270 ;
        RECT 2182.930 3447.490 2184.110 3448.670 ;
        RECT 2200.930 3467.090 2202.110 3468.270 ;
        RECT 2200.930 3465.490 2202.110 3466.670 ;
        RECT 2200.930 3287.090 2202.110 3288.270 ;
        RECT 2200.930 3285.490 2202.110 3286.670 ;
        RECT 2398.930 3551.210 2400.110 3552.390 ;
        RECT 2398.930 3549.610 2400.110 3550.790 ;
        RECT 2380.930 3541.810 2382.110 3542.990 ;
        RECT 2380.930 3540.210 2382.110 3541.390 ;
        RECT 2362.930 3532.410 2364.110 3533.590 ;
        RECT 2362.930 3530.810 2364.110 3531.990 ;
        RECT 2218.930 3485.090 2220.110 3486.270 ;
        RECT 2218.930 3483.490 2220.110 3484.670 ;
        RECT 2218.930 3305.090 2220.110 3306.270 ;
        RECT 2218.930 3303.490 2220.110 3304.670 ;
        RECT 2344.930 3523.010 2346.110 3524.190 ;
        RECT 2344.930 3521.410 2346.110 3522.590 ;
        RECT 2344.930 3431.090 2346.110 3432.270 ;
        RECT 2344.930 3429.490 2346.110 3430.670 ;
        RECT 2362.930 3449.090 2364.110 3450.270 ;
        RECT 2362.930 3447.490 2364.110 3448.670 ;
        RECT 2380.930 3467.090 2382.110 3468.270 ;
        RECT 2380.930 3465.490 2382.110 3466.670 ;
        RECT 2380.930 3287.090 2382.110 3288.270 ;
        RECT 2380.930 3285.490 2382.110 3286.670 ;
        RECT 2578.930 3551.210 2580.110 3552.390 ;
        RECT 2578.930 3549.610 2580.110 3550.790 ;
        RECT 2560.930 3541.810 2562.110 3542.990 ;
        RECT 2560.930 3540.210 2562.110 3541.390 ;
        RECT 2542.930 3532.410 2544.110 3533.590 ;
        RECT 2542.930 3530.810 2544.110 3531.990 ;
        RECT 2398.930 3485.090 2400.110 3486.270 ;
        RECT 2398.930 3483.490 2400.110 3484.670 ;
        RECT 2398.930 3305.090 2400.110 3306.270 ;
        RECT 2398.930 3303.490 2400.110 3304.670 ;
        RECT 2524.930 3523.010 2526.110 3524.190 ;
        RECT 2524.930 3521.410 2526.110 3522.590 ;
        RECT 2524.930 3431.090 2526.110 3432.270 ;
        RECT 2524.930 3429.490 2526.110 3430.670 ;
        RECT 2542.930 3449.090 2544.110 3450.270 ;
        RECT 2542.930 3447.490 2544.110 3448.670 ;
        RECT 2560.930 3467.090 2562.110 3468.270 ;
        RECT 2560.930 3465.490 2562.110 3466.670 ;
        RECT 2560.930 3287.090 2562.110 3288.270 ;
        RECT 2560.930 3285.490 2562.110 3286.670 ;
        RECT 2758.930 3551.210 2760.110 3552.390 ;
        RECT 2758.930 3549.610 2760.110 3550.790 ;
        RECT 2740.930 3541.810 2742.110 3542.990 ;
        RECT 2740.930 3540.210 2742.110 3541.390 ;
        RECT 2722.930 3532.410 2724.110 3533.590 ;
        RECT 2722.930 3530.810 2724.110 3531.990 ;
        RECT 2578.930 3485.090 2580.110 3486.270 ;
        RECT 2578.930 3483.490 2580.110 3484.670 ;
        RECT 2578.930 3305.090 2580.110 3306.270 ;
        RECT 2578.930 3303.490 2580.110 3304.670 ;
        RECT 2704.930 3523.010 2706.110 3524.190 ;
        RECT 2704.930 3521.410 2706.110 3522.590 ;
        RECT 2704.930 3431.090 2706.110 3432.270 ;
        RECT 2704.930 3429.490 2706.110 3430.670 ;
        RECT 2164.930 3251.090 2166.110 3252.270 ;
        RECT 2164.930 3249.490 2166.110 3250.670 ;
        RECT 2704.930 3251.090 2706.110 3252.270 ;
        RECT 2704.930 3249.490 2706.110 3250.670 ;
        RECT 2164.930 3071.090 2166.110 3072.270 ;
        RECT 2164.930 3069.490 2166.110 3070.670 ;
        RECT 2164.930 2891.090 2166.110 2892.270 ;
        RECT 2164.930 2889.490 2166.110 2890.670 ;
        RECT 2582.680 3125.090 2583.860 3126.270 ;
        RECT 2582.680 3123.490 2583.860 3124.670 ;
        RECT 2582.680 3107.090 2583.860 3108.270 ;
        RECT 2582.680 3105.490 2583.860 3106.670 ;
        RECT 2582.680 3089.090 2583.860 3090.270 ;
        RECT 2582.680 3087.490 2583.860 3088.670 ;
        RECT 2582.680 3071.090 2583.860 3072.270 ;
        RECT 2582.680 3069.490 2583.860 3070.670 ;
        RECT 2582.680 2945.090 2583.860 2946.270 ;
        RECT 2582.680 2943.490 2583.860 2944.670 ;
        RECT 2582.680 2927.090 2583.860 2928.270 ;
        RECT 2582.680 2925.490 2583.860 2926.670 ;
        RECT 2582.680 2909.090 2583.860 2910.270 ;
        RECT 2582.680 2907.490 2583.860 2908.670 ;
        RECT 2582.680 2891.090 2583.860 2892.270 ;
        RECT 2582.680 2889.490 2583.860 2890.670 ;
        RECT 2704.930 3071.090 2706.110 3072.270 ;
        RECT 2704.930 3069.490 2706.110 3070.670 ;
        RECT 2704.930 2891.090 2706.110 2892.270 ;
        RECT 2704.930 2889.490 2706.110 2890.670 ;
        RECT 2164.930 2711.090 2166.110 2712.270 ;
        RECT 2164.930 2709.490 2166.110 2710.670 ;
        RECT 2164.930 2531.090 2166.110 2532.270 ;
        RECT 2164.930 2529.490 2166.110 2530.670 ;
        RECT 2164.930 2351.090 2166.110 2352.270 ;
        RECT 2164.930 2349.490 2166.110 2350.670 ;
        RECT 2164.930 2171.090 2166.110 2172.270 ;
        RECT 2164.930 2169.490 2166.110 2170.670 ;
        RECT 2164.930 1991.090 2166.110 1992.270 ;
        RECT 2164.930 1989.490 2166.110 1990.670 ;
        RECT 2164.930 1811.090 2166.110 1812.270 ;
        RECT 2164.930 1809.490 2166.110 1810.670 ;
        RECT 2164.930 1631.090 2166.110 1632.270 ;
        RECT 2164.930 1629.490 2166.110 1630.670 ;
        RECT 2164.930 1451.090 2166.110 1452.270 ;
        RECT 2164.930 1449.490 2166.110 1450.670 ;
        RECT 2164.930 1271.090 2166.110 1272.270 ;
        RECT 2164.930 1269.490 2166.110 1270.670 ;
        RECT 2164.930 1091.090 2166.110 1092.270 ;
        RECT 2164.930 1089.490 2166.110 1090.670 ;
        RECT 2164.930 911.090 2166.110 912.270 ;
        RECT 2164.930 909.490 2166.110 910.670 ;
        RECT 2164.930 731.090 2166.110 732.270 ;
        RECT 2164.930 729.490 2166.110 730.670 ;
        RECT 2164.930 551.090 2166.110 552.270 ;
        RECT 2164.930 549.490 2166.110 550.670 ;
        RECT 2164.930 371.090 2166.110 372.270 ;
        RECT 2164.930 369.490 2166.110 370.670 ;
        RECT 2164.930 191.090 2166.110 192.270 ;
        RECT 2164.930 189.490 2166.110 190.670 ;
        RECT 2164.930 11.090 2166.110 12.270 ;
        RECT 2164.930 9.490 2166.110 10.670 ;
        RECT 2164.930 -2.910 2166.110 -1.730 ;
        RECT 2164.930 -4.510 2166.110 -3.330 ;
        RECT 2182.930 2729.090 2184.110 2730.270 ;
        RECT 2182.930 2727.490 2184.110 2728.670 ;
        RECT 2182.930 2549.090 2184.110 2550.270 ;
        RECT 2182.930 2547.490 2184.110 2548.670 ;
        RECT 2182.930 2369.090 2184.110 2370.270 ;
        RECT 2182.930 2367.490 2184.110 2368.670 ;
        RECT 2182.930 2189.090 2184.110 2190.270 ;
        RECT 2182.930 2187.490 2184.110 2188.670 ;
        RECT 2182.930 2009.090 2184.110 2010.270 ;
        RECT 2182.930 2007.490 2184.110 2008.670 ;
        RECT 2182.930 1829.090 2184.110 1830.270 ;
        RECT 2182.930 1827.490 2184.110 1828.670 ;
        RECT 2182.930 1649.090 2184.110 1650.270 ;
        RECT 2182.930 1647.490 2184.110 1648.670 ;
        RECT 2182.930 1469.090 2184.110 1470.270 ;
        RECT 2182.930 1467.490 2184.110 1468.670 ;
        RECT 2182.930 1289.090 2184.110 1290.270 ;
        RECT 2182.930 1287.490 2184.110 1288.670 ;
        RECT 2182.930 1109.090 2184.110 1110.270 ;
        RECT 2182.930 1107.490 2184.110 1108.670 ;
        RECT 2182.930 929.090 2184.110 930.270 ;
        RECT 2182.930 927.490 2184.110 928.670 ;
        RECT 2182.930 749.090 2184.110 750.270 ;
        RECT 2182.930 747.490 2184.110 748.670 ;
        RECT 2182.930 569.090 2184.110 570.270 ;
        RECT 2182.930 567.490 2184.110 568.670 ;
        RECT 2182.930 389.090 2184.110 390.270 ;
        RECT 2182.930 387.490 2184.110 388.670 ;
        RECT 2182.930 209.090 2184.110 210.270 ;
        RECT 2182.930 207.490 2184.110 208.670 ;
        RECT 2182.930 29.090 2184.110 30.270 ;
        RECT 2182.930 27.490 2184.110 28.670 ;
        RECT 2182.930 -12.310 2184.110 -11.130 ;
        RECT 2182.930 -13.910 2184.110 -12.730 ;
        RECT 2200.930 2747.090 2202.110 2748.270 ;
        RECT 2200.930 2745.490 2202.110 2746.670 ;
        RECT 2200.930 2567.090 2202.110 2568.270 ;
        RECT 2200.930 2565.490 2202.110 2566.670 ;
        RECT 2200.930 2387.090 2202.110 2388.270 ;
        RECT 2200.930 2385.490 2202.110 2386.670 ;
        RECT 2200.930 2207.090 2202.110 2208.270 ;
        RECT 2200.930 2205.490 2202.110 2206.670 ;
        RECT 2200.930 2027.090 2202.110 2028.270 ;
        RECT 2200.930 2025.490 2202.110 2026.670 ;
        RECT 2200.930 1847.090 2202.110 1848.270 ;
        RECT 2200.930 1845.490 2202.110 1846.670 ;
        RECT 2200.930 1667.090 2202.110 1668.270 ;
        RECT 2200.930 1665.490 2202.110 1666.670 ;
        RECT 2200.930 1487.090 2202.110 1488.270 ;
        RECT 2200.930 1485.490 2202.110 1486.670 ;
        RECT 2200.930 1307.090 2202.110 1308.270 ;
        RECT 2200.930 1305.490 2202.110 1306.670 ;
        RECT 2200.930 1127.090 2202.110 1128.270 ;
        RECT 2200.930 1125.490 2202.110 1126.670 ;
        RECT 2200.930 947.090 2202.110 948.270 ;
        RECT 2200.930 945.490 2202.110 946.670 ;
        RECT 2200.930 767.090 2202.110 768.270 ;
        RECT 2200.930 765.490 2202.110 766.670 ;
        RECT 2200.930 587.090 2202.110 588.270 ;
        RECT 2200.930 585.490 2202.110 586.670 ;
        RECT 2200.930 407.090 2202.110 408.270 ;
        RECT 2200.930 405.490 2202.110 406.670 ;
        RECT 2200.930 227.090 2202.110 228.270 ;
        RECT 2200.930 225.490 2202.110 226.670 ;
        RECT 2200.930 47.090 2202.110 48.270 ;
        RECT 2200.930 45.490 2202.110 46.670 ;
        RECT 2200.930 -21.710 2202.110 -20.530 ;
        RECT 2200.930 -23.310 2202.110 -22.130 ;
        RECT 2218.930 2765.090 2220.110 2766.270 ;
        RECT 2218.930 2763.490 2220.110 2764.670 ;
        RECT 2218.930 2585.090 2220.110 2586.270 ;
        RECT 2218.930 2583.490 2220.110 2584.670 ;
        RECT 2218.930 2405.090 2220.110 2406.270 ;
        RECT 2218.930 2403.490 2220.110 2404.670 ;
        RECT 2218.930 2225.090 2220.110 2226.270 ;
        RECT 2218.930 2223.490 2220.110 2224.670 ;
        RECT 2218.930 2045.090 2220.110 2046.270 ;
        RECT 2218.930 2043.490 2220.110 2044.670 ;
        RECT 2218.930 1865.090 2220.110 1866.270 ;
        RECT 2218.930 1863.490 2220.110 1864.670 ;
        RECT 2218.930 1685.090 2220.110 1686.270 ;
        RECT 2218.930 1683.490 2220.110 1684.670 ;
        RECT 2218.930 1505.090 2220.110 1506.270 ;
        RECT 2218.930 1503.490 2220.110 1504.670 ;
        RECT 2218.930 1325.090 2220.110 1326.270 ;
        RECT 2218.930 1323.490 2220.110 1324.670 ;
        RECT 2218.930 1145.090 2220.110 1146.270 ;
        RECT 2218.930 1143.490 2220.110 1144.670 ;
        RECT 2218.930 965.090 2220.110 966.270 ;
        RECT 2218.930 963.490 2220.110 964.670 ;
        RECT 2218.930 785.090 2220.110 786.270 ;
        RECT 2218.930 783.490 2220.110 784.670 ;
        RECT 2218.930 605.090 2220.110 606.270 ;
        RECT 2218.930 603.490 2220.110 604.670 ;
        RECT 2218.930 425.090 2220.110 426.270 ;
        RECT 2218.930 423.490 2220.110 424.670 ;
        RECT 2218.930 245.090 2220.110 246.270 ;
        RECT 2218.930 243.490 2220.110 244.670 ;
        RECT 2218.930 65.090 2220.110 66.270 ;
        RECT 2218.930 63.490 2220.110 64.670 ;
        RECT 2038.930 -31.110 2040.110 -29.930 ;
        RECT 2038.930 -32.710 2040.110 -31.530 ;
        RECT 2344.930 2711.090 2346.110 2712.270 ;
        RECT 2344.930 2709.490 2346.110 2710.670 ;
        RECT 2344.930 2531.090 2346.110 2532.270 ;
        RECT 2344.930 2529.490 2346.110 2530.670 ;
        RECT 2344.930 2351.090 2346.110 2352.270 ;
        RECT 2344.930 2349.490 2346.110 2350.670 ;
        RECT 2344.930 2171.090 2346.110 2172.270 ;
        RECT 2344.930 2169.490 2346.110 2170.670 ;
        RECT 2344.930 1991.090 2346.110 1992.270 ;
        RECT 2344.930 1989.490 2346.110 1990.670 ;
        RECT 2344.930 1811.090 2346.110 1812.270 ;
        RECT 2344.930 1809.490 2346.110 1810.670 ;
        RECT 2344.930 1631.090 2346.110 1632.270 ;
        RECT 2344.930 1629.490 2346.110 1630.670 ;
        RECT 2344.930 1451.090 2346.110 1452.270 ;
        RECT 2344.930 1449.490 2346.110 1450.670 ;
        RECT 2344.930 1271.090 2346.110 1272.270 ;
        RECT 2344.930 1269.490 2346.110 1270.670 ;
        RECT 2344.930 1091.090 2346.110 1092.270 ;
        RECT 2344.930 1089.490 2346.110 1090.670 ;
        RECT 2344.930 911.090 2346.110 912.270 ;
        RECT 2344.930 909.490 2346.110 910.670 ;
        RECT 2344.930 731.090 2346.110 732.270 ;
        RECT 2344.930 729.490 2346.110 730.670 ;
        RECT 2344.930 551.090 2346.110 552.270 ;
        RECT 2344.930 549.490 2346.110 550.670 ;
        RECT 2344.930 371.090 2346.110 372.270 ;
        RECT 2344.930 369.490 2346.110 370.670 ;
        RECT 2344.930 191.090 2346.110 192.270 ;
        RECT 2344.930 189.490 2346.110 190.670 ;
        RECT 2344.930 11.090 2346.110 12.270 ;
        RECT 2344.930 9.490 2346.110 10.670 ;
        RECT 2344.930 -2.910 2346.110 -1.730 ;
        RECT 2344.930 -4.510 2346.110 -3.330 ;
        RECT 2362.930 2729.090 2364.110 2730.270 ;
        RECT 2362.930 2727.490 2364.110 2728.670 ;
        RECT 2362.930 2549.090 2364.110 2550.270 ;
        RECT 2362.930 2547.490 2364.110 2548.670 ;
        RECT 2362.930 2369.090 2364.110 2370.270 ;
        RECT 2362.930 2367.490 2364.110 2368.670 ;
        RECT 2362.930 2189.090 2364.110 2190.270 ;
        RECT 2362.930 2187.490 2364.110 2188.670 ;
        RECT 2362.930 2009.090 2364.110 2010.270 ;
        RECT 2362.930 2007.490 2364.110 2008.670 ;
        RECT 2362.930 1829.090 2364.110 1830.270 ;
        RECT 2362.930 1827.490 2364.110 1828.670 ;
        RECT 2362.930 1649.090 2364.110 1650.270 ;
        RECT 2362.930 1647.490 2364.110 1648.670 ;
        RECT 2362.930 1469.090 2364.110 1470.270 ;
        RECT 2362.930 1467.490 2364.110 1468.670 ;
        RECT 2362.930 1289.090 2364.110 1290.270 ;
        RECT 2362.930 1287.490 2364.110 1288.670 ;
        RECT 2362.930 1109.090 2364.110 1110.270 ;
        RECT 2362.930 1107.490 2364.110 1108.670 ;
        RECT 2362.930 929.090 2364.110 930.270 ;
        RECT 2362.930 927.490 2364.110 928.670 ;
        RECT 2362.930 749.090 2364.110 750.270 ;
        RECT 2362.930 747.490 2364.110 748.670 ;
        RECT 2362.930 569.090 2364.110 570.270 ;
        RECT 2362.930 567.490 2364.110 568.670 ;
        RECT 2362.930 389.090 2364.110 390.270 ;
        RECT 2362.930 387.490 2364.110 388.670 ;
        RECT 2362.930 209.090 2364.110 210.270 ;
        RECT 2362.930 207.490 2364.110 208.670 ;
        RECT 2362.930 29.090 2364.110 30.270 ;
        RECT 2362.930 27.490 2364.110 28.670 ;
        RECT 2362.930 -12.310 2364.110 -11.130 ;
        RECT 2362.930 -13.910 2364.110 -12.730 ;
        RECT 2380.930 2747.090 2382.110 2748.270 ;
        RECT 2380.930 2745.490 2382.110 2746.670 ;
        RECT 2380.930 2567.090 2382.110 2568.270 ;
        RECT 2380.930 2565.490 2382.110 2566.670 ;
        RECT 2380.930 2387.090 2382.110 2388.270 ;
        RECT 2380.930 2385.490 2382.110 2386.670 ;
        RECT 2380.930 2207.090 2382.110 2208.270 ;
        RECT 2380.930 2205.490 2382.110 2206.670 ;
        RECT 2380.930 2027.090 2382.110 2028.270 ;
        RECT 2380.930 2025.490 2382.110 2026.670 ;
        RECT 2380.930 1847.090 2382.110 1848.270 ;
        RECT 2380.930 1845.490 2382.110 1846.670 ;
        RECT 2380.930 1667.090 2382.110 1668.270 ;
        RECT 2380.930 1665.490 2382.110 1666.670 ;
        RECT 2380.930 1487.090 2382.110 1488.270 ;
        RECT 2380.930 1485.490 2382.110 1486.670 ;
        RECT 2380.930 1307.090 2382.110 1308.270 ;
        RECT 2380.930 1305.490 2382.110 1306.670 ;
        RECT 2380.930 1127.090 2382.110 1128.270 ;
        RECT 2380.930 1125.490 2382.110 1126.670 ;
        RECT 2380.930 947.090 2382.110 948.270 ;
        RECT 2380.930 945.490 2382.110 946.670 ;
        RECT 2380.930 767.090 2382.110 768.270 ;
        RECT 2380.930 765.490 2382.110 766.670 ;
        RECT 2380.930 587.090 2382.110 588.270 ;
        RECT 2380.930 585.490 2382.110 586.670 ;
        RECT 2380.930 407.090 2382.110 408.270 ;
        RECT 2380.930 405.490 2382.110 406.670 ;
        RECT 2380.930 227.090 2382.110 228.270 ;
        RECT 2380.930 225.490 2382.110 226.670 ;
        RECT 2380.930 47.090 2382.110 48.270 ;
        RECT 2380.930 45.490 2382.110 46.670 ;
        RECT 2380.930 -21.710 2382.110 -20.530 ;
        RECT 2380.930 -23.310 2382.110 -22.130 ;
        RECT 2398.930 2765.090 2400.110 2766.270 ;
        RECT 2398.930 2763.490 2400.110 2764.670 ;
        RECT 2398.930 2585.090 2400.110 2586.270 ;
        RECT 2398.930 2583.490 2400.110 2584.670 ;
        RECT 2398.930 2405.090 2400.110 2406.270 ;
        RECT 2398.930 2403.490 2400.110 2404.670 ;
        RECT 2398.930 2225.090 2400.110 2226.270 ;
        RECT 2398.930 2223.490 2400.110 2224.670 ;
        RECT 2398.930 2045.090 2400.110 2046.270 ;
        RECT 2398.930 2043.490 2400.110 2044.670 ;
        RECT 2398.930 1865.090 2400.110 1866.270 ;
        RECT 2398.930 1863.490 2400.110 1864.670 ;
        RECT 2398.930 1685.090 2400.110 1686.270 ;
        RECT 2398.930 1683.490 2400.110 1684.670 ;
        RECT 2398.930 1505.090 2400.110 1506.270 ;
        RECT 2398.930 1503.490 2400.110 1504.670 ;
        RECT 2398.930 1325.090 2400.110 1326.270 ;
        RECT 2398.930 1323.490 2400.110 1324.670 ;
        RECT 2398.930 1145.090 2400.110 1146.270 ;
        RECT 2398.930 1143.490 2400.110 1144.670 ;
        RECT 2398.930 965.090 2400.110 966.270 ;
        RECT 2398.930 963.490 2400.110 964.670 ;
        RECT 2398.930 785.090 2400.110 786.270 ;
        RECT 2398.930 783.490 2400.110 784.670 ;
        RECT 2398.930 605.090 2400.110 606.270 ;
        RECT 2398.930 603.490 2400.110 604.670 ;
        RECT 2398.930 425.090 2400.110 426.270 ;
        RECT 2398.930 423.490 2400.110 424.670 ;
        RECT 2398.930 245.090 2400.110 246.270 ;
        RECT 2398.930 243.490 2400.110 244.670 ;
        RECT 2398.930 65.090 2400.110 66.270 ;
        RECT 2398.930 63.490 2400.110 64.670 ;
        RECT 2218.930 -31.110 2220.110 -29.930 ;
        RECT 2218.930 -32.710 2220.110 -31.530 ;
        RECT 2524.930 2711.090 2526.110 2712.270 ;
        RECT 2524.930 2709.490 2526.110 2710.670 ;
        RECT 2524.930 2531.090 2526.110 2532.270 ;
        RECT 2524.930 2529.490 2526.110 2530.670 ;
        RECT 2524.930 2351.090 2526.110 2352.270 ;
        RECT 2524.930 2349.490 2526.110 2350.670 ;
        RECT 2524.930 2171.090 2526.110 2172.270 ;
        RECT 2524.930 2169.490 2526.110 2170.670 ;
        RECT 2524.930 1991.090 2526.110 1992.270 ;
        RECT 2524.930 1989.490 2526.110 1990.670 ;
        RECT 2524.930 1811.090 2526.110 1812.270 ;
        RECT 2524.930 1809.490 2526.110 1810.670 ;
        RECT 2524.930 1631.090 2526.110 1632.270 ;
        RECT 2524.930 1629.490 2526.110 1630.670 ;
        RECT 2524.930 1451.090 2526.110 1452.270 ;
        RECT 2524.930 1449.490 2526.110 1450.670 ;
        RECT 2524.930 1271.090 2526.110 1272.270 ;
        RECT 2524.930 1269.490 2526.110 1270.670 ;
        RECT 2524.930 1091.090 2526.110 1092.270 ;
        RECT 2524.930 1089.490 2526.110 1090.670 ;
        RECT 2524.930 911.090 2526.110 912.270 ;
        RECT 2524.930 909.490 2526.110 910.670 ;
        RECT 2524.930 731.090 2526.110 732.270 ;
        RECT 2524.930 729.490 2526.110 730.670 ;
        RECT 2524.930 551.090 2526.110 552.270 ;
        RECT 2524.930 549.490 2526.110 550.670 ;
        RECT 2524.930 371.090 2526.110 372.270 ;
        RECT 2524.930 369.490 2526.110 370.670 ;
        RECT 2524.930 191.090 2526.110 192.270 ;
        RECT 2524.930 189.490 2526.110 190.670 ;
        RECT 2524.930 11.090 2526.110 12.270 ;
        RECT 2524.930 9.490 2526.110 10.670 ;
        RECT 2524.930 -2.910 2526.110 -1.730 ;
        RECT 2524.930 -4.510 2526.110 -3.330 ;
        RECT 2542.930 2729.090 2544.110 2730.270 ;
        RECT 2542.930 2727.490 2544.110 2728.670 ;
        RECT 2542.930 2549.090 2544.110 2550.270 ;
        RECT 2542.930 2547.490 2544.110 2548.670 ;
        RECT 2542.930 2369.090 2544.110 2370.270 ;
        RECT 2542.930 2367.490 2544.110 2368.670 ;
        RECT 2542.930 2189.090 2544.110 2190.270 ;
        RECT 2542.930 2187.490 2544.110 2188.670 ;
        RECT 2542.930 2009.090 2544.110 2010.270 ;
        RECT 2542.930 2007.490 2544.110 2008.670 ;
        RECT 2542.930 1829.090 2544.110 1830.270 ;
        RECT 2542.930 1827.490 2544.110 1828.670 ;
        RECT 2542.930 1649.090 2544.110 1650.270 ;
        RECT 2542.930 1647.490 2544.110 1648.670 ;
        RECT 2542.930 1469.090 2544.110 1470.270 ;
        RECT 2542.930 1467.490 2544.110 1468.670 ;
        RECT 2542.930 1289.090 2544.110 1290.270 ;
        RECT 2542.930 1287.490 2544.110 1288.670 ;
        RECT 2542.930 1109.090 2544.110 1110.270 ;
        RECT 2542.930 1107.490 2544.110 1108.670 ;
        RECT 2542.930 929.090 2544.110 930.270 ;
        RECT 2542.930 927.490 2544.110 928.670 ;
        RECT 2542.930 749.090 2544.110 750.270 ;
        RECT 2542.930 747.490 2544.110 748.670 ;
        RECT 2542.930 569.090 2544.110 570.270 ;
        RECT 2542.930 567.490 2544.110 568.670 ;
        RECT 2542.930 389.090 2544.110 390.270 ;
        RECT 2542.930 387.490 2544.110 388.670 ;
        RECT 2542.930 209.090 2544.110 210.270 ;
        RECT 2542.930 207.490 2544.110 208.670 ;
        RECT 2542.930 29.090 2544.110 30.270 ;
        RECT 2542.930 27.490 2544.110 28.670 ;
        RECT 2542.930 -12.310 2544.110 -11.130 ;
        RECT 2542.930 -13.910 2544.110 -12.730 ;
        RECT 2560.930 2747.090 2562.110 2748.270 ;
        RECT 2560.930 2745.490 2562.110 2746.670 ;
        RECT 2560.930 2567.090 2562.110 2568.270 ;
        RECT 2560.930 2565.490 2562.110 2566.670 ;
        RECT 2560.930 2387.090 2562.110 2388.270 ;
        RECT 2560.930 2385.490 2562.110 2386.670 ;
        RECT 2560.930 2207.090 2562.110 2208.270 ;
        RECT 2560.930 2205.490 2562.110 2206.670 ;
        RECT 2560.930 2027.090 2562.110 2028.270 ;
        RECT 2560.930 2025.490 2562.110 2026.670 ;
        RECT 2560.930 1847.090 2562.110 1848.270 ;
        RECT 2560.930 1845.490 2562.110 1846.670 ;
        RECT 2560.930 1667.090 2562.110 1668.270 ;
        RECT 2560.930 1665.490 2562.110 1666.670 ;
        RECT 2560.930 1487.090 2562.110 1488.270 ;
        RECT 2560.930 1485.490 2562.110 1486.670 ;
        RECT 2560.930 1307.090 2562.110 1308.270 ;
        RECT 2560.930 1305.490 2562.110 1306.670 ;
        RECT 2560.930 1127.090 2562.110 1128.270 ;
        RECT 2560.930 1125.490 2562.110 1126.670 ;
        RECT 2560.930 947.090 2562.110 948.270 ;
        RECT 2560.930 945.490 2562.110 946.670 ;
        RECT 2560.930 767.090 2562.110 768.270 ;
        RECT 2560.930 765.490 2562.110 766.670 ;
        RECT 2560.930 587.090 2562.110 588.270 ;
        RECT 2560.930 585.490 2562.110 586.670 ;
        RECT 2560.930 407.090 2562.110 408.270 ;
        RECT 2560.930 405.490 2562.110 406.670 ;
        RECT 2560.930 227.090 2562.110 228.270 ;
        RECT 2560.930 225.490 2562.110 226.670 ;
        RECT 2560.930 47.090 2562.110 48.270 ;
        RECT 2560.930 45.490 2562.110 46.670 ;
        RECT 2560.930 -21.710 2562.110 -20.530 ;
        RECT 2560.930 -23.310 2562.110 -22.130 ;
        RECT 2578.930 2765.090 2580.110 2766.270 ;
        RECT 2578.930 2763.490 2580.110 2764.670 ;
        RECT 2578.930 2585.090 2580.110 2586.270 ;
        RECT 2578.930 2583.490 2580.110 2584.670 ;
        RECT 2578.930 2405.090 2580.110 2406.270 ;
        RECT 2578.930 2403.490 2580.110 2404.670 ;
        RECT 2578.930 2225.090 2580.110 2226.270 ;
        RECT 2578.930 2223.490 2580.110 2224.670 ;
        RECT 2578.930 2045.090 2580.110 2046.270 ;
        RECT 2578.930 2043.490 2580.110 2044.670 ;
        RECT 2578.930 1865.090 2580.110 1866.270 ;
        RECT 2578.930 1863.490 2580.110 1864.670 ;
        RECT 2578.930 1685.090 2580.110 1686.270 ;
        RECT 2578.930 1683.490 2580.110 1684.670 ;
        RECT 2578.930 1505.090 2580.110 1506.270 ;
        RECT 2578.930 1503.490 2580.110 1504.670 ;
        RECT 2578.930 1325.090 2580.110 1326.270 ;
        RECT 2578.930 1323.490 2580.110 1324.670 ;
        RECT 2578.930 1145.090 2580.110 1146.270 ;
        RECT 2578.930 1143.490 2580.110 1144.670 ;
        RECT 2578.930 965.090 2580.110 966.270 ;
        RECT 2578.930 963.490 2580.110 964.670 ;
        RECT 2578.930 785.090 2580.110 786.270 ;
        RECT 2578.930 783.490 2580.110 784.670 ;
        RECT 2578.930 605.090 2580.110 606.270 ;
        RECT 2578.930 603.490 2580.110 604.670 ;
        RECT 2578.930 425.090 2580.110 426.270 ;
        RECT 2578.930 423.490 2580.110 424.670 ;
        RECT 2578.930 245.090 2580.110 246.270 ;
        RECT 2578.930 243.490 2580.110 244.670 ;
        RECT 2578.930 65.090 2580.110 66.270 ;
        RECT 2578.930 63.490 2580.110 64.670 ;
        RECT 2398.930 -31.110 2400.110 -29.930 ;
        RECT 2398.930 -32.710 2400.110 -31.530 ;
        RECT 2704.930 2711.090 2706.110 2712.270 ;
        RECT 2704.930 2709.490 2706.110 2710.670 ;
        RECT 2704.930 2531.090 2706.110 2532.270 ;
        RECT 2704.930 2529.490 2706.110 2530.670 ;
        RECT 2704.930 2351.090 2706.110 2352.270 ;
        RECT 2704.930 2349.490 2706.110 2350.670 ;
        RECT 2704.930 2171.090 2706.110 2172.270 ;
        RECT 2704.930 2169.490 2706.110 2170.670 ;
        RECT 2704.930 1991.090 2706.110 1992.270 ;
        RECT 2704.930 1989.490 2706.110 1990.670 ;
        RECT 2704.930 1811.090 2706.110 1812.270 ;
        RECT 2704.930 1809.490 2706.110 1810.670 ;
        RECT 2704.930 1631.090 2706.110 1632.270 ;
        RECT 2704.930 1629.490 2706.110 1630.670 ;
        RECT 2704.930 1451.090 2706.110 1452.270 ;
        RECT 2704.930 1449.490 2706.110 1450.670 ;
        RECT 2704.930 1271.090 2706.110 1272.270 ;
        RECT 2704.930 1269.490 2706.110 1270.670 ;
        RECT 2704.930 1091.090 2706.110 1092.270 ;
        RECT 2704.930 1089.490 2706.110 1090.670 ;
        RECT 2704.930 911.090 2706.110 912.270 ;
        RECT 2704.930 909.490 2706.110 910.670 ;
        RECT 2704.930 731.090 2706.110 732.270 ;
        RECT 2704.930 729.490 2706.110 730.670 ;
        RECT 2704.930 551.090 2706.110 552.270 ;
        RECT 2704.930 549.490 2706.110 550.670 ;
        RECT 2704.930 371.090 2706.110 372.270 ;
        RECT 2704.930 369.490 2706.110 370.670 ;
        RECT 2704.930 191.090 2706.110 192.270 ;
        RECT 2704.930 189.490 2706.110 190.670 ;
        RECT 2704.930 11.090 2706.110 12.270 ;
        RECT 2704.930 9.490 2706.110 10.670 ;
        RECT 2704.930 -2.910 2706.110 -1.730 ;
        RECT 2704.930 -4.510 2706.110 -3.330 ;
        RECT 2722.930 3449.090 2724.110 3450.270 ;
        RECT 2722.930 3447.490 2724.110 3448.670 ;
        RECT 2722.930 3269.090 2724.110 3270.270 ;
        RECT 2722.930 3267.490 2724.110 3268.670 ;
        RECT 2722.930 3089.090 2724.110 3090.270 ;
        RECT 2722.930 3087.490 2724.110 3088.670 ;
        RECT 2722.930 2909.090 2724.110 2910.270 ;
        RECT 2722.930 2907.490 2724.110 2908.670 ;
        RECT 2722.930 2729.090 2724.110 2730.270 ;
        RECT 2722.930 2727.490 2724.110 2728.670 ;
        RECT 2722.930 2549.090 2724.110 2550.270 ;
        RECT 2722.930 2547.490 2724.110 2548.670 ;
        RECT 2722.930 2369.090 2724.110 2370.270 ;
        RECT 2722.930 2367.490 2724.110 2368.670 ;
        RECT 2722.930 2189.090 2724.110 2190.270 ;
        RECT 2722.930 2187.490 2724.110 2188.670 ;
        RECT 2722.930 2009.090 2724.110 2010.270 ;
        RECT 2722.930 2007.490 2724.110 2008.670 ;
        RECT 2722.930 1829.090 2724.110 1830.270 ;
        RECT 2722.930 1827.490 2724.110 1828.670 ;
        RECT 2722.930 1649.090 2724.110 1650.270 ;
        RECT 2722.930 1647.490 2724.110 1648.670 ;
        RECT 2722.930 1469.090 2724.110 1470.270 ;
        RECT 2722.930 1467.490 2724.110 1468.670 ;
        RECT 2722.930 1289.090 2724.110 1290.270 ;
        RECT 2722.930 1287.490 2724.110 1288.670 ;
        RECT 2722.930 1109.090 2724.110 1110.270 ;
        RECT 2722.930 1107.490 2724.110 1108.670 ;
        RECT 2722.930 929.090 2724.110 930.270 ;
        RECT 2722.930 927.490 2724.110 928.670 ;
        RECT 2722.930 749.090 2724.110 750.270 ;
        RECT 2722.930 747.490 2724.110 748.670 ;
        RECT 2722.930 569.090 2724.110 570.270 ;
        RECT 2722.930 567.490 2724.110 568.670 ;
        RECT 2722.930 389.090 2724.110 390.270 ;
        RECT 2722.930 387.490 2724.110 388.670 ;
        RECT 2722.930 209.090 2724.110 210.270 ;
        RECT 2722.930 207.490 2724.110 208.670 ;
        RECT 2722.930 29.090 2724.110 30.270 ;
        RECT 2722.930 27.490 2724.110 28.670 ;
        RECT 2722.930 -12.310 2724.110 -11.130 ;
        RECT 2722.930 -13.910 2724.110 -12.730 ;
        RECT 2740.930 3467.090 2742.110 3468.270 ;
        RECT 2740.930 3465.490 2742.110 3466.670 ;
        RECT 2740.930 3287.090 2742.110 3288.270 ;
        RECT 2740.930 3285.490 2742.110 3286.670 ;
        RECT 2740.930 3107.090 2742.110 3108.270 ;
        RECT 2740.930 3105.490 2742.110 3106.670 ;
        RECT 2740.930 2927.090 2742.110 2928.270 ;
        RECT 2740.930 2925.490 2742.110 2926.670 ;
        RECT 2740.930 2747.090 2742.110 2748.270 ;
        RECT 2740.930 2745.490 2742.110 2746.670 ;
        RECT 2740.930 2567.090 2742.110 2568.270 ;
        RECT 2740.930 2565.490 2742.110 2566.670 ;
        RECT 2740.930 2387.090 2742.110 2388.270 ;
        RECT 2740.930 2385.490 2742.110 2386.670 ;
        RECT 2740.930 2207.090 2742.110 2208.270 ;
        RECT 2740.930 2205.490 2742.110 2206.670 ;
        RECT 2740.930 2027.090 2742.110 2028.270 ;
        RECT 2740.930 2025.490 2742.110 2026.670 ;
        RECT 2740.930 1847.090 2742.110 1848.270 ;
        RECT 2740.930 1845.490 2742.110 1846.670 ;
        RECT 2740.930 1667.090 2742.110 1668.270 ;
        RECT 2740.930 1665.490 2742.110 1666.670 ;
        RECT 2740.930 1487.090 2742.110 1488.270 ;
        RECT 2740.930 1485.490 2742.110 1486.670 ;
        RECT 2740.930 1307.090 2742.110 1308.270 ;
        RECT 2740.930 1305.490 2742.110 1306.670 ;
        RECT 2740.930 1127.090 2742.110 1128.270 ;
        RECT 2740.930 1125.490 2742.110 1126.670 ;
        RECT 2740.930 947.090 2742.110 948.270 ;
        RECT 2740.930 945.490 2742.110 946.670 ;
        RECT 2740.930 767.090 2742.110 768.270 ;
        RECT 2740.930 765.490 2742.110 766.670 ;
        RECT 2740.930 587.090 2742.110 588.270 ;
        RECT 2740.930 585.490 2742.110 586.670 ;
        RECT 2740.930 407.090 2742.110 408.270 ;
        RECT 2740.930 405.490 2742.110 406.670 ;
        RECT 2740.930 227.090 2742.110 228.270 ;
        RECT 2740.930 225.490 2742.110 226.670 ;
        RECT 2740.930 47.090 2742.110 48.270 ;
        RECT 2740.930 45.490 2742.110 46.670 ;
        RECT 2740.930 -21.710 2742.110 -20.530 ;
        RECT 2740.930 -23.310 2742.110 -22.130 ;
        RECT 2955.710 3551.210 2956.890 3552.390 ;
        RECT 2955.710 3549.610 2956.890 3550.790 ;
        RECT 2946.310 3541.810 2947.490 3542.990 ;
        RECT 2946.310 3540.210 2947.490 3541.390 ;
        RECT 2902.930 3532.410 2904.110 3533.590 ;
        RECT 2902.930 3530.810 2904.110 3531.990 ;
        RECT 2758.930 3485.090 2760.110 3486.270 ;
        RECT 2758.930 3483.490 2760.110 3484.670 ;
        RECT 2758.930 3305.090 2760.110 3306.270 ;
        RECT 2758.930 3303.490 2760.110 3304.670 ;
        RECT 2758.930 3125.090 2760.110 3126.270 ;
        RECT 2758.930 3123.490 2760.110 3124.670 ;
        RECT 2758.930 2945.090 2760.110 2946.270 ;
        RECT 2758.930 2943.490 2760.110 2944.670 ;
        RECT 2758.930 2765.090 2760.110 2766.270 ;
        RECT 2758.930 2763.490 2760.110 2764.670 ;
        RECT 2758.930 2585.090 2760.110 2586.270 ;
        RECT 2758.930 2583.490 2760.110 2584.670 ;
        RECT 2758.930 2405.090 2760.110 2406.270 ;
        RECT 2758.930 2403.490 2760.110 2404.670 ;
        RECT 2758.930 2225.090 2760.110 2226.270 ;
        RECT 2758.930 2223.490 2760.110 2224.670 ;
        RECT 2758.930 2045.090 2760.110 2046.270 ;
        RECT 2758.930 2043.490 2760.110 2044.670 ;
        RECT 2758.930 1865.090 2760.110 1866.270 ;
        RECT 2758.930 1863.490 2760.110 1864.670 ;
        RECT 2758.930 1685.090 2760.110 1686.270 ;
        RECT 2758.930 1683.490 2760.110 1684.670 ;
        RECT 2758.930 1505.090 2760.110 1506.270 ;
        RECT 2758.930 1503.490 2760.110 1504.670 ;
        RECT 2758.930 1325.090 2760.110 1326.270 ;
        RECT 2758.930 1323.490 2760.110 1324.670 ;
        RECT 2758.930 1145.090 2760.110 1146.270 ;
        RECT 2758.930 1143.490 2760.110 1144.670 ;
        RECT 2758.930 965.090 2760.110 966.270 ;
        RECT 2758.930 963.490 2760.110 964.670 ;
        RECT 2758.930 785.090 2760.110 786.270 ;
        RECT 2758.930 783.490 2760.110 784.670 ;
        RECT 2758.930 605.090 2760.110 606.270 ;
        RECT 2758.930 603.490 2760.110 604.670 ;
        RECT 2758.930 425.090 2760.110 426.270 ;
        RECT 2758.930 423.490 2760.110 424.670 ;
        RECT 2758.930 245.090 2760.110 246.270 ;
        RECT 2758.930 243.490 2760.110 244.670 ;
        RECT 2758.930 65.090 2760.110 66.270 ;
        RECT 2758.930 63.490 2760.110 64.670 ;
        RECT 2578.930 -31.110 2580.110 -29.930 ;
        RECT 2578.930 -32.710 2580.110 -31.530 ;
        RECT 2884.930 3523.010 2886.110 3524.190 ;
        RECT 2884.930 3521.410 2886.110 3522.590 ;
        RECT 2884.930 3431.090 2886.110 3432.270 ;
        RECT 2884.930 3429.490 2886.110 3430.670 ;
        RECT 2884.930 3251.090 2886.110 3252.270 ;
        RECT 2884.930 3249.490 2886.110 3250.670 ;
        RECT 2884.930 3071.090 2886.110 3072.270 ;
        RECT 2884.930 3069.490 2886.110 3070.670 ;
        RECT 2884.930 2891.090 2886.110 2892.270 ;
        RECT 2884.930 2889.490 2886.110 2890.670 ;
        RECT 2884.930 2711.090 2886.110 2712.270 ;
        RECT 2884.930 2709.490 2886.110 2710.670 ;
        RECT 2884.930 2531.090 2886.110 2532.270 ;
        RECT 2884.930 2529.490 2886.110 2530.670 ;
        RECT 2884.930 2351.090 2886.110 2352.270 ;
        RECT 2884.930 2349.490 2886.110 2350.670 ;
        RECT 2884.930 2171.090 2886.110 2172.270 ;
        RECT 2884.930 2169.490 2886.110 2170.670 ;
        RECT 2884.930 1991.090 2886.110 1992.270 ;
        RECT 2884.930 1989.490 2886.110 1990.670 ;
        RECT 2884.930 1811.090 2886.110 1812.270 ;
        RECT 2884.930 1809.490 2886.110 1810.670 ;
        RECT 2884.930 1631.090 2886.110 1632.270 ;
        RECT 2884.930 1629.490 2886.110 1630.670 ;
        RECT 2884.930 1451.090 2886.110 1452.270 ;
        RECT 2884.930 1449.490 2886.110 1450.670 ;
        RECT 2884.930 1271.090 2886.110 1272.270 ;
        RECT 2884.930 1269.490 2886.110 1270.670 ;
        RECT 2884.930 1091.090 2886.110 1092.270 ;
        RECT 2884.930 1089.490 2886.110 1090.670 ;
        RECT 2884.930 911.090 2886.110 912.270 ;
        RECT 2884.930 909.490 2886.110 910.670 ;
        RECT 2884.930 731.090 2886.110 732.270 ;
        RECT 2884.930 729.490 2886.110 730.670 ;
        RECT 2884.930 551.090 2886.110 552.270 ;
        RECT 2884.930 549.490 2886.110 550.670 ;
        RECT 2884.930 371.090 2886.110 372.270 ;
        RECT 2884.930 369.490 2886.110 370.670 ;
        RECT 2884.930 191.090 2886.110 192.270 ;
        RECT 2884.930 189.490 2886.110 190.670 ;
        RECT 2884.930 11.090 2886.110 12.270 ;
        RECT 2884.930 9.490 2886.110 10.670 ;
        RECT 2884.930 -2.910 2886.110 -1.730 ;
        RECT 2884.930 -4.510 2886.110 -3.330 ;
        RECT 2936.910 3532.410 2938.090 3533.590 ;
        RECT 2936.910 3530.810 2938.090 3531.990 ;
        RECT 2902.930 3449.090 2904.110 3450.270 ;
        RECT 2902.930 3447.490 2904.110 3448.670 ;
        RECT 2902.930 3269.090 2904.110 3270.270 ;
        RECT 2902.930 3267.490 2904.110 3268.670 ;
        RECT 2902.930 3089.090 2904.110 3090.270 ;
        RECT 2902.930 3087.490 2904.110 3088.670 ;
        RECT 2902.930 2909.090 2904.110 2910.270 ;
        RECT 2902.930 2907.490 2904.110 2908.670 ;
        RECT 2902.930 2729.090 2904.110 2730.270 ;
        RECT 2902.930 2727.490 2904.110 2728.670 ;
        RECT 2902.930 2549.090 2904.110 2550.270 ;
        RECT 2902.930 2547.490 2904.110 2548.670 ;
        RECT 2902.930 2369.090 2904.110 2370.270 ;
        RECT 2902.930 2367.490 2904.110 2368.670 ;
        RECT 2902.930 2189.090 2904.110 2190.270 ;
        RECT 2902.930 2187.490 2904.110 2188.670 ;
        RECT 2902.930 2009.090 2904.110 2010.270 ;
        RECT 2902.930 2007.490 2904.110 2008.670 ;
        RECT 2902.930 1829.090 2904.110 1830.270 ;
        RECT 2902.930 1827.490 2904.110 1828.670 ;
        RECT 2902.930 1649.090 2904.110 1650.270 ;
        RECT 2902.930 1647.490 2904.110 1648.670 ;
        RECT 2902.930 1469.090 2904.110 1470.270 ;
        RECT 2902.930 1467.490 2904.110 1468.670 ;
        RECT 2902.930 1289.090 2904.110 1290.270 ;
        RECT 2902.930 1287.490 2904.110 1288.670 ;
        RECT 2902.930 1109.090 2904.110 1110.270 ;
        RECT 2902.930 1107.490 2904.110 1108.670 ;
        RECT 2902.930 929.090 2904.110 930.270 ;
        RECT 2902.930 927.490 2904.110 928.670 ;
        RECT 2902.930 749.090 2904.110 750.270 ;
        RECT 2902.930 747.490 2904.110 748.670 ;
        RECT 2902.930 569.090 2904.110 570.270 ;
        RECT 2902.930 567.490 2904.110 568.670 ;
        RECT 2902.930 389.090 2904.110 390.270 ;
        RECT 2902.930 387.490 2904.110 388.670 ;
        RECT 2902.930 209.090 2904.110 210.270 ;
        RECT 2902.930 207.490 2904.110 208.670 ;
        RECT 2902.930 29.090 2904.110 30.270 ;
        RECT 2902.930 27.490 2904.110 28.670 ;
        RECT 2927.510 3523.010 2928.690 3524.190 ;
        RECT 2927.510 3521.410 2928.690 3522.590 ;
        RECT 2927.510 3431.090 2928.690 3432.270 ;
        RECT 2927.510 3429.490 2928.690 3430.670 ;
        RECT 2927.510 3251.090 2928.690 3252.270 ;
        RECT 2927.510 3249.490 2928.690 3250.670 ;
        RECT 2927.510 3071.090 2928.690 3072.270 ;
        RECT 2927.510 3069.490 2928.690 3070.670 ;
        RECT 2927.510 2891.090 2928.690 2892.270 ;
        RECT 2927.510 2889.490 2928.690 2890.670 ;
        RECT 2927.510 2711.090 2928.690 2712.270 ;
        RECT 2927.510 2709.490 2928.690 2710.670 ;
        RECT 2927.510 2531.090 2928.690 2532.270 ;
        RECT 2927.510 2529.490 2928.690 2530.670 ;
        RECT 2927.510 2351.090 2928.690 2352.270 ;
        RECT 2927.510 2349.490 2928.690 2350.670 ;
        RECT 2927.510 2171.090 2928.690 2172.270 ;
        RECT 2927.510 2169.490 2928.690 2170.670 ;
        RECT 2927.510 1991.090 2928.690 1992.270 ;
        RECT 2927.510 1989.490 2928.690 1990.670 ;
        RECT 2927.510 1811.090 2928.690 1812.270 ;
        RECT 2927.510 1809.490 2928.690 1810.670 ;
        RECT 2927.510 1631.090 2928.690 1632.270 ;
        RECT 2927.510 1629.490 2928.690 1630.670 ;
        RECT 2927.510 1451.090 2928.690 1452.270 ;
        RECT 2927.510 1449.490 2928.690 1450.670 ;
        RECT 2927.510 1271.090 2928.690 1272.270 ;
        RECT 2927.510 1269.490 2928.690 1270.670 ;
        RECT 2927.510 1091.090 2928.690 1092.270 ;
        RECT 2927.510 1089.490 2928.690 1090.670 ;
        RECT 2927.510 911.090 2928.690 912.270 ;
        RECT 2927.510 909.490 2928.690 910.670 ;
        RECT 2927.510 731.090 2928.690 732.270 ;
        RECT 2927.510 729.490 2928.690 730.670 ;
        RECT 2927.510 551.090 2928.690 552.270 ;
        RECT 2927.510 549.490 2928.690 550.670 ;
        RECT 2927.510 371.090 2928.690 372.270 ;
        RECT 2927.510 369.490 2928.690 370.670 ;
        RECT 2927.510 191.090 2928.690 192.270 ;
        RECT 2927.510 189.490 2928.690 190.670 ;
        RECT 2927.510 11.090 2928.690 12.270 ;
        RECT 2927.510 9.490 2928.690 10.670 ;
        RECT 2927.510 -2.910 2928.690 -1.730 ;
        RECT 2927.510 -4.510 2928.690 -3.330 ;
        RECT 2936.910 3449.090 2938.090 3450.270 ;
        RECT 2936.910 3447.490 2938.090 3448.670 ;
        RECT 2936.910 3269.090 2938.090 3270.270 ;
        RECT 2936.910 3267.490 2938.090 3268.670 ;
        RECT 2936.910 3089.090 2938.090 3090.270 ;
        RECT 2936.910 3087.490 2938.090 3088.670 ;
        RECT 2936.910 2909.090 2938.090 2910.270 ;
        RECT 2936.910 2907.490 2938.090 2908.670 ;
        RECT 2936.910 2729.090 2938.090 2730.270 ;
        RECT 2936.910 2727.490 2938.090 2728.670 ;
        RECT 2936.910 2549.090 2938.090 2550.270 ;
        RECT 2936.910 2547.490 2938.090 2548.670 ;
        RECT 2936.910 2369.090 2938.090 2370.270 ;
        RECT 2936.910 2367.490 2938.090 2368.670 ;
        RECT 2936.910 2189.090 2938.090 2190.270 ;
        RECT 2936.910 2187.490 2938.090 2188.670 ;
        RECT 2936.910 2009.090 2938.090 2010.270 ;
        RECT 2936.910 2007.490 2938.090 2008.670 ;
        RECT 2936.910 1829.090 2938.090 1830.270 ;
        RECT 2936.910 1827.490 2938.090 1828.670 ;
        RECT 2936.910 1649.090 2938.090 1650.270 ;
        RECT 2936.910 1647.490 2938.090 1648.670 ;
        RECT 2936.910 1469.090 2938.090 1470.270 ;
        RECT 2936.910 1467.490 2938.090 1468.670 ;
        RECT 2936.910 1289.090 2938.090 1290.270 ;
        RECT 2936.910 1287.490 2938.090 1288.670 ;
        RECT 2936.910 1109.090 2938.090 1110.270 ;
        RECT 2936.910 1107.490 2938.090 1108.670 ;
        RECT 2936.910 929.090 2938.090 930.270 ;
        RECT 2936.910 927.490 2938.090 928.670 ;
        RECT 2936.910 749.090 2938.090 750.270 ;
        RECT 2936.910 747.490 2938.090 748.670 ;
        RECT 2936.910 569.090 2938.090 570.270 ;
        RECT 2936.910 567.490 2938.090 568.670 ;
        RECT 2936.910 389.090 2938.090 390.270 ;
        RECT 2936.910 387.490 2938.090 388.670 ;
        RECT 2936.910 209.090 2938.090 210.270 ;
        RECT 2936.910 207.490 2938.090 208.670 ;
        RECT 2936.910 29.090 2938.090 30.270 ;
        RECT 2936.910 27.490 2938.090 28.670 ;
        RECT 2902.930 -12.310 2904.110 -11.130 ;
        RECT 2902.930 -13.910 2904.110 -12.730 ;
        RECT 2936.910 -12.310 2938.090 -11.130 ;
        RECT 2936.910 -13.910 2938.090 -12.730 ;
        RECT 2946.310 3467.090 2947.490 3468.270 ;
        RECT 2946.310 3465.490 2947.490 3466.670 ;
        RECT 2946.310 3287.090 2947.490 3288.270 ;
        RECT 2946.310 3285.490 2947.490 3286.670 ;
        RECT 2946.310 3107.090 2947.490 3108.270 ;
        RECT 2946.310 3105.490 2947.490 3106.670 ;
        RECT 2946.310 2927.090 2947.490 2928.270 ;
        RECT 2946.310 2925.490 2947.490 2926.670 ;
        RECT 2946.310 2747.090 2947.490 2748.270 ;
        RECT 2946.310 2745.490 2947.490 2746.670 ;
        RECT 2946.310 2567.090 2947.490 2568.270 ;
        RECT 2946.310 2565.490 2947.490 2566.670 ;
        RECT 2946.310 2387.090 2947.490 2388.270 ;
        RECT 2946.310 2385.490 2947.490 2386.670 ;
        RECT 2946.310 2207.090 2947.490 2208.270 ;
        RECT 2946.310 2205.490 2947.490 2206.670 ;
        RECT 2946.310 2027.090 2947.490 2028.270 ;
        RECT 2946.310 2025.490 2947.490 2026.670 ;
        RECT 2946.310 1847.090 2947.490 1848.270 ;
        RECT 2946.310 1845.490 2947.490 1846.670 ;
        RECT 2946.310 1667.090 2947.490 1668.270 ;
        RECT 2946.310 1665.490 2947.490 1666.670 ;
        RECT 2946.310 1487.090 2947.490 1488.270 ;
        RECT 2946.310 1485.490 2947.490 1486.670 ;
        RECT 2946.310 1307.090 2947.490 1308.270 ;
        RECT 2946.310 1305.490 2947.490 1306.670 ;
        RECT 2946.310 1127.090 2947.490 1128.270 ;
        RECT 2946.310 1125.490 2947.490 1126.670 ;
        RECT 2946.310 947.090 2947.490 948.270 ;
        RECT 2946.310 945.490 2947.490 946.670 ;
        RECT 2946.310 767.090 2947.490 768.270 ;
        RECT 2946.310 765.490 2947.490 766.670 ;
        RECT 2946.310 587.090 2947.490 588.270 ;
        RECT 2946.310 585.490 2947.490 586.670 ;
        RECT 2946.310 407.090 2947.490 408.270 ;
        RECT 2946.310 405.490 2947.490 406.670 ;
        RECT 2946.310 227.090 2947.490 228.270 ;
        RECT 2946.310 225.490 2947.490 226.670 ;
        RECT 2946.310 47.090 2947.490 48.270 ;
        RECT 2946.310 45.490 2947.490 46.670 ;
        RECT 2946.310 -21.710 2947.490 -20.530 ;
        RECT 2946.310 -23.310 2947.490 -22.130 ;
        RECT 2955.710 3485.090 2956.890 3486.270 ;
        RECT 2955.710 3483.490 2956.890 3484.670 ;
        RECT 2955.710 3305.090 2956.890 3306.270 ;
        RECT 2955.710 3303.490 2956.890 3304.670 ;
        RECT 2955.710 3125.090 2956.890 3126.270 ;
        RECT 2955.710 3123.490 2956.890 3124.670 ;
        RECT 2955.710 2945.090 2956.890 2946.270 ;
        RECT 2955.710 2943.490 2956.890 2944.670 ;
        RECT 2955.710 2765.090 2956.890 2766.270 ;
        RECT 2955.710 2763.490 2956.890 2764.670 ;
        RECT 2955.710 2585.090 2956.890 2586.270 ;
        RECT 2955.710 2583.490 2956.890 2584.670 ;
        RECT 2955.710 2405.090 2956.890 2406.270 ;
        RECT 2955.710 2403.490 2956.890 2404.670 ;
        RECT 2955.710 2225.090 2956.890 2226.270 ;
        RECT 2955.710 2223.490 2956.890 2224.670 ;
        RECT 2955.710 2045.090 2956.890 2046.270 ;
        RECT 2955.710 2043.490 2956.890 2044.670 ;
        RECT 2955.710 1865.090 2956.890 1866.270 ;
        RECT 2955.710 1863.490 2956.890 1864.670 ;
        RECT 2955.710 1685.090 2956.890 1686.270 ;
        RECT 2955.710 1683.490 2956.890 1684.670 ;
        RECT 2955.710 1505.090 2956.890 1506.270 ;
        RECT 2955.710 1503.490 2956.890 1504.670 ;
        RECT 2955.710 1325.090 2956.890 1326.270 ;
        RECT 2955.710 1323.490 2956.890 1324.670 ;
        RECT 2955.710 1145.090 2956.890 1146.270 ;
        RECT 2955.710 1143.490 2956.890 1144.670 ;
        RECT 2955.710 965.090 2956.890 966.270 ;
        RECT 2955.710 963.490 2956.890 964.670 ;
        RECT 2955.710 785.090 2956.890 786.270 ;
        RECT 2955.710 783.490 2956.890 784.670 ;
        RECT 2955.710 605.090 2956.890 606.270 ;
        RECT 2955.710 603.490 2956.890 604.670 ;
        RECT 2955.710 425.090 2956.890 426.270 ;
        RECT 2955.710 423.490 2956.890 424.670 ;
        RECT 2955.710 245.090 2956.890 246.270 ;
        RECT 2955.710 243.490 2956.890 244.670 ;
        RECT 2955.710 65.090 2956.890 66.270 ;
        RECT 2955.710 63.490 2956.890 64.670 ;
        RECT 2758.930 -31.110 2760.110 -29.930 ;
        RECT 2758.930 -32.710 2760.110 -31.530 ;
        RECT 2955.710 -31.110 2956.890 -29.930 ;
        RECT 2955.710 -32.710 2956.890 -31.530 ;
      LAYER met5 ;
        RECT -38.180 3552.500 -35.180 3552.510 ;
        RECT 58.020 3552.500 61.020 3552.510 ;
        RECT 238.020 3552.500 241.020 3552.510 ;
        RECT 418.020 3552.500 421.020 3552.510 ;
        RECT 598.020 3552.500 601.020 3552.510 ;
        RECT 778.020 3552.500 781.020 3552.510 ;
        RECT 958.020 3552.500 961.020 3552.510 ;
        RECT 1138.020 3552.500 1141.020 3552.510 ;
        RECT 1318.020 3552.500 1321.020 3552.510 ;
        RECT 1498.020 3552.500 1501.020 3552.510 ;
        RECT 1678.020 3552.500 1681.020 3552.510 ;
        RECT 1858.020 3552.500 1861.020 3552.510 ;
        RECT 2038.020 3552.500 2041.020 3552.510 ;
        RECT 2218.020 3552.500 2221.020 3552.510 ;
        RECT 2398.020 3552.500 2401.020 3552.510 ;
        RECT 2578.020 3552.500 2581.020 3552.510 ;
        RECT 2758.020 3552.500 2761.020 3552.510 ;
        RECT 2954.800 3552.500 2957.800 3552.510 ;
        RECT -38.180 3549.500 2957.800 3552.500 ;
        RECT -38.180 3549.490 -35.180 3549.500 ;
        RECT 58.020 3549.490 61.020 3549.500 ;
        RECT 238.020 3549.490 241.020 3549.500 ;
        RECT 418.020 3549.490 421.020 3549.500 ;
        RECT 598.020 3549.490 601.020 3549.500 ;
        RECT 778.020 3549.490 781.020 3549.500 ;
        RECT 958.020 3549.490 961.020 3549.500 ;
        RECT 1138.020 3549.490 1141.020 3549.500 ;
        RECT 1318.020 3549.490 1321.020 3549.500 ;
        RECT 1498.020 3549.490 1501.020 3549.500 ;
        RECT 1678.020 3549.490 1681.020 3549.500 ;
        RECT 1858.020 3549.490 1861.020 3549.500 ;
        RECT 2038.020 3549.490 2041.020 3549.500 ;
        RECT 2218.020 3549.490 2221.020 3549.500 ;
        RECT 2398.020 3549.490 2401.020 3549.500 ;
        RECT 2578.020 3549.490 2581.020 3549.500 ;
        RECT 2758.020 3549.490 2761.020 3549.500 ;
        RECT 2954.800 3549.490 2957.800 3549.500 ;
        RECT -28.780 3543.100 -25.780 3543.110 ;
        RECT 40.020 3543.100 43.020 3543.110 ;
        RECT 220.020 3543.100 223.020 3543.110 ;
        RECT 400.020 3543.100 403.020 3543.110 ;
        RECT 580.020 3543.100 583.020 3543.110 ;
        RECT 760.020 3543.100 763.020 3543.110 ;
        RECT 940.020 3543.100 943.020 3543.110 ;
        RECT 1120.020 3543.100 1123.020 3543.110 ;
        RECT 1300.020 3543.100 1303.020 3543.110 ;
        RECT 1480.020 3543.100 1483.020 3543.110 ;
        RECT 1660.020 3543.100 1663.020 3543.110 ;
        RECT 1840.020 3543.100 1843.020 3543.110 ;
        RECT 2020.020 3543.100 2023.020 3543.110 ;
        RECT 2200.020 3543.100 2203.020 3543.110 ;
        RECT 2380.020 3543.100 2383.020 3543.110 ;
        RECT 2560.020 3543.100 2563.020 3543.110 ;
        RECT 2740.020 3543.100 2743.020 3543.110 ;
        RECT 2945.400 3543.100 2948.400 3543.110 ;
        RECT -28.780 3540.100 2948.400 3543.100 ;
        RECT -28.780 3540.090 -25.780 3540.100 ;
        RECT 40.020 3540.090 43.020 3540.100 ;
        RECT 220.020 3540.090 223.020 3540.100 ;
        RECT 400.020 3540.090 403.020 3540.100 ;
        RECT 580.020 3540.090 583.020 3540.100 ;
        RECT 760.020 3540.090 763.020 3540.100 ;
        RECT 940.020 3540.090 943.020 3540.100 ;
        RECT 1120.020 3540.090 1123.020 3540.100 ;
        RECT 1300.020 3540.090 1303.020 3540.100 ;
        RECT 1480.020 3540.090 1483.020 3540.100 ;
        RECT 1660.020 3540.090 1663.020 3540.100 ;
        RECT 1840.020 3540.090 1843.020 3540.100 ;
        RECT 2020.020 3540.090 2023.020 3540.100 ;
        RECT 2200.020 3540.090 2203.020 3540.100 ;
        RECT 2380.020 3540.090 2383.020 3540.100 ;
        RECT 2560.020 3540.090 2563.020 3540.100 ;
        RECT 2740.020 3540.090 2743.020 3540.100 ;
        RECT 2945.400 3540.090 2948.400 3540.100 ;
        RECT -19.380 3533.700 -16.380 3533.710 ;
        RECT 22.020 3533.700 25.020 3533.710 ;
        RECT 202.020 3533.700 205.020 3533.710 ;
        RECT 382.020 3533.700 385.020 3533.710 ;
        RECT 562.020 3533.700 565.020 3533.710 ;
        RECT 742.020 3533.700 745.020 3533.710 ;
        RECT 922.020 3533.700 925.020 3533.710 ;
        RECT 1102.020 3533.700 1105.020 3533.710 ;
        RECT 1282.020 3533.700 1285.020 3533.710 ;
        RECT 1462.020 3533.700 1465.020 3533.710 ;
        RECT 1642.020 3533.700 1645.020 3533.710 ;
        RECT 1822.020 3533.700 1825.020 3533.710 ;
        RECT 2002.020 3533.700 2005.020 3533.710 ;
        RECT 2182.020 3533.700 2185.020 3533.710 ;
        RECT 2362.020 3533.700 2365.020 3533.710 ;
        RECT 2542.020 3533.700 2545.020 3533.710 ;
        RECT 2722.020 3533.700 2725.020 3533.710 ;
        RECT 2902.020 3533.700 2905.020 3533.710 ;
        RECT 2936.000 3533.700 2939.000 3533.710 ;
        RECT -19.380 3530.700 2939.000 3533.700 ;
        RECT -19.380 3530.690 -16.380 3530.700 ;
        RECT 22.020 3530.690 25.020 3530.700 ;
        RECT 202.020 3530.690 205.020 3530.700 ;
        RECT 382.020 3530.690 385.020 3530.700 ;
        RECT 562.020 3530.690 565.020 3530.700 ;
        RECT 742.020 3530.690 745.020 3530.700 ;
        RECT 922.020 3530.690 925.020 3530.700 ;
        RECT 1102.020 3530.690 1105.020 3530.700 ;
        RECT 1282.020 3530.690 1285.020 3530.700 ;
        RECT 1462.020 3530.690 1465.020 3530.700 ;
        RECT 1642.020 3530.690 1645.020 3530.700 ;
        RECT 1822.020 3530.690 1825.020 3530.700 ;
        RECT 2002.020 3530.690 2005.020 3530.700 ;
        RECT 2182.020 3530.690 2185.020 3530.700 ;
        RECT 2362.020 3530.690 2365.020 3530.700 ;
        RECT 2542.020 3530.690 2545.020 3530.700 ;
        RECT 2722.020 3530.690 2725.020 3530.700 ;
        RECT 2902.020 3530.690 2905.020 3530.700 ;
        RECT 2936.000 3530.690 2939.000 3530.700 ;
        RECT -9.980 3524.300 -6.980 3524.310 ;
        RECT 4.020 3524.300 7.020 3524.310 ;
        RECT 184.020 3524.300 187.020 3524.310 ;
        RECT 364.020 3524.300 367.020 3524.310 ;
        RECT 544.020 3524.300 547.020 3524.310 ;
        RECT 724.020 3524.300 727.020 3524.310 ;
        RECT 904.020 3524.300 907.020 3524.310 ;
        RECT 1084.020 3524.300 1087.020 3524.310 ;
        RECT 1264.020 3524.300 1267.020 3524.310 ;
        RECT 1444.020 3524.300 1447.020 3524.310 ;
        RECT 1624.020 3524.300 1627.020 3524.310 ;
        RECT 1804.020 3524.300 1807.020 3524.310 ;
        RECT 1984.020 3524.300 1987.020 3524.310 ;
        RECT 2164.020 3524.300 2167.020 3524.310 ;
        RECT 2344.020 3524.300 2347.020 3524.310 ;
        RECT 2524.020 3524.300 2527.020 3524.310 ;
        RECT 2704.020 3524.300 2707.020 3524.310 ;
        RECT 2884.020 3524.300 2887.020 3524.310 ;
        RECT 2926.600 3524.300 2929.600 3524.310 ;
        RECT -9.980 3521.300 2929.600 3524.300 ;
        RECT -9.980 3521.290 -6.980 3521.300 ;
        RECT 4.020 3521.290 7.020 3521.300 ;
        RECT 184.020 3521.290 187.020 3521.300 ;
        RECT 364.020 3521.290 367.020 3521.300 ;
        RECT 544.020 3521.290 547.020 3521.300 ;
        RECT 724.020 3521.290 727.020 3521.300 ;
        RECT 904.020 3521.290 907.020 3521.300 ;
        RECT 1084.020 3521.290 1087.020 3521.300 ;
        RECT 1264.020 3521.290 1267.020 3521.300 ;
        RECT 1444.020 3521.290 1447.020 3521.300 ;
        RECT 1624.020 3521.290 1627.020 3521.300 ;
        RECT 1804.020 3521.290 1807.020 3521.300 ;
        RECT 1984.020 3521.290 1987.020 3521.300 ;
        RECT 2164.020 3521.290 2167.020 3521.300 ;
        RECT 2344.020 3521.290 2347.020 3521.300 ;
        RECT 2524.020 3521.290 2527.020 3521.300 ;
        RECT 2704.020 3521.290 2707.020 3521.300 ;
        RECT 2884.020 3521.290 2887.020 3521.300 ;
        RECT 2926.600 3521.290 2929.600 3521.300 ;
        RECT -38.180 3486.380 -35.180 3486.390 ;
        RECT 58.020 3486.380 61.020 3486.390 ;
        RECT 238.020 3486.380 241.020 3486.390 ;
        RECT 418.020 3486.380 421.020 3486.390 ;
        RECT 598.020 3486.380 601.020 3486.390 ;
        RECT 778.020 3486.380 781.020 3486.390 ;
        RECT 958.020 3486.380 961.020 3486.390 ;
        RECT 1138.020 3486.380 1141.020 3486.390 ;
        RECT 1318.020 3486.380 1321.020 3486.390 ;
        RECT 1498.020 3486.380 1501.020 3486.390 ;
        RECT 1678.020 3486.380 1681.020 3486.390 ;
        RECT 1858.020 3486.380 1861.020 3486.390 ;
        RECT 2038.020 3486.380 2041.020 3486.390 ;
        RECT 2218.020 3486.380 2221.020 3486.390 ;
        RECT 2398.020 3486.380 2401.020 3486.390 ;
        RECT 2578.020 3486.380 2581.020 3486.390 ;
        RECT 2758.020 3486.380 2761.020 3486.390 ;
        RECT 2954.800 3486.380 2957.800 3486.390 ;
        RECT -42.880 3483.380 2962.500 3486.380 ;
        RECT -38.180 3483.370 -35.180 3483.380 ;
        RECT 58.020 3483.370 61.020 3483.380 ;
        RECT 238.020 3483.370 241.020 3483.380 ;
        RECT 418.020 3483.370 421.020 3483.380 ;
        RECT 598.020 3483.370 601.020 3483.380 ;
        RECT 778.020 3483.370 781.020 3483.380 ;
        RECT 958.020 3483.370 961.020 3483.380 ;
        RECT 1138.020 3483.370 1141.020 3483.380 ;
        RECT 1318.020 3483.370 1321.020 3483.380 ;
        RECT 1498.020 3483.370 1501.020 3483.380 ;
        RECT 1678.020 3483.370 1681.020 3483.380 ;
        RECT 1858.020 3483.370 1861.020 3483.380 ;
        RECT 2038.020 3483.370 2041.020 3483.380 ;
        RECT 2218.020 3483.370 2221.020 3483.380 ;
        RECT 2398.020 3483.370 2401.020 3483.380 ;
        RECT 2578.020 3483.370 2581.020 3483.380 ;
        RECT 2758.020 3483.370 2761.020 3483.380 ;
        RECT 2954.800 3483.370 2957.800 3483.380 ;
        RECT -28.780 3468.380 -25.780 3468.390 ;
        RECT 40.020 3468.380 43.020 3468.390 ;
        RECT 220.020 3468.380 223.020 3468.390 ;
        RECT 400.020 3468.380 403.020 3468.390 ;
        RECT 580.020 3468.380 583.020 3468.390 ;
        RECT 760.020 3468.380 763.020 3468.390 ;
        RECT 940.020 3468.380 943.020 3468.390 ;
        RECT 1120.020 3468.380 1123.020 3468.390 ;
        RECT 1300.020 3468.380 1303.020 3468.390 ;
        RECT 1480.020 3468.380 1483.020 3468.390 ;
        RECT 1660.020 3468.380 1663.020 3468.390 ;
        RECT 1840.020 3468.380 1843.020 3468.390 ;
        RECT 2020.020 3468.380 2023.020 3468.390 ;
        RECT 2200.020 3468.380 2203.020 3468.390 ;
        RECT 2380.020 3468.380 2383.020 3468.390 ;
        RECT 2560.020 3468.380 2563.020 3468.390 ;
        RECT 2740.020 3468.380 2743.020 3468.390 ;
        RECT 2945.400 3468.380 2948.400 3468.390 ;
        RECT -33.480 3465.380 2953.100 3468.380 ;
        RECT -28.780 3465.370 -25.780 3465.380 ;
        RECT 40.020 3465.370 43.020 3465.380 ;
        RECT 220.020 3465.370 223.020 3465.380 ;
        RECT 400.020 3465.370 403.020 3465.380 ;
        RECT 580.020 3465.370 583.020 3465.380 ;
        RECT 760.020 3465.370 763.020 3465.380 ;
        RECT 940.020 3465.370 943.020 3465.380 ;
        RECT 1120.020 3465.370 1123.020 3465.380 ;
        RECT 1300.020 3465.370 1303.020 3465.380 ;
        RECT 1480.020 3465.370 1483.020 3465.380 ;
        RECT 1660.020 3465.370 1663.020 3465.380 ;
        RECT 1840.020 3465.370 1843.020 3465.380 ;
        RECT 2020.020 3465.370 2023.020 3465.380 ;
        RECT 2200.020 3465.370 2203.020 3465.380 ;
        RECT 2380.020 3465.370 2383.020 3465.380 ;
        RECT 2560.020 3465.370 2563.020 3465.380 ;
        RECT 2740.020 3465.370 2743.020 3465.380 ;
        RECT 2945.400 3465.370 2948.400 3465.380 ;
        RECT -19.380 3450.380 -16.380 3450.390 ;
        RECT 22.020 3450.380 25.020 3450.390 ;
        RECT 202.020 3450.380 205.020 3450.390 ;
        RECT 382.020 3450.380 385.020 3450.390 ;
        RECT 562.020 3450.380 565.020 3450.390 ;
        RECT 742.020 3450.380 745.020 3450.390 ;
        RECT 922.020 3450.380 925.020 3450.390 ;
        RECT 1102.020 3450.380 1105.020 3450.390 ;
        RECT 1282.020 3450.380 1285.020 3450.390 ;
        RECT 1462.020 3450.380 1465.020 3450.390 ;
        RECT 1642.020 3450.380 1645.020 3450.390 ;
        RECT 1822.020 3450.380 1825.020 3450.390 ;
        RECT 2002.020 3450.380 2005.020 3450.390 ;
        RECT 2182.020 3450.380 2185.020 3450.390 ;
        RECT 2362.020 3450.380 2365.020 3450.390 ;
        RECT 2542.020 3450.380 2545.020 3450.390 ;
        RECT 2722.020 3450.380 2725.020 3450.390 ;
        RECT 2902.020 3450.380 2905.020 3450.390 ;
        RECT 2936.000 3450.380 2939.000 3450.390 ;
        RECT -24.080 3447.380 2943.700 3450.380 ;
        RECT -19.380 3447.370 -16.380 3447.380 ;
        RECT 22.020 3447.370 25.020 3447.380 ;
        RECT 202.020 3447.370 205.020 3447.380 ;
        RECT 382.020 3447.370 385.020 3447.380 ;
        RECT 562.020 3447.370 565.020 3447.380 ;
        RECT 742.020 3447.370 745.020 3447.380 ;
        RECT 922.020 3447.370 925.020 3447.380 ;
        RECT 1102.020 3447.370 1105.020 3447.380 ;
        RECT 1282.020 3447.370 1285.020 3447.380 ;
        RECT 1462.020 3447.370 1465.020 3447.380 ;
        RECT 1642.020 3447.370 1645.020 3447.380 ;
        RECT 1822.020 3447.370 1825.020 3447.380 ;
        RECT 2002.020 3447.370 2005.020 3447.380 ;
        RECT 2182.020 3447.370 2185.020 3447.380 ;
        RECT 2362.020 3447.370 2365.020 3447.380 ;
        RECT 2542.020 3447.370 2545.020 3447.380 ;
        RECT 2722.020 3447.370 2725.020 3447.380 ;
        RECT 2902.020 3447.370 2905.020 3447.380 ;
        RECT 2936.000 3447.370 2939.000 3447.380 ;
        RECT -9.980 3432.380 -6.980 3432.390 ;
        RECT 4.020 3432.380 7.020 3432.390 ;
        RECT 184.020 3432.380 187.020 3432.390 ;
        RECT 364.020 3432.380 367.020 3432.390 ;
        RECT 544.020 3432.380 547.020 3432.390 ;
        RECT 724.020 3432.380 727.020 3432.390 ;
        RECT 904.020 3432.380 907.020 3432.390 ;
        RECT 1084.020 3432.380 1087.020 3432.390 ;
        RECT 1264.020 3432.380 1267.020 3432.390 ;
        RECT 1444.020 3432.380 1447.020 3432.390 ;
        RECT 1624.020 3432.380 1627.020 3432.390 ;
        RECT 1804.020 3432.380 1807.020 3432.390 ;
        RECT 1984.020 3432.380 1987.020 3432.390 ;
        RECT 2164.020 3432.380 2167.020 3432.390 ;
        RECT 2344.020 3432.380 2347.020 3432.390 ;
        RECT 2524.020 3432.380 2527.020 3432.390 ;
        RECT 2704.020 3432.380 2707.020 3432.390 ;
        RECT 2884.020 3432.380 2887.020 3432.390 ;
        RECT 2926.600 3432.380 2929.600 3432.390 ;
        RECT -14.680 3429.380 2934.300 3432.380 ;
        RECT -9.980 3429.370 -6.980 3429.380 ;
        RECT 4.020 3429.370 7.020 3429.380 ;
        RECT 184.020 3429.370 187.020 3429.380 ;
        RECT 364.020 3429.370 367.020 3429.380 ;
        RECT 544.020 3429.370 547.020 3429.380 ;
        RECT 724.020 3429.370 727.020 3429.380 ;
        RECT 904.020 3429.370 907.020 3429.380 ;
        RECT 1084.020 3429.370 1087.020 3429.380 ;
        RECT 1264.020 3429.370 1267.020 3429.380 ;
        RECT 1444.020 3429.370 1447.020 3429.380 ;
        RECT 1624.020 3429.370 1627.020 3429.380 ;
        RECT 1804.020 3429.370 1807.020 3429.380 ;
        RECT 1984.020 3429.370 1987.020 3429.380 ;
        RECT 2164.020 3429.370 2167.020 3429.380 ;
        RECT 2344.020 3429.370 2347.020 3429.380 ;
        RECT 2524.020 3429.370 2527.020 3429.380 ;
        RECT 2704.020 3429.370 2707.020 3429.380 ;
        RECT 2884.020 3429.370 2887.020 3429.380 ;
        RECT 2926.600 3429.370 2929.600 3429.380 ;
        RECT -38.180 3306.380 -35.180 3306.390 ;
        RECT 58.020 3306.380 61.020 3306.390 ;
        RECT 238.020 3306.380 241.020 3306.390 ;
        RECT 418.020 3306.380 421.020 3306.390 ;
        RECT 598.020 3306.380 601.020 3306.390 ;
        RECT 778.020 3306.380 781.020 3306.390 ;
        RECT 958.020 3306.380 961.020 3306.390 ;
        RECT 1138.020 3306.380 1141.020 3306.390 ;
        RECT 1318.020 3306.380 1321.020 3306.390 ;
        RECT 1498.020 3306.380 1501.020 3306.390 ;
        RECT 1678.020 3306.380 1681.020 3306.390 ;
        RECT 1858.020 3306.380 1861.020 3306.390 ;
        RECT 2038.020 3306.380 2041.020 3306.390 ;
        RECT 2218.020 3306.380 2221.020 3306.390 ;
        RECT 2398.020 3306.380 2401.020 3306.390 ;
        RECT 2578.020 3306.380 2581.020 3306.390 ;
        RECT 2758.020 3306.380 2761.020 3306.390 ;
        RECT 2954.800 3306.380 2957.800 3306.390 ;
        RECT -42.880 3303.380 2962.500 3306.380 ;
        RECT -38.180 3303.370 -35.180 3303.380 ;
        RECT 58.020 3303.370 61.020 3303.380 ;
        RECT 238.020 3303.370 241.020 3303.380 ;
        RECT 418.020 3303.370 421.020 3303.380 ;
        RECT 598.020 3303.370 601.020 3303.380 ;
        RECT 778.020 3303.370 781.020 3303.380 ;
        RECT 958.020 3303.370 961.020 3303.380 ;
        RECT 1138.020 3303.370 1141.020 3303.380 ;
        RECT 1318.020 3303.370 1321.020 3303.380 ;
        RECT 1498.020 3303.370 1501.020 3303.380 ;
        RECT 1678.020 3303.370 1681.020 3303.380 ;
        RECT 1858.020 3303.370 1861.020 3303.380 ;
        RECT 2038.020 3303.370 2041.020 3303.380 ;
        RECT 2218.020 3303.370 2221.020 3303.380 ;
        RECT 2398.020 3303.370 2401.020 3303.380 ;
        RECT 2578.020 3303.370 2581.020 3303.380 ;
        RECT 2758.020 3303.370 2761.020 3303.380 ;
        RECT 2954.800 3303.370 2957.800 3303.380 ;
        RECT -28.780 3288.380 -25.780 3288.390 ;
        RECT 40.020 3288.380 43.020 3288.390 ;
        RECT 220.020 3288.380 223.020 3288.390 ;
        RECT 400.020 3288.380 403.020 3288.390 ;
        RECT 580.020 3288.380 583.020 3288.390 ;
        RECT 760.020 3288.380 763.020 3288.390 ;
        RECT 940.020 3288.380 943.020 3288.390 ;
        RECT 1120.020 3288.380 1123.020 3288.390 ;
        RECT 1300.020 3288.380 1303.020 3288.390 ;
        RECT 1480.020 3288.380 1483.020 3288.390 ;
        RECT 1660.020 3288.380 1663.020 3288.390 ;
        RECT 1840.020 3288.380 1843.020 3288.390 ;
        RECT 2020.020 3288.380 2023.020 3288.390 ;
        RECT 2200.020 3288.380 2203.020 3288.390 ;
        RECT 2380.020 3288.380 2383.020 3288.390 ;
        RECT 2560.020 3288.380 2563.020 3288.390 ;
        RECT 2740.020 3288.380 2743.020 3288.390 ;
        RECT 2945.400 3288.380 2948.400 3288.390 ;
        RECT -33.480 3285.380 2953.100 3288.380 ;
        RECT -28.780 3285.370 -25.780 3285.380 ;
        RECT 40.020 3285.370 43.020 3285.380 ;
        RECT 220.020 3285.370 223.020 3285.380 ;
        RECT 400.020 3285.370 403.020 3285.380 ;
        RECT 580.020 3285.370 583.020 3285.380 ;
        RECT 760.020 3285.370 763.020 3285.380 ;
        RECT 940.020 3285.370 943.020 3285.380 ;
        RECT 1120.020 3285.370 1123.020 3285.380 ;
        RECT 1300.020 3285.370 1303.020 3285.380 ;
        RECT 1480.020 3285.370 1483.020 3285.380 ;
        RECT 1660.020 3285.370 1663.020 3285.380 ;
        RECT 1840.020 3285.370 1843.020 3285.380 ;
        RECT 2020.020 3285.370 2023.020 3285.380 ;
        RECT 2200.020 3285.370 2203.020 3285.380 ;
        RECT 2380.020 3285.370 2383.020 3285.380 ;
        RECT 2560.020 3285.370 2563.020 3285.380 ;
        RECT 2740.020 3285.370 2743.020 3285.380 ;
        RECT 2945.400 3285.370 2948.400 3285.380 ;
        RECT -19.380 3270.380 -16.380 3270.390 ;
        RECT 22.020 3270.380 25.020 3270.390 ;
        RECT 202.020 3270.380 205.020 3270.390 ;
        RECT 742.020 3270.380 745.020 3270.390 ;
        RECT 922.020 3270.380 925.020 3270.390 ;
        RECT 1462.020 3270.380 1465.020 3270.390 ;
        RECT 2002.020 3270.380 2005.020 3270.390 ;
        RECT 2722.020 3270.380 2725.020 3270.390 ;
        RECT 2902.020 3270.380 2905.020 3270.390 ;
        RECT 2936.000 3270.380 2939.000 3270.390 ;
        RECT -24.080 3267.380 2943.700 3270.380 ;
        RECT -19.380 3267.370 -16.380 3267.380 ;
        RECT 22.020 3267.370 25.020 3267.380 ;
        RECT 202.020 3267.370 205.020 3267.380 ;
        RECT 742.020 3267.370 745.020 3267.380 ;
        RECT 922.020 3267.370 925.020 3267.380 ;
        RECT 1462.020 3267.370 1465.020 3267.380 ;
        RECT 2002.020 3267.370 2005.020 3267.380 ;
        RECT 2722.020 3267.370 2725.020 3267.380 ;
        RECT 2902.020 3267.370 2905.020 3267.380 ;
        RECT 2936.000 3267.370 2939.000 3267.380 ;
        RECT -9.980 3252.380 -6.980 3252.390 ;
        RECT 4.020 3252.380 7.020 3252.390 ;
        RECT 184.020 3252.380 187.020 3252.390 ;
        RECT 724.020 3252.380 727.020 3252.390 ;
        RECT 904.020 3252.380 907.020 3252.390 ;
        RECT 1444.020 3252.380 1447.020 3252.390 ;
        RECT 1984.020 3252.380 1987.020 3252.390 ;
        RECT 2164.020 3252.380 2167.020 3252.390 ;
        RECT 2704.020 3252.380 2707.020 3252.390 ;
        RECT 2884.020 3252.380 2887.020 3252.390 ;
        RECT 2926.600 3252.380 2929.600 3252.390 ;
        RECT -14.680 3249.380 2934.300 3252.380 ;
        RECT -9.980 3249.370 -6.980 3249.380 ;
        RECT 4.020 3249.370 7.020 3249.380 ;
        RECT 184.020 3249.370 187.020 3249.380 ;
        RECT 724.020 3249.370 727.020 3249.380 ;
        RECT 904.020 3249.370 907.020 3249.380 ;
        RECT 1444.020 3249.370 1447.020 3249.380 ;
        RECT 1984.020 3249.370 1987.020 3249.380 ;
        RECT 2164.020 3249.370 2167.020 3249.380 ;
        RECT 2704.020 3249.370 2707.020 3249.380 ;
        RECT 2884.020 3249.370 2887.020 3249.380 ;
        RECT 2926.600 3249.370 2929.600 3249.380 ;
        RECT -38.180 3126.380 -35.180 3126.390 ;
        RECT 58.020 3126.380 61.020 3126.390 ;
        RECT 238.020 3126.380 241.020 3126.390 ;
        RECT 682.470 3126.380 684.070 3126.390 ;
        RECT 778.020 3126.380 781.020 3126.390 ;
        RECT 1332.470 3126.380 1334.070 3126.390 ;
        RECT 1498.020 3126.380 1501.020 3126.390 ;
        RECT 1932.470 3126.380 1934.070 3126.390 ;
        RECT 2038.020 3126.380 2041.020 3126.390 ;
        RECT 2582.470 3126.380 2584.070 3126.390 ;
        RECT 2758.020 3126.380 2761.020 3126.390 ;
        RECT 2954.800 3126.380 2957.800 3126.390 ;
        RECT -42.880 3123.380 2962.500 3126.380 ;
        RECT -38.180 3123.370 -35.180 3123.380 ;
        RECT 58.020 3123.370 61.020 3123.380 ;
        RECT 238.020 3123.370 241.020 3123.380 ;
        RECT 682.470 3123.370 684.070 3123.380 ;
        RECT 778.020 3123.370 781.020 3123.380 ;
        RECT 1332.470 3123.370 1334.070 3123.380 ;
        RECT 1498.020 3123.370 1501.020 3123.380 ;
        RECT 1932.470 3123.370 1934.070 3123.380 ;
        RECT 2038.020 3123.370 2041.020 3123.380 ;
        RECT 2582.470 3123.370 2584.070 3123.380 ;
        RECT 2758.020 3123.370 2761.020 3123.380 ;
        RECT 2954.800 3123.370 2957.800 3123.380 ;
        RECT -28.780 3108.380 -25.780 3108.390 ;
        RECT 40.020 3108.380 43.020 3108.390 ;
        RECT 220.020 3108.380 223.020 3108.390 ;
        RECT 682.470 3108.380 684.070 3108.390 ;
        RECT 760.020 3108.380 763.020 3108.390 ;
        RECT 1332.470 3108.380 1334.070 3108.390 ;
        RECT 1480.020 3108.380 1483.020 3108.390 ;
        RECT 1932.470 3108.380 1934.070 3108.390 ;
        RECT 2020.020 3108.380 2023.020 3108.390 ;
        RECT 2582.470 3108.380 2584.070 3108.390 ;
        RECT 2740.020 3108.380 2743.020 3108.390 ;
        RECT 2945.400 3108.380 2948.400 3108.390 ;
        RECT -33.480 3105.380 2953.100 3108.380 ;
        RECT -28.780 3105.370 -25.780 3105.380 ;
        RECT 40.020 3105.370 43.020 3105.380 ;
        RECT 220.020 3105.370 223.020 3105.380 ;
        RECT 682.470 3105.370 684.070 3105.380 ;
        RECT 760.020 3105.370 763.020 3105.380 ;
        RECT 1332.470 3105.370 1334.070 3105.380 ;
        RECT 1480.020 3105.370 1483.020 3105.380 ;
        RECT 1932.470 3105.370 1934.070 3105.380 ;
        RECT 2020.020 3105.370 2023.020 3105.380 ;
        RECT 2582.470 3105.370 2584.070 3105.380 ;
        RECT 2740.020 3105.370 2743.020 3105.380 ;
        RECT 2945.400 3105.370 2948.400 3105.380 ;
        RECT -19.380 3090.380 -16.380 3090.390 ;
        RECT 22.020 3090.380 25.020 3090.390 ;
        RECT 202.020 3090.380 205.020 3090.390 ;
        RECT 682.470 3090.380 684.070 3090.390 ;
        RECT 742.020 3090.380 745.020 3090.390 ;
        RECT 922.020 3090.380 925.020 3090.390 ;
        RECT 1332.470 3090.380 1334.070 3090.390 ;
        RECT 1462.020 3090.380 1465.020 3090.390 ;
        RECT 1932.470 3090.380 1934.070 3090.390 ;
        RECT 2002.020 3090.380 2005.020 3090.390 ;
        RECT 2582.470 3090.380 2584.070 3090.390 ;
        RECT 2722.020 3090.380 2725.020 3090.390 ;
        RECT 2902.020 3090.380 2905.020 3090.390 ;
        RECT 2936.000 3090.380 2939.000 3090.390 ;
        RECT -24.080 3087.380 2943.700 3090.380 ;
        RECT -19.380 3087.370 -16.380 3087.380 ;
        RECT 22.020 3087.370 25.020 3087.380 ;
        RECT 202.020 3087.370 205.020 3087.380 ;
        RECT 682.470 3087.370 684.070 3087.380 ;
        RECT 742.020 3087.370 745.020 3087.380 ;
        RECT 922.020 3087.370 925.020 3087.380 ;
        RECT 1332.470 3087.370 1334.070 3087.380 ;
        RECT 1462.020 3087.370 1465.020 3087.380 ;
        RECT 1932.470 3087.370 1934.070 3087.380 ;
        RECT 2002.020 3087.370 2005.020 3087.380 ;
        RECT 2582.470 3087.370 2584.070 3087.380 ;
        RECT 2722.020 3087.370 2725.020 3087.380 ;
        RECT 2902.020 3087.370 2905.020 3087.380 ;
        RECT 2936.000 3087.370 2939.000 3087.380 ;
        RECT -9.980 3072.380 -6.980 3072.390 ;
        RECT 4.020 3072.380 7.020 3072.390 ;
        RECT 184.020 3072.380 187.020 3072.390 ;
        RECT 682.470 3072.380 684.070 3072.390 ;
        RECT 724.020 3072.380 727.020 3072.390 ;
        RECT 904.020 3072.380 907.020 3072.390 ;
        RECT 1332.470 3072.380 1334.070 3072.390 ;
        RECT 1444.020 3072.380 1447.020 3072.390 ;
        RECT 1932.470 3072.380 1934.070 3072.390 ;
        RECT 1984.020 3072.380 1987.020 3072.390 ;
        RECT 2164.020 3072.380 2167.020 3072.390 ;
        RECT 2582.470 3072.380 2584.070 3072.390 ;
        RECT 2704.020 3072.380 2707.020 3072.390 ;
        RECT 2884.020 3072.380 2887.020 3072.390 ;
        RECT 2926.600 3072.380 2929.600 3072.390 ;
        RECT -14.680 3069.380 2934.300 3072.380 ;
        RECT -9.980 3069.370 -6.980 3069.380 ;
        RECT 4.020 3069.370 7.020 3069.380 ;
        RECT 184.020 3069.370 187.020 3069.380 ;
        RECT 682.470 3069.370 684.070 3069.380 ;
        RECT 724.020 3069.370 727.020 3069.380 ;
        RECT 904.020 3069.370 907.020 3069.380 ;
        RECT 1332.470 3069.370 1334.070 3069.380 ;
        RECT 1444.020 3069.370 1447.020 3069.380 ;
        RECT 1932.470 3069.370 1934.070 3069.380 ;
        RECT 1984.020 3069.370 1987.020 3069.380 ;
        RECT 2164.020 3069.370 2167.020 3069.380 ;
        RECT 2582.470 3069.370 2584.070 3069.380 ;
        RECT 2704.020 3069.370 2707.020 3069.380 ;
        RECT 2884.020 3069.370 2887.020 3069.380 ;
        RECT 2926.600 3069.370 2929.600 3069.380 ;
        RECT -38.180 2946.380 -35.180 2946.390 ;
        RECT 58.020 2946.380 61.020 2946.390 ;
        RECT 238.020 2946.380 241.020 2946.390 ;
        RECT 682.470 2946.380 684.070 2946.390 ;
        RECT 778.020 2946.380 781.020 2946.390 ;
        RECT 1332.470 2946.380 1334.070 2946.390 ;
        RECT 1498.020 2946.380 1501.020 2946.390 ;
        RECT 1932.470 2946.380 1934.070 2946.390 ;
        RECT 2038.020 2946.380 2041.020 2946.390 ;
        RECT 2582.470 2946.380 2584.070 2946.390 ;
        RECT 2758.020 2946.380 2761.020 2946.390 ;
        RECT 2954.800 2946.380 2957.800 2946.390 ;
        RECT -42.880 2943.380 2962.500 2946.380 ;
        RECT -38.180 2943.370 -35.180 2943.380 ;
        RECT 58.020 2943.370 61.020 2943.380 ;
        RECT 238.020 2943.370 241.020 2943.380 ;
        RECT 682.470 2943.370 684.070 2943.380 ;
        RECT 778.020 2943.370 781.020 2943.380 ;
        RECT 1332.470 2943.370 1334.070 2943.380 ;
        RECT 1498.020 2943.370 1501.020 2943.380 ;
        RECT 1932.470 2943.370 1934.070 2943.380 ;
        RECT 2038.020 2943.370 2041.020 2943.380 ;
        RECT 2582.470 2943.370 2584.070 2943.380 ;
        RECT 2758.020 2943.370 2761.020 2943.380 ;
        RECT 2954.800 2943.370 2957.800 2943.380 ;
        RECT -28.780 2928.380 -25.780 2928.390 ;
        RECT 40.020 2928.380 43.020 2928.390 ;
        RECT 220.020 2928.380 223.020 2928.390 ;
        RECT 682.470 2928.380 684.070 2928.390 ;
        RECT 760.020 2928.380 763.020 2928.390 ;
        RECT 1332.470 2928.380 1334.070 2928.390 ;
        RECT 1480.020 2928.380 1483.020 2928.390 ;
        RECT 1932.470 2928.380 1934.070 2928.390 ;
        RECT 2020.020 2928.380 2023.020 2928.390 ;
        RECT 2582.470 2928.380 2584.070 2928.390 ;
        RECT 2740.020 2928.380 2743.020 2928.390 ;
        RECT 2945.400 2928.380 2948.400 2928.390 ;
        RECT -33.480 2925.380 2953.100 2928.380 ;
        RECT -28.780 2925.370 -25.780 2925.380 ;
        RECT 40.020 2925.370 43.020 2925.380 ;
        RECT 220.020 2925.370 223.020 2925.380 ;
        RECT 682.470 2925.370 684.070 2925.380 ;
        RECT 760.020 2925.370 763.020 2925.380 ;
        RECT 1332.470 2925.370 1334.070 2925.380 ;
        RECT 1480.020 2925.370 1483.020 2925.380 ;
        RECT 1932.470 2925.370 1934.070 2925.380 ;
        RECT 2020.020 2925.370 2023.020 2925.380 ;
        RECT 2582.470 2925.370 2584.070 2925.380 ;
        RECT 2740.020 2925.370 2743.020 2925.380 ;
        RECT 2945.400 2925.370 2948.400 2925.380 ;
        RECT -19.380 2910.380 -16.380 2910.390 ;
        RECT 22.020 2910.380 25.020 2910.390 ;
        RECT 202.020 2910.380 205.020 2910.390 ;
        RECT 682.470 2910.380 684.070 2910.390 ;
        RECT 742.020 2910.380 745.020 2910.390 ;
        RECT 922.020 2910.380 925.020 2910.390 ;
        RECT 1332.470 2910.380 1334.070 2910.390 ;
        RECT 1462.020 2910.380 1465.020 2910.390 ;
        RECT 1932.470 2910.380 1934.070 2910.390 ;
        RECT 2002.020 2910.380 2005.020 2910.390 ;
        RECT 2582.470 2910.380 2584.070 2910.390 ;
        RECT 2722.020 2910.380 2725.020 2910.390 ;
        RECT 2902.020 2910.380 2905.020 2910.390 ;
        RECT 2936.000 2910.380 2939.000 2910.390 ;
        RECT -24.080 2907.380 2943.700 2910.380 ;
        RECT -19.380 2907.370 -16.380 2907.380 ;
        RECT 22.020 2907.370 25.020 2907.380 ;
        RECT 202.020 2907.370 205.020 2907.380 ;
        RECT 682.470 2907.370 684.070 2907.380 ;
        RECT 742.020 2907.370 745.020 2907.380 ;
        RECT 922.020 2907.370 925.020 2907.380 ;
        RECT 1332.470 2907.370 1334.070 2907.380 ;
        RECT 1462.020 2907.370 1465.020 2907.380 ;
        RECT 1932.470 2907.370 1934.070 2907.380 ;
        RECT 2002.020 2907.370 2005.020 2907.380 ;
        RECT 2582.470 2907.370 2584.070 2907.380 ;
        RECT 2722.020 2907.370 2725.020 2907.380 ;
        RECT 2902.020 2907.370 2905.020 2907.380 ;
        RECT 2936.000 2907.370 2939.000 2907.380 ;
        RECT -9.980 2892.380 -6.980 2892.390 ;
        RECT 4.020 2892.380 7.020 2892.390 ;
        RECT 184.020 2892.380 187.020 2892.390 ;
        RECT 682.470 2892.380 684.070 2892.390 ;
        RECT 724.020 2892.380 727.020 2892.390 ;
        RECT 904.020 2892.380 907.020 2892.390 ;
        RECT 1332.470 2892.380 1334.070 2892.390 ;
        RECT 1444.020 2892.380 1447.020 2892.390 ;
        RECT 1932.470 2892.380 1934.070 2892.390 ;
        RECT 1984.020 2892.380 1987.020 2892.390 ;
        RECT 2164.020 2892.380 2167.020 2892.390 ;
        RECT 2582.470 2892.380 2584.070 2892.390 ;
        RECT 2704.020 2892.380 2707.020 2892.390 ;
        RECT 2884.020 2892.380 2887.020 2892.390 ;
        RECT 2926.600 2892.380 2929.600 2892.390 ;
        RECT -14.680 2889.380 2934.300 2892.380 ;
        RECT -9.980 2889.370 -6.980 2889.380 ;
        RECT 4.020 2889.370 7.020 2889.380 ;
        RECT 184.020 2889.370 187.020 2889.380 ;
        RECT 682.470 2889.370 684.070 2889.380 ;
        RECT 724.020 2889.370 727.020 2889.380 ;
        RECT 904.020 2889.370 907.020 2889.380 ;
        RECT 1332.470 2889.370 1334.070 2889.380 ;
        RECT 1444.020 2889.370 1447.020 2889.380 ;
        RECT 1932.470 2889.370 1934.070 2889.380 ;
        RECT 1984.020 2889.370 1987.020 2889.380 ;
        RECT 2164.020 2889.370 2167.020 2889.380 ;
        RECT 2582.470 2889.370 2584.070 2889.380 ;
        RECT 2704.020 2889.370 2707.020 2889.380 ;
        RECT 2884.020 2889.370 2887.020 2889.380 ;
        RECT 2926.600 2889.370 2929.600 2889.380 ;
        RECT -38.180 2766.380 -35.180 2766.390 ;
        RECT 58.020 2766.380 61.020 2766.390 ;
        RECT 238.020 2766.380 241.020 2766.390 ;
        RECT 418.020 2766.380 421.020 2766.390 ;
        RECT 598.020 2766.380 601.020 2766.390 ;
        RECT 778.020 2766.380 781.020 2766.390 ;
        RECT 958.020 2766.380 961.020 2766.390 ;
        RECT 1138.020 2766.380 1141.020 2766.390 ;
        RECT 1318.020 2766.380 1321.020 2766.390 ;
        RECT 1498.020 2766.380 1501.020 2766.390 ;
        RECT 1678.020 2766.380 1681.020 2766.390 ;
        RECT 1858.020 2766.380 1861.020 2766.390 ;
        RECT 2038.020 2766.380 2041.020 2766.390 ;
        RECT 2218.020 2766.380 2221.020 2766.390 ;
        RECT 2398.020 2766.380 2401.020 2766.390 ;
        RECT 2578.020 2766.380 2581.020 2766.390 ;
        RECT 2758.020 2766.380 2761.020 2766.390 ;
        RECT 2954.800 2766.380 2957.800 2766.390 ;
        RECT -42.880 2763.380 2962.500 2766.380 ;
        RECT -38.180 2763.370 -35.180 2763.380 ;
        RECT 58.020 2763.370 61.020 2763.380 ;
        RECT 238.020 2763.370 241.020 2763.380 ;
        RECT 418.020 2763.370 421.020 2763.380 ;
        RECT 598.020 2763.370 601.020 2763.380 ;
        RECT 778.020 2763.370 781.020 2763.380 ;
        RECT 958.020 2763.370 961.020 2763.380 ;
        RECT 1138.020 2763.370 1141.020 2763.380 ;
        RECT 1318.020 2763.370 1321.020 2763.380 ;
        RECT 1498.020 2763.370 1501.020 2763.380 ;
        RECT 1678.020 2763.370 1681.020 2763.380 ;
        RECT 1858.020 2763.370 1861.020 2763.380 ;
        RECT 2038.020 2763.370 2041.020 2763.380 ;
        RECT 2218.020 2763.370 2221.020 2763.380 ;
        RECT 2398.020 2763.370 2401.020 2763.380 ;
        RECT 2578.020 2763.370 2581.020 2763.380 ;
        RECT 2758.020 2763.370 2761.020 2763.380 ;
        RECT 2954.800 2763.370 2957.800 2763.380 ;
        RECT -28.780 2748.380 -25.780 2748.390 ;
        RECT 40.020 2748.380 43.020 2748.390 ;
        RECT 220.020 2748.380 223.020 2748.390 ;
        RECT 400.020 2748.380 403.020 2748.390 ;
        RECT 580.020 2748.380 583.020 2748.390 ;
        RECT 760.020 2748.380 763.020 2748.390 ;
        RECT 940.020 2748.380 943.020 2748.390 ;
        RECT 1120.020 2748.380 1123.020 2748.390 ;
        RECT 1300.020 2748.380 1303.020 2748.390 ;
        RECT 1480.020 2748.380 1483.020 2748.390 ;
        RECT 1660.020 2748.380 1663.020 2748.390 ;
        RECT 1840.020 2748.380 1843.020 2748.390 ;
        RECT 2020.020 2748.380 2023.020 2748.390 ;
        RECT 2200.020 2748.380 2203.020 2748.390 ;
        RECT 2380.020 2748.380 2383.020 2748.390 ;
        RECT 2560.020 2748.380 2563.020 2748.390 ;
        RECT 2740.020 2748.380 2743.020 2748.390 ;
        RECT 2945.400 2748.380 2948.400 2748.390 ;
        RECT -33.480 2745.380 2953.100 2748.380 ;
        RECT -28.780 2745.370 -25.780 2745.380 ;
        RECT 40.020 2745.370 43.020 2745.380 ;
        RECT 220.020 2745.370 223.020 2745.380 ;
        RECT 400.020 2745.370 403.020 2745.380 ;
        RECT 580.020 2745.370 583.020 2745.380 ;
        RECT 760.020 2745.370 763.020 2745.380 ;
        RECT 940.020 2745.370 943.020 2745.380 ;
        RECT 1120.020 2745.370 1123.020 2745.380 ;
        RECT 1300.020 2745.370 1303.020 2745.380 ;
        RECT 1480.020 2745.370 1483.020 2745.380 ;
        RECT 1660.020 2745.370 1663.020 2745.380 ;
        RECT 1840.020 2745.370 1843.020 2745.380 ;
        RECT 2020.020 2745.370 2023.020 2745.380 ;
        RECT 2200.020 2745.370 2203.020 2745.380 ;
        RECT 2380.020 2745.370 2383.020 2745.380 ;
        RECT 2560.020 2745.370 2563.020 2745.380 ;
        RECT 2740.020 2745.370 2743.020 2745.380 ;
        RECT 2945.400 2745.370 2948.400 2745.380 ;
        RECT -19.380 2730.380 -16.380 2730.390 ;
        RECT 22.020 2730.380 25.020 2730.390 ;
        RECT 202.020 2730.380 205.020 2730.390 ;
        RECT 382.020 2730.380 385.020 2730.390 ;
        RECT 562.020 2730.380 565.020 2730.390 ;
        RECT 742.020 2730.380 745.020 2730.390 ;
        RECT 922.020 2730.380 925.020 2730.390 ;
        RECT 1102.020 2730.380 1105.020 2730.390 ;
        RECT 1282.020 2730.380 1285.020 2730.390 ;
        RECT 1462.020 2730.380 1465.020 2730.390 ;
        RECT 1642.020 2730.380 1645.020 2730.390 ;
        RECT 1822.020 2730.380 1825.020 2730.390 ;
        RECT 2002.020 2730.380 2005.020 2730.390 ;
        RECT 2182.020 2730.380 2185.020 2730.390 ;
        RECT 2362.020 2730.380 2365.020 2730.390 ;
        RECT 2542.020 2730.380 2545.020 2730.390 ;
        RECT 2722.020 2730.380 2725.020 2730.390 ;
        RECT 2902.020 2730.380 2905.020 2730.390 ;
        RECT 2936.000 2730.380 2939.000 2730.390 ;
        RECT -24.080 2727.380 2943.700 2730.380 ;
        RECT -19.380 2727.370 -16.380 2727.380 ;
        RECT 22.020 2727.370 25.020 2727.380 ;
        RECT 202.020 2727.370 205.020 2727.380 ;
        RECT 382.020 2727.370 385.020 2727.380 ;
        RECT 562.020 2727.370 565.020 2727.380 ;
        RECT 742.020 2727.370 745.020 2727.380 ;
        RECT 922.020 2727.370 925.020 2727.380 ;
        RECT 1102.020 2727.370 1105.020 2727.380 ;
        RECT 1282.020 2727.370 1285.020 2727.380 ;
        RECT 1462.020 2727.370 1465.020 2727.380 ;
        RECT 1642.020 2727.370 1645.020 2727.380 ;
        RECT 1822.020 2727.370 1825.020 2727.380 ;
        RECT 2002.020 2727.370 2005.020 2727.380 ;
        RECT 2182.020 2727.370 2185.020 2727.380 ;
        RECT 2362.020 2727.370 2365.020 2727.380 ;
        RECT 2542.020 2727.370 2545.020 2727.380 ;
        RECT 2722.020 2727.370 2725.020 2727.380 ;
        RECT 2902.020 2727.370 2905.020 2727.380 ;
        RECT 2936.000 2727.370 2939.000 2727.380 ;
        RECT -9.980 2712.380 -6.980 2712.390 ;
        RECT 4.020 2712.380 7.020 2712.390 ;
        RECT 184.020 2712.380 187.020 2712.390 ;
        RECT 1444.020 2712.380 1447.020 2712.390 ;
        RECT 1624.020 2712.380 1627.020 2712.390 ;
        RECT 1804.020 2712.380 1807.020 2712.390 ;
        RECT 1984.020 2712.380 1987.020 2712.390 ;
        RECT 2164.020 2712.380 2167.020 2712.390 ;
        RECT 2344.020 2712.380 2347.020 2712.390 ;
        RECT 2524.020 2712.380 2527.020 2712.390 ;
        RECT 2704.020 2712.380 2707.020 2712.390 ;
        RECT 2884.020 2712.380 2887.020 2712.390 ;
        RECT 2926.600 2712.380 2929.600 2712.390 ;
        RECT -14.680 2709.380 2934.300 2712.380 ;
        RECT -9.980 2709.370 -6.980 2709.380 ;
        RECT 4.020 2709.370 7.020 2709.380 ;
        RECT 184.020 2709.370 187.020 2709.380 ;
        RECT 1444.020 2709.370 1447.020 2709.380 ;
        RECT 1624.020 2709.370 1627.020 2709.380 ;
        RECT 1804.020 2709.370 1807.020 2709.380 ;
        RECT 1984.020 2709.370 1987.020 2709.380 ;
        RECT 2164.020 2709.370 2167.020 2709.380 ;
        RECT 2344.020 2709.370 2347.020 2709.380 ;
        RECT 2524.020 2709.370 2527.020 2709.380 ;
        RECT 2704.020 2709.370 2707.020 2709.380 ;
        RECT 2884.020 2709.370 2887.020 2709.380 ;
        RECT 2926.600 2709.370 2929.600 2709.380 ;
        RECT -38.180 2586.380 -35.180 2586.390 ;
        RECT 58.020 2586.380 61.020 2586.390 ;
        RECT 238.020 2586.380 241.020 2586.390 ;
        RECT 321.040 2586.380 322.640 2586.390 ;
        RECT 1498.020 2586.380 1501.020 2586.390 ;
        RECT 1678.020 2586.380 1681.020 2586.390 ;
        RECT 1858.020 2586.380 1861.020 2586.390 ;
        RECT 2038.020 2586.380 2041.020 2586.390 ;
        RECT 2218.020 2586.380 2221.020 2586.390 ;
        RECT 2398.020 2586.380 2401.020 2586.390 ;
        RECT 2578.020 2586.380 2581.020 2586.390 ;
        RECT 2758.020 2586.380 2761.020 2586.390 ;
        RECT 2954.800 2586.380 2957.800 2586.390 ;
        RECT -42.880 2583.380 2962.500 2586.380 ;
        RECT -38.180 2583.370 -35.180 2583.380 ;
        RECT 58.020 2583.370 61.020 2583.380 ;
        RECT 238.020 2583.370 241.020 2583.380 ;
        RECT 321.040 2583.370 322.640 2583.380 ;
        RECT 1498.020 2583.370 1501.020 2583.380 ;
        RECT 1678.020 2583.370 1681.020 2583.380 ;
        RECT 1858.020 2583.370 1861.020 2583.380 ;
        RECT 2038.020 2583.370 2041.020 2583.380 ;
        RECT 2218.020 2583.370 2221.020 2583.380 ;
        RECT 2398.020 2583.370 2401.020 2583.380 ;
        RECT 2578.020 2583.370 2581.020 2583.380 ;
        RECT 2758.020 2583.370 2761.020 2583.380 ;
        RECT 2954.800 2583.370 2957.800 2583.380 ;
        RECT -28.780 2568.380 -25.780 2568.390 ;
        RECT 40.020 2568.380 43.020 2568.390 ;
        RECT 220.020 2568.380 223.020 2568.390 ;
        RECT 321.040 2568.380 322.640 2568.390 ;
        RECT 1480.020 2568.380 1483.020 2568.390 ;
        RECT 1660.020 2568.380 1663.020 2568.390 ;
        RECT 1840.020 2568.380 1843.020 2568.390 ;
        RECT 2020.020 2568.380 2023.020 2568.390 ;
        RECT 2200.020 2568.380 2203.020 2568.390 ;
        RECT 2380.020 2568.380 2383.020 2568.390 ;
        RECT 2560.020 2568.380 2563.020 2568.390 ;
        RECT 2740.020 2568.380 2743.020 2568.390 ;
        RECT 2945.400 2568.380 2948.400 2568.390 ;
        RECT -33.480 2565.380 2953.100 2568.380 ;
        RECT -28.780 2565.370 -25.780 2565.380 ;
        RECT 40.020 2565.370 43.020 2565.380 ;
        RECT 220.020 2565.370 223.020 2565.380 ;
        RECT 321.040 2565.370 322.640 2565.380 ;
        RECT 1480.020 2565.370 1483.020 2565.380 ;
        RECT 1660.020 2565.370 1663.020 2565.380 ;
        RECT 1840.020 2565.370 1843.020 2565.380 ;
        RECT 2020.020 2565.370 2023.020 2565.380 ;
        RECT 2200.020 2565.370 2203.020 2565.380 ;
        RECT 2380.020 2565.370 2383.020 2565.380 ;
        RECT 2560.020 2565.370 2563.020 2565.380 ;
        RECT 2740.020 2565.370 2743.020 2565.380 ;
        RECT 2945.400 2565.370 2948.400 2565.380 ;
        RECT -19.380 2550.380 -16.380 2550.390 ;
        RECT 22.020 2550.380 25.020 2550.390 ;
        RECT 202.020 2550.380 205.020 2550.390 ;
        RECT 321.040 2550.380 322.640 2550.390 ;
        RECT 1462.020 2550.380 1465.020 2550.390 ;
        RECT 1642.020 2550.380 1645.020 2550.390 ;
        RECT 1822.020 2550.380 1825.020 2550.390 ;
        RECT 2002.020 2550.380 2005.020 2550.390 ;
        RECT 2182.020 2550.380 2185.020 2550.390 ;
        RECT 2362.020 2550.380 2365.020 2550.390 ;
        RECT 2542.020 2550.380 2545.020 2550.390 ;
        RECT 2722.020 2550.380 2725.020 2550.390 ;
        RECT 2902.020 2550.380 2905.020 2550.390 ;
        RECT 2936.000 2550.380 2939.000 2550.390 ;
        RECT -24.080 2547.380 2943.700 2550.380 ;
        RECT -19.380 2547.370 -16.380 2547.380 ;
        RECT 22.020 2547.370 25.020 2547.380 ;
        RECT 202.020 2547.370 205.020 2547.380 ;
        RECT 321.040 2547.370 322.640 2547.380 ;
        RECT 1462.020 2547.370 1465.020 2547.380 ;
        RECT 1642.020 2547.370 1645.020 2547.380 ;
        RECT 1822.020 2547.370 1825.020 2547.380 ;
        RECT 2002.020 2547.370 2005.020 2547.380 ;
        RECT 2182.020 2547.370 2185.020 2547.380 ;
        RECT 2362.020 2547.370 2365.020 2547.380 ;
        RECT 2542.020 2547.370 2545.020 2547.380 ;
        RECT 2722.020 2547.370 2725.020 2547.380 ;
        RECT 2902.020 2547.370 2905.020 2547.380 ;
        RECT 2936.000 2547.370 2939.000 2547.380 ;
        RECT -9.980 2532.380 -6.980 2532.390 ;
        RECT 4.020 2532.380 7.020 2532.390 ;
        RECT 184.020 2532.380 187.020 2532.390 ;
        RECT 321.040 2532.380 322.640 2532.390 ;
        RECT 1444.020 2532.380 1447.020 2532.390 ;
        RECT 1624.020 2532.380 1627.020 2532.390 ;
        RECT 1804.020 2532.380 1807.020 2532.390 ;
        RECT 1984.020 2532.380 1987.020 2532.390 ;
        RECT 2164.020 2532.380 2167.020 2532.390 ;
        RECT 2344.020 2532.380 2347.020 2532.390 ;
        RECT 2524.020 2532.380 2527.020 2532.390 ;
        RECT 2704.020 2532.380 2707.020 2532.390 ;
        RECT 2884.020 2532.380 2887.020 2532.390 ;
        RECT 2926.600 2532.380 2929.600 2532.390 ;
        RECT -14.680 2529.380 2934.300 2532.380 ;
        RECT -9.980 2529.370 -6.980 2529.380 ;
        RECT 4.020 2529.370 7.020 2529.380 ;
        RECT 184.020 2529.370 187.020 2529.380 ;
        RECT 321.040 2529.370 322.640 2529.380 ;
        RECT 1444.020 2529.370 1447.020 2529.380 ;
        RECT 1624.020 2529.370 1627.020 2529.380 ;
        RECT 1804.020 2529.370 1807.020 2529.380 ;
        RECT 1984.020 2529.370 1987.020 2529.380 ;
        RECT 2164.020 2529.370 2167.020 2529.380 ;
        RECT 2344.020 2529.370 2347.020 2529.380 ;
        RECT 2524.020 2529.370 2527.020 2529.380 ;
        RECT 2704.020 2529.370 2707.020 2529.380 ;
        RECT 2884.020 2529.370 2887.020 2529.380 ;
        RECT 2926.600 2529.370 2929.600 2529.380 ;
        RECT -38.180 2406.380 -35.180 2406.390 ;
        RECT 58.020 2406.380 61.020 2406.390 ;
        RECT 238.020 2406.380 241.020 2406.390 ;
        RECT 321.040 2406.380 322.640 2406.390 ;
        RECT 1498.020 2406.380 1501.020 2406.390 ;
        RECT 1678.020 2406.380 1681.020 2406.390 ;
        RECT 1858.020 2406.380 1861.020 2406.390 ;
        RECT 2038.020 2406.380 2041.020 2406.390 ;
        RECT 2218.020 2406.380 2221.020 2406.390 ;
        RECT 2398.020 2406.380 2401.020 2406.390 ;
        RECT 2578.020 2406.380 2581.020 2406.390 ;
        RECT 2758.020 2406.380 2761.020 2406.390 ;
        RECT 2954.800 2406.380 2957.800 2406.390 ;
        RECT -42.880 2403.380 2962.500 2406.380 ;
        RECT -38.180 2403.370 -35.180 2403.380 ;
        RECT 58.020 2403.370 61.020 2403.380 ;
        RECT 238.020 2403.370 241.020 2403.380 ;
        RECT 321.040 2403.370 322.640 2403.380 ;
        RECT 1498.020 2403.370 1501.020 2403.380 ;
        RECT 1678.020 2403.370 1681.020 2403.380 ;
        RECT 1858.020 2403.370 1861.020 2403.380 ;
        RECT 2038.020 2403.370 2041.020 2403.380 ;
        RECT 2218.020 2403.370 2221.020 2403.380 ;
        RECT 2398.020 2403.370 2401.020 2403.380 ;
        RECT 2578.020 2403.370 2581.020 2403.380 ;
        RECT 2758.020 2403.370 2761.020 2403.380 ;
        RECT 2954.800 2403.370 2957.800 2403.380 ;
        RECT -28.780 2388.380 -25.780 2388.390 ;
        RECT 40.020 2388.380 43.020 2388.390 ;
        RECT 220.020 2388.380 223.020 2388.390 ;
        RECT 321.040 2388.380 322.640 2388.390 ;
        RECT 1480.020 2388.380 1483.020 2388.390 ;
        RECT 1660.020 2388.380 1663.020 2388.390 ;
        RECT 1840.020 2388.380 1843.020 2388.390 ;
        RECT 2020.020 2388.380 2023.020 2388.390 ;
        RECT 2200.020 2388.380 2203.020 2388.390 ;
        RECT 2380.020 2388.380 2383.020 2388.390 ;
        RECT 2560.020 2388.380 2563.020 2388.390 ;
        RECT 2740.020 2388.380 2743.020 2388.390 ;
        RECT 2945.400 2388.380 2948.400 2388.390 ;
        RECT -33.480 2385.380 2953.100 2388.380 ;
        RECT -28.780 2385.370 -25.780 2385.380 ;
        RECT 40.020 2385.370 43.020 2385.380 ;
        RECT 220.020 2385.370 223.020 2385.380 ;
        RECT 321.040 2385.370 322.640 2385.380 ;
        RECT 1480.020 2385.370 1483.020 2385.380 ;
        RECT 1660.020 2385.370 1663.020 2385.380 ;
        RECT 1840.020 2385.370 1843.020 2385.380 ;
        RECT 2020.020 2385.370 2023.020 2385.380 ;
        RECT 2200.020 2385.370 2203.020 2385.380 ;
        RECT 2380.020 2385.370 2383.020 2385.380 ;
        RECT 2560.020 2385.370 2563.020 2385.380 ;
        RECT 2740.020 2385.370 2743.020 2385.380 ;
        RECT 2945.400 2385.370 2948.400 2385.380 ;
        RECT -19.380 2370.380 -16.380 2370.390 ;
        RECT 22.020 2370.380 25.020 2370.390 ;
        RECT 202.020 2370.380 205.020 2370.390 ;
        RECT 321.040 2370.380 322.640 2370.390 ;
        RECT 1462.020 2370.380 1465.020 2370.390 ;
        RECT 1642.020 2370.380 1645.020 2370.390 ;
        RECT 1822.020 2370.380 1825.020 2370.390 ;
        RECT 2002.020 2370.380 2005.020 2370.390 ;
        RECT 2182.020 2370.380 2185.020 2370.390 ;
        RECT 2362.020 2370.380 2365.020 2370.390 ;
        RECT 2542.020 2370.380 2545.020 2370.390 ;
        RECT 2722.020 2370.380 2725.020 2370.390 ;
        RECT 2902.020 2370.380 2905.020 2370.390 ;
        RECT 2936.000 2370.380 2939.000 2370.390 ;
        RECT -24.080 2367.380 2943.700 2370.380 ;
        RECT -19.380 2367.370 -16.380 2367.380 ;
        RECT 22.020 2367.370 25.020 2367.380 ;
        RECT 202.020 2367.370 205.020 2367.380 ;
        RECT 321.040 2367.370 322.640 2367.380 ;
        RECT 1462.020 2367.370 1465.020 2367.380 ;
        RECT 1642.020 2367.370 1645.020 2367.380 ;
        RECT 1822.020 2367.370 1825.020 2367.380 ;
        RECT 2002.020 2367.370 2005.020 2367.380 ;
        RECT 2182.020 2367.370 2185.020 2367.380 ;
        RECT 2362.020 2367.370 2365.020 2367.380 ;
        RECT 2542.020 2367.370 2545.020 2367.380 ;
        RECT 2722.020 2367.370 2725.020 2367.380 ;
        RECT 2902.020 2367.370 2905.020 2367.380 ;
        RECT 2936.000 2367.370 2939.000 2367.380 ;
        RECT -9.980 2352.380 -6.980 2352.390 ;
        RECT 4.020 2352.380 7.020 2352.390 ;
        RECT 184.020 2352.380 187.020 2352.390 ;
        RECT 321.040 2352.380 322.640 2352.390 ;
        RECT 1444.020 2352.380 1447.020 2352.390 ;
        RECT 1624.020 2352.380 1627.020 2352.390 ;
        RECT 1804.020 2352.380 1807.020 2352.390 ;
        RECT 1984.020 2352.380 1987.020 2352.390 ;
        RECT 2164.020 2352.380 2167.020 2352.390 ;
        RECT 2344.020 2352.380 2347.020 2352.390 ;
        RECT 2524.020 2352.380 2527.020 2352.390 ;
        RECT 2704.020 2352.380 2707.020 2352.390 ;
        RECT 2884.020 2352.380 2887.020 2352.390 ;
        RECT 2926.600 2352.380 2929.600 2352.390 ;
        RECT -14.680 2349.380 2934.300 2352.380 ;
        RECT -9.980 2349.370 -6.980 2349.380 ;
        RECT 4.020 2349.370 7.020 2349.380 ;
        RECT 184.020 2349.370 187.020 2349.380 ;
        RECT 321.040 2349.370 322.640 2349.380 ;
        RECT 1444.020 2349.370 1447.020 2349.380 ;
        RECT 1624.020 2349.370 1627.020 2349.380 ;
        RECT 1804.020 2349.370 1807.020 2349.380 ;
        RECT 1984.020 2349.370 1987.020 2349.380 ;
        RECT 2164.020 2349.370 2167.020 2349.380 ;
        RECT 2344.020 2349.370 2347.020 2349.380 ;
        RECT 2524.020 2349.370 2527.020 2349.380 ;
        RECT 2704.020 2349.370 2707.020 2349.380 ;
        RECT 2884.020 2349.370 2887.020 2349.380 ;
        RECT 2926.600 2349.370 2929.600 2349.380 ;
        RECT -38.180 2226.380 -35.180 2226.390 ;
        RECT 58.020 2226.380 61.020 2226.390 ;
        RECT 238.020 2226.380 241.020 2226.390 ;
        RECT 321.040 2226.380 322.640 2226.390 ;
        RECT 1498.020 2226.380 1501.020 2226.390 ;
        RECT 1678.020 2226.380 1681.020 2226.390 ;
        RECT 1858.020 2226.380 1861.020 2226.390 ;
        RECT 2038.020 2226.380 2041.020 2226.390 ;
        RECT 2218.020 2226.380 2221.020 2226.390 ;
        RECT 2398.020 2226.380 2401.020 2226.390 ;
        RECT 2578.020 2226.380 2581.020 2226.390 ;
        RECT 2758.020 2226.380 2761.020 2226.390 ;
        RECT 2954.800 2226.380 2957.800 2226.390 ;
        RECT -42.880 2223.380 2962.500 2226.380 ;
        RECT -38.180 2223.370 -35.180 2223.380 ;
        RECT 58.020 2223.370 61.020 2223.380 ;
        RECT 238.020 2223.370 241.020 2223.380 ;
        RECT 321.040 2223.370 322.640 2223.380 ;
        RECT 1498.020 2223.370 1501.020 2223.380 ;
        RECT 1678.020 2223.370 1681.020 2223.380 ;
        RECT 1858.020 2223.370 1861.020 2223.380 ;
        RECT 2038.020 2223.370 2041.020 2223.380 ;
        RECT 2218.020 2223.370 2221.020 2223.380 ;
        RECT 2398.020 2223.370 2401.020 2223.380 ;
        RECT 2578.020 2223.370 2581.020 2223.380 ;
        RECT 2758.020 2223.370 2761.020 2223.380 ;
        RECT 2954.800 2223.370 2957.800 2223.380 ;
        RECT -28.780 2208.380 -25.780 2208.390 ;
        RECT 40.020 2208.380 43.020 2208.390 ;
        RECT 220.020 2208.380 223.020 2208.390 ;
        RECT 321.040 2208.380 322.640 2208.390 ;
        RECT 1480.020 2208.380 1483.020 2208.390 ;
        RECT 1660.020 2208.380 1663.020 2208.390 ;
        RECT 1840.020 2208.380 1843.020 2208.390 ;
        RECT 2020.020 2208.380 2023.020 2208.390 ;
        RECT 2200.020 2208.380 2203.020 2208.390 ;
        RECT 2380.020 2208.380 2383.020 2208.390 ;
        RECT 2560.020 2208.380 2563.020 2208.390 ;
        RECT 2740.020 2208.380 2743.020 2208.390 ;
        RECT 2945.400 2208.380 2948.400 2208.390 ;
        RECT -33.480 2205.380 2953.100 2208.380 ;
        RECT -28.780 2205.370 -25.780 2205.380 ;
        RECT 40.020 2205.370 43.020 2205.380 ;
        RECT 220.020 2205.370 223.020 2205.380 ;
        RECT 321.040 2205.370 322.640 2205.380 ;
        RECT 1480.020 2205.370 1483.020 2205.380 ;
        RECT 1660.020 2205.370 1663.020 2205.380 ;
        RECT 1840.020 2205.370 1843.020 2205.380 ;
        RECT 2020.020 2205.370 2023.020 2205.380 ;
        RECT 2200.020 2205.370 2203.020 2205.380 ;
        RECT 2380.020 2205.370 2383.020 2205.380 ;
        RECT 2560.020 2205.370 2563.020 2205.380 ;
        RECT 2740.020 2205.370 2743.020 2205.380 ;
        RECT 2945.400 2205.370 2948.400 2205.380 ;
        RECT -19.380 2190.380 -16.380 2190.390 ;
        RECT 22.020 2190.380 25.020 2190.390 ;
        RECT 202.020 2190.380 205.020 2190.390 ;
        RECT 321.040 2190.380 322.640 2190.390 ;
        RECT 1462.020 2190.380 1465.020 2190.390 ;
        RECT 1642.020 2190.380 1645.020 2190.390 ;
        RECT 1822.020 2190.380 1825.020 2190.390 ;
        RECT 2002.020 2190.380 2005.020 2190.390 ;
        RECT 2182.020 2190.380 2185.020 2190.390 ;
        RECT 2362.020 2190.380 2365.020 2190.390 ;
        RECT 2542.020 2190.380 2545.020 2190.390 ;
        RECT 2722.020 2190.380 2725.020 2190.390 ;
        RECT 2902.020 2190.380 2905.020 2190.390 ;
        RECT 2936.000 2190.380 2939.000 2190.390 ;
        RECT -24.080 2187.380 2943.700 2190.380 ;
        RECT -19.380 2187.370 -16.380 2187.380 ;
        RECT 22.020 2187.370 25.020 2187.380 ;
        RECT 202.020 2187.370 205.020 2187.380 ;
        RECT 321.040 2187.370 322.640 2187.380 ;
        RECT 1462.020 2187.370 1465.020 2187.380 ;
        RECT 1642.020 2187.370 1645.020 2187.380 ;
        RECT 1822.020 2187.370 1825.020 2187.380 ;
        RECT 2002.020 2187.370 2005.020 2187.380 ;
        RECT 2182.020 2187.370 2185.020 2187.380 ;
        RECT 2362.020 2187.370 2365.020 2187.380 ;
        RECT 2542.020 2187.370 2545.020 2187.380 ;
        RECT 2722.020 2187.370 2725.020 2187.380 ;
        RECT 2902.020 2187.370 2905.020 2187.380 ;
        RECT 2936.000 2187.370 2939.000 2187.380 ;
        RECT -9.980 2172.380 -6.980 2172.390 ;
        RECT 4.020 2172.380 7.020 2172.390 ;
        RECT 184.020 2172.380 187.020 2172.390 ;
        RECT 321.040 2172.380 322.640 2172.390 ;
        RECT 1444.020 2172.380 1447.020 2172.390 ;
        RECT 1624.020 2172.380 1627.020 2172.390 ;
        RECT 1804.020 2172.380 1807.020 2172.390 ;
        RECT 1984.020 2172.380 1987.020 2172.390 ;
        RECT 2164.020 2172.380 2167.020 2172.390 ;
        RECT 2344.020 2172.380 2347.020 2172.390 ;
        RECT 2524.020 2172.380 2527.020 2172.390 ;
        RECT 2704.020 2172.380 2707.020 2172.390 ;
        RECT 2884.020 2172.380 2887.020 2172.390 ;
        RECT 2926.600 2172.380 2929.600 2172.390 ;
        RECT -14.680 2169.380 2934.300 2172.380 ;
        RECT -9.980 2169.370 -6.980 2169.380 ;
        RECT 4.020 2169.370 7.020 2169.380 ;
        RECT 184.020 2169.370 187.020 2169.380 ;
        RECT 321.040 2169.370 322.640 2169.380 ;
        RECT 1444.020 2169.370 1447.020 2169.380 ;
        RECT 1624.020 2169.370 1627.020 2169.380 ;
        RECT 1804.020 2169.370 1807.020 2169.380 ;
        RECT 1984.020 2169.370 1987.020 2169.380 ;
        RECT 2164.020 2169.370 2167.020 2169.380 ;
        RECT 2344.020 2169.370 2347.020 2169.380 ;
        RECT 2524.020 2169.370 2527.020 2169.380 ;
        RECT 2704.020 2169.370 2707.020 2169.380 ;
        RECT 2884.020 2169.370 2887.020 2169.380 ;
        RECT 2926.600 2169.370 2929.600 2169.380 ;
        RECT -38.180 2046.380 -35.180 2046.390 ;
        RECT 58.020 2046.380 61.020 2046.390 ;
        RECT 238.020 2046.380 241.020 2046.390 ;
        RECT 321.040 2046.380 322.640 2046.390 ;
        RECT 1498.020 2046.380 1501.020 2046.390 ;
        RECT 1678.020 2046.380 1681.020 2046.390 ;
        RECT 1858.020 2046.380 1861.020 2046.390 ;
        RECT 2038.020 2046.380 2041.020 2046.390 ;
        RECT 2218.020 2046.380 2221.020 2046.390 ;
        RECT 2398.020 2046.380 2401.020 2046.390 ;
        RECT 2578.020 2046.380 2581.020 2046.390 ;
        RECT 2758.020 2046.380 2761.020 2046.390 ;
        RECT 2954.800 2046.380 2957.800 2046.390 ;
        RECT -42.880 2043.380 2962.500 2046.380 ;
        RECT -38.180 2043.370 -35.180 2043.380 ;
        RECT 58.020 2043.370 61.020 2043.380 ;
        RECT 238.020 2043.370 241.020 2043.380 ;
        RECT 321.040 2043.370 322.640 2043.380 ;
        RECT 1498.020 2043.370 1501.020 2043.380 ;
        RECT 1678.020 2043.370 1681.020 2043.380 ;
        RECT 1858.020 2043.370 1861.020 2043.380 ;
        RECT 2038.020 2043.370 2041.020 2043.380 ;
        RECT 2218.020 2043.370 2221.020 2043.380 ;
        RECT 2398.020 2043.370 2401.020 2043.380 ;
        RECT 2578.020 2043.370 2581.020 2043.380 ;
        RECT 2758.020 2043.370 2761.020 2043.380 ;
        RECT 2954.800 2043.370 2957.800 2043.380 ;
        RECT -28.780 2028.380 -25.780 2028.390 ;
        RECT 40.020 2028.380 43.020 2028.390 ;
        RECT 220.020 2028.380 223.020 2028.390 ;
        RECT 321.040 2028.380 322.640 2028.390 ;
        RECT 1480.020 2028.380 1483.020 2028.390 ;
        RECT 1660.020 2028.380 1663.020 2028.390 ;
        RECT 1840.020 2028.380 1843.020 2028.390 ;
        RECT 2020.020 2028.380 2023.020 2028.390 ;
        RECT 2200.020 2028.380 2203.020 2028.390 ;
        RECT 2380.020 2028.380 2383.020 2028.390 ;
        RECT 2560.020 2028.380 2563.020 2028.390 ;
        RECT 2740.020 2028.380 2743.020 2028.390 ;
        RECT 2945.400 2028.380 2948.400 2028.390 ;
        RECT -33.480 2025.380 2953.100 2028.380 ;
        RECT -28.780 2025.370 -25.780 2025.380 ;
        RECT 40.020 2025.370 43.020 2025.380 ;
        RECT 220.020 2025.370 223.020 2025.380 ;
        RECT 321.040 2025.370 322.640 2025.380 ;
        RECT 1480.020 2025.370 1483.020 2025.380 ;
        RECT 1660.020 2025.370 1663.020 2025.380 ;
        RECT 1840.020 2025.370 1843.020 2025.380 ;
        RECT 2020.020 2025.370 2023.020 2025.380 ;
        RECT 2200.020 2025.370 2203.020 2025.380 ;
        RECT 2380.020 2025.370 2383.020 2025.380 ;
        RECT 2560.020 2025.370 2563.020 2025.380 ;
        RECT 2740.020 2025.370 2743.020 2025.380 ;
        RECT 2945.400 2025.370 2948.400 2025.380 ;
        RECT -19.380 2010.380 -16.380 2010.390 ;
        RECT 22.020 2010.380 25.020 2010.390 ;
        RECT 202.020 2010.380 205.020 2010.390 ;
        RECT 321.040 2010.380 322.640 2010.390 ;
        RECT 1462.020 2010.380 1465.020 2010.390 ;
        RECT 1642.020 2010.380 1645.020 2010.390 ;
        RECT 1822.020 2010.380 1825.020 2010.390 ;
        RECT 2002.020 2010.380 2005.020 2010.390 ;
        RECT 2182.020 2010.380 2185.020 2010.390 ;
        RECT 2362.020 2010.380 2365.020 2010.390 ;
        RECT 2542.020 2010.380 2545.020 2010.390 ;
        RECT 2722.020 2010.380 2725.020 2010.390 ;
        RECT 2902.020 2010.380 2905.020 2010.390 ;
        RECT 2936.000 2010.380 2939.000 2010.390 ;
        RECT -24.080 2007.380 2943.700 2010.380 ;
        RECT -19.380 2007.370 -16.380 2007.380 ;
        RECT 22.020 2007.370 25.020 2007.380 ;
        RECT 202.020 2007.370 205.020 2007.380 ;
        RECT 321.040 2007.370 322.640 2007.380 ;
        RECT 1462.020 2007.370 1465.020 2007.380 ;
        RECT 1642.020 2007.370 1645.020 2007.380 ;
        RECT 1822.020 2007.370 1825.020 2007.380 ;
        RECT 2002.020 2007.370 2005.020 2007.380 ;
        RECT 2182.020 2007.370 2185.020 2007.380 ;
        RECT 2362.020 2007.370 2365.020 2007.380 ;
        RECT 2542.020 2007.370 2545.020 2007.380 ;
        RECT 2722.020 2007.370 2725.020 2007.380 ;
        RECT 2902.020 2007.370 2905.020 2007.380 ;
        RECT 2936.000 2007.370 2939.000 2007.380 ;
        RECT -9.980 1992.380 -6.980 1992.390 ;
        RECT 4.020 1992.380 7.020 1992.390 ;
        RECT 184.020 1992.380 187.020 1992.390 ;
        RECT 321.040 1992.380 322.640 1992.390 ;
        RECT 1444.020 1992.380 1447.020 1992.390 ;
        RECT 1624.020 1992.380 1627.020 1992.390 ;
        RECT 1804.020 1992.380 1807.020 1992.390 ;
        RECT 1984.020 1992.380 1987.020 1992.390 ;
        RECT 2164.020 1992.380 2167.020 1992.390 ;
        RECT 2344.020 1992.380 2347.020 1992.390 ;
        RECT 2524.020 1992.380 2527.020 1992.390 ;
        RECT 2704.020 1992.380 2707.020 1992.390 ;
        RECT 2884.020 1992.380 2887.020 1992.390 ;
        RECT 2926.600 1992.380 2929.600 1992.390 ;
        RECT -14.680 1989.380 2934.300 1992.380 ;
        RECT -9.980 1989.370 -6.980 1989.380 ;
        RECT 4.020 1989.370 7.020 1989.380 ;
        RECT 184.020 1989.370 187.020 1989.380 ;
        RECT 321.040 1989.370 322.640 1989.380 ;
        RECT 1444.020 1989.370 1447.020 1989.380 ;
        RECT 1624.020 1989.370 1627.020 1989.380 ;
        RECT 1804.020 1989.370 1807.020 1989.380 ;
        RECT 1984.020 1989.370 1987.020 1989.380 ;
        RECT 2164.020 1989.370 2167.020 1989.380 ;
        RECT 2344.020 1989.370 2347.020 1989.380 ;
        RECT 2524.020 1989.370 2527.020 1989.380 ;
        RECT 2704.020 1989.370 2707.020 1989.380 ;
        RECT 2884.020 1989.370 2887.020 1989.380 ;
        RECT 2926.600 1989.370 2929.600 1989.380 ;
        RECT -38.180 1866.380 -35.180 1866.390 ;
        RECT 58.020 1866.380 61.020 1866.390 ;
        RECT 238.020 1866.380 241.020 1866.390 ;
        RECT 321.040 1866.380 322.640 1866.390 ;
        RECT 1498.020 1866.380 1501.020 1866.390 ;
        RECT 1678.020 1866.380 1681.020 1866.390 ;
        RECT 1858.020 1866.380 1861.020 1866.390 ;
        RECT 2038.020 1866.380 2041.020 1866.390 ;
        RECT 2218.020 1866.380 2221.020 1866.390 ;
        RECT 2398.020 1866.380 2401.020 1866.390 ;
        RECT 2578.020 1866.380 2581.020 1866.390 ;
        RECT 2758.020 1866.380 2761.020 1866.390 ;
        RECT 2954.800 1866.380 2957.800 1866.390 ;
        RECT -42.880 1863.380 2962.500 1866.380 ;
        RECT -38.180 1863.370 -35.180 1863.380 ;
        RECT 58.020 1863.370 61.020 1863.380 ;
        RECT 238.020 1863.370 241.020 1863.380 ;
        RECT 321.040 1863.370 322.640 1863.380 ;
        RECT 1498.020 1863.370 1501.020 1863.380 ;
        RECT 1678.020 1863.370 1681.020 1863.380 ;
        RECT 1858.020 1863.370 1861.020 1863.380 ;
        RECT 2038.020 1863.370 2041.020 1863.380 ;
        RECT 2218.020 1863.370 2221.020 1863.380 ;
        RECT 2398.020 1863.370 2401.020 1863.380 ;
        RECT 2578.020 1863.370 2581.020 1863.380 ;
        RECT 2758.020 1863.370 2761.020 1863.380 ;
        RECT 2954.800 1863.370 2957.800 1863.380 ;
        RECT -28.780 1848.380 -25.780 1848.390 ;
        RECT 40.020 1848.380 43.020 1848.390 ;
        RECT 220.020 1848.380 223.020 1848.390 ;
        RECT 321.040 1848.380 322.640 1848.390 ;
        RECT 1480.020 1848.380 1483.020 1848.390 ;
        RECT 1660.020 1848.380 1663.020 1848.390 ;
        RECT 1840.020 1848.380 1843.020 1848.390 ;
        RECT 2020.020 1848.380 2023.020 1848.390 ;
        RECT 2200.020 1848.380 2203.020 1848.390 ;
        RECT 2380.020 1848.380 2383.020 1848.390 ;
        RECT 2560.020 1848.380 2563.020 1848.390 ;
        RECT 2740.020 1848.380 2743.020 1848.390 ;
        RECT 2945.400 1848.380 2948.400 1848.390 ;
        RECT -33.480 1845.380 2953.100 1848.380 ;
        RECT -28.780 1845.370 -25.780 1845.380 ;
        RECT 40.020 1845.370 43.020 1845.380 ;
        RECT 220.020 1845.370 223.020 1845.380 ;
        RECT 321.040 1845.370 322.640 1845.380 ;
        RECT 1480.020 1845.370 1483.020 1845.380 ;
        RECT 1660.020 1845.370 1663.020 1845.380 ;
        RECT 1840.020 1845.370 1843.020 1845.380 ;
        RECT 2020.020 1845.370 2023.020 1845.380 ;
        RECT 2200.020 1845.370 2203.020 1845.380 ;
        RECT 2380.020 1845.370 2383.020 1845.380 ;
        RECT 2560.020 1845.370 2563.020 1845.380 ;
        RECT 2740.020 1845.370 2743.020 1845.380 ;
        RECT 2945.400 1845.370 2948.400 1845.380 ;
        RECT -19.380 1830.380 -16.380 1830.390 ;
        RECT 22.020 1830.380 25.020 1830.390 ;
        RECT 202.020 1830.380 205.020 1830.390 ;
        RECT 321.040 1830.380 322.640 1830.390 ;
        RECT 1462.020 1830.380 1465.020 1830.390 ;
        RECT 1642.020 1830.380 1645.020 1830.390 ;
        RECT 1822.020 1830.380 1825.020 1830.390 ;
        RECT 2002.020 1830.380 2005.020 1830.390 ;
        RECT 2182.020 1830.380 2185.020 1830.390 ;
        RECT 2362.020 1830.380 2365.020 1830.390 ;
        RECT 2542.020 1830.380 2545.020 1830.390 ;
        RECT 2722.020 1830.380 2725.020 1830.390 ;
        RECT 2902.020 1830.380 2905.020 1830.390 ;
        RECT 2936.000 1830.380 2939.000 1830.390 ;
        RECT -24.080 1827.380 2943.700 1830.380 ;
        RECT -19.380 1827.370 -16.380 1827.380 ;
        RECT 22.020 1827.370 25.020 1827.380 ;
        RECT 202.020 1827.370 205.020 1827.380 ;
        RECT 321.040 1827.370 322.640 1827.380 ;
        RECT 1462.020 1827.370 1465.020 1827.380 ;
        RECT 1642.020 1827.370 1645.020 1827.380 ;
        RECT 1822.020 1827.370 1825.020 1827.380 ;
        RECT 2002.020 1827.370 2005.020 1827.380 ;
        RECT 2182.020 1827.370 2185.020 1827.380 ;
        RECT 2362.020 1827.370 2365.020 1827.380 ;
        RECT 2542.020 1827.370 2545.020 1827.380 ;
        RECT 2722.020 1827.370 2725.020 1827.380 ;
        RECT 2902.020 1827.370 2905.020 1827.380 ;
        RECT 2936.000 1827.370 2939.000 1827.380 ;
        RECT -9.980 1812.380 -6.980 1812.390 ;
        RECT 4.020 1812.380 7.020 1812.390 ;
        RECT 184.020 1812.380 187.020 1812.390 ;
        RECT 321.040 1812.380 322.640 1812.390 ;
        RECT 1444.020 1812.380 1447.020 1812.390 ;
        RECT 1624.020 1812.380 1627.020 1812.390 ;
        RECT 1804.020 1812.380 1807.020 1812.390 ;
        RECT 1984.020 1812.380 1987.020 1812.390 ;
        RECT 2164.020 1812.380 2167.020 1812.390 ;
        RECT 2344.020 1812.380 2347.020 1812.390 ;
        RECT 2524.020 1812.380 2527.020 1812.390 ;
        RECT 2704.020 1812.380 2707.020 1812.390 ;
        RECT 2884.020 1812.380 2887.020 1812.390 ;
        RECT 2926.600 1812.380 2929.600 1812.390 ;
        RECT -14.680 1809.380 2934.300 1812.380 ;
        RECT -9.980 1809.370 -6.980 1809.380 ;
        RECT 4.020 1809.370 7.020 1809.380 ;
        RECT 184.020 1809.370 187.020 1809.380 ;
        RECT 321.040 1809.370 322.640 1809.380 ;
        RECT 1444.020 1809.370 1447.020 1809.380 ;
        RECT 1624.020 1809.370 1627.020 1809.380 ;
        RECT 1804.020 1809.370 1807.020 1809.380 ;
        RECT 1984.020 1809.370 1987.020 1809.380 ;
        RECT 2164.020 1809.370 2167.020 1809.380 ;
        RECT 2344.020 1809.370 2347.020 1809.380 ;
        RECT 2524.020 1809.370 2527.020 1809.380 ;
        RECT 2704.020 1809.370 2707.020 1809.380 ;
        RECT 2884.020 1809.370 2887.020 1809.380 ;
        RECT 2926.600 1809.370 2929.600 1809.380 ;
        RECT -38.180 1686.380 -35.180 1686.390 ;
        RECT 58.020 1686.380 61.020 1686.390 ;
        RECT 238.020 1686.380 241.020 1686.390 ;
        RECT 321.040 1686.380 322.640 1686.390 ;
        RECT 1498.020 1686.380 1501.020 1686.390 ;
        RECT 1678.020 1686.380 1681.020 1686.390 ;
        RECT 1858.020 1686.380 1861.020 1686.390 ;
        RECT 2038.020 1686.380 2041.020 1686.390 ;
        RECT 2218.020 1686.380 2221.020 1686.390 ;
        RECT 2398.020 1686.380 2401.020 1686.390 ;
        RECT 2578.020 1686.380 2581.020 1686.390 ;
        RECT 2758.020 1686.380 2761.020 1686.390 ;
        RECT 2954.800 1686.380 2957.800 1686.390 ;
        RECT -42.880 1683.380 2962.500 1686.380 ;
        RECT -38.180 1683.370 -35.180 1683.380 ;
        RECT 58.020 1683.370 61.020 1683.380 ;
        RECT 238.020 1683.370 241.020 1683.380 ;
        RECT 321.040 1683.370 322.640 1683.380 ;
        RECT 1498.020 1683.370 1501.020 1683.380 ;
        RECT 1678.020 1683.370 1681.020 1683.380 ;
        RECT 1858.020 1683.370 1861.020 1683.380 ;
        RECT 2038.020 1683.370 2041.020 1683.380 ;
        RECT 2218.020 1683.370 2221.020 1683.380 ;
        RECT 2398.020 1683.370 2401.020 1683.380 ;
        RECT 2578.020 1683.370 2581.020 1683.380 ;
        RECT 2758.020 1683.370 2761.020 1683.380 ;
        RECT 2954.800 1683.370 2957.800 1683.380 ;
        RECT -28.780 1668.380 -25.780 1668.390 ;
        RECT 40.020 1668.380 43.020 1668.390 ;
        RECT 220.020 1668.380 223.020 1668.390 ;
        RECT 321.040 1668.380 322.640 1668.390 ;
        RECT 1480.020 1668.380 1483.020 1668.390 ;
        RECT 1660.020 1668.380 1663.020 1668.390 ;
        RECT 1840.020 1668.380 1843.020 1668.390 ;
        RECT 2020.020 1668.380 2023.020 1668.390 ;
        RECT 2200.020 1668.380 2203.020 1668.390 ;
        RECT 2380.020 1668.380 2383.020 1668.390 ;
        RECT 2560.020 1668.380 2563.020 1668.390 ;
        RECT 2740.020 1668.380 2743.020 1668.390 ;
        RECT 2945.400 1668.380 2948.400 1668.390 ;
        RECT -33.480 1665.380 2953.100 1668.380 ;
        RECT -28.780 1665.370 -25.780 1665.380 ;
        RECT 40.020 1665.370 43.020 1665.380 ;
        RECT 220.020 1665.370 223.020 1665.380 ;
        RECT 321.040 1665.370 322.640 1665.380 ;
        RECT 1480.020 1665.370 1483.020 1665.380 ;
        RECT 1660.020 1665.370 1663.020 1665.380 ;
        RECT 1840.020 1665.370 1843.020 1665.380 ;
        RECT 2020.020 1665.370 2023.020 1665.380 ;
        RECT 2200.020 1665.370 2203.020 1665.380 ;
        RECT 2380.020 1665.370 2383.020 1665.380 ;
        RECT 2560.020 1665.370 2563.020 1665.380 ;
        RECT 2740.020 1665.370 2743.020 1665.380 ;
        RECT 2945.400 1665.370 2948.400 1665.380 ;
        RECT -19.380 1650.380 -16.380 1650.390 ;
        RECT 22.020 1650.380 25.020 1650.390 ;
        RECT 202.020 1650.380 205.020 1650.390 ;
        RECT 321.040 1650.380 322.640 1650.390 ;
        RECT 1462.020 1650.380 1465.020 1650.390 ;
        RECT 1642.020 1650.380 1645.020 1650.390 ;
        RECT 1822.020 1650.380 1825.020 1650.390 ;
        RECT 2002.020 1650.380 2005.020 1650.390 ;
        RECT 2182.020 1650.380 2185.020 1650.390 ;
        RECT 2362.020 1650.380 2365.020 1650.390 ;
        RECT 2542.020 1650.380 2545.020 1650.390 ;
        RECT 2722.020 1650.380 2725.020 1650.390 ;
        RECT 2902.020 1650.380 2905.020 1650.390 ;
        RECT 2936.000 1650.380 2939.000 1650.390 ;
        RECT -24.080 1647.380 2943.700 1650.380 ;
        RECT -19.380 1647.370 -16.380 1647.380 ;
        RECT 22.020 1647.370 25.020 1647.380 ;
        RECT 202.020 1647.370 205.020 1647.380 ;
        RECT 321.040 1647.370 322.640 1647.380 ;
        RECT 1462.020 1647.370 1465.020 1647.380 ;
        RECT 1642.020 1647.370 1645.020 1647.380 ;
        RECT 1822.020 1647.370 1825.020 1647.380 ;
        RECT 2002.020 1647.370 2005.020 1647.380 ;
        RECT 2182.020 1647.370 2185.020 1647.380 ;
        RECT 2362.020 1647.370 2365.020 1647.380 ;
        RECT 2542.020 1647.370 2545.020 1647.380 ;
        RECT 2722.020 1647.370 2725.020 1647.380 ;
        RECT 2902.020 1647.370 2905.020 1647.380 ;
        RECT 2936.000 1647.370 2939.000 1647.380 ;
        RECT -9.980 1632.380 -6.980 1632.390 ;
        RECT 4.020 1632.380 7.020 1632.390 ;
        RECT 184.020 1632.380 187.020 1632.390 ;
        RECT 321.040 1632.380 322.640 1632.390 ;
        RECT 1444.020 1632.380 1447.020 1632.390 ;
        RECT 1624.020 1632.380 1627.020 1632.390 ;
        RECT 1804.020 1632.380 1807.020 1632.390 ;
        RECT 1984.020 1632.380 1987.020 1632.390 ;
        RECT 2164.020 1632.380 2167.020 1632.390 ;
        RECT 2344.020 1632.380 2347.020 1632.390 ;
        RECT 2524.020 1632.380 2527.020 1632.390 ;
        RECT 2704.020 1632.380 2707.020 1632.390 ;
        RECT 2884.020 1632.380 2887.020 1632.390 ;
        RECT 2926.600 1632.380 2929.600 1632.390 ;
        RECT -14.680 1629.380 2934.300 1632.380 ;
        RECT -9.980 1629.370 -6.980 1629.380 ;
        RECT 4.020 1629.370 7.020 1629.380 ;
        RECT 184.020 1629.370 187.020 1629.380 ;
        RECT 321.040 1629.370 322.640 1629.380 ;
        RECT 1444.020 1629.370 1447.020 1629.380 ;
        RECT 1624.020 1629.370 1627.020 1629.380 ;
        RECT 1804.020 1629.370 1807.020 1629.380 ;
        RECT 1984.020 1629.370 1987.020 1629.380 ;
        RECT 2164.020 1629.370 2167.020 1629.380 ;
        RECT 2344.020 1629.370 2347.020 1629.380 ;
        RECT 2524.020 1629.370 2527.020 1629.380 ;
        RECT 2704.020 1629.370 2707.020 1629.380 ;
        RECT 2884.020 1629.370 2887.020 1629.380 ;
        RECT 2926.600 1629.370 2929.600 1629.380 ;
        RECT -38.180 1506.380 -35.180 1506.390 ;
        RECT 58.020 1506.380 61.020 1506.390 ;
        RECT 238.020 1506.380 241.020 1506.390 ;
        RECT 1498.020 1506.380 1501.020 1506.390 ;
        RECT 1678.020 1506.380 1681.020 1506.390 ;
        RECT 1858.020 1506.380 1861.020 1506.390 ;
        RECT 2038.020 1506.380 2041.020 1506.390 ;
        RECT 2218.020 1506.380 2221.020 1506.390 ;
        RECT 2398.020 1506.380 2401.020 1506.390 ;
        RECT 2578.020 1506.380 2581.020 1506.390 ;
        RECT 2758.020 1506.380 2761.020 1506.390 ;
        RECT 2954.800 1506.380 2957.800 1506.390 ;
        RECT -42.880 1503.380 2962.500 1506.380 ;
        RECT -38.180 1503.370 -35.180 1503.380 ;
        RECT 58.020 1503.370 61.020 1503.380 ;
        RECT 238.020 1503.370 241.020 1503.380 ;
        RECT 1498.020 1503.370 1501.020 1503.380 ;
        RECT 1678.020 1503.370 1681.020 1503.380 ;
        RECT 1858.020 1503.370 1861.020 1503.380 ;
        RECT 2038.020 1503.370 2041.020 1503.380 ;
        RECT 2218.020 1503.370 2221.020 1503.380 ;
        RECT 2398.020 1503.370 2401.020 1503.380 ;
        RECT 2578.020 1503.370 2581.020 1503.380 ;
        RECT 2758.020 1503.370 2761.020 1503.380 ;
        RECT 2954.800 1503.370 2957.800 1503.380 ;
        RECT -28.780 1488.380 -25.780 1488.390 ;
        RECT 40.020 1488.380 43.020 1488.390 ;
        RECT 220.020 1488.380 223.020 1488.390 ;
        RECT 1480.020 1488.380 1483.020 1488.390 ;
        RECT 1660.020 1488.380 1663.020 1488.390 ;
        RECT 1840.020 1488.380 1843.020 1488.390 ;
        RECT 2020.020 1488.380 2023.020 1488.390 ;
        RECT 2200.020 1488.380 2203.020 1488.390 ;
        RECT 2380.020 1488.380 2383.020 1488.390 ;
        RECT 2560.020 1488.380 2563.020 1488.390 ;
        RECT 2740.020 1488.380 2743.020 1488.390 ;
        RECT 2945.400 1488.380 2948.400 1488.390 ;
        RECT -33.480 1485.380 2953.100 1488.380 ;
        RECT -28.780 1485.370 -25.780 1485.380 ;
        RECT 40.020 1485.370 43.020 1485.380 ;
        RECT 220.020 1485.370 223.020 1485.380 ;
        RECT 1480.020 1485.370 1483.020 1485.380 ;
        RECT 1660.020 1485.370 1663.020 1485.380 ;
        RECT 1840.020 1485.370 1843.020 1485.380 ;
        RECT 2020.020 1485.370 2023.020 1485.380 ;
        RECT 2200.020 1485.370 2203.020 1485.380 ;
        RECT 2380.020 1485.370 2383.020 1485.380 ;
        RECT 2560.020 1485.370 2563.020 1485.380 ;
        RECT 2740.020 1485.370 2743.020 1485.380 ;
        RECT 2945.400 1485.370 2948.400 1485.380 ;
        RECT -19.380 1470.380 -16.380 1470.390 ;
        RECT 22.020 1470.380 25.020 1470.390 ;
        RECT 202.020 1470.380 205.020 1470.390 ;
        RECT 382.020 1470.380 385.020 1470.390 ;
        RECT 562.020 1470.380 565.020 1470.390 ;
        RECT 742.020 1470.380 745.020 1470.390 ;
        RECT 922.020 1470.380 925.020 1470.390 ;
        RECT 1102.020 1470.380 1105.020 1470.390 ;
        RECT 1282.020 1470.380 1285.020 1470.390 ;
        RECT 1462.020 1470.380 1465.020 1470.390 ;
        RECT 1642.020 1470.380 1645.020 1470.390 ;
        RECT 1822.020 1470.380 1825.020 1470.390 ;
        RECT 2002.020 1470.380 2005.020 1470.390 ;
        RECT 2182.020 1470.380 2185.020 1470.390 ;
        RECT 2362.020 1470.380 2365.020 1470.390 ;
        RECT 2542.020 1470.380 2545.020 1470.390 ;
        RECT 2722.020 1470.380 2725.020 1470.390 ;
        RECT 2902.020 1470.380 2905.020 1470.390 ;
        RECT 2936.000 1470.380 2939.000 1470.390 ;
        RECT -24.080 1467.380 2943.700 1470.380 ;
        RECT -19.380 1467.370 -16.380 1467.380 ;
        RECT 22.020 1467.370 25.020 1467.380 ;
        RECT 202.020 1467.370 205.020 1467.380 ;
        RECT 382.020 1467.370 385.020 1467.380 ;
        RECT 562.020 1467.370 565.020 1467.380 ;
        RECT 742.020 1467.370 745.020 1467.380 ;
        RECT 922.020 1467.370 925.020 1467.380 ;
        RECT 1102.020 1467.370 1105.020 1467.380 ;
        RECT 1282.020 1467.370 1285.020 1467.380 ;
        RECT 1462.020 1467.370 1465.020 1467.380 ;
        RECT 1642.020 1467.370 1645.020 1467.380 ;
        RECT 1822.020 1467.370 1825.020 1467.380 ;
        RECT 2002.020 1467.370 2005.020 1467.380 ;
        RECT 2182.020 1467.370 2185.020 1467.380 ;
        RECT 2362.020 1467.370 2365.020 1467.380 ;
        RECT 2542.020 1467.370 2545.020 1467.380 ;
        RECT 2722.020 1467.370 2725.020 1467.380 ;
        RECT 2902.020 1467.370 2905.020 1467.380 ;
        RECT 2936.000 1467.370 2939.000 1467.380 ;
        RECT -9.980 1452.380 -6.980 1452.390 ;
        RECT 4.020 1452.380 7.020 1452.390 ;
        RECT 184.020 1452.380 187.020 1452.390 ;
        RECT 364.020 1452.380 367.020 1452.390 ;
        RECT 544.020 1452.380 547.020 1452.390 ;
        RECT 724.020 1452.380 727.020 1452.390 ;
        RECT 904.020 1452.380 907.020 1452.390 ;
        RECT 1084.020 1452.380 1087.020 1452.390 ;
        RECT 1264.020 1452.380 1267.020 1452.390 ;
        RECT 1444.020 1452.380 1447.020 1452.390 ;
        RECT 1624.020 1452.380 1627.020 1452.390 ;
        RECT 1804.020 1452.380 1807.020 1452.390 ;
        RECT 1984.020 1452.380 1987.020 1452.390 ;
        RECT 2164.020 1452.380 2167.020 1452.390 ;
        RECT 2344.020 1452.380 2347.020 1452.390 ;
        RECT 2524.020 1452.380 2527.020 1452.390 ;
        RECT 2704.020 1452.380 2707.020 1452.390 ;
        RECT 2884.020 1452.380 2887.020 1452.390 ;
        RECT 2926.600 1452.380 2929.600 1452.390 ;
        RECT -14.680 1449.380 2934.300 1452.380 ;
        RECT -9.980 1449.370 -6.980 1449.380 ;
        RECT 4.020 1449.370 7.020 1449.380 ;
        RECT 184.020 1449.370 187.020 1449.380 ;
        RECT 364.020 1449.370 367.020 1449.380 ;
        RECT 544.020 1449.370 547.020 1449.380 ;
        RECT 724.020 1449.370 727.020 1449.380 ;
        RECT 904.020 1449.370 907.020 1449.380 ;
        RECT 1084.020 1449.370 1087.020 1449.380 ;
        RECT 1264.020 1449.370 1267.020 1449.380 ;
        RECT 1444.020 1449.370 1447.020 1449.380 ;
        RECT 1624.020 1449.370 1627.020 1449.380 ;
        RECT 1804.020 1449.370 1807.020 1449.380 ;
        RECT 1984.020 1449.370 1987.020 1449.380 ;
        RECT 2164.020 1449.370 2167.020 1449.380 ;
        RECT 2344.020 1449.370 2347.020 1449.380 ;
        RECT 2524.020 1449.370 2527.020 1449.380 ;
        RECT 2704.020 1449.370 2707.020 1449.380 ;
        RECT 2884.020 1449.370 2887.020 1449.380 ;
        RECT 2926.600 1449.370 2929.600 1449.380 ;
        RECT -38.180 1326.380 -35.180 1326.390 ;
        RECT 58.020 1326.380 61.020 1326.390 ;
        RECT 238.020 1326.380 241.020 1326.390 ;
        RECT 418.020 1326.380 421.020 1326.390 ;
        RECT 598.020 1326.380 601.020 1326.390 ;
        RECT 778.020 1326.380 781.020 1326.390 ;
        RECT 958.020 1326.380 961.020 1326.390 ;
        RECT 1138.020 1326.380 1141.020 1326.390 ;
        RECT 1318.020 1326.380 1321.020 1326.390 ;
        RECT 1498.020 1326.380 1501.020 1326.390 ;
        RECT 1678.020 1326.380 1681.020 1326.390 ;
        RECT 1858.020 1326.380 1861.020 1326.390 ;
        RECT 2038.020 1326.380 2041.020 1326.390 ;
        RECT 2218.020 1326.380 2221.020 1326.390 ;
        RECT 2398.020 1326.380 2401.020 1326.390 ;
        RECT 2578.020 1326.380 2581.020 1326.390 ;
        RECT 2758.020 1326.380 2761.020 1326.390 ;
        RECT 2954.800 1326.380 2957.800 1326.390 ;
        RECT -42.880 1323.380 2962.500 1326.380 ;
        RECT -38.180 1323.370 -35.180 1323.380 ;
        RECT 58.020 1323.370 61.020 1323.380 ;
        RECT 238.020 1323.370 241.020 1323.380 ;
        RECT 418.020 1323.370 421.020 1323.380 ;
        RECT 598.020 1323.370 601.020 1323.380 ;
        RECT 778.020 1323.370 781.020 1323.380 ;
        RECT 958.020 1323.370 961.020 1323.380 ;
        RECT 1138.020 1323.370 1141.020 1323.380 ;
        RECT 1318.020 1323.370 1321.020 1323.380 ;
        RECT 1498.020 1323.370 1501.020 1323.380 ;
        RECT 1678.020 1323.370 1681.020 1323.380 ;
        RECT 1858.020 1323.370 1861.020 1323.380 ;
        RECT 2038.020 1323.370 2041.020 1323.380 ;
        RECT 2218.020 1323.370 2221.020 1323.380 ;
        RECT 2398.020 1323.370 2401.020 1323.380 ;
        RECT 2578.020 1323.370 2581.020 1323.380 ;
        RECT 2758.020 1323.370 2761.020 1323.380 ;
        RECT 2954.800 1323.370 2957.800 1323.380 ;
        RECT -28.780 1308.380 -25.780 1308.390 ;
        RECT 40.020 1308.380 43.020 1308.390 ;
        RECT 220.020 1308.380 223.020 1308.390 ;
        RECT 400.020 1308.380 403.020 1308.390 ;
        RECT 580.020 1308.380 583.020 1308.390 ;
        RECT 760.020 1308.380 763.020 1308.390 ;
        RECT 940.020 1308.380 943.020 1308.390 ;
        RECT 1120.020 1308.380 1123.020 1308.390 ;
        RECT 1300.020 1308.380 1303.020 1308.390 ;
        RECT 1480.020 1308.380 1483.020 1308.390 ;
        RECT 1660.020 1308.380 1663.020 1308.390 ;
        RECT 1840.020 1308.380 1843.020 1308.390 ;
        RECT 2020.020 1308.380 2023.020 1308.390 ;
        RECT 2200.020 1308.380 2203.020 1308.390 ;
        RECT 2380.020 1308.380 2383.020 1308.390 ;
        RECT 2560.020 1308.380 2563.020 1308.390 ;
        RECT 2740.020 1308.380 2743.020 1308.390 ;
        RECT 2945.400 1308.380 2948.400 1308.390 ;
        RECT -33.480 1305.380 2953.100 1308.380 ;
        RECT -28.780 1305.370 -25.780 1305.380 ;
        RECT 40.020 1305.370 43.020 1305.380 ;
        RECT 220.020 1305.370 223.020 1305.380 ;
        RECT 400.020 1305.370 403.020 1305.380 ;
        RECT 580.020 1305.370 583.020 1305.380 ;
        RECT 760.020 1305.370 763.020 1305.380 ;
        RECT 940.020 1305.370 943.020 1305.380 ;
        RECT 1120.020 1305.370 1123.020 1305.380 ;
        RECT 1300.020 1305.370 1303.020 1305.380 ;
        RECT 1480.020 1305.370 1483.020 1305.380 ;
        RECT 1660.020 1305.370 1663.020 1305.380 ;
        RECT 1840.020 1305.370 1843.020 1305.380 ;
        RECT 2020.020 1305.370 2023.020 1305.380 ;
        RECT 2200.020 1305.370 2203.020 1305.380 ;
        RECT 2380.020 1305.370 2383.020 1305.380 ;
        RECT 2560.020 1305.370 2563.020 1305.380 ;
        RECT 2740.020 1305.370 2743.020 1305.380 ;
        RECT 2945.400 1305.370 2948.400 1305.380 ;
        RECT -19.380 1290.380 -16.380 1290.390 ;
        RECT 22.020 1290.380 25.020 1290.390 ;
        RECT 202.020 1290.380 205.020 1290.390 ;
        RECT 382.020 1290.380 385.020 1290.390 ;
        RECT 562.020 1290.380 565.020 1290.390 ;
        RECT 742.020 1290.380 745.020 1290.390 ;
        RECT 922.020 1290.380 925.020 1290.390 ;
        RECT 1102.020 1290.380 1105.020 1290.390 ;
        RECT 1282.020 1290.380 1285.020 1290.390 ;
        RECT 1462.020 1290.380 1465.020 1290.390 ;
        RECT 1642.020 1290.380 1645.020 1290.390 ;
        RECT 1822.020 1290.380 1825.020 1290.390 ;
        RECT 2002.020 1290.380 2005.020 1290.390 ;
        RECT 2182.020 1290.380 2185.020 1290.390 ;
        RECT 2362.020 1290.380 2365.020 1290.390 ;
        RECT 2542.020 1290.380 2545.020 1290.390 ;
        RECT 2722.020 1290.380 2725.020 1290.390 ;
        RECT 2902.020 1290.380 2905.020 1290.390 ;
        RECT 2936.000 1290.380 2939.000 1290.390 ;
        RECT -24.080 1287.380 2943.700 1290.380 ;
        RECT -19.380 1287.370 -16.380 1287.380 ;
        RECT 22.020 1287.370 25.020 1287.380 ;
        RECT 202.020 1287.370 205.020 1287.380 ;
        RECT 382.020 1287.370 385.020 1287.380 ;
        RECT 562.020 1287.370 565.020 1287.380 ;
        RECT 742.020 1287.370 745.020 1287.380 ;
        RECT 922.020 1287.370 925.020 1287.380 ;
        RECT 1102.020 1287.370 1105.020 1287.380 ;
        RECT 1282.020 1287.370 1285.020 1287.380 ;
        RECT 1462.020 1287.370 1465.020 1287.380 ;
        RECT 1642.020 1287.370 1645.020 1287.380 ;
        RECT 1822.020 1287.370 1825.020 1287.380 ;
        RECT 2002.020 1287.370 2005.020 1287.380 ;
        RECT 2182.020 1287.370 2185.020 1287.380 ;
        RECT 2362.020 1287.370 2365.020 1287.380 ;
        RECT 2542.020 1287.370 2545.020 1287.380 ;
        RECT 2722.020 1287.370 2725.020 1287.380 ;
        RECT 2902.020 1287.370 2905.020 1287.380 ;
        RECT 2936.000 1287.370 2939.000 1287.380 ;
        RECT -9.980 1272.380 -6.980 1272.390 ;
        RECT 4.020 1272.380 7.020 1272.390 ;
        RECT 184.020 1272.380 187.020 1272.390 ;
        RECT 364.020 1272.380 367.020 1272.390 ;
        RECT 544.020 1272.380 547.020 1272.390 ;
        RECT 724.020 1272.380 727.020 1272.390 ;
        RECT 904.020 1272.380 907.020 1272.390 ;
        RECT 1084.020 1272.380 1087.020 1272.390 ;
        RECT 1264.020 1272.380 1267.020 1272.390 ;
        RECT 1444.020 1272.380 1447.020 1272.390 ;
        RECT 1624.020 1272.380 1627.020 1272.390 ;
        RECT 1804.020 1272.380 1807.020 1272.390 ;
        RECT 1984.020 1272.380 1987.020 1272.390 ;
        RECT 2164.020 1272.380 2167.020 1272.390 ;
        RECT 2344.020 1272.380 2347.020 1272.390 ;
        RECT 2524.020 1272.380 2527.020 1272.390 ;
        RECT 2704.020 1272.380 2707.020 1272.390 ;
        RECT 2884.020 1272.380 2887.020 1272.390 ;
        RECT 2926.600 1272.380 2929.600 1272.390 ;
        RECT -14.680 1269.380 2934.300 1272.380 ;
        RECT -9.980 1269.370 -6.980 1269.380 ;
        RECT 4.020 1269.370 7.020 1269.380 ;
        RECT 184.020 1269.370 187.020 1269.380 ;
        RECT 364.020 1269.370 367.020 1269.380 ;
        RECT 544.020 1269.370 547.020 1269.380 ;
        RECT 724.020 1269.370 727.020 1269.380 ;
        RECT 904.020 1269.370 907.020 1269.380 ;
        RECT 1084.020 1269.370 1087.020 1269.380 ;
        RECT 1264.020 1269.370 1267.020 1269.380 ;
        RECT 1444.020 1269.370 1447.020 1269.380 ;
        RECT 1624.020 1269.370 1627.020 1269.380 ;
        RECT 1804.020 1269.370 1807.020 1269.380 ;
        RECT 1984.020 1269.370 1987.020 1269.380 ;
        RECT 2164.020 1269.370 2167.020 1269.380 ;
        RECT 2344.020 1269.370 2347.020 1269.380 ;
        RECT 2524.020 1269.370 2527.020 1269.380 ;
        RECT 2704.020 1269.370 2707.020 1269.380 ;
        RECT 2884.020 1269.370 2887.020 1269.380 ;
        RECT 2926.600 1269.370 2929.600 1269.380 ;
        RECT -38.180 1146.380 -35.180 1146.390 ;
        RECT 58.020 1146.380 61.020 1146.390 ;
        RECT 238.020 1146.380 241.020 1146.390 ;
        RECT 418.020 1146.380 421.020 1146.390 ;
        RECT 598.020 1146.380 601.020 1146.390 ;
        RECT 778.020 1146.380 781.020 1146.390 ;
        RECT 958.020 1146.380 961.020 1146.390 ;
        RECT 1138.020 1146.380 1141.020 1146.390 ;
        RECT 1318.020 1146.380 1321.020 1146.390 ;
        RECT 1498.020 1146.380 1501.020 1146.390 ;
        RECT 1678.020 1146.380 1681.020 1146.390 ;
        RECT 1858.020 1146.380 1861.020 1146.390 ;
        RECT 2038.020 1146.380 2041.020 1146.390 ;
        RECT 2218.020 1146.380 2221.020 1146.390 ;
        RECT 2398.020 1146.380 2401.020 1146.390 ;
        RECT 2578.020 1146.380 2581.020 1146.390 ;
        RECT 2758.020 1146.380 2761.020 1146.390 ;
        RECT 2954.800 1146.380 2957.800 1146.390 ;
        RECT -42.880 1143.380 2962.500 1146.380 ;
        RECT -38.180 1143.370 -35.180 1143.380 ;
        RECT 58.020 1143.370 61.020 1143.380 ;
        RECT 238.020 1143.370 241.020 1143.380 ;
        RECT 418.020 1143.370 421.020 1143.380 ;
        RECT 598.020 1143.370 601.020 1143.380 ;
        RECT 778.020 1143.370 781.020 1143.380 ;
        RECT 958.020 1143.370 961.020 1143.380 ;
        RECT 1138.020 1143.370 1141.020 1143.380 ;
        RECT 1318.020 1143.370 1321.020 1143.380 ;
        RECT 1498.020 1143.370 1501.020 1143.380 ;
        RECT 1678.020 1143.370 1681.020 1143.380 ;
        RECT 1858.020 1143.370 1861.020 1143.380 ;
        RECT 2038.020 1143.370 2041.020 1143.380 ;
        RECT 2218.020 1143.370 2221.020 1143.380 ;
        RECT 2398.020 1143.370 2401.020 1143.380 ;
        RECT 2578.020 1143.370 2581.020 1143.380 ;
        RECT 2758.020 1143.370 2761.020 1143.380 ;
        RECT 2954.800 1143.370 2957.800 1143.380 ;
        RECT -28.780 1128.380 -25.780 1128.390 ;
        RECT 40.020 1128.380 43.020 1128.390 ;
        RECT 220.020 1128.380 223.020 1128.390 ;
        RECT 400.020 1128.380 403.020 1128.390 ;
        RECT 580.020 1128.380 583.020 1128.390 ;
        RECT 760.020 1128.380 763.020 1128.390 ;
        RECT 940.020 1128.380 943.020 1128.390 ;
        RECT 1120.020 1128.380 1123.020 1128.390 ;
        RECT 1300.020 1128.380 1303.020 1128.390 ;
        RECT 1480.020 1128.380 1483.020 1128.390 ;
        RECT 1660.020 1128.380 1663.020 1128.390 ;
        RECT 1840.020 1128.380 1843.020 1128.390 ;
        RECT 2020.020 1128.380 2023.020 1128.390 ;
        RECT 2200.020 1128.380 2203.020 1128.390 ;
        RECT 2380.020 1128.380 2383.020 1128.390 ;
        RECT 2560.020 1128.380 2563.020 1128.390 ;
        RECT 2740.020 1128.380 2743.020 1128.390 ;
        RECT 2945.400 1128.380 2948.400 1128.390 ;
        RECT -33.480 1125.380 2953.100 1128.380 ;
        RECT -28.780 1125.370 -25.780 1125.380 ;
        RECT 40.020 1125.370 43.020 1125.380 ;
        RECT 220.020 1125.370 223.020 1125.380 ;
        RECT 400.020 1125.370 403.020 1125.380 ;
        RECT 580.020 1125.370 583.020 1125.380 ;
        RECT 760.020 1125.370 763.020 1125.380 ;
        RECT 940.020 1125.370 943.020 1125.380 ;
        RECT 1120.020 1125.370 1123.020 1125.380 ;
        RECT 1300.020 1125.370 1303.020 1125.380 ;
        RECT 1480.020 1125.370 1483.020 1125.380 ;
        RECT 1660.020 1125.370 1663.020 1125.380 ;
        RECT 1840.020 1125.370 1843.020 1125.380 ;
        RECT 2020.020 1125.370 2023.020 1125.380 ;
        RECT 2200.020 1125.370 2203.020 1125.380 ;
        RECT 2380.020 1125.370 2383.020 1125.380 ;
        RECT 2560.020 1125.370 2563.020 1125.380 ;
        RECT 2740.020 1125.370 2743.020 1125.380 ;
        RECT 2945.400 1125.370 2948.400 1125.380 ;
        RECT -19.380 1110.380 -16.380 1110.390 ;
        RECT 22.020 1110.380 25.020 1110.390 ;
        RECT 202.020 1110.380 205.020 1110.390 ;
        RECT 382.020 1110.380 385.020 1110.390 ;
        RECT 562.020 1110.380 565.020 1110.390 ;
        RECT 742.020 1110.380 745.020 1110.390 ;
        RECT 922.020 1110.380 925.020 1110.390 ;
        RECT 1102.020 1110.380 1105.020 1110.390 ;
        RECT 1282.020 1110.380 1285.020 1110.390 ;
        RECT 1462.020 1110.380 1465.020 1110.390 ;
        RECT 1642.020 1110.380 1645.020 1110.390 ;
        RECT 1822.020 1110.380 1825.020 1110.390 ;
        RECT 2002.020 1110.380 2005.020 1110.390 ;
        RECT 2182.020 1110.380 2185.020 1110.390 ;
        RECT 2362.020 1110.380 2365.020 1110.390 ;
        RECT 2542.020 1110.380 2545.020 1110.390 ;
        RECT 2722.020 1110.380 2725.020 1110.390 ;
        RECT 2902.020 1110.380 2905.020 1110.390 ;
        RECT 2936.000 1110.380 2939.000 1110.390 ;
        RECT -24.080 1107.380 2943.700 1110.380 ;
        RECT -19.380 1107.370 -16.380 1107.380 ;
        RECT 22.020 1107.370 25.020 1107.380 ;
        RECT 202.020 1107.370 205.020 1107.380 ;
        RECT 382.020 1107.370 385.020 1107.380 ;
        RECT 562.020 1107.370 565.020 1107.380 ;
        RECT 742.020 1107.370 745.020 1107.380 ;
        RECT 922.020 1107.370 925.020 1107.380 ;
        RECT 1102.020 1107.370 1105.020 1107.380 ;
        RECT 1282.020 1107.370 1285.020 1107.380 ;
        RECT 1462.020 1107.370 1465.020 1107.380 ;
        RECT 1642.020 1107.370 1645.020 1107.380 ;
        RECT 1822.020 1107.370 1825.020 1107.380 ;
        RECT 2002.020 1107.370 2005.020 1107.380 ;
        RECT 2182.020 1107.370 2185.020 1107.380 ;
        RECT 2362.020 1107.370 2365.020 1107.380 ;
        RECT 2542.020 1107.370 2545.020 1107.380 ;
        RECT 2722.020 1107.370 2725.020 1107.380 ;
        RECT 2902.020 1107.370 2905.020 1107.380 ;
        RECT 2936.000 1107.370 2939.000 1107.380 ;
        RECT -9.980 1092.380 -6.980 1092.390 ;
        RECT 4.020 1092.380 7.020 1092.390 ;
        RECT 184.020 1092.380 187.020 1092.390 ;
        RECT 364.020 1092.380 367.020 1092.390 ;
        RECT 544.020 1092.380 547.020 1092.390 ;
        RECT 724.020 1092.380 727.020 1092.390 ;
        RECT 904.020 1092.380 907.020 1092.390 ;
        RECT 1084.020 1092.380 1087.020 1092.390 ;
        RECT 1264.020 1092.380 1267.020 1092.390 ;
        RECT 1444.020 1092.380 1447.020 1092.390 ;
        RECT 1624.020 1092.380 1627.020 1092.390 ;
        RECT 1804.020 1092.380 1807.020 1092.390 ;
        RECT 1984.020 1092.380 1987.020 1092.390 ;
        RECT 2164.020 1092.380 2167.020 1092.390 ;
        RECT 2344.020 1092.380 2347.020 1092.390 ;
        RECT 2524.020 1092.380 2527.020 1092.390 ;
        RECT 2704.020 1092.380 2707.020 1092.390 ;
        RECT 2884.020 1092.380 2887.020 1092.390 ;
        RECT 2926.600 1092.380 2929.600 1092.390 ;
        RECT -14.680 1089.380 2934.300 1092.380 ;
        RECT -9.980 1089.370 -6.980 1089.380 ;
        RECT 4.020 1089.370 7.020 1089.380 ;
        RECT 184.020 1089.370 187.020 1089.380 ;
        RECT 364.020 1089.370 367.020 1089.380 ;
        RECT 544.020 1089.370 547.020 1089.380 ;
        RECT 724.020 1089.370 727.020 1089.380 ;
        RECT 904.020 1089.370 907.020 1089.380 ;
        RECT 1084.020 1089.370 1087.020 1089.380 ;
        RECT 1264.020 1089.370 1267.020 1089.380 ;
        RECT 1444.020 1089.370 1447.020 1089.380 ;
        RECT 1624.020 1089.370 1627.020 1089.380 ;
        RECT 1804.020 1089.370 1807.020 1089.380 ;
        RECT 1984.020 1089.370 1987.020 1089.380 ;
        RECT 2164.020 1089.370 2167.020 1089.380 ;
        RECT 2344.020 1089.370 2347.020 1089.380 ;
        RECT 2524.020 1089.370 2527.020 1089.380 ;
        RECT 2704.020 1089.370 2707.020 1089.380 ;
        RECT 2884.020 1089.370 2887.020 1089.380 ;
        RECT 2926.600 1089.370 2929.600 1089.380 ;
        RECT -38.180 966.380 -35.180 966.390 ;
        RECT 58.020 966.380 61.020 966.390 ;
        RECT 238.020 966.380 241.020 966.390 ;
        RECT 418.020 966.380 421.020 966.390 ;
        RECT 598.020 966.380 601.020 966.390 ;
        RECT 778.020 966.380 781.020 966.390 ;
        RECT 958.020 966.380 961.020 966.390 ;
        RECT 1138.020 966.380 1141.020 966.390 ;
        RECT 1318.020 966.380 1321.020 966.390 ;
        RECT 1498.020 966.380 1501.020 966.390 ;
        RECT 1678.020 966.380 1681.020 966.390 ;
        RECT 1858.020 966.380 1861.020 966.390 ;
        RECT 2038.020 966.380 2041.020 966.390 ;
        RECT 2218.020 966.380 2221.020 966.390 ;
        RECT 2398.020 966.380 2401.020 966.390 ;
        RECT 2578.020 966.380 2581.020 966.390 ;
        RECT 2758.020 966.380 2761.020 966.390 ;
        RECT 2954.800 966.380 2957.800 966.390 ;
        RECT -42.880 963.380 2962.500 966.380 ;
        RECT -38.180 963.370 -35.180 963.380 ;
        RECT 58.020 963.370 61.020 963.380 ;
        RECT 238.020 963.370 241.020 963.380 ;
        RECT 418.020 963.370 421.020 963.380 ;
        RECT 598.020 963.370 601.020 963.380 ;
        RECT 778.020 963.370 781.020 963.380 ;
        RECT 958.020 963.370 961.020 963.380 ;
        RECT 1138.020 963.370 1141.020 963.380 ;
        RECT 1318.020 963.370 1321.020 963.380 ;
        RECT 1498.020 963.370 1501.020 963.380 ;
        RECT 1678.020 963.370 1681.020 963.380 ;
        RECT 1858.020 963.370 1861.020 963.380 ;
        RECT 2038.020 963.370 2041.020 963.380 ;
        RECT 2218.020 963.370 2221.020 963.380 ;
        RECT 2398.020 963.370 2401.020 963.380 ;
        RECT 2578.020 963.370 2581.020 963.380 ;
        RECT 2758.020 963.370 2761.020 963.380 ;
        RECT 2954.800 963.370 2957.800 963.380 ;
        RECT -28.780 948.380 -25.780 948.390 ;
        RECT 40.020 948.380 43.020 948.390 ;
        RECT 220.020 948.380 223.020 948.390 ;
        RECT 400.020 948.380 403.020 948.390 ;
        RECT 580.020 948.380 583.020 948.390 ;
        RECT 760.020 948.380 763.020 948.390 ;
        RECT 940.020 948.380 943.020 948.390 ;
        RECT 1120.020 948.380 1123.020 948.390 ;
        RECT 1300.020 948.380 1303.020 948.390 ;
        RECT 1480.020 948.380 1483.020 948.390 ;
        RECT 1660.020 948.380 1663.020 948.390 ;
        RECT 1840.020 948.380 1843.020 948.390 ;
        RECT 2020.020 948.380 2023.020 948.390 ;
        RECT 2200.020 948.380 2203.020 948.390 ;
        RECT 2380.020 948.380 2383.020 948.390 ;
        RECT 2560.020 948.380 2563.020 948.390 ;
        RECT 2740.020 948.380 2743.020 948.390 ;
        RECT 2945.400 948.380 2948.400 948.390 ;
        RECT -33.480 945.380 2953.100 948.380 ;
        RECT -28.780 945.370 -25.780 945.380 ;
        RECT 40.020 945.370 43.020 945.380 ;
        RECT 220.020 945.370 223.020 945.380 ;
        RECT 400.020 945.370 403.020 945.380 ;
        RECT 580.020 945.370 583.020 945.380 ;
        RECT 760.020 945.370 763.020 945.380 ;
        RECT 940.020 945.370 943.020 945.380 ;
        RECT 1120.020 945.370 1123.020 945.380 ;
        RECT 1300.020 945.370 1303.020 945.380 ;
        RECT 1480.020 945.370 1483.020 945.380 ;
        RECT 1660.020 945.370 1663.020 945.380 ;
        RECT 1840.020 945.370 1843.020 945.380 ;
        RECT 2020.020 945.370 2023.020 945.380 ;
        RECT 2200.020 945.370 2203.020 945.380 ;
        RECT 2380.020 945.370 2383.020 945.380 ;
        RECT 2560.020 945.370 2563.020 945.380 ;
        RECT 2740.020 945.370 2743.020 945.380 ;
        RECT 2945.400 945.370 2948.400 945.380 ;
        RECT -19.380 930.380 -16.380 930.390 ;
        RECT 22.020 930.380 25.020 930.390 ;
        RECT 202.020 930.380 205.020 930.390 ;
        RECT 382.020 930.380 385.020 930.390 ;
        RECT 562.020 930.380 565.020 930.390 ;
        RECT 742.020 930.380 745.020 930.390 ;
        RECT 922.020 930.380 925.020 930.390 ;
        RECT 1102.020 930.380 1105.020 930.390 ;
        RECT 1282.020 930.380 1285.020 930.390 ;
        RECT 1462.020 930.380 1465.020 930.390 ;
        RECT 1642.020 930.380 1645.020 930.390 ;
        RECT 1822.020 930.380 1825.020 930.390 ;
        RECT 2002.020 930.380 2005.020 930.390 ;
        RECT 2182.020 930.380 2185.020 930.390 ;
        RECT 2362.020 930.380 2365.020 930.390 ;
        RECT 2542.020 930.380 2545.020 930.390 ;
        RECT 2722.020 930.380 2725.020 930.390 ;
        RECT 2902.020 930.380 2905.020 930.390 ;
        RECT 2936.000 930.380 2939.000 930.390 ;
        RECT -24.080 927.380 2943.700 930.380 ;
        RECT -19.380 927.370 -16.380 927.380 ;
        RECT 22.020 927.370 25.020 927.380 ;
        RECT 202.020 927.370 205.020 927.380 ;
        RECT 382.020 927.370 385.020 927.380 ;
        RECT 562.020 927.370 565.020 927.380 ;
        RECT 742.020 927.370 745.020 927.380 ;
        RECT 922.020 927.370 925.020 927.380 ;
        RECT 1102.020 927.370 1105.020 927.380 ;
        RECT 1282.020 927.370 1285.020 927.380 ;
        RECT 1462.020 927.370 1465.020 927.380 ;
        RECT 1642.020 927.370 1645.020 927.380 ;
        RECT 1822.020 927.370 1825.020 927.380 ;
        RECT 2002.020 927.370 2005.020 927.380 ;
        RECT 2182.020 927.370 2185.020 927.380 ;
        RECT 2362.020 927.370 2365.020 927.380 ;
        RECT 2542.020 927.370 2545.020 927.380 ;
        RECT 2722.020 927.370 2725.020 927.380 ;
        RECT 2902.020 927.370 2905.020 927.380 ;
        RECT 2936.000 927.370 2939.000 927.380 ;
        RECT -9.980 912.380 -6.980 912.390 ;
        RECT 4.020 912.380 7.020 912.390 ;
        RECT 184.020 912.380 187.020 912.390 ;
        RECT 364.020 912.380 367.020 912.390 ;
        RECT 544.020 912.380 547.020 912.390 ;
        RECT 724.020 912.380 727.020 912.390 ;
        RECT 904.020 912.380 907.020 912.390 ;
        RECT 1084.020 912.380 1087.020 912.390 ;
        RECT 1264.020 912.380 1267.020 912.390 ;
        RECT 1444.020 912.380 1447.020 912.390 ;
        RECT 1624.020 912.380 1627.020 912.390 ;
        RECT 1804.020 912.380 1807.020 912.390 ;
        RECT 1984.020 912.380 1987.020 912.390 ;
        RECT 2164.020 912.380 2167.020 912.390 ;
        RECT 2344.020 912.380 2347.020 912.390 ;
        RECT 2524.020 912.380 2527.020 912.390 ;
        RECT 2704.020 912.380 2707.020 912.390 ;
        RECT 2884.020 912.380 2887.020 912.390 ;
        RECT 2926.600 912.380 2929.600 912.390 ;
        RECT -14.680 909.380 2934.300 912.380 ;
        RECT -9.980 909.370 -6.980 909.380 ;
        RECT 4.020 909.370 7.020 909.380 ;
        RECT 184.020 909.370 187.020 909.380 ;
        RECT 364.020 909.370 367.020 909.380 ;
        RECT 544.020 909.370 547.020 909.380 ;
        RECT 724.020 909.370 727.020 909.380 ;
        RECT 904.020 909.370 907.020 909.380 ;
        RECT 1084.020 909.370 1087.020 909.380 ;
        RECT 1264.020 909.370 1267.020 909.380 ;
        RECT 1444.020 909.370 1447.020 909.380 ;
        RECT 1624.020 909.370 1627.020 909.380 ;
        RECT 1804.020 909.370 1807.020 909.380 ;
        RECT 1984.020 909.370 1987.020 909.380 ;
        RECT 2164.020 909.370 2167.020 909.380 ;
        RECT 2344.020 909.370 2347.020 909.380 ;
        RECT 2524.020 909.370 2527.020 909.380 ;
        RECT 2704.020 909.370 2707.020 909.380 ;
        RECT 2884.020 909.370 2887.020 909.380 ;
        RECT 2926.600 909.370 2929.600 909.380 ;
        RECT -38.180 786.380 -35.180 786.390 ;
        RECT 58.020 786.380 61.020 786.390 ;
        RECT 238.020 786.380 241.020 786.390 ;
        RECT 418.020 786.380 421.020 786.390 ;
        RECT 598.020 786.380 601.020 786.390 ;
        RECT 778.020 786.380 781.020 786.390 ;
        RECT 958.020 786.380 961.020 786.390 ;
        RECT 1138.020 786.380 1141.020 786.390 ;
        RECT 1318.020 786.380 1321.020 786.390 ;
        RECT 1498.020 786.380 1501.020 786.390 ;
        RECT 1678.020 786.380 1681.020 786.390 ;
        RECT 1858.020 786.380 1861.020 786.390 ;
        RECT 2038.020 786.380 2041.020 786.390 ;
        RECT 2218.020 786.380 2221.020 786.390 ;
        RECT 2398.020 786.380 2401.020 786.390 ;
        RECT 2578.020 786.380 2581.020 786.390 ;
        RECT 2758.020 786.380 2761.020 786.390 ;
        RECT 2954.800 786.380 2957.800 786.390 ;
        RECT -42.880 783.380 2962.500 786.380 ;
        RECT -38.180 783.370 -35.180 783.380 ;
        RECT 58.020 783.370 61.020 783.380 ;
        RECT 238.020 783.370 241.020 783.380 ;
        RECT 418.020 783.370 421.020 783.380 ;
        RECT 598.020 783.370 601.020 783.380 ;
        RECT 778.020 783.370 781.020 783.380 ;
        RECT 958.020 783.370 961.020 783.380 ;
        RECT 1138.020 783.370 1141.020 783.380 ;
        RECT 1318.020 783.370 1321.020 783.380 ;
        RECT 1498.020 783.370 1501.020 783.380 ;
        RECT 1678.020 783.370 1681.020 783.380 ;
        RECT 1858.020 783.370 1861.020 783.380 ;
        RECT 2038.020 783.370 2041.020 783.380 ;
        RECT 2218.020 783.370 2221.020 783.380 ;
        RECT 2398.020 783.370 2401.020 783.380 ;
        RECT 2578.020 783.370 2581.020 783.380 ;
        RECT 2758.020 783.370 2761.020 783.380 ;
        RECT 2954.800 783.370 2957.800 783.380 ;
        RECT -28.780 768.380 -25.780 768.390 ;
        RECT 40.020 768.380 43.020 768.390 ;
        RECT 220.020 768.380 223.020 768.390 ;
        RECT 400.020 768.380 403.020 768.390 ;
        RECT 580.020 768.380 583.020 768.390 ;
        RECT 760.020 768.380 763.020 768.390 ;
        RECT 940.020 768.380 943.020 768.390 ;
        RECT 1120.020 768.380 1123.020 768.390 ;
        RECT 1300.020 768.380 1303.020 768.390 ;
        RECT 1480.020 768.380 1483.020 768.390 ;
        RECT 1660.020 768.380 1663.020 768.390 ;
        RECT 1840.020 768.380 1843.020 768.390 ;
        RECT 2020.020 768.380 2023.020 768.390 ;
        RECT 2200.020 768.380 2203.020 768.390 ;
        RECT 2380.020 768.380 2383.020 768.390 ;
        RECT 2560.020 768.380 2563.020 768.390 ;
        RECT 2740.020 768.380 2743.020 768.390 ;
        RECT 2945.400 768.380 2948.400 768.390 ;
        RECT -33.480 765.380 2953.100 768.380 ;
        RECT -28.780 765.370 -25.780 765.380 ;
        RECT 40.020 765.370 43.020 765.380 ;
        RECT 220.020 765.370 223.020 765.380 ;
        RECT 400.020 765.370 403.020 765.380 ;
        RECT 580.020 765.370 583.020 765.380 ;
        RECT 760.020 765.370 763.020 765.380 ;
        RECT 940.020 765.370 943.020 765.380 ;
        RECT 1120.020 765.370 1123.020 765.380 ;
        RECT 1300.020 765.370 1303.020 765.380 ;
        RECT 1480.020 765.370 1483.020 765.380 ;
        RECT 1660.020 765.370 1663.020 765.380 ;
        RECT 1840.020 765.370 1843.020 765.380 ;
        RECT 2020.020 765.370 2023.020 765.380 ;
        RECT 2200.020 765.370 2203.020 765.380 ;
        RECT 2380.020 765.370 2383.020 765.380 ;
        RECT 2560.020 765.370 2563.020 765.380 ;
        RECT 2740.020 765.370 2743.020 765.380 ;
        RECT 2945.400 765.370 2948.400 765.380 ;
        RECT -19.380 750.380 -16.380 750.390 ;
        RECT 22.020 750.380 25.020 750.390 ;
        RECT 202.020 750.380 205.020 750.390 ;
        RECT 382.020 750.380 385.020 750.390 ;
        RECT 562.020 750.380 565.020 750.390 ;
        RECT 742.020 750.380 745.020 750.390 ;
        RECT 922.020 750.380 925.020 750.390 ;
        RECT 1102.020 750.380 1105.020 750.390 ;
        RECT 1282.020 750.380 1285.020 750.390 ;
        RECT 1462.020 750.380 1465.020 750.390 ;
        RECT 1642.020 750.380 1645.020 750.390 ;
        RECT 1822.020 750.380 1825.020 750.390 ;
        RECT 2002.020 750.380 2005.020 750.390 ;
        RECT 2182.020 750.380 2185.020 750.390 ;
        RECT 2362.020 750.380 2365.020 750.390 ;
        RECT 2542.020 750.380 2545.020 750.390 ;
        RECT 2722.020 750.380 2725.020 750.390 ;
        RECT 2902.020 750.380 2905.020 750.390 ;
        RECT 2936.000 750.380 2939.000 750.390 ;
        RECT -24.080 747.380 2943.700 750.380 ;
        RECT -19.380 747.370 -16.380 747.380 ;
        RECT 22.020 747.370 25.020 747.380 ;
        RECT 202.020 747.370 205.020 747.380 ;
        RECT 382.020 747.370 385.020 747.380 ;
        RECT 562.020 747.370 565.020 747.380 ;
        RECT 742.020 747.370 745.020 747.380 ;
        RECT 922.020 747.370 925.020 747.380 ;
        RECT 1102.020 747.370 1105.020 747.380 ;
        RECT 1282.020 747.370 1285.020 747.380 ;
        RECT 1462.020 747.370 1465.020 747.380 ;
        RECT 1642.020 747.370 1645.020 747.380 ;
        RECT 1822.020 747.370 1825.020 747.380 ;
        RECT 2002.020 747.370 2005.020 747.380 ;
        RECT 2182.020 747.370 2185.020 747.380 ;
        RECT 2362.020 747.370 2365.020 747.380 ;
        RECT 2542.020 747.370 2545.020 747.380 ;
        RECT 2722.020 747.370 2725.020 747.380 ;
        RECT 2902.020 747.370 2905.020 747.380 ;
        RECT 2936.000 747.370 2939.000 747.380 ;
        RECT -9.980 732.380 -6.980 732.390 ;
        RECT 4.020 732.380 7.020 732.390 ;
        RECT 184.020 732.380 187.020 732.390 ;
        RECT 364.020 732.380 367.020 732.390 ;
        RECT 544.020 732.380 547.020 732.390 ;
        RECT 724.020 732.380 727.020 732.390 ;
        RECT 904.020 732.380 907.020 732.390 ;
        RECT 1084.020 732.380 1087.020 732.390 ;
        RECT 1264.020 732.380 1267.020 732.390 ;
        RECT 1444.020 732.380 1447.020 732.390 ;
        RECT 1624.020 732.380 1627.020 732.390 ;
        RECT 1804.020 732.380 1807.020 732.390 ;
        RECT 1984.020 732.380 1987.020 732.390 ;
        RECT 2164.020 732.380 2167.020 732.390 ;
        RECT 2344.020 732.380 2347.020 732.390 ;
        RECT 2524.020 732.380 2527.020 732.390 ;
        RECT 2704.020 732.380 2707.020 732.390 ;
        RECT 2884.020 732.380 2887.020 732.390 ;
        RECT 2926.600 732.380 2929.600 732.390 ;
        RECT -14.680 729.380 2934.300 732.380 ;
        RECT -9.980 729.370 -6.980 729.380 ;
        RECT 4.020 729.370 7.020 729.380 ;
        RECT 184.020 729.370 187.020 729.380 ;
        RECT 364.020 729.370 367.020 729.380 ;
        RECT 544.020 729.370 547.020 729.380 ;
        RECT 724.020 729.370 727.020 729.380 ;
        RECT 904.020 729.370 907.020 729.380 ;
        RECT 1084.020 729.370 1087.020 729.380 ;
        RECT 1264.020 729.370 1267.020 729.380 ;
        RECT 1444.020 729.370 1447.020 729.380 ;
        RECT 1624.020 729.370 1627.020 729.380 ;
        RECT 1804.020 729.370 1807.020 729.380 ;
        RECT 1984.020 729.370 1987.020 729.380 ;
        RECT 2164.020 729.370 2167.020 729.380 ;
        RECT 2344.020 729.370 2347.020 729.380 ;
        RECT 2524.020 729.370 2527.020 729.380 ;
        RECT 2704.020 729.370 2707.020 729.380 ;
        RECT 2884.020 729.370 2887.020 729.380 ;
        RECT 2926.600 729.370 2929.600 729.380 ;
        RECT -38.180 606.380 -35.180 606.390 ;
        RECT 58.020 606.380 61.020 606.390 ;
        RECT 238.020 606.380 241.020 606.390 ;
        RECT 418.020 606.380 421.020 606.390 ;
        RECT 598.020 606.380 601.020 606.390 ;
        RECT 778.020 606.380 781.020 606.390 ;
        RECT 958.020 606.380 961.020 606.390 ;
        RECT 1138.020 606.380 1141.020 606.390 ;
        RECT 1318.020 606.380 1321.020 606.390 ;
        RECT 1498.020 606.380 1501.020 606.390 ;
        RECT 1678.020 606.380 1681.020 606.390 ;
        RECT 1858.020 606.380 1861.020 606.390 ;
        RECT 2038.020 606.380 2041.020 606.390 ;
        RECT 2218.020 606.380 2221.020 606.390 ;
        RECT 2398.020 606.380 2401.020 606.390 ;
        RECT 2578.020 606.380 2581.020 606.390 ;
        RECT 2758.020 606.380 2761.020 606.390 ;
        RECT 2954.800 606.380 2957.800 606.390 ;
        RECT -42.880 603.380 2962.500 606.380 ;
        RECT -38.180 603.370 -35.180 603.380 ;
        RECT 58.020 603.370 61.020 603.380 ;
        RECT 238.020 603.370 241.020 603.380 ;
        RECT 418.020 603.370 421.020 603.380 ;
        RECT 598.020 603.370 601.020 603.380 ;
        RECT 778.020 603.370 781.020 603.380 ;
        RECT 958.020 603.370 961.020 603.380 ;
        RECT 1138.020 603.370 1141.020 603.380 ;
        RECT 1318.020 603.370 1321.020 603.380 ;
        RECT 1498.020 603.370 1501.020 603.380 ;
        RECT 1678.020 603.370 1681.020 603.380 ;
        RECT 1858.020 603.370 1861.020 603.380 ;
        RECT 2038.020 603.370 2041.020 603.380 ;
        RECT 2218.020 603.370 2221.020 603.380 ;
        RECT 2398.020 603.370 2401.020 603.380 ;
        RECT 2578.020 603.370 2581.020 603.380 ;
        RECT 2758.020 603.370 2761.020 603.380 ;
        RECT 2954.800 603.370 2957.800 603.380 ;
        RECT -28.780 588.380 -25.780 588.390 ;
        RECT 40.020 588.380 43.020 588.390 ;
        RECT 220.020 588.380 223.020 588.390 ;
        RECT 400.020 588.380 403.020 588.390 ;
        RECT 580.020 588.380 583.020 588.390 ;
        RECT 760.020 588.380 763.020 588.390 ;
        RECT 940.020 588.380 943.020 588.390 ;
        RECT 1120.020 588.380 1123.020 588.390 ;
        RECT 1300.020 588.380 1303.020 588.390 ;
        RECT 1480.020 588.380 1483.020 588.390 ;
        RECT 1660.020 588.380 1663.020 588.390 ;
        RECT 1840.020 588.380 1843.020 588.390 ;
        RECT 2020.020 588.380 2023.020 588.390 ;
        RECT 2200.020 588.380 2203.020 588.390 ;
        RECT 2380.020 588.380 2383.020 588.390 ;
        RECT 2560.020 588.380 2563.020 588.390 ;
        RECT 2740.020 588.380 2743.020 588.390 ;
        RECT 2945.400 588.380 2948.400 588.390 ;
        RECT -33.480 585.380 2953.100 588.380 ;
        RECT -28.780 585.370 -25.780 585.380 ;
        RECT 40.020 585.370 43.020 585.380 ;
        RECT 220.020 585.370 223.020 585.380 ;
        RECT 400.020 585.370 403.020 585.380 ;
        RECT 580.020 585.370 583.020 585.380 ;
        RECT 760.020 585.370 763.020 585.380 ;
        RECT 940.020 585.370 943.020 585.380 ;
        RECT 1120.020 585.370 1123.020 585.380 ;
        RECT 1300.020 585.370 1303.020 585.380 ;
        RECT 1480.020 585.370 1483.020 585.380 ;
        RECT 1660.020 585.370 1663.020 585.380 ;
        RECT 1840.020 585.370 1843.020 585.380 ;
        RECT 2020.020 585.370 2023.020 585.380 ;
        RECT 2200.020 585.370 2203.020 585.380 ;
        RECT 2380.020 585.370 2383.020 585.380 ;
        RECT 2560.020 585.370 2563.020 585.380 ;
        RECT 2740.020 585.370 2743.020 585.380 ;
        RECT 2945.400 585.370 2948.400 585.380 ;
        RECT -19.380 570.380 -16.380 570.390 ;
        RECT 22.020 570.380 25.020 570.390 ;
        RECT 202.020 570.380 205.020 570.390 ;
        RECT 382.020 570.380 385.020 570.390 ;
        RECT 562.020 570.380 565.020 570.390 ;
        RECT 742.020 570.380 745.020 570.390 ;
        RECT 922.020 570.380 925.020 570.390 ;
        RECT 1102.020 570.380 1105.020 570.390 ;
        RECT 1282.020 570.380 1285.020 570.390 ;
        RECT 1462.020 570.380 1465.020 570.390 ;
        RECT 1642.020 570.380 1645.020 570.390 ;
        RECT 1822.020 570.380 1825.020 570.390 ;
        RECT 2002.020 570.380 2005.020 570.390 ;
        RECT 2182.020 570.380 2185.020 570.390 ;
        RECT 2362.020 570.380 2365.020 570.390 ;
        RECT 2542.020 570.380 2545.020 570.390 ;
        RECT 2722.020 570.380 2725.020 570.390 ;
        RECT 2902.020 570.380 2905.020 570.390 ;
        RECT 2936.000 570.380 2939.000 570.390 ;
        RECT -24.080 567.380 2943.700 570.380 ;
        RECT -19.380 567.370 -16.380 567.380 ;
        RECT 22.020 567.370 25.020 567.380 ;
        RECT 202.020 567.370 205.020 567.380 ;
        RECT 382.020 567.370 385.020 567.380 ;
        RECT 562.020 567.370 565.020 567.380 ;
        RECT 742.020 567.370 745.020 567.380 ;
        RECT 922.020 567.370 925.020 567.380 ;
        RECT 1102.020 567.370 1105.020 567.380 ;
        RECT 1282.020 567.370 1285.020 567.380 ;
        RECT 1462.020 567.370 1465.020 567.380 ;
        RECT 1642.020 567.370 1645.020 567.380 ;
        RECT 1822.020 567.370 1825.020 567.380 ;
        RECT 2002.020 567.370 2005.020 567.380 ;
        RECT 2182.020 567.370 2185.020 567.380 ;
        RECT 2362.020 567.370 2365.020 567.380 ;
        RECT 2542.020 567.370 2545.020 567.380 ;
        RECT 2722.020 567.370 2725.020 567.380 ;
        RECT 2902.020 567.370 2905.020 567.380 ;
        RECT 2936.000 567.370 2939.000 567.380 ;
        RECT -9.980 552.380 -6.980 552.390 ;
        RECT 4.020 552.380 7.020 552.390 ;
        RECT 184.020 552.380 187.020 552.390 ;
        RECT 364.020 552.380 367.020 552.390 ;
        RECT 544.020 552.380 547.020 552.390 ;
        RECT 724.020 552.380 727.020 552.390 ;
        RECT 904.020 552.380 907.020 552.390 ;
        RECT 1084.020 552.380 1087.020 552.390 ;
        RECT 1264.020 552.380 1267.020 552.390 ;
        RECT 1444.020 552.380 1447.020 552.390 ;
        RECT 1624.020 552.380 1627.020 552.390 ;
        RECT 1804.020 552.380 1807.020 552.390 ;
        RECT 1984.020 552.380 1987.020 552.390 ;
        RECT 2164.020 552.380 2167.020 552.390 ;
        RECT 2344.020 552.380 2347.020 552.390 ;
        RECT 2524.020 552.380 2527.020 552.390 ;
        RECT 2704.020 552.380 2707.020 552.390 ;
        RECT 2884.020 552.380 2887.020 552.390 ;
        RECT 2926.600 552.380 2929.600 552.390 ;
        RECT -14.680 549.380 2934.300 552.380 ;
        RECT -9.980 549.370 -6.980 549.380 ;
        RECT 4.020 549.370 7.020 549.380 ;
        RECT 184.020 549.370 187.020 549.380 ;
        RECT 364.020 549.370 367.020 549.380 ;
        RECT 544.020 549.370 547.020 549.380 ;
        RECT 724.020 549.370 727.020 549.380 ;
        RECT 904.020 549.370 907.020 549.380 ;
        RECT 1084.020 549.370 1087.020 549.380 ;
        RECT 1264.020 549.370 1267.020 549.380 ;
        RECT 1444.020 549.370 1447.020 549.380 ;
        RECT 1624.020 549.370 1627.020 549.380 ;
        RECT 1804.020 549.370 1807.020 549.380 ;
        RECT 1984.020 549.370 1987.020 549.380 ;
        RECT 2164.020 549.370 2167.020 549.380 ;
        RECT 2344.020 549.370 2347.020 549.380 ;
        RECT 2524.020 549.370 2527.020 549.380 ;
        RECT 2704.020 549.370 2707.020 549.380 ;
        RECT 2884.020 549.370 2887.020 549.380 ;
        RECT 2926.600 549.370 2929.600 549.380 ;
        RECT -38.180 426.380 -35.180 426.390 ;
        RECT 58.020 426.380 61.020 426.390 ;
        RECT 238.020 426.380 241.020 426.390 ;
        RECT 418.020 426.380 421.020 426.390 ;
        RECT 598.020 426.380 601.020 426.390 ;
        RECT 778.020 426.380 781.020 426.390 ;
        RECT 958.020 426.380 961.020 426.390 ;
        RECT 1138.020 426.380 1141.020 426.390 ;
        RECT 1318.020 426.380 1321.020 426.390 ;
        RECT 1498.020 426.380 1501.020 426.390 ;
        RECT 1678.020 426.380 1681.020 426.390 ;
        RECT 1858.020 426.380 1861.020 426.390 ;
        RECT 2038.020 426.380 2041.020 426.390 ;
        RECT 2218.020 426.380 2221.020 426.390 ;
        RECT 2398.020 426.380 2401.020 426.390 ;
        RECT 2578.020 426.380 2581.020 426.390 ;
        RECT 2758.020 426.380 2761.020 426.390 ;
        RECT 2954.800 426.380 2957.800 426.390 ;
        RECT -42.880 423.380 2962.500 426.380 ;
        RECT -38.180 423.370 -35.180 423.380 ;
        RECT 58.020 423.370 61.020 423.380 ;
        RECT 238.020 423.370 241.020 423.380 ;
        RECT 418.020 423.370 421.020 423.380 ;
        RECT 598.020 423.370 601.020 423.380 ;
        RECT 778.020 423.370 781.020 423.380 ;
        RECT 958.020 423.370 961.020 423.380 ;
        RECT 1138.020 423.370 1141.020 423.380 ;
        RECT 1318.020 423.370 1321.020 423.380 ;
        RECT 1498.020 423.370 1501.020 423.380 ;
        RECT 1678.020 423.370 1681.020 423.380 ;
        RECT 1858.020 423.370 1861.020 423.380 ;
        RECT 2038.020 423.370 2041.020 423.380 ;
        RECT 2218.020 423.370 2221.020 423.380 ;
        RECT 2398.020 423.370 2401.020 423.380 ;
        RECT 2578.020 423.370 2581.020 423.380 ;
        RECT 2758.020 423.370 2761.020 423.380 ;
        RECT 2954.800 423.370 2957.800 423.380 ;
        RECT -28.780 408.380 -25.780 408.390 ;
        RECT 40.020 408.380 43.020 408.390 ;
        RECT 220.020 408.380 223.020 408.390 ;
        RECT 400.020 408.380 403.020 408.390 ;
        RECT 580.020 408.380 583.020 408.390 ;
        RECT 760.020 408.380 763.020 408.390 ;
        RECT 940.020 408.380 943.020 408.390 ;
        RECT 1120.020 408.380 1123.020 408.390 ;
        RECT 1300.020 408.380 1303.020 408.390 ;
        RECT 1480.020 408.380 1483.020 408.390 ;
        RECT 1660.020 408.380 1663.020 408.390 ;
        RECT 1840.020 408.380 1843.020 408.390 ;
        RECT 2020.020 408.380 2023.020 408.390 ;
        RECT 2200.020 408.380 2203.020 408.390 ;
        RECT 2380.020 408.380 2383.020 408.390 ;
        RECT 2560.020 408.380 2563.020 408.390 ;
        RECT 2740.020 408.380 2743.020 408.390 ;
        RECT 2945.400 408.380 2948.400 408.390 ;
        RECT -33.480 405.380 2953.100 408.380 ;
        RECT -28.780 405.370 -25.780 405.380 ;
        RECT 40.020 405.370 43.020 405.380 ;
        RECT 220.020 405.370 223.020 405.380 ;
        RECT 400.020 405.370 403.020 405.380 ;
        RECT 580.020 405.370 583.020 405.380 ;
        RECT 760.020 405.370 763.020 405.380 ;
        RECT 940.020 405.370 943.020 405.380 ;
        RECT 1120.020 405.370 1123.020 405.380 ;
        RECT 1300.020 405.370 1303.020 405.380 ;
        RECT 1480.020 405.370 1483.020 405.380 ;
        RECT 1660.020 405.370 1663.020 405.380 ;
        RECT 1840.020 405.370 1843.020 405.380 ;
        RECT 2020.020 405.370 2023.020 405.380 ;
        RECT 2200.020 405.370 2203.020 405.380 ;
        RECT 2380.020 405.370 2383.020 405.380 ;
        RECT 2560.020 405.370 2563.020 405.380 ;
        RECT 2740.020 405.370 2743.020 405.380 ;
        RECT 2945.400 405.370 2948.400 405.380 ;
        RECT -19.380 390.380 -16.380 390.390 ;
        RECT 22.020 390.380 25.020 390.390 ;
        RECT 202.020 390.380 205.020 390.390 ;
        RECT 382.020 390.380 385.020 390.390 ;
        RECT 562.020 390.380 565.020 390.390 ;
        RECT 742.020 390.380 745.020 390.390 ;
        RECT 922.020 390.380 925.020 390.390 ;
        RECT 1102.020 390.380 1105.020 390.390 ;
        RECT 1282.020 390.380 1285.020 390.390 ;
        RECT 1462.020 390.380 1465.020 390.390 ;
        RECT 1642.020 390.380 1645.020 390.390 ;
        RECT 1822.020 390.380 1825.020 390.390 ;
        RECT 2002.020 390.380 2005.020 390.390 ;
        RECT 2182.020 390.380 2185.020 390.390 ;
        RECT 2362.020 390.380 2365.020 390.390 ;
        RECT 2542.020 390.380 2545.020 390.390 ;
        RECT 2722.020 390.380 2725.020 390.390 ;
        RECT 2902.020 390.380 2905.020 390.390 ;
        RECT 2936.000 390.380 2939.000 390.390 ;
        RECT -24.080 387.380 2943.700 390.380 ;
        RECT -19.380 387.370 -16.380 387.380 ;
        RECT 22.020 387.370 25.020 387.380 ;
        RECT 202.020 387.370 205.020 387.380 ;
        RECT 382.020 387.370 385.020 387.380 ;
        RECT 562.020 387.370 565.020 387.380 ;
        RECT 742.020 387.370 745.020 387.380 ;
        RECT 922.020 387.370 925.020 387.380 ;
        RECT 1102.020 387.370 1105.020 387.380 ;
        RECT 1282.020 387.370 1285.020 387.380 ;
        RECT 1462.020 387.370 1465.020 387.380 ;
        RECT 1642.020 387.370 1645.020 387.380 ;
        RECT 1822.020 387.370 1825.020 387.380 ;
        RECT 2002.020 387.370 2005.020 387.380 ;
        RECT 2182.020 387.370 2185.020 387.380 ;
        RECT 2362.020 387.370 2365.020 387.380 ;
        RECT 2542.020 387.370 2545.020 387.380 ;
        RECT 2722.020 387.370 2725.020 387.380 ;
        RECT 2902.020 387.370 2905.020 387.380 ;
        RECT 2936.000 387.370 2939.000 387.380 ;
        RECT -9.980 372.380 -6.980 372.390 ;
        RECT 4.020 372.380 7.020 372.390 ;
        RECT 184.020 372.380 187.020 372.390 ;
        RECT 364.020 372.380 367.020 372.390 ;
        RECT 544.020 372.380 547.020 372.390 ;
        RECT 724.020 372.380 727.020 372.390 ;
        RECT 904.020 372.380 907.020 372.390 ;
        RECT 1084.020 372.380 1087.020 372.390 ;
        RECT 1264.020 372.380 1267.020 372.390 ;
        RECT 1444.020 372.380 1447.020 372.390 ;
        RECT 1624.020 372.380 1627.020 372.390 ;
        RECT 1804.020 372.380 1807.020 372.390 ;
        RECT 1984.020 372.380 1987.020 372.390 ;
        RECT 2164.020 372.380 2167.020 372.390 ;
        RECT 2344.020 372.380 2347.020 372.390 ;
        RECT 2524.020 372.380 2527.020 372.390 ;
        RECT 2704.020 372.380 2707.020 372.390 ;
        RECT 2884.020 372.380 2887.020 372.390 ;
        RECT 2926.600 372.380 2929.600 372.390 ;
        RECT -14.680 369.380 2934.300 372.380 ;
        RECT -9.980 369.370 -6.980 369.380 ;
        RECT 4.020 369.370 7.020 369.380 ;
        RECT 184.020 369.370 187.020 369.380 ;
        RECT 364.020 369.370 367.020 369.380 ;
        RECT 544.020 369.370 547.020 369.380 ;
        RECT 724.020 369.370 727.020 369.380 ;
        RECT 904.020 369.370 907.020 369.380 ;
        RECT 1084.020 369.370 1087.020 369.380 ;
        RECT 1264.020 369.370 1267.020 369.380 ;
        RECT 1444.020 369.370 1447.020 369.380 ;
        RECT 1624.020 369.370 1627.020 369.380 ;
        RECT 1804.020 369.370 1807.020 369.380 ;
        RECT 1984.020 369.370 1987.020 369.380 ;
        RECT 2164.020 369.370 2167.020 369.380 ;
        RECT 2344.020 369.370 2347.020 369.380 ;
        RECT 2524.020 369.370 2527.020 369.380 ;
        RECT 2704.020 369.370 2707.020 369.380 ;
        RECT 2884.020 369.370 2887.020 369.380 ;
        RECT 2926.600 369.370 2929.600 369.380 ;
        RECT -38.180 246.380 -35.180 246.390 ;
        RECT 58.020 246.380 61.020 246.390 ;
        RECT 238.020 246.380 241.020 246.390 ;
        RECT 418.020 246.380 421.020 246.390 ;
        RECT 598.020 246.380 601.020 246.390 ;
        RECT 778.020 246.380 781.020 246.390 ;
        RECT 958.020 246.380 961.020 246.390 ;
        RECT 1138.020 246.380 1141.020 246.390 ;
        RECT 1318.020 246.380 1321.020 246.390 ;
        RECT 1498.020 246.380 1501.020 246.390 ;
        RECT 1678.020 246.380 1681.020 246.390 ;
        RECT 1858.020 246.380 1861.020 246.390 ;
        RECT 2038.020 246.380 2041.020 246.390 ;
        RECT 2218.020 246.380 2221.020 246.390 ;
        RECT 2398.020 246.380 2401.020 246.390 ;
        RECT 2578.020 246.380 2581.020 246.390 ;
        RECT 2758.020 246.380 2761.020 246.390 ;
        RECT 2954.800 246.380 2957.800 246.390 ;
        RECT -42.880 243.380 2962.500 246.380 ;
        RECT -38.180 243.370 -35.180 243.380 ;
        RECT 58.020 243.370 61.020 243.380 ;
        RECT 238.020 243.370 241.020 243.380 ;
        RECT 418.020 243.370 421.020 243.380 ;
        RECT 598.020 243.370 601.020 243.380 ;
        RECT 778.020 243.370 781.020 243.380 ;
        RECT 958.020 243.370 961.020 243.380 ;
        RECT 1138.020 243.370 1141.020 243.380 ;
        RECT 1318.020 243.370 1321.020 243.380 ;
        RECT 1498.020 243.370 1501.020 243.380 ;
        RECT 1678.020 243.370 1681.020 243.380 ;
        RECT 1858.020 243.370 1861.020 243.380 ;
        RECT 2038.020 243.370 2041.020 243.380 ;
        RECT 2218.020 243.370 2221.020 243.380 ;
        RECT 2398.020 243.370 2401.020 243.380 ;
        RECT 2578.020 243.370 2581.020 243.380 ;
        RECT 2758.020 243.370 2761.020 243.380 ;
        RECT 2954.800 243.370 2957.800 243.380 ;
        RECT -28.780 228.380 -25.780 228.390 ;
        RECT 40.020 228.380 43.020 228.390 ;
        RECT 220.020 228.380 223.020 228.390 ;
        RECT 400.020 228.380 403.020 228.390 ;
        RECT 580.020 228.380 583.020 228.390 ;
        RECT 760.020 228.380 763.020 228.390 ;
        RECT 940.020 228.380 943.020 228.390 ;
        RECT 1120.020 228.380 1123.020 228.390 ;
        RECT 1300.020 228.380 1303.020 228.390 ;
        RECT 1480.020 228.380 1483.020 228.390 ;
        RECT 1660.020 228.380 1663.020 228.390 ;
        RECT 1840.020 228.380 1843.020 228.390 ;
        RECT 2020.020 228.380 2023.020 228.390 ;
        RECT 2200.020 228.380 2203.020 228.390 ;
        RECT 2380.020 228.380 2383.020 228.390 ;
        RECT 2560.020 228.380 2563.020 228.390 ;
        RECT 2740.020 228.380 2743.020 228.390 ;
        RECT 2945.400 228.380 2948.400 228.390 ;
        RECT -33.480 225.380 2953.100 228.380 ;
        RECT -28.780 225.370 -25.780 225.380 ;
        RECT 40.020 225.370 43.020 225.380 ;
        RECT 220.020 225.370 223.020 225.380 ;
        RECT 400.020 225.370 403.020 225.380 ;
        RECT 580.020 225.370 583.020 225.380 ;
        RECT 760.020 225.370 763.020 225.380 ;
        RECT 940.020 225.370 943.020 225.380 ;
        RECT 1120.020 225.370 1123.020 225.380 ;
        RECT 1300.020 225.370 1303.020 225.380 ;
        RECT 1480.020 225.370 1483.020 225.380 ;
        RECT 1660.020 225.370 1663.020 225.380 ;
        RECT 1840.020 225.370 1843.020 225.380 ;
        RECT 2020.020 225.370 2023.020 225.380 ;
        RECT 2200.020 225.370 2203.020 225.380 ;
        RECT 2380.020 225.370 2383.020 225.380 ;
        RECT 2560.020 225.370 2563.020 225.380 ;
        RECT 2740.020 225.370 2743.020 225.380 ;
        RECT 2945.400 225.370 2948.400 225.380 ;
        RECT -19.380 210.380 -16.380 210.390 ;
        RECT 22.020 210.380 25.020 210.390 ;
        RECT 202.020 210.380 205.020 210.390 ;
        RECT 382.020 210.380 385.020 210.390 ;
        RECT 562.020 210.380 565.020 210.390 ;
        RECT 742.020 210.380 745.020 210.390 ;
        RECT 922.020 210.380 925.020 210.390 ;
        RECT 1102.020 210.380 1105.020 210.390 ;
        RECT 1282.020 210.380 1285.020 210.390 ;
        RECT 1462.020 210.380 1465.020 210.390 ;
        RECT 1642.020 210.380 1645.020 210.390 ;
        RECT 1822.020 210.380 1825.020 210.390 ;
        RECT 2002.020 210.380 2005.020 210.390 ;
        RECT 2182.020 210.380 2185.020 210.390 ;
        RECT 2362.020 210.380 2365.020 210.390 ;
        RECT 2542.020 210.380 2545.020 210.390 ;
        RECT 2722.020 210.380 2725.020 210.390 ;
        RECT 2902.020 210.380 2905.020 210.390 ;
        RECT 2936.000 210.380 2939.000 210.390 ;
        RECT -24.080 207.380 2943.700 210.380 ;
        RECT -19.380 207.370 -16.380 207.380 ;
        RECT 22.020 207.370 25.020 207.380 ;
        RECT 202.020 207.370 205.020 207.380 ;
        RECT 382.020 207.370 385.020 207.380 ;
        RECT 562.020 207.370 565.020 207.380 ;
        RECT 742.020 207.370 745.020 207.380 ;
        RECT 922.020 207.370 925.020 207.380 ;
        RECT 1102.020 207.370 1105.020 207.380 ;
        RECT 1282.020 207.370 1285.020 207.380 ;
        RECT 1462.020 207.370 1465.020 207.380 ;
        RECT 1642.020 207.370 1645.020 207.380 ;
        RECT 1822.020 207.370 1825.020 207.380 ;
        RECT 2002.020 207.370 2005.020 207.380 ;
        RECT 2182.020 207.370 2185.020 207.380 ;
        RECT 2362.020 207.370 2365.020 207.380 ;
        RECT 2542.020 207.370 2545.020 207.380 ;
        RECT 2722.020 207.370 2725.020 207.380 ;
        RECT 2902.020 207.370 2905.020 207.380 ;
        RECT 2936.000 207.370 2939.000 207.380 ;
        RECT -9.980 192.380 -6.980 192.390 ;
        RECT 4.020 192.380 7.020 192.390 ;
        RECT 184.020 192.380 187.020 192.390 ;
        RECT 364.020 192.380 367.020 192.390 ;
        RECT 544.020 192.380 547.020 192.390 ;
        RECT 724.020 192.380 727.020 192.390 ;
        RECT 904.020 192.380 907.020 192.390 ;
        RECT 1084.020 192.380 1087.020 192.390 ;
        RECT 1264.020 192.380 1267.020 192.390 ;
        RECT 1444.020 192.380 1447.020 192.390 ;
        RECT 1624.020 192.380 1627.020 192.390 ;
        RECT 1804.020 192.380 1807.020 192.390 ;
        RECT 1984.020 192.380 1987.020 192.390 ;
        RECT 2164.020 192.380 2167.020 192.390 ;
        RECT 2344.020 192.380 2347.020 192.390 ;
        RECT 2524.020 192.380 2527.020 192.390 ;
        RECT 2704.020 192.380 2707.020 192.390 ;
        RECT 2884.020 192.380 2887.020 192.390 ;
        RECT 2926.600 192.380 2929.600 192.390 ;
        RECT -14.680 189.380 2934.300 192.380 ;
        RECT -9.980 189.370 -6.980 189.380 ;
        RECT 4.020 189.370 7.020 189.380 ;
        RECT 184.020 189.370 187.020 189.380 ;
        RECT 364.020 189.370 367.020 189.380 ;
        RECT 544.020 189.370 547.020 189.380 ;
        RECT 724.020 189.370 727.020 189.380 ;
        RECT 904.020 189.370 907.020 189.380 ;
        RECT 1084.020 189.370 1087.020 189.380 ;
        RECT 1264.020 189.370 1267.020 189.380 ;
        RECT 1444.020 189.370 1447.020 189.380 ;
        RECT 1624.020 189.370 1627.020 189.380 ;
        RECT 1804.020 189.370 1807.020 189.380 ;
        RECT 1984.020 189.370 1987.020 189.380 ;
        RECT 2164.020 189.370 2167.020 189.380 ;
        RECT 2344.020 189.370 2347.020 189.380 ;
        RECT 2524.020 189.370 2527.020 189.380 ;
        RECT 2704.020 189.370 2707.020 189.380 ;
        RECT 2884.020 189.370 2887.020 189.380 ;
        RECT 2926.600 189.370 2929.600 189.380 ;
        RECT -38.180 66.380 -35.180 66.390 ;
        RECT 58.020 66.380 61.020 66.390 ;
        RECT 238.020 66.380 241.020 66.390 ;
        RECT 418.020 66.380 421.020 66.390 ;
        RECT 598.020 66.380 601.020 66.390 ;
        RECT 778.020 66.380 781.020 66.390 ;
        RECT 958.020 66.380 961.020 66.390 ;
        RECT 1138.020 66.380 1141.020 66.390 ;
        RECT 1318.020 66.380 1321.020 66.390 ;
        RECT 1498.020 66.380 1501.020 66.390 ;
        RECT 1678.020 66.380 1681.020 66.390 ;
        RECT 1858.020 66.380 1861.020 66.390 ;
        RECT 2038.020 66.380 2041.020 66.390 ;
        RECT 2218.020 66.380 2221.020 66.390 ;
        RECT 2398.020 66.380 2401.020 66.390 ;
        RECT 2578.020 66.380 2581.020 66.390 ;
        RECT 2758.020 66.380 2761.020 66.390 ;
        RECT 2954.800 66.380 2957.800 66.390 ;
        RECT -42.880 63.380 2962.500 66.380 ;
        RECT -38.180 63.370 -35.180 63.380 ;
        RECT 58.020 63.370 61.020 63.380 ;
        RECT 238.020 63.370 241.020 63.380 ;
        RECT 418.020 63.370 421.020 63.380 ;
        RECT 598.020 63.370 601.020 63.380 ;
        RECT 778.020 63.370 781.020 63.380 ;
        RECT 958.020 63.370 961.020 63.380 ;
        RECT 1138.020 63.370 1141.020 63.380 ;
        RECT 1318.020 63.370 1321.020 63.380 ;
        RECT 1498.020 63.370 1501.020 63.380 ;
        RECT 1678.020 63.370 1681.020 63.380 ;
        RECT 1858.020 63.370 1861.020 63.380 ;
        RECT 2038.020 63.370 2041.020 63.380 ;
        RECT 2218.020 63.370 2221.020 63.380 ;
        RECT 2398.020 63.370 2401.020 63.380 ;
        RECT 2578.020 63.370 2581.020 63.380 ;
        RECT 2758.020 63.370 2761.020 63.380 ;
        RECT 2954.800 63.370 2957.800 63.380 ;
        RECT -28.780 48.380 -25.780 48.390 ;
        RECT 40.020 48.380 43.020 48.390 ;
        RECT 220.020 48.380 223.020 48.390 ;
        RECT 400.020 48.380 403.020 48.390 ;
        RECT 580.020 48.380 583.020 48.390 ;
        RECT 760.020 48.380 763.020 48.390 ;
        RECT 940.020 48.380 943.020 48.390 ;
        RECT 1120.020 48.380 1123.020 48.390 ;
        RECT 1300.020 48.380 1303.020 48.390 ;
        RECT 1480.020 48.380 1483.020 48.390 ;
        RECT 1660.020 48.380 1663.020 48.390 ;
        RECT 1840.020 48.380 1843.020 48.390 ;
        RECT 2020.020 48.380 2023.020 48.390 ;
        RECT 2200.020 48.380 2203.020 48.390 ;
        RECT 2380.020 48.380 2383.020 48.390 ;
        RECT 2560.020 48.380 2563.020 48.390 ;
        RECT 2740.020 48.380 2743.020 48.390 ;
        RECT 2945.400 48.380 2948.400 48.390 ;
        RECT -33.480 45.380 2953.100 48.380 ;
        RECT -28.780 45.370 -25.780 45.380 ;
        RECT 40.020 45.370 43.020 45.380 ;
        RECT 220.020 45.370 223.020 45.380 ;
        RECT 400.020 45.370 403.020 45.380 ;
        RECT 580.020 45.370 583.020 45.380 ;
        RECT 760.020 45.370 763.020 45.380 ;
        RECT 940.020 45.370 943.020 45.380 ;
        RECT 1120.020 45.370 1123.020 45.380 ;
        RECT 1300.020 45.370 1303.020 45.380 ;
        RECT 1480.020 45.370 1483.020 45.380 ;
        RECT 1660.020 45.370 1663.020 45.380 ;
        RECT 1840.020 45.370 1843.020 45.380 ;
        RECT 2020.020 45.370 2023.020 45.380 ;
        RECT 2200.020 45.370 2203.020 45.380 ;
        RECT 2380.020 45.370 2383.020 45.380 ;
        RECT 2560.020 45.370 2563.020 45.380 ;
        RECT 2740.020 45.370 2743.020 45.380 ;
        RECT 2945.400 45.370 2948.400 45.380 ;
        RECT -19.380 30.380 -16.380 30.390 ;
        RECT 22.020 30.380 25.020 30.390 ;
        RECT 202.020 30.380 205.020 30.390 ;
        RECT 382.020 30.380 385.020 30.390 ;
        RECT 562.020 30.380 565.020 30.390 ;
        RECT 742.020 30.380 745.020 30.390 ;
        RECT 922.020 30.380 925.020 30.390 ;
        RECT 1102.020 30.380 1105.020 30.390 ;
        RECT 1282.020 30.380 1285.020 30.390 ;
        RECT 1462.020 30.380 1465.020 30.390 ;
        RECT 1642.020 30.380 1645.020 30.390 ;
        RECT 1822.020 30.380 1825.020 30.390 ;
        RECT 2002.020 30.380 2005.020 30.390 ;
        RECT 2182.020 30.380 2185.020 30.390 ;
        RECT 2362.020 30.380 2365.020 30.390 ;
        RECT 2542.020 30.380 2545.020 30.390 ;
        RECT 2722.020 30.380 2725.020 30.390 ;
        RECT 2902.020 30.380 2905.020 30.390 ;
        RECT 2936.000 30.380 2939.000 30.390 ;
        RECT -24.080 27.380 2943.700 30.380 ;
        RECT -19.380 27.370 -16.380 27.380 ;
        RECT 22.020 27.370 25.020 27.380 ;
        RECT 202.020 27.370 205.020 27.380 ;
        RECT 382.020 27.370 385.020 27.380 ;
        RECT 562.020 27.370 565.020 27.380 ;
        RECT 742.020 27.370 745.020 27.380 ;
        RECT 922.020 27.370 925.020 27.380 ;
        RECT 1102.020 27.370 1105.020 27.380 ;
        RECT 1282.020 27.370 1285.020 27.380 ;
        RECT 1462.020 27.370 1465.020 27.380 ;
        RECT 1642.020 27.370 1645.020 27.380 ;
        RECT 1822.020 27.370 1825.020 27.380 ;
        RECT 2002.020 27.370 2005.020 27.380 ;
        RECT 2182.020 27.370 2185.020 27.380 ;
        RECT 2362.020 27.370 2365.020 27.380 ;
        RECT 2542.020 27.370 2545.020 27.380 ;
        RECT 2722.020 27.370 2725.020 27.380 ;
        RECT 2902.020 27.370 2905.020 27.380 ;
        RECT 2936.000 27.370 2939.000 27.380 ;
        RECT -9.980 12.380 -6.980 12.390 ;
        RECT 4.020 12.380 7.020 12.390 ;
        RECT 184.020 12.380 187.020 12.390 ;
        RECT 364.020 12.380 367.020 12.390 ;
        RECT 544.020 12.380 547.020 12.390 ;
        RECT 724.020 12.380 727.020 12.390 ;
        RECT 904.020 12.380 907.020 12.390 ;
        RECT 1084.020 12.380 1087.020 12.390 ;
        RECT 1264.020 12.380 1267.020 12.390 ;
        RECT 1444.020 12.380 1447.020 12.390 ;
        RECT 1624.020 12.380 1627.020 12.390 ;
        RECT 1804.020 12.380 1807.020 12.390 ;
        RECT 1984.020 12.380 1987.020 12.390 ;
        RECT 2164.020 12.380 2167.020 12.390 ;
        RECT 2344.020 12.380 2347.020 12.390 ;
        RECT 2524.020 12.380 2527.020 12.390 ;
        RECT 2704.020 12.380 2707.020 12.390 ;
        RECT 2884.020 12.380 2887.020 12.390 ;
        RECT 2926.600 12.380 2929.600 12.390 ;
        RECT -14.680 9.380 2934.300 12.380 ;
        RECT -9.980 9.370 -6.980 9.380 ;
        RECT 4.020 9.370 7.020 9.380 ;
        RECT 184.020 9.370 187.020 9.380 ;
        RECT 364.020 9.370 367.020 9.380 ;
        RECT 544.020 9.370 547.020 9.380 ;
        RECT 724.020 9.370 727.020 9.380 ;
        RECT 904.020 9.370 907.020 9.380 ;
        RECT 1084.020 9.370 1087.020 9.380 ;
        RECT 1264.020 9.370 1267.020 9.380 ;
        RECT 1444.020 9.370 1447.020 9.380 ;
        RECT 1624.020 9.370 1627.020 9.380 ;
        RECT 1804.020 9.370 1807.020 9.380 ;
        RECT 1984.020 9.370 1987.020 9.380 ;
        RECT 2164.020 9.370 2167.020 9.380 ;
        RECT 2344.020 9.370 2347.020 9.380 ;
        RECT 2524.020 9.370 2527.020 9.380 ;
        RECT 2704.020 9.370 2707.020 9.380 ;
        RECT 2884.020 9.370 2887.020 9.380 ;
        RECT 2926.600 9.370 2929.600 9.380 ;
        RECT -9.980 -1.620 -6.980 -1.610 ;
        RECT 4.020 -1.620 7.020 -1.610 ;
        RECT 184.020 -1.620 187.020 -1.610 ;
        RECT 364.020 -1.620 367.020 -1.610 ;
        RECT 544.020 -1.620 547.020 -1.610 ;
        RECT 724.020 -1.620 727.020 -1.610 ;
        RECT 904.020 -1.620 907.020 -1.610 ;
        RECT 1084.020 -1.620 1087.020 -1.610 ;
        RECT 1264.020 -1.620 1267.020 -1.610 ;
        RECT 1444.020 -1.620 1447.020 -1.610 ;
        RECT 1624.020 -1.620 1627.020 -1.610 ;
        RECT 1804.020 -1.620 1807.020 -1.610 ;
        RECT 1984.020 -1.620 1987.020 -1.610 ;
        RECT 2164.020 -1.620 2167.020 -1.610 ;
        RECT 2344.020 -1.620 2347.020 -1.610 ;
        RECT 2524.020 -1.620 2527.020 -1.610 ;
        RECT 2704.020 -1.620 2707.020 -1.610 ;
        RECT 2884.020 -1.620 2887.020 -1.610 ;
        RECT 2926.600 -1.620 2929.600 -1.610 ;
        RECT -9.980 -4.620 2929.600 -1.620 ;
        RECT -9.980 -4.630 -6.980 -4.620 ;
        RECT 4.020 -4.630 7.020 -4.620 ;
        RECT 184.020 -4.630 187.020 -4.620 ;
        RECT 364.020 -4.630 367.020 -4.620 ;
        RECT 544.020 -4.630 547.020 -4.620 ;
        RECT 724.020 -4.630 727.020 -4.620 ;
        RECT 904.020 -4.630 907.020 -4.620 ;
        RECT 1084.020 -4.630 1087.020 -4.620 ;
        RECT 1264.020 -4.630 1267.020 -4.620 ;
        RECT 1444.020 -4.630 1447.020 -4.620 ;
        RECT 1624.020 -4.630 1627.020 -4.620 ;
        RECT 1804.020 -4.630 1807.020 -4.620 ;
        RECT 1984.020 -4.630 1987.020 -4.620 ;
        RECT 2164.020 -4.630 2167.020 -4.620 ;
        RECT 2344.020 -4.630 2347.020 -4.620 ;
        RECT 2524.020 -4.630 2527.020 -4.620 ;
        RECT 2704.020 -4.630 2707.020 -4.620 ;
        RECT 2884.020 -4.630 2887.020 -4.620 ;
        RECT 2926.600 -4.630 2929.600 -4.620 ;
        RECT -19.380 -11.020 -16.380 -11.010 ;
        RECT 22.020 -11.020 25.020 -11.010 ;
        RECT 202.020 -11.020 205.020 -11.010 ;
        RECT 382.020 -11.020 385.020 -11.010 ;
        RECT 562.020 -11.020 565.020 -11.010 ;
        RECT 742.020 -11.020 745.020 -11.010 ;
        RECT 922.020 -11.020 925.020 -11.010 ;
        RECT 1102.020 -11.020 1105.020 -11.010 ;
        RECT 1282.020 -11.020 1285.020 -11.010 ;
        RECT 1462.020 -11.020 1465.020 -11.010 ;
        RECT 1642.020 -11.020 1645.020 -11.010 ;
        RECT 1822.020 -11.020 1825.020 -11.010 ;
        RECT 2002.020 -11.020 2005.020 -11.010 ;
        RECT 2182.020 -11.020 2185.020 -11.010 ;
        RECT 2362.020 -11.020 2365.020 -11.010 ;
        RECT 2542.020 -11.020 2545.020 -11.010 ;
        RECT 2722.020 -11.020 2725.020 -11.010 ;
        RECT 2902.020 -11.020 2905.020 -11.010 ;
        RECT 2936.000 -11.020 2939.000 -11.010 ;
        RECT -19.380 -14.020 2939.000 -11.020 ;
        RECT -19.380 -14.030 -16.380 -14.020 ;
        RECT 22.020 -14.030 25.020 -14.020 ;
        RECT 202.020 -14.030 205.020 -14.020 ;
        RECT 382.020 -14.030 385.020 -14.020 ;
        RECT 562.020 -14.030 565.020 -14.020 ;
        RECT 742.020 -14.030 745.020 -14.020 ;
        RECT 922.020 -14.030 925.020 -14.020 ;
        RECT 1102.020 -14.030 1105.020 -14.020 ;
        RECT 1282.020 -14.030 1285.020 -14.020 ;
        RECT 1462.020 -14.030 1465.020 -14.020 ;
        RECT 1642.020 -14.030 1645.020 -14.020 ;
        RECT 1822.020 -14.030 1825.020 -14.020 ;
        RECT 2002.020 -14.030 2005.020 -14.020 ;
        RECT 2182.020 -14.030 2185.020 -14.020 ;
        RECT 2362.020 -14.030 2365.020 -14.020 ;
        RECT 2542.020 -14.030 2545.020 -14.020 ;
        RECT 2722.020 -14.030 2725.020 -14.020 ;
        RECT 2902.020 -14.030 2905.020 -14.020 ;
        RECT 2936.000 -14.030 2939.000 -14.020 ;
        RECT -28.780 -20.420 -25.780 -20.410 ;
        RECT 40.020 -20.420 43.020 -20.410 ;
        RECT 220.020 -20.420 223.020 -20.410 ;
        RECT 400.020 -20.420 403.020 -20.410 ;
        RECT 580.020 -20.420 583.020 -20.410 ;
        RECT 760.020 -20.420 763.020 -20.410 ;
        RECT 940.020 -20.420 943.020 -20.410 ;
        RECT 1120.020 -20.420 1123.020 -20.410 ;
        RECT 1300.020 -20.420 1303.020 -20.410 ;
        RECT 1480.020 -20.420 1483.020 -20.410 ;
        RECT 1660.020 -20.420 1663.020 -20.410 ;
        RECT 1840.020 -20.420 1843.020 -20.410 ;
        RECT 2020.020 -20.420 2023.020 -20.410 ;
        RECT 2200.020 -20.420 2203.020 -20.410 ;
        RECT 2380.020 -20.420 2383.020 -20.410 ;
        RECT 2560.020 -20.420 2563.020 -20.410 ;
        RECT 2740.020 -20.420 2743.020 -20.410 ;
        RECT 2945.400 -20.420 2948.400 -20.410 ;
        RECT -28.780 -23.420 2948.400 -20.420 ;
        RECT -28.780 -23.430 -25.780 -23.420 ;
        RECT 40.020 -23.430 43.020 -23.420 ;
        RECT 220.020 -23.430 223.020 -23.420 ;
        RECT 400.020 -23.430 403.020 -23.420 ;
        RECT 580.020 -23.430 583.020 -23.420 ;
        RECT 760.020 -23.430 763.020 -23.420 ;
        RECT 940.020 -23.430 943.020 -23.420 ;
        RECT 1120.020 -23.430 1123.020 -23.420 ;
        RECT 1300.020 -23.430 1303.020 -23.420 ;
        RECT 1480.020 -23.430 1483.020 -23.420 ;
        RECT 1660.020 -23.430 1663.020 -23.420 ;
        RECT 1840.020 -23.430 1843.020 -23.420 ;
        RECT 2020.020 -23.430 2023.020 -23.420 ;
        RECT 2200.020 -23.430 2203.020 -23.420 ;
        RECT 2380.020 -23.430 2383.020 -23.420 ;
        RECT 2560.020 -23.430 2563.020 -23.420 ;
        RECT 2740.020 -23.430 2743.020 -23.420 ;
        RECT 2945.400 -23.430 2948.400 -23.420 ;
        RECT -38.180 -29.820 -35.180 -29.810 ;
        RECT 58.020 -29.820 61.020 -29.810 ;
        RECT 238.020 -29.820 241.020 -29.810 ;
        RECT 418.020 -29.820 421.020 -29.810 ;
        RECT 598.020 -29.820 601.020 -29.810 ;
        RECT 778.020 -29.820 781.020 -29.810 ;
        RECT 958.020 -29.820 961.020 -29.810 ;
        RECT 1138.020 -29.820 1141.020 -29.810 ;
        RECT 1318.020 -29.820 1321.020 -29.810 ;
        RECT 1498.020 -29.820 1501.020 -29.810 ;
        RECT 1678.020 -29.820 1681.020 -29.810 ;
        RECT 1858.020 -29.820 1861.020 -29.810 ;
        RECT 2038.020 -29.820 2041.020 -29.810 ;
        RECT 2218.020 -29.820 2221.020 -29.810 ;
        RECT 2398.020 -29.820 2401.020 -29.810 ;
        RECT 2578.020 -29.820 2581.020 -29.810 ;
        RECT 2758.020 -29.820 2761.020 -29.810 ;
        RECT 2954.800 -29.820 2957.800 -29.810 ;
        RECT -38.180 -32.820 2957.800 -29.820 ;
        RECT -38.180 -32.830 -35.180 -32.820 ;
        RECT 58.020 -32.830 61.020 -32.820 ;
        RECT 238.020 -32.830 241.020 -32.820 ;
        RECT 418.020 -32.830 421.020 -32.820 ;
        RECT 598.020 -32.830 601.020 -32.820 ;
        RECT 778.020 -32.830 781.020 -32.820 ;
        RECT 958.020 -32.830 961.020 -32.820 ;
        RECT 1138.020 -32.830 1141.020 -32.820 ;
        RECT 1318.020 -32.830 1321.020 -32.820 ;
        RECT 1498.020 -32.830 1501.020 -32.820 ;
        RECT 1678.020 -32.830 1681.020 -32.820 ;
        RECT 1858.020 -32.830 1861.020 -32.820 ;
        RECT 2038.020 -32.830 2041.020 -32.820 ;
        RECT 2218.020 -32.830 2221.020 -32.820 ;
        RECT 2398.020 -32.830 2401.020 -32.820 ;
        RECT 2578.020 -32.830 2581.020 -32.820 ;
        RECT 2758.020 -32.830 2761.020 -32.820 ;
        RECT 2954.800 -32.830 2957.800 -32.820 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 681.040 3251.235 686.300 3252.140 ;
        RECT 1331.040 3251.235 1336.300 3252.140 ;
        RECT 1931.040 3251.235 1936.300 3252.140 ;
        RECT 2581.040 3251.235 2586.300 3252.140 ;
        RECT 681.480 3250.400 686.300 3251.235 ;
        RECT 1331.480 3250.400 1336.300 3251.235 ;
        RECT 1931.480 3250.400 1936.300 3251.235 ;
        RECT 2581.480 3250.400 2586.300 3251.235 ;
      LAYER via3 ;
        RECT 684.720 3250.440 686.240 3252.050 ;
        RECT 1334.720 3250.440 1336.240 3252.050 ;
        RECT 1934.720 3250.440 1936.240 3252.050 ;
        RECT 2584.720 3250.440 2586.240 3252.050 ;
      LAYER met4 ;
        RECT -42.880 -37.520 -39.880 3557.200 ;
        RECT -33.480 -28.120 -30.480 3547.800 ;
        RECT -24.080 -18.720 -21.080 3538.400 ;
        RECT -14.680 -9.320 -11.680 3529.000 ;
        RECT 94.020 -9.320 97.020 3529.000 ;
        RECT 112.020 -18.720 115.020 3538.400 ;
        RECT 130.020 -28.120 133.020 3547.800 ;
        RECT 148.020 -37.520 151.020 3557.200 ;
        RECT 274.020 -9.320 277.020 3529.000 ;
        RECT 292.020 3271.235 295.020 3538.400 ;
        RECT 310.020 3271.235 313.020 3547.800 ;
        RECT 328.020 3271.235 331.020 3557.200 ;
        RECT 454.020 3271.235 457.020 3529.000 ;
        RECT 472.020 3271.235 475.020 3538.400 ;
        RECT 490.020 3271.235 493.020 3547.800 ;
        RECT 508.020 3271.235 511.020 3557.200 ;
        RECT 634.020 3271.235 637.020 3529.000 ;
        RECT 652.020 3271.235 655.020 3538.400 ;
        RECT 670.020 3271.235 673.020 3547.800 ;
        RECT 688.020 3271.235 691.020 3557.200 ;
        RECT 684.690 2804.060 686.310 3252.140 ;
        RECT 814.020 2715.000 817.020 3529.000 ;
        RECT 832.020 2715.000 835.020 3538.400 ;
        RECT 850.020 2715.000 853.020 3547.800 ;
        RECT 868.020 2715.000 871.020 3557.200 ;
        RECT 994.020 3271.235 997.020 3529.000 ;
        RECT 1012.020 3271.235 1015.020 3538.400 ;
        RECT 1030.020 3271.235 1033.020 3547.800 ;
        RECT 1048.020 3271.235 1051.020 3557.200 ;
        RECT 1174.020 3271.235 1177.020 3529.000 ;
        RECT 1192.020 3271.235 1195.020 3538.400 ;
        RECT 1210.020 3271.235 1213.020 3547.800 ;
        RECT 1228.020 3271.235 1231.020 3557.200 ;
        RECT 1334.690 2804.060 1336.310 3252.140 ;
        RECT 1354.020 2715.000 1357.020 3529.000 ;
        RECT 1372.020 2715.000 1375.020 3538.400 ;
        RECT 1390.020 2715.000 1393.020 3547.800 ;
        RECT 1408.020 2715.000 1411.020 3557.200 ;
        RECT 1534.020 3271.235 1537.020 3529.000 ;
        RECT 1552.020 3271.235 1555.020 3538.400 ;
        RECT 1570.020 3271.235 1573.020 3547.800 ;
        RECT 1588.020 3271.235 1591.020 3557.200 ;
        RECT 1714.020 3271.235 1717.020 3529.000 ;
        RECT 1732.020 3271.235 1735.020 3538.400 ;
        RECT 1750.020 3271.235 1753.020 3547.800 ;
        RECT 1768.020 3271.235 1771.020 3557.200 ;
        RECT 1894.020 3271.235 1897.020 3529.000 ;
        RECT 1912.020 3271.235 1915.020 3538.400 ;
        RECT 1930.020 3271.235 1933.020 3547.800 ;
        RECT 1948.020 3271.235 1951.020 3557.200 ;
        RECT 1934.690 2804.060 1936.310 3252.140 ;
        RECT 397.840 1510.640 399.440 2688.880 ;
        RECT 292.020 -18.720 295.020 1485.000 ;
        RECT 310.020 -28.120 313.020 1485.000 ;
        RECT 328.020 -37.520 331.020 1485.000 ;
        RECT 454.020 -9.320 457.020 1485.000 ;
        RECT 472.020 -18.720 475.020 1485.000 ;
        RECT 490.020 -28.120 493.020 1485.000 ;
        RECT 508.020 -37.520 511.020 1485.000 ;
        RECT 634.020 -9.320 637.020 1485.000 ;
        RECT 652.020 -18.720 655.020 1485.000 ;
        RECT 670.020 -28.120 673.020 1485.000 ;
        RECT 688.020 -37.520 691.020 1485.000 ;
        RECT 814.020 -9.320 817.020 1485.000 ;
        RECT 832.020 -18.720 835.020 1485.000 ;
        RECT 850.020 -28.120 853.020 1485.000 ;
        RECT 868.020 -37.520 871.020 1485.000 ;
        RECT 994.020 -9.320 997.020 1485.000 ;
        RECT 1012.020 -18.720 1015.020 1485.000 ;
        RECT 1030.020 -28.120 1033.020 1485.000 ;
        RECT 1048.020 -37.520 1051.020 1485.000 ;
        RECT 1174.020 -9.320 1177.020 1485.000 ;
        RECT 1192.020 -18.720 1195.020 1485.000 ;
        RECT 1210.020 -28.120 1213.020 1485.000 ;
        RECT 1228.020 -37.520 1231.020 1485.000 ;
        RECT 1354.020 -9.320 1357.020 1485.000 ;
        RECT 1372.020 -18.720 1375.020 1485.000 ;
        RECT 1390.020 -28.120 1393.020 1485.000 ;
        RECT 1408.020 -37.520 1411.020 1485.000 ;
        RECT 1534.020 -9.320 1537.020 2785.000 ;
        RECT 1552.020 -18.720 1555.020 2785.000 ;
        RECT 1570.020 -28.120 1573.020 2785.000 ;
        RECT 1588.020 -37.520 1591.020 2785.000 ;
        RECT 1714.020 -9.320 1717.020 2785.000 ;
        RECT 1732.020 -18.720 1735.020 2785.000 ;
        RECT 1750.020 -28.120 1753.020 2785.000 ;
        RECT 1768.020 -37.520 1771.020 2785.000 ;
        RECT 1894.020 -9.320 1897.020 2785.000 ;
        RECT 1912.020 -18.720 1915.020 2785.000 ;
        RECT 1930.020 -28.120 1933.020 2785.000 ;
        RECT 1948.020 -37.520 1951.020 2785.000 ;
        RECT 2074.020 -9.320 2077.020 3529.000 ;
        RECT 2092.020 -18.720 2095.020 3538.400 ;
        RECT 2110.020 -28.120 2113.020 3547.800 ;
        RECT 2128.020 -37.520 2131.020 3557.200 ;
        RECT 2254.020 3271.235 2257.020 3529.000 ;
        RECT 2272.020 3271.235 2275.020 3538.400 ;
        RECT 2290.020 3271.235 2293.020 3547.800 ;
        RECT 2308.020 3271.235 2311.020 3557.200 ;
        RECT 2434.020 3271.235 2437.020 3529.000 ;
        RECT 2452.020 3271.235 2455.020 3538.400 ;
        RECT 2470.020 3271.235 2473.020 3547.800 ;
        RECT 2488.020 3271.235 2491.020 3557.200 ;
        RECT 2584.690 2804.060 2586.310 3252.140 ;
        RECT 2254.020 -9.320 2257.020 2785.000 ;
        RECT 2272.020 -18.720 2275.020 2785.000 ;
        RECT 2290.020 -28.120 2293.020 2785.000 ;
        RECT 2308.020 -37.520 2311.020 2785.000 ;
        RECT 2434.020 -9.320 2437.020 2785.000 ;
        RECT 2452.020 -18.720 2455.020 2785.000 ;
        RECT 2470.020 -28.120 2473.020 2785.000 ;
        RECT 2488.020 -37.520 2491.020 2785.000 ;
        RECT 2614.020 -9.320 2617.020 3529.000 ;
        RECT 2632.020 -18.720 2635.020 3538.400 ;
        RECT 2650.020 -28.120 2653.020 3547.800 ;
        RECT 2668.020 -37.520 2671.020 3557.200 ;
        RECT 2794.020 -9.320 2797.020 3529.000 ;
        RECT 2812.020 -18.720 2815.020 3538.400 ;
        RECT 2830.020 -28.120 2833.020 3547.800 ;
        RECT 2848.020 -37.520 2851.020 3557.200 ;
        RECT 2931.300 -9.320 2934.300 3529.000 ;
        RECT 2940.700 -18.720 2943.700 3538.400 ;
        RECT 2950.100 -28.120 2953.100 3547.800 ;
        RECT 2959.500 -37.520 2962.500 3557.200 ;
      LAYER via4 ;
        RECT -41.970 3555.910 -40.790 3557.090 ;
        RECT -41.970 3554.310 -40.790 3555.490 ;
        RECT 148.930 3555.910 150.110 3557.090 ;
        RECT 148.930 3554.310 150.110 3555.490 ;
        RECT -41.970 3395.090 -40.790 3396.270 ;
        RECT -41.970 3393.490 -40.790 3394.670 ;
        RECT -41.970 3215.090 -40.790 3216.270 ;
        RECT -41.970 3213.490 -40.790 3214.670 ;
        RECT -41.970 3035.090 -40.790 3036.270 ;
        RECT -41.970 3033.490 -40.790 3034.670 ;
        RECT -41.970 2855.090 -40.790 2856.270 ;
        RECT -41.970 2853.490 -40.790 2854.670 ;
        RECT -41.970 2675.090 -40.790 2676.270 ;
        RECT -41.970 2673.490 -40.790 2674.670 ;
        RECT -41.970 2495.090 -40.790 2496.270 ;
        RECT -41.970 2493.490 -40.790 2494.670 ;
        RECT -41.970 2315.090 -40.790 2316.270 ;
        RECT -41.970 2313.490 -40.790 2314.670 ;
        RECT -41.970 2135.090 -40.790 2136.270 ;
        RECT -41.970 2133.490 -40.790 2134.670 ;
        RECT -41.970 1955.090 -40.790 1956.270 ;
        RECT -41.970 1953.490 -40.790 1954.670 ;
        RECT -41.970 1775.090 -40.790 1776.270 ;
        RECT -41.970 1773.490 -40.790 1774.670 ;
        RECT -41.970 1595.090 -40.790 1596.270 ;
        RECT -41.970 1593.490 -40.790 1594.670 ;
        RECT -41.970 1415.090 -40.790 1416.270 ;
        RECT -41.970 1413.490 -40.790 1414.670 ;
        RECT -41.970 1235.090 -40.790 1236.270 ;
        RECT -41.970 1233.490 -40.790 1234.670 ;
        RECT -41.970 1055.090 -40.790 1056.270 ;
        RECT -41.970 1053.490 -40.790 1054.670 ;
        RECT -41.970 875.090 -40.790 876.270 ;
        RECT -41.970 873.490 -40.790 874.670 ;
        RECT -41.970 695.090 -40.790 696.270 ;
        RECT -41.970 693.490 -40.790 694.670 ;
        RECT -41.970 515.090 -40.790 516.270 ;
        RECT -41.970 513.490 -40.790 514.670 ;
        RECT -41.970 335.090 -40.790 336.270 ;
        RECT -41.970 333.490 -40.790 334.670 ;
        RECT -41.970 155.090 -40.790 156.270 ;
        RECT -41.970 153.490 -40.790 154.670 ;
        RECT -32.570 3546.510 -31.390 3547.690 ;
        RECT -32.570 3544.910 -31.390 3546.090 ;
        RECT 130.930 3546.510 132.110 3547.690 ;
        RECT 130.930 3544.910 132.110 3546.090 ;
        RECT -32.570 3377.090 -31.390 3378.270 ;
        RECT -32.570 3375.490 -31.390 3376.670 ;
        RECT -32.570 3197.090 -31.390 3198.270 ;
        RECT -32.570 3195.490 -31.390 3196.670 ;
        RECT -32.570 3017.090 -31.390 3018.270 ;
        RECT -32.570 3015.490 -31.390 3016.670 ;
        RECT -32.570 2837.090 -31.390 2838.270 ;
        RECT -32.570 2835.490 -31.390 2836.670 ;
        RECT -32.570 2657.090 -31.390 2658.270 ;
        RECT -32.570 2655.490 -31.390 2656.670 ;
        RECT -32.570 2477.090 -31.390 2478.270 ;
        RECT -32.570 2475.490 -31.390 2476.670 ;
        RECT -32.570 2297.090 -31.390 2298.270 ;
        RECT -32.570 2295.490 -31.390 2296.670 ;
        RECT -32.570 2117.090 -31.390 2118.270 ;
        RECT -32.570 2115.490 -31.390 2116.670 ;
        RECT -32.570 1937.090 -31.390 1938.270 ;
        RECT -32.570 1935.490 -31.390 1936.670 ;
        RECT -32.570 1757.090 -31.390 1758.270 ;
        RECT -32.570 1755.490 -31.390 1756.670 ;
        RECT -32.570 1577.090 -31.390 1578.270 ;
        RECT -32.570 1575.490 -31.390 1576.670 ;
        RECT -32.570 1397.090 -31.390 1398.270 ;
        RECT -32.570 1395.490 -31.390 1396.670 ;
        RECT -32.570 1217.090 -31.390 1218.270 ;
        RECT -32.570 1215.490 -31.390 1216.670 ;
        RECT -32.570 1037.090 -31.390 1038.270 ;
        RECT -32.570 1035.490 -31.390 1036.670 ;
        RECT -32.570 857.090 -31.390 858.270 ;
        RECT -32.570 855.490 -31.390 856.670 ;
        RECT -32.570 677.090 -31.390 678.270 ;
        RECT -32.570 675.490 -31.390 676.670 ;
        RECT -32.570 497.090 -31.390 498.270 ;
        RECT -32.570 495.490 -31.390 496.670 ;
        RECT -32.570 317.090 -31.390 318.270 ;
        RECT -32.570 315.490 -31.390 316.670 ;
        RECT -32.570 137.090 -31.390 138.270 ;
        RECT -32.570 135.490 -31.390 136.670 ;
        RECT -23.170 3537.110 -21.990 3538.290 ;
        RECT -23.170 3535.510 -21.990 3536.690 ;
        RECT 112.930 3537.110 114.110 3538.290 ;
        RECT 112.930 3535.510 114.110 3536.690 ;
        RECT -23.170 3359.090 -21.990 3360.270 ;
        RECT -23.170 3357.490 -21.990 3358.670 ;
        RECT -23.170 3179.090 -21.990 3180.270 ;
        RECT -23.170 3177.490 -21.990 3178.670 ;
        RECT -23.170 2999.090 -21.990 3000.270 ;
        RECT -23.170 2997.490 -21.990 2998.670 ;
        RECT -23.170 2819.090 -21.990 2820.270 ;
        RECT -23.170 2817.490 -21.990 2818.670 ;
        RECT -23.170 2639.090 -21.990 2640.270 ;
        RECT -23.170 2637.490 -21.990 2638.670 ;
        RECT -23.170 2459.090 -21.990 2460.270 ;
        RECT -23.170 2457.490 -21.990 2458.670 ;
        RECT -23.170 2279.090 -21.990 2280.270 ;
        RECT -23.170 2277.490 -21.990 2278.670 ;
        RECT -23.170 2099.090 -21.990 2100.270 ;
        RECT -23.170 2097.490 -21.990 2098.670 ;
        RECT -23.170 1919.090 -21.990 1920.270 ;
        RECT -23.170 1917.490 -21.990 1918.670 ;
        RECT -23.170 1739.090 -21.990 1740.270 ;
        RECT -23.170 1737.490 -21.990 1738.670 ;
        RECT -23.170 1559.090 -21.990 1560.270 ;
        RECT -23.170 1557.490 -21.990 1558.670 ;
        RECT -23.170 1379.090 -21.990 1380.270 ;
        RECT -23.170 1377.490 -21.990 1378.670 ;
        RECT -23.170 1199.090 -21.990 1200.270 ;
        RECT -23.170 1197.490 -21.990 1198.670 ;
        RECT -23.170 1019.090 -21.990 1020.270 ;
        RECT -23.170 1017.490 -21.990 1018.670 ;
        RECT -23.170 839.090 -21.990 840.270 ;
        RECT -23.170 837.490 -21.990 838.670 ;
        RECT -23.170 659.090 -21.990 660.270 ;
        RECT -23.170 657.490 -21.990 658.670 ;
        RECT -23.170 479.090 -21.990 480.270 ;
        RECT -23.170 477.490 -21.990 478.670 ;
        RECT -23.170 299.090 -21.990 300.270 ;
        RECT -23.170 297.490 -21.990 298.670 ;
        RECT -23.170 119.090 -21.990 120.270 ;
        RECT -23.170 117.490 -21.990 118.670 ;
        RECT -13.770 3527.710 -12.590 3528.890 ;
        RECT -13.770 3526.110 -12.590 3527.290 ;
        RECT -13.770 3341.090 -12.590 3342.270 ;
        RECT -13.770 3339.490 -12.590 3340.670 ;
        RECT -13.770 3161.090 -12.590 3162.270 ;
        RECT -13.770 3159.490 -12.590 3160.670 ;
        RECT -13.770 2981.090 -12.590 2982.270 ;
        RECT -13.770 2979.490 -12.590 2980.670 ;
        RECT -13.770 2801.090 -12.590 2802.270 ;
        RECT -13.770 2799.490 -12.590 2800.670 ;
        RECT -13.770 2621.090 -12.590 2622.270 ;
        RECT -13.770 2619.490 -12.590 2620.670 ;
        RECT -13.770 2441.090 -12.590 2442.270 ;
        RECT -13.770 2439.490 -12.590 2440.670 ;
        RECT -13.770 2261.090 -12.590 2262.270 ;
        RECT -13.770 2259.490 -12.590 2260.670 ;
        RECT -13.770 2081.090 -12.590 2082.270 ;
        RECT -13.770 2079.490 -12.590 2080.670 ;
        RECT -13.770 1901.090 -12.590 1902.270 ;
        RECT -13.770 1899.490 -12.590 1900.670 ;
        RECT -13.770 1721.090 -12.590 1722.270 ;
        RECT -13.770 1719.490 -12.590 1720.670 ;
        RECT -13.770 1541.090 -12.590 1542.270 ;
        RECT -13.770 1539.490 -12.590 1540.670 ;
        RECT -13.770 1361.090 -12.590 1362.270 ;
        RECT -13.770 1359.490 -12.590 1360.670 ;
        RECT -13.770 1181.090 -12.590 1182.270 ;
        RECT -13.770 1179.490 -12.590 1180.670 ;
        RECT -13.770 1001.090 -12.590 1002.270 ;
        RECT -13.770 999.490 -12.590 1000.670 ;
        RECT -13.770 821.090 -12.590 822.270 ;
        RECT -13.770 819.490 -12.590 820.670 ;
        RECT -13.770 641.090 -12.590 642.270 ;
        RECT -13.770 639.490 -12.590 640.670 ;
        RECT -13.770 461.090 -12.590 462.270 ;
        RECT -13.770 459.490 -12.590 460.670 ;
        RECT -13.770 281.090 -12.590 282.270 ;
        RECT -13.770 279.490 -12.590 280.670 ;
        RECT -13.770 101.090 -12.590 102.270 ;
        RECT -13.770 99.490 -12.590 100.670 ;
        RECT -13.770 -7.610 -12.590 -6.430 ;
        RECT -13.770 -9.210 -12.590 -8.030 ;
        RECT 94.930 3527.710 96.110 3528.890 ;
        RECT 94.930 3526.110 96.110 3527.290 ;
        RECT 94.930 3341.090 96.110 3342.270 ;
        RECT 94.930 3339.490 96.110 3340.670 ;
        RECT 94.930 3161.090 96.110 3162.270 ;
        RECT 94.930 3159.490 96.110 3160.670 ;
        RECT 94.930 2981.090 96.110 2982.270 ;
        RECT 94.930 2979.490 96.110 2980.670 ;
        RECT 94.930 2801.090 96.110 2802.270 ;
        RECT 94.930 2799.490 96.110 2800.670 ;
        RECT 94.930 2621.090 96.110 2622.270 ;
        RECT 94.930 2619.490 96.110 2620.670 ;
        RECT 94.930 2441.090 96.110 2442.270 ;
        RECT 94.930 2439.490 96.110 2440.670 ;
        RECT 94.930 2261.090 96.110 2262.270 ;
        RECT 94.930 2259.490 96.110 2260.670 ;
        RECT 94.930 2081.090 96.110 2082.270 ;
        RECT 94.930 2079.490 96.110 2080.670 ;
        RECT 94.930 1901.090 96.110 1902.270 ;
        RECT 94.930 1899.490 96.110 1900.670 ;
        RECT 94.930 1721.090 96.110 1722.270 ;
        RECT 94.930 1719.490 96.110 1720.670 ;
        RECT 94.930 1541.090 96.110 1542.270 ;
        RECT 94.930 1539.490 96.110 1540.670 ;
        RECT 94.930 1361.090 96.110 1362.270 ;
        RECT 94.930 1359.490 96.110 1360.670 ;
        RECT 94.930 1181.090 96.110 1182.270 ;
        RECT 94.930 1179.490 96.110 1180.670 ;
        RECT 94.930 1001.090 96.110 1002.270 ;
        RECT 94.930 999.490 96.110 1000.670 ;
        RECT 94.930 821.090 96.110 822.270 ;
        RECT 94.930 819.490 96.110 820.670 ;
        RECT 94.930 641.090 96.110 642.270 ;
        RECT 94.930 639.490 96.110 640.670 ;
        RECT 94.930 461.090 96.110 462.270 ;
        RECT 94.930 459.490 96.110 460.670 ;
        RECT 94.930 281.090 96.110 282.270 ;
        RECT 94.930 279.490 96.110 280.670 ;
        RECT 94.930 101.090 96.110 102.270 ;
        RECT 94.930 99.490 96.110 100.670 ;
        RECT 94.930 -7.610 96.110 -6.430 ;
        RECT 94.930 -9.210 96.110 -8.030 ;
        RECT 112.930 3359.090 114.110 3360.270 ;
        RECT 112.930 3357.490 114.110 3358.670 ;
        RECT 112.930 3179.090 114.110 3180.270 ;
        RECT 112.930 3177.490 114.110 3178.670 ;
        RECT 112.930 2999.090 114.110 3000.270 ;
        RECT 112.930 2997.490 114.110 2998.670 ;
        RECT 112.930 2819.090 114.110 2820.270 ;
        RECT 112.930 2817.490 114.110 2818.670 ;
        RECT 112.930 2639.090 114.110 2640.270 ;
        RECT 112.930 2637.490 114.110 2638.670 ;
        RECT 112.930 2459.090 114.110 2460.270 ;
        RECT 112.930 2457.490 114.110 2458.670 ;
        RECT 112.930 2279.090 114.110 2280.270 ;
        RECT 112.930 2277.490 114.110 2278.670 ;
        RECT 112.930 2099.090 114.110 2100.270 ;
        RECT 112.930 2097.490 114.110 2098.670 ;
        RECT 112.930 1919.090 114.110 1920.270 ;
        RECT 112.930 1917.490 114.110 1918.670 ;
        RECT 112.930 1739.090 114.110 1740.270 ;
        RECT 112.930 1737.490 114.110 1738.670 ;
        RECT 112.930 1559.090 114.110 1560.270 ;
        RECT 112.930 1557.490 114.110 1558.670 ;
        RECT 112.930 1379.090 114.110 1380.270 ;
        RECT 112.930 1377.490 114.110 1378.670 ;
        RECT 112.930 1199.090 114.110 1200.270 ;
        RECT 112.930 1197.490 114.110 1198.670 ;
        RECT 112.930 1019.090 114.110 1020.270 ;
        RECT 112.930 1017.490 114.110 1018.670 ;
        RECT 112.930 839.090 114.110 840.270 ;
        RECT 112.930 837.490 114.110 838.670 ;
        RECT 112.930 659.090 114.110 660.270 ;
        RECT 112.930 657.490 114.110 658.670 ;
        RECT 112.930 479.090 114.110 480.270 ;
        RECT 112.930 477.490 114.110 478.670 ;
        RECT 112.930 299.090 114.110 300.270 ;
        RECT 112.930 297.490 114.110 298.670 ;
        RECT 112.930 119.090 114.110 120.270 ;
        RECT 112.930 117.490 114.110 118.670 ;
        RECT -23.170 -17.010 -21.990 -15.830 ;
        RECT -23.170 -18.610 -21.990 -17.430 ;
        RECT 112.930 -17.010 114.110 -15.830 ;
        RECT 112.930 -18.610 114.110 -17.430 ;
        RECT 130.930 3377.090 132.110 3378.270 ;
        RECT 130.930 3375.490 132.110 3376.670 ;
        RECT 130.930 3197.090 132.110 3198.270 ;
        RECT 130.930 3195.490 132.110 3196.670 ;
        RECT 130.930 3017.090 132.110 3018.270 ;
        RECT 130.930 3015.490 132.110 3016.670 ;
        RECT 130.930 2837.090 132.110 2838.270 ;
        RECT 130.930 2835.490 132.110 2836.670 ;
        RECT 130.930 2657.090 132.110 2658.270 ;
        RECT 130.930 2655.490 132.110 2656.670 ;
        RECT 130.930 2477.090 132.110 2478.270 ;
        RECT 130.930 2475.490 132.110 2476.670 ;
        RECT 130.930 2297.090 132.110 2298.270 ;
        RECT 130.930 2295.490 132.110 2296.670 ;
        RECT 130.930 2117.090 132.110 2118.270 ;
        RECT 130.930 2115.490 132.110 2116.670 ;
        RECT 130.930 1937.090 132.110 1938.270 ;
        RECT 130.930 1935.490 132.110 1936.670 ;
        RECT 130.930 1757.090 132.110 1758.270 ;
        RECT 130.930 1755.490 132.110 1756.670 ;
        RECT 130.930 1577.090 132.110 1578.270 ;
        RECT 130.930 1575.490 132.110 1576.670 ;
        RECT 130.930 1397.090 132.110 1398.270 ;
        RECT 130.930 1395.490 132.110 1396.670 ;
        RECT 130.930 1217.090 132.110 1218.270 ;
        RECT 130.930 1215.490 132.110 1216.670 ;
        RECT 130.930 1037.090 132.110 1038.270 ;
        RECT 130.930 1035.490 132.110 1036.670 ;
        RECT 130.930 857.090 132.110 858.270 ;
        RECT 130.930 855.490 132.110 856.670 ;
        RECT 130.930 677.090 132.110 678.270 ;
        RECT 130.930 675.490 132.110 676.670 ;
        RECT 130.930 497.090 132.110 498.270 ;
        RECT 130.930 495.490 132.110 496.670 ;
        RECT 130.930 317.090 132.110 318.270 ;
        RECT 130.930 315.490 132.110 316.670 ;
        RECT 130.930 137.090 132.110 138.270 ;
        RECT 130.930 135.490 132.110 136.670 ;
        RECT -32.570 -26.410 -31.390 -25.230 ;
        RECT -32.570 -28.010 -31.390 -26.830 ;
        RECT 130.930 -26.410 132.110 -25.230 ;
        RECT 130.930 -28.010 132.110 -26.830 ;
        RECT 328.930 3555.910 330.110 3557.090 ;
        RECT 328.930 3554.310 330.110 3555.490 ;
        RECT 310.930 3546.510 312.110 3547.690 ;
        RECT 310.930 3544.910 312.110 3546.090 ;
        RECT 292.930 3537.110 294.110 3538.290 ;
        RECT 292.930 3535.510 294.110 3536.690 ;
        RECT 148.930 3395.090 150.110 3396.270 ;
        RECT 148.930 3393.490 150.110 3394.670 ;
        RECT 148.930 3215.090 150.110 3216.270 ;
        RECT 148.930 3213.490 150.110 3214.670 ;
        RECT 148.930 3035.090 150.110 3036.270 ;
        RECT 148.930 3033.490 150.110 3034.670 ;
        RECT 148.930 2855.090 150.110 2856.270 ;
        RECT 148.930 2853.490 150.110 2854.670 ;
        RECT 148.930 2675.090 150.110 2676.270 ;
        RECT 148.930 2673.490 150.110 2674.670 ;
        RECT 148.930 2495.090 150.110 2496.270 ;
        RECT 148.930 2493.490 150.110 2494.670 ;
        RECT 148.930 2315.090 150.110 2316.270 ;
        RECT 148.930 2313.490 150.110 2314.670 ;
        RECT 148.930 2135.090 150.110 2136.270 ;
        RECT 148.930 2133.490 150.110 2134.670 ;
        RECT 148.930 1955.090 150.110 1956.270 ;
        RECT 148.930 1953.490 150.110 1954.670 ;
        RECT 148.930 1775.090 150.110 1776.270 ;
        RECT 148.930 1773.490 150.110 1774.670 ;
        RECT 148.930 1595.090 150.110 1596.270 ;
        RECT 148.930 1593.490 150.110 1594.670 ;
        RECT 148.930 1415.090 150.110 1416.270 ;
        RECT 148.930 1413.490 150.110 1414.670 ;
        RECT 148.930 1235.090 150.110 1236.270 ;
        RECT 148.930 1233.490 150.110 1234.670 ;
        RECT 148.930 1055.090 150.110 1056.270 ;
        RECT 148.930 1053.490 150.110 1054.670 ;
        RECT 148.930 875.090 150.110 876.270 ;
        RECT 148.930 873.490 150.110 874.670 ;
        RECT 148.930 695.090 150.110 696.270 ;
        RECT 148.930 693.490 150.110 694.670 ;
        RECT 148.930 515.090 150.110 516.270 ;
        RECT 148.930 513.490 150.110 514.670 ;
        RECT 148.930 335.090 150.110 336.270 ;
        RECT 148.930 333.490 150.110 334.670 ;
        RECT 148.930 155.090 150.110 156.270 ;
        RECT 148.930 153.490 150.110 154.670 ;
        RECT -41.970 -35.810 -40.790 -34.630 ;
        RECT -41.970 -37.410 -40.790 -36.230 ;
        RECT 274.930 3527.710 276.110 3528.890 ;
        RECT 274.930 3526.110 276.110 3527.290 ;
        RECT 274.930 3341.090 276.110 3342.270 ;
        RECT 274.930 3339.490 276.110 3340.670 ;
        RECT 292.930 3359.090 294.110 3360.270 ;
        RECT 292.930 3357.490 294.110 3358.670 ;
        RECT 310.930 3377.090 312.110 3378.270 ;
        RECT 310.930 3375.490 312.110 3376.670 ;
        RECT 508.930 3555.910 510.110 3557.090 ;
        RECT 508.930 3554.310 510.110 3555.490 ;
        RECT 490.930 3546.510 492.110 3547.690 ;
        RECT 490.930 3544.910 492.110 3546.090 ;
        RECT 472.930 3537.110 474.110 3538.290 ;
        RECT 472.930 3535.510 474.110 3536.690 ;
        RECT 328.930 3395.090 330.110 3396.270 ;
        RECT 328.930 3393.490 330.110 3394.670 ;
        RECT 454.930 3527.710 456.110 3528.890 ;
        RECT 454.930 3526.110 456.110 3527.290 ;
        RECT 454.930 3341.090 456.110 3342.270 ;
        RECT 454.930 3339.490 456.110 3340.670 ;
        RECT 472.930 3359.090 474.110 3360.270 ;
        RECT 472.930 3357.490 474.110 3358.670 ;
        RECT 490.930 3377.090 492.110 3378.270 ;
        RECT 490.930 3375.490 492.110 3376.670 ;
        RECT 688.930 3555.910 690.110 3557.090 ;
        RECT 688.930 3554.310 690.110 3555.490 ;
        RECT 670.930 3546.510 672.110 3547.690 ;
        RECT 670.930 3544.910 672.110 3546.090 ;
        RECT 652.930 3537.110 654.110 3538.290 ;
        RECT 652.930 3535.510 654.110 3536.690 ;
        RECT 508.930 3395.090 510.110 3396.270 ;
        RECT 508.930 3393.490 510.110 3394.670 ;
        RECT 634.930 3527.710 636.110 3528.890 ;
        RECT 634.930 3526.110 636.110 3527.290 ;
        RECT 634.930 3341.090 636.110 3342.270 ;
        RECT 634.930 3339.490 636.110 3340.670 ;
        RECT 652.930 3359.090 654.110 3360.270 ;
        RECT 652.930 3357.490 654.110 3358.670 ;
        RECT 670.930 3377.090 672.110 3378.270 ;
        RECT 670.930 3375.490 672.110 3376.670 ;
        RECT 868.930 3555.910 870.110 3557.090 ;
        RECT 868.930 3554.310 870.110 3555.490 ;
        RECT 850.930 3546.510 852.110 3547.690 ;
        RECT 850.930 3544.910 852.110 3546.090 ;
        RECT 832.930 3537.110 834.110 3538.290 ;
        RECT 832.930 3535.510 834.110 3536.690 ;
        RECT 688.930 3395.090 690.110 3396.270 ;
        RECT 688.930 3393.490 690.110 3394.670 ;
        RECT 814.930 3527.710 816.110 3528.890 ;
        RECT 814.930 3526.110 816.110 3527.290 ;
        RECT 814.930 3341.090 816.110 3342.270 ;
        RECT 814.930 3339.490 816.110 3340.670 ;
        RECT 274.930 3161.090 276.110 3162.270 ;
        RECT 274.930 3159.490 276.110 3160.670 ;
        RECT 274.930 2981.090 276.110 2982.270 ;
        RECT 274.930 2979.490 276.110 2980.670 ;
        RECT 684.910 3215.090 686.090 3216.270 ;
        RECT 684.910 3213.490 686.090 3214.670 ;
        RECT 684.910 3197.090 686.090 3198.270 ;
        RECT 684.910 3195.490 686.090 3196.670 ;
        RECT 684.910 3179.090 686.090 3180.270 ;
        RECT 684.910 3177.490 686.090 3178.670 ;
        RECT 684.910 3161.090 686.090 3162.270 ;
        RECT 684.910 3159.490 686.090 3160.670 ;
        RECT 684.910 3035.090 686.090 3036.270 ;
        RECT 684.910 3033.490 686.090 3034.670 ;
        RECT 684.910 3017.090 686.090 3018.270 ;
        RECT 684.910 3015.490 686.090 3016.670 ;
        RECT 684.910 2999.090 686.090 3000.270 ;
        RECT 684.910 2997.490 686.090 2998.670 ;
        RECT 684.910 2981.090 686.090 2982.270 ;
        RECT 684.910 2979.490 686.090 2980.670 ;
        RECT 684.910 2855.090 686.090 2856.270 ;
        RECT 684.910 2853.490 686.090 2854.670 ;
        RECT 684.910 2837.090 686.090 2838.270 ;
        RECT 684.910 2835.490 686.090 2836.670 ;
        RECT 684.910 2819.090 686.090 2820.270 ;
        RECT 684.910 2817.490 686.090 2818.670 ;
        RECT 814.930 3161.090 816.110 3162.270 ;
        RECT 814.930 3159.490 816.110 3160.670 ;
        RECT 814.930 2981.090 816.110 2982.270 ;
        RECT 814.930 2979.490 816.110 2980.670 ;
        RECT 274.930 2801.090 276.110 2802.270 ;
        RECT 274.930 2799.490 276.110 2800.670 ;
        RECT 814.930 2801.090 816.110 2802.270 ;
        RECT 814.930 2799.490 816.110 2800.670 ;
        RECT 832.930 3359.090 834.110 3360.270 ;
        RECT 832.930 3357.490 834.110 3358.670 ;
        RECT 832.930 3179.090 834.110 3180.270 ;
        RECT 832.930 3177.490 834.110 3178.670 ;
        RECT 832.930 2999.090 834.110 3000.270 ;
        RECT 832.930 2997.490 834.110 2998.670 ;
        RECT 832.930 2819.090 834.110 2820.270 ;
        RECT 832.930 2817.490 834.110 2818.670 ;
        RECT 850.930 3377.090 852.110 3378.270 ;
        RECT 850.930 3375.490 852.110 3376.670 ;
        RECT 850.930 3197.090 852.110 3198.270 ;
        RECT 850.930 3195.490 852.110 3196.670 ;
        RECT 850.930 3017.090 852.110 3018.270 ;
        RECT 850.930 3015.490 852.110 3016.670 ;
        RECT 850.930 2837.090 852.110 2838.270 ;
        RECT 850.930 2835.490 852.110 2836.670 ;
        RECT 1048.930 3555.910 1050.110 3557.090 ;
        RECT 1048.930 3554.310 1050.110 3555.490 ;
        RECT 1030.930 3546.510 1032.110 3547.690 ;
        RECT 1030.930 3544.910 1032.110 3546.090 ;
        RECT 1012.930 3537.110 1014.110 3538.290 ;
        RECT 1012.930 3535.510 1014.110 3536.690 ;
        RECT 868.930 3395.090 870.110 3396.270 ;
        RECT 868.930 3393.490 870.110 3394.670 ;
        RECT 994.930 3527.710 996.110 3528.890 ;
        RECT 994.930 3526.110 996.110 3527.290 ;
        RECT 994.930 3341.090 996.110 3342.270 ;
        RECT 994.930 3339.490 996.110 3340.670 ;
        RECT 1012.930 3359.090 1014.110 3360.270 ;
        RECT 1012.930 3357.490 1014.110 3358.670 ;
        RECT 1030.930 3377.090 1032.110 3378.270 ;
        RECT 1030.930 3375.490 1032.110 3376.670 ;
        RECT 1228.930 3555.910 1230.110 3557.090 ;
        RECT 1228.930 3554.310 1230.110 3555.490 ;
        RECT 1210.930 3546.510 1212.110 3547.690 ;
        RECT 1210.930 3544.910 1212.110 3546.090 ;
        RECT 1192.930 3537.110 1194.110 3538.290 ;
        RECT 1192.930 3535.510 1194.110 3536.690 ;
        RECT 1048.930 3395.090 1050.110 3396.270 ;
        RECT 1048.930 3393.490 1050.110 3394.670 ;
        RECT 1174.930 3527.710 1176.110 3528.890 ;
        RECT 1174.930 3526.110 1176.110 3527.290 ;
        RECT 1174.930 3341.090 1176.110 3342.270 ;
        RECT 1174.930 3339.490 1176.110 3340.670 ;
        RECT 1192.930 3359.090 1194.110 3360.270 ;
        RECT 1192.930 3357.490 1194.110 3358.670 ;
        RECT 1210.930 3377.090 1212.110 3378.270 ;
        RECT 1210.930 3375.490 1212.110 3376.670 ;
        RECT 1408.930 3555.910 1410.110 3557.090 ;
        RECT 1408.930 3554.310 1410.110 3555.490 ;
        RECT 1390.930 3546.510 1392.110 3547.690 ;
        RECT 1390.930 3544.910 1392.110 3546.090 ;
        RECT 1372.930 3537.110 1374.110 3538.290 ;
        RECT 1372.930 3535.510 1374.110 3536.690 ;
        RECT 1228.930 3395.090 1230.110 3396.270 ;
        RECT 1228.930 3393.490 1230.110 3394.670 ;
        RECT 1354.930 3527.710 1356.110 3528.890 ;
        RECT 1354.930 3526.110 1356.110 3527.290 ;
        RECT 1354.930 3341.090 1356.110 3342.270 ;
        RECT 1354.930 3339.490 1356.110 3340.670 ;
        RECT 868.930 3215.090 870.110 3216.270 ;
        RECT 868.930 3213.490 870.110 3214.670 ;
        RECT 868.930 3035.090 870.110 3036.270 ;
        RECT 868.930 3033.490 870.110 3034.670 ;
        RECT 868.930 2855.090 870.110 2856.270 ;
        RECT 868.930 2853.490 870.110 2854.670 ;
        RECT 1334.910 3215.090 1336.090 3216.270 ;
        RECT 1334.910 3213.490 1336.090 3214.670 ;
        RECT 1334.910 3197.090 1336.090 3198.270 ;
        RECT 1334.910 3195.490 1336.090 3196.670 ;
        RECT 1334.910 3179.090 1336.090 3180.270 ;
        RECT 1334.910 3177.490 1336.090 3178.670 ;
        RECT 1334.910 3161.090 1336.090 3162.270 ;
        RECT 1334.910 3159.490 1336.090 3160.670 ;
        RECT 1334.910 3035.090 1336.090 3036.270 ;
        RECT 1334.910 3033.490 1336.090 3034.670 ;
        RECT 1334.910 3017.090 1336.090 3018.270 ;
        RECT 1334.910 3015.490 1336.090 3016.670 ;
        RECT 1334.910 2999.090 1336.090 3000.270 ;
        RECT 1334.910 2997.490 1336.090 2998.670 ;
        RECT 1334.910 2981.090 1336.090 2982.270 ;
        RECT 1334.910 2979.490 1336.090 2980.670 ;
        RECT 1334.910 2855.090 1336.090 2856.270 ;
        RECT 1334.910 2853.490 1336.090 2854.670 ;
        RECT 1334.910 2837.090 1336.090 2838.270 ;
        RECT 1334.910 2835.490 1336.090 2836.670 ;
        RECT 1334.910 2819.090 1336.090 2820.270 ;
        RECT 1334.910 2817.490 1336.090 2818.670 ;
        RECT 1354.930 3161.090 1356.110 3162.270 ;
        RECT 1354.930 3159.490 1356.110 3160.670 ;
        RECT 1354.930 2981.090 1356.110 2982.270 ;
        RECT 1354.930 2979.490 1356.110 2980.670 ;
        RECT 1354.930 2801.090 1356.110 2802.270 ;
        RECT 1354.930 2799.490 1356.110 2800.670 ;
        RECT 1372.930 3359.090 1374.110 3360.270 ;
        RECT 1372.930 3357.490 1374.110 3358.670 ;
        RECT 1372.930 3179.090 1374.110 3180.270 ;
        RECT 1372.930 3177.490 1374.110 3178.670 ;
        RECT 1372.930 2999.090 1374.110 3000.270 ;
        RECT 1372.930 2997.490 1374.110 2998.670 ;
        RECT 1372.930 2819.090 1374.110 2820.270 ;
        RECT 1372.930 2817.490 1374.110 2818.670 ;
        RECT 1390.930 3377.090 1392.110 3378.270 ;
        RECT 1390.930 3375.490 1392.110 3376.670 ;
        RECT 1390.930 3197.090 1392.110 3198.270 ;
        RECT 1390.930 3195.490 1392.110 3196.670 ;
        RECT 1390.930 3017.090 1392.110 3018.270 ;
        RECT 1390.930 3015.490 1392.110 3016.670 ;
        RECT 1390.930 2837.090 1392.110 2838.270 ;
        RECT 1390.930 2835.490 1392.110 2836.670 ;
        RECT 1588.930 3555.910 1590.110 3557.090 ;
        RECT 1588.930 3554.310 1590.110 3555.490 ;
        RECT 1570.930 3546.510 1572.110 3547.690 ;
        RECT 1570.930 3544.910 1572.110 3546.090 ;
        RECT 1552.930 3537.110 1554.110 3538.290 ;
        RECT 1552.930 3535.510 1554.110 3536.690 ;
        RECT 1408.930 3395.090 1410.110 3396.270 ;
        RECT 1408.930 3393.490 1410.110 3394.670 ;
        RECT 1534.930 3527.710 1536.110 3528.890 ;
        RECT 1534.930 3526.110 1536.110 3527.290 ;
        RECT 1534.930 3341.090 1536.110 3342.270 ;
        RECT 1534.930 3339.490 1536.110 3340.670 ;
        RECT 1552.930 3359.090 1554.110 3360.270 ;
        RECT 1552.930 3357.490 1554.110 3358.670 ;
        RECT 1570.930 3377.090 1572.110 3378.270 ;
        RECT 1570.930 3375.490 1572.110 3376.670 ;
        RECT 1768.930 3555.910 1770.110 3557.090 ;
        RECT 1768.930 3554.310 1770.110 3555.490 ;
        RECT 1750.930 3546.510 1752.110 3547.690 ;
        RECT 1750.930 3544.910 1752.110 3546.090 ;
        RECT 1732.930 3537.110 1734.110 3538.290 ;
        RECT 1732.930 3535.510 1734.110 3536.690 ;
        RECT 1588.930 3395.090 1590.110 3396.270 ;
        RECT 1588.930 3393.490 1590.110 3394.670 ;
        RECT 1714.930 3527.710 1716.110 3528.890 ;
        RECT 1714.930 3526.110 1716.110 3527.290 ;
        RECT 1714.930 3341.090 1716.110 3342.270 ;
        RECT 1714.930 3339.490 1716.110 3340.670 ;
        RECT 1732.930 3359.090 1734.110 3360.270 ;
        RECT 1732.930 3357.490 1734.110 3358.670 ;
        RECT 1750.930 3377.090 1752.110 3378.270 ;
        RECT 1750.930 3375.490 1752.110 3376.670 ;
        RECT 1948.930 3555.910 1950.110 3557.090 ;
        RECT 1948.930 3554.310 1950.110 3555.490 ;
        RECT 1930.930 3546.510 1932.110 3547.690 ;
        RECT 1930.930 3544.910 1932.110 3546.090 ;
        RECT 1912.930 3537.110 1914.110 3538.290 ;
        RECT 1912.930 3535.510 1914.110 3536.690 ;
        RECT 1768.930 3395.090 1770.110 3396.270 ;
        RECT 1768.930 3393.490 1770.110 3394.670 ;
        RECT 1894.930 3527.710 1896.110 3528.890 ;
        RECT 1894.930 3526.110 1896.110 3527.290 ;
        RECT 1894.930 3341.090 1896.110 3342.270 ;
        RECT 1894.930 3339.490 1896.110 3340.670 ;
        RECT 1912.930 3359.090 1914.110 3360.270 ;
        RECT 1912.930 3357.490 1914.110 3358.670 ;
        RECT 1930.930 3377.090 1932.110 3378.270 ;
        RECT 1930.930 3375.490 1932.110 3376.670 ;
        RECT 2128.930 3555.910 2130.110 3557.090 ;
        RECT 2128.930 3554.310 2130.110 3555.490 ;
        RECT 2110.930 3546.510 2112.110 3547.690 ;
        RECT 2110.930 3544.910 2112.110 3546.090 ;
        RECT 2092.930 3537.110 2094.110 3538.290 ;
        RECT 2092.930 3535.510 2094.110 3536.690 ;
        RECT 1948.930 3395.090 1950.110 3396.270 ;
        RECT 1948.930 3393.490 1950.110 3394.670 ;
        RECT 2074.930 3527.710 2076.110 3528.890 ;
        RECT 2074.930 3526.110 2076.110 3527.290 ;
        RECT 2074.930 3341.090 2076.110 3342.270 ;
        RECT 2074.930 3339.490 2076.110 3340.670 ;
        RECT 1408.930 3215.090 1410.110 3216.270 ;
        RECT 1408.930 3213.490 1410.110 3214.670 ;
        RECT 1408.930 3035.090 1410.110 3036.270 ;
        RECT 1408.930 3033.490 1410.110 3034.670 ;
        RECT 1408.930 2855.090 1410.110 2856.270 ;
        RECT 1408.930 2853.490 1410.110 2854.670 ;
        RECT 1934.910 3215.090 1936.090 3216.270 ;
        RECT 1934.910 3213.490 1936.090 3214.670 ;
        RECT 1934.910 3197.090 1936.090 3198.270 ;
        RECT 1934.910 3195.490 1936.090 3196.670 ;
        RECT 1934.910 3179.090 1936.090 3180.270 ;
        RECT 1934.910 3177.490 1936.090 3178.670 ;
        RECT 1934.910 3161.090 1936.090 3162.270 ;
        RECT 1934.910 3159.490 1936.090 3160.670 ;
        RECT 1934.910 3035.090 1936.090 3036.270 ;
        RECT 1934.910 3033.490 1936.090 3034.670 ;
        RECT 1934.910 3017.090 1936.090 3018.270 ;
        RECT 1934.910 3015.490 1936.090 3016.670 ;
        RECT 1934.910 2999.090 1936.090 3000.270 ;
        RECT 1934.910 2997.490 1936.090 2998.670 ;
        RECT 1934.910 2981.090 1936.090 2982.270 ;
        RECT 1934.910 2979.490 1936.090 2980.670 ;
        RECT 1934.910 2855.090 1936.090 2856.270 ;
        RECT 1934.910 2853.490 1936.090 2854.670 ;
        RECT 1934.910 2837.090 1936.090 2838.270 ;
        RECT 1934.910 2835.490 1936.090 2836.670 ;
        RECT 1934.910 2819.090 1936.090 2820.270 ;
        RECT 1934.910 2817.490 1936.090 2818.670 ;
        RECT 2074.930 3161.090 2076.110 3162.270 ;
        RECT 2074.930 3159.490 2076.110 3160.670 ;
        RECT 2074.930 2981.090 2076.110 2982.270 ;
        RECT 2074.930 2979.490 2076.110 2980.670 ;
        RECT 2074.930 2801.090 2076.110 2802.270 ;
        RECT 2074.930 2799.490 2076.110 2800.670 ;
        RECT 274.930 2621.090 276.110 2622.270 ;
        RECT 274.930 2619.490 276.110 2620.670 ;
        RECT 274.930 2441.090 276.110 2442.270 ;
        RECT 274.930 2439.490 276.110 2440.670 ;
        RECT 274.930 2261.090 276.110 2262.270 ;
        RECT 274.930 2259.490 276.110 2260.670 ;
        RECT 274.930 2081.090 276.110 2082.270 ;
        RECT 274.930 2079.490 276.110 2080.670 ;
        RECT 274.930 1901.090 276.110 1902.270 ;
        RECT 274.930 1899.490 276.110 1900.670 ;
        RECT 274.930 1721.090 276.110 1722.270 ;
        RECT 274.930 1719.490 276.110 1720.670 ;
        RECT 274.930 1541.090 276.110 1542.270 ;
        RECT 274.930 1539.490 276.110 1540.670 ;
        RECT 398.050 2675.090 399.230 2676.270 ;
        RECT 398.050 2673.490 399.230 2674.670 ;
        RECT 398.050 2657.090 399.230 2658.270 ;
        RECT 398.050 2655.490 399.230 2656.670 ;
        RECT 398.050 2639.090 399.230 2640.270 ;
        RECT 398.050 2637.490 399.230 2638.670 ;
        RECT 398.050 2621.090 399.230 2622.270 ;
        RECT 398.050 2619.490 399.230 2620.670 ;
        RECT 398.050 2495.090 399.230 2496.270 ;
        RECT 398.050 2493.490 399.230 2494.670 ;
        RECT 398.050 2477.090 399.230 2478.270 ;
        RECT 398.050 2475.490 399.230 2476.670 ;
        RECT 398.050 2459.090 399.230 2460.270 ;
        RECT 398.050 2457.490 399.230 2458.670 ;
        RECT 398.050 2441.090 399.230 2442.270 ;
        RECT 398.050 2439.490 399.230 2440.670 ;
        RECT 398.050 2315.090 399.230 2316.270 ;
        RECT 398.050 2313.490 399.230 2314.670 ;
        RECT 398.050 2297.090 399.230 2298.270 ;
        RECT 398.050 2295.490 399.230 2296.670 ;
        RECT 398.050 2279.090 399.230 2280.270 ;
        RECT 398.050 2277.490 399.230 2278.670 ;
        RECT 398.050 2261.090 399.230 2262.270 ;
        RECT 398.050 2259.490 399.230 2260.670 ;
        RECT 398.050 2135.090 399.230 2136.270 ;
        RECT 398.050 2133.490 399.230 2134.670 ;
        RECT 398.050 2117.090 399.230 2118.270 ;
        RECT 398.050 2115.490 399.230 2116.670 ;
        RECT 398.050 2099.090 399.230 2100.270 ;
        RECT 398.050 2097.490 399.230 2098.670 ;
        RECT 398.050 2081.090 399.230 2082.270 ;
        RECT 398.050 2079.490 399.230 2080.670 ;
        RECT 398.050 1955.090 399.230 1956.270 ;
        RECT 398.050 1953.490 399.230 1954.670 ;
        RECT 398.050 1937.090 399.230 1938.270 ;
        RECT 398.050 1935.490 399.230 1936.670 ;
        RECT 398.050 1919.090 399.230 1920.270 ;
        RECT 398.050 1917.490 399.230 1918.670 ;
        RECT 398.050 1901.090 399.230 1902.270 ;
        RECT 398.050 1899.490 399.230 1900.670 ;
        RECT 398.050 1775.090 399.230 1776.270 ;
        RECT 398.050 1773.490 399.230 1774.670 ;
        RECT 398.050 1757.090 399.230 1758.270 ;
        RECT 398.050 1755.490 399.230 1756.670 ;
        RECT 398.050 1739.090 399.230 1740.270 ;
        RECT 398.050 1737.490 399.230 1738.670 ;
        RECT 398.050 1721.090 399.230 1722.270 ;
        RECT 398.050 1719.490 399.230 1720.670 ;
        RECT 398.050 1595.090 399.230 1596.270 ;
        RECT 398.050 1593.490 399.230 1594.670 ;
        RECT 398.050 1577.090 399.230 1578.270 ;
        RECT 398.050 1575.490 399.230 1576.670 ;
        RECT 398.050 1559.090 399.230 1560.270 ;
        RECT 398.050 1557.490 399.230 1558.670 ;
        RECT 398.050 1541.090 399.230 1542.270 ;
        RECT 398.050 1539.490 399.230 1540.670 ;
        RECT 1534.930 2621.090 1536.110 2622.270 ;
        RECT 1534.930 2619.490 1536.110 2620.670 ;
        RECT 1534.930 2441.090 1536.110 2442.270 ;
        RECT 1534.930 2439.490 1536.110 2440.670 ;
        RECT 1534.930 2261.090 1536.110 2262.270 ;
        RECT 1534.930 2259.490 1536.110 2260.670 ;
        RECT 1534.930 2081.090 1536.110 2082.270 ;
        RECT 1534.930 2079.490 1536.110 2080.670 ;
        RECT 1534.930 1901.090 1536.110 1902.270 ;
        RECT 1534.930 1899.490 1536.110 1900.670 ;
        RECT 1534.930 1721.090 1536.110 1722.270 ;
        RECT 1534.930 1719.490 1536.110 1720.670 ;
        RECT 1534.930 1541.090 1536.110 1542.270 ;
        RECT 1534.930 1539.490 1536.110 1540.670 ;
        RECT 274.930 1361.090 276.110 1362.270 ;
        RECT 274.930 1359.490 276.110 1360.670 ;
        RECT 274.930 1181.090 276.110 1182.270 ;
        RECT 274.930 1179.490 276.110 1180.670 ;
        RECT 274.930 1001.090 276.110 1002.270 ;
        RECT 274.930 999.490 276.110 1000.670 ;
        RECT 274.930 821.090 276.110 822.270 ;
        RECT 274.930 819.490 276.110 820.670 ;
        RECT 274.930 641.090 276.110 642.270 ;
        RECT 274.930 639.490 276.110 640.670 ;
        RECT 274.930 461.090 276.110 462.270 ;
        RECT 274.930 459.490 276.110 460.670 ;
        RECT 274.930 281.090 276.110 282.270 ;
        RECT 274.930 279.490 276.110 280.670 ;
        RECT 274.930 101.090 276.110 102.270 ;
        RECT 274.930 99.490 276.110 100.670 ;
        RECT 274.930 -7.610 276.110 -6.430 ;
        RECT 274.930 -9.210 276.110 -8.030 ;
        RECT 292.930 1379.090 294.110 1380.270 ;
        RECT 292.930 1377.490 294.110 1378.670 ;
        RECT 292.930 1199.090 294.110 1200.270 ;
        RECT 292.930 1197.490 294.110 1198.670 ;
        RECT 292.930 1019.090 294.110 1020.270 ;
        RECT 292.930 1017.490 294.110 1018.670 ;
        RECT 292.930 839.090 294.110 840.270 ;
        RECT 292.930 837.490 294.110 838.670 ;
        RECT 292.930 659.090 294.110 660.270 ;
        RECT 292.930 657.490 294.110 658.670 ;
        RECT 292.930 479.090 294.110 480.270 ;
        RECT 292.930 477.490 294.110 478.670 ;
        RECT 292.930 299.090 294.110 300.270 ;
        RECT 292.930 297.490 294.110 298.670 ;
        RECT 292.930 119.090 294.110 120.270 ;
        RECT 292.930 117.490 294.110 118.670 ;
        RECT 292.930 -17.010 294.110 -15.830 ;
        RECT 292.930 -18.610 294.110 -17.430 ;
        RECT 310.930 1397.090 312.110 1398.270 ;
        RECT 310.930 1395.490 312.110 1396.670 ;
        RECT 310.930 1217.090 312.110 1218.270 ;
        RECT 310.930 1215.490 312.110 1216.670 ;
        RECT 310.930 1037.090 312.110 1038.270 ;
        RECT 310.930 1035.490 312.110 1036.670 ;
        RECT 310.930 857.090 312.110 858.270 ;
        RECT 310.930 855.490 312.110 856.670 ;
        RECT 310.930 677.090 312.110 678.270 ;
        RECT 310.930 675.490 312.110 676.670 ;
        RECT 310.930 497.090 312.110 498.270 ;
        RECT 310.930 495.490 312.110 496.670 ;
        RECT 310.930 317.090 312.110 318.270 ;
        RECT 310.930 315.490 312.110 316.670 ;
        RECT 310.930 137.090 312.110 138.270 ;
        RECT 310.930 135.490 312.110 136.670 ;
        RECT 310.930 -26.410 312.110 -25.230 ;
        RECT 310.930 -28.010 312.110 -26.830 ;
        RECT 328.930 1415.090 330.110 1416.270 ;
        RECT 328.930 1413.490 330.110 1414.670 ;
        RECT 328.930 1235.090 330.110 1236.270 ;
        RECT 328.930 1233.490 330.110 1234.670 ;
        RECT 328.930 1055.090 330.110 1056.270 ;
        RECT 328.930 1053.490 330.110 1054.670 ;
        RECT 328.930 875.090 330.110 876.270 ;
        RECT 328.930 873.490 330.110 874.670 ;
        RECT 328.930 695.090 330.110 696.270 ;
        RECT 328.930 693.490 330.110 694.670 ;
        RECT 328.930 515.090 330.110 516.270 ;
        RECT 328.930 513.490 330.110 514.670 ;
        RECT 328.930 335.090 330.110 336.270 ;
        RECT 328.930 333.490 330.110 334.670 ;
        RECT 328.930 155.090 330.110 156.270 ;
        RECT 328.930 153.490 330.110 154.670 ;
        RECT 148.930 -35.810 150.110 -34.630 ;
        RECT 148.930 -37.410 150.110 -36.230 ;
        RECT 454.930 1361.090 456.110 1362.270 ;
        RECT 454.930 1359.490 456.110 1360.670 ;
        RECT 454.930 1181.090 456.110 1182.270 ;
        RECT 454.930 1179.490 456.110 1180.670 ;
        RECT 454.930 1001.090 456.110 1002.270 ;
        RECT 454.930 999.490 456.110 1000.670 ;
        RECT 454.930 821.090 456.110 822.270 ;
        RECT 454.930 819.490 456.110 820.670 ;
        RECT 454.930 641.090 456.110 642.270 ;
        RECT 454.930 639.490 456.110 640.670 ;
        RECT 454.930 461.090 456.110 462.270 ;
        RECT 454.930 459.490 456.110 460.670 ;
        RECT 454.930 281.090 456.110 282.270 ;
        RECT 454.930 279.490 456.110 280.670 ;
        RECT 454.930 101.090 456.110 102.270 ;
        RECT 454.930 99.490 456.110 100.670 ;
        RECT 454.930 -7.610 456.110 -6.430 ;
        RECT 454.930 -9.210 456.110 -8.030 ;
        RECT 472.930 1379.090 474.110 1380.270 ;
        RECT 472.930 1377.490 474.110 1378.670 ;
        RECT 472.930 1199.090 474.110 1200.270 ;
        RECT 472.930 1197.490 474.110 1198.670 ;
        RECT 472.930 1019.090 474.110 1020.270 ;
        RECT 472.930 1017.490 474.110 1018.670 ;
        RECT 472.930 839.090 474.110 840.270 ;
        RECT 472.930 837.490 474.110 838.670 ;
        RECT 472.930 659.090 474.110 660.270 ;
        RECT 472.930 657.490 474.110 658.670 ;
        RECT 472.930 479.090 474.110 480.270 ;
        RECT 472.930 477.490 474.110 478.670 ;
        RECT 472.930 299.090 474.110 300.270 ;
        RECT 472.930 297.490 474.110 298.670 ;
        RECT 472.930 119.090 474.110 120.270 ;
        RECT 472.930 117.490 474.110 118.670 ;
        RECT 472.930 -17.010 474.110 -15.830 ;
        RECT 472.930 -18.610 474.110 -17.430 ;
        RECT 490.930 1397.090 492.110 1398.270 ;
        RECT 490.930 1395.490 492.110 1396.670 ;
        RECT 490.930 1217.090 492.110 1218.270 ;
        RECT 490.930 1215.490 492.110 1216.670 ;
        RECT 490.930 1037.090 492.110 1038.270 ;
        RECT 490.930 1035.490 492.110 1036.670 ;
        RECT 490.930 857.090 492.110 858.270 ;
        RECT 490.930 855.490 492.110 856.670 ;
        RECT 490.930 677.090 492.110 678.270 ;
        RECT 490.930 675.490 492.110 676.670 ;
        RECT 490.930 497.090 492.110 498.270 ;
        RECT 490.930 495.490 492.110 496.670 ;
        RECT 490.930 317.090 492.110 318.270 ;
        RECT 490.930 315.490 492.110 316.670 ;
        RECT 490.930 137.090 492.110 138.270 ;
        RECT 490.930 135.490 492.110 136.670 ;
        RECT 490.930 -26.410 492.110 -25.230 ;
        RECT 490.930 -28.010 492.110 -26.830 ;
        RECT 508.930 1415.090 510.110 1416.270 ;
        RECT 508.930 1413.490 510.110 1414.670 ;
        RECT 508.930 1235.090 510.110 1236.270 ;
        RECT 508.930 1233.490 510.110 1234.670 ;
        RECT 508.930 1055.090 510.110 1056.270 ;
        RECT 508.930 1053.490 510.110 1054.670 ;
        RECT 508.930 875.090 510.110 876.270 ;
        RECT 508.930 873.490 510.110 874.670 ;
        RECT 508.930 695.090 510.110 696.270 ;
        RECT 508.930 693.490 510.110 694.670 ;
        RECT 508.930 515.090 510.110 516.270 ;
        RECT 508.930 513.490 510.110 514.670 ;
        RECT 508.930 335.090 510.110 336.270 ;
        RECT 508.930 333.490 510.110 334.670 ;
        RECT 508.930 155.090 510.110 156.270 ;
        RECT 508.930 153.490 510.110 154.670 ;
        RECT 328.930 -35.810 330.110 -34.630 ;
        RECT 328.930 -37.410 330.110 -36.230 ;
        RECT 634.930 1361.090 636.110 1362.270 ;
        RECT 634.930 1359.490 636.110 1360.670 ;
        RECT 634.930 1181.090 636.110 1182.270 ;
        RECT 634.930 1179.490 636.110 1180.670 ;
        RECT 634.930 1001.090 636.110 1002.270 ;
        RECT 634.930 999.490 636.110 1000.670 ;
        RECT 634.930 821.090 636.110 822.270 ;
        RECT 634.930 819.490 636.110 820.670 ;
        RECT 634.930 641.090 636.110 642.270 ;
        RECT 634.930 639.490 636.110 640.670 ;
        RECT 634.930 461.090 636.110 462.270 ;
        RECT 634.930 459.490 636.110 460.670 ;
        RECT 634.930 281.090 636.110 282.270 ;
        RECT 634.930 279.490 636.110 280.670 ;
        RECT 634.930 101.090 636.110 102.270 ;
        RECT 634.930 99.490 636.110 100.670 ;
        RECT 634.930 -7.610 636.110 -6.430 ;
        RECT 634.930 -9.210 636.110 -8.030 ;
        RECT 652.930 1379.090 654.110 1380.270 ;
        RECT 652.930 1377.490 654.110 1378.670 ;
        RECT 652.930 1199.090 654.110 1200.270 ;
        RECT 652.930 1197.490 654.110 1198.670 ;
        RECT 652.930 1019.090 654.110 1020.270 ;
        RECT 652.930 1017.490 654.110 1018.670 ;
        RECT 652.930 839.090 654.110 840.270 ;
        RECT 652.930 837.490 654.110 838.670 ;
        RECT 652.930 659.090 654.110 660.270 ;
        RECT 652.930 657.490 654.110 658.670 ;
        RECT 652.930 479.090 654.110 480.270 ;
        RECT 652.930 477.490 654.110 478.670 ;
        RECT 652.930 299.090 654.110 300.270 ;
        RECT 652.930 297.490 654.110 298.670 ;
        RECT 652.930 119.090 654.110 120.270 ;
        RECT 652.930 117.490 654.110 118.670 ;
        RECT 652.930 -17.010 654.110 -15.830 ;
        RECT 652.930 -18.610 654.110 -17.430 ;
        RECT 670.930 1397.090 672.110 1398.270 ;
        RECT 670.930 1395.490 672.110 1396.670 ;
        RECT 670.930 1217.090 672.110 1218.270 ;
        RECT 670.930 1215.490 672.110 1216.670 ;
        RECT 670.930 1037.090 672.110 1038.270 ;
        RECT 670.930 1035.490 672.110 1036.670 ;
        RECT 670.930 857.090 672.110 858.270 ;
        RECT 670.930 855.490 672.110 856.670 ;
        RECT 670.930 677.090 672.110 678.270 ;
        RECT 670.930 675.490 672.110 676.670 ;
        RECT 670.930 497.090 672.110 498.270 ;
        RECT 670.930 495.490 672.110 496.670 ;
        RECT 670.930 317.090 672.110 318.270 ;
        RECT 670.930 315.490 672.110 316.670 ;
        RECT 670.930 137.090 672.110 138.270 ;
        RECT 670.930 135.490 672.110 136.670 ;
        RECT 670.930 -26.410 672.110 -25.230 ;
        RECT 670.930 -28.010 672.110 -26.830 ;
        RECT 688.930 1415.090 690.110 1416.270 ;
        RECT 688.930 1413.490 690.110 1414.670 ;
        RECT 688.930 1235.090 690.110 1236.270 ;
        RECT 688.930 1233.490 690.110 1234.670 ;
        RECT 688.930 1055.090 690.110 1056.270 ;
        RECT 688.930 1053.490 690.110 1054.670 ;
        RECT 688.930 875.090 690.110 876.270 ;
        RECT 688.930 873.490 690.110 874.670 ;
        RECT 688.930 695.090 690.110 696.270 ;
        RECT 688.930 693.490 690.110 694.670 ;
        RECT 688.930 515.090 690.110 516.270 ;
        RECT 688.930 513.490 690.110 514.670 ;
        RECT 688.930 335.090 690.110 336.270 ;
        RECT 688.930 333.490 690.110 334.670 ;
        RECT 688.930 155.090 690.110 156.270 ;
        RECT 688.930 153.490 690.110 154.670 ;
        RECT 508.930 -35.810 510.110 -34.630 ;
        RECT 508.930 -37.410 510.110 -36.230 ;
        RECT 814.930 1361.090 816.110 1362.270 ;
        RECT 814.930 1359.490 816.110 1360.670 ;
        RECT 814.930 1181.090 816.110 1182.270 ;
        RECT 814.930 1179.490 816.110 1180.670 ;
        RECT 814.930 1001.090 816.110 1002.270 ;
        RECT 814.930 999.490 816.110 1000.670 ;
        RECT 814.930 821.090 816.110 822.270 ;
        RECT 814.930 819.490 816.110 820.670 ;
        RECT 814.930 641.090 816.110 642.270 ;
        RECT 814.930 639.490 816.110 640.670 ;
        RECT 814.930 461.090 816.110 462.270 ;
        RECT 814.930 459.490 816.110 460.670 ;
        RECT 814.930 281.090 816.110 282.270 ;
        RECT 814.930 279.490 816.110 280.670 ;
        RECT 814.930 101.090 816.110 102.270 ;
        RECT 814.930 99.490 816.110 100.670 ;
        RECT 814.930 -7.610 816.110 -6.430 ;
        RECT 814.930 -9.210 816.110 -8.030 ;
        RECT 832.930 1379.090 834.110 1380.270 ;
        RECT 832.930 1377.490 834.110 1378.670 ;
        RECT 832.930 1199.090 834.110 1200.270 ;
        RECT 832.930 1197.490 834.110 1198.670 ;
        RECT 832.930 1019.090 834.110 1020.270 ;
        RECT 832.930 1017.490 834.110 1018.670 ;
        RECT 832.930 839.090 834.110 840.270 ;
        RECT 832.930 837.490 834.110 838.670 ;
        RECT 832.930 659.090 834.110 660.270 ;
        RECT 832.930 657.490 834.110 658.670 ;
        RECT 832.930 479.090 834.110 480.270 ;
        RECT 832.930 477.490 834.110 478.670 ;
        RECT 832.930 299.090 834.110 300.270 ;
        RECT 832.930 297.490 834.110 298.670 ;
        RECT 832.930 119.090 834.110 120.270 ;
        RECT 832.930 117.490 834.110 118.670 ;
        RECT 832.930 -17.010 834.110 -15.830 ;
        RECT 832.930 -18.610 834.110 -17.430 ;
        RECT 850.930 1397.090 852.110 1398.270 ;
        RECT 850.930 1395.490 852.110 1396.670 ;
        RECT 850.930 1217.090 852.110 1218.270 ;
        RECT 850.930 1215.490 852.110 1216.670 ;
        RECT 850.930 1037.090 852.110 1038.270 ;
        RECT 850.930 1035.490 852.110 1036.670 ;
        RECT 850.930 857.090 852.110 858.270 ;
        RECT 850.930 855.490 852.110 856.670 ;
        RECT 850.930 677.090 852.110 678.270 ;
        RECT 850.930 675.490 852.110 676.670 ;
        RECT 850.930 497.090 852.110 498.270 ;
        RECT 850.930 495.490 852.110 496.670 ;
        RECT 850.930 317.090 852.110 318.270 ;
        RECT 850.930 315.490 852.110 316.670 ;
        RECT 850.930 137.090 852.110 138.270 ;
        RECT 850.930 135.490 852.110 136.670 ;
        RECT 850.930 -26.410 852.110 -25.230 ;
        RECT 850.930 -28.010 852.110 -26.830 ;
        RECT 868.930 1415.090 870.110 1416.270 ;
        RECT 868.930 1413.490 870.110 1414.670 ;
        RECT 868.930 1235.090 870.110 1236.270 ;
        RECT 868.930 1233.490 870.110 1234.670 ;
        RECT 868.930 1055.090 870.110 1056.270 ;
        RECT 868.930 1053.490 870.110 1054.670 ;
        RECT 868.930 875.090 870.110 876.270 ;
        RECT 868.930 873.490 870.110 874.670 ;
        RECT 868.930 695.090 870.110 696.270 ;
        RECT 868.930 693.490 870.110 694.670 ;
        RECT 868.930 515.090 870.110 516.270 ;
        RECT 868.930 513.490 870.110 514.670 ;
        RECT 868.930 335.090 870.110 336.270 ;
        RECT 868.930 333.490 870.110 334.670 ;
        RECT 868.930 155.090 870.110 156.270 ;
        RECT 868.930 153.490 870.110 154.670 ;
        RECT 688.930 -35.810 690.110 -34.630 ;
        RECT 688.930 -37.410 690.110 -36.230 ;
        RECT 994.930 1361.090 996.110 1362.270 ;
        RECT 994.930 1359.490 996.110 1360.670 ;
        RECT 994.930 1181.090 996.110 1182.270 ;
        RECT 994.930 1179.490 996.110 1180.670 ;
        RECT 994.930 1001.090 996.110 1002.270 ;
        RECT 994.930 999.490 996.110 1000.670 ;
        RECT 994.930 821.090 996.110 822.270 ;
        RECT 994.930 819.490 996.110 820.670 ;
        RECT 994.930 641.090 996.110 642.270 ;
        RECT 994.930 639.490 996.110 640.670 ;
        RECT 994.930 461.090 996.110 462.270 ;
        RECT 994.930 459.490 996.110 460.670 ;
        RECT 994.930 281.090 996.110 282.270 ;
        RECT 994.930 279.490 996.110 280.670 ;
        RECT 994.930 101.090 996.110 102.270 ;
        RECT 994.930 99.490 996.110 100.670 ;
        RECT 994.930 -7.610 996.110 -6.430 ;
        RECT 994.930 -9.210 996.110 -8.030 ;
        RECT 1012.930 1379.090 1014.110 1380.270 ;
        RECT 1012.930 1377.490 1014.110 1378.670 ;
        RECT 1012.930 1199.090 1014.110 1200.270 ;
        RECT 1012.930 1197.490 1014.110 1198.670 ;
        RECT 1012.930 1019.090 1014.110 1020.270 ;
        RECT 1012.930 1017.490 1014.110 1018.670 ;
        RECT 1012.930 839.090 1014.110 840.270 ;
        RECT 1012.930 837.490 1014.110 838.670 ;
        RECT 1012.930 659.090 1014.110 660.270 ;
        RECT 1012.930 657.490 1014.110 658.670 ;
        RECT 1012.930 479.090 1014.110 480.270 ;
        RECT 1012.930 477.490 1014.110 478.670 ;
        RECT 1012.930 299.090 1014.110 300.270 ;
        RECT 1012.930 297.490 1014.110 298.670 ;
        RECT 1012.930 119.090 1014.110 120.270 ;
        RECT 1012.930 117.490 1014.110 118.670 ;
        RECT 1012.930 -17.010 1014.110 -15.830 ;
        RECT 1012.930 -18.610 1014.110 -17.430 ;
        RECT 1030.930 1397.090 1032.110 1398.270 ;
        RECT 1030.930 1395.490 1032.110 1396.670 ;
        RECT 1030.930 1217.090 1032.110 1218.270 ;
        RECT 1030.930 1215.490 1032.110 1216.670 ;
        RECT 1030.930 1037.090 1032.110 1038.270 ;
        RECT 1030.930 1035.490 1032.110 1036.670 ;
        RECT 1030.930 857.090 1032.110 858.270 ;
        RECT 1030.930 855.490 1032.110 856.670 ;
        RECT 1030.930 677.090 1032.110 678.270 ;
        RECT 1030.930 675.490 1032.110 676.670 ;
        RECT 1030.930 497.090 1032.110 498.270 ;
        RECT 1030.930 495.490 1032.110 496.670 ;
        RECT 1030.930 317.090 1032.110 318.270 ;
        RECT 1030.930 315.490 1032.110 316.670 ;
        RECT 1030.930 137.090 1032.110 138.270 ;
        RECT 1030.930 135.490 1032.110 136.670 ;
        RECT 1030.930 -26.410 1032.110 -25.230 ;
        RECT 1030.930 -28.010 1032.110 -26.830 ;
        RECT 1048.930 1415.090 1050.110 1416.270 ;
        RECT 1048.930 1413.490 1050.110 1414.670 ;
        RECT 1048.930 1235.090 1050.110 1236.270 ;
        RECT 1048.930 1233.490 1050.110 1234.670 ;
        RECT 1048.930 1055.090 1050.110 1056.270 ;
        RECT 1048.930 1053.490 1050.110 1054.670 ;
        RECT 1048.930 875.090 1050.110 876.270 ;
        RECT 1048.930 873.490 1050.110 874.670 ;
        RECT 1048.930 695.090 1050.110 696.270 ;
        RECT 1048.930 693.490 1050.110 694.670 ;
        RECT 1048.930 515.090 1050.110 516.270 ;
        RECT 1048.930 513.490 1050.110 514.670 ;
        RECT 1048.930 335.090 1050.110 336.270 ;
        RECT 1048.930 333.490 1050.110 334.670 ;
        RECT 1048.930 155.090 1050.110 156.270 ;
        RECT 1048.930 153.490 1050.110 154.670 ;
        RECT 868.930 -35.810 870.110 -34.630 ;
        RECT 868.930 -37.410 870.110 -36.230 ;
        RECT 1174.930 1361.090 1176.110 1362.270 ;
        RECT 1174.930 1359.490 1176.110 1360.670 ;
        RECT 1174.930 1181.090 1176.110 1182.270 ;
        RECT 1174.930 1179.490 1176.110 1180.670 ;
        RECT 1174.930 1001.090 1176.110 1002.270 ;
        RECT 1174.930 999.490 1176.110 1000.670 ;
        RECT 1174.930 821.090 1176.110 822.270 ;
        RECT 1174.930 819.490 1176.110 820.670 ;
        RECT 1174.930 641.090 1176.110 642.270 ;
        RECT 1174.930 639.490 1176.110 640.670 ;
        RECT 1174.930 461.090 1176.110 462.270 ;
        RECT 1174.930 459.490 1176.110 460.670 ;
        RECT 1174.930 281.090 1176.110 282.270 ;
        RECT 1174.930 279.490 1176.110 280.670 ;
        RECT 1174.930 101.090 1176.110 102.270 ;
        RECT 1174.930 99.490 1176.110 100.670 ;
        RECT 1174.930 -7.610 1176.110 -6.430 ;
        RECT 1174.930 -9.210 1176.110 -8.030 ;
        RECT 1192.930 1379.090 1194.110 1380.270 ;
        RECT 1192.930 1377.490 1194.110 1378.670 ;
        RECT 1192.930 1199.090 1194.110 1200.270 ;
        RECT 1192.930 1197.490 1194.110 1198.670 ;
        RECT 1192.930 1019.090 1194.110 1020.270 ;
        RECT 1192.930 1017.490 1194.110 1018.670 ;
        RECT 1192.930 839.090 1194.110 840.270 ;
        RECT 1192.930 837.490 1194.110 838.670 ;
        RECT 1192.930 659.090 1194.110 660.270 ;
        RECT 1192.930 657.490 1194.110 658.670 ;
        RECT 1192.930 479.090 1194.110 480.270 ;
        RECT 1192.930 477.490 1194.110 478.670 ;
        RECT 1192.930 299.090 1194.110 300.270 ;
        RECT 1192.930 297.490 1194.110 298.670 ;
        RECT 1192.930 119.090 1194.110 120.270 ;
        RECT 1192.930 117.490 1194.110 118.670 ;
        RECT 1192.930 -17.010 1194.110 -15.830 ;
        RECT 1192.930 -18.610 1194.110 -17.430 ;
        RECT 1210.930 1397.090 1212.110 1398.270 ;
        RECT 1210.930 1395.490 1212.110 1396.670 ;
        RECT 1210.930 1217.090 1212.110 1218.270 ;
        RECT 1210.930 1215.490 1212.110 1216.670 ;
        RECT 1210.930 1037.090 1212.110 1038.270 ;
        RECT 1210.930 1035.490 1212.110 1036.670 ;
        RECT 1210.930 857.090 1212.110 858.270 ;
        RECT 1210.930 855.490 1212.110 856.670 ;
        RECT 1210.930 677.090 1212.110 678.270 ;
        RECT 1210.930 675.490 1212.110 676.670 ;
        RECT 1210.930 497.090 1212.110 498.270 ;
        RECT 1210.930 495.490 1212.110 496.670 ;
        RECT 1210.930 317.090 1212.110 318.270 ;
        RECT 1210.930 315.490 1212.110 316.670 ;
        RECT 1210.930 137.090 1212.110 138.270 ;
        RECT 1210.930 135.490 1212.110 136.670 ;
        RECT 1210.930 -26.410 1212.110 -25.230 ;
        RECT 1210.930 -28.010 1212.110 -26.830 ;
        RECT 1228.930 1415.090 1230.110 1416.270 ;
        RECT 1228.930 1413.490 1230.110 1414.670 ;
        RECT 1228.930 1235.090 1230.110 1236.270 ;
        RECT 1228.930 1233.490 1230.110 1234.670 ;
        RECT 1228.930 1055.090 1230.110 1056.270 ;
        RECT 1228.930 1053.490 1230.110 1054.670 ;
        RECT 1228.930 875.090 1230.110 876.270 ;
        RECT 1228.930 873.490 1230.110 874.670 ;
        RECT 1228.930 695.090 1230.110 696.270 ;
        RECT 1228.930 693.490 1230.110 694.670 ;
        RECT 1228.930 515.090 1230.110 516.270 ;
        RECT 1228.930 513.490 1230.110 514.670 ;
        RECT 1228.930 335.090 1230.110 336.270 ;
        RECT 1228.930 333.490 1230.110 334.670 ;
        RECT 1228.930 155.090 1230.110 156.270 ;
        RECT 1228.930 153.490 1230.110 154.670 ;
        RECT 1048.930 -35.810 1050.110 -34.630 ;
        RECT 1048.930 -37.410 1050.110 -36.230 ;
        RECT 1354.930 1361.090 1356.110 1362.270 ;
        RECT 1354.930 1359.490 1356.110 1360.670 ;
        RECT 1354.930 1181.090 1356.110 1182.270 ;
        RECT 1354.930 1179.490 1356.110 1180.670 ;
        RECT 1354.930 1001.090 1356.110 1002.270 ;
        RECT 1354.930 999.490 1356.110 1000.670 ;
        RECT 1354.930 821.090 1356.110 822.270 ;
        RECT 1354.930 819.490 1356.110 820.670 ;
        RECT 1354.930 641.090 1356.110 642.270 ;
        RECT 1354.930 639.490 1356.110 640.670 ;
        RECT 1354.930 461.090 1356.110 462.270 ;
        RECT 1354.930 459.490 1356.110 460.670 ;
        RECT 1354.930 281.090 1356.110 282.270 ;
        RECT 1354.930 279.490 1356.110 280.670 ;
        RECT 1354.930 101.090 1356.110 102.270 ;
        RECT 1354.930 99.490 1356.110 100.670 ;
        RECT 1354.930 -7.610 1356.110 -6.430 ;
        RECT 1354.930 -9.210 1356.110 -8.030 ;
        RECT 1372.930 1379.090 1374.110 1380.270 ;
        RECT 1372.930 1377.490 1374.110 1378.670 ;
        RECT 1372.930 1199.090 1374.110 1200.270 ;
        RECT 1372.930 1197.490 1374.110 1198.670 ;
        RECT 1372.930 1019.090 1374.110 1020.270 ;
        RECT 1372.930 1017.490 1374.110 1018.670 ;
        RECT 1372.930 839.090 1374.110 840.270 ;
        RECT 1372.930 837.490 1374.110 838.670 ;
        RECT 1372.930 659.090 1374.110 660.270 ;
        RECT 1372.930 657.490 1374.110 658.670 ;
        RECT 1372.930 479.090 1374.110 480.270 ;
        RECT 1372.930 477.490 1374.110 478.670 ;
        RECT 1372.930 299.090 1374.110 300.270 ;
        RECT 1372.930 297.490 1374.110 298.670 ;
        RECT 1372.930 119.090 1374.110 120.270 ;
        RECT 1372.930 117.490 1374.110 118.670 ;
        RECT 1372.930 -17.010 1374.110 -15.830 ;
        RECT 1372.930 -18.610 1374.110 -17.430 ;
        RECT 1390.930 1397.090 1392.110 1398.270 ;
        RECT 1390.930 1395.490 1392.110 1396.670 ;
        RECT 1390.930 1217.090 1392.110 1218.270 ;
        RECT 1390.930 1215.490 1392.110 1216.670 ;
        RECT 1390.930 1037.090 1392.110 1038.270 ;
        RECT 1390.930 1035.490 1392.110 1036.670 ;
        RECT 1390.930 857.090 1392.110 858.270 ;
        RECT 1390.930 855.490 1392.110 856.670 ;
        RECT 1390.930 677.090 1392.110 678.270 ;
        RECT 1390.930 675.490 1392.110 676.670 ;
        RECT 1390.930 497.090 1392.110 498.270 ;
        RECT 1390.930 495.490 1392.110 496.670 ;
        RECT 1390.930 317.090 1392.110 318.270 ;
        RECT 1390.930 315.490 1392.110 316.670 ;
        RECT 1390.930 137.090 1392.110 138.270 ;
        RECT 1390.930 135.490 1392.110 136.670 ;
        RECT 1390.930 -26.410 1392.110 -25.230 ;
        RECT 1390.930 -28.010 1392.110 -26.830 ;
        RECT 1408.930 1415.090 1410.110 1416.270 ;
        RECT 1408.930 1413.490 1410.110 1414.670 ;
        RECT 1408.930 1235.090 1410.110 1236.270 ;
        RECT 1408.930 1233.490 1410.110 1234.670 ;
        RECT 1408.930 1055.090 1410.110 1056.270 ;
        RECT 1408.930 1053.490 1410.110 1054.670 ;
        RECT 1408.930 875.090 1410.110 876.270 ;
        RECT 1408.930 873.490 1410.110 874.670 ;
        RECT 1408.930 695.090 1410.110 696.270 ;
        RECT 1408.930 693.490 1410.110 694.670 ;
        RECT 1408.930 515.090 1410.110 516.270 ;
        RECT 1408.930 513.490 1410.110 514.670 ;
        RECT 1408.930 335.090 1410.110 336.270 ;
        RECT 1408.930 333.490 1410.110 334.670 ;
        RECT 1408.930 155.090 1410.110 156.270 ;
        RECT 1408.930 153.490 1410.110 154.670 ;
        RECT 1228.930 -35.810 1230.110 -34.630 ;
        RECT 1228.930 -37.410 1230.110 -36.230 ;
        RECT 1534.930 1361.090 1536.110 1362.270 ;
        RECT 1534.930 1359.490 1536.110 1360.670 ;
        RECT 1534.930 1181.090 1536.110 1182.270 ;
        RECT 1534.930 1179.490 1536.110 1180.670 ;
        RECT 1534.930 1001.090 1536.110 1002.270 ;
        RECT 1534.930 999.490 1536.110 1000.670 ;
        RECT 1534.930 821.090 1536.110 822.270 ;
        RECT 1534.930 819.490 1536.110 820.670 ;
        RECT 1534.930 641.090 1536.110 642.270 ;
        RECT 1534.930 639.490 1536.110 640.670 ;
        RECT 1534.930 461.090 1536.110 462.270 ;
        RECT 1534.930 459.490 1536.110 460.670 ;
        RECT 1534.930 281.090 1536.110 282.270 ;
        RECT 1534.930 279.490 1536.110 280.670 ;
        RECT 1534.930 101.090 1536.110 102.270 ;
        RECT 1534.930 99.490 1536.110 100.670 ;
        RECT 1534.930 -7.610 1536.110 -6.430 ;
        RECT 1534.930 -9.210 1536.110 -8.030 ;
        RECT 1552.930 2639.090 1554.110 2640.270 ;
        RECT 1552.930 2637.490 1554.110 2638.670 ;
        RECT 1552.930 2459.090 1554.110 2460.270 ;
        RECT 1552.930 2457.490 1554.110 2458.670 ;
        RECT 1552.930 2279.090 1554.110 2280.270 ;
        RECT 1552.930 2277.490 1554.110 2278.670 ;
        RECT 1552.930 2099.090 1554.110 2100.270 ;
        RECT 1552.930 2097.490 1554.110 2098.670 ;
        RECT 1552.930 1919.090 1554.110 1920.270 ;
        RECT 1552.930 1917.490 1554.110 1918.670 ;
        RECT 1552.930 1739.090 1554.110 1740.270 ;
        RECT 1552.930 1737.490 1554.110 1738.670 ;
        RECT 1552.930 1559.090 1554.110 1560.270 ;
        RECT 1552.930 1557.490 1554.110 1558.670 ;
        RECT 1552.930 1379.090 1554.110 1380.270 ;
        RECT 1552.930 1377.490 1554.110 1378.670 ;
        RECT 1552.930 1199.090 1554.110 1200.270 ;
        RECT 1552.930 1197.490 1554.110 1198.670 ;
        RECT 1552.930 1019.090 1554.110 1020.270 ;
        RECT 1552.930 1017.490 1554.110 1018.670 ;
        RECT 1552.930 839.090 1554.110 840.270 ;
        RECT 1552.930 837.490 1554.110 838.670 ;
        RECT 1552.930 659.090 1554.110 660.270 ;
        RECT 1552.930 657.490 1554.110 658.670 ;
        RECT 1552.930 479.090 1554.110 480.270 ;
        RECT 1552.930 477.490 1554.110 478.670 ;
        RECT 1552.930 299.090 1554.110 300.270 ;
        RECT 1552.930 297.490 1554.110 298.670 ;
        RECT 1552.930 119.090 1554.110 120.270 ;
        RECT 1552.930 117.490 1554.110 118.670 ;
        RECT 1552.930 -17.010 1554.110 -15.830 ;
        RECT 1552.930 -18.610 1554.110 -17.430 ;
        RECT 1570.930 2657.090 1572.110 2658.270 ;
        RECT 1570.930 2655.490 1572.110 2656.670 ;
        RECT 1570.930 2477.090 1572.110 2478.270 ;
        RECT 1570.930 2475.490 1572.110 2476.670 ;
        RECT 1570.930 2297.090 1572.110 2298.270 ;
        RECT 1570.930 2295.490 1572.110 2296.670 ;
        RECT 1570.930 2117.090 1572.110 2118.270 ;
        RECT 1570.930 2115.490 1572.110 2116.670 ;
        RECT 1570.930 1937.090 1572.110 1938.270 ;
        RECT 1570.930 1935.490 1572.110 1936.670 ;
        RECT 1570.930 1757.090 1572.110 1758.270 ;
        RECT 1570.930 1755.490 1572.110 1756.670 ;
        RECT 1570.930 1577.090 1572.110 1578.270 ;
        RECT 1570.930 1575.490 1572.110 1576.670 ;
        RECT 1570.930 1397.090 1572.110 1398.270 ;
        RECT 1570.930 1395.490 1572.110 1396.670 ;
        RECT 1570.930 1217.090 1572.110 1218.270 ;
        RECT 1570.930 1215.490 1572.110 1216.670 ;
        RECT 1570.930 1037.090 1572.110 1038.270 ;
        RECT 1570.930 1035.490 1572.110 1036.670 ;
        RECT 1570.930 857.090 1572.110 858.270 ;
        RECT 1570.930 855.490 1572.110 856.670 ;
        RECT 1570.930 677.090 1572.110 678.270 ;
        RECT 1570.930 675.490 1572.110 676.670 ;
        RECT 1570.930 497.090 1572.110 498.270 ;
        RECT 1570.930 495.490 1572.110 496.670 ;
        RECT 1570.930 317.090 1572.110 318.270 ;
        RECT 1570.930 315.490 1572.110 316.670 ;
        RECT 1570.930 137.090 1572.110 138.270 ;
        RECT 1570.930 135.490 1572.110 136.670 ;
        RECT 1570.930 -26.410 1572.110 -25.230 ;
        RECT 1570.930 -28.010 1572.110 -26.830 ;
        RECT 1588.930 2675.090 1590.110 2676.270 ;
        RECT 1588.930 2673.490 1590.110 2674.670 ;
        RECT 1588.930 2495.090 1590.110 2496.270 ;
        RECT 1588.930 2493.490 1590.110 2494.670 ;
        RECT 1588.930 2315.090 1590.110 2316.270 ;
        RECT 1588.930 2313.490 1590.110 2314.670 ;
        RECT 1588.930 2135.090 1590.110 2136.270 ;
        RECT 1588.930 2133.490 1590.110 2134.670 ;
        RECT 1588.930 1955.090 1590.110 1956.270 ;
        RECT 1588.930 1953.490 1590.110 1954.670 ;
        RECT 1588.930 1775.090 1590.110 1776.270 ;
        RECT 1588.930 1773.490 1590.110 1774.670 ;
        RECT 1588.930 1595.090 1590.110 1596.270 ;
        RECT 1588.930 1593.490 1590.110 1594.670 ;
        RECT 1588.930 1415.090 1590.110 1416.270 ;
        RECT 1588.930 1413.490 1590.110 1414.670 ;
        RECT 1588.930 1235.090 1590.110 1236.270 ;
        RECT 1588.930 1233.490 1590.110 1234.670 ;
        RECT 1588.930 1055.090 1590.110 1056.270 ;
        RECT 1588.930 1053.490 1590.110 1054.670 ;
        RECT 1588.930 875.090 1590.110 876.270 ;
        RECT 1588.930 873.490 1590.110 874.670 ;
        RECT 1588.930 695.090 1590.110 696.270 ;
        RECT 1588.930 693.490 1590.110 694.670 ;
        RECT 1588.930 515.090 1590.110 516.270 ;
        RECT 1588.930 513.490 1590.110 514.670 ;
        RECT 1588.930 335.090 1590.110 336.270 ;
        RECT 1588.930 333.490 1590.110 334.670 ;
        RECT 1588.930 155.090 1590.110 156.270 ;
        RECT 1588.930 153.490 1590.110 154.670 ;
        RECT 1408.930 -35.810 1410.110 -34.630 ;
        RECT 1408.930 -37.410 1410.110 -36.230 ;
        RECT 1714.930 2621.090 1716.110 2622.270 ;
        RECT 1714.930 2619.490 1716.110 2620.670 ;
        RECT 1714.930 2441.090 1716.110 2442.270 ;
        RECT 1714.930 2439.490 1716.110 2440.670 ;
        RECT 1714.930 2261.090 1716.110 2262.270 ;
        RECT 1714.930 2259.490 1716.110 2260.670 ;
        RECT 1714.930 2081.090 1716.110 2082.270 ;
        RECT 1714.930 2079.490 1716.110 2080.670 ;
        RECT 1714.930 1901.090 1716.110 1902.270 ;
        RECT 1714.930 1899.490 1716.110 1900.670 ;
        RECT 1714.930 1721.090 1716.110 1722.270 ;
        RECT 1714.930 1719.490 1716.110 1720.670 ;
        RECT 1714.930 1541.090 1716.110 1542.270 ;
        RECT 1714.930 1539.490 1716.110 1540.670 ;
        RECT 1714.930 1361.090 1716.110 1362.270 ;
        RECT 1714.930 1359.490 1716.110 1360.670 ;
        RECT 1714.930 1181.090 1716.110 1182.270 ;
        RECT 1714.930 1179.490 1716.110 1180.670 ;
        RECT 1714.930 1001.090 1716.110 1002.270 ;
        RECT 1714.930 999.490 1716.110 1000.670 ;
        RECT 1714.930 821.090 1716.110 822.270 ;
        RECT 1714.930 819.490 1716.110 820.670 ;
        RECT 1714.930 641.090 1716.110 642.270 ;
        RECT 1714.930 639.490 1716.110 640.670 ;
        RECT 1714.930 461.090 1716.110 462.270 ;
        RECT 1714.930 459.490 1716.110 460.670 ;
        RECT 1714.930 281.090 1716.110 282.270 ;
        RECT 1714.930 279.490 1716.110 280.670 ;
        RECT 1714.930 101.090 1716.110 102.270 ;
        RECT 1714.930 99.490 1716.110 100.670 ;
        RECT 1714.930 -7.610 1716.110 -6.430 ;
        RECT 1714.930 -9.210 1716.110 -8.030 ;
        RECT 1732.930 2639.090 1734.110 2640.270 ;
        RECT 1732.930 2637.490 1734.110 2638.670 ;
        RECT 1732.930 2459.090 1734.110 2460.270 ;
        RECT 1732.930 2457.490 1734.110 2458.670 ;
        RECT 1732.930 2279.090 1734.110 2280.270 ;
        RECT 1732.930 2277.490 1734.110 2278.670 ;
        RECT 1732.930 2099.090 1734.110 2100.270 ;
        RECT 1732.930 2097.490 1734.110 2098.670 ;
        RECT 1732.930 1919.090 1734.110 1920.270 ;
        RECT 1732.930 1917.490 1734.110 1918.670 ;
        RECT 1732.930 1739.090 1734.110 1740.270 ;
        RECT 1732.930 1737.490 1734.110 1738.670 ;
        RECT 1732.930 1559.090 1734.110 1560.270 ;
        RECT 1732.930 1557.490 1734.110 1558.670 ;
        RECT 1732.930 1379.090 1734.110 1380.270 ;
        RECT 1732.930 1377.490 1734.110 1378.670 ;
        RECT 1732.930 1199.090 1734.110 1200.270 ;
        RECT 1732.930 1197.490 1734.110 1198.670 ;
        RECT 1732.930 1019.090 1734.110 1020.270 ;
        RECT 1732.930 1017.490 1734.110 1018.670 ;
        RECT 1732.930 839.090 1734.110 840.270 ;
        RECT 1732.930 837.490 1734.110 838.670 ;
        RECT 1732.930 659.090 1734.110 660.270 ;
        RECT 1732.930 657.490 1734.110 658.670 ;
        RECT 1732.930 479.090 1734.110 480.270 ;
        RECT 1732.930 477.490 1734.110 478.670 ;
        RECT 1732.930 299.090 1734.110 300.270 ;
        RECT 1732.930 297.490 1734.110 298.670 ;
        RECT 1732.930 119.090 1734.110 120.270 ;
        RECT 1732.930 117.490 1734.110 118.670 ;
        RECT 1732.930 -17.010 1734.110 -15.830 ;
        RECT 1732.930 -18.610 1734.110 -17.430 ;
        RECT 1750.930 2657.090 1752.110 2658.270 ;
        RECT 1750.930 2655.490 1752.110 2656.670 ;
        RECT 1750.930 2477.090 1752.110 2478.270 ;
        RECT 1750.930 2475.490 1752.110 2476.670 ;
        RECT 1750.930 2297.090 1752.110 2298.270 ;
        RECT 1750.930 2295.490 1752.110 2296.670 ;
        RECT 1750.930 2117.090 1752.110 2118.270 ;
        RECT 1750.930 2115.490 1752.110 2116.670 ;
        RECT 1750.930 1937.090 1752.110 1938.270 ;
        RECT 1750.930 1935.490 1752.110 1936.670 ;
        RECT 1750.930 1757.090 1752.110 1758.270 ;
        RECT 1750.930 1755.490 1752.110 1756.670 ;
        RECT 1750.930 1577.090 1752.110 1578.270 ;
        RECT 1750.930 1575.490 1752.110 1576.670 ;
        RECT 1750.930 1397.090 1752.110 1398.270 ;
        RECT 1750.930 1395.490 1752.110 1396.670 ;
        RECT 1750.930 1217.090 1752.110 1218.270 ;
        RECT 1750.930 1215.490 1752.110 1216.670 ;
        RECT 1750.930 1037.090 1752.110 1038.270 ;
        RECT 1750.930 1035.490 1752.110 1036.670 ;
        RECT 1750.930 857.090 1752.110 858.270 ;
        RECT 1750.930 855.490 1752.110 856.670 ;
        RECT 1750.930 677.090 1752.110 678.270 ;
        RECT 1750.930 675.490 1752.110 676.670 ;
        RECT 1750.930 497.090 1752.110 498.270 ;
        RECT 1750.930 495.490 1752.110 496.670 ;
        RECT 1750.930 317.090 1752.110 318.270 ;
        RECT 1750.930 315.490 1752.110 316.670 ;
        RECT 1750.930 137.090 1752.110 138.270 ;
        RECT 1750.930 135.490 1752.110 136.670 ;
        RECT 1750.930 -26.410 1752.110 -25.230 ;
        RECT 1750.930 -28.010 1752.110 -26.830 ;
        RECT 1768.930 2675.090 1770.110 2676.270 ;
        RECT 1768.930 2673.490 1770.110 2674.670 ;
        RECT 1768.930 2495.090 1770.110 2496.270 ;
        RECT 1768.930 2493.490 1770.110 2494.670 ;
        RECT 1768.930 2315.090 1770.110 2316.270 ;
        RECT 1768.930 2313.490 1770.110 2314.670 ;
        RECT 1768.930 2135.090 1770.110 2136.270 ;
        RECT 1768.930 2133.490 1770.110 2134.670 ;
        RECT 1768.930 1955.090 1770.110 1956.270 ;
        RECT 1768.930 1953.490 1770.110 1954.670 ;
        RECT 1768.930 1775.090 1770.110 1776.270 ;
        RECT 1768.930 1773.490 1770.110 1774.670 ;
        RECT 1768.930 1595.090 1770.110 1596.270 ;
        RECT 1768.930 1593.490 1770.110 1594.670 ;
        RECT 1768.930 1415.090 1770.110 1416.270 ;
        RECT 1768.930 1413.490 1770.110 1414.670 ;
        RECT 1768.930 1235.090 1770.110 1236.270 ;
        RECT 1768.930 1233.490 1770.110 1234.670 ;
        RECT 1768.930 1055.090 1770.110 1056.270 ;
        RECT 1768.930 1053.490 1770.110 1054.670 ;
        RECT 1768.930 875.090 1770.110 876.270 ;
        RECT 1768.930 873.490 1770.110 874.670 ;
        RECT 1768.930 695.090 1770.110 696.270 ;
        RECT 1768.930 693.490 1770.110 694.670 ;
        RECT 1768.930 515.090 1770.110 516.270 ;
        RECT 1768.930 513.490 1770.110 514.670 ;
        RECT 1768.930 335.090 1770.110 336.270 ;
        RECT 1768.930 333.490 1770.110 334.670 ;
        RECT 1768.930 155.090 1770.110 156.270 ;
        RECT 1768.930 153.490 1770.110 154.670 ;
        RECT 1588.930 -35.810 1590.110 -34.630 ;
        RECT 1588.930 -37.410 1590.110 -36.230 ;
        RECT 1894.930 2621.090 1896.110 2622.270 ;
        RECT 1894.930 2619.490 1896.110 2620.670 ;
        RECT 1894.930 2441.090 1896.110 2442.270 ;
        RECT 1894.930 2439.490 1896.110 2440.670 ;
        RECT 1894.930 2261.090 1896.110 2262.270 ;
        RECT 1894.930 2259.490 1896.110 2260.670 ;
        RECT 1894.930 2081.090 1896.110 2082.270 ;
        RECT 1894.930 2079.490 1896.110 2080.670 ;
        RECT 1894.930 1901.090 1896.110 1902.270 ;
        RECT 1894.930 1899.490 1896.110 1900.670 ;
        RECT 1894.930 1721.090 1896.110 1722.270 ;
        RECT 1894.930 1719.490 1896.110 1720.670 ;
        RECT 1894.930 1541.090 1896.110 1542.270 ;
        RECT 1894.930 1539.490 1896.110 1540.670 ;
        RECT 1894.930 1361.090 1896.110 1362.270 ;
        RECT 1894.930 1359.490 1896.110 1360.670 ;
        RECT 1894.930 1181.090 1896.110 1182.270 ;
        RECT 1894.930 1179.490 1896.110 1180.670 ;
        RECT 1894.930 1001.090 1896.110 1002.270 ;
        RECT 1894.930 999.490 1896.110 1000.670 ;
        RECT 1894.930 821.090 1896.110 822.270 ;
        RECT 1894.930 819.490 1896.110 820.670 ;
        RECT 1894.930 641.090 1896.110 642.270 ;
        RECT 1894.930 639.490 1896.110 640.670 ;
        RECT 1894.930 461.090 1896.110 462.270 ;
        RECT 1894.930 459.490 1896.110 460.670 ;
        RECT 1894.930 281.090 1896.110 282.270 ;
        RECT 1894.930 279.490 1896.110 280.670 ;
        RECT 1894.930 101.090 1896.110 102.270 ;
        RECT 1894.930 99.490 1896.110 100.670 ;
        RECT 1894.930 -7.610 1896.110 -6.430 ;
        RECT 1894.930 -9.210 1896.110 -8.030 ;
        RECT 1912.930 2639.090 1914.110 2640.270 ;
        RECT 1912.930 2637.490 1914.110 2638.670 ;
        RECT 1912.930 2459.090 1914.110 2460.270 ;
        RECT 1912.930 2457.490 1914.110 2458.670 ;
        RECT 1912.930 2279.090 1914.110 2280.270 ;
        RECT 1912.930 2277.490 1914.110 2278.670 ;
        RECT 1912.930 2099.090 1914.110 2100.270 ;
        RECT 1912.930 2097.490 1914.110 2098.670 ;
        RECT 1912.930 1919.090 1914.110 1920.270 ;
        RECT 1912.930 1917.490 1914.110 1918.670 ;
        RECT 1912.930 1739.090 1914.110 1740.270 ;
        RECT 1912.930 1737.490 1914.110 1738.670 ;
        RECT 1912.930 1559.090 1914.110 1560.270 ;
        RECT 1912.930 1557.490 1914.110 1558.670 ;
        RECT 1912.930 1379.090 1914.110 1380.270 ;
        RECT 1912.930 1377.490 1914.110 1378.670 ;
        RECT 1912.930 1199.090 1914.110 1200.270 ;
        RECT 1912.930 1197.490 1914.110 1198.670 ;
        RECT 1912.930 1019.090 1914.110 1020.270 ;
        RECT 1912.930 1017.490 1914.110 1018.670 ;
        RECT 1912.930 839.090 1914.110 840.270 ;
        RECT 1912.930 837.490 1914.110 838.670 ;
        RECT 1912.930 659.090 1914.110 660.270 ;
        RECT 1912.930 657.490 1914.110 658.670 ;
        RECT 1912.930 479.090 1914.110 480.270 ;
        RECT 1912.930 477.490 1914.110 478.670 ;
        RECT 1912.930 299.090 1914.110 300.270 ;
        RECT 1912.930 297.490 1914.110 298.670 ;
        RECT 1912.930 119.090 1914.110 120.270 ;
        RECT 1912.930 117.490 1914.110 118.670 ;
        RECT 1912.930 -17.010 1914.110 -15.830 ;
        RECT 1912.930 -18.610 1914.110 -17.430 ;
        RECT 1930.930 2657.090 1932.110 2658.270 ;
        RECT 1930.930 2655.490 1932.110 2656.670 ;
        RECT 1930.930 2477.090 1932.110 2478.270 ;
        RECT 1930.930 2475.490 1932.110 2476.670 ;
        RECT 1930.930 2297.090 1932.110 2298.270 ;
        RECT 1930.930 2295.490 1932.110 2296.670 ;
        RECT 1930.930 2117.090 1932.110 2118.270 ;
        RECT 1930.930 2115.490 1932.110 2116.670 ;
        RECT 1930.930 1937.090 1932.110 1938.270 ;
        RECT 1930.930 1935.490 1932.110 1936.670 ;
        RECT 1930.930 1757.090 1932.110 1758.270 ;
        RECT 1930.930 1755.490 1932.110 1756.670 ;
        RECT 1930.930 1577.090 1932.110 1578.270 ;
        RECT 1930.930 1575.490 1932.110 1576.670 ;
        RECT 1930.930 1397.090 1932.110 1398.270 ;
        RECT 1930.930 1395.490 1932.110 1396.670 ;
        RECT 1930.930 1217.090 1932.110 1218.270 ;
        RECT 1930.930 1215.490 1932.110 1216.670 ;
        RECT 1930.930 1037.090 1932.110 1038.270 ;
        RECT 1930.930 1035.490 1932.110 1036.670 ;
        RECT 1930.930 857.090 1932.110 858.270 ;
        RECT 1930.930 855.490 1932.110 856.670 ;
        RECT 1930.930 677.090 1932.110 678.270 ;
        RECT 1930.930 675.490 1932.110 676.670 ;
        RECT 1930.930 497.090 1932.110 498.270 ;
        RECT 1930.930 495.490 1932.110 496.670 ;
        RECT 1930.930 317.090 1932.110 318.270 ;
        RECT 1930.930 315.490 1932.110 316.670 ;
        RECT 1930.930 137.090 1932.110 138.270 ;
        RECT 1930.930 135.490 1932.110 136.670 ;
        RECT 1930.930 -26.410 1932.110 -25.230 ;
        RECT 1930.930 -28.010 1932.110 -26.830 ;
        RECT 1948.930 2675.090 1950.110 2676.270 ;
        RECT 1948.930 2673.490 1950.110 2674.670 ;
        RECT 1948.930 2495.090 1950.110 2496.270 ;
        RECT 1948.930 2493.490 1950.110 2494.670 ;
        RECT 1948.930 2315.090 1950.110 2316.270 ;
        RECT 1948.930 2313.490 1950.110 2314.670 ;
        RECT 1948.930 2135.090 1950.110 2136.270 ;
        RECT 1948.930 2133.490 1950.110 2134.670 ;
        RECT 1948.930 1955.090 1950.110 1956.270 ;
        RECT 1948.930 1953.490 1950.110 1954.670 ;
        RECT 1948.930 1775.090 1950.110 1776.270 ;
        RECT 1948.930 1773.490 1950.110 1774.670 ;
        RECT 1948.930 1595.090 1950.110 1596.270 ;
        RECT 1948.930 1593.490 1950.110 1594.670 ;
        RECT 1948.930 1415.090 1950.110 1416.270 ;
        RECT 1948.930 1413.490 1950.110 1414.670 ;
        RECT 1948.930 1235.090 1950.110 1236.270 ;
        RECT 1948.930 1233.490 1950.110 1234.670 ;
        RECT 1948.930 1055.090 1950.110 1056.270 ;
        RECT 1948.930 1053.490 1950.110 1054.670 ;
        RECT 1948.930 875.090 1950.110 876.270 ;
        RECT 1948.930 873.490 1950.110 874.670 ;
        RECT 1948.930 695.090 1950.110 696.270 ;
        RECT 1948.930 693.490 1950.110 694.670 ;
        RECT 1948.930 515.090 1950.110 516.270 ;
        RECT 1948.930 513.490 1950.110 514.670 ;
        RECT 1948.930 335.090 1950.110 336.270 ;
        RECT 1948.930 333.490 1950.110 334.670 ;
        RECT 1948.930 155.090 1950.110 156.270 ;
        RECT 1948.930 153.490 1950.110 154.670 ;
        RECT 1768.930 -35.810 1770.110 -34.630 ;
        RECT 1768.930 -37.410 1770.110 -36.230 ;
        RECT 2074.930 2621.090 2076.110 2622.270 ;
        RECT 2074.930 2619.490 2076.110 2620.670 ;
        RECT 2074.930 2441.090 2076.110 2442.270 ;
        RECT 2074.930 2439.490 2076.110 2440.670 ;
        RECT 2074.930 2261.090 2076.110 2262.270 ;
        RECT 2074.930 2259.490 2076.110 2260.670 ;
        RECT 2074.930 2081.090 2076.110 2082.270 ;
        RECT 2074.930 2079.490 2076.110 2080.670 ;
        RECT 2074.930 1901.090 2076.110 1902.270 ;
        RECT 2074.930 1899.490 2076.110 1900.670 ;
        RECT 2074.930 1721.090 2076.110 1722.270 ;
        RECT 2074.930 1719.490 2076.110 1720.670 ;
        RECT 2074.930 1541.090 2076.110 1542.270 ;
        RECT 2074.930 1539.490 2076.110 1540.670 ;
        RECT 2074.930 1361.090 2076.110 1362.270 ;
        RECT 2074.930 1359.490 2076.110 1360.670 ;
        RECT 2074.930 1181.090 2076.110 1182.270 ;
        RECT 2074.930 1179.490 2076.110 1180.670 ;
        RECT 2074.930 1001.090 2076.110 1002.270 ;
        RECT 2074.930 999.490 2076.110 1000.670 ;
        RECT 2074.930 821.090 2076.110 822.270 ;
        RECT 2074.930 819.490 2076.110 820.670 ;
        RECT 2074.930 641.090 2076.110 642.270 ;
        RECT 2074.930 639.490 2076.110 640.670 ;
        RECT 2074.930 461.090 2076.110 462.270 ;
        RECT 2074.930 459.490 2076.110 460.670 ;
        RECT 2074.930 281.090 2076.110 282.270 ;
        RECT 2074.930 279.490 2076.110 280.670 ;
        RECT 2074.930 101.090 2076.110 102.270 ;
        RECT 2074.930 99.490 2076.110 100.670 ;
        RECT 2074.930 -7.610 2076.110 -6.430 ;
        RECT 2074.930 -9.210 2076.110 -8.030 ;
        RECT 2092.930 3359.090 2094.110 3360.270 ;
        RECT 2092.930 3357.490 2094.110 3358.670 ;
        RECT 2092.930 3179.090 2094.110 3180.270 ;
        RECT 2092.930 3177.490 2094.110 3178.670 ;
        RECT 2092.930 2999.090 2094.110 3000.270 ;
        RECT 2092.930 2997.490 2094.110 2998.670 ;
        RECT 2092.930 2819.090 2094.110 2820.270 ;
        RECT 2092.930 2817.490 2094.110 2818.670 ;
        RECT 2092.930 2639.090 2094.110 2640.270 ;
        RECT 2092.930 2637.490 2094.110 2638.670 ;
        RECT 2092.930 2459.090 2094.110 2460.270 ;
        RECT 2092.930 2457.490 2094.110 2458.670 ;
        RECT 2092.930 2279.090 2094.110 2280.270 ;
        RECT 2092.930 2277.490 2094.110 2278.670 ;
        RECT 2092.930 2099.090 2094.110 2100.270 ;
        RECT 2092.930 2097.490 2094.110 2098.670 ;
        RECT 2092.930 1919.090 2094.110 1920.270 ;
        RECT 2092.930 1917.490 2094.110 1918.670 ;
        RECT 2092.930 1739.090 2094.110 1740.270 ;
        RECT 2092.930 1737.490 2094.110 1738.670 ;
        RECT 2092.930 1559.090 2094.110 1560.270 ;
        RECT 2092.930 1557.490 2094.110 1558.670 ;
        RECT 2092.930 1379.090 2094.110 1380.270 ;
        RECT 2092.930 1377.490 2094.110 1378.670 ;
        RECT 2092.930 1199.090 2094.110 1200.270 ;
        RECT 2092.930 1197.490 2094.110 1198.670 ;
        RECT 2092.930 1019.090 2094.110 1020.270 ;
        RECT 2092.930 1017.490 2094.110 1018.670 ;
        RECT 2092.930 839.090 2094.110 840.270 ;
        RECT 2092.930 837.490 2094.110 838.670 ;
        RECT 2092.930 659.090 2094.110 660.270 ;
        RECT 2092.930 657.490 2094.110 658.670 ;
        RECT 2092.930 479.090 2094.110 480.270 ;
        RECT 2092.930 477.490 2094.110 478.670 ;
        RECT 2092.930 299.090 2094.110 300.270 ;
        RECT 2092.930 297.490 2094.110 298.670 ;
        RECT 2092.930 119.090 2094.110 120.270 ;
        RECT 2092.930 117.490 2094.110 118.670 ;
        RECT 2092.930 -17.010 2094.110 -15.830 ;
        RECT 2092.930 -18.610 2094.110 -17.430 ;
        RECT 2110.930 3377.090 2112.110 3378.270 ;
        RECT 2110.930 3375.490 2112.110 3376.670 ;
        RECT 2110.930 3197.090 2112.110 3198.270 ;
        RECT 2110.930 3195.490 2112.110 3196.670 ;
        RECT 2110.930 3017.090 2112.110 3018.270 ;
        RECT 2110.930 3015.490 2112.110 3016.670 ;
        RECT 2110.930 2837.090 2112.110 2838.270 ;
        RECT 2110.930 2835.490 2112.110 2836.670 ;
        RECT 2110.930 2657.090 2112.110 2658.270 ;
        RECT 2110.930 2655.490 2112.110 2656.670 ;
        RECT 2110.930 2477.090 2112.110 2478.270 ;
        RECT 2110.930 2475.490 2112.110 2476.670 ;
        RECT 2110.930 2297.090 2112.110 2298.270 ;
        RECT 2110.930 2295.490 2112.110 2296.670 ;
        RECT 2110.930 2117.090 2112.110 2118.270 ;
        RECT 2110.930 2115.490 2112.110 2116.670 ;
        RECT 2110.930 1937.090 2112.110 1938.270 ;
        RECT 2110.930 1935.490 2112.110 1936.670 ;
        RECT 2110.930 1757.090 2112.110 1758.270 ;
        RECT 2110.930 1755.490 2112.110 1756.670 ;
        RECT 2110.930 1577.090 2112.110 1578.270 ;
        RECT 2110.930 1575.490 2112.110 1576.670 ;
        RECT 2110.930 1397.090 2112.110 1398.270 ;
        RECT 2110.930 1395.490 2112.110 1396.670 ;
        RECT 2110.930 1217.090 2112.110 1218.270 ;
        RECT 2110.930 1215.490 2112.110 1216.670 ;
        RECT 2110.930 1037.090 2112.110 1038.270 ;
        RECT 2110.930 1035.490 2112.110 1036.670 ;
        RECT 2110.930 857.090 2112.110 858.270 ;
        RECT 2110.930 855.490 2112.110 856.670 ;
        RECT 2110.930 677.090 2112.110 678.270 ;
        RECT 2110.930 675.490 2112.110 676.670 ;
        RECT 2110.930 497.090 2112.110 498.270 ;
        RECT 2110.930 495.490 2112.110 496.670 ;
        RECT 2110.930 317.090 2112.110 318.270 ;
        RECT 2110.930 315.490 2112.110 316.670 ;
        RECT 2110.930 137.090 2112.110 138.270 ;
        RECT 2110.930 135.490 2112.110 136.670 ;
        RECT 2110.930 -26.410 2112.110 -25.230 ;
        RECT 2110.930 -28.010 2112.110 -26.830 ;
        RECT 2308.930 3555.910 2310.110 3557.090 ;
        RECT 2308.930 3554.310 2310.110 3555.490 ;
        RECT 2290.930 3546.510 2292.110 3547.690 ;
        RECT 2290.930 3544.910 2292.110 3546.090 ;
        RECT 2272.930 3537.110 2274.110 3538.290 ;
        RECT 2272.930 3535.510 2274.110 3536.690 ;
        RECT 2128.930 3395.090 2130.110 3396.270 ;
        RECT 2128.930 3393.490 2130.110 3394.670 ;
        RECT 2254.930 3527.710 2256.110 3528.890 ;
        RECT 2254.930 3526.110 2256.110 3527.290 ;
        RECT 2254.930 3341.090 2256.110 3342.270 ;
        RECT 2254.930 3339.490 2256.110 3340.670 ;
        RECT 2272.930 3359.090 2274.110 3360.270 ;
        RECT 2272.930 3357.490 2274.110 3358.670 ;
        RECT 2290.930 3377.090 2292.110 3378.270 ;
        RECT 2290.930 3375.490 2292.110 3376.670 ;
        RECT 2488.930 3555.910 2490.110 3557.090 ;
        RECT 2488.930 3554.310 2490.110 3555.490 ;
        RECT 2470.930 3546.510 2472.110 3547.690 ;
        RECT 2470.930 3544.910 2472.110 3546.090 ;
        RECT 2452.930 3537.110 2454.110 3538.290 ;
        RECT 2452.930 3535.510 2454.110 3536.690 ;
        RECT 2308.930 3395.090 2310.110 3396.270 ;
        RECT 2308.930 3393.490 2310.110 3394.670 ;
        RECT 2434.930 3527.710 2436.110 3528.890 ;
        RECT 2434.930 3526.110 2436.110 3527.290 ;
        RECT 2434.930 3341.090 2436.110 3342.270 ;
        RECT 2434.930 3339.490 2436.110 3340.670 ;
        RECT 2452.930 3359.090 2454.110 3360.270 ;
        RECT 2452.930 3357.490 2454.110 3358.670 ;
        RECT 2470.930 3377.090 2472.110 3378.270 ;
        RECT 2470.930 3375.490 2472.110 3376.670 ;
        RECT 2668.930 3555.910 2670.110 3557.090 ;
        RECT 2668.930 3554.310 2670.110 3555.490 ;
        RECT 2650.930 3546.510 2652.110 3547.690 ;
        RECT 2650.930 3544.910 2652.110 3546.090 ;
        RECT 2632.930 3537.110 2634.110 3538.290 ;
        RECT 2632.930 3535.510 2634.110 3536.690 ;
        RECT 2488.930 3395.090 2490.110 3396.270 ;
        RECT 2488.930 3393.490 2490.110 3394.670 ;
        RECT 2614.930 3527.710 2616.110 3528.890 ;
        RECT 2614.930 3526.110 2616.110 3527.290 ;
        RECT 2614.930 3341.090 2616.110 3342.270 ;
        RECT 2614.930 3339.490 2616.110 3340.670 ;
        RECT 2128.930 3215.090 2130.110 3216.270 ;
        RECT 2128.930 3213.490 2130.110 3214.670 ;
        RECT 2128.930 3035.090 2130.110 3036.270 ;
        RECT 2128.930 3033.490 2130.110 3034.670 ;
        RECT 2128.930 2855.090 2130.110 2856.270 ;
        RECT 2128.930 2853.490 2130.110 2854.670 ;
        RECT 2584.910 3215.090 2586.090 3216.270 ;
        RECT 2584.910 3213.490 2586.090 3214.670 ;
        RECT 2584.910 3197.090 2586.090 3198.270 ;
        RECT 2584.910 3195.490 2586.090 3196.670 ;
        RECT 2584.910 3179.090 2586.090 3180.270 ;
        RECT 2584.910 3177.490 2586.090 3178.670 ;
        RECT 2584.910 3161.090 2586.090 3162.270 ;
        RECT 2584.910 3159.490 2586.090 3160.670 ;
        RECT 2584.910 3035.090 2586.090 3036.270 ;
        RECT 2584.910 3033.490 2586.090 3034.670 ;
        RECT 2584.910 3017.090 2586.090 3018.270 ;
        RECT 2584.910 3015.490 2586.090 3016.670 ;
        RECT 2584.910 2999.090 2586.090 3000.270 ;
        RECT 2584.910 2997.490 2586.090 2998.670 ;
        RECT 2584.910 2981.090 2586.090 2982.270 ;
        RECT 2584.910 2979.490 2586.090 2980.670 ;
        RECT 2584.910 2855.090 2586.090 2856.270 ;
        RECT 2584.910 2853.490 2586.090 2854.670 ;
        RECT 2584.910 2837.090 2586.090 2838.270 ;
        RECT 2584.910 2835.490 2586.090 2836.670 ;
        RECT 2584.910 2819.090 2586.090 2820.270 ;
        RECT 2584.910 2817.490 2586.090 2818.670 ;
        RECT 2614.930 3161.090 2616.110 3162.270 ;
        RECT 2614.930 3159.490 2616.110 3160.670 ;
        RECT 2614.930 2981.090 2616.110 2982.270 ;
        RECT 2614.930 2979.490 2616.110 2980.670 ;
        RECT 2614.930 2801.090 2616.110 2802.270 ;
        RECT 2614.930 2799.490 2616.110 2800.670 ;
        RECT 2128.930 2675.090 2130.110 2676.270 ;
        RECT 2128.930 2673.490 2130.110 2674.670 ;
        RECT 2128.930 2495.090 2130.110 2496.270 ;
        RECT 2128.930 2493.490 2130.110 2494.670 ;
        RECT 2128.930 2315.090 2130.110 2316.270 ;
        RECT 2128.930 2313.490 2130.110 2314.670 ;
        RECT 2128.930 2135.090 2130.110 2136.270 ;
        RECT 2128.930 2133.490 2130.110 2134.670 ;
        RECT 2128.930 1955.090 2130.110 1956.270 ;
        RECT 2128.930 1953.490 2130.110 1954.670 ;
        RECT 2128.930 1775.090 2130.110 1776.270 ;
        RECT 2128.930 1773.490 2130.110 1774.670 ;
        RECT 2128.930 1595.090 2130.110 1596.270 ;
        RECT 2128.930 1593.490 2130.110 1594.670 ;
        RECT 2128.930 1415.090 2130.110 1416.270 ;
        RECT 2128.930 1413.490 2130.110 1414.670 ;
        RECT 2128.930 1235.090 2130.110 1236.270 ;
        RECT 2128.930 1233.490 2130.110 1234.670 ;
        RECT 2128.930 1055.090 2130.110 1056.270 ;
        RECT 2128.930 1053.490 2130.110 1054.670 ;
        RECT 2128.930 875.090 2130.110 876.270 ;
        RECT 2128.930 873.490 2130.110 874.670 ;
        RECT 2128.930 695.090 2130.110 696.270 ;
        RECT 2128.930 693.490 2130.110 694.670 ;
        RECT 2128.930 515.090 2130.110 516.270 ;
        RECT 2128.930 513.490 2130.110 514.670 ;
        RECT 2128.930 335.090 2130.110 336.270 ;
        RECT 2128.930 333.490 2130.110 334.670 ;
        RECT 2128.930 155.090 2130.110 156.270 ;
        RECT 2128.930 153.490 2130.110 154.670 ;
        RECT 1948.930 -35.810 1950.110 -34.630 ;
        RECT 1948.930 -37.410 1950.110 -36.230 ;
        RECT 2254.930 2621.090 2256.110 2622.270 ;
        RECT 2254.930 2619.490 2256.110 2620.670 ;
        RECT 2254.930 2441.090 2256.110 2442.270 ;
        RECT 2254.930 2439.490 2256.110 2440.670 ;
        RECT 2254.930 2261.090 2256.110 2262.270 ;
        RECT 2254.930 2259.490 2256.110 2260.670 ;
        RECT 2254.930 2081.090 2256.110 2082.270 ;
        RECT 2254.930 2079.490 2256.110 2080.670 ;
        RECT 2254.930 1901.090 2256.110 1902.270 ;
        RECT 2254.930 1899.490 2256.110 1900.670 ;
        RECT 2254.930 1721.090 2256.110 1722.270 ;
        RECT 2254.930 1719.490 2256.110 1720.670 ;
        RECT 2254.930 1541.090 2256.110 1542.270 ;
        RECT 2254.930 1539.490 2256.110 1540.670 ;
        RECT 2254.930 1361.090 2256.110 1362.270 ;
        RECT 2254.930 1359.490 2256.110 1360.670 ;
        RECT 2254.930 1181.090 2256.110 1182.270 ;
        RECT 2254.930 1179.490 2256.110 1180.670 ;
        RECT 2254.930 1001.090 2256.110 1002.270 ;
        RECT 2254.930 999.490 2256.110 1000.670 ;
        RECT 2254.930 821.090 2256.110 822.270 ;
        RECT 2254.930 819.490 2256.110 820.670 ;
        RECT 2254.930 641.090 2256.110 642.270 ;
        RECT 2254.930 639.490 2256.110 640.670 ;
        RECT 2254.930 461.090 2256.110 462.270 ;
        RECT 2254.930 459.490 2256.110 460.670 ;
        RECT 2254.930 281.090 2256.110 282.270 ;
        RECT 2254.930 279.490 2256.110 280.670 ;
        RECT 2254.930 101.090 2256.110 102.270 ;
        RECT 2254.930 99.490 2256.110 100.670 ;
        RECT 2254.930 -7.610 2256.110 -6.430 ;
        RECT 2254.930 -9.210 2256.110 -8.030 ;
        RECT 2272.930 2639.090 2274.110 2640.270 ;
        RECT 2272.930 2637.490 2274.110 2638.670 ;
        RECT 2272.930 2459.090 2274.110 2460.270 ;
        RECT 2272.930 2457.490 2274.110 2458.670 ;
        RECT 2272.930 2279.090 2274.110 2280.270 ;
        RECT 2272.930 2277.490 2274.110 2278.670 ;
        RECT 2272.930 2099.090 2274.110 2100.270 ;
        RECT 2272.930 2097.490 2274.110 2098.670 ;
        RECT 2272.930 1919.090 2274.110 1920.270 ;
        RECT 2272.930 1917.490 2274.110 1918.670 ;
        RECT 2272.930 1739.090 2274.110 1740.270 ;
        RECT 2272.930 1737.490 2274.110 1738.670 ;
        RECT 2272.930 1559.090 2274.110 1560.270 ;
        RECT 2272.930 1557.490 2274.110 1558.670 ;
        RECT 2272.930 1379.090 2274.110 1380.270 ;
        RECT 2272.930 1377.490 2274.110 1378.670 ;
        RECT 2272.930 1199.090 2274.110 1200.270 ;
        RECT 2272.930 1197.490 2274.110 1198.670 ;
        RECT 2272.930 1019.090 2274.110 1020.270 ;
        RECT 2272.930 1017.490 2274.110 1018.670 ;
        RECT 2272.930 839.090 2274.110 840.270 ;
        RECT 2272.930 837.490 2274.110 838.670 ;
        RECT 2272.930 659.090 2274.110 660.270 ;
        RECT 2272.930 657.490 2274.110 658.670 ;
        RECT 2272.930 479.090 2274.110 480.270 ;
        RECT 2272.930 477.490 2274.110 478.670 ;
        RECT 2272.930 299.090 2274.110 300.270 ;
        RECT 2272.930 297.490 2274.110 298.670 ;
        RECT 2272.930 119.090 2274.110 120.270 ;
        RECT 2272.930 117.490 2274.110 118.670 ;
        RECT 2272.930 -17.010 2274.110 -15.830 ;
        RECT 2272.930 -18.610 2274.110 -17.430 ;
        RECT 2290.930 2657.090 2292.110 2658.270 ;
        RECT 2290.930 2655.490 2292.110 2656.670 ;
        RECT 2290.930 2477.090 2292.110 2478.270 ;
        RECT 2290.930 2475.490 2292.110 2476.670 ;
        RECT 2290.930 2297.090 2292.110 2298.270 ;
        RECT 2290.930 2295.490 2292.110 2296.670 ;
        RECT 2290.930 2117.090 2292.110 2118.270 ;
        RECT 2290.930 2115.490 2292.110 2116.670 ;
        RECT 2290.930 1937.090 2292.110 1938.270 ;
        RECT 2290.930 1935.490 2292.110 1936.670 ;
        RECT 2290.930 1757.090 2292.110 1758.270 ;
        RECT 2290.930 1755.490 2292.110 1756.670 ;
        RECT 2290.930 1577.090 2292.110 1578.270 ;
        RECT 2290.930 1575.490 2292.110 1576.670 ;
        RECT 2290.930 1397.090 2292.110 1398.270 ;
        RECT 2290.930 1395.490 2292.110 1396.670 ;
        RECT 2290.930 1217.090 2292.110 1218.270 ;
        RECT 2290.930 1215.490 2292.110 1216.670 ;
        RECT 2290.930 1037.090 2292.110 1038.270 ;
        RECT 2290.930 1035.490 2292.110 1036.670 ;
        RECT 2290.930 857.090 2292.110 858.270 ;
        RECT 2290.930 855.490 2292.110 856.670 ;
        RECT 2290.930 677.090 2292.110 678.270 ;
        RECT 2290.930 675.490 2292.110 676.670 ;
        RECT 2290.930 497.090 2292.110 498.270 ;
        RECT 2290.930 495.490 2292.110 496.670 ;
        RECT 2290.930 317.090 2292.110 318.270 ;
        RECT 2290.930 315.490 2292.110 316.670 ;
        RECT 2290.930 137.090 2292.110 138.270 ;
        RECT 2290.930 135.490 2292.110 136.670 ;
        RECT 2290.930 -26.410 2292.110 -25.230 ;
        RECT 2290.930 -28.010 2292.110 -26.830 ;
        RECT 2308.930 2675.090 2310.110 2676.270 ;
        RECT 2308.930 2673.490 2310.110 2674.670 ;
        RECT 2308.930 2495.090 2310.110 2496.270 ;
        RECT 2308.930 2493.490 2310.110 2494.670 ;
        RECT 2308.930 2315.090 2310.110 2316.270 ;
        RECT 2308.930 2313.490 2310.110 2314.670 ;
        RECT 2308.930 2135.090 2310.110 2136.270 ;
        RECT 2308.930 2133.490 2310.110 2134.670 ;
        RECT 2308.930 1955.090 2310.110 1956.270 ;
        RECT 2308.930 1953.490 2310.110 1954.670 ;
        RECT 2308.930 1775.090 2310.110 1776.270 ;
        RECT 2308.930 1773.490 2310.110 1774.670 ;
        RECT 2308.930 1595.090 2310.110 1596.270 ;
        RECT 2308.930 1593.490 2310.110 1594.670 ;
        RECT 2308.930 1415.090 2310.110 1416.270 ;
        RECT 2308.930 1413.490 2310.110 1414.670 ;
        RECT 2308.930 1235.090 2310.110 1236.270 ;
        RECT 2308.930 1233.490 2310.110 1234.670 ;
        RECT 2308.930 1055.090 2310.110 1056.270 ;
        RECT 2308.930 1053.490 2310.110 1054.670 ;
        RECT 2308.930 875.090 2310.110 876.270 ;
        RECT 2308.930 873.490 2310.110 874.670 ;
        RECT 2308.930 695.090 2310.110 696.270 ;
        RECT 2308.930 693.490 2310.110 694.670 ;
        RECT 2308.930 515.090 2310.110 516.270 ;
        RECT 2308.930 513.490 2310.110 514.670 ;
        RECT 2308.930 335.090 2310.110 336.270 ;
        RECT 2308.930 333.490 2310.110 334.670 ;
        RECT 2308.930 155.090 2310.110 156.270 ;
        RECT 2308.930 153.490 2310.110 154.670 ;
        RECT 2128.930 -35.810 2130.110 -34.630 ;
        RECT 2128.930 -37.410 2130.110 -36.230 ;
        RECT 2434.930 2621.090 2436.110 2622.270 ;
        RECT 2434.930 2619.490 2436.110 2620.670 ;
        RECT 2434.930 2441.090 2436.110 2442.270 ;
        RECT 2434.930 2439.490 2436.110 2440.670 ;
        RECT 2434.930 2261.090 2436.110 2262.270 ;
        RECT 2434.930 2259.490 2436.110 2260.670 ;
        RECT 2434.930 2081.090 2436.110 2082.270 ;
        RECT 2434.930 2079.490 2436.110 2080.670 ;
        RECT 2434.930 1901.090 2436.110 1902.270 ;
        RECT 2434.930 1899.490 2436.110 1900.670 ;
        RECT 2434.930 1721.090 2436.110 1722.270 ;
        RECT 2434.930 1719.490 2436.110 1720.670 ;
        RECT 2434.930 1541.090 2436.110 1542.270 ;
        RECT 2434.930 1539.490 2436.110 1540.670 ;
        RECT 2434.930 1361.090 2436.110 1362.270 ;
        RECT 2434.930 1359.490 2436.110 1360.670 ;
        RECT 2434.930 1181.090 2436.110 1182.270 ;
        RECT 2434.930 1179.490 2436.110 1180.670 ;
        RECT 2434.930 1001.090 2436.110 1002.270 ;
        RECT 2434.930 999.490 2436.110 1000.670 ;
        RECT 2434.930 821.090 2436.110 822.270 ;
        RECT 2434.930 819.490 2436.110 820.670 ;
        RECT 2434.930 641.090 2436.110 642.270 ;
        RECT 2434.930 639.490 2436.110 640.670 ;
        RECT 2434.930 461.090 2436.110 462.270 ;
        RECT 2434.930 459.490 2436.110 460.670 ;
        RECT 2434.930 281.090 2436.110 282.270 ;
        RECT 2434.930 279.490 2436.110 280.670 ;
        RECT 2434.930 101.090 2436.110 102.270 ;
        RECT 2434.930 99.490 2436.110 100.670 ;
        RECT 2434.930 -7.610 2436.110 -6.430 ;
        RECT 2434.930 -9.210 2436.110 -8.030 ;
        RECT 2452.930 2639.090 2454.110 2640.270 ;
        RECT 2452.930 2637.490 2454.110 2638.670 ;
        RECT 2452.930 2459.090 2454.110 2460.270 ;
        RECT 2452.930 2457.490 2454.110 2458.670 ;
        RECT 2452.930 2279.090 2454.110 2280.270 ;
        RECT 2452.930 2277.490 2454.110 2278.670 ;
        RECT 2452.930 2099.090 2454.110 2100.270 ;
        RECT 2452.930 2097.490 2454.110 2098.670 ;
        RECT 2452.930 1919.090 2454.110 1920.270 ;
        RECT 2452.930 1917.490 2454.110 1918.670 ;
        RECT 2452.930 1739.090 2454.110 1740.270 ;
        RECT 2452.930 1737.490 2454.110 1738.670 ;
        RECT 2452.930 1559.090 2454.110 1560.270 ;
        RECT 2452.930 1557.490 2454.110 1558.670 ;
        RECT 2452.930 1379.090 2454.110 1380.270 ;
        RECT 2452.930 1377.490 2454.110 1378.670 ;
        RECT 2452.930 1199.090 2454.110 1200.270 ;
        RECT 2452.930 1197.490 2454.110 1198.670 ;
        RECT 2452.930 1019.090 2454.110 1020.270 ;
        RECT 2452.930 1017.490 2454.110 1018.670 ;
        RECT 2452.930 839.090 2454.110 840.270 ;
        RECT 2452.930 837.490 2454.110 838.670 ;
        RECT 2452.930 659.090 2454.110 660.270 ;
        RECT 2452.930 657.490 2454.110 658.670 ;
        RECT 2452.930 479.090 2454.110 480.270 ;
        RECT 2452.930 477.490 2454.110 478.670 ;
        RECT 2452.930 299.090 2454.110 300.270 ;
        RECT 2452.930 297.490 2454.110 298.670 ;
        RECT 2452.930 119.090 2454.110 120.270 ;
        RECT 2452.930 117.490 2454.110 118.670 ;
        RECT 2452.930 -17.010 2454.110 -15.830 ;
        RECT 2452.930 -18.610 2454.110 -17.430 ;
        RECT 2470.930 2657.090 2472.110 2658.270 ;
        RECT 2470.930 2655.490 2472.110 2656.670 ;
        RECT 2470.930 2477.090 2472.110 2478.270 ;
        RECT 2470.930 2475.490 2472.110 2476.670 ;
        RECT 2470.930 2297.090 2472.110 2298.270 ;
        RECT 2470.930 2295.490 2472.110 2296.670 ;
        RECT 2470.930 2117.090 2472.110 2118.270 ;
        RECT 2470.930 2115.490 2472.110 2116.670 ;
        RECT 2470.930 1937.090 2472.110 1938.270 ;
        RECT 2470.930 1935.490 2472.110 1936.670 ;
        RECT 2470.930 1757.090 2472.110 1758.270 ;
        RECT 2470.930 1755.490 2472.110 1756.670 ;
        RECT 2470.930 1577.090 2472.110 1578.270 ;
        RECT 2470.930 1575.490 2472.110 1576.670 ;
        RECT 2470.930 1397.090 2472.110 1398.270 ;
        RECT 2470.930 1395.490 2472.110 1396.670 ;
        RECT 2470.930 1217.090 2472.110 1218.270 ;
        RECT 2470.930 1215.490 2472.110 1216.670 ;
        RECT 2470.930 1037.090 2472.110 1038.270 ;
        RECT 2470.930 1035.490 2472.110 1036.670 ;
        RECT 2470.930 857.090 2472.110 858.270 ;
        RECT 2470.930 855.490 2472.110 856.670 ;
        RECT 2470.930 677.090 2472.110 678.270 ;
        RECT 2470.930 675.490 2472.110 676.670 ;
        RECT 2470.930 497.090 2472.110 498.270 ;
        RECT 2470.930 495.490 2472.110 496.670 ;
        RECT 2470.930 317.090 2472.110 318.270 ;
        RECT 2470.930 315.490 2472.110 316.670 ;
        RECT 2470.930 137.090 2472.110 138.270 ;
        RECT 2470.930 135.490 2472.110 136.670 ;
        RECT 2470.930 -26.410 2472.110 -25.230 ;
        RECT 2470.930 -28.010 2472.110 -26.830 ;
        RECT 2488.930 2675.090 2490.110 2676.270 ;
        RECT 2488.930 2673.490 2490.110 2674.670 ;
        RECT 2488.930 2495.090 2490.110 2496.270 ;
        RECT 2488.930 2493.490 2490.110 2494.670 ;
        RECT 2488.930 2315.090 2490.110 2316.270 ;
        RECT 2488.930 2313.490 2490.110 2314.670 ;
        RECT 2488.930 2135.090 2490.110 2136.270 ;
        RECT 2488.930 2133.490 2490.110 2134.670 ;
        RECT 2488.930 1955.090 2490.110 1956.270 ;
        RECT 2488.930 1953.490 2490.110 1954.670 ;
        RECT 2488.930 1775.090 2490.110 1776.270 ;
        RECT 2488.930 1773.490 2490.110 1774.670 ;
        RECT 2488.930 1595.090 2490.110 1596.270 ;
        RECT 2488.930 1593.490 2490.110 1594.670 ;
        RECT 2488.930 1415.090 2490.110 1416.270 ;
        RECT 2488.930 1413.490 2490.110 1414.670 ;
        RECT 2488.930 1235.090 2490.110 1236.270 ;
        RECT 2488.930 1233.490 2490.110 1234.670 ;
        RECT 2488.930 1055.090 2490.110 1056.270 ;
        RECT 2488.930 1053.490 2490.110 1054.670 ;
        RECT 2488.930 875.090 2490.110 876.270 ;
        RECT 2488.930 873.490 2490.110 874.670 ;
        RECT 2488.930 695.090 2490.110 696.270 ;
        RECT 2488.930 693.490 2490.110 694.670 ;
        RECT 2488.930 515.090 2490.110 516.270 ;
        RECT 2488.930 513.490 2490.110 514.670 ;
        RECT 2488.930 335.090 2490.110 336.270 ;
        RECT 2488.930 333.490 2490.110 334.670 ;
        RECT 2488.930 155.090 2490.110 156.270 ;
        RECT 2488.930 153.490 2490.110 154.670 ;
        RECT 2308.930 -35.810 2310.110 -34.630 ;
        RECT 2308.930 -37.410 2310.110 -36.230 ;
        RECT 2614.930 2621.090 2616.110 2622.270 ;
        RECT 2614.930 2619.490 2616.110 2620.670 ;
        RECT 2614.930 2441.090 2616.110 2442.270 ;
        RECT 2614.930 2439.490 2616.110 2440.670 ;
        RECT 2614.930 2261.090 2616.110 2262.270 ;
        RECT 2614.930 2259.490 2616.110 2260.670 ;
        RECT 2614.930 2081.090 2616.110 2082.270 ;
        RECT 2614.930 2079.490 2616.110 2080.670 ;
        RECT 2614.930 1901.090 2616.110 1902.270 ;
        RECT 2614.930 1899.490 2616.110 1900.670 ;
        RECT 2614.930 1721.090 2616.110 1722.270 ;
        RECT 2614.930 1719.490 2616.110 1720.670 ;
        RECT 2614.930 1541.090 2616.110 1542.270 ;
        RECT 2614.930 1539.490 2616.110 1540.670 ;
        RECT 2614.930 1361.090 2616.110 1362.270 ;
        RECT 2614.930 1359.490 2616.110 1360.670 ;
        RECT 2614.930 1181.090 2616.110 1182.270 ;
        RECT 2614.930 1179.490 2616.110 1180.670 ;
        RECT 2614.930 1001.090 2616.110 1002.270 ;
        RECT 2614.930 999.490 2616.110 1000.670 ;
        RECT 2614.930 821.090 2616.110 822.270 ;
        RECT 2614.930 819.490 2616.110 820.670 ;
        RECT 2614.930 641.090 2616.110 642.270 ;
        RECT 2614.930 639.490 2616.110 640.670 ;
        RECT 2614.930 461.090 2616.110 462.270 ;
        RECT 2614.930 459.490 2616.110 460.670 ;
        RECT 2614.930 281.090 2616.110 282.270 ;
        RECT 2614.930 279.490 2616.110 280.670 ;
        RECT 2614.930 101.090 2616.110 102.270 ;
        RECT 2614.930 99.490 2616.110 100.670 ;
        RECT 2614.930 -7.610 2616.110 -6.430 ;
        RECT 2614.930 -9.210 2616.110 -8.030 ;
        RECT 2632.930 3359.090 2634.110 3360.270 ;
        RECT 2632.930 3357.490 2634.110 3358.670 ;
        RECT 2632.930 3179.090 2634.110 3180.270 ;
        RECT 2632.930 3177.490 2634.110 3178.670 ;
        RECT 2632.930 2999.090 2634.110 3000.270 ;
        RECT 2632.930 2997.490 2634.110 2998.670 ;
        RECT 2632.930 2819.090 2634.110 2820.270 ;
        RECT 2632.930 2817.490 2634.110 2818.670 ;
        RECT 2632.930 2639.090 2634.110 2640.270 ;
        RECT 2632.930 2637.490 2634.110 2638.670 ;
        RECT 2632.930 2459.090 2634.110 2460.270 ;
        RECT 2632.930 2457.490 2634.110 2458.670 ;
        RECT 2632.930 2279.090 2634.110 2280.270 ;
        RECT 2632.930 2277.490 2634.110 2278.670 ;
        RECT 2632.930 2099.090 2634.110 2100.270 ;
        RECT 2632.930 2097.490 2634.110 2098.670 ;
        RECT 2632.930 1919.090 2634.110 1920.270 ;
        RECT 2632.930 1917.490 2634.110 1918.670 ;
        RECT 2632.930 1739.090 2634.110 1740.270 ;
        RECT 2632.930 1737.490 2634.110 1738.670 ;
        RECT 2632.930 1559.090 2634.110 1560.270 ;
        RECT 2632.930 1557.490 2634.110 1558.670 ;
        RECT 2632.930 1379.090 2634.110 1380.270 ;
        RECT 2632.930 1377.490 2634.110 1378.670 ;
        RECT 2632.930 1199.090 2634.110 1200.270 ;
        RECT 2632.930 1197.490 2634.110 1198.670 ;
        RECT 2632.930 1019.090 2634.110 1020.270 ;
        RECT 2632.930 1017.490 2634.110 1018.670 ;
        RECT 2632.930 839.090 2634.110 840.270 ;
        RECT 2632.930 837.490 2634.110 838.670 ;
        RECT 2632.930 659.090 2634.110 660.270 ;
        RECT 2632.930 657.490 2634.110 658.670 ;
        RECT 2632.930 479.090 2634.110 480.270 ;
        RECT 2632.930 477.490 2634.110 478.670 ;
        RECT 2632.930 299.090 2634.110 300.270 ;
        RECT 2632.930 297.490 2634.110 298.670 ;
        RECT 2632.930 119.090 2634.110 120.270 ;
        RECT 2632.930 117.490 2634.110 118.670 ;
        RECT 2632.930 -17.010 2634.110 -15.830 ;
        RECT 2632.930 -18.610 2634.110 -17.430 ;
        RECT 2650.930 3377.090 2652.110 3378.270 ;
        RECT 2650.930 3375.490 2652.110 3376.670 ;
        RECT 2650.930 3197.090 2652.110 3198.270 ;
        RECT 2650.930 3195.490 2652.110 3196.670 ;
        RECT 2650.930 3017.090 2652.110 3018.270 ;
        RECT 2650.930 3015.490 2652.110 3016.670 ;
        RECT 2650.930 2837.090 2652.110 2838.270 ;
        RECT 2650.930 2835.490 2652.110 2836.670 ;
        RECT 2650.930 2657.090 2652.110 2658.270 ;
        RECT 2650.930 2655.490 2652.110 2656.670 ;
        RECT 2650.930 2477.090 2652.110 2478.270 ;
        RECT 2650.930 2475.490 2652.110 2476.670 ;
        RECT 2650.930 2297.090 2652.110 2298.270 ;
        RECT 2650.930 2295.490 2652.110 2296.670 ;
        RECT 2650.930 2117.090 2652.110 2118.270 ;
        RECT 2650.930 2115.490 2652.110 2116.670 ;
        RECT 2650.930 1937.090 2652.110 1938.270 ;
        RECT 2650.930 1935.490 2652.110 1936.670 ;
        RECT 2650.930 1757.090 2652.110 1758.270 ;
        RECT 2650.930 1755.490 2652.110 1756.670 ;
        RECT 2650.930 1577.090 2652.110 1578.270 ;
        RECT 2650.930 1575.490 2652.110 1576.670 ;
        RECT 2650.930 1397.090 2652.110 1398.270 ;
        RECT 2650.930 1395.490 2652.110 1396.670 ;
        RECT 2650.930 1217.090 2652.110 1218.270 ;
        RECT 2650.930 1215.490 2652.110 1216.670 ;
        RECT 2650.930 1037.090 2652.110 1038.270 ;
        RECT 2650.930 1035.490 2652.110 1036.670 ;
        RECT 2650.930 857.090 2652.110 858.270 ;
        RECT 2650.930 855.490 2652.110 856.670 ;
        RECT 2650.930 677.090 2652.110 678.270 ;
        RECT 2650.930 675.490 2652.110 676.670 ;
        RECT 2650.930 497.090 2652.110 498.270 ;
        RECT 2650.930 495.490 2652.110 496.670 ;
        RECT 2650.930 317.090 2652.110 318.270 ;
        RECT 2650.930 315.490 2652.110 316.670 ;
        RECT 2650.930 137.090 2652.110 138.270 ;
        RECT 2650.930 135.490 2652.110 136.670 ;
        RECT 2650.930 -26.410 2652.110 -25.230 ;
        RECT 2650.930 -28.010 2652.110 -26.830 ;
        RECT 2848.930 3555.910 2850.110 3557.090 ;
        RECT 2848.930 3554.310 2850.110 3555.490 ;
        RECT 2830.930 3546.510 2832.110 3547.690 ;
        RECT 2830.930 3544.910 2832.110 3546.090 ;
        RECT 2812.930 3537.110 2814.110 3538.290 ;
        RECT 2812.930 3535.510 2814.110 3536.690 ;
        RECT 2668.930 3395.090 2670.110 3396.270 ;
        RECT 2668.930 3393.490 2670.110 3394.670 ;
        RECT 2668.930 3215.090 2670.110 3216.270 ;
        RECT 2668.930 3213.490 2670.110 3214.670 ;
        RECT 2668.930 3035.090 2670.110 3036.270 ;
        RECT 2668.930 3033.490 2670.110 3034.670 ;
        RECT 2668.930 2855.090 2670.110 2856.270 ;
        RECT 2668.930 2853.490 2670.110 2854.670 ;
        RECT 2668.930 2675.090 2670.110 2676.270 ;
        RECT 2668.930 2673.490 2670.110 2674.670 ;
        RECT 2668.930 2495.090 2670.110 2496.270 ;
        RECT 2668.930 2493.490 2670.110 2494.670 ;
        RECT 2668.930 2315.090 2670.110 2316.270 ;
        RECT 2668.930 2313.490 2670.110 2314.670 ;
        RECT 2668.930 2135.090 2670.110 2136.270 ;
        RECT 2668.930 2133.490 2670.110 2134.670 ;
        RECT 2668.930 1955.090 2670.110 1956.270 ;
        RECT 2668.930 1953.490 2670.110 1954.670 ;
        RECT 2668.930 1775.090 2670.110 1776.270 ;
        RECT 2668.930 1773.490 2670.110 1774.670 ;
        RECT 2668.930 1595.090 2670.110 1596.270 ;
        RECT 2668.930 1593.490 2670.110 1594.670 ;
        RECT 2668.930 1415.090 2670.110 1416.270 ;
        RECT 2668.930 1413.490 2670.110 1414.670 ;
        RECT 2668.930 1235.090 2670.110 1236.270 ;
        RECT 2668.930 1233.490 2670.110 1234.670 ;
        RECT 2668.930 1055.090 2670.110 1056.270 ;
        RECT 2668.930 1053.490 2670.110 1054.670 ;
        RECT 2668.930 875.090 2670.110 876.270 ;
        RECT 2668.930 873.490 2670.110 874.670 ;
        RECT 2668.930 695.090 2670.110 696.270 ;
        RECT 2668.930 693.490 2670.110 694.670 ;
        RECT 2668.930 515.090 2670.110 516.270 ;
        RECT 2668.930 513.490 2670.110 514.670 ;
        RECT 2668.930 335.090 2670.110 336.270 ;
        RECT 2668.930 333.490 2670.110 334.670 ;
        RECT 2668.930 155.090 2670.110 156.270 ;
        RECT 2668.930 153.490 2670.110 154.670 ;
        RECT 2488.930 -35.810 2490.110 -34.630 ;
        RECT 2488.930 -37.410 2490.110 -36.230 ;
        RECT 2794.930 3527.710 2796.110 3528.890 ;
        RECT 2794.930 3526.110 2796.110 3527.290 ;
        RECT 2794.930 3341.090 2796.110 3342.270 ;
        RECT 2794.930 3339.490 2796.110 3340.670 ;
        RECT 2794.930 3161.090 2796.110 3162.270 ;
        RECT 2794.930 3159.490 2796.110 3160.670 ;
        RECT 2794.930 2981.090 2796.110 2982.270 ;
        RECT 2794.930 2979.490 2796.110 2980.670 ;
        RECT 2794.930 2801.090 2796.110 2802.270 ;
        RECT 2794.930 2799.490 2796.110 2800.670 ;
        RECT 2794.930 2621.090 2796.110 2622.270 ;
        RECT 2794.930 2619.490 2796.110 2620.670 ;
        RECT 2794.930 2441.090 2796.110 2442.270 ;
        RECT 2794.930 2439.490 2796.110 2440.670 ;
        RECT 2794.930 2261.090 2796.110 2262.270 ;
        RECT 2794.930 2259.490 2796.110 2260.670 ;
        RECT 2794.930 2081.090 2796.110 2082.270 ;
        RECT 2794.930 2079.490 2796.110 2080.670 ;
        RECT 2794.930 1901.090 2796.110 1902.270 ;
        RECT 2794.930 1899.490 2796.110 1900.670 ;
        RECT 2794.930 1721.090 2796.110 1722.270 ;
        RECT 2794.930 1719.490 2796.110 1720.670 ;
        RECT 2794.930 1541.090 2796.110 1542.270 ;
        RECT 2794.930 1539.490 2796.110 1540.670 ;
        RECT 2794.930 1361.090 2796.110 1362.270 ;
        RECT 2794.930 1359.490 2796.110 1360.670 ;
        RECT 2794.930 1181.090 2796.110 1182.270 ;
        RECT 2794.930 1179.490 2796.110 1180.670 ;
        RECT 2794.930 1001.090 2796.110 1002.270 ;
        RECT 2794.930 999.490 2796.110 1000.670 ;
        RECT 2794.930 821.090 2796.110 822.270 ;
        RECT 2794.930 819.490 2796.110 820.670 ;
        RECT 2794.930 641.090 2796.110 642.270 ;
        RECT 2794.930 639.490 2796.110 640.670 ;
        RECT 2794.930 461.090 2796.110 462.270 ;
        RECT 2794.930 459.490 2796.110 460.670 ;
        RECT 2794.930 281.090 2796.110 282.270 ;
        RECT 2794.930 279.490 2796.110 280.670 ;
        RECT 2794.930 101.090 2796.110 102.270 ;
        RECT 2794.930 99.490 2796.110 100.670 ;
        RECT 2794.930 -7.610 2796.110 -6.430 ;
        RECT 2794.930 -9.210 2796.110 -8.030 ;
        RECT 2812.930 3359.090 2814.110 3360.270 ;
        RECT 2812.930 3357.490 2814.110 3358.670 ;
        RECT 2812.930 3179.090 2814.110 3180.270 ;
        RECT 2812.930 3177.490 2814.110 3178.670 ;
        RECT 2812.930 2999.090 2814.110 3000.270 ;
        RECT 2812.930 2997.490 2814.110 2998.670 ;
        RECT 2812.930 2819.090 2814.110 2820.270 ;
        RECT 2812.930 2817.490 2814.110 2818.670 ;
        RECT 2812.930 2639.090 2814.110 2640.270 ;
        RECT 2812.930 2637.490 2814.110 2638.670 ;
        RECT 2812.930 2459.090 2814.110 2460.270 ;
        RECT 2812.930 2457.490 2814.110 2458.670 ;
        RECT 2812.930 2279.090 2814.110 2280.270 ;
        RECT 2812.930 2277.490 2814.110 2278.670 ;
        RECT 2812.930 2099.090 2814.110 2100.270 ;
        RECT 2812.930 2097.490 2814.110 2098.670 ;
        RECT 2812.930 1919.090 2814.110 1920.270 ;
        RECT 2812.930 1917.490 2814.110 1918.670 ;
        RECT 2812.930 1739.090 2814.110 1740.270 ;
        RECT 2812.930 1737.490 2814.110 1738.670 ;
        RECT 2812.930 1559.090 2814.110 1560.270 ;
        RECT 2812.930 1557.490 2814.110 1558.670 ;
        RECT 2812.930 1379.090 2814.110 1380.270 ;
        RECT 2812.930 1377.490 2814.110 1378.670 ;
        RECT 2812.930 1199.090 2814.110 1200.270 ;
        RECT 2812.930 1197.490 2814.110 1198.670 ;
        RECT 2812.930 1019.090 2814.110 1020.270 ;
        RECT 2812.930 1017.490 2814.110 1018.670 ;
        RECT 2812.930 839.090 2814.110 840.270 ;
        RECT 2812.930 837.490 2814.110 838.670 ;
        RECT 2812.930 659.090 2814.110 660.270 ;
        RECT 2812.930 657.490 2814.110 658.670 ;
        RECT 2812.930 479.090 2814.110 480.270 ;
        RECT 2812.930 477.490 2814.110 478.670 ;
        RECT 2812.930 299.090 2814.110 300.270 ;
        RECT 2812.930 297.490 2814.110 298.670 ;
        RECT 2812.930 119.090 2814.110 120.270 ;
        RECT 2812.930 117.490 2814.110 118.670 ;
        RECT 2812.930 -17.010 2814.110 -15.830 ;
        RECT 2812.930 -18.610 2814.110 -17.430 ;
        RECT 2830.930 3377.090 2832.110 3378.270 ;
        RECT 2830.930 3375.490 2832.110 3376.670 ;
        RECT 2830.930 3197.090 2832.110 3198.270 ;
        RECT 2830.930 3195.490 2832.110 3196.670 ;
        RECT 2830.930 3017.090 2832.110 3018.270 ;
        RECT 2830.930 3015.490 2832.110 3016.670 ;
        RECT 2830.930 2837.090 2832.110 2838.270 ;
        RECT 2830.930 2835.490 2832.110 2836.670 ;
        RECT 2830.930 2657.090 2832.110 2658.270 ;
        RECT 2830.930 2655.490 2832.110 2656.670 ;
        RECT 2830.930 2477.090 2832.110 2478.270 ;
        RECT 2830.930 2475.490 2832.110 2476.670 ;
        RECT 2830.930 2297.090 2832.110 2298.270 ;
        RECT 2830.930 2295.490 2832.110 2296.670 ;
        RECT 2830.930 2117.090 2832.110 2118.270 ;
        RECT 2830.930 2115.490 2832.110 2116.670 ;
        RECT 2830.930 1937.090 2832.110 1938.270 ;
        RECT 2830.930 1935.490 2832.110 1936.670 ;
        RECT 2830.930 1757.090 2832.110 1758.270 ;
        RECT 2830.930 1755.490 2832.110 1756.670 ;
        RECT 2830.930 1577.090 2832.110 1578.270 ;
        RECT 2830.930 1575.490 2832.110 1576.670 ;
        RECT 2830.930 1397.090 2832.110 1398.270 ;
        RECT 2830.930 1395.490 2832.110 1396.670 ;
        RECT 2830.930 1217.090 2832.110 1218.270 ;
        RECT 2830.930 1215.490 2832.110 1216.670 ;
        RECT 2830.930 1037.090 2832.110 1038.270 ;
        RECT 2830.930 1035.490 2832.110 1036.670 ;
        RECT 2830.930 857.090 2832.110 858.270 ;
        RECT 2830.930 855.490 2832.110 856.670 ;
        RECT 2830.930 677.090 2832.110 678.270 ;
        RECT 2830.930 675.490 2832.110 676.670 ;
        RECT 2830.930 497.090 2832.110 498.270 ;
        RECT 2830.930 495.490 2832.110 496.670 ;
        RECT 2830.930 317.090 2832.110 318.270 ;
        RECT 2830.930 315.490 2832.110 316.670 ;
        RECT 2830.930 137.090 2832.110 138.270 ;
        RECT 2830.930 135.490 2832.110 136.670 ;
        RECT 2830.930 -26.410 2832.110 -25.230 ;
        RECT 2830.930 -28.010 2832.110 -26.830 ;
        RECT 2960.410 3555.910 2961.590 3557.090 ;
        RECT 2960.410 3554.310 2961.590 3555.490 ;
        RECT 2951.010 3546.510 2952.190 3547.690 ;
        RECT 2951.010 3544.910 2952.190 3546.090 ;
        RECT 2941.610 3537.110 2942.790 3538.290 ;
        RECT 2941.610 3535.510 2942.790 3536.690 ;
        RECT 2848.930 3395.090 2850.110 3396.270 ;
        RECT 2848.930 3393.490 2850.110 3394.670 ;
        RECT 2848.930 3215.090 2850.110 3216.270 ;
        RECT 2848.930 3213.490 2850.110 3214.670 ;
        RECT 2848.930 3035.090 2850.110 3036.270 ;
        RECT 2848.930 3033.490 2850.110 3034.670 ;
        RECT 2848.930 2855.090 2850.110 2856.270 ;
        RECT 2848.930 2853.490 2850.110 2854.670 ;
        RECT 2848.930 2675.090 2850.110 2676.270 ;
        RECT 2848.930 2673.490 2850.110 2674.670 ;
        RECT 2848.930 2495.090 2850.110 2496.270 ;
        RECT 2848.930 2493.490 2850.110 2494.670 ;
        RECT 2848.930 2315.090 2850.110 2316.270 ;
        RECT 2848.930 2313.490 2850.110 2314.670 ;
        RECT 2848.930 2135.090 2850.110 2136.270 ;
        RECT 2848.930 2133.490 2850.110 2134.670 ;
        RECT 2848.930 1955.090 2850.110 1956.270 ;
        RECT 2848.930 1953.490 2850.110 1954.670 ;
        RECT 2848.930 1775.090 2850.110 1776.270 ;
        RECT 2848.930 1773.490 2850.110 1774.670 ;
        RECT 2848.930 1595.090 2850.110 1596.270 ;
        RECT 2848.930 1593.490 2850.110 1594.670 ;
        RECT 2848.930 1415.090 2850.110 1416.270 ;
        RECT 2848.930 1413.490 2850.110 1414.670 ;
        RECT 2848.930 1235.090 2850.110 1236.270 ;
        RECT 2848.930 1233.490 2850.110 1234.670 ;
        RECT 2848.930 1055.090 2850.110 1056.270 ;
        RECT 2848.930 1053.490 2850.110 1054.670 ;
        RECT 2848.930 875.090 2850.110 876.270 ;
        RECT 2848.930 873.490 2850.110 874.670 ;
        RECT 2848.930 695.090 2850.110 696.270 ;
        RECT 2848.930 693.490 2850.110 694.670 ;
        RECT 2848.930 515.090 2850.110 516.270 ;
        RECT 2848.930 513.490 2850.110 514.670 ;
        RECT 2848.930 335.090 2850.110 336.270 ;
        RECT 2848.930 333.490 2850.110 334.670 ;
        RECT 2848.930 155.090 2850.110 156.270 ;
        RECT 2848.930 153.490 2850.110 154.670 ;
        RECT 2668.930 -35.810 2670.110 -34.630 ;
        RECT 2668.930 -37.410 2670.110 -36.230 ;
        RECT 2932.210 3527.710 2933.390 3528.890 ;
        RECT 2932.210 3526.110 2933.390 3527.290 ;
        RECT 2932.210 3341.090 2933.390 3342.270 ;
        RECT 2932.210 3339.490 2933.390 3340.670 ;
        RECT 2932.210 3161.090 2933.390 3162.270 ;
        RECT 2932.210 3159.490 2933.390 3160.670 ;
        RECT 2932.210 2981.090 2933.390 2982.270 ;
        RECT 2932.210 2979.490 2933.390 2980.670 ;
        RECT 2932.210 2801.090 2933.390 2802.270 ;
        RECT 2932.210 2799.490 2933.390 2800.670 ;
        RECT 2932.210 2621.090 2933.390 2622.270 ;
        RECT 2932.210 2619.490 2933.390 2620.670 ;
        RECT 2932.210 2441.090 2933.390 2442.270 ;
        RECT 2932.210 2439.490 2933.390 2440.670 ;
        RECT 2932.210 2261.090 2933.390 2262.270 ;
        RECT 2932.210 2259.490 2933.390 2260.670 ;
        RECT 2932.210 2081.090 2933.390 2082.270 ;
        RECT 2932.210 2079.490 2933.390 2080.670 ;
        RECT 2932.210 1901.090 2933.390 1902.270 ;
        RECT 2932.210 1899.490 2933.390 1900.670 ;
        RECT 2932.210 1721.090 2933.390 1722.270 ;
        RECT 2932.210 1719.490 2933.390 1720.670 ;
        RECT 2932.210 1541.090 2933.390 1542.270 ;
        RECT 2932.210 1539.490 2933.390 1540.670 ;
        RECT 2932.210 1361.090 2933.390 1362.270 ;
        RECT 2932.210 1359.490 2933.390 1360.670 ;
        RECT 2932.210 1181.090 2933.390 1182.270 ;
        RECT 2932.210 1179.490 2933.390 1180.670 ;
        RECT 2932.210 1001.090 2933.390 1002.270 ;
        RECT 2932.210 999.490 2933.390 1000.670 ;
        RECT 2932.210 821.090 2933.390 822.270 ;
        RECT 2932.210 819.490 2933.390 820.670 ;
        RECT 2932.210 641.090 2933.390 642.270 ;
        RECT 2932.210 639.490 2933.390 640.670 ;
        RECT 2932.210 461.090 2933.390 462.270 ;
        RECT 2932.210 459.490 2933.390 460.670 ;
        RECT 2932.210 281.090 2933.390 282.270 ;
        RECT 2932.210 279.490 2933.390 280.670 ;
        RECT 2932.210 101.090 2933.390 102.270 ;
        RECT 2932.210 99.490 2933.390 100.670 ;
        RECT 2932.210 -7.610 2933.390 -6.430 ;
        RECT 2932.210 -9.210 2933.390 -8.030 ;
        RECT 2941.610 3359.090 2942.790 3360.270 ;
        RECT 2941.610 3357.490 2942.790 3358.670 ;
        RECT 2941.610 3179.090 2942.790 3180.270 ;
        RECT 2941.610 3177.490 2942.790 3178.670 ;
        RECT 2941.610 2999.090 2942.790 3000.270 ;
        RECT 2941.610 2997.490 2942.790 2998.670 ;
        RECT 2941.610 2819.090 2942.790 2820.270 ;
        RECT 2941.610 2817.490 2942.790 2818.670 ;
        RECT 2941.610 2639.090 2942.790 2640.270 ;
        RECT 2941.610 2637.490 2942.790 2638.670 ;
        RECT 2941.610 2459.090 2942.790 2460.270 ;
        RECT 2941.610 2457.490 2942.790 2458.670 ;
        RECT 2941.610 2279.090 2942.790 2280.270 ;
        RECT 2941.610 2277.490 2942.790 2278.670 ;
        RECT 2941.610 2099.090 2942.790 2100.270 ;
        RECT 2941.610 2097.490 2942.790 2098.670 ;
        RECT 2941.610 1919.090 2942.790 1920.270 ;
        RECT 2941.610 1917.490 2942.790 1918.670 ;
        RECT 2941.610 1739.090 2942.790 1740.270 ;
        RECT 2941.610 1737.490 2942.790 1738.670 ;
        RECT 2941.610 1559.090 2942.790 1560.270 ;
        RECT 2941.610 1557.490 2942.790 1558.670 ;
        RECT 2941.610 1379.090 2942.790 1380.270 ;
        RECT 2941.610 1377.490 2942.790 1378.670 ;
        RECT 2941.610 1199.090 2942.790 1200.270 ;
        RECT 2941.610 1197.490 2942.790 1198.670 ;
        RECT 2941.610 1019.090 2942.790 1020.270 ;
        RECT 2941.610 1017.490 2942.790 1018.670 ;
        RECT 2941.610 839.090 2942.790 840.270 ;
        RECT 2941.610 837.490 2942.790 838.670 ;
        RECT 2941.610 659.090 2942.790 660.270 ;
        RECT 2941.610 657.490 2942.790 658.670 ;
        RECT 2941.610 479.090 2942.790 480.270 ;
        RECT 2941.610 477.490 2942.790 478.670 ;
        RECT 2941.610 299.090 2942.790 300.270 ;
        RECT 2941.610 297.490 2942.790 298.670 ;
        RECT 2941.610 119.090 2942.790 120.270 ;
        RECT 2941.610 117.490 2942.790 118.670 ;
        RECT 2941.610 -17.010 2942.790 -15.830 ;
        RECT 2941.610 -18.610 2942.790 -17.430 ;
        RECT 2951.010 3377.090 2952.190 3378.270 ;
        RECT 2951.010 3375.490 2952.190 3376.670 ;
        RECT 2951.010 3197.090 2952.190 3198.270 ;
        RECT 2951.010 3195.490 2952.190 3196.670 ;
        RECT 2951.010 3017.090 2952.190 3018.270 ;
        RECT 2951.010 3015.490 2952.190 3016.670 ;
        RECT 2951.010 2837.090 2952.190 2838.270 ;
        RECT 2951.010 2835.490 2952.190 2836.670 ;
        RECT 2951.010 2657.090 2952.190 2658.270 ;
        RECT 2951.010 2655.490 2952.190 2656.670 ;
        RECT 2951.010 2477.090 2952.190 2478.270 ;
        RECT 2951.010 2475.490 2952.190 2476.670 ;
        RECT 2951.010 2297.090 2952.190 2298.270 ;
        RECT 2951.010 2295.490 2952.190 2296.670 ;
        RECT 2951.010 2117.090 2952.190 2118.270 ;
        RECT 2951.010 2115.490 2952.190 2116.670 ;
        RECT 2951.010 1937.090 2952.190 1938.270 ;
        RECT 2951.010 1935.490 2952.190 1936.670 ;
        RECT 2951.010 1757.090 2952.190 1758.270 ;
        RECT 2951.010 1755.490 2952.190 1756.670 ;
        RECT 2951.010 1577.090 2952.190 1578.270 ;
        RECT 2951.010 1575.490 2952.190 1576.670 ;
        RECT 2951.010 1397.090 2952.190 1398.270 ;
        RECT 2951.010 1395.490 2952.190 1396.670 ;
        RECT 2951.010 1217.090 2952.190 1218.270 ;
        RECT 2951.010 1215.490 2952.190 1216.670 ;
        RECT 2951.010 1037.090 2952.190 1038.270 ;
        RECT 2951.010 1035.490 2952.190 1036.670 ;
        RECT 2951.010 857.090 2952.190 858.270 ;
        RECT 2951.010 855.490 2952.190 856.670 ;
        RECT 2951.010 677.090 2952.190 678.270 ;
        RECT 2951.010 675.490 2952.190 676.670 ;
        RECT 2951.010 497.090 2952.190 498.270 ;
        RECT 2951.010 495.490 2952.190 496.670 ;
        RECT 2951.010 317.090 2952.190 318.270 ;
        RECT 2951.010 315.490 2952.190 316.670 ;
        RECT 2951.010 137.090 2952.190 138.270 ;
        RECT 2951.010 135.490 2952.190 136.670 ;
        RECT 2951.010 -26.410 2952.190 -25.230 ;
        RECT 2951.010 -28.010 2952.190 -26.830 ;
        RECT 2960.410 3395.090 2961.590 3396.270 ;
        RECT 2960.410 3393.490 2961.590 3394.670 ;
        RECT 2960.410 3215.090 2961.590 3216.270 ;
        RECT 2960.410 3213.490 2961.590 3214.670 ;
        RECT 2960.410 3035.090 2961.590 3036.270 ;
        RECT 2960.410 3033.490 2961.590 3034.670 ;
        RECT 2960.410 2855.090 2961.590 2856.270 ;
        RECT 2960.410 2853.490 2961.590 2854.670 ;
        RECT 2960.410 2675.090 2961.590 2676.270 ;
        RECT 2960.410 2673.490 2961.590 2674.670 ;
        RECT 2960.410 2495.090 2961.590 2496.270 ;
        RECT 2960.410 2493.490 2961.590 2494.670 ;
        RECT 2960.410 2315.090 2961.590 2316.270 ;
        RECT 2960.410 2313.490 2961.590 2314.670 ;
        RECT 2960.410 2135.090 2961.590 2136.270 ;
        RECT 2960.410 2133.490 2961.590 2134.670 ;
        RECT 2960.410 1955.090 2961.590 1956.270 ;
        RECT 2960.410 1953.490 2961.590 1954.670 ;
        RECT 2960.410 1775.090 2961.590 1776.270 ;
        RECT 2960.410 1773.490 2961.590 1774.670 ;
        RECT 2960.410 1595.090 2961.590 1596.270 ;
        RECT 2960.410 1593.490 2961.590 1594.670 ;
        RECT 2960.410 1415.090 2961.590 1416.270 ;
        RECT 2960.410 1413.490 2961.590 1414.670 ;
        RECT 2960.410 1235.090 2961.590 1236.270 ;
        RECT 2960.410 1233.490 2961.590 1234.670 ;
        RECT 2960.410 1055.090 2961.590 1056.270 ;
        RECT 2960.410 1053.490 2961.590 1054.670 ;
        RECT 2960.410 875.090 2961.590 876.270 ;
        RECT 2960.410 873.490 2961.590 874.670 ;
        RECT 2960.410 695.090 2961.590 696.270 ;
        RECT 2960.410 693.490 2961.590 694.670 ;
        RECT 2960.410 515.090 2961.590 516.270 ;
        RECT 2960.410 513.490 2961.590 514.670 ;
        RECT 2960.410 335.090 2961.590 336.270 ;
        RECT 2960.410 333.490 2961.590 334.670 ;
        RECT 2960.410 155.090 2961.590 156.270 ;
        RECT 2960.410 153.490 2961.590 154.670 ;
        RECT 2848.930 -35.810 2850.110 -34.630 ;
        RECT 2848.930 -37.410 2850.110 -36.230 ;
        RECT 2960.410 -35.810 2961.590 -34.630 ;
        RECT 2960.410 -37.410 2961.590 -36.230 ;
      LAYER met5 ;
        RECT -42.880 3557.200 -39.880 3557.210 ;
        RECT 148.020 3557.200 151.020 3557.210 ;
        RECT 328.020 3557.200 331.020 3557.210 ;
        RECT 508.020 3557.200 511.020 3557.210 ;
        RECT 688.020 3557.200 691.020 3557.210 ;
        RECT 868.020 3557.200 871.020 3557.210 ;
        RECT 1048.020 3557.200 1051.020 3557.210 ;
        RECT 1228.020 3557.200 1231.020 3557.210 ;
        RECT 1408.020 3557.200 1411.020 3557.210 ;
        RECT 1588.020 3557.200 1591.020 3557.210 ;
        RECT 1768.020 3557.200 1771.020 3557.210 ;
        RECT 1948.020 3557.200 1951.020 3557.210 ;
        RECT 2128.020 3557.200 2131.020 3557.210 ;
        RECT 2308.020 3557.200 2311.020 3557.210 ;
        RECT 2488.020 3557.200 2491.020 3557.210 ;
        RECT 2668.020 3557.200 2671.020 3557.210 ;
        RECT 2848.020 3557.200 2851.020 3557.210 ;
        RECT 2959.500 3557.200 2962.500 3557.210 ;
        RECT -42.880 3554.200 2962.500 3557.200 ;
        RECT -42.880 3554.190 -39.880 3554.200 ;
        RECT 148.020 3554.190 151.020 3554.200 ;
        RECT 328.020 3554.190 331.020 3554.200 ;
        RECT 508.020 3554.190 511.020 3554.200 ;
        RECT 688.020 3554.190 691.020 3554.200 ;
        RECT 868.020 3554.190 871.020 3554.200 ;
        RECT 1048.020 3554.190 1051.020 3554.200 ;
        RECT 1228.020 3554.190 1231.020 3554.200 ;
        RECT 1408.020 3554.190 1411.020 3554.200 ;
        RECT 1588.020 3554.190 1591.020 3554.200 ;
        RECT 1768.020 3554.190 1771.020 3554.200 ;
        RECT 1948.020 3554.190 1951.020 3554.200 ;
        RECT 2128.020 3554.190 2131.020 3554.200 ;
        RECT 2308.020 3554.190 2311.020 3554.200 ;
        RECT 2488.020 3554.190 2491.020 3554.200 ;
        RECT 2668.020 3554.190 2671.020 3554.200 ;
        RECT 2848.020 3554.190 2851.020 3554.200 ;
        RECT 2959.500 3554.190 2962.500 3554.200 ;
        RECT -33.480 3547.800 -30.480 3547.810 ;
        RECT 130.020 3547.800 133.020 3547.810 ;
        RECT 310.020 3547.800 313.020 3547.810 ;
        RECT 490.020 3547.800 493.020 3547.810 ;
        RECT 670.020 3547.800 673.020 3547.810 ;
        RECT 850.020 3547.800 853.020 3547.810 ;
        RECT 1030.020 3547.800 1033.020 3547.810 ;
        RECT 1210.020 3547.800 1213.020 3547.810 ;
        RECT 1390.020 3547.800 1393.020 3547.810 ;
        RECT 1570.020 3547.800 1573.020 3547.810 ;
        RECT 1750.020 3547.800 1753.020 3547.810 ;
        RECT 1930.020 3547.800 1933.020 3547.810 ;
        RECT 2110.020 3547.800 2113.020 3547.810 ;
        RECT 2290.020 3547.800 2293.020 3547.810 ;
        RECT 2470.020 3547.800 2473.020 3547.810 ;
        RECT 2650.020 3547.800 2653.020 3547.810 ;
        RECT 2830.020 3547.800 2833.020 3547.810 ;
        RECT 2950.100 3547.800 2953.100 3547.810 ;
        RECT -33.480 3544.800 2953.100 3547.800 ;
        RECT -33.480 3544.790 -30.480 3544.800 ;
        RECT 130.020 3544.790 133.020 3544.800 ;
        RECT 310.020 3544.790 313.020 3544.800 ;
        RECT 490.020 3544.790 493.020 3544.800 ;
        RECT 670.020 3544.790 673.020 3544.800 ;
        RECT 850.020 3544.790 853.020 3544.800 ;
        RECT 1030.020 3544.790 1033.020 3544.800 ;
        RECT 1210.020 3544.790 1213.020 3544.800 ;
        RECT 1390.020 3544.790 1393.020 3544.800 ;
        RECT 1570.020 3544.790 1573.020 3544.800 ;
        RECT 1750.020 3544.790 1753.020 3544.800 ;
        RECT 1930.020 3544.790 1933.020 3544.800 ;
        RECT 2110.020 3544.790 2113.020 3544.800 ;
        RECT 2290.020 3544.790 2293.020 3544.800 ;
        RECT 2470.020 3544.790 2473.020 3544.800 ;
        RECT 2650.020 3544.790 2653.020 3544.800 ;
        RECT 2830.020 3544.790 2833.020 3544.800 ;
        RECT 2950.100 3544.790 2953.100 3544.800 ;
        RECT -24.080 3538.400 -21.080 3538.410 ;
        RECT 112.020 3538.400 115.020 3538.410 ;
        RECT 292.020 3538.400 295.020 3538.410 ;
        RECT 472.020 3538.400 475.020 3538.410 ;
        RECT 652.020 3538.400 655.020 3538.410 ;
        RECT 832.020 3538.400 835.020 3538.410 ;
        RECT 1012.020 3538.400 1015.020 3538.410 ;
        RECT 1192.020 3538.400 1195.020 3538.410 ;
        RECT 1372.020 3538.400 1375.020 3538.410 ;
        RECT 1552.020 3538.400 1555.020 3538.410 ;
        RECT 1732.020 3538.400 1735.020 3538.410 ;
        RECT 1912.020 3538.400 1915.020 3538.410 ;
        RECT 2092.020 3538.400 2095.020 3538.410 ;
        RECT 2272.020 3538.400 2275.020 3538.410 ;
        RECT 2452.020 3538.400 2455.020 3538.410 ;
        RECT 2632.020 3538.400 2635.020 3538.410 ;
        RECT 2812.020 3538.400 2815.020 3538.410 ;
        RECT 2940.700 3538.400 2943.700 3538.410 ;
        RECT -24.080 3535.400 2943.700 3538.400 ;
        RECT -24.080 3535.390 -21.080 3535.400 ;
        RECT 112.020 3535.390 115.020 3535.400 ;
        RECT 292.020 3535.390 295.020 3535.400 ;
        RECT 472.020 3535.390 475.020 3535.400 ;
        RECT 652.020 3535.390 655.020 3535.400 ;
        RECT 832.020 3535.390 835.020 3535.400 ;
        RECT 1012.020 3535.390 1015.020 3535.400 ;
        RECT 1192.020 3535.390 1195.020 3535.400 ;
        RECT 1372.020 3535.390 1375.020 3535.400 ;
        RECT 1552.020 3535.390 1555.020 3535.400 ;
        RECT 1732.020 3535.390 1735.020 3535.400 ;
        RECT 1912.020 3535.390 1915.020 3535.400 ;
        RECT 2092.020 3535.390 2095.020 3535.400 ;
        RECT 2272.020 3535.390 2275.020 3535.400 ;
        RECT 2452.020 3535.390 2455.020 3535.400 ;
        RECT 2632.020 3535.390 2635.020 3535.400 ;
        RECT 2812.020 3535.390 2815.020 3535.400 ;
        RECT 2940.700 3535.390 2943.700 3535.400 ;
        RECT -14.680 3529.000 -11.680 3529.010 ;
        RECT 94.020 3529.000 97.020 3529.010 ;
        RECT 274.020 3529.000 277.020 3529.010 ;
        RECT 454.020 3529.000 457.020 3529.010 ;
        RECT 634.020 3529.000 637.020 3529.010 ;
        RECT 814.020 3529.000 817.020 3529.010 ;
        RECT 994.020 3529.000 997.020 3529.010 ;
        RECT 1174.020 3529.000 1177.020 3529.010 ;
        RECT 1354.020 3529.000 1357.020 3529.010 ;
        RECT 1534.020 3529.000 1537.020 3529.010 ;
        RECT 1714.020 3529.000 1717.020 3529.010 ;
        RECT 1894.020 3529.000 1897.020 3529.010 ;
        RECT 2074.020 3529.000 2077.020 3529.010 ;
        RECT 2254.020 3529.000 2257.020 3529.010 ;
        RECT 2434.020 3529.000 2437.020 3529.010 ;
        RECT 2614.020 3529.000 2617.020 3529.010 ;
        RECT 2794.020 3529.000 2797.020 3529.010 ;
        RECT 2931.300 3529.000 2934.300 3529.010 ;
        RECT -14.680 3526.000 2934.300 3529.000 ;
        RECT -14.680 3525.990 -11.680 3526.000 ;
        RECT 94.020 3525.990 97.020 3526.000 ;
        RECT 274.020 3525.990 277.020 3526.000 ;
        RECT 454.020 3525.990 457.020 3526.000 ;
        RECT 634.020 3525.990 637.020 3526.000 ;
        RECT 814.020 3525.990 817.020 3526.000 ;
        RECT 994.020 3525.990 997.020 3526.000 ;
        RECT 1174.020 3525.990 1177.020 3526.000 ;
        RECT 1354.020 3525.990 1357.020 3526.000 ;
        RECT 1534.020 3525.990 1537.020 3526.000 ;
        RECT 1714.020 3525.990 1717.020 3526.000 ;
        RECT 1894.020 3525.990 1897.020 3526.000 ;
        RECT 2074.020 3525.990 2077.020 3526.000 ;
        RECT 2254.020 3525.990 2257.020 3526.000 ;
        RECT 2434.020 3525.990 2437.020 3526.000 ;
        RECT 2614.020 3525.990 2617.020 3526.000 ;
        RECT 2794.020 3525.990 2797.020 3526.000 ;
        RECT 2931.300 3525.990 2934.300 3526.000 ;
        RECT -42.880 3396.380 -39.880 3396.390 ;
        RECT 148.020 3396.380 151.020 3396.390 ;
        RECT 328.020 3396.380 331.020 3396.390 ;
        RECT 508.020 3396.380 511.020 3396.390 ;
        RECT 688.020 3396.380 691.020 3396.390 ;
        RECT 868.020 3396.380 871.020 3396.390 ;
        RECT 1048.020 3396.380 1051.020 3396.390 ;
        RECT 1228.020 3396.380 1231.020 3396.390 ;
        RECT 1408.020 3396.380 1411.020 3396.390 ;
        RECT 1588.020 3396.380 1591.020 3396.390 ;
        RECT 1768.020 3396.380 1771.020 3396.390 ;
        RECT 1948.020 3396.380 1951.020 3396.390 ;
        RECT 2128.020 3396.380 2131.020 3396.390 ;
        RECT 2308.020 3396.380 2311.020 3396.390 ;
        RECT 2488.020 3396.380 2491.020 3396.390 ;
        RECT 2668.020 3396.380 2671.020 3396.390 ;
        RECT 2848.020 3396.380 2851.020 3396.390 ;
        RECT 2959.500 3396.380 2962.500 3396.390 ;
        RECT -42.880 3393.380 2962.500 3396.380 ;
        RECT -42.880 3393.370 -39.880 3393.380 ;
        RECT 148.020 3393.370 151.020 3393.380 ;
        RECT 328.020 3393.370 331.020 3393.380 ;
        RECT 508.020 3393.370 511.020 3393.380 ;
        RECT 688.020 3393.370 691.020 3393.380 ;
        RECT 868.020 3393.370 871.020 3393.380 ;
        RECT 1048.020 3393.370 1051.020 3393.380 ;
        RECT 1228.020 3393.370 1231.020 3393.380 ;
        RECT 1408.020 3393.370 1411.020 3393.380 ;
        RECT 1588.020 3393.370 1591.020 3393.380 ;
        RECT 1768.020 3393.370 1771.020 3393.380 ;
        RECT 1948.020 3393.370 1951.020 3393.380 ;
        RECT 2128.020 3393.370 2131.020 3393.380 ;
        RECT 2308.020 3393.370 2311.020 3393.380 ;
        RECT 2488.020 3393.370 2491.020 3393.380 ;
        RECT 2668.020 3393.370 2671.020 3393.380 ;
        RECT 2848.020 3393.370 2851.020 3393.380 ;
        RECT 2959.500 3393.370 2962.500 3393.380 ;
        RECT -33.480 3378.380 -30.480 3378.390 ;
        RECT 130.020 3378.380 133.020 3378.390 ;
        RECT 310.020 3378.380 313.020 3378.390 ;
        RECT 490.020 3378.380 493.020 3378.390 ;
        RECT 670.020 3378.380 673.020 3378.390 ;
        RECT 850.020 3378.380 853.020 3378.390 ;
        RECT 1030.020 3378.380 1033.020 3378.390 ;
        RECT 1210.020 3378.380 1213.020 3378.390 ;
        RECT 1390.020 3378.380 1393.020 3378.390 ;
        RECT 1570.020 3378.380 1573.020 3378.390 ;
        RECT 1750.020 3378.380 1753.020 3378.390 ;
        RECT 1930.020 3378.380 1933.020 3378.390 ;
        RECT 2110.020 3378.380 2113.020 3378.390 ;
        RECT 2290.020 3378.380 2293.020 3378.390 ;
        RECT 2470.020 3378.380 2473.020 3378.390 ;
        RECT 2650.020 3378.380 2653.020 3378.390 ;
        RECT 2830.020 3378.380 2833.020 3378.390 ;
        RECT 2950.100 3378.380 2953.100 3378.390 ;
        RECT -33.480 3375.380 2953.100 3378.380 ;
        RECT -33.480 3375.370 -30.480 3375.380 ;
        RECT 130.020 3375.370 133.020 3375.380 ;
        RECT 310.020 3375.370 313.020 3375.380 ;
        RECT 490.020 3375.370 493.020 3375.380 ;
        RECT 670.020 3375.370 673.020 3375.380 ;
        RECT 850.020 3375.370 853.020 3375.380 ;
        RECT 1030.020 3375.370 1033.020 3375.380 ;
        RECT 1210.020 3375.370 1213.020 3375.380 ;
        RECT 1390.020 3375.370 1393.020 3375.380 ;
        RECT 1570.020 3375.370 1573.020 3375.380 ;
        RECT 1750.020 3375.370 1753.020 3375.380 ;
        RECT 1930.020 3375.370 1933.020 3375.380 ;
        RECT 2110.020 3375.370 2113.020 3375.380 ;
        RECT 2290.020 3375.370 2293.020 3375.380 ;
        RECT 2470.020 3375.370 2473.020 3375.380 ;
        RECT 2650.020 3375.370 2653.020 3375.380 ;
        RECT 2830.020 3375.370 2833.020 3375.380 ;
        RECT 2950.100 3375.370 2953.100 3375.380 ;
        RECT -24.080 3360.380 -21.080 3360.390 ;
        RECT 112.020 3360.380 115.020 3360.390 ;
        RECT 292.020 3360.380 295.020 3360.390 ;
        RECT 472.020 3360.380 475.020 3360.390 ;
        RECT 652.020 3360.380 655.020 3360.390 ;
        RECT 832.020 3360.380 835.020 3360.390 ;
        RECT 1012.020 3360.380 1015.020 3360.390 ;
        RECT 1192.020 3360.380 1195.020 3360.390 ;
        RECT 1372.020 3360.380 1375.020 3360.390 ;
        RECT 1552.020 3360.380 1555.020 3360.390 ;
        RECT 1732.020 3360.380 1735.020 3360.390 ;
        RECT 1912.020 3360.380 1915.020 3360.390 ;
        RECT 2092.020 3360.380 2095.020 3360.390 ;
        RECT 2272.020 3360.380 2275.020 3360.390 ;
        RECT 2452.020 3360.380 2455.020 3360.390 ;
        RECT 2632.020 3360.380 2635.020 3360.390 ;
        RECT 2812.020 3360.380 2815.020 3360.390 ;
        RECT 2940.700 3360.380 2943.700 3360.390 ;
        RECT -24.080 3357.380 2943.700 3360.380 ;
        RECT -24.080 3357.370 -21.080 3357.380 ;
        RECT 112.020 3357.370 115.020 3357.380 ;
        RECT 292.020 3357.370 295.020 3357.380 ;
        RECT 472.020 3357.370 475.020 3357.380 ;
        RECT 652.020 3357.370 655.020 3357.380 ;
        RECT 832.020 3357.370 835.020 3357.380 ;
        RECT 1012.020 3357.370 1015.020 3357.380 ;
        RECT 1192.020 3357.370 1195.020 3357.380 ;
        RECT 1372.020 3357.370 1375.020 3357.380 ;
        RECT 1552.020 3357.370 1555.020 3357.380 ;
        RECT 1732.020 3357.370 1735.020 3357.380 ;
        RECT 1912.020 3357.370 1915.020 3357.380 ;
        RECT 2092.020 3357.370 2095.020 3357.380 ;
        RECT 2272.020 3357.370 2275.020 3357.380 ;
        RECT 2452.020 3357.370 2455.020 3357.380 ;
        RECT 2632.020 3357.370 2635.020 3357.380 ;
        RECT 2812.020 3357.370 2815.020 3357.380 ;
        RECT 2940.700 3357.370 2943.700 3357.380 ;
        RECT -14.680 3342.380 -11.680 3342.390 ;
        RECT 94.020 3342.380 97.020 3342.390 ;
        RECT 274.020 3342.380 277.020 3342.390 ;
        RECT 454.020 3342.380 457.020 3342.390 ;
        RECT 634.020 3342.380 637.020 3342.390 ;
        RECT 814.020 3342.380 817.020 3342.390 ;
        RECT 994.020 3342.380 997.020 3342.390 ;
        RECT 1174.020 3342.380 1177.020 3342.390 ;
        RECT 1354.020 3342.380 1357.020 3342.390 ;
        RECT 1534.020 3342.380 1537.020 3342.390 ;
        RECT 1714.020 3342.380 1717.020 3342.390 ;
        RECT 1894.020 3342.380 1897.020 3342.390 ;
        RECT 2074.020 3342.380 2077.020 3342.390 ;
        RECT 2254.020 3342.380 2257.020 3342.390 ;
        RECT 2434.020 3342.380 2437.020 3342.390 ;
        RECT 2614.020 3342.380 2617.020 3342.390 ;
        RECT 2794.020 3342.380 2797.020 3342.390 ;
        RECT 2931.300 3342.380 2934.300 3342.390 ;
        RECT -14.680 3339.380 2934.300 3342.380 ;
        RECT -14.680 3339.370 -11.680 3339.380 ;
        RECT 94.020 3339.370 97.020 3339.380 ;
        RECT 274.020 3339.370 277.020 3339.380 ;
        RECT 454.020 3339.370 457.020 3339.380 ;
        RECT 634.020 3339.370 637.020 3339.380 ;
        RECT 814.020 3339.370 817.020 3339.380 ;
        RECT 994.020 3339.370 997.020 3339.380 ;
        RECT 1174.020 3339.370 1177.020 3339.380 ;
        RECT 1354.020 3339.370 1357.020 3339.380 ;
        RECT 1534.020 3339.370 1537.020 3339.380 ;
        RECT 1714.020 3339.370 1717.020 3339.380 ;
        RECT 1894.020 3339.370 1897.020 3339.380 ;
        RECT 2074.020 3339.370 2077.020 3339.380 ;
        RECT 2254.020 3339.370 2257.020 3339.380 ;
        RECT 2434.020 3339.370 2437.020 3339.380 ;
        RECT 2614.020 3339.370 2617.020 3339.380 ;
        RECT 2794.020 3339.370 2797.020 3339.380 ;
        RECT 2931.300 3339.370 2934.300 3339.380 ;
        RECT -42.880 3216.380 -39.880 3216.390 ;
        RECT 148.020 3216.380 151.020 3216.390 ;
        RECT 684.690 3216.380 686.310 3216.390 ;
        RECT 868.020 3216.380 871.020 3216.390 ;
        RECT 1334.690 3216.380 1336.310 3216.390 ;
        RECT 1408.020 3216.380 1411.020 3216.390 ;
        RECT 1934.690 3216.380 1936.310 3216.390 ;
        RECT 2128.020 3216.380 2131.020 3216.390 ;
        RECT 2584.690 3216.380 2586.310 3216.390 ;
        RECT 2668.020 3216.380 2671.020 3216.390 ;
        RECT 2848.020 3216.380 2851.020 3216.390 ;
        RECT 2959.500 3216.380 2962.500 3216.390 ;
        RECT -42.880 3213.380 2962.500 3216.380 ;
        RECT -42.880 3213.370 -39.880 3213.380 ;
        RECT 148.020 3213.370 151.020 3213.380 ;
        RECT 684.690 3213.370 686.310 3213.380 ;
        RECT 868.020 3213.370 871.020 3213.380 ;
        RECT 1334.690 3213.370 1336.310 3213.380 ;
        RECT 1408.020 3213.370 1411.020 3213.380 ;
        RECT 1934.690 3213.370 1936.310 3213.380 ;
        RECT 2128.020 3213.370 2131.020 3213.380 ;
        RECT 2584.690 3213.370 2586.310 3213.380 ;
        RECT 2668.020 3213.370 2671.020 3213.380 ;
        RECT 2848.020 3213.370 2851.020 3213.380 ;
        RECT 2959.500 3213.370 2962.500 3213.380 ;
        RECT -33.480 3198.380 -30.480 3198.390 ;
        RECT 130.020 3198.380 133.020 3198.390 ;
        RECT 684.690 3198.380 686.310 3198.390 ;
        RECT 850.020 3198.380 853.020 3198.390 ;
        RECT 1334.690 3198.380 1336.310 3198.390 ;
        RECT 1390.020 3198.380 1393.020 3198.390 ;
        RECT 1934.690 3198.380 1936.310 3198.390 ;
        RECT 2110.020 3198.380 2113.020 3198.390 ;
        RECT 2584.690 3198.380 2586.310 3198.390 ;
        RECT 2650.020 3198.380 2653.020 3198.390 ;
        RECT 2830.020 3198.380 2833.020 3198.390 ;
        RECT 2950.100 3198.380 2953.100 3198.390 ;
        RECT -33.480 3195.380 2953.100 3198.380 ;
        RECT -33.480 3195.370 -30.480 3195.380 ;
        RECT 130.020 3195.370 133.020 3195.380 ;
        RECT 684.690 3195.370 686.310 3195.380 ;
        RECT 850.020 3195.370 853.020 3195.380 ;
        RECT 1334.690 3195.370 1336.310 3195.380 ;
        RECT 1390.020 3195.370 1393.020 3195.380 ;
        RECT 1934.690 3195.370 1936.310 3195.380 ;
        RECT 2110.020 3195.370 2113.020 3195.380 ;
        RECT 2584.690 3195.370 2586.310 3195.380 ;
        RECT 2650.020 3195.370 2653.020 3195.380 ;
        RECT 2830.020 3195.370 2833.020 3195.380 ;
        RECT 2950.100 3195.370 2953.100 3195.380 ;
        RECT -24.080 3180.380 -21.080 3180.390 ;
        RECT 112.020 3180.380 115.020 3180.390 ;
        RECT 684.690 3180.380 686.310 3180.390 ;
        RECT 832.020 3180.380 835.020 3180.390 ;
        RECT 1334.690 3180.380 1336.310 3180.390 ;
        RECT 1372.020 3180.380 1375.020 3180.390 ;
        RECT 1934.690 3180.380 1936.310 3180.390 ;
        RECT 2092.020 3180.380 2095.020 3180.390 ;
        RECT 2584.690 3180.380 2586.310 3180.390 ;
        RECT 2632.020 3180.380 2635.020 3180.390 ;
        RECT 2812.020 3180.380 2815.020 3180.390 ;
        RECT 2940.700 3180.380 2943.700 3180.390 ;
        RECT -24.080 3177.380 2943.700 3180.380 ;
        RECT -24.080 3177.370 -21.080 3177.380 ;
        RECT 112.020 3177.370 115.020 3177.380 ;
        RECT 684.690 3177.370 686.310 3177.380 ;
        RECT 832.020 3177.370 835.020 3177.380 ;
        RECT 1334.690 3177.370 1336.310 3177.380 ;
        RECT 1372.020 3177.370 1375.020 3177.380 ;
        RECT 1934.690 3177.370 1936.310 3177.380 ;
        RECT 2092.020 3177.370 2095.020 3177.380 ;
        RECT 2584.690 3177.370 2586.310 3177.380 ;
        RECT 2632.020 3177.370 2635.020 3177.380 ;
        RECT 2812.020 3177.370 2815.020 3177.380 ;
        RECT 2940.700 3177.370 2943.700 3177.380 ;
        RECT -14.680 3162.380 -11.680 3162.390 ;
        RECT 94.020 3162.380 97.020 3162.390 ;
        RECT 274.020 3162.380 277.020 3162.390 ;
        RECT 684.690 3162.380 686.310 3162.390 ;
        RECT 814.020 3162.380 817.020 3162.390 ;
        RECT 1334.690 3162.380 1336.310 3162.390 ;
        RECT 1354.020 3162.380 1357.020 3162.390 ;
        RECT 1934.690 3162.380 1936.310 3162.390 ;
        RECT 2074.020 3162.380 2077.020 3162.390 ;
        RECT 2584.690 3162.380 2586.310 3162.390 ;
        RECT 2614.020 3162.380 2617.020 3162.390 ;
        RECT 2794.020 3162.380 2797.020 3162.390 ;
        RECT 2931.300 3162.380 2934.300 3162.390 ;
        RECT -14.680 3159.380 2934.300 3162.380 ;
        RECT -14.680 3159.370 -11.680 3159.380 ;
        RECT 94.020 3159.370 97.020 3159.380 ;
        RECT 274.020 3159.370 277.020 3159.380 ;
        RECT 684.690 3159.370 686.310 3159.380 ;
        RECT 814.020 3159.370 817.020 3159.380 ;
        RECT 1334.690 3159.370 1336.310 3159.380 ;
        RECT 1354.020 3159.370 1357.020 3159.380 ;
        RECT 1934.690 3159.370 1936.310 3159.380 ;
        RECT 2074.020 3159.370 2077.020 3159.380 ;
        RECT 2584.690 3159.370 2586.310 3159.380 ;
        RECT 2614.020 3159.370 2617.020 3159.380 ;
        RECT 2794.020 3159.370 2797.020 3159.380 ;
        RECT 2931.300 3159.370 2934.300 3159.380 ;
        RECT -42.880 3036.380 -39.880 3036.390 ;
        RECT 148.020 3036.380 151.020 3036.390 ;
        RECT 684.690 3036.380 686.310 3036.390 ;
        RECT 868.020 3036.380 871.020 3036.390 ;
        RECT 1334.690 3036.380 1336.310 3036.390 ;
        RECT 1408.020 3036.380 1411.020 3036.390 ;
        RECT 1934.690 3036.380 1936.310 3036.390 ;
        RECT 2128.020 3036.380 2131.020 3036.390 ;
        RECT 2584.690 3036.380 2586.310 3036.390 ;
        RECT 2668.020 3036.380 2671.020 3036.390 ;
        RECT 2848.020 3036.380 2851.020 3036.390 ;
        RECT 2959.500 3036.380 2962.500 3036.390 ;
        RECT -42.880 3033.380 2962.500 3036.380 ;
        RECT -42.880 3033.370 -39.880 3033.380 ;
        RECT 148.020 3033.370 151.020 3033.380 ;
        RECT 684.690 3033.370 686.310 3033.380 ;
        RECT 868.020 3033.370 871.020 3033.380 ;
        RECT 1334.690 3033.370 1336.310 3033.380 ;
        RECT 1408.020 3033.370 1411.020 3033.380 ;
        RECT 1934.690 3033.370 1936.310 3033.380 ;
        RECT 2128.020 3033.370 2131.020 3033.380 ;
        RECT 2584.690 3033.370 2586.310 3033.380 ;
        RECT 2668.020 3033.370 2671.020 3033.380 ;
        RECT 2848.020 3033.370 2851.020 3033.380 ;
        RECT 2959.500 3033.370 2962.500 3033.380 ;
        RECT -33.480 3018.380 -30.480 3018.390 ;
        RECT 130.020 3018.380 133.020 3018.390 ;
        RECT 684.690 3018.380 686.310 3018.390 ;
        RECT 850.020 3018.380 853.020 3018.390 ;
        RECT 1334.690 3018.380 1336.310 3018.390 ;
        RECT 1390.020 3018.380 1393.020 3018.390 ;
        RECT 1934.690 3018.380 1936.310 3018.390 ;
        RECT 2110.020 3018.380 2113.020 3018.390 ;
        RECT 2584.690 3018.380 2586.310 3018.390 ;
        RECT 2650.020 3018.380 2653.020 3018.390 ;
        RECT 2830.020 3018.380 2833.020 3018.390 ;
        RECT 2950.100 3018.380 2953.100 3018.390 ;
        RECT -33.480 3015.380 2953.100 3018.380 ;
        RECT -33.480 3015.370 -30.480 3015.380 ;
        RECT 130.020 3015.370 133.020 3015.380 ;
        RECT 684.690 3015.370 686.310 3015.380 ;
        RECT 850.020 3015.370 853.020 3015.380 ;
        RECT 1334.690 3015.370 1336.310 3015.380 ;
        RECT 1390.020 3015.370 1393.020 3015.380 ;
        RECT 1934.690 3015.370 1936.310 3015.380 ;
        RECT 2110.020 3015.370 2113.020 3015.380 ;
        RECT 2584.690 3015.370 2586.310 3015.380 ;
        RECT 2650.020 3015.370 2653.020 3015.380 ;
        RECT 2830.020 3015.370 2833.020 3015.380 ;
        RECT 2950.100 3015.370 2953.100 3015.380 ;
        RECT -24.080 3000.380 -21.080 3000.390 ;
        RECT 112.020 3000.380 115.020 3000.390 ;
        RECT 684.690 3000.380 686.310 3000.390 ;
        RECT 832.020 3000.380 835.020 3000.390 ;
        RECT 1334.690 3000.380 1336.310 3000.390 ;
        RECT 1372.020 3000.380 1375.020 3000.390 ;
        RECT 1934.690 3000.380 1936.310 3000.390 ;
        RECT 2092.020 3000.380 2095.020 3000.390 ;
        RECT 2584.690 3000.380 2586.310 3000.390 ;
        RECT 2632.020 3000.380 2635.020 3000.390 ;
        RECT 2812.020 3000.380 2815.020 3000.390 ;
        RECT 2940.700 3000.380 2943.700 3000.390 ;
        RECT -24.080 2997.380 2943.700 3000.380 ;
        RECT -24.080 2997.370 -21.080 2997.380 ;
        RECT 112.020 2997.370 115.020 2997.380 ;
        RECT 684.690 2997.370 686.310 2997.380 ;
        RECT 832.020 2997.370 835.020 2997.380 ;
        RECT 1334.690 2997.370 1336.310 2997.380 ;
        RECT 1372.020 2997.370 1375.020 2997.380 ;
        RECT 1934.690 2997.370 1936.310 2997.380 ;
        RECT 2092.020 2997.370 2095.020 2997.380 ;
        RECT 2584.690 2997.370 2586.310 2997.380 ;
        RECT 2632.020 2997.370 2635.020 2997.380 ;
        RECT 2812.020 2997.370 2815.020 2997.380 ;
        RECT 2940.700 2997.370 2943.700 2997.380 ;
        RECT -14.680 2982.380 -11.680 2982.390 ;
        RECT 94.020 2982.380 97.020 2982.390 ;
        RECT 274.020 2982.380 277.020 2982.390 ;
        RECT 684.690 2982.380 686.310 2982.390 ;
        RECT 814.020 2982.380 817.020 2982.390 ;
        RECT 1334.690 2982.380 1336.310 2982.390 ;
        RECT 1354.020 2982.380 1357.020 2982.390 ;
        RECT 1934.690 2982.380 1936.310 2982.390 ;
        RECT 2074.020 2982.380 2077.020 2982.390 ;
        RECT 2584.690 2982.380 2586.310 2982.390 ;
        RECT 2614.020 2982.380 2617.020 2982.390 ;
        RECT 2794.020 2982.380 2797.020 2982.390 ;
        RECT 2931.300 2982.380 2934.300 2982.390 ;
        RECT -14.680 2979.380 2934.300 2982.380 ;
        RECT -14.680 2979.370 -11.680 2979.380 ;
        RECT 94.020 2979.370 97.020 2979.380 ;
        RECT 274.020 2979.370 277.020 2979.380 ;
        RECT 684.690 2979.370 686.310 2979.380 ;
        RECT 814.020 2979.370 817.020 2979.380 ;
        RECT 1334.690 2979.370 1336.310 2979.380 ;
        RECT 1354.020 2979.370 1357.020 2979.380 ;
        RECT 1934.690 2979.370 1936.310 2979.380 ;
        RECT 2074.020 2979.370 2077.020 2979.380 ;
        RECT 2584.690 2979.370 2586.310 2979.380 ;
        RECT 2614.020 2979.370 2617.020 2979.380 ;
        RECT 2794.020 2979.370 2797.020 2979.380 ;
        RECT 2931.300 2979.370 2934.300 2979.380 ;
        RECT -42.880 2856.380 -39.880 2856.390 ;
        RECT 148.020 2856.380 151.020 2856.390 ;
        RECT 684.690 2856.380 686.310 2856.390 ;
        RECT 868.020 2856.380 871.020 2856.390 ;
        RECT 1334.690 2856.380 1336.310 2856.390 ;
        RECT 1408.020 2856.380 1411.020 2856.390 ;
        RECT 1934.690 2856.380 1936.310 2856.390 ;
        RECT 2128.020 2856.380 2131.020 2856.390 ;
        RECT 2584.690 2856.380 2586.310 2856.390 ;
        RECT 2668.020 2856.380 2671.020 2856.390 ;
        RECT 2848.020 2856.380 2851.020 2856.390 ;
        RECT 2959.500 2856.380 2962.500 2856.390 ;
        RECT -42.880 2853.380 2962.500 2856.380 ;
        RECT -42.880 2853.370 -39.880 2853.380 ;
        RECT 148.020 2853.370 151.020 2853.380 ;
        RECT 684.690 2853.370 686.310 2853.380 ;
        RECT 868.020 2853.370 871.020 2853.380 ;
        RECT 1334.690 2853.370 1336.310 2853.380 ;
        RECT 1408.020 2853.370 1411.020 2853.380 ;
        RECT 1934.690 2853.370 1936.310 2853.380 ;
        RECT 2128.020 2853.370 2131.020 2853.380 ;
        RECT 2584.690 2853.370 2586.310 2853.380 ;
        RECT 2668.020 2853.370 2671.020 2853.380 ;
        RECT 2848.020 2853.370 2851.020 2853.380 ;
        RECT 2959.500 2853.370 2962.500 2853.380 ;
        RECT -33.480 2838.380 -30.480 2838.390 ;
        RECT 130.020 2838.380 133.020 2838.390 ;
        RECT 684.690 2838.380 686.310 2838.390 ;
        RECT 850.020 2838.380 853.020 2838.390 ;
        RECT 1334.690 2838.380 1336.310 2838.390 ;
        RECT 1390.020 2838.380 1393.020 2838.390 ;
        RECT 1934.690 2838.380 1936.310 2838.390 ;
        RECT 2110.020 2838.380 2113.020 2838.390 ;
        RECT 2584.690 2838.380 2586.310 2838.390 ;
        RECT 2650.020 2838.380 2653.020 2838.390 ;
        RECT 2830.020 2838.380 2833.020 2838.390 ;
        RECT 2950.100 2838.380 2953.100 2838.390 ;
        RECT -33.480 2835.380 2953.100 2838.380 ;
        RECT -33.480 2835.370 -30.480 2835.380 ;
        RECT 130.020 2835.370 133.020 2835.380 ;
        RECT 684.690 2835.370 686.310 2835.380 ;
        RECT 850.020 2835.370 853.020 2835.380 ;
        RECT 1334.690 2835.370 1336.310 2835.380 ;
        RECT 1390.020 2835.370 1393.020 2835.380 ;
        RECT 1934.690 2835.370 1936.310 2835.380 ;
        RECT 2110.020 2835.370 2113.020 2835.380 ;
        RECT 2584.690 2835.370 2586.310 2835.380 ;
        RECT 2650.020 2835.370 2653.020 2835.380 ;
        RECT 2830.020 2835.370 2833.020 2835.380 ;
        RECT 2950.100 2835.370 2953.100 2835.380 ;
        RECT -24.080 2820.380 -21.080 2820.390 ;
        RECT 112.020 2820.380 115.020 2820.390 ;
        RECT 684.690 2820.380 686.310 2820.390 ;
        RECT 832.020 2820.380 835.020 2820.390 ;
        RECT 1334.690 2820.380 1336.310 2820.390 ;
        RECT 1372.020 2820.380 1375.020 2820.390 ;
        RECT 1934.690 2820.380 1936.310 2820.390 ;
        RECT 2092.020 2820.380 2095.020 2820.390 ;
        RECT 2584.690 2820.380 2586.310 2820.390 ;
        RECT 2632.020 2820.380 2635.020 2820.390 ;
        RECT 2812.020 2820.380 2815.020 2820.390 ;
        RECT 2940.700 2820.380 2943.700 2820.390 ;
        RECT -24.080 2817.380 2943.700 2820.380 ;
        RECT -24.080 2817.370 -21.080 2817.380 ;
        RECT 112.020 2817.370 115.020 2817.380 ;
        RECT 684.690 2817.370 686.310 2817.380 ;
        RECT 832.020 2817.370 835.020 2817.380 ;
        RECT 1334.690 2817.370 1336.310 2817.380 ;
        RECT 1372.020 2817.370 1375.020 2817.380 ;
        RECT 1934.690 2817.370 1936.310 2817.380 ;
        RECT 2092.020 2817.370 2095.020 2817.380 ;
        RECT 2584.690 2817.370 2586.310 2817.380 ;
        RECT 2632.020 2817.370 2635.020 2817.380 ;
        RECT 2812.020 2817.370 2815.020 2817.380 ;
        RECT 2940.700 2817.370 2943.700 2817.380 ;
        RECT -14.680 2802.380 -11.680 2802.390 ;
        RECT 94.020 2802.380 97.020 2802.390 ;
        RECT 274.020 2802.380 277.020 2802.390 ;
        RECT 814.020 2802.380 817.020 2802.390 ;
        RECT 1354.020 2802.380 1357.020 2802.390 ;
        RECT 2074.020 2802.380 2077.020 2802.390 ;
        RECT 2614.020 2802.380 2617.020 2802.390 ;
        RECT 2794.020 2802.380 2797.020 2802.390 ;
        RECT 2931.300 2802.380 2934.300 2802.390 ;
        RECT -14.680 2799.380 2934.300 2802.380 ;
        RECT -14.680 2799.370 -11.680 2799.380 ;
        RECT 94.020 2799.370 97.020 2799.380 ;
        RECT 274.020 2799.370 277.020 2799.380 ;
        RECT 814.020 2799.370 817.020 2799.380 ;
        RECT 1354.020 2799.370 1357.020 2799.380 ;
        RECT 2074.020 2799.370 2077.020 2799.380 ;
        RECT 2614.020 2799.370 2617.020 2799.380 ;
        RECT 2794.020 2799.370 2797.020 2799.380 ;
        RECT 2931.300 2799.370 2934.300 2799.380 ;
        RECT -42.880 2676.380 -39.880 2676.390 ;
        RECT 148.020 2676.380 151.020 2676.390 ;
        RECT 397.840 2676.380 399.440 2676.390 ;
        RECT 1588.020 2676.380 1591.020 2676.390 ;
        RECT 1768.020 2676.380 1771.020 2676.390 ;
        RECT 1948.020 2676.380 1951.020 2676.390 ;
        RECT 2128.020 2676.380 2131.020 2676.390 ;
        RECT 2308.020 2676.380 2311.020 2676.390 ;
        RECT 2488.020 2676.380 2491.020 2676.390 ;
        RECT 2668.020 2676.380 2671.020 2676.390 ;
        RECT 2848.020 2676.380 2851.020 2676.390 ;
        RECT 2959.500 2676.380 2962.500 2676.390 ;
        RECT -42.880 2673.380 2962.500 2676.380 ;
        RECT -42.880 2673.370 -39.880 2673.380 ;
        RECT 148.020 2673.370 151.020 2673.380 ;
        RECT 397.840 2673.370 399.440 2673.380 ;
        RECT 1588.020 2673.370 1591.020 2673.380 ;
        RECT 1768.020 2673.370 1771.020 2673.380 ;
        RECT 1948.020 2673.370 1951.020 2673.380 ;
        RECT 2128.020 2673.370 2131.020 2673.380 ;
        RECT 2308.020 2673.370 2311.020 2673.380 ;
        RECT 2488.020 2673.370 2491.020 2673.380 ;
        RECT 2668.020 2673.370 2671.020 2673.380 ;
        RECT 2848.020 2673.370 2851.020 2673.380 ;
        RECT 2959.500 2673.370 2962.500 2673.380 ;
        RECT -33.480 2658.380 -30.480 2658.390 ;
        RECT 130.020 2658.380 133.020 2658.390 ;
        RECT 397.840 2658.380 399.440 2658.390 ;
        RECT 1570.020 2658.380 1573.020 2658.390 ;
        RECT 1750.020 2658.380 1753.020 2658.390 ;
        RECT 1930.020 2658.380 1933.020 2658.390 ;
        RECT 2110.020 2658.380 2113.020 2658.390 ;
        RECT 2290.020 2658.380 2293.020 2658.390 ;
        RECT 2470.020 2658.380 2473.020 2658.390 ;
        RECT 2650.020 2658.380 2653.020 2658.390 ;
        RECT 2830.020 2658.380 2833.020 2658.390 ;
        RECT 2950.100 2658.380 2953.100 2658.390 ;
        RECT -33.480 2655.380 2953.100 2658.380 ;
        RECT -33.480 2655.370 -30.480 2655.380 ;
        RECT 130.020 2655.370 133.020 2655.380 ;
        RECT 397.840 2655.370 399.440 2655.380 ;
        RECT 1570.020 2655.370 1573.020 2655.380 ;
        RECT 1750.020 2655.370 1753.020 2655.380 ;
        RECT 1930.020 2655.370 1933.020 2655.380 ;
        RECT 2110.020 2655.370 2113.020 2655.380 ;
        RECT 2290.020 2655.370 2293.020 2655.380 ;
        RECT 2470.020 2655.370 2473.020 2655.380 ;
        RECT 2650.020 2655.370 2653.020 2655.380 ;
        RECT 2830.020 2655.370 2833.020 2655.380 ;
        RECT 2950.100 2655.370 2953.100 2655.380 ;
        RECT -24.080 2640.380 -21.080 2640.390 ;
        RECT 112.020 2640.380 115.020 2640.390 ;
        RECT 397.840 2640.380 399.440 2640.390 ;
        RECT 1552.020 2640.380 1555.020 2640.390 ;
        RECT 1732.020 2640.380 1735.020 2640.390 ;
        RECT 1912.020 2640.380 1915.020 2640.390 ;
        RECT 2092.020 2640.380 2095.020 2640.390 ;
        RECT 2272.020 2640.380 2275.020 2640.390 ;
        RECT 2452.020 2640.380 2455.020 2640.390 ;
        RECT 2632.020 2640.380 2635.020 2640.390 ;
        RECT 2812.020 2640.380 2815.020 2640.390 ;
        RECT 2940.700 2640.380 2943.700 2640.390 ;
        RECT -24.080 2637.380 2943.700 2640.380 ;
        RECT -24.080 2637.370 -21.080 2637.380 ;
        RECT 112.020 2637.370 115.020 2637.380 ;
        RECT 397.840 2637.370 399.440 2637.380 ;
        RECT 1552.020 2637.370 1555.020 2637.380 ;
        RECT 1732.020 2637.370 1735.020 2637.380 ;
        RECT 1912.020 2637.370 1915.020 2637.380 ;
        RECT 2092.020 2637.370 2095.020 2637.380 ;
        RECT 2272.020 2637.370 2275.020 2637.380 ;
        RECT 2452.020 2637.370 2455.020 2637.380 ;
        RECT 2632.020 2637.370 2635.020 2637.380 ;
        RECT 2812.020 2637.370 2815.020 2637.380 ;
        RECT 2940.700 2637.370 2943.700 2637.380 ;
        RECT -14.680 2622.380 -11.680 2622.390 ;
        RECT 94.020 2622.380 97.020 2622.390 ;
        RECT 274.020 2622.380 277.020 2622.390 ;
        RECT 397.840 2622.380 399.440 2622.390 ;
        RECT 1534.020 2622.380 1537.020 2622.390 ;
        RECT 1714.020 2622.380 1717.020 2622.390 ;
        RECT 1894.020 2622.380 1897.020 2622.390 ;
        RECT 2074.020 2622.380 2077.020 2622.390 ;
        RECT 2254.020 2622.380 2257.020 2622.390 ;
        RECT 2434.020 2622.380 2437.020 2622.390 ;
        RECT 2614.020 2622.380 2617.020 2622.390 ;
        RECT 2794.020 2622.380 2797.020 2622.390 ;
        RECT 2931.300 2622.380 2934.300 2622.390 ;
        RECT -14.680 2619.380 2934.300 2622.380 ;
        RECT -14.680 2619.370 -11.680 2619.380 ;
        RECT 94.020 2619.370 97.020 2619.380 ;
        RECT 274.020 2619.370 277.020 2619.380 ;
        RECT 397.840 2619.370 399.440 2619.380 ;
        RECT 1534.020 2619.370 1537.020 2619.380 ;
        RECT 1714.020 2619.370 1717.020 2619.380 ;
        RECT 1894.020 2619.370 1897.020 2619.380 ;
        RECT 2074.020 2619.370 2077.020 2619.380 ;
        RECT 2254.020 2619.370 2257.020 2619.380 ;
        RECT 2434.020 2619.370 2437.020 2619.380 ;
        RECT 2614.020 2619.370 2617.020 2619.380 ;
        RECT 2794.020 2619.370 2797.020 2619.380 ;
        RECT 2931.300 2619.370 2934.300 2619.380 ;
        RECT -42.880 2496.380 -39.880 2496.390 ;
        RECT 148.020 2496.380 151.020 2496.390 ;
        RECT 397.840 2496.380 399.440 2496.390 ;
        RECT 1588.020 2496.380 1591.020 2496.390 ;
        RECT 1768.020 2496.380 1771.020 2496.390 ;
        RECT 1948.020 2496.380 1951.020 2496.390 ;
        RECT 2128.020 2496.380 2131.020 2496.390 ;
        RECT 2308.020 2496.380 2311.020 2496.390 ;
        RECT 2488.020 2496.380 2491.020 2496.390 ;
        RECT 2668.020 2496.380 2671.020 2496.390 ;
        RECT 2848.020 2496.380 2851.020 2496.390 ;
        RECT 2959.500 2496.380 2962.500 2496.390 ;
        RECT -42.880 2493.380 2962.500 2496.380 ;
        RECT -42.880 2493.370 -39.880 2493.380 ;
        RECT 148.020 2493.370 151.020 2493.380 ;
        RECT 397.840 2493.370 399.440 2493.380 ;
        RECT 1588.020 2493.370 1591.020 2493.380 ;
        RECT 1768.020 2493.370 1771.020 2493.380 ;
        RECT 1948.020 2493.370 1951.020 2493.380 ;
        RECT 2128.020 2493.370 2131.020 2493.380 ;
        RECT 2308.020 2493.370 2311.020 2493.380 ;
        RECT 2488.020 2493.370 2491.020 2493.380 ;
        RECT 2668.020 2493.370 2671.020 2493.380 ;
        RECT 2848.020 2493.370 2851.020 2493.380 ;
        RECT 2959.500 2493.370 2962.500 2493.380 ;
        RECT -33.480 2478.380 -30.480 2478.390 ;
        RECT 130.020 2478.380 133.020 2478.390 ;
        RECT 397.840 2478.380 399.440 2478.390 ;
        RECT 1570.020 2478.380 1573.020 2478.390 ;
        RECT 1750.020 2478.380 1753.020 2478.390 ;
        RECT 1930.020 2478.380 1933.020 2478.390 ;
        RECT 2110.020 2478.380 2113.020 2478.390 ;
        RECT 2290.020 2478.380 2293.020 2478.390 ;
        RECT 2470.020 2478.380 2473.020 2478.390 ;
        RECT 2650.020 2478.380 2653.020 2478.390 ;
        RECT 2830.020 2478.380 2833.020 2478.390 ;
        RECT 2950.100 2478.380 2953.100 2478.390 ;
        RECT -33.480 2475.380 2953.100 2478.380 ;
        RECT -33.480 2475.370 -30.480 2475.380 ;
        RECT 130.020 2475.370 133.020 2475.380 ;
        RECT 397.840 2475.370 399.440 2475.380 ;
        RECT 1570.020 2475.370 1573.020 2475.380 ;
        RECT 1750.020 2475.370 1753.020 2475.380 ;
        RECT 1930.020 2475.370 1933.020 2475.380 ;
        RECT 2110.020 2475.370 2113.020 2475.380 ;
        RECT 2290.020 2475.370 2293.020 2475.380 ;
        RECT 2470.020 2475.370 2473.020 2475.380 ;
        RECT 2650.020 2475.370 2653.020 2475.380 ;
        RECT 2830.020 2475.370 2833.020 2475.380 ;
        RECT 2950.100 2475.370 2953.100 2475.380 ;
        RECT -24.080 2460.380 -21.080 2460.390 ;
        RECT 112.020 2460.380 115.020 2460.390 ;
        RECT 397.840 2460.380 399.440 2460.390 ;
        RECT 1552.020 2460.380 1555.020 2460.390 ;
        RECT 1732.020 2460.380 1735.020 2460.390 ;
        RECT 1912.020 2460.380 1915.020 2460.390 ;
        RECT 2092.020 2460.380 2095.020 2460.390 ;
        RECT 2272.020 2460.380 2275.020 2460.390 ;
        RECT 2452.020 2460.380 2455.020 2460.390 ;
        RECT 2632.020 2460.380 2635.020 2460.390 ;
        RECT 2812.020 2460.380 2815.020 2460.390 ;
        RECT 2940.700 2460.380 2943.700 2460.390 ;
        RECT -24.080 2457.380 2943.700 2460.380 ;
        RECT -24.080 2457.370 -21.080 2457.380 ;
        RECT 112.020 2457.370 115.020 2457.380 ;
        RECT 397.840 2457.370 399.440 2457.380 ;
        RECT 1552.020 2457.370 1555.020 2457.380 ;
        RECT 1732.020 2457.370 1735.020 2457.380 ;
        RECT 1912.020 2457.370 1915.020 2457.380 ;
        RECT 2092.020 2457.370 2095.020 2457.380 ;
        RECT 2272.020 2457.370 2275.020 2457.380 ;
        RECT 2452.020 2457.370 2455.020 2457.380 ;
        RECT 2632.020 2457.370 2635.020 2457.380 ;
        RECT 2812.020 2457.370 2815.020 2457.380 ;
        RECT 2940.700 2457.370 2943.700 2457.380 ;
        RECT -14.680 2442.380 -11.680 2442.390 ;
        RECT 94.020 2442.380 97.020 2442.390 ;
        RECT 274.020 2442.380 277.020 2442.390 ;
        RECT 397.840 2442.380 399.440 2442.390 ;
        RECT 1534.020 2442.380 1537.020 2442.390 ;
        RECT 1714.020 2442.380 1717.020 2442.390 ;
        RECT 1894.020 2442.380 1897.020 2442.390 ;
        RECT 2074.020 2442.380 2077.020 2442.390 ;
        RECT 2254.020 2442.380 2257.020 2442.390 ;
        RECT 2434.020 2442.380 2437.020 2442.390 ;
        RECT 2614.020 2442.380 2617.020 2442.390 ;
        RECT 2794.020 2442.380 2797.020 2442.390 ;
        RECT 2931.300 2442.380 2934.300 2442.390 ;
        RECT -14.680 2439.380 2934.300 2442.380 ;
        RECT -14.680 2439.370 -11.680 2439.380 ;
        RECT 94.020 2439.370 97.020 2439.380 ;
        RECT 274.020 2439.370 277.020 2439.380 ;
        RECT 397.840 2439.370 399.440 2439.380 ;
        RECT 1534.020 2439.370 1537.020 2439.380 ;
        RECT 1714.020 2439.370 1717.020 2439.380 ;
        RECT 1894.020 2439.370 1897.020 2439.380 ;
        RECT 2074.020 2439.370 2077.020 2439.380 ;
        RECT 2254.020 2439.370 2257.020 2439.380 ;
        RECT 2434.020 2439.370 2437.020 2439.380 ;
        RECT 2614.020 2439.370 2617.020 2439.380 ;
        RECT 2794.020 2439.370 2797.020 2439.380 ;
        RECT 2931.300 2439.370 2934.300 2439.380 ;
        RECT -42.880 2316.380 -39.880 2316.390 ;
        RECT 148.020 2316.380 151.020 2316.390 ;
        RECT 397.840 2316.380 399.440 2316.390 ;
        RECT 1588.020 2316.380 1591.020 2316.390 ;
        RECT 1768.020 2316.380 1771.020 2316.390 ;
        RECT 1948.020 2316.380 1951.020 2316.390 ;
        RECT 2128.020 2316.380 2131.020 2316.390 ;
        RECT 2308.020 2316.380 2311.020 2316.390 ;
        RECT 2488.020 2316.380 2491.020 2316.390 ;
        RECT 2668.020 2316.380 2671.020 2316.390 ;
        RECT 2848.020 2316.380 2851.020 2316.390 ;
        RECT 2959.500 2316.380 2962.500 2316.390 ;
        RECT -42.880 2313.380 2962.500 2316.380 ;
        RECT -42.880 2313.370 -39.880 2313.380 ;
        RECT 148.020 2313.370 151.020 2313.380 ;
        RECT 397.840 2313.370 399.440 2313.380 ;
        RECT 1588.020 2313.370 1591.020 2313.380 ;
        RECT 1768.020 2313.370 1771.020 2313.380 ;
        RECT 1948.020 2313.370 1951.020 2313.380 ;
        RECT 2128.020 2313.370 2131.020 2313.380 ;
        RECT 2308.020 2313.370 2311.020 2313.380 ;
        RECT 2488.020 2313.370 2491.020 2313.380 ;
        RECT 2668.020 2313.370 2671.020 2313.380 ;
        RECT 2848.020 2313.370 2851.020 2313.380 ;
        RECT 2959.500 2313.370 2962.500 2313.380 ;
        RECT -33.480 2298.380 -30.480 2298.390 ;
        RECT 130.020 2298.380 133.020 2298.390 ;
        RECT 397.840 2298.380 399.440 2298.390 ;
        RECT 1570.020 2298.380 1573.020 2298.390 ;
        RECT 1750.020 2298.380 1753.020 2298.390 ;
        RECT 1930.020 2298.380 1933.020 2298.390 ;
        RECT 2110.020 2298.380 2113.020 2298.390 ;
        RECT 2290.020 2298.380 2293.020 2298.390 ;
        RECT 2470.020 2298.380 2473.020 2298.390 ;
        RECT 2650.020 2298.380 2653.020 2298.390 ;
        RECT 2830.020 2298.380 2833.020 2298.390 ;
        RECT 2950.100 2298.380 2953.100 2298.390 ;
        RECT -33.480 2295.380 2953.100 2298.380 ;
        RECT -33.480 2295.370 -30.480 2295.380 ;
        RECT 130.020 2295.370 133.020 2295.380 ;
        RECT 397.840 2295.370 399.440 2295.380 ;
        RECT 1570.020 2295.370 1573.020 2295.380 ;
        RECT 1750.020 2295.370 1753.020 2295.380 ;
        RECT 1930.020 2295.370 1933.020 2295.380 ;
        RECT 2110.020 2295.370 2113.020 2295.380 ;
        RECT 2290.020 2295.370 2293.020 2295.380 ;
        RECT 2470.020 2295.370 2473.020 2295.380 ;
        RECT 2650.020 2295.370 2653.020 2295.380 ;
        RECT 2830.020 2295.370 2833.020 2295.380 ;
        RECT 2950.100 2295.370 2953.100 2295.380 ;
        RECT -24.080 2280.380 -21.080 2280.390 ;
        RECT 112.020 2280.380 115.020 2280.390 ;
        RECT 397.840 2280.380 399.440 2280.390 ;
        RECT 1552.020 2280.380 1555.020 2280.390 ;
        RECT 1732.020 2280.380 1735.020 2280.390 ;
        RECT 1912.020 2280.380 1915.020 2280.390 ;
        RECT 2092.020 2280.380 2095.020 2280.390 ;
        RECT 2272.020 2280.380 2275.020 2280.390 ;
        RECT 2452.020 2280.380 2455.020 2280.390 ;
        RECT 2632.020 2280.380 2635.020 2280.390 ;
        RECT 2812.020 2280.380 2815.020 2280.390 ;
        RECT 2940.700 2280.380 2943.700 2280.390 ;
        RECT -24.080 2277.380 2943.700 2280.380 ;
        RECT -24.080 2277.370 -21.080 2277.380 ;
        RECT 112.020 2277.370 115.020 2277.380 ;
        RECT 397.840 2277.370 399.440 2277.380 ;
        RECT 1552.020 2277.370 1555.020 2277.380 ;
        RECT 1732.020 2277.370 1735.020 2277.380 ;
        RECT 1912.020 2277.370 1915.020 2277.380 ;
        RECT 2092.020 2277.370 2095.020 2277.380 ;
        RECT 2272.020 2277.370 2275.020 2277.380 ;
        RECT 2452.020 2277.370 2455.020 2277.380 ;
        RECT 2632.020 2277.370 2635.020 2277.380 ;
        RECT 2812.020 2277.370 2815.020 2277.380 ;
        RECT 2940.700 2277.370 2943.700 2277.380 ;
        RECT -14.680 2262.380 -11.680 2262.390 ;
        RECT 94.020 2262.380 97.020 2262.390 ;
        RECT 274.020 2262.380 277.020 2262.390 ;
        RECT 397.840 2262.380 399.440 2262.390 ;
        RECT 1534.020 2262.380 1537.020 2262.390 ;
        RECT 1714.020 2262.380 1717.020 2262.390 ;
        RECT 1894.020 2262.380 1897.020 2262.390 ;
        RECT 2074.020 2262.380 2077.020 2262.390 ;
        RECT 2254.020 2262.380 2257.020 2262.390 ;
        RECT 2434.020 2262.380 2437.020 2262.390 ;
        RECT 2614.020 2262.380 2617.020 2262.390 ;
        RECT 2794.020 2262.380 2797.020 2262.390 ;
        RECT 2931.300 2262.380 2934.300 2262.390 ;
        RECT -14.680 2259.380 2934.300 2262.380 ;
        RECT -14.680 2259.370 -11.680 2259.380 ;
        RECT 94.020 2259.370 97.020 2259.380 ;
        RECT 274.020 2259.370 277.020 2259.380 ;
        RECT 397.840 2259.370 399.440 2259.380 ;
        RECT 1534.020 2259.370 1537.020 2259.380 ;
        RECT 1714.020 2259.370 1717.020 2259.380 ;
        RECT 1894.020 2259.370 1897.020 2259.380 ;
        RECT 2074.020 2259.370 2077.020 2259.380 ;
        RECT 2254.020 2259.370 2257.020 2259.380 ;
        RECT 2434.020 2259.370 2437.020 2259.380 ;
        RECT 2614.020 2259.370 2617.020 2259.380 ;
        RECT 2794.020 2259.370 2797.020 2259.380 ;
        RECT 2931.300 2259.370 2934.300 2259.380 ;
        RECT -42.880 2136.380 -39.880 2136.390 ;
        RECT 148.020 2136.380 151.020 2136.390 ;
        RECT 397.840 2136.380 399.440 2136.390 ;
        RECT 1588.020 2136.380 1591.020 2136.390 ;
        RECT 1768.020 2136.380 1771.020 2136.390 ;
        RECT 1948.020 2136.380 1951.020 2136.390 ;
        RECT 2128.020 2136.380 2131.020 2136.390 ;
        RECT 2308.020 2136.380 2311.020 2136.390 ;
        RECT 2488.020 2136.380 2491.020 2136.390 ;
        RECT 2668.020 2136.380 2671.020 2136.390 ;
        RECT 2848.020 2136.380 2851.020 2136.390 ;
        RECT 2959.500 2136.380 2962.500 2136.390 ;
        RECT -42.880 2133.380 2962.500 2136.380 ;
        RECT -42.880 2133.370 -39.880 2133.380 ;
        RECT 148.020 2133.370 151.020 2133.380 ;
        RECT 397.840 2133.370 399.440 2133.380 ;
        RECT 1588.020 2133.370 1591.020 2133.380 ;
        RECT 1768.020 2133.370 1771.020 2133.380 ;
        RECT 1948.020 2133.370 1951.020 2133.380 ;
        RECT 2128.020 2133.370 2131.020 2133.380 ;
        RECT 2308.020 2133.370 2311.020 2133.380 ;
        RECT 2488.020 2133.370 2491.020 2133.380 ;
        RECT 2668.020 2133.370 2671.020 2133.380 ;
        RECT 2848.020 2133.370 2851.020 2133.380 ;
        RECT 2959.500 2133.370 2962.500 2133.380 ;
        RECT -33.480 2118.380 -30.480 2118.390 ;
        RECT 130.020 2118.380 133.020 2118.390 ;
        RECT 397.840 2118.380 399.440 2118.390 ;
        RECT 1570.020 2118.380 1573.020 2118.390 ;
        RECT 1750.020 2118.380 1753.020 2118.390 ;
        RECT 1930.020 2118.380 1933.020 2118.390 ;
        RECT 2110.020 2118.380 2113.020 2118.390 ;
        RECT 2290.020 2118.380 2293.020 2118.390 ;
        RECT 2470.020 2118.380 2473.020 2118.390 ;
        RECT 2650.020 2118.380 2653.020 2118.390 ;
        RECT 2830.020 2118.380 2833.020 2118.390 ;
        RECT 2950.100 2118.380 2953.100 2118.390 ;
        RECT -33.480 2115.380 2953.100 2118.380 ;
        RECT -33.480 2115.370 -30.480 2115.380 ;
        RECT 130.020 2115.370 133.020 2115.380 ;
        RECT 397.840 2115.370 399.440 2115.380 ;
        RECT 1570.020 2115.370 1573.020 2115.380 ;
        RECT 1750.020 2115.370 1753.020 2115.380 ;
        RECT 1930.020 2115.370 1933.020 2115.380 ;
        RECT 2110.020 2115.370 2113.020 2115.380 ;
        RECT 2290.020 2115.370 2293.020 2115.380 ;
        RECT 2470.020 2115.370 2473.020 2115.380 ;
        RECT 2650.020 2115.370 2653.020 2115.380 ;
        RECT 2830.020 2115.370 2833.020 2115.380 ;
        RECT 2950.100 2115.370 2953.100 2115.380 ;
        RECT -24.080 2100.380 -21.080 2100.390 ;
        RECT 112.020 2100.380 115.020 2100.390 ;
        RECT 397.840 2100.380 399.440 2100.390 ;
        RECT 1552.020 2100.380 1555.020 2100.390 ;
        RECT 1732.020 2100.380 1735.020 2100.390 ;
        RECT 1912.020 2100.380 1915.020 2100.390 ;
        RECT 2092.020 2100.380 2095.020 2100.390 ;
        RECT 2272.020 2100.380 2275.020 2100.390 ;
        RECT 2452.020 2100.380 2455.020 2100.390 ;
        RECT 2632.020 2100.380 2635.020 2100.390 ;
        RECT 2812.020 2100.380 2815.020 2100.390 ;
        RECT 2940.700 2100.380 2943.700 2100.390 ;
        RECT -24.080 2097.380 2943.700 2100.380 ;
        RECT -24.080 2097.370 -21.080 2097.380 ;
        RECT 112.020 2097.370 115.020 2097.380 ;
        RECT 397.840 2097.370 399.440 2097.380 ;
        RECT 1552.020 2097.370 1555.020 2097.380 ;
        RECT 1732.020 2097.370 1735.020 2097.380 ;
        RECT 1912.020 2097.370 1915.020 2097.380 ;
        RECT 2092.020 2097.370 2095.020 2097.380 ;
        RECT 2272.020 2097.370 2275.020 2097.380 ;
        RECT 2452.020 2097.370 2455.020 2097.380 ;
        RECT 2632.020 2097.370 2635.020 2097.380 ;
        RECT 2812.020 2097.370 2815.020 2097.380 ;
        RECT 2940.700 2097.370 2943.700 2097.380 ;
        RECT -14.680 2082.380 -11.680 2082.390 ;
        RECT 94.020 2082.380 97.020 2082.390 ;
        RECT 274.020 2082.380 277.020 2082.390 ;
        RECT 397.840 2082.380 399.440 2082.390 ;
        RECT 1534.020 2082.380 1537.020 2082.390 ;
        RECT 1714.020 2082.380 1717.020 2082.390 ;
        RECT 1894.020 2082.380 1897.020 2082.390 ;
        RECT 2074.020 2082.380 2077.020 2082.390 ;
        RECT 2254.020 2082.380 2257.020 2082.390 ;
        RECT 2434.020 2082.380 2437.020 2082.390 ;
        RECT 2614.020 2082.380 2617.020 2082.390 ;
        RECT 2794.020 2082.380 2797.020 2082.390 ;
        RECT 2931.300 2082.380 2934.300 2082.390 ;
        RECT -14.680 2079.380 2934.300 2082.380 ;
        RECT -14.680 2079.370 -11.680 2079.380 ;
        RECT 94.020 2079.370 97.020 2079.380 ;
        RECT 274.020 2079.370 277.020 2079.380 ;
        RECT 397.840 2079.370 399.440 2079.380 ;
        RECT 1534.020 2079.370 1537.020 2079.380 ;
        RECT 1714.020 2079.370 1717.020 2079.380 ;
        RECT 1894.020 2079.370 1897.020 2079.380 ;
        RECT 2074.020 2079.370 2077.020 2079.380 ;
        RECT 2254.020 2079.370 2257.020 2079.380 ;
        RECT 2434.020 2079.370 2437.020 2079.380 ;
        RECT 2614.020 2079.370 2617.020 2079.380 ;
        RECT 2794.020 2079.370 2797.020 2079.380 ;
        RECT 2931.300 2079.370 2934.300 2079.380 ;
        RECT -42.880 1956.380 -39.880 1956.390 ;
        RECT 148.020 1956.380 151.020 1956.390 ;
        RECT 397.840 1956.380 399.440 1956.390 ;
        RECT 1588.020 1956.380 1591.020 1956.390 ;
        RECT 1768.020 1956.380 1771.020 1956.390 ;
        RECT 1948.020 1956.380 1951.020 1956.390 ;
        RECT 2128.020 1956.380 2131.020 1956.390 ;
        RECT 2308.020 1956.380 2311.020 1956.390 ;
        RECT 2488.020 1956.380 2491.020 1956.390 ;
        RECT 2668.020 1956.380 2671.020 1956.390 ;
        RECT 2848.020 1956.380 2851.020 1956.390 ;
        RECT 2959.500 1956.380 2962.500 1956.390 ;
        RECT -42.880 1953.380 2962.500 1956.380 ;
        RECT -42.880 1953.370 -39.880 1953.380 ;
        RECT 148.020 1953.370 151.020 1953.380 ;
        RECT 397.840 1953.370 399.440 1953.380 ;
        RECT 1588.020 1953.370 1591.020 1953.380 ;
        RECT 1768.020 1953.370 1771.020 1953.380 ;
        RECT 1948.020 1953.370 1951.020 1953.380 ;
        RECT 2128.020 1953.370 2131.020 1953.380 ;
        RECT 2308.020 1953.370 2311.020 1953.380 ;
        RECT 2488.020 1953.370 2491.020 1953.380 ;
        RECT 2668.020 1953.370 2671.020 1953.380 ;
        RECT 2848.020 1953.370 2851.020 1953.380 ;
        RECT 2959.500 1953.370 2962.500 1953.380 ;
        RECT -33.480 1938.380 -30.480 1938.390 ;
        RECT 130.020 1938.380 133.020 1938.390 ;
        RECT 397.840 1938.380 399.440 1938.390 ;
        RECT 1570.020 1938.380 1573.020 1938.390 ;
        RECT 1750.020 1938.380 1753.020 1938.390 ;
        RECT 1930.020 1938.380 1933.020 1938.390 ;
        RECT 2110.020 1938.380 2113.020 1938.390 ;
        RECT 2290.020 1938.380 2293.020 1938.390 ;
        RECT 2470.020 1938.380 2473.020 1938.390 ;
        RECT 2650.020 1938.380 2653.020 1938.390 ;
        RECT 2830.020 1938.380 2833.020 1938.390 ;
        RECT 2950.100 1938.380 2953.100 1938.390 ;
        RECT -33.480 1935.380 2953.100 1938.380 ;
        RECT -33.480 1935.370 -30.480 1935.380 ;
        RECT 130.020 1935.370 133.020 1935.380 ;
        RECT 397.840 1935.370 399.440 1935.380 ;
        RECT 1570.020 1935.370 1573.020 1935.380 ;
        RECT 1750.020 1935.370 1753.020 1935.380 ;
        RECT 1930.020 1935.370 1933.020 1935.380 ;
        RECT 2110.020 1935.370 2113.020 1935.380 ;
        RECT 2290.020 1935.370 2293.020 1935.380 ;
        RECT 2470.020 1935.370 2473.020 1935.380 ;
        RECT 2650.020 1935.370 2653.020 1935.380 ;
        RECT 2830.020 1935.370 2833.020 1935.380 ;
        RECT 2950.100 1935.370 2953.100 1935.380 ;
        RECT -24.080 1920.380 -21.080 1920.390 ;
        RECT 112.020 1920.380 115.020 1920.390 ;
        RECT 397.840 1920.380 399.440 1920.390 ;
        RECT 1552.020 1920.380 1555.020 1920.390 ;
        RECT 1732.020 1920.380 1735.020 1920.390 ;
        RECT 1912.020 1920.380 1915.020 1920.390 ;
        RECT 2092.020 1920.380 2095.020 1920.390 ;
        RECT 2272.020 1920.380 2275.020 1920.390 ;
        RECT 2452.020 1920.380 2455.020 1920.390 ;
        RECT 2632.020 1920.380 2635.020 1920.390 ;
        RECT 2812.020 1920.380 2815.020 1920.390 ;
        RECT 2940.700 1920.380 2943.700 1920.390 ;
        RECT -24.080 1917.380 2943.700 1920.380 ;
        RECT -24.080 1917.370 -21.080 1917.380 ;
        RECT 112.020 1917.370 115.020 1917.380 ;
        RECT 397.840 1917.370 399.440 1917.380 ;
        RECT 1552.020 1917.370 1555.020 1917.380 ;
        RECT 1732.020 1917.370 1735.020 1917.380 ;
        RECT 1912.020 1917.370 1915.020 1917.380 ;
        RECT 2092.020 1917.370 2095.020 1917.380 ;
        RECT 2272.020 1917.370 2275.020 1917.380 ;
        RECT 2452.020 1917.370 2455.020 1917.380 ;
        RECT 2632.020 1917.370 2635.020 1917.380 ;
        RECT 2812.020 1917.370 2815.020 1917.380 ;
        RECT 2940.700 1917.370 2943.700 1917.380 ;
        RECT -14.680 1902.380 -11.680 1902.390 ;
        RECT 94.020 1902.380 97.020 1902.390 ;
        RECT 274.020 1902.380 277.020 1902.390 ;
        RECT 397.840 1902.380 399.440 1902.390 ;
        RECT 1534.020 1902.380 1537.020 1902.390 ;
        RECT 1714.020 1902.380 1717.020 1902.390 ;
        RECT 1894.020 1902.380 1897.020 1902.390 ;
        RECT 2074.020 1902.380 2077.020 1902.390 ;
        RECT 2254.020 1902.380 2257.020 1902.390 ;
        RECT 2434.020 1902.380 2437.020 1902.390 ;
        RECT 2614.020 1902.380 2617.020 1902.390 ;
        RECT 2794.020 1902.380 2797.020 1902.390 ;
        RECT 2931.300 1902.380 2934.300 1902.390 ;
        RECT -14.680 1899.380 2934.300 1902.380 ;
        RECT -14.680 1899.370 -11.680 1899.380 ;
        RECT 94.020 1899.370 97.020 1899.380 ;
        RECT 274.020 1899.370 277.020 1899.380 ;
        RECT 397.840 1899.370 399.440 1899.380 ;
        RECT 1534.020 1899.370 1537.020 1899.380 ;
        RECT 1714.020 1899.370 1717.020 1899.380 ;
        RECT 1894.020 1899.370 1897.020 1899.380 ;
        RECT 2074.020 1899.370 2077.020 1899.380 ;
        RECT 2254.020 1899.370 2257.020 1899.380 ;
        RECT 2434.020 1899.370 2437.020 1899.380 ;
        RECT 2614.020 1899.370 2617.020 1899.380 ;
        RECT 2794.020 1899.370 2797.020 1899.380 ;
        RECT 2931.300 1899.370 2934.300 1899.380 ;
        RECT -42.880 1776.380 -39.880 1776.390 ;
        RECT 148.020 1776.380 151.020 1776.390 ;
        RECT 397.840 1776.380 399.440 1776.390 ;
        RECT 1588.020 1776.380 1591.020 1776.390 ;
        RECT 1768.020 1776.380 1771.020 1776.390 ;
        RECT 1948.020 1776.380 1951.020 1776.390 ;
        RECT 2128.020 1776.380 2131.020 1776.390 ;
        RECT 2308.020 1776.380 2311.020 1776.390 ;
        RECT 2488.020 1776.380 2491.020 1776.390 ;
        RECT 2668.020 1776.380 2671.020 1776.390 ;
        RECT 2848.020 1776.380 2851.020 1776.390 ;
        RECT 2959.500 1776.380 2962.500 1776.390 ;
        RECT -42.880 1773.380 2962.500 1776.380 ;
        RECT -42.880 1773.370 -39.880 1773.380 ;
        RECT 148.020 1773.370 151.020 1773.380 ;
        RECT 397.840 1773.370 399.440 1773.380 ;
        RECT 1588.020 1773.370 1591.020 1773.380 ;
        RECT 1768.020 1773.370 1771.020 1773.380 ;
        RECT 1948.020 1773.370 1951.020 1773.380 ;
        RECT 2128.020 1773.370 2131.020 1773.380 ;
        RECT 2308.020 1773.370 2311.020 1773.380 ;
        RECT 2488.020 1773.370 2491.020 1773.380 ;
        RECT 2668.020 1773.370 2671.020 1773.380 ;
        RECT 2848.020 1773.370 2851.020 1773.380 ;
        RECT 2959.500 1773.370 2962.500 1773.380 ;
        RECT -33.480 1758.380 -30.480 1758.390 ;
        RECT 130.020 1758.380 133.020 1758.390 ;
        RECT 397.840 1758.380 399.440 1758.390 ;
        RECT 1570.020 1758.380 1573.020 1758.390 ;
        RECT 1750.020 1758.380 1753.020 1758.390 ;
        RECT 1930.020 1758.380 1933.020 1758.390 ;
        RECT 2110.020 1758.380 2113.020 1758.390 ;
        RECT 2290.020 1758.380 2293.020 1758.390 ;
        RECT 2470.020 1758.380 2473.020 1758.390 ;
        RECT 2650.020 1758.380 2653.020 1758.390 ;
        RECT 2830.020 1758.380 2833.020 1758.390 ;
        RECT 2950.100 1758.380 2953.100 1758.390 ;
        RECT -33.480 1755.380 2953.100 1758.380 ;
        RECT -33.480 1755.370 -30.480 1755.380 ;
        RECT 130.020 1755.370 133.020 1755.380 ;
        RECT 397.840 1755.370 399.440 1755.380 ;
        RECT 1570.020 1755.370 1573.020 1755.380 ;
        RECT 1750.020 1755.370 1753.020 1755.380 ;
        RECT 1930.020 1755.370 1933.020 1755.380 ;
        RECT 2110.020 1755.370 2113.020 1755.380 ;
        RECT 2290.020 1755.370 2293.020 1755.380 ;
        RECT 2470.020 1755.370 2473.020 1755.380 ;
        RECT 2650.020 1755.370 2653.020 1755.380 ;
        RECT 2830.020 1755.370 2833.020 1755.380 ;
        RECT 2950.100 1755.370 2953.100 1755.380 ;
        RECT -24.080 1740.380 -21.080 1740.390 ;
        RECT 112.020 1740.380 115.020 1740.390 ;
        RECT 397.840 1740.380 399.440 1740.390 ;
        RECT 1552.020 1740.380 1555.020 1740.390 ;
        RECT 1732.020 1740.380 1735.020 1740.390 ;
        RECT 1912.020 1740.380 1915.020 1740.390 ;
        RECT 2092.020 1740.380 2095.020 1740.390 ;
        RECT 2272.020 1740.380 2275.020 1740.390 ;
        RECT 2452.020 1740.380 2455.020 1740.390 ;
        RECT 2632.020 1740.380 2635.020 1740.390 ;
        RECT 2812.020 1740.380 2815.020 1740.390 ;
        RECT 2940.700 1740.380 2943.700 1740.390 ;
        RECT -24.080 1737.380 2943.700 1740.380 ;
        RECT -24.080 1737.370 -21.080 1737.380 ;
        RECT 112.020 1737.370 115.020 1737.380 ;
        RECT 397.840 1737.370 399.440 1737.380 ;
        RECT 1552.020 1737.370 1555.020 1737.380 ;
        RECT 1732.020 1737.370 1735.020 1737.380 ;
        RECT 1912.020 1737.370 1915.020 1737.380 ;
        RECT 2092.020 1737.370 2095.020 1737.380 ;
        RECT 2272.020 1737.370 2275.020 1737.380 ;
        RECT 2452.020 1737.370 2455.020 1737.380 ;
        RECT 2632.020 1737.370 2635.020 1737.380 ;
        RECT 2812.020 1737.370 2815.020 1737.380 ;
        RECT 2940.700 1737.370 2943.700 1737.380 ;
        RECT -14.680 1722.380 -11.680 1722.390 ;
        RECT 94.020 1722.380 97.020 1722.390 ;
        RECT 274.020 1722.380 277.020 1722.390 ;
        RECT 397.840 1722.380 399.440 1722.390 ;
        RECT 1534.020 1722.380 1537.020 1722.390 ;
        RECT 1714.020 1722.380 1717.020 1722.390 ;
        RECT 1894.020 1722.380 1897.020 1722.390 ;
        RECT 2074.020 1722.380 2077.020 1722.390 ;
        RECT 2254.020 1722.380 2257.020 1722.390 ;
        RECT 2434.020 1722.380 2437.020 1722.390 ;
        RECT 2614.020 1722.380 2617.020 1722.390 ;
        RECT 2794.020 1722.380 2797.020 1722.390 ;
        RECT 2931.300 1722.380 2934.300 1722.390 ;
        RECT -14.680 1719.380 2934.300 1722.380 ;
        RECT -14.680 1719.370 -11.680 1719.380 ;
        RECT 94.020 1719.370 97.020 1719.380 ;
        RECT 274.020 1719.370 277.020 1719.380 ;
        RECT 397.840 1719.370 399.440 1719.380 ;
        RECT 1534.020 1719.370 1537.020 1719.380 ;
        RECT 1714.020 1719.370 1717.020 1719.380 ;
        RECT 1894.020 1719.370 1897.020 1719.380 ;
        RECT 2074.020 1719.370 2077.020 1719.380 ;
        RECT 2254.020 1719.370 2257.020 1719.380 ;
        RECT 2434.020 1719.370 2437.020 1719.380 ;
        RECT 2614.020 1719.370 2617.020 1719.380 ;
        RECT 2794.020 1719.370 2797.020 1719.380 ;
        RECT 2931.300 1719.370 2934.300 1719.380 ;
        RECT -42.880 1596.380 -39.880 1596.390 ;
        RECT 148.020 1596.380 151.020 1596.390 ;
        RECT 397.840 1596.380 399.440 1596.390 ;
        RECT 1588.020 1596.380 1591.020 1596.390 ;
        RECT 1768.020 1596.380 1771.020 1596.390 ;
        RECT 1948.020 1596.380 1951.020 1596.390 ;
        RECT 2128.020 1596.380 2131.020 1596.390 ;
        RECT 2308.020 1596.380 2311.020 1596.390 ;
        RECT 2488.020 1596.380 2491.020 1596.390 ;
        RECT 2668.020 1596.380 2671.020 1596.390 ;
        RECT 2848.020 1596.380 2851.020 1596.390 ;
        RECT 2959.500 1596.380 2962.500 1596.390 ;
        RECT -42.880 1593.380 2962.500 1596.380 ;
        RECT -42.880 1593.370 -39.880 1593.380 ;
        RECT 148.020 1593.370 151.020 1593.380 ;
        RECT 397.840 1593.370 399.440 1593.380 ;
        RECT 1588.020 1593.370 1591.020 1593.380 ;
        RECT 1768.020 1593.370 1771.020 1593.380 ;
        RECT 1948.020 1593.370 1951.020 1593.380 ;
        RECT 2128.020 1593.370 2131.020 1593.380 ;
        RECT 2308.020 1593.370 2311.020 1593.380 ;
        RECT 2488.020 1593.370 2491.020 1593.380 ;
        RECT 2668.020 1593.370 2671.020 1593.380 ;
        RECT 2848.020 1593.370 2851.020 1593.380 ;
        RECT 2959.500 1593.370 2962.500 1593.380 ;
        RECT -33.480 1578.380 -30.480 1578.390 ;
        RECT 130.020 1578.380 133.020 1578.390 ;
        RECT 397.840 1578.380 399.440 1578.390 ;
        RECT 1570.020 1578.380 1573.020 1578.390 ;
        RECT 1750.020 1578.380 1753.020 1578.390 ;
        RECT 1930.020 1578.380 1933.020 1578.390 ;
        RECT 2110.020 1578.380 2113.020 1578.390 ;
        RECT 2290.020 1578.380 2293.020 1578.390 ;
        RECT 2470.020 1578.380 2473.020 1578.390 ;
        RECT 2650.020 1578.380 2653.020 1578.390 ;
        RECT 2830.020 1578.380 2833.020 1578.390 ;
        RECT 2950.100 1578.380 2953.100 1578.390 ;
        RECT -33.480 1575.380 2953.100 1578.380 ;
        RECT -33.480 1575.370 -30.480 1575.380 ;
        RECT 130.020 1575.370 133.020 1575.380 ;
        RECT 397.840 1575.370 399.440 1575.380 ;
        RECT 1570.020 1575.370 1573.020 1575.380 ;
        RECT 1750.020 1575.370 1753.020 1575.380 ;
        RECT 1930.020 1575.370 1933.020 1575.380 ;
        RECT 2110.020 1575.370 2113.020 1575.380 ;
        RECT 2290.020 1575.370 2293.020 1575.380 ;
        RECT 2470.020 1575.370 2473.020 1575.380 ;
        RECT 2650.020 1575.370 2653.020 1575.380 ;
        RECT 2830.020 1575.370 2833.020 1575.380 ;
        RECT 2950.100 1575.370 2953.100 1575.380 ;
        RECT -24.080 1560.380 -21.080 1560.390 ;
        RECT 112.020 1560.380 115.020 1560.390 ;
        RECT 397.840 1560.380 399.440 1560.390 ;
        RECT 1552.020 1560.380 1555.020 1560.390 ;
        RECT 1732.020 1560.380 1735.020 1560.390 ;
        RECT 1912.020 1560.380 1915.020 1560.390 ;
        RECT 2092.020 1560.380 2095.020 1560.390 ;
        RECT 2272.020 1560.380 2275.020 1560.390 ;
        RECT 2452.020 1560.380 2455.020 1560.390 ;
        RECT 2632.020 1560.380 2635.020 1560.390 ;
        RECT 2812.020 1560.380 2815.020 1560.390 ;
        RECT 2940.700 1560.380 2943.700 1560.390 ;
        RECT -24.080 1557.380 2943.700 1560.380 ;
        RECT -24.080 1557.370 -21.080 1557.380 ;
        RECT 112.020 1557.370 115.020 1557.380 ;
        RECT 397.840 1557.370 399.440 1557.380 ;
        RECT 1552.020 1557.370 1555.020 1557.380 ;
        RECT 1732.020 1557.370 1735.020 1557.380 ;
        RECT 1912.020 1557.370 1915.020 1557.380 ;
        RECT 2092.020 1557.370 2095.020 1557.380 ;
        RECT 2272.020 1557.370 2275.020 1557.380 ;
        RECT 2452.020 1557.370 2455.020 1557.380 ;
        RECT 2632.020 1557.370 2635.020 1557.380 ;
        RECT 2812.020 1557.370 2815.020 1557.380 ;
        RECT 2940.700 1557.370 2943.700 1557.380 ;
        RECT -14.680 1542.380 -11.680 1542.390 ;
        RECT 94.020 1542.380 97.020 1542.390 ;
        RECT 274.020 1542.380 277.020 1542.390 ;
        RECT 397.840 1542.380 399.440 1542.390 ;
        RECT 1534.020 1542.380 1537.020 1542.390 ;
        RECT 1714.020 1542.380 1717.020 1542.390 ;
        RECT 1894.020 1542.380 1897.020 1542.390 ;
        RECT 2074.020 1542.380 2077.020 1542.390 ;
        RECT 2254.020 1542.380 2257.020 1542.390 ;
        RECT 2434.020 1542.380 2437.020 1542.390 ;
        RECT 2614.020 1542.380 2617.020 1542.390 ;
        RECT 2794.020 1542.380 2797.020 1542.390 ;
        RECT 2931.300 1542.380 2934.300 1542.390 ;
        RECT -14.680 1539.380 2934.300 1542.380 ;
        RECT -14.680 1539.370 -11.680 1539.380 ;
        RECT 94.020 1539.370 97.020 1539.380 ;
        RECT 274.020 1539.370 277.020 1539.380 ;
        RECT 397.840 1539.370 399.440 1539.380 ;
        RECT 1534.020 1539.370 1537.020 1539.380 ;
        RECT 1714.020 1539.370 1717.020 1539.380 ;
        RECT 1894.020 1539.370 1897.020 1539.380 ;
        RECT 2074.020 1539.370 2077.020 1539.380 ;
        RECT 2254.020 1539.370 2257.020 1539.380 ;
        RECT 2434.020 1539.370 2437.020 1539.380 ;
        RECT 2614.020 1539.370 2617.020 1539.380 ;
        RECT 2794.020 1539.370 2797.020 1539.380 ;
        RECT 2931.300 1539.370 2934.300 1539.380 ;
        RECT -42.880 1416.380 -39.880 1416.390 ;
        RECT 148.020 1416.380 151.020 1416.390 ;
        RECT 328.020 1416.380 331.020 1416.390 ;
        RECT 508.020 1416.380 511.020 1416.390 ;
        RECT 688.020 1416.380 691.020 1416.390 ;
        RECT 868.020 1416.380 871.020 1416.390 ;
        RECT 1048.020 1416.380 1051.020 1416.390 ;
        RECT 1228.020 1416.380 1231.020 1416.390 ;
        RECT 1408.020 1416.380 1411.020 1416.390 ;
        RECT 1588.020 1416.380 1591.020 1416.390 ;
        RECT 1768.020 1416.380 1771.020 1416.390 ;
        RECT 1948.020 1416.380 1951.020 1416.390 ;
        RECT 2128.020 1416.380 2131.020 1416.390 ;
        RECT 2308.020 1416.380 2311.020 1416.390 ;
        RECT 2488.020 1416.380 2491.020 1416.390 ;
        RECT 2668.020 1416.380 2671.020 1416.390 ;
        RECT 2848.020 1416.380 2851.020 1416.390 ;
        RECT 2959.500 1416.380 2962.500 1416.390 ;
        RECT -42.880 1413.380 2962.500 1416.380 ;
        RECT -42.880 1413.370 -39.880 1413.380 ;
        RECT 148.020 1413.370 151.020 1413.380 ;
        RECT 328.020 1413.370 331.020 1413.380 ;
        RECT 508.020 1413.370 511.020 1413.380 ;
        RECT 688.020 1413.370 691.020 1413.380 ;
        RECT 868.020 1413.370 871.020 1413.380 ;
        RECT 1048.020 1413.370 1051.020 1413.380 ;
        RECT 1228.020 1413.370 1231.020 1413.380 ;
        RECT 1408.020 1413.370 1411.020 1413.380 ;
        RECT 1588.020 1413.370 1591.020 1413.380 ;
        RECT 1768.020 1413.370 1771.020 1413.380 ;
        RECT 1948.020 1413.370 1951.020 1413.380 ;
        RECT 2128.020 1413.370 2131.020 1413.380 ;
        RECT 2308.020 1413.370 2311.020 1413.380 ;
        RECT 2488.020 1413.370 2491.020 1413.380 ;
        RECT 2668.020 1413.370 2671.020 1413.380 ;
        RECT 2848.020 1413.370 2851.020 1413.380 ;
        RECT 2959.500 1413.370 2962.500 1413.380 ;
        RECT -33.480 1398.380 -30.480 1398.390 ;
        RECT 130.020 1398.380 133.020 1398.390 ;
        RECT 310.020 1398.380 313.020 1398.390 ;
        RECT 490.020 1398.380 493.020 1398.390 ;
        RECT 670.020 1398.380 673.020 1398.390 ;
        RECT 850.020 1398.380 853.020 1398.390 ;
        RECT 1030.020 1398.380 1033.020 1398.390 ;
        RECT 1210.020 1398.380 1213.020 1398.390 ;
        RECT 1390.020 1398.380 1393.020 1398.390 ;
        RECT 1570.020 1398.380 1573.020 1398.390 ;
        RECT 1750.020 1398.380 1753.020 1398.390 ;
        RECT 1930.020 1398.380 1933.020 1398.390 ;
        RECT 2110.020 1398.380 2113.020 1398.390 ;
        RECT 2290.020 1398.380 2293.020 1398.390 ;
        RECT 2470.020 1398.380 2473.020 1398.390 ;
        RECT 2650.020 1398.380 2653.020 1398.390 ;
        RECT 2830.020 1398.380 2833.020 1398.390 ;
        RECT 2950.100 1398.380 2953.100 1398.390 ;
        RECT -33.480 1395.380 2953.100 1398.380 ;
        RECT -33.480 1395.370 -30.480 1395.380 ;
        RECT 130.020 1395.370 133.020 1395.380 ;
        RECT 310.020 1395.370 313.020 1395.380 ;
        RECT 490.020 1395.370 493.020 1395.380 ;
        RECT 670.020 1395.370 673.020 1395.380 ;
        RECT 850.020 1395.370 853.020 1395.380 ;
        RECT 1030.020 1395.370 1033.020 1395.380 ;
        RECT 1210.020 1395.370 1213.020 1395.380 ;
        RECT 1390.020 1395.370 1393.020 1395.380 ;
        RECT 1570.020 1395.370 1573.020 1395.380 ;
        RECT 1750.020 1395.370 1753.020 1395.380 ;
        RECT 1930.020 1395.370 1933.020 1395.380 ;
        RECT 2110.020 1395.370 2113.020 1395.380 ;
        RECT 2290.020 1395.370 2293.020 1395.380 ;
        RECT 2470.020 1395.370 2473.020 1395.380 ;
        RECT 2650.020 1395.370 2653.020 1395.380 ;
        RECT 2830.020 1395.370 2833.020 1395.380 ;
        RECT 2950.100 1395.370 2953.100 1395.380 ;
        RECT -24.080 1380.380 -21.080 1380.390 ;
        RECT 112.020 1380.380 115.020 1380.390 ;
        RECT 292.020 1380.380 295.020 1380.390 ;
        RECT 472.020 1380.380 475.020 1380.390 ;
        RECT 652.020 1380.380 655.020 1380.390 ;
        RECT 832.020 1380.380 835.020 1380.390 ;
        RECT 1012.020 1380.380 1015.020 1380.390 ;
        RECT 1192.020 1380.380 1195.020 1380.390 ;
        RECT 1372.020 1380.380 1375.020 1380.390 ;
        RECT 1552.020 1380.380 1555.020 1380.390 ;
        RECT 1732.020 1380.380 1735.020 1380.390 ;
        RECT 1912.020 1380.380 1915.020 1380.390 ;
        RECT 2092.020 1380.380 2095.020 1380.390 ;
        RECT 2272.020 1380.380 2275.020 1380.390 ;
        RECT 2452.020 1380.380 2455.020 1380.390 ;
        RECT 2632.020 1380.380 2635.020 1380.390 ;
        RECT 2812.020 1380.380 2815.020 1380.390 ;
        RECT 2940.700 1380.380 2943.700 1380.390 ;
        RECT -24.080 1377.380 2943.700 1380.380 ;
        RECT -24.080 1377.370 -21.080 1377.380 ;
        RECT 112.020 1377.370 115.020 1377.380 ;
        RECT 292.020 1377.370 295.020 1377.380 ;
        RECT 472.020 1377.370 475.020 1377.380 ;
        RECT 652.020 1377.370 655.020 1377.380 ;
        RECT 832.020 1377.370 835.020 1377.380 ;
        RECT 1012.020 1377.370 1015.020 1377.380 ;
        RECT 1192.020 1377.370 1195.020 1377.380 ;
        RECT 1372.020 1377.370 1375.020 1377.380 ;
        RECT 1552.020 1377.370 1555.020 1377.380 ;
        RECT 1732.020 1377.370 1735.020 1377.380 ;
        RECT 1912.020 1377.370 1915.020 1377.380 ;
        RECT 2092.020 1377.370 2095.020 1377.380 ;
        RECT 2272.020 1377.370 2275.020 1377.380 ;
        RECT 2452.020 1377.370 2455.020 1377.380 ;
        RECT 2632.020 1377.370 2635.020 1377.380 ;
        RECT 2812.020 1377.370 2815.020 1377.380 ;
        RECT 2940.700 1377.370 2943.700 1377.380 ;
        RECT -14.680 1362.380 -11.680 1362.390 ;
        RECT 94.020 1362.380 97.020 1362.390 ;
        RECT 274.020 1362.380 277.020 1362.390 ;
        RECT 454.020 1362.380 457.020 1362.390 ;
        RECT 634.020 1362.380 637.020 1362.390 ;
        RECT 814.020 1362.380 817.020 1362.390 ;
        RECT 994.020 1362.380 997.020 1362.390 ;
        RECT 1174.020 1362.380 1177.020 1362.390 ;
        RECT 1354.020 1362.380 1357.020 1362.390 ;
        RECT 1534.020 1362.380 1537.020 1362.390 ;
        RECT 1714.020 1362.380 1717.020 1362.390 ;
        RECT 1894.020 1362.380 1897.020 1362.390 ;
        RECT 2074.020 1362.380 2077.020 1362.390 ;
        RECT 2254.020 1362.380 2257.020 1362.390 ;
        RECT 2434.020 1362.380 2437.020 1362.390 ;
        RECT 2614.020 1362.380 2617.020 1362.390 ;
        RECT 2794.020 1362.380 2797.020 1362.390 ;
        RECT 2931.300 1362.380 2934.300 1362.390 ;
        RECT -14.680 1359.380 2934.300 1362.380 ;
        RECT -14.680 1359.370 -11.680 1359.380 ;
        RECT 94.020 1359.370 97.020 1359.380 ;
        RECT 274.020 1359.370 277.020 1359.380 ;
        RECT 454.020 1359.370 457.020 1359.380 ;
        RECT 634.020 1359.370 637.020 1359.380 ;
        RECT 814.020 1359.370 817.020 1359.380 ;
        RECT 994.020 1359.370 997.020 1359.380 ;
        RECT 1174.020 1359.370 1177.020 1359.380 ;
        RECT 1354.020 1359.370 1357.020 1359.380 ;
        RECT 1534.020 1359.370 1537.020 1359.380 ;
        RECT 1714.020 1359.370 1717.020 1359.380 ;
        RECT 1894.020 1359.370 1897.020 1359.380 ;
        RECT 2074.020 1359.370 2077.020 1359.380 ;
        RECT 2254.020 1359.370 2257.020 1359.380 ;
        RECT 2434.020 1359.370 2437.020 1359.380 ;
        RECT 2614.020 1359.370 2617.020 1359.380 ;
        RECT 2794.020 1359.370 2797.020 1359.380 ;
        RECT 2931.300 1359.370 2934.300 1359.380 ;
        RECT -42.880 1236.380 -39.880 1236.390 ;
        RECT 148.020 1236.380 151.020 1236.390 ;
        RECT 328.020 1236.380 331.020 1236.390 ;
        RECT 508.020 1236.380 511.020 1236.390 ;
        RECT 688.020 1236.380 691.020 1236.390 ;
        RECT 868.020 1236.380 871.020 1236.390 ;
        RECT 1048.020 1236.380 1051.020 1236.390 ;
        RECT 1228.020 1236.380 1231.020 1236.390 ;
        RECT 1408.020 1236.380 1411.020 1236.390 ;
        RECT 1588.020 1236.380 1591.020 1236.390 ;
        RECT 1768.020 1236.380 1771.020 1236.390 ;
        RECT 1948.020 1236.380 1951.020 1236.390 ;
        RECT 2128.020 1236.380 2131.020 1236.390 ;
        RECT 2308.020 1236.380 2311.020 1236.390 ;
        RECT 2488.020 1236.380 2491.020 1236.390 ;
        RECT 2668.020 1236.380 2671.020 1236.390 ;
        RECT 2848.020 1236.380 2851.020 1236.390 ;
        RECT 2959.500 1236.380 2962.500 1236.390 ;
        RECT -42.880 1233.380 2962.500 1236.380 ;
        RECT -42.880 1233.370 -39.880 1233.380 ;
        RECT 148.020 1233.370 151.020 1233.380 ;
        RECT 328.020 1233.370 331.020 1233.380 ;
        RECT 508.020 1233.370 511.020 1233.380 ;
        RECT 688.020 1233.370 691.020 1233.380 ;
        RECT 868.020 1233.370 871.020 1233.380 ;
        RECT 1048.020 1233.370 1051.020 1233.380 ;
        RECT 1228.020 1233.370 1231.020 1233.380 ;
        RECT 1408.020 1233.370 1411.020 1233.380 ;
        RECT 1588.020 1233.370 1591.020 1233.380 ;
        RECT 1768.020 1233.370 1771.020 1233.380 ;
        RECT 1948.020 1233.370 1951.020 1233.380 ;
        RECT 2128.020 1233.370 2131.020 1233.380 ;
        RECT 2308.020 1233.370 2311.020 1233.380 ;
        RECT 2488.020 1233.370 2491.020 1233.380 ;
        RECT 2668.020 1233.370 2671.020 1233.380 ;
        RECT 2848.020 1233.370 2851.020 1233.380 ;
        RECT 2959.500 1233.370 2962.500 1233.380 ;
        RECT -33.480 1218.380 -30.480 1218.390 ;
        RECT 130.020 1218.380 133.020 1218.390 ;
        RECT 310.020 1218.380 313.020 1218.390 ;
        RECT 490.020 1218.380 493.020 1218.390 ;
        RECT 670.020 1218.380 673.020 1218.390 ;
        RECT 850.020 1218.380 853.020 1218.390 ;
        RECT 1030.020 1218.380 1033.020 1218.390 ;
        RECT 1210.020 1218.380 1213.020 1218.390 ;
        RECT 1390.020 1218.380 1393.020 1218.390 ;
        RECT 1570.020 1218.380 1573.020 1218.390 ;
        RECT 1750.020 1218.380 1753.020 1218.390 ;
        RECT 1930.020 1218.380 1933.020 1218.390 ;
        RECT 2110.020 1218.380 2113.020 1218.390 ;
        RECT 2290.020 1218.380 2293.020 1218.390 ;
        RECT 2470.020 1218.380 2473.020 1218.390 ;
        RECT 2650.020 1218.380 2653.020 1218.390 ;
        RECT 2830.020 1218.380 2833.020 1218.390 ;
        RECT 2950.100 1218.380 2953.100 1218.390 ;
        RECT -33.480 1215.380 2953.100 1218.380 ;
        RECT -33.480 1215.370 -30.480 1215.380 ;
        RECT 130.020 1215.370 133.020 1215.380 ;
        RECT 310.020 1215.370 313.020 1215.380 ;
        RECT 490.020 1215.370 493.020 1215.380 ;
        RECT 670.020 1215.370 673.020 1215.380 ;
        RECT 850.020 1215.370 853.020 1215.380 ;
        RECT 1030.020 1215.370 1033.020 1215.380 ;
        RECT 1210.020 1215.370 1213.020 1215.380 ;
        RECT 1390.020 1215.370 1393.020 1215.380 ;
        RECT 1570.020 1215.370 1573.020 1215.380 ;
        RECT 1750.020 1215.370 1753.020 1215.380 ;
        RECT 1930.020 1215.370 1933.020 1215.380 ;
        RECT 2110.020 1215.370 2113.020 1215.380 ;
        RECT 2290.020 1215.370 2293.020 1215.380 ;
        RECT 2470.020 1215.370 2473.020 1215.380 ;
        RECT 2650.020 1215.370 2653.020 1215.380 ;
        RECT 2830.020 1215.370 2833.020 1215.380 ;
        RECT 2950.100 1215.370 2953.100 1215.380 ;
        RECT -24.080 1200.380 -21.080 1200.390 ;
        RECT 112.020 1200.380 115.020 1200.390 ;
        RECT 292.020 1200.380 295.020 1200.390 ;
        RECT 472.020 1200.380 475.020 1200.390 ;
        RECT 652.020 1200.380 655.020 1200.390 ;
        RECT 832.020 1200.380 835.020 1200.390 ;
        RECT 1012.020 1200.380 1015.020 1200.390 ;
        RECT 1192.020 1200.380 1195.020 1200.390 ;
        RECT 1372.020 1200.380 1375.020 1200.390 ;
        RECT 1552.020 1200.380 1555.020 1200.390 ;
        RECT 1732.020 1200.380 1735.020 1200.390 ;
        RECT 1912.020 1200.380 1915.020 1200.390 ;
        RECT 2092.020 1200.380 2095.020 1200.390 ;
        RECT 2272.020 1200.380 2275.020 1200.390 ;
        RECT 2452.020 1200.380 2455.020 1200.390 ;
        RECT 2632.020 1200.380 2635.020 1200.390 ;
        RECT 2812.020 1200.380 2815.020 1200.390 ;
        RECT 2940.700 1200.380 2943.700 1200.390 ;
        RECT -24.080 1197.380 2943.700 1200.380 ;
        RECT -24.080 1197.370 -21.080 1197.380 ;
        RECT 112.020 1197.370 115.020 1197.380 ;
        RECT 292.020 1197.370 295.020 1197.380 ;
        RECT 472.020 1197.370 475.020 1197.380 ;
        RECT 652.020 1197.370 655.020 1197.380 ;
        RECT 832.020 1197.370 835.020 1197.380 ;
        RECT 1012.020 1197.370 1015.020 1197.380 ;
        RECT 1192.020 1197.370 1195.020 1197.380 ;
        RECT 1372.020 1197.370 1375.020 1197.380 ;
        RECT 1552.020 1197.370 1555.020 1197.380 ;
        RECT 1732.020 1197.370 1735.020 1197.380 ;
        RECT 1912.020 1197.370 1915.020 1197.380 ;
        RECT 2092.020 1197.370 2095.020 1197.380 ;
        RECT 2272.020 1197.370 2275.020 1197.380 ;
        RECT 2452.020 1197.370 2455.020 1197.380 ;
        RECT 2632.020 1197.370 2635.020 1197.380 ;
        RECT 2812.020 1197.370 2815.020 1197.380 ;
        RECT 2940.700 1197.370 2943.700 1197.380 ;
        RECT -14.680 1182.380 -11.680 1182.390 ;
        RECT 94.020 1182.380 97.020 1182.390 ;
        RECT 274.020 1182.380 277.020 1182.390 ;
        RECT 454.020 1182.380 457.020 1182.390 ;
        RECT 634.020 1182.380 637.020 1182.390 ;
        RECT 814.020 1182.380 817.020 1182.390 ;
        RECT 994.020 1182.380 997.020 1182.390 ;
        RECT 1174.020 1182.380 1177.020 1182.390 ;
        RECT 1354.020 1182.380 1357.020 1182.390 ;
        RECT 1534.020 1182.380 1537.020 1182.390 ;
        RECT 1714.020 1182.380 1717.020 1182.390 ;
        RECT 1894.020 1182.380 1897.020 1182.390 ;
        RECT 2074.020 1182.380 2077.020 1182.390 ;
        RECT 2254.020 1182.380 2257.020 1182.390 ;
        RECT 2434.020 1182.380 2437.020 1182.390 ;
        RECT 2614.020 1182.380 2617.020 1182.390 ;
        RECT 2794.020 1182.380 2797.020 1182.390 ;
        RECT 2931.300 1182.380 2934.300 1182.390 ;
        RECT -14.680 1179.380 2934.300 1182.380 ;
        RECT -14.680 1179.370 -11.680 1179.380 ;
        RECT 94.020 1179.370 97.020 1179.380 ;
        RECT 274.020 1179.370 277.020 1179.380 ;
        RECT 454.020 1179.370 457.020 1179.380 ;
        RECT 634.020 1179.370 637.020 1179.380 ;
        RECT 814.020 1179.370 817.020 1179.380 ;
        RECT 994.020 1179.370 997.020 1179.380 ;
        RECT 1174.020 1179.370 1177.020 1179.380 ;
        RECT 1354.020 1179.370 1357.020 1179.380 ;
        RECT 1534.020 1179.370 1537.020 1179.380 ;
        RECT 1714.020 1179.370 1717.020 1179.380 ;
        RECT 1894.020 1179.370 1897.020 1179.380 ;
        RECT 2074.020 1179.370 2077.020 1179.380 ;
        RECT 2254.020 1179.370 2257.020 1179.380 ;
        RECT 2434.020 1179.370 2437.020 1179.380 ;
        RECT 2614.020 1179.370 2617.020 1179.380 ;
        RECT 2794.020 1179.370 2797.020 1179.380 ;
        RECT 2931.300 1179.370 2934.300 1179.380 ;
        RECT -42.880 1056.380 -39.880 1056.390 ;
        RECT 148.020 1056.380 151.020 1056.390 ;
        RECT 328.020 1056.380 331.020 1056.390 ;
        RECT 508.020 1056.380 511.020 1056.390 ;
        RECT 688.020 1056.380 691.020 1056.390 ;
        RECT 868.020 1056.380 871.020 1056.390 ;
        RECT 1048.020 1056.380 1051.020 1056.390 ;
        RECT 1228.020 1056.380 1231.020 1056.390 ;
        RECT 1408.020 1056.380 1411.020 1056.390 ;
        RECT 1588.020 1056.380 1591.020 1056.390 ;
        RECT 1768.020 1056.380 1771.020 1056.390 ;
        RECT 1948.020 1056.380 1951.020 1056.390 ;
        RECT 2128.020 1056.380 2131.020 1056.390 ;
        RECT 2308.020 1056.380 2311.020 1056.390 ;
        RECT 2488.020 1056.380 2491.020 1056.390 ;
        RECT 2668.020 1056.380 2671.020 1056.390 ;
        RECT 2848.020 1056.380 2851.020 1056.390 ;
        RECT 2959.500 1056.380 2962.500 1056.390 ;
        RECT -42.880 1053.380 2962.500 1056.380 ;
        RECT -42.880 1053.370 -39.880 1053.380 ;
        RECT 148.020 1053.370 151.020 1053.380 ;
        RECT 328.020 1053.370 331.020 1053.380 ;
        RECT 508.020 1053.370 511.020 1053.380 ;
        RECT 688.020 1053.370 691.020 1053.380 ;
        RECT 868.020 1053.370 871.020 1053.380 ;
        RECT 1048.020 1053.370 1051.020 1053.380 ;
        RECT 1228.020 1053.370 1231.020 1053.380 ;
        RECT 1408.020 1053.370 1411.020 1053.380 ;
        RECT 1588.020 1053.370 1591.020 1053.380 ;
        RECT 1768.020 1053.370 1771.020 1053.380 ;
        RECT 1948.020 1053.370 1951.020 1053.380 ;
        RECT 2128.020 1053.370 2131.020 1053.380 ;
        RECT 2308.020 1053.370 2311.020 1053.380 ;
        RECT 2488.020 1053.370 2491.020 1053.380 ;
        RECT 2668.020 1053.370 2671.020 1053.380 ;
        RECT 2848.020 1053.370 2851.020 1053.380 ;
        RECT 2959.500 1053.370 2962.500 1053.380 ;
        RECT -33.480 1038.380 -30.480 1038.390 ;
        RECT 130.020 1038.380 133.020 1038.390 ;
        RECT 310.020 1038.380 313.020 1038.390 ;
        RECT 490.020 1038.380 493.020 1038.390 ;
        RECT 670.020 1038.380 673.020 1038.390 ;
        RECT 850.020 1038.380 853.020 1038.390 ;
        RECT 1030.020 1038.380 1033.020 1038.390 ;
        RECT 1210.020 1038.380 1213.020 1038.390 ;
        RECT 1390.020 1038.380 1393.020 1038.390 ;
        RECT 1570.020 1038.380 1573.020 1038.390 ;
        RECT 1750.020 1038.380 1753.020 1038.390 ;
        RECT 1930.020 1038.380 1933.020 1038.390 ;
        RECT 2110.020 1038.380 2113.020 1038.390 ;
        RECT 2290.020 1038.380 2293.020 1038.390 ;
        RECT 2470.020 1038.380 2473.020 1038.390 ;
        RECT 2650.020 1038.380 2653.020 1038.390 ;
        RECT 2830.020 1038.380 2833.020 1038.390 ;
        RECT 2950.100 1038.380 2953.100 1038.390 ;
        RECT -33.480 1035.380 2953.100 1038.380 ;
        RECT -33.480 1035.370 -30.480 1035.380 ;
        RECT 130.020 1035.370 133.020 1035.380 ;
        RECT 310.020 1035.370 313.020 1035.380 ;
        RECT 490.020 1035.370 493.020 1035.380 ;
        RECT 670.020 1035.370 673.020 1035.380 ;
        RECT 850.020 1035.370 853.020 1035.380 ;
        RECT 1030.020 1035.370 1033.020 1035.380 ;
        RECT 1210.020 1035.370 1213.020 1035.380 ;
        RECT 1390.020 1035.370 1393.020 1035.380 ;
        RECT 1570.020 1035.370 1573.020 1035.380 ;
        RECT 1750.020 1035.370 1753.020 1035.380 ;
        RECT 1930.020 1035.370 1933.020 1035.380 ;
        RECT 2110.020 1035.370 2113.020 1035.380 ;
        RECT 2290.020 1035.370 2293.020 1035.380 ;
        RECT 2470.020 1035.370 2473.020 1035.380 ;
        RECT 2650.020 1035.370 2653.020 1035.380 ;
        RECT 2830.020 1035.370 2833.020 1035.380 ;
        RECT 2950.100 1035.370 2953.100 1035.380 ;
        RECT -24.080 1020.380 -21.080 1020.390 ;
        RECT 112.020 1020.380 115.020 1020.390 ;
        RECT 292.020 1020.380 295.020 1020.390 ;
        RECT 472.020 1020.380 475.020 1020.390 ;
        RECT 652.020 1020.380 655.020 1020.390 ;
        RECT 832.020 1020.380 835.020 1020.390 ;
        RECT 1012.020 1020.380 1015.020 1020.390 ;
        RECT 1192.020 1020.380 1195.020 1020.390 ;
        RECT 1372.020 1020.380 1375.020 1020.390 ;
        RECT 1552.020 1020.380 1555.020 1020.390 ;
        RECT 1732.020 1020.380 1735.020 1020.390 ;
        RECT 1912.020 1020.380 1915.020 1020.390 ;
        RECT 2092.020 1020.380 2095.020 1020.390 ;
        RECT 2272.020 1020.380 2275.020 1020.390 ;
        RECT 2452.020 1020.380 2455.020 1020.390 ;
        RECT 2632.020 1020.380 2635.020 1020.390 ;
        RECT 2812.020 1020.380 2815.020 1020.390 ;
        RECT 2940.700 1020.380 2943.700 1020.390 ;
        RECT -24.080 1017.380 2943.700 1020.380 ;
        RECT -24.080 1017.370 -21.080 1017.380 ;
        RECT 112.020 1017.370 115.020 1017.380 ;
        RECT 292.020 1017.370 295.020 1017.380 ;
        RECT 472.020 1017.370 475.020 1017.380 ;
        RECT 652.020 1017.370 655.020 1017.380 ;
        RECT 832.020 1017.370 835.020 1017.380 ;
        RECT 1012.020 1017.370 1015.020 1017.380 ;
        RECT 1192.020 1017.370 1195.020 1017.380 ;
        RECT 1372.020 1017.370 1375.020 1017.380 ;
        RECT 1552.020 1017.370 1555.020 1017.380 ;
        RECT 1732.020 1017.370 1735.020 1017.380 ;
        RECT 1912.020 1017.370 1915.020 1017.380 ;
        RECT 2092.020 1017.370 2095.020 1017.380 ;
        RECT 2272.020 1017.370 2275.020 1017.380 ;
        RECT 2452.020 1017.370 2455.020 1017.380 ;
        RECT 2632.020 1017.370 2635.020 1017.380 ;
        RECT 2812.020 1017.370 2815.020 1017.380 ;
        RECT 2940.700 1017.370 2943.700 1017.380 ;
        RECT -14.680 1002.380 -11.680 1002.390 ;
        RECT 94.020 1002.380 97.020 1002.390 ;
        RECT 274.020 1002.380 277.020 1002.390 ;
        RECT 454.020 1002.380 457.020 1002.390 ;
        RECT 634.020 1002.380 637.020 1002.390 ;
        RECT 814.020 1002.380 817.020 1002.390 ;
        RECT 994.020 1002.380 997.020 1002.390 ;
        RECT 1174.020 1002.380 1177.020 1002.390 ;
        RECT 1354.020 1002.380 1357.020 1002.390 ;
        RECT 1534.020 1002.380 1537.020 1002.390 ;
        RECT 1714.020 1002.380 1717.020 1002.390 ;
        RECT 1894.020 1002.380 1897.020 1002.390 ;
        RECT 2074.020 1002.380 2077.020 1002.390 ;
        RECT 2254.020 1002.380 2257.020 1002.390 ;
        RECT 2434.020 1002.380 2437.020 1002.390 ;
        RECT 2614.020 1002.380 2617.020 1002.390 ;
        RECT 2794.020 1002.380 2797.020 1002.390 ;
        RECT 2931.300 1002.380 2934.300 1002.390 ;
        RECT -14.680 999.380 2934.300 1002.380 ;
        RECT -14.680 999.370 -11.680 999.380 ;
        RECT 94.020 999.370 97.020 999.380 ;
        RECT 274.020 999.370 277.020 999.380 ;
        RECT 454.020 999.370 457.020 999.380 ;
        RECT 634.020 999.370 637.020 999.380 ;
        RECT 814.020 999.370 817.020 999.380 ;
        RECT 994.020 999.370 997.020 999.380 ;
        RECT 1174.020 999.370 1177.020 999.380 ;
        RECT 1354.020 999.370 1357.020 999.380 ;
        RECT 1534.020 999.370 1537.020 999.380 ;
        RECT 1714.020 999.370 1717.020 999.380 ;
        RECT 1894.020 999.370 1897.020 999.380 ;
        RECT 2074.020 999.370 2077.020 999.380 ;
        RECT 2254.020 999.370 2257.020 999.380 ;
        RECT 2434.020 999.370 2437.020 999.380 ;
        RECT 2614.020 999.370 2617.020 999.380 ;
        RECT 2794.020 999.370 2797.020 999.380 ;
        RECT 2931.300 999.370 2934.300 999.380 ;
        RECT -42.880 876.380 -39.880 876.390 ;
        RECT 148.020 876.380 151.020 876.390 ;
        RECT 328.020 876.380 331.020 876.390 ;
        RECT 508.020 876.380 511.020 876.390 ;
        RECT 688.020 876.380 691.020 876.390 ;
        RECT 868.020 876.380 871.020 876.390 ;
        RECT 1048.020 876.380 1051.020 876.390 ;
        RECT 1228.020 876.380 1231.020 876.390 ;
        RECT 1408.020 876.380 1411.020 876.390 ;
        RECT 1588.020 876.380 1591.020 876.390 ;
        RECT 1768.020 876.380 1771.020 876.390 ;
        RECT 1948.020 876.380 1951.020 876.390 ;
        RECT 2128.020 876.380 2131.020 876.390 ;
        RECT 2308.020 876.380 2311.020 876.390 ;
        RECT 2488.020 876.380 2491.020 876.390 ;
        RECT 2668.020 876.380 2671.020 876.390 ;
        RECT 2848.020 876.380 2851.020 876.390 ;
        RECT 2959.500 876.380 2962.500 876.390 ;
        RECT -42.880 873.380 2962.500 876.380 ;
        RECT -42.880 873.370 -39.880 873.380 ;
        RECT 148.020 873.370 151.020 873.380 ;
        RECT 328.020 873.370 331.020 873.380 ;
        RECT 508.020 873.370 511.020 873.380 ;
        RECT 688.020 873.370 691.020 873.380 ;
        RECT 868.020 873.370 871.020 873.380 ;
        RECT 1048.020 873.370 1051.020 873.380 ;
        RECT 1228.020 873.370 1231.020 873.380 ;
        RECT 1408.020 873.370 1411.020 873.380 ;
        RECT 1588.020 873.370 1591.020 873.380 ;
        RECT 1768.020 873.370 1771.020 873.380 ;
        RECT 1948.020 873.370 1951.020 873.380 ;
        RECT 2128.020 873.370 2131.020 873.380 ;
        RECT 2308.020 873.370 2311.020 873.380 ;
        RECT 2488.020 873.370 2491.020 873.380 ;
        RECT 2668.020 873.370 2671.020 873.380 ;
        RECT 2848.020 873.370 2851.020 873.380 ;
        RECT 2959.500 873.370 2962.500 873.380 ;
        RECT -33.480 858.380 -30.480 858.390 ;
        RECT 130.020 858.380 133.020 858.390 ;
        RECT 310.020 858.380 313.020 858.390 ;
        RECT 490.020 858.380 493.020 858.390 ;
        RECT 670.020 858.380 673.020 858.390 ;
        RECT 850.020 858.380 853.020 858.390 ;
        RECT 1030.020 858.380 1033.020 858.390 ;
        RECT 1210.020 858.380 1213.020 858.390 ;
        RECT 1390.020 858.380 1393.020 858.390 ;
        RECT 1570.020 858.380 1573.020 858.390 ;
        RECT 1750.020 858.380 1753.020 858.390 ;
        RECT 1930.020 858.380 1933.020 858.390 ;
        RECT 2110.020 858.380 2113.020 858.390 ;
        RECT 2290.020 858.380 2293.020 858.390 ;
        RECT 2470.020 858.380 2473.020 858.390 ;
        RECT 2650.020 858.380 2653.020 858.390 ;
        RECT 2830.020 858.380 2833.020 858.390 ;
        RECT 2950.100 858.380 2953.100 858.390 ;
        RECT -33.480 855.380 2953.100 858.380 ;
        RECT -33.480 855.370 -30.480 855.380 ;
        RECT 130.020 855.370 133.020 855.380 ;
        RECT 310.020 855.370 313.020 855.380 ;
        RECT 490.020 855.370 493.020 855.380 ;
        RECT 670.020 855.370 673.020 855.380 ;
        RECT 850.020 855.370 853.020 855.380 ;
        RECT 1030.020 855.370 1033.020 855.380 ;
        RECT 1210.020 855.370 1213.020 855.380 ;
        RECT 1390.020 855.370 1393.020 855.380 ;
        RECT 1570.020 855.370 1573.020 855.380 ;
        RECT 1750.020 855.370 1753.020 855.380 ;
        RECT 1930.020 855.370 1933.020 855.380 ;
        RECT 2110.020 855.370 2113.020 855.380 ;
        RECT 2290.020 855.370 2293.020 855.380 ;
        RECT 2470.020 855.370 2473.020 855.380 ;
        RECT 2650.020 855.370 2653.020 855.380 ;
        RECT 2830.020 855.370 2833.020 855.380 ;
        RECT 2950.100 855.370 2953.100 855.380 ;
        RECT -24.080 840.380 -21.080 840.390 ;
        RECT 112.020 840.380 115.020 840.390 ;
        RECT 292.020 840.380 295.020 840.390 ;
        RECT 472.020 840.380 475.020 840.390 ;
        RECT 652.020 840.380 655.020 840.390 ;
        RECT 832.020 840.380 835.020 840.390 ;
        RECT 1012.020 840.380 1015.020 840.390 ;
        RECT 1192.020 840.380 1195.020 840.390 ;
        RECT 1372.020 840.380 1375.020 840.390 ;
        RECT 1552.020 840.380 1555.020 840.390 ;
        RECT 1732.020 840.380 1735.020 840.390 ;
        RECT 1912.020 840.380 1915.020 840.390 ;
        RECT 2092.020 840.380 2095.020 840.390 ;
        RECT 2272.020 840.380 2275.020 840.390 ;
        RECT 2452.020 840.380 2455.020 840.390 ;
        RECT 2632.020 840.380 2635.020 840.390 ;
        RECT 2812.020 840.380 2815.020 840.390 ;
        RECT 2940.700 840.380 2943.700 840.390 ;
        RECT -24.080 837.380 2943.700 840.380 ;
        RECT -24.080 837.370 -21.080 837.380 ;
        RECT 112.020 837.370 115.020 837.380 ;
        RECT 292.020 837.370 295.020 837.380 ;
        RECT 472.020 837.370 475.020 837.380 ;
        RECT 652.020 837.370 655.020 837.380 ;
        RECT 832.020 837.370 835.020 837.380 ;
        RECT 1012.020 837.370 1015.020 837.380 ;
        RECT 1192.020 837.370 1195.020 837.380 ;
        RECT 1372.020 837.370 1375.020 837.380 ;
        RECT 1552.020 837.370 1555.020 837.380 ;
        RECT 1732.020 837.370 1735.020 837.380 ;
        RECT 1912.020 837.370 1915.020 837.380 ;
        RECT 2092.020 837.370 2095.020 837.380 ;
        RECT 2272.020 837.370 2275.020 837.380 ;
        RECT 2452.020 837.370 2455.020 837.380 ;
        RECT 2632.020 837.370 2635.020 837.380 ;
        RECT 2812.020 837.370 2815.020 837.380 ;
        RECT 2940.700 837.370 2943.700 837.380 ;
        RECT -14.680 822.380 -11.680 822.390 ;
        RECT 94.020 822.380 97.020 822.390 ;
        RECT 274.020 822.380 277.020 822.390 ;
        RECT 454.020 822.380 457.020 822.390 ;
        RECT 634.020 822.380 637.020 822.390 ;
        RECT 814.020 822.380 817.020 822.390 ;
        RECT 994.020 822.380 997.020 822.390 ;
        RECT 1174.020 822.380 1177.020 822.390 ;
        RECT 1354.020 822.380 1357.020 822.390 ;
        RECT 1534.020 822.380 1537.020 822.390 ;
        RECT 1714.020 822.380 1717.020 822.390 ;
        RECT 1894.020 822.380 1897.020 822.390 ;
        RECT 2074.020 822.380 2077.020 822.390 ;
        RECT 2254.020 822.380 2257.020 822.390 ;
        RECT 2434.020 822.380 2437.020 822.390 ;
        RECT 2614.020 822.380 2617.020 822.390 ;
        RECT 2794.020 822.380 2797.020 822.390 ;
        RECT 2931.300 822.380 2934.300 822.390 ;
        RECT -14.680 819.380 2934.300 822.380 ;
        RECT -14.680 819.370 -11.680 819.380 ;
        RECT 94.020 819.370 97.020 819.380 ;
        RECT 274.020 819.370 277.020 819.380 ;
        RECT 454.020 819.370 457.020 819.380 ;
        RECT 634.020 819.370 637.020 819.380 ;
        RECT 814.020 819.370 817.020 819.380 ;
        RECT 994.020 819.370 997.020 819.380 ;
        RECT 1174.020 819.370 1177.020 819.380 ;
        RECT 1354.020 819.370 1357.020 819.380 ;
        RECT 1534.020 819.370 1537.020 819.380 ;
        RECT 1714.020 819.370 1717.020 819.380 ;
        RECT 1894.020 819.370 1897.020 819.380 ;
        RECT 2074.020 819.370 2077.020 819.380 ;
        RECT 2254.020 819.370 2257.020 819.380 ;
        RECT 2434.020 819.370 2437.020 819.380 ;
        RECT 2614.020 819.370 2617.020 819.380 ;
        RECT 2794.020 819.370 2797.020 819.380 ;
        RECT 2931.300 819.370 2934.300 819.380 ;
        RECT -42.880 696.380 -39.880 696.390 ;
        RECT 148.020 696.380 151.020 696.390 ;
        RECT 328.020 696.380 331.020 696.390 ;
        RECT 508.020 696.380 511.020 696.390 ;
        RECT 688.020 696.380 691.020 696.390 ;
        RECT 868.020 696.380 871.020 696.390 ;
        RECT 1048.020 696.380 1051.020 696.390 ;
        RECT 1228.020 696.380 1231.020 696.390 ;
        RECT 1408.020 696.380 1411.020 696.390 ;
        RECT 1588.020 696.380 1591.020 696.390 ;
        RECT 1768.020 696.380 1771.020 696.390 ;
        RECT 1948.020 696.380 1951.020 696.390 ;
        RECT 2128.020 696.380 2131.020 696.390 ;
        RECT 2308.020 696.380 2311.020 696.390 ;
        RECT 2488.020 696.380 2491.020 696.390 ;
        RECT 2668.020 696.380 2671.020 696.390 ;
        RECT 2848.020 696.380 2851.020 696.390 ;
        RECT 2959.500 696.380 2962.500 696.390 ;
        RECT -42.880 693.380 2962.500 696.380 ;
        RECT -42.880 693.370 -39.880 693.380 ;
        RECT 148.020 693.370 151.020 693.380 ;
        RECT 328.020 693.370 331.020 693.380 ;
        RECT 508.020 693.370 511.020 693.380 ;
        RECT 688.020 693.370 691.020 693.380 ;
        RECT 868.020 693.370 871.020 693.380 ;
        RECT 1048.020 693.370 1051.020 693.380 ;
        RECT 1228.020 693.370 1231.020 693.380 ;
        RECT 1408.020 693.370 1411.020 693.380 ;
        RECT 1588.020 693.370 1591.020 693.380 ;
        RECT 1768.020 693.370 1771.020 693.380 ;
        RECT 1948.020 693.370 1951.020 693.380 ;
        RECT 2128.020 693.370 2131.020 693.380 ;
        RECT 2308.020 693.370 2311.020 693.380 ;
        RECT 2488.020 693.370 2491.020 693.380 ;
        RECT 2668.020 693.370 2671.020 693.380 ;
        RECT 2848.020 693.370 2851.020 693.380 ;
        RECT 2959.500 693.370 2962.500 693.380 ;
        RECT -33.480 678.380 -30.480 678.390 ;
        RECT 130.020 678.380 133.020 678.390 ;
        RECT 310.020 678.380 313.020 678.390 ;
        RECT 490.020 678.380 493.020 678.390 ;
        RECT 670.020 678.380 673.020 678.390 ;
        RECT 850.020 678.380 853.020 678.390 ;
        RECT 1030.020 678.380 1033.020 678.390 ;
        RECT 1210.020 678.380 1213.020 678.390 ;
        RECT 1390.020 678.380 1393.020 678.390 ;
        RECT 1570.020 678.380 1573.020 678.390 ;
        RECT 1750.020 678.380 1753.020 678.390 ;
        RECT 1930.020 678.380 1933.020 678.390 ;
        RECT 2110.020 678.380 2113.020 678.390 ;
        RECT 2290.020 678.380 2293.020 678.390 ;
        RECT 2470.020 678.380 2473.020 678.390 ;
        RECT 2650.020 678.380 2653.020 678.390 ;
        RECT 2830.020 678.380 2833.020 678.390 ;
        RECT 2950.100 678.380 2953.100 678.390 ;
        RECT -33.480 675.380 2953.100 678.380 ;
        RECT -33.480 675.370 -30.480 675.380 ;
        RECT 130.020 675.370 133.020 675.380 ;
        RECT 310.020 675.370 313.020 675.380 ;
        RECT 490.020 675.370 493.020 675.380 ;
        RECT 670.020 675.370 673.020 675.380 ;
        RECT 850.020 675.370 853.020 675.380 ;
        RECT 1030.020 675.370 1033.020 675.380 ;
        RECT 1210.020 675.370 1213.020 675.380 ;
        RECT 1390.020 675.370 1393.020 675.380 ;
        RECT 1570.020 675.370 1573.020 675.380 ;
        RECT 1750.020 675.370 1753.020 675.380 ;
        RECT 1930.020 675.370 1933.020 675.380 ;
        RECT 2110.020 675.370 2113.020 675.380 ;
        RECT 2290.020 675.370 2293.020 675.380 ;
        RECT 2470.020 675.370 2473.020 675.380 ;
        RECT 2650.020 675.370 2653.020 675.380 ;
        RECT 2830.020 675.370 2833.020 675.380 ;
        RECT 2950.100 675.370 2953.100 675.380 ;
        RECT -24.080 660.380 -21.080 660.390 ;
        RECT 112.020 660.380 115.020 660.390 ;
        RECT 292.020 660.380 295.020 660.390 ;
        RECT 472.020 660.380 475.020 660.390 ;
        RECT 652.020 660.380 655.020 660.390 ;
        RECT 832.020 660.380 835.020 660.390 ;
        RECT 1012.020 660.380 1015.020 660.390 ;
        RECT 1192.020 660.380 1195.020 660.390 ;
        RECT 1372.020 660.380 1375.020 660.390 ;
        RECT 1552.020 660.380 1555.020 660.390 ;
        RECT 1732.020 660.380 1735.020 660.390 ;
        RECT 1912.020 660.380 1915.020 660.390 ;
        RECT 2092.020 660.380 2095.020 660.390 ;
        RECT 2272.020 660.380 2275.020 660.390 ;
        RECT 2452.020 660.380 2455.020 660.390 ;
        RECT 2632.020 660.380 2635.020 660.390 ;
        RECT 2812.020 660.380 2815.020 660.390 ;
        RECT 2940.700 660.380 2943.700 660.390 ;
        RECT -24.080 657.380 2943.700 660.380 ;
        RECT -24.080 657.370 -21.080 657.380 ;
        RECT 112.020 657.370 115.020 657.380 ;
        RECT 292.020 657.370 295.020 657.380 ;
        RECT 472.020 657.370 475.020 657.380 ;
        RECT 652.020 657.370 655.020 657.380 ;
        RECT 832.020 657.370 835.020 657.380 ;
        RECT 1012.020 657.370 1015.020 657.380 ;
        RECT 1192.020 657.370 1195.020 657.380 ;
        RECT 1372.020 657.370 1375.020 657.380 ;
        RECT 1552.020 657.370 1555.020 657.380 ;
        RECT 1732.020 657.370 1735.020 657.380 ;
        RECT 1912.020 657.370 1915.020 657.380 ;
        RECT 2092.020 657.370 2095.020 657.380 ;
        RECT 2272.020 657.370 2275.020 657.380 ;
        RECT 2452.020 657.370 2455.020 657.380 ;
        RECT 2632.020 657.370 2635.020 657.380 ;
        RECT 2812.020 657.370 2815.020 657.380 ;
        RECT 2940.700 657.370 2943.700 657.380 ;
        RECT -14.680 642.380 -11.680 642.390 ;
        RECT 94.020 642.380 97.020 642.390 ;
        RECT 274.020 642.380 277.020 642.390 ;
        RECT 454.020 642.380 457.020 642.390 ;
        RECT 634.020 642.380 637.020 642.390 ;
        RECT 814.020 642.380 817.020 642.390 ;
        RECT 994.020 642.380 997.020 642.390 ;
        RECT 1174.020 642.380 1177.020 642.390 ;
        RECT 1354.020 642.380 1357.020 642.390 ;
        RECT 1534.020 642.380 1537.020 642.390 ;
        RECT 1714.020 642.380 1717.020 642.390 ;
        RECT 1894.020 642.380 1897.020 642.390 ;
        RECT 2074.020 642.380 2077.020 642.390 ;
        RECT 2254.020 642.380 2257.020 642.390 ;
        RECT 2434.020 642.380 2437.020 642.390 ;
        RECT 2614.020 642.380 2617.020 642.390 ;
        RECT 2794.020 642.380 2797.020 642.390 ;
        RECT 2931.300 642.380 2934.300 642.390 ;
        RECT -14.680 639.380 2934.300 642.380 ;
        RECT -14.680 639.370 -11.680 639.380 ;
        RECT 94.020 639.370 97.020 639.380 ;
        RECT 274.020 639.370 277.020 639.380 ;
        RECT 454.020 639.370 457.020 639.380 ;
        RECT 634.020 639.370 637.020 639.380 ;
        RECT 814.020 639.370 817.020 639.380 ;
        RECT 994.020 639.370 997.020 639.380 ;
        RECT 1174.020 639.370 1177.020 639.380 ;
        RECT 1354.020 639.370 1357.020 639.380 ;
        RECT 1534.020 639.370 1537.020 639.380 ;
        RECT 1714.020 639.370 1717.020 639.380 ;
        RECT 1894.020 639.370 1897.020 639.380 ;
        RECT 2074.020 639.370 2077.020 639.380 ;
        RECT 2254.020 639.370 2257.020 639.380 ;
        RECT 2434.020 639.370 2437.020 639.380 ;
        RECT 2614.020 639.370 2617.020 639.380 ;
        RECT 2794.020 639.370 2797.020 639.380 ;
        RECT 2931.300 639.370 2934.300 639.380 ;
        RECT -42.880 516.380 -39.880 516.390 ;
        RECT 148.020 516.380 151.020 516.390 ;
        RECT 328.020 516.380 331.020 516.390 ;
        RECT 508.020 516.380 511.020 516.390 ;
        RECT 688.020 516.380 691.020 516.390 ;
        RECT 868.020 516.380 871.020 516.390 ;
        RECT 1048.020 516.380 1051.020 516.390 ;
        RECT 1228.020 516.380 1231.020 516.390 ;
        RECT 1408.020 516.380 1411.020 516.390 ;
        RECT 1588.020 516.380 1591.020 516.390 ;
        RECT 1768.020 516.380 1771.020 516.390 ;
        RECT 1948.020 516.380 1951.020 516.390 ;
        RECT 2128.020 516.380 2131.020 516.390 ;
        RECT 2308.020 516.380 2311.020 516.390 ;
        RECT 2488.020 516.380 2491.020 516.390 ;
        RECT 2668.020 516.380 2671.020 516.390 ;
        RECT 2848.020 516.380 2851.020 516.390 ;
        RECT 2959.500 516.380 2962.500 516.390 ;
        RECT -42.880 513.380 2962.500 516.380 ;
        RECT -42.880 513.370 -39.880 513.380 ;
        RECT 148.020 513.370 151.020 513.380 ;
        RECT 328.020 513.370 331.020 513.380 ;
        RECT 508.020 513.370 511.020 513.380 ;
        RECT 688.020 513.370 691.020 513.380 ;
        RECT 868.020 513.370 871.020 513.380 ;
        RECT 1048.020 513.370 1051.020 513.380 ;
        RECT 1228.020 513.370 1231.020 513.380 ;
        RECT 1408.020 513.370 1411.020 513.380 ;
        RECT 1588.020 513.370 1591.020 513.380 ;
        RECT 1768.020 513.370 1771.020 513.380 ;
        RECT 1948.020 513.370 1951.020 513.380 ;
        RECT 2128.020 513.370 2131.020 513.380 ;
        RECT 2308.020 513.370 2311.020 513.380 ;
        RECT 2488.020 513.370 2491.020 513.380 ;
        RECT 2668.020 513.370 2671.020 513.380 ;
        RECT 2848.020 513.370 2851.020 513.380 ;
        RECT 2959.500 513.370 2962.500 513.380 ;
        RECT -33.480 498.380 -30.480 498.390 ;
        RECT 130.020 498.380 133.020 498.390 ;
        RECT 310.020 498.380 313.020 498.390 ;
        RECT 490.020 498.380 493.020 498.390 ;
        RECT 670.020 498.380 673.020 498.390 ;
        RECT 850.020 498.380 853.020 498.390 ;
        RECT 1030.020 498.380 1033.020 498.390 ;
        RECT 1210.020 498.380 1213.020 498.390 ;
        RECT 1390.020 498.380 1393.020 498.390 ;
        RECT 1570.020 498.380 1573.020 498.390 ;
        RECT 1750.020 498.380 1753.020 498.390 ;
        RECT 1930.020 498.380 1933.020 498.390 ;
        RECT 2110.020 498.380 2113.020 498.390 ;
        RECT 2290.020 498.380 2293.020 498.390 ;
        RECT 2470.020 498.380 2473.020 498.390 ;
        RECT 2650.020 498.380 2653.020 498.390 ;
        RECT 2830.020 498.380 2833.020 498.390 ;
        RECT 2950.100 498.380 2953.100 498.390 ;
        RECT -33.480 495.380 2953.100 498.380 ;
        RECT -33.480 495.370 -30.480 495.380 ;
        RECT 130.020 495.370 133.020 495.380 ;
        RECT 310.020 495.370 313.020 495.380 ;
        RECT 490.020 495.370 493.020 495.380 ;
        RECT 670.020 495.370 673.020 495.380 ;
        RECT 850.020 495.370 853.020 495.380 ;
        RECT 1030.020 495.370 1033.020 495.380 ;
        RECT 1210.020 495.370 1213.020 495.380 ;
        RECT 1390.020 495.370 1393.020 495.380 ;
        RECT 1570.020 495.370 1573.020 495.380 ;
        RECT 1750.020 495.370 1753.020 495.380 ;
        RECT 1930.020 495.370 1933.020 495.380 ;
        RECT 2110.020 495.370 2113.020 495.380 ;
        RECT 2290.020 495.370 2293.020 495.380 ;
        RECT 2470.020 495.370 2473.020 495.380 ;
        RECT 2650.020 495.370 2653.020 495.380 ;
        RECT 2830.020 495.370 2833.020 495.380 ;
        RECT 2950.100 495.370 2953.100 495.380 ;
        RECT -24.080 480.380 -21.080 480.390 ;
        RECT 112.020 480.380 115.020 480.390 ;
        RECT 292.020 480.380 295.020 480.390 ;
        RECT 472.020 480.380 475.020 480.390 ;
        RECT 652.020 480.380 655.020 480.390 ;
        RECT 832.020 480.380 835.020 480.390 ;
        RECT 1012.020 480.380 1015.020 480.390 ;
        RECT 1192.020 480.380 1195.020 480.390 ;
        RECT 1372.020 480.380 1375.020 480.390 ;
        RECT 1552.020 480.380 1555.020 480.390 ;
        RECT 1732.020 480.380 1735.020 480.390 ;
        RECT 1912.020 480.380 1915.020 480.390 ;
        RECT 2092.020 480.380 2095.020 480.390 ;
        RECT 2272.020 480.380 2275.020 480.390 ;
        RECT 2452.020 480.380 2455.020 480.390 ;
        RECT 2632.020 480.380 2635.020 480.390 ;
        RECT 2812.020 480.380 2815.020 480.390 ;
        RECT 2940.700 480.380 2943.700 480.390 ;
        RECT -24.080 477.380 2943.700 480.380 ;
        RECT -24.080 477.370 -21.080 477.380 ;
        RECT 112.020 477.370 115.020 477.380 ;
        RECT 292.020 477.370 295.020 477.380 ;
        RECT 472.020 477.370 475.020 477.380 ;
        RECT 652.020 477.370 655.020 477.380 ;
        RECT 832.020 477.370 835.020 477.380 ;
        RECT 1012.020 477.370 1015.020 477.380 ;
        RECT 1192.020 477.370 1195.020 477.380 ;
        RECT 1372.020 477.370 1375.020 477.380 ;
        RECT 1552.020 477.370 1555.020 477.380 ;
        RECT 1732.020 477.370 1735.020 477.380 ;
        RECT 1912.020 477.370 1915.020 477.380 ;
        RECT 2092.020 477.370 2095.020 477.380 ;
        RECT 2272.020 477.370 2275.020 477.380 ;
        RECT 2452.020 477.370 2455.020 477.380 ;
        RECT 2632.020 477.370 2635.020 477.380 ;
        RECT 2812.020 477.370 2815.020 477.380 ;
        RECT 2940.700 477.370 2943.700 477.380 ;
        RECT -14.680 462.380 -11.680 462.390 ;
        RECT 94.020 462.380 97.020 462.390 ;
        RECT 274.020 462.380 277.020 462.390 ;
        RECT 454.020 462.380 457.020 462.390 ;
        RECT 634.020 462.380 637.020 462.390 ;
        RECT 814.020 462.380 817.020 462.390 ;
        RECT 994.020 462.380 997.020 462.390 ;
        RECT 1174.020 462.380 1177.020 462.390 ;
        RECT 1354.020 462.380 1357.020 462.390 ;
        RECT 1534.020 462.380 1537.020 462.390 ;
        RECT 1714.020 462.380 1717.020 462.390 ;
        RECT 1894.020 462.380 1897.020 462.390 ;
        RECT 2074.020 462.380 2077.020 462.390 ;
        RECT 2254.020 462.380 2257.020 462.390 ;
        RECT 2434.020 462.380 2437.020 462.390 ;
        RECT 2614.020 462.380 2617.020 462.390 ;
        RECT 2794.020 462.380 2797.020 462.390 ;
        RECT 2931.300 462.380 2934.300 462.390 ;
        RECT -14.680 459.380 2934.300 462.380 ;
        RECT -14.680 459.370 -11.680 459.380 ;
        RECT 94.020 459.370 97.020 459.380 ;
        RECT 274.020 459.370 277.020 459.380 ;
        RECT 454.020 459.370 457.020 459.380 ;
        RECT 634.020 459.370 637.020 459.380 ;
        RECT 814.020 459.370 817.020 459.380 ;
        RECT 994.020 459.370 997.020 459.380 ;
        RECT 1174.020 459.370 1177.020 459.380 ;
        RECT 1354.020 459.370 1357.020 459.380 ;
        RECT 1534.020 459.370 1537.020 459.380 ;
        RECT 1714.020 459.370 1717.020 459.380 ;
        RECT 1894.020 459.370 1897.020 459.380 ;
        RECT 2074.020 459.370 2077.020 459.380 ;
        RECT 2254.020 459.370 2257.020 459.380 ;
        RECT 2434.020 459.370 2437.020 459.380 ;
        RECT 2614.020 459.370 2617.020 459.380 ;
        RECT 2794.020 459.370 2797.020 459.380 ;
        RECT 2931.300 459.370 2934.300 459.380 ;
        RECT -42.880 336.380 -39.880 336.390 ;
        RECT 148.020 336.380 151.020 336.390 ;
        RECT 328.020 336.380 331.020 336.390 ;
        RECT 508.020 336.380 511.020 336.390 ;
        RECT 688.020 336.380 691.020 336.390 ;
        RECT 868.020 336.380 871.020 336.390 ;
        RECT 1048.020 336.380 1051.020 336.390 ;
        RECT 1228.020 336.380 1231.020 336.390 ;
        RECT 1408.020 336.380 1411.020 336.390 ;
        RECT 1588.020 336.380 1591.020 336.390 ;
        RECT 1768.020 336.380 1771.020 336.390 ;
        RECT 1948.020 336.380 1951.020 336.390 ;
        RECT 2128.020 336.380 2131.020 336.390 ;
        RECT 2308.020 336.380 2311.020 336.390 ;
        RECT 2488.020 336.380 2491.020 336.390 ;
        RECT 2668.020 336.380 2671.020 336.390 ;
        RECT 2848.020 336.380 2851.020 336.390 ;
        RECT 2959.500 336.380 2962.500 336.390 ;
        RECT -42.880 333.380 2962.500 336.380 ;
        RECT -42.880 333.370 -39.880 333.380 ;
        RECT 148.020 333.370 151.020 333.380 ;
        RECT 328.020 333.370 331.020 333.380 ;
        RECT 508.020 333.370 511.020 333.380 ;
        RECT 688.020 333.370 691.020 333.380 ;
        RECT 868.020 333.370 871.020 333.380 ;
        RECT 1048.020 333.370 1051.020 333.380 ;
        RECT 1228.020 333.370 1231.020 333.380 ;
        RECT 1408.020 333.370 1411.020 333.380 ;
        RECT 1588.020 333.370 1591.020 333.380 ;
        RECT 1768.020 333.370 1771.020 333.380 ;
        RECT 1948.020 333.370 1951.020 333.380 ;
        RECT 2128.020 333.370 2131.020 333.380 ;
        RECT 2308.020 333.370 2311.020 333.380 ;
        RECT 2488.020 333.370 2491.020 333.380 ;
        RECT 2668.020 333.370 2671.020 333.380 ;
        RECT 2848.020 333.370 2851.020 333.380 ;
        RECT 2959.500 333.370 2962.500 333.380 ;
        RECT -33.480 318.380 -30.480 318.390 ;
        RECT 130.020 318.380 133.020 318.390 ;
        RECT 310.020 318.380 313.020 318.390 ;
        RECT 490.020 318.380 493.020 318.390 ;
        RECT 670.020 318.380 673.020 318.390 ;
        RECT 850.020 318.380 853.020 318.390 ;
        RECT 1030.020 318.380 1033.020 318.390 ;
        RECT 1210.020 318.380 1213.020 318.390 ;
        RECT 1390.020 318.380 1393.020 318.390 ;
        RECT 1570.020 318.380 1573.020 318.390 ;
        RECT 1750.020 318.380 1753.020 318.390 ;
        RECT 1930.020 318.380 1933.020 318.390 ;
        RECT 2110.020 318.380 2113.020 318.390 ;
        RECT 2290.020 318.380 2293.020 318.390 ;
        RECT 2470.020 318.380 2473.020 318.390 ;
        RECT 2650.020 318.380 2653.020 318.390 ;
        RECT 2830.020 318.380 2833.020 318.390 ;
        RECT 2950.100 318.380 2953.100 318.390 ;
        RECT -33.480 315.380 2953.100 318.380 ;
        RECT -33.480 315.370 -30.480 315.380 ;
        RECT 130.020 315.370 133.020 315.380 ;
        RECT 310.020 315.370 313.020 315.380 ;
        RECT 490.020 315.370 493.020 315.380 ;
        RECT 670.020 315.370 673.020 315.380 ;
        RECT 850.020 315.370 853.020 315.380 ;
        RECT 1030.020 315.370 1033.020 315.380 ;
        RECT 1210.020 315.370 1213.020 315.380 ;
        RECT 1390.020 315.370 1393.020 315.380 ;
        RECT 1570.020 315.370 1573.020 315.380 ;
        RECT 1750.020 315.370 1753.020 315.380 ;
        RECT 1930.020 315.370 1933.020 315.380 ;
        RECT 2110.020 315.370 2113.020 315.380 ;
        RECT 2290.020 315.370 2293.020 315.380 ;
        RECT 2470.020 315.370 2473.020 315.380 ;
        RECT 2650.020 315.370 2653.020 315.380 ;
        RECT 2830.020 315.370 2833.020 315.380 ;
        RECT 2950.100 315.370 2953.100 315.380 ;
        RECT -24.080 300.380 -21.080 300.390 ;
        RECT 112.020 300.380 115.020 300.390 ;
        RECT 292.020 300.380 295.020 300.390 ;
        RECT 472.020 300.380 475.020 300.390 ;
        RECT 652.020 300.380 655.020 300.390 ;
        RECT 832.020 300.380 835.020 300.390 ;
        RECT 1012.020 300.380 1015.020 300.390 ;
        RECT 1192.020 300.380 1195.020 300.390 ;
        RECT 1372.020 300.380 1375.020 300.390 ;
        RECT 1552.020 300.380 1555.020 300.390 ;
        RECT 1732.020 300.380 1735.020 300.390 ;
        RECT 1912.020 300.380 1915.020 300.390 ;
        RECT 2092.020 300.380 2095.020 300.390 ;
        RECT 2272.020 300.380 2275.020 300.390 ;
        RECT 2452.020 300.380 2455.020 300.390 ;
        RECT 2632.020 300.380 2635.020 300.390 ;
        RECT 2812.020 300.380 2815.020 300.390 ;
        RECT 2940.700 300.380 2943.700 300.390 ;
        RECT -24.080 297.380 2943.700 300.380 ;
        RECT -24.080 297.370 -21.080 297.380 ;
        RECT 112.020 297.370 115.020 297.380 ;
        RECT 292.020 297.370 295.020 297.380 ;
        RECT 472.020 297.370 475.020 297.380 ;
        RECT 652.020 297.370 655.020 297.380 ;
        RECT 832.020 297.370 835.020 297.380 ;
        RECT 1012.020 297.370 1015.020 297.380 ;
        RECT 1192.020 297.370 1195.020 297.380 ;
        RECT 1372.020 297.370 1375.020 297.380 ;
        RECT 1552.020 297.370 1555.020 297.380 ;
        RECT 1732.020 297.370 1735.020 297.380 ;
        RECT 1912.020 297.370 1915.020 297.380 ;
        RECT 2092.020 297.370 2095.020 297.380 ;
        RECT 2272.020 297.370 2275.020 297.380 ;
        RECT 2452.020 297.370 2455.020 297.380 ;
        RECT 2632.020 297.370 2635.020 297.380 ;
        RECT 2812.020 297.370 2815.020 297.380 ;
        RECT 2940.700 297.370 2943.700 297.380 ;
        RECT -14.680 282.380 -11.680 282.390 ;
        RECT 94.020 282.380 97.020 282.390 ;
        RECT 274.020 282.380 277.020 282.390 ;
        RECT 454.020 282.380 457.020 282.390 ;
        RECT 634.020 282.380 637.020 282.390 ;
        RECT 814.020 282.380 817.020 282.390 ;
        RECT 994.020 282.380 997.020 282.390 ;
        RECT 1174.020 282.380 1177.020 282.390 ;
        RECT 1354.020 282.380 1357.020 282.390 ;
        RECT 1534.020 282.380 1537.020 282.390 ;
        RECT 1714.020 282.380 1717.020 282.390 ;
        RECT 1894.020 282.380 1897.020 282.390 ;
        RECT 2074.020 282.380 2077.020 282.390 ;
        RECT 2254.020 282.380 2257.020 282.390 ;
        RECT 2434.020 282.380 2437.020 282.390 ;
        RECT 2614.020 282.380 2617.020 282.390 ;
        RECT 2794.020 282.380 2797.020 282.390 ;
        RECT 2931.300 282.380 2934.300 282.390 ;
        RECT -14.680 279.380 2934.300 282.380 ;
        RECT -14.680 279.370 -11.680 279.380 ;
        RECT 94.020 279.370 97.020 279.380 ;
        RECT 274.020 279.370 277.020 279.380 ;
        RECT 454.020 279.370 457.020 279.380 ;
        RECT 634.020 279.370 637.020 279.380 ;
        RECT 814.020 279.370 817.020 279.380 ;
        RECT 994.020 279.370 997.020 279.380 ;
        RECT 1174.020 279.370 1177.020 279.380 ;
        RECT 1354.020 279.370 1357.020 279.380 ;
        RECT 1534.020 279.370 1537.020 279.380 ;
        RECT 1714.020 279.370 1717.020 279.380 ;
        RECT 1894.020 279.370 1897.020 279.380 ;
        RECT 2074.020 279.370 2077.020 279.380 ;
        RECT 2254.020 279.370 2257.020 279.380 ;
        RECT 2434.020 279.370 2437.020 279.380 ;
        RECT 2614.020 279.370 2617.020 279.380 ;
        RECT 2794.020 279.370 2797.020 279.380 ;
        RECT 2931.300 279.370 2934.300 279.380 ;
        RECT -42.880 156.380 -39.880 156.390 ;
        RECT 148.020 156.380 151.020 156.390 ;
        RECT 328.020 156.380 331.020 156.390 ;
        RECT 508.020 156.380 511.020 156.390 ;
        RECT 688.020 156.380 691.020 156.390 ;
        RECT 868.020 156.380 871.020 156.390 ;
        RECT 1048.020 156.380 1051.020 156.390 ;
        RECT 1228.020 156.380 1231.020 156.390 ;
        RECT 1408.020 156.380 1411.020 156.390 ;
        RECT 1588.020 156.380 1591.020 156.390 ;
        RECT 1768.020 156.380 1771.020 156.390 ;
        RECT 1948.020 156.380 1951.020 156.390 ;
        RECT 2128.020 156.380 2131.020 156.390 ;
        RECT 2308.020 156.380 2311.020 156.390 ;
        RECT 2488.020 156.380 2491.020 156.390 ;
        RECT 2668.020 156.380 2671.020 156.390 ;
        RECT 2848.020 156.380 2851.020 156.390 ;
        RECT 2959.500 156.380 2962.500 156.390 ;
        RECT -42.880 153.380 2962.500 156.380 ;
        RECT -42.880 153.370 -39.880 153.380 ;
        RECT 148.020 153.370 151.020 153.380 ;
        RECT 328.020 153.370 331.020 153.380 ;
        RECT 508.020 153.370 511.020 153.380 ;
        RECT 688.020 153.370 691.020 153.380 ;
        RECT 868.020 153.370 871.020 153.380 ;
        RECT 1048.020 153.370 1051.020 153.380 ;
        RECT 1228.020 153.370 1231.020 153.380 ;
        RECT 1408.020 153.370 1411.020 153.380 ;
        RECT 1588.020 153.370 1591.020 153.380 ;
        RECT 1768.020 153.370 1771.020 153.380 ;
        RECT 1948.020 153.370 1951.020 153.380 ;
        RECT 2128.020 153.370 2131.020 153.380 ;
        RECT 2308.020 153.370 2311.020 153.380 ;
        RECT 2488.020 153.370 2491.020 153.380 ;
        RECT 2668.020 153.370 2671.020 153.380 ;
        RECT 2848.020 153.370 2851.020 153.380 ;
        RECT 2959.500 153.370 2962.500 153.380 ;
        RECT -33.480 138.380 -30.480 138.390 ;
        RECT 130.020 138.380 133.020 138.390 ;
        RECT 310.020 138.380 313.020 138.390 ;
        RECT 490.020 138.380 493.020 138.390 ;
        RECT 670.020 138.380 673.020 138.390 ;
        RECT 850.020 138.380 853.020 138.390 ;
        RECT 1030.020 138.380 1033.020 138.390 ;
        RECT 1210.020 138.380 1213.020 138.390 ;
        RECT 1390.020 138.380 1393.020 138.390 ;
        RECT 1570.020 138.380 1573.020 138.390 ;
        RECT 1750.020 138.380 1753.020 138.390 ;
        RECT 1930.020 138.380 1933.020 138.390 ;
        RECT 2110.020 138.380 2113.020 138.390 ;
        RECT 2290.020 138.380 2293.020 138.390 ;
        RECT 2470.020 138.380 2473.020 138.390 ;
        RECT 2650.020 138.380 2653.020 138.390 ;
        RECT 2830.020 138.380 2833.020 138.390 ;
        RECT 2950.100 138.380 2953.100 138.390 ;
        RECT -33.480 135.380 2953.100 138.380 ;
        RECT -33.480 135.370 -30.480 135.380 ;
        RECT 130.020 135.370 133.020 135.380 ;
        RECT 310.020 135.370 313.020 135.380 ;
        RECT 490.020 135.370 493.020 135.380 ;
        RECT 670.020 135.370 673.020 135.380 ;
        RECT 850.020 135.370 853.020 135.380 ;
        RECT 1030.020 135.370 1033.020 135.380 ;
        RECT 1210.020 135.370 1213.020 135.380 ;
        RECT 1390.020 135.370 1393.020 135.380 ;
        RECT 1570.020 135.370 1573.020 135.380 ;
        RECT 1750.020 135.370 1753.020 135.380 ;
        RECT 1930.020 135.370 1933.020 135.380 ;
        RECT 2110.020 135.370 2113.020 135.380 ;
        RECT 2290.020 135.370 2293.020 135.380 ;
        RECT 2470.020 135.370 2473.020 135.380 ;
        RECT 2650.020 135.370 2653.020 135.380 ;
        RECT 2830.020 135.370 2833.020 135.380 ;
        RECT 2950.100 135.370 2953.100 135.380 ;
        RECT -24.080 120.380 -21.080 120.390 ;
        RECT 112.020 120.380 115.020 120.390 ;
        RECT 292.020 120.380 295.020 120.390 ;
        RECT 472.020 120.380 475.020 120.390 ;
        RECT 652.020 120.380 655.020 120.390 ;
        RECT 832.020 120.380 835.020 120.390 ;
        RECT 1012.020 120.380 1015.020 120.390 ;
        RECT 1192.020 120.380 1195.020 120.390 ;
        RECT 1372.020 120.380 1375.020 120.390 ;
        RECT 1552.020 120.380 1555.020 120.390 ;
        RECT 1732.020 120.380 1735.020 120.390 ;
        RECT 1912.020 120.380 1915.020 120.390 ;
        RECT 2092.020 120.380 2095.020 120.390 ;
        RECT 2272.020 120.380 2275.020 120.390 ;
        RECT 2452.020 120.380 2455.020 120.390 ;
        RECT 2632.020 120.380 2635.020 120.390 ;
        RECT 2812.020 120.380 2815.020 120.390 ;
        RECT 2940.700 120.380 2943.700 120.390 ;
        RECT -24.080 117.380 2943.700 120.380 ;
        RECT -24.080 117.370 -21.080 117.380 ;
        RECT 112.020 117.370 115.020 117.380 ;
        RECT 292.020 117.370 295.020 117.380 ;
        RECT 472.020 117.370 475.020 117.380 ;
        RECT 652.020 117.370 655.020 117.380 ;
        RECT 832.020 117.370 835.020 117.380 ;
        RECT 1012.020 117.370 1015.020 117.380 ;
        RECT 1192.020 117.370 1195.020 117.380 ;
        RECT 1372.020 117.370 1375.020 117.380 ;
        RECT 1552.020 117.370 1555.020 117.380 ;
        RECT 1732.020 117.370 1735.020 117.380 ;
        RECT 1912.020 117.370 1915.020 117.380 ;
        RECT 2092.020 117.370 2095.020 117.380 ;
        RECT 2272.020 117.370 2275.020 117.380 ;
        RECT 2452.020 117.370 2455.020 117.380 ;
        RECT 2632.020 117.370 2635.020 117.380 ;
        RECT 2812.020 117.370 2815.020 117.380 ;
        RECT 2940.700 117.370 2943.700 117.380 ;
        RECT -14.680 102.380 -11.680 102.390 ;
        RECT 94.020 102.380 97.020 102.390 ;
        RECT 274.020 102.380 277.020 102.390 ;
        RECT 454.020 102.380 457.020 102.390 ;
        RECT 634.020 102.380 637.020 102.390 ;
        RECT 814.020 102.380 817.020 102.390 ;
        RECT 994.020 102.380 997.020 102.390 ;
        RECT 1174.020 102.380 1177.020 102.390 ;
        RECT 1354.020 102.380 1357.020 102.390 ;
        RECT 1534.020 102.380 1537.020 102.390 ;
        RECT 1714.020 102.380 1717.020 102.390 ;
        RECT 1894.020 102.380 1897.020 102.390 ;
        RECT 2074.020 102.380 2077.020 102.390 ;
        RECT 2254.020 102.380 2257.020 102.390 ;
        RECT 2434.020 102.380 2437.020 102.390 ;
        RECT 2614.020 102.380 2617.020 102.390 ;
        RECT 2794.020 102.380 2797.020 102.390 ;
        RECT 2931.300 102.380 2934.300 102.390 ;
        RECT -14.680 99.380 2934.300 102.380 ;
        RECT -14.680 99.370 -11.680 99.380 ;
        RECT 94.020 99.370 97.020 99.380 ;
        RECT 274.020 99.370 277.020 99.380 ;
        RECT 454.020 99.370 457.020 99.380 ;
        RECT 634.020 99.370 637.020 99.380 ;
        RECT 814.020 99.370 817.020 99.380 ;
        RECT 994.020 99.370 997.020 99.380 ;
        RECT 1174.020 99.370 1177.020 99.380 ;
        RECT 1354.020 99.370 1357.020 99.380 ;
        RECT 1534.020 99.370 1537.020 99.380 ;
        RECT 1714.020 99.370 1717.020 99.380 ;
        RECT 1894.020 99.370 1897.020 99.380 ;
        RECT 2074.020 99.370 2077.020 99.380 ;
        RECT 2254.020 99.370 2257.020 99.380 ;
        RECT 2434.020 99.370 2437.020 99.380 ;
        RECT 2614.020 99.370 2617.020 99.380 ;
        RECT 2794.020 99.370 2797.020 99.380 ;
        RECT 2931.300 99.370 2934.300 99.380 ;
        RECT -14.680 -6.320 -11.680 -6.310 ;
        RECT 94.020 -6.320 97.020 -6.310 ;
        RECT 274.020 -6.320 277.020 -6.310 ;
        RECT 454.020 -6.320 457.020 -6.310 ;
        RECT 634.020 -6.320 637.020 -6.310 ;
        RECT 814.020 -6.320 817.020 -6.310 ;
        RECT 994.020 -6.320 997.020 -6.310 ;
        RECT 1174.020 -6.320 1177.020 -6.310 ;
        RECT 1354.020 -6.320 1357.020 -6.310 ;
        RECT 1534.020 -6.320 1537.020 -6.310 ;
        RECT 1714.020 -6.320 1717.020 -6.310 ;
        RECT 1894.020 -6.320 1897.020 -6.310 ;
        RECT 2074.020 -6.320 2077.020 -6.310 ;
        RECT 2254.020 -6.320 2257.020 -6.310 ;
        RECT 2434.020 -6.320 2437.020 -6.310 ;
        RECT 2614.020 -6.320 2617.020 -6.310 ;
        RECT 2794.020 -6.320 2797.020 -6.310 ;
        RECT 2931.300 -6.320 2934.300 -6.310 ;
        RECT -14.680 -9.320 2934.300 -6.320 ;
        RECT -14.680 -9.330 -11.680 -9.320 ;
        RECT 94.020 -9.330 97.020 -9.320 ;
        RECT 274.020 -9.330 277.020 -9.320 ;
        RECT 454.020 -9.330 457.020 -9.320 ;
        RECT 634.020 -9.330 637.020 -9.320 ;
        RECT 814.020 -9.330 817.020 -9.320 ;
        RECT 994.020 -9.330 997.020 -9.320 ;
        RECT 1174.020 -9.330 1177.020 -9.320 ;
        RECT 1354.020 -9.330 1357.020 -9.320 ;
        RECT 1534.020 -9.330 1537.020 -9.320 ;
        RECT 1714.020 -9.330 1717.020 -9.320 ;
        RECT 1894.020 -9.330 1897.020 -9.320 ;
        RECT 2074.020 -9.330 2077.020 -9.320 ;
        RECT 2254.020 -9.330 2257.020 -9.320 ;
        RECT 2434.020 -9.330 2437.020 -9.320 ;
        RECT 2614.020 -9.330 2617.020 -9.320 ;
        RECT 2794.020 -9.330 2797.020 -9.320 ;
        RECT 2931.300 -9.330 2934.300 -9.320 ;
        RECT -24.080 -15.720 -21.080 -15.710 ;
        RECT 112.020 -15.720 115.020 -15.710 ;
        RECT 292.020 -15.720 295.020 -15.710 ;
        RECT 472.020 -15.720 475.020 -15.710 ;
        RECT 652.020 -15.720 655.020 -15.710 ;
        RECT 832.020 -15.720 835.020 -15.710 ;
        RECT 1012.020 -15.720 1015.020 -15.710 ;
        RECT 1192.020 -15.720 1195.020 -15.710 ;
        RECT 1372.020 -15.720 1375.020 -15.710 ;
        RECT 1552.020 -15.720 1555.020 -15.710 ;
        RECT 1732.020 -15.720 1735.020 -15.710 ;
        RECT 1912.020 -15.720 1915.020 -15.710 ;
        RECT 2092.020 -15.720 2095.020 -15.710 ;
        RECT 2272.020 -15.720 2275.020 -15.710 ;
        RECT 2452.020 -15.720 2455.020 -15.710 ;
        RECT 2632.020 -15.720 2635.020 -15.710 ;
        RECT 2812.020 -15.720 2815.020 -15.710 ;
        RECT 2940.700 -15.720 2943.700 -15.710 ;
        RECT -24.080 -18.720 2943.700 -15.720 ;
        RECT -24.080 -18.730 -21.080 -18.720 ;
        RECT 112.020 -18.730 115.020 -18.720 ;
        RECT 292.020 -18.730 295.020 -18.720 ;
        RECT 472.020 -18.730 475.020 -18.720 ;
        RECT 652.020 -18.730 655.020 -18.720 ;
        RECT 832.020 -18.730 835.020 -18.720 ;
        RECT 1012.020 -18.730 1015.020 -18.720 ;
        RECT 1192.020 -18.730 1195.020 -18.720 ;
        RECT 1372.020 -18.730 1375.020 -18.720 ;
        RECT 1552.020 -18.730 1555.020 -18.720 ;
        RECT 1732.020 -18.730 1735.020 -18.720 ;
        RECT 1912.020 -18.730 1915.020 -18.720 ;
        RECT 2092.020 -18.730 2095.020 -18.720 ;
        RECT 2272.020 -18.730 2275.020 -18.720 ;
        RECT 2452.020 -18.730 2455.020 -18.720 ;
        RECT 2632.020 -18.730 2635.020 -18.720 ;
        RECT 2812.020 -18.730 2815.020 -18.720 ;
        RECT 2940.700 -18.730 2943.700 -18.720 ;
        RECT -33.480 -25.120 -30.480 -25.110 ;
        RECT 130.020 -25.120 133.020 -25.110 ;
        RECT 310.020 -25.120 313.020 -25.110 ;
        RECT 490.020 -25.120 493.020 -25.110 ;
        RECT 670.020 -25.120 673.020 -25.110 ;
        RECT 850.020 -25.120 853.020 -25.110 ;
        RECT 1030.020 -25.120 1033.020 -25.110 ;
        RECT 1210.020 -25.120 1213.020 -25.110 ;
        RECT 1390.020 -25.120 1393.020 -25.110 ;
        RECT 1570.020 -25.120 1573.020 -25.110 ;
        RECT 1750.020 -25.120 1753.020 -25.110 ;
        RECT 1930.020 -25.120 1933.020 -25.110 ;
        RECT 2110.020 -25.120 2113.020 -25.110 ;
        RECT 2290.020 -25.120 2293.020 -25.110 ;
        RECT 2470.020 -25.120 2473.020 -25.110 ;
        RECT 2650.020 -25.120 2653.020 -25.110 ;
        RECT 2830.020 -25.120 2833.020 -25.110 ;
        RECT 2950.100 -25.120 2953.100 -25.110 ;
        RECT -33.480 -28.120 2953.100 -25.120 ;
        RECT -33.480 -28.130 -30.480 -28.120 ;
        RECT 130.020 -28.130 133.020 -28.120 ;
        RECT 310.020 -28.130 313.020 -28.120 ;
        RECT 490.020 -28.130 493.020 -28.120 ;
        RECT 670.020 -28.130 673.020 -28.120 ;
        RECT 850.020 -28.130 853.020 -28.120 ;
        RECT 1030.020 -28.130 1033.020 -28.120 ;
        RECT 1210.020 -28.130 1213.020 -28.120 ;
        RECT 1390.020 -28.130 1393.020 -28.120 ;
        RECT 1570.020 -28.130 1573.020 -28.120 ;
        RECT 1750.020 -28.130 1753.020 -28.120 ;
        RECT 1930.020 -28.130 1933.020 -28.120 ;
        RECT 2110.020 -28.130 2113.020 -28.120 ;
        RECT 2290.020 -28.130 2293.020 -28.120 ;
        RECT 2470.020 -28.130 2473.020 -28.120 ;
        RECT 2650.020 -28.130 2653.020 -28.120 ;
        RECT 2830.020 -28.130 2833.020 -28.120 ;
        RECT 2950.100 -28.130 2953.100 -28.120 ;
        RECT -42.880 -34.520 -39.880 -34.510 ;
        RECT 148.020 -34.520 151.020 -34.510 ;
        RECT 328.020 -34.520 331.020 -34.510 ;
        RECT 508.020 -34.520 511.020 -34.510 ;
        RECT 688.020 -34.520 691.020 -34.510 ;
        RECT 868.020 -34.520 871.020 -34.510 ;
        RECT 1048.020 -34.520 1051.020 -34.510 ;
        RECT 1228.020 -34.520 1231.020 -34.510 ;
        RECT 1408.020 -34.520 1411.020 -34.510 ;
        RECT 1588.020 -34.520 1591.020 -34.510 ;
        RECT 1768.020 -34.520 1771.020 -34.510 ;
        RECT 1948.020 -34.520 1951.020 -34.510 ;
        RECT 2128.020 -34.520 2131.020 -34.510 ;
        RECT 2308.020 -34.520 2311.020 -34.510 ;
        RECT 2488.020 -34.520 2491.020 -34.510 ;
        RECT 2668.020 -34.520 2671.020 -34.510 ;
        RECT 2848.020 -34.520 2851.020 -34.510 ;
        RECT 2959.500 -34.520 2962.500 -34.510 ;
        RECT -42.880 -37.520 2962.500 -34.520 ;
        RECT -42.880 -37.530 -39.880 -37.520 ;
        RECT 148.020 -37.530 151.020 -37.520 ;
        RECT 328.020 -37.530 331.020 -37.520 ;
        RECT 508.020 -37.530 511.020 -37.520 ;
        RECT 688.020 -37.530 691.020 -37.520 ;
        RECT 868.020 -37.530 871.020 -37.520 ;
        RECT 1048.020 -37.530 1051.020 -37.520 ;
        RECT 1228.020 -37.530 1231.020 -37.520 ;
        RECT 1408.020 -37.530 1411.020 -37.520 ;
        RECT 1588.020 -37.530 1591.020 -37.520 ;
        RECT 1768.020 -37.530 1771.020 -37.520 ;
        RECT 1948.020 -37.530 1951.020 -37.520 ;
        RECT 2128.020 -37.530 2131.020 -37.520 ;
        RECT 2308.020 -37.530 2311.020 -37.520 ;
        RECT 2488.020 -37.530 2491.020 -37.520 ;
        RECT 2668.020 -37.530 2671.020 -37.520 ;
        RECT 2848.020 -37.530 2851.020 -37.520 ;
        RECT 2959.500 -37.530 2962.500 -37.520 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 305.000 2805.000 681.480 3251.235 ;
        RECT 955.000 2805.000 1331.480 3251.235 ;
        RECT 1555.000 2805.000 1931.480 3251.235 ;
        RECT 2205.000 2805.000 2581.480 3251.235 ;
        RECT 305.520 1510.795 1394.340 2688.725 ;
      LAYER met1 ;
        RECT 2539.270 3266.960 2539.590 3267.020 ;
        RECT 2566.870 3266.960 2567.190 3267.020 ;
        RECT 2539.270 3266.820 2567.190 3266.960 ;
        RECT 2539.270 3266.760 2539.590 3266.820 ;
        RECT 2566.870 3266.760 2567.190 3266.820 ;
        RECT 2566.870 3264.240 2567.190 3264.300 ;
        RECT 2594.470 3264.240 2594.790 3264.300 ;
        RECT 2566.870 3264.100 2594.790 3264.240 ;
        RECT 2566.870 3264.040 2567.190 3264.100 ;
        RECT 2594.470 3264.040 2594.790 3264.100 ;
        RECT 646.370 3263.900 646.690 3263.960 ;
        RECT 667.990 3263.900 668.310 3263.960 ;
        RECT 697.890 3263.900 698.210 3263.960 ;
        RECT 1295.890 3263.900 1296.210 3263.960 ;
        RECT 1318.890 3263.900 1319.210 3263.960 ;
        RECT 1345.570 3263.900 1345.890 3263.960 ;
        RECT 1892.510 3263.900 1892.830 3263.960 ;
        RECT 1917.350 3263.900 1917.670 3263.960 ;
        RECT 1946.790 3263.900 1947.110 3263.960 ;
        RECT 2539.270 3263.900 2539.590 3263.960 ;
        RECT 646.370 3263.760 2539.590 3263.900 ;
        RECT 646.370 3263.700 646.690 3263.760 ;
        RECT 667.990 3263.700 668.310 3263.760 ;
        RECT 697.890 3263.700 698.210 3263.760 ;
        RECT 1295.890 3263.700 1296.210 3263.760 ;
        RECT 1318.890 3263.700 1319.210 3263.760 ;
        RECT 1345.570 3263.700 1345.890 3263.760 ;
        RECT 1892.510 3263.700 1892.830 3263.760 ;
        RECT 1917.350 3263.700 1917.670 3263.760 ;
        RECT 1946.790 3263.700 1947.110 3263.760 ;
        RECT 2539.270 3263.700 2539.590 3263.760 ;
        RECT 696.970 3252.000 697.290 3252.060 ;
        RECT 1331.770 3252.000 1332.090 3252.060 ;
        RECT 696.970 3251.860 1332.090 3252.000 ;
        RECT 696.970 3251.800 697.290 3251.860 ;
        RECT 1331.770 3251.800 1332.090 3251.860 ;
        RECT 1409.970 3252.000 1410.290 3252.060 ;
        RECT 1945.870 3252.000 1946.190 3252.060 ;
        RECT 2582.050 3252.000 2582.370 3252.060 ;
        RECT 1409.970 3251.860 2582.370 3252.000 ;
        RECT 1409.970 3251.800 1410.290 3251.860 ;
        RECT 1945.870 3251.800 1946.190 3251.860 ;
        RECT 2582.050 3251.800 2582.370 3251.860 ;
      LAYER met1 ;
        RECT 305.000 2805.000 681.480 3251.235 ;
      LAYER met1 ;
        RECT 710.310 3229.560 710.630 3229.620 ;
        RECT 938.470 3229.560 938.790 3229.620 ;
        RECT 710.310 3229.420 938.790 3229.560 ;
        RECT 710.310 3229.360 710.630 3229.420 ;
        RECT 938.470 3229.360 938.790 3229.420 ;
        RECT 703.410 3222.420 703.730 3222.480 ;
        RECT 938.470 3222.420 938.790 3222.480 ;
        RECT 703.410 3222.280 938.790 3222.420 ;
        RECT 703.410 3222.220 703.730 3222.280 ;
        RECT 938.470 3222.220 938.790 3222.280 ;
        RECT 689.610 3215.620 689.930 3215.680 ;
        RECT 938.470 3215.620 938.790 3215.680 ;
        RECT 689.610 3215.480 938.790 3215.620 ;
        RECT 689.610 3215.420 689.930 3215.480 ;
        RECT 938.470 3215.420 938.790 3215.480 ;
        RECT 803.690 3208.820 804.010 3208.880 ;
        RECT 938.470 3208.820 938.790 3208.880 ;
        RECT 803.690 3208.680 938.790 3208.820 ;
        RECT 803.690 3208.620 804.010 3208.680 ;
        RECT 938.470 3208.620 938.790 3208.680 ;
        RECT 796.790 3201.680 797.110 3201.740 ;
        RECT 938.470 3201.680 938.790 3201.740 ;
        RECT 796.790 3201.540 938.790 3201.680 ;
        RECT 796.790 3201.480 797.110 3201.540 ;
        RECT 938.470 3201.480 938.790 3201.540 ;
        RECT 889.710 2898.400 890.030 2898.460 ;
        RECT 938.470 2898.400 938.790 2898.460 ;
        RECT 889.710 2898.260 938.790 2898.400 ;
        RECT 889.710 2898.200 890.030 2898.260 ;
        RECT 938.470 2898.200 938.790 2898.260 ;
      LAYER met1 ;
        RECT 955.000 2805.000 1331.480 3251.235 ;
      LAYER met1 ;
        RECT 1331.770 3250.300 1332.090 3250.360 ;
        RECT 1407.670 3250.300 1407.990 3250.360 ;
        RECT 1409.970 3250.300 1410.290 3250.360 ;
        RECT 1331.770 3250.160 1410.290 3250.300 ;
        RECT 1331.770 3250.100 1332.090 3250.160 ;
        RECT 1407.670 3250.100 1407.990 3250.160 ;
        RECT 1409.970 3250.100 1410.290 3250.160 ;
        RECT 1459.650 3229.560 1459.970 3229.620 ;
        RECT 1536.930 3229.560 1537.250 3229.620 ;
        RECT 1459.650 3229.420 1537.250 3229.560 ;
        RECT 1459.650 3229.360 1459.970 3229.420 ;
        RECT 1536.930 3229.360 1537.250 3229.420 ;
        RECT 1452.750 3222.420 1453.070 3222.480 ;
        RECT 1535.550 3222.420 1535.870 3222.480 ;
        RECT 1452.750 3222.280 1535.870 3222.420 ;
        RECT 1452.750 3222.220 1453.070 3222.280 ;
        RECT 1535.550 3222.220 1535.870 3222.280 ;
        RECT 1438.490 3215.620 1438.810 3215.680 ;
        RECT 1535.550 3215.620 1535.870 3215.680 ;
        RECT 1438.490 3215.480 1535.870 3215.620 ;
        RECT 1438.490 3215.420 1438.810 3215.480 ;
        RECT 1535.550 3215.420 1535.870 3215.480 ;
        RECT 1431.590 3208.820 1431.910 3208.880 ;
        RECT 1538.310 3208.820 1538.630 3208.880 ;
        RECT 1431.590 3208.680 1538.630 3208.820 ;
        RECT 1431.590 3208.620 1431.910 3208.680 ;
        RECT 1538.310 3208.620 1538.630 3208.680 ;
        RECT 1424.690 3201.680 1425.010 3201.740 ;
        RECT 1538.310 3201.680 1538.630 3201.740 ;
        RECT 1424.690 3201.540 1538.630 3201.680 ;
        RECT 1424.690 3201.480 1425.010 3201.540 ;
        RECT 1538.310 3201.480 1538.630 3201.540 ;
        RECT 1417.790 3194.880 1418.110 3194.940 ;
        RECT 1533.250 3194.880 1533.570 3194.940 ;
        RECT 1417.790 3194.740 1533.570 3194.880 ;
        RECT 1417.790 3194.680 1418.110 3194.740 ;
        RECT 1533.250 3194.680 1533.570 3194.740 ;
        RECT 1472.990 3188.080 1473.310 3188.140 ;
        RECT 1497.830 3188.080 1498.150 3188.140 ;
        RECT 1472.990 3187.940 1498.150 3188.080 ;
        RECT 1472.990 3187.880 1473.310 3187.940 ;
        RECT 1497.830 3187.880 1498.150 3187.940 ;
        RECT 1350.170 2901.460 1350.490 2901.520 ;
        RECT 1408.130 2901.460 1408.450 2901.520 ;
        RECT 1350.170 2901.320 1408.450 2901.460 ;
        RECT 1350.170 2901.260 1350.490 2901.320 ;
        RECT 1408.130 2901.260 1408.450 2901.320 ;
        RECT 1425.150 2898.400 1425.470 2898.460 ;
        RECT 1534.630 2898.400 1534.950 2898.460 ;
        RECT 1425.150 2898.260 1534.950 2898.400 ;
        RECT 1425.150 2898.200 1425.470 2898.260 ;
        RECT 1534.630 2898.200 1534.950 2898.260 ;
        RECT 1410.890 2891.260 1411.210 2891.320 ;
        RECT 1531.870 2891.260 1532.190 2891.320 ;
        RECT 1410.890 2891.120 1532.190 2891.260 ;
        RECT 1410.890 2891.060 1411.210 2891.120 ;
        RECT 1531.870 2891.060 1532.190 2891.120 ;
        RECT 1408.590 2808.300 1408.910 2808.360 ;
        RECT 1410.890 2808.300 1411.210 2808.360 ;
        RECT 1408.590 2808.160 1411.210 2808.300 ;
        RECT 1408.590 2808.100 1408.910 2808.160 ;
        RECT 1410.890 2808.100 1411.210 2808.160 ;
      LAYER met1 ;
        RECT 1555.000 2805.000 1931.480 3251.235 ;
      LAYER met1 ;
        RECT 1997.390 3229.560 1997.710 3229.620 ;
        RECT 2187.370 3229.560 2187.690 3229.620 ;
        RECT 1997.390 3229.420 2187.690 3229.560 ;
        RECT 1997.390 3229.360 1997.710 3229.420 ;
        RECT 2187.370 3229.360 2187.690 3229.420 ;
        RECT 1990.490 3222.420 1990.810 3222.480 ;
        RECT 2187.370 3222.420 2187.690 3222.480 ;
        RECT 1990.490 3222.280 2187.690 3222.420 ;
        RECT 1990.490 3222.220 1990.810 3222.280 ;
        RECT 2187.370 3222.220 2187.690 3222.280 ;
        RECT 1976.690 3215.620 1977.010 3215.680 ;
        RECT 2187.370 3215.620 2187.690 3215.680 ;
        RECT 1976.690 3215.480 2187.690 3215.620 ;
        RECT 1976.690 3215.420 1977.010 3215.480 ;
        RECT 2187.370 3215.420 2187.690 3215.480 ;
        RECT 1969.790 3208.820 1970.110 3208.880 ;
        RECT 2187.370 3208.820 2187.690 3208.880 ;
        RECT 1969.790 3208.680 2187.690 3208.820 ;
        RECT 1969.790 3208.620 1970.110 3208.680 ;
        RECT 2187.370 3208.620 2187.690 3208.680 ;
        RECT 1962.890 3201.680 1963.210 3201.740 ;
        RECT 2187.370 3201.680 2187.690 3201.740 ;
        RECT 1962.890 3201.540 2187.690 3201.680 ;
        RECT 1962.890 3201.480 1963.210 3201.540 ;
        RECT 2187.370 3201.480 2187.690 3201.540 ;
        RECT 1955.990 3194.880 1956.310 3194.940 ;
        RECT 2187.370 3194.880 2187.690 3194.940 ;
        RECT 1955.990 3194.740 2187.690 3194.880 ;
        RECT 1955.990 3194.680 1956.310 3194.740 ;
        RECT 2187.370 3194.680 2187.690 3194.740 ;
        RECT 2125.360 3188.280 2147.580 3188.420 ;
        RECT 1942.190 3188.080 1942.510 3188.140 ;
        RECT 2125.360 3188.080 2125.500 3188.280 ;
        RECT 1942.190 3187.940 2125.500 3188.080 ;
        RECT 2147.440 3188.080 2147.580 3188.280 ;
        RECT 2187.370 3188.080 2187.690 3188.140 ;
        RECT 2147.440 3187.940 2187.690 3188.080 ;
        RECT 1942.190 3187.880 1942.510 3187.940 ;
        RECT 2187.370 3187.880 2187.690 3187.940 ;
        RECT 2011.190 2898.400 2011.510 2898.460 ;
        RECT 2187.370 2898.400 2187.690 2898.460 ;
        RECT 2011.190 2898.260 2187.690 2898.400 ;
        RECT 2011.190 2898.200 2011.510 2898.260 ;
        RECT 2187.370 2898.200 2187.690 2898.260 ;
      LAYER met1 ;
        RECT 2205.000 2805.000 2581.480 3251.235 ;
      LAYER met1 ;
        RECT 298.150 2804.560 298.470 2804.620 ;
        RECT 944.910 2804.560 945.230 2804.620 ;
        RECT 1408.590 2804.560 1408.910 2804.620 ;
        RECT 298.150 2804.420 1408.910 2804.560 ;
        RECT 298.150 2804.360 298.470 2804.420 ;
        RECT 944.910 2804.360 945.230 2804.420 ;
        RECT 1408.590 2804.360 1408.910 2804.420 ;
        RECT 1531.410 2804.560 1531.730 2804.620 ;
        RECT 2190.590 2804.560 2190.910 2804.620 ;
        RECT 1531.410 2804.420 2190.910 2804.560 ;
        RECT 1531.410 2804.360 1531.730 2804.420 ;
        RECT 2190.590 2804.360 2190.910 2804.420 ;
        RECT 396.590 2794.360 396.910 2794.420 ;
        RECT 407.170 2794.360 407.490 2794.420 ;
        RECT 396.590 2794.220 407.490 2794.360 ;
        RECT 396.590 2794.160 396.910 2794.220 ;
        RECT 407.170 2794.160 407.490 2794.220 ;
        RECT 407.630 2794.360 407.950 2794.420 ;
        RECT 434.310 2794.360 434.630 2794.420 ;
        RECT 450.410 2794.360 450.730 2794.420 ;
        RECT 455.010 2794.360 455.330 2794.420 ;
        RECT 407.630 2794.220 434.630 2794.360 ;
        RECT 407.630 2794.160 407.950 2794.220 ;
        RECT 434.310 2794.160 434.630 2794.220 ;
        RECT 439.000 2794.220 455.330 2794.360 ;
        RECT 403.490 2794.020 403.810 2794.080 ;
        RECT 439.000 2794.020 439.140 2794.220 ;
        RECT 450.410 2794.160 450.730 2794.220 ;
        RECT 455.010 2794.160 455.330 2794.220 ;
        RECT 1677.230 2794.360 1677.550 2794.420 ;
        RECT 1721.390 2794.360 1721.710 2794.420 ;
        RECT 1677.230 2794.220 1721.710 2794.360 ;
        RECT 1677.230 2794.160 1677.550 2794.220 ;
        RECT 1721.390 2794.160 1721.710 2794.220 ;
        RECT 1776.590 2794.360 1776.910 2794.420 ;
        RECT 2415.070 2794.360 2415.390 2794.420 ;
        RECT 1776.590 2794.220 2415.390 2794.360 ;
        RECT 1776.590 2794.160 1776.910 2794.220 ;
        RECT 2415.070 2794.160 2415.390 2794.220 ;
        RECT 403.490 2793.880 439.140 2794.020 ;
        RECT 439.370 2794.020 439.690 2794.080 ;
        RECT 483.070 2794.020 483.390 2794.080 ;
        RECT 439.370 2793.880 483.390 2794.020 ;
        RECT 403.490 2793.820 403.810 2793.880 ;
        RECT 439.370 2793.820 439.690 2793.880 ;
        RECT 483.070 2793.820 483.390 2793.880 ;
        RECT 1117.870 2794.020 1118.190 2794.080 ;
        RECT 1159.730 2794.020 1160.050 2794.080 ;
        RECT 1117.870 2793.880 1160.050 2794.020 ;
        RECT 1117.870 2793.820 1118.190 2793.880 ;
        RECT 1159.730 2793.820 1160.050 2793.880 ;
        RECT 1718.630 2794.020 1718.950 2794.080 ;
        RECT 1759.570 2794.020 1759.890 2794.080 ;
        RECT 1718.630 2793.880 1759.890 2794.020 ;
        RECT 1718.630 2793.820 1718.950 2793.880 ;
        RECT 1759.570 2793.820 1759.890 2793.880 ;
        RECT 2294.090 2794.020 2294.410 2794.080 ;
        RECT 2340.090 2794.020 2340.410 2794.080 ;
        RECT 2385.630 2794.020 2385.950 2794.080 ;
        RECT 2428.870 2794.020 2429.190 2794.080 ;
        RECT 2294.090 2793.880 2429.190 2794.020 ;
        RECT 2294.090 2793.820 2294.410 2793.880 ;
        RECT 2340.090 2793.820 2340.410 2793.880 ;
        RECT 2385.630 2793.820 2385.950 2793.880 ;
        RECT 2428.870 2793.820 2429.190 2793.880 ;
        RECT 397.510 2793.680 397.830 2793.740 ;
        RECT 444.890 2793.680 445.210 2793.740 ;
        RECT 501.470 2793.680 501.790 2793.740 ;
        RECT 397.510 2793.540 445.210 2793.680 ;
        RECT 397.510 2793.480 397.830 2793.540 ;
        RECT 444.890 2793.480 445.210 2793.540 ;
        RECT 467.520 2793.540 501.790 2793.680 ;
        RECT 386.930 2793.340 387.250 2793.400 ;
        RECT 407.630 2793.340 407.950 2793.400 ;
        RECT 386.930 2793.200 407.950 2793.340 ;
        RECT 386.930 2793.140 387.250 2793.200 ;
        RECT 407.630 2793.140 407.950 2793.200 ;
        RECT 408.090 2793.340 408.410 2793.400 ;
        RECT 456.850 2793.340 457.170 2793.400 ;
        RECT 467.520 2793.340 467.660 2793.540 ;
        RECT 501.470 2793.480 501.790 2793.540 ;
        RECT 1083.830 2793.680 1084.150 2793.740 ;
        RECT 1128.910 2793.680 1129.230 2793.740 ;
        RECT 1083.830 2793.540 1129.230 2793.680 ;
        RECT 1083.830 2793.480 1084.150 2793.540 ;
        RECT 1128.910 2793.480 1129.230 2793.540 ;
        RECT 1131.670 2793.680 1131.990 2793.740 ;
        RECT 1135.810 2793.680 1136.130 2793.740 ;
        RECT 1179.970 2793.680 1180.290 2793.740 ;
        RECT 1131.670 2793.540 1180.290 2793.680 ;
        RECT 1131.670 2793.480 1131.990 2793.540 ;
        RECT 1135.810 2793.480 1136.130 2793.540 ;
        RECT 1179.970 2793.480 1180.290 2793.540 ;
        RECT 1721.390 2793.680 1721.710 2793.740 ;
        RECT 1766.470 2793.680 1766.790 2793.740 ;
        RECT 1721.390 2793.540 1766.790 2793.680 ;
        RECT 1721.390 2793.480 1721.710 2793.540 ;
        RECT 1766.470 2793.480 1766.790 2793.540 ;
        RECT 2303.290 2793.680 2303.610 2793.740 ;
        RECT 2342.850 2793.680 2343.170 2793.740 ;
        RECT 2303.290 2793.540 2343.170 2793.680 ;
        RECT 2303.290 2793.480 2303.610 2793.540 ;
        RECT 2342.850 2793.480 2343.170 2793.540 ;
        RECT 2377.810 2793.680 2378.130 2793.740 ;
        RECT 2421.970 2793.680 2422.290 2793.740 ;
        RECT 2377.810 2793.540 2422.290 2793.680 ;
        RECT 2377.810 2793.480 2378.130 2793.540 ;
        RECT 2421.970 2793.480 2422.290 2793.540 ;
        RECT 408.090 2793.200 467.660 2793.340 ;
        RECT 476.630 2793.340 476.950 2793.400 ;
        RECT 526.770 2793.340 527.090 2793.400 ;
        RECT 530.450 2793.340 530.770 2793.400 ;
        RECT 476.630 2793.200 530.770 2793.340 ;
        RECT 408.090 2793.140 408.410 2793.200 ;
        RECT 456.850 2793.140 457.170 2793.200 ;
        RECT 476.630 2793.140 476.950 2793.200 ;
        RECT 526.770 2793.140 527.090 2793.200 ;
        RECT 530.450 2793.140 530.770 2793.200 ;
        RECT 1076.470 2793.340 1076.790 2793.400 ;
        RECT 1122.010 2793.340 1122.330 2793.400 ;
        RECT 1166.170 2793.340 1166.490 2793.400 ;
        RECT 1076.470 2793.200 1166.490 2793.340 ;
        RECT 1076.470 2793.140 1076.790 2793.200 ;
        RECT 1122.010 2793.140 1122.330 2793.200 ;
        RECT 1166.170 2793.140 1166.490 2793.200 ;
        RECT 1694.710 2793.340 1695.030 2793.400 ;
        RECT 1741.630 2793.340 1741.950 2793.400 ;
        RECT 1787.170 2793.340 1787.490 2793.400 ;
        RECT 2422.430 2793.340 2422.750 2793.400 ;
        RECT 1694.710 2793.200 1787.490 2793.340 ;
        RECT 1694.710 2793.140 1695.030 2793.200 ;
        RECT 1741.630 2793.140 1741.950 2793.200 ;
        RECT 1787.170 2793.140 1787.490 2793.200 ;
        RECT 1787.720 2793.200 2422.750 2793.340 ;
        RECT 378.650 2793.000 378.970 2793.060 ;
        RECT 421.430 2793.000 421.750 2793.060 ;
        RECT 467.890 2793.000 468.210 2793.060 ;
        RECT 378.650 2792.860 468.210 2793.000 ;
        RECT 378.650 2792.800 378.970 2792.860 ;
        RECT 421.430 2792.800 421.750 2792.860 ;
        RECT 467.890 2792.800 468.210 2792.860 ;
        RECT 542.870 2793.000 543.190 2793.060 ;
        RECT 1056.690 2793.000 1057.010 2793.060 ;
        RECT 542.870 2792.860 1057.010 2793.000 ;
        RECT 542.870 2792.800 543.190 2792.860 ;
        RECT 1056.690 2792.800 1057.010 2792.860 ;
        RECT 1062.670 2793.000 1062.990 2793.060 ;
        RECT 1065.890 2793.000 1066.210 2793.060 ;
        RECT 1111.430 2793.000 1111.750 2793.060 ;
        RECT 1159.270 2793.000 1159.590 2793.060 ;
        RECT 1062.670 2792.860 1159.590 2793.000 ;
        RECT 1062.670 2792.800 1062.990 2792.860 ;
        RECT 1065.890 2792.800 1066.210 2792.860 ;
        RECT 1111.430 2792.800 1111.750 2792.860 ;
        RECT 1159.270 2792.800 1159.590 2792.860 ;
        RECT 1683.210 2793.000 1683.530 2793.060 ;
        RECT 1731.510 2793.000 1731.830 2793.060 ;
        RECT 1734.730 2793.000 1735.050 2793.060 ;
        RECT 1780.270 2793.000 1780.590 2793.060 ;
        RECT 1683.210 2792.860 1731.830 2793.000 ;
        RECT 1734.295 2792.860 1780.590 2793.000 ;
        RECT 1683.210 2792.800 1683.530 2792.860 ;
        RECT 1731.510 2792.800 1731.830 2792.860 ;
        RECT 1734.730 2792.800 1735.050 2792.860 ;
        RECT 1780.270 2792.800 1780.590 2792.860 ;
        RECT 1783.950 2793.000 1784.270 2793.060 ;
        RECT 1787.720 2793.000 1787.860 2793.200 ;
        RECT 2422.430 2793.140 2422.750 2793.200 ;
        RECT 1783.950 2792.860 1787.860 2793.000 ;
        RECT 2267.410 2793.000 2267.730 2793.060 ;
        RECT 2314.790 2793.000 2315.110 2793.060 ;
        RECT 2318.010 2793.000 2318.330 2793.060 ;
        RECT 2267.410 2792.860 2318.330 2793.000 ;
        RECT 1783.950 2792.800 1784.270 2792.860 ;
        RECT 2267.410 2792.800 2267.730 2792.860 ;
        RECT 2314.790 2792.800 2315.110 2792.860 ;
        RECT 2318.010 2792.800 2318.330 2792.860 ;
        RECT 2321.690 2793.000 2322.010 2793.060 ;
        RECT 2367.690 2793.000 2368.010 2793.060 ;
        RECT 2415.070 2793.000 2415.390 2793.060 ;
        RECT 2321.690 2792.860 2415.390 2793.000 ;
        RECT 2321.690 2792.800 2322.010 2792.860 ;
        RECT 2367.690 2792.800 2368.010 2792.860 ;
        RECT 2415.070 2792.800 2415.390 2792.860 ;
        RECT 362.090 2792.660 362.410 2792.720 ;
        RECT 408.090 2792.660 408.410 2792.720 ;
        RECT 362.090 2792.520 408.410 2792.660 ;
        RECT 362.090 2792.460 362.410 2792.520 ;
        RECT 408.090 2792.460 408.410 2792.520 ;
        RECT 434.310 2792.660 434.630 2792.720 ;
        RECT 476.630 2792.660 476.950 2792.720 ;
        RECT 434.310 2792.520 476.950 2792.660 ;
        RECT 434.310 2792.460 434.630 2792.520 ;
        RECT 476.630 2792.460 476.950 2792.520 ;
        RECT 483.070 2792.660 483.390 2792.720 ;
        RECT 531.370 2792.660 531.690 2792.720 ;
        RECT 537.350 2792.660 537.670 2792.720 ;
        RECT 483.070 2792.520 537.670 2792.660 ;
        RECT 483.070 2792.460 483.390 2792.520 ;
        RECT 531.370 2792.460 531.690 2792.520 ;
        RECT 537.350 2792.460 537.670 2792.520 ;
        RECT 539.190 2792.660 539.510 2792.720 ;
        RECT 1048.870 2792.660 1049.190 2792.720 ;
        RECT 539.190 2792.520 1049.190 2792.660 ;
        RECT 539.190 2792.460 539.510 2792.520 ;
        RECT 1048.870 2792.460 1049.190 2792.520 ;
        RECT 1055.770 2792.660 1056.090 2792.720 ;
        RECT 1059.450 2792.660 1059.770 2792.720 ;
        RECT 1105.450 2792.660 1105.770 2792.720 ;
        RECT 1152.370 2792.660 1152.690 2792.720 ;
        RECT 1055.770 2792.520 1152.690 2792.660 ;
        RECT 1055.770 2792.460 1056.090 2792.520 ;
        RECT 1059.450 2792.460 1059.770 2792.520 ;
        RECT 1105.450 2792.460 1105.770 2792.520 ;
        RECT 1152.370 2792.460 1152.690 2792.520 ;
        RECT 1686.890 2792.660 1687.210 2792.720 ;
        RECT 1734.820 2792.660 1734.960 2792.800 ;
        RECT 1686.890 2792.520 1734.960 2792.660 ;
        RECT 2301.910 2792.660 2302.230 2792.720 ;
        RECT 2304.210 2792.660 2304.530 2792.720 ;
        RECT 2350.210 2792.660 2350.530 2792.720 ;
        RECT 2397.130 2792.660 2397.450 2792.720 ;
        RECT 2442.670 2792.660 2442.990 2792.720 ;
        RECT 2301.910 2792.520 2442.990 2792.660 ;
        RECT 1686.890 2792.460 1687.210 2792.520 ;
        RECT 2301.910 2792.460 2302.230 2792.520 ;
        RECT 2304.210 2792.460 2304.530 2792.520 ;
        RECT 2350.210 2792.460 2350.530 2792.520 ;
        RECT 2397.130 2792.460 2397.450 2792.520 ;
        RECT 2442.670 2792.460 2442.990 2792.520 ;
        RECT 380.030 2792.320 380.350 2792.380 ;
        RECT 426.950 2792.320 427.270 2792.380 ;
        RECT 472.950 2792.320 473.270 2792.380 ;
        RECT 519.870 2792.320 520.190 2792.380 ;
        RECT 523.550 2792.320 523.870 2792.380 ;
        RECT 380.030 2792.180 523.870 2792.320 ;
        RECT 380.030 2792.120 380.350 2792.180 ;
        RECT 426.950 2792.120 427.270 2792.180 ;
        RECT 472.950 2792.120 473.270 2792.180 ;
        RECT 519.870 2792.120 520.190 2792.180 ;
        RECT 523.550 2792.120 523.870 2792.180 ;
        RECT 834.510 2792.320 834.830 2792.380 ;
        RECT 1007.470 2792.320 1007.790 2792.380 ;
        RECT 834.510 2792.180 1007.790 2792.320 ;
        RECT 834.510 2792.120 834.830 2792.180 ;
        RECT 1007.470 2792.120 1007.790 2792.180 ;
        RECT 1656.530 2792.320 1656.850 2792.380 ;
        RECT 1658.830 2792.320 1659.150 2792.380 ;
        RECT 1704.830 2792.320 1705.150 2792.380 ;
        RECT 1752.670 2792.320 1752.990 2792.380 ;
        RECT 1656.530 2792.180 1752.990 2792.320 ;
        RECT 1656.530 2792.120 1656.850 2792.180 ;
        RECT 1658.830 2792.120 1659.150 2792.180 ;
        RECT 1704.830 2792.120 1705.150 2792.180 ;
        RECT 1752.670 2792.120 1752.990 2792.180 ;
        RECT 2266.490 2792.320 2266.810 2792.380 ;
        RECT 2308.810 2792.320 2309.130 2792.380 ;
        RECT 2356.190 2792.320 2356.510 2792.380 ;
        RECT 2402.190 2792.320 2402.510 2792.380 ;
        RECT 2266.490 2792.180 2402.510 2792.320 ;
        RECT 2266.490 2792.120 2266.810 2792.180 ;
        RECT 2308.810 2792.120 2309.130 2792.180 ;
        RECT 2356.190 2792.120 2356.510 2792.180 ;
        RECT 2402.190 2792.120 2402.510 2792.180 ;
        RECT 368.530 2791.980 368.850 2792.040 ;
        RECT 414.530 2791.980 414.850 2792.040 ;
        RECT 462.370 2791.980 462.690 2792.040 ;
        RECT 503.770 2791.980 504.090 2792.040 ;
        RECT 368.530 2791.840 504.090 2791.980 ;
        RECT 368.530 2791.780 368.850 2791.840 ;
        RECT 414.530 2791.780 414.850 2791.840 ;
        RECT 462.370 2791.780 462.690 2791.840 ;
        RECT 503.770 2791.780 504.090 2791.840 ;
        RECT 827.610 2791.980 827.930 2792.040 ;
        RECT 1001.030 2791.980 1001.350 2792.040 ;
        RECT 827.610 2791.840 1001.350 2791.980 ;
        RECT 827.610 2791.780 827.930 2791.840 ;
        RECT 1001.030 2791.780 1001.350 2791.840 ;
        RECT 1090.270 2791.980 1090.590 2792.040 ;
        RECT 1094.410 2791.980 1094.730 2792.040 ;
        RECT 1138.570 2791.980 1138.890 2792.040 ;
        RECT 1090.270 2791.840 1138.890 2791.980 ;
        RECT 1090.270 2791.780 1090.590 2791.840 ;
        RECT 1094.410 2791.780 1094.730 2791.840 ;
        RECT 1138.570 2791.780 1138.890 2791.840 ;
        RECT 1139.030 2791.980 1139.350 2792.040 ;
        RECT 1147.310 2791.980 1147.630 2792.040 ;
        RECT 1193.770 2791.980 1194.090 2792.040 ;
        RECT 1139.030 2791.840 1194.090 2791.980 ;
        RECT 1139.030 2791.780 1139.350 2791.840 ;
        RECT 1147.310 2791.780 1147.630 2791.840 ;
        RECT 1193.770 2791.780 1194.090 2791.840 ;
        RECT 1663.430 2791.980 1663.750 2792.040 ;
        RECT 1712.650 2791.980 1712.970 2792.040 ;
        RECT 1739.790 2791.980 1740.110 2792.040 ;
        RECT 1663.430 2791.840 1740.110 2791.980 ;
        RECT 1663.430 2791.780 1663.750 2791.840 ;
        RECT 1712.650 2791.780 1712.970 2791.840 ;
        RECT 1739.790 2791.780 1740.110 2791.840 ;
        RECT 1790.850 2791.980 1791.170 2792.040 ;
        RECT 2277.070 2791.980 2277.390 2792.040 ;
        RECT 1790.850 2791.840 2277.390 2791.980 ;
        RECT 1790.850 2791.780 1791.170 2791.840 ;
        RECT 2277.070 2791.780 2277.390 2791.840 ;
        RECT 2318.010 2791.980 2318.330 2792.040 ;
        RECT 2361.250 2791.980 2361.570 2792.040 ;
        RECT 2408.170 2791.980 2408.490 2792.040 ;
        RECT 2318.010 2791.840 2408.490 2791.980 ;
        RECT 2318.010 2791.780 2318.330 2791.840 ;
        RECT 2361.250 2791.780 2361.570 2791.840 ;
        RECT 2408.170 2791.780 2408.490 2791.840 ;
        RECT 379.110 2791.640 379.430 2791.700 ;
        RECT 400.270 2791.640 400.590 2791.700 ;
        RECT 379.110 2791.500 400.590 2791.640 ;
        RECT 379.110 2791.440 379.430 2791.500 ;
        RECT 400.270 2791.440 400.590 2791.500 ;
        RECT 444.890 2791.640 445.210 2791.700 ;
        RECT 491.350 2791.640 491.670 2791.700 ;
        RECT 539.190 2791.640 539.510 2791.700 ;
        RECT 444.890 2791.500 539.510 2791.640 ;
        RECT 444.890 2791.440 445.210 2791.500 ;
        RECT 491.350 2791.440 491.670 2791.500 ;
        RECT 539.190 2791.440 539.510 2791.500 ;
        RECT 813.810 2791.640 814.130 2791.700 ;
        RECT 993.670 2791.640 993.990 2791.700 ;
        RECT 813.810 2791.500 993.990 2791.640 ;
        RECT 813.810 2791.440 814.130 2791.500 ;
        RECT 993.670 2791.440 993.990 2791.500 ;
        RECT 1069.570 2791.640 1069.890 2791.700 ;
        RECT 1117.870 2791.640 1118.190 2791.700 ;
        RECT 1069.570 2791.500 1118.190 2791.640 ;
        RECT 1069.570 2791.440 1069.890 2791.500 ;
        RECT 1117.870 2791.440 1118.190 2791.500 ;
        RECT 1128.910 2791.640 1129.230 2791.700 ;
        RECT 1173.070 2791.640 1173.390 2791.700 ;
        RECT 1128.910 2791.500 1173.390 2791.640 ;
        RECT 1128.910 2791.440 1129.230 2791.500 ;
        RECT 1173.070 2791.440 1173.390 2791.500 ;
        RECT 1699.310 2791.640 1699.630 2791.700 ;
        RECT 1747.610 2791.640 1747.930 2791.700 ;
        RECT 1788.550 2791.640 1788.870 2791.700 ;
        RECT 1699.310 2791.500 1788.870 2791.640 ;
        RECT 1699.310 2791.440 1699.630 2791.500 ;
        RECT 1747.610 2791.440 1747.930 2791.500 ;
        RECT 1788.550 2791.440 1788.870 2791.500 ;
        RECT 1797.290 2791.640 1797.610 2791.700 ;
        RECT 2283.970 2791.640 2284.290 2791.700 ;
        RECT 1797.290 2791.500 2284.290 2791.640 ;
        RECT 1797.290 2791.440 1797.610 2791.500 ;
        RECT 2283.970 2791.440 2284.290 2791.500 ;
        RECT 2325.830 2791.640 2326.150 2791.700 ;
        RECT 2374.130 2791.640 2374.450 2791.700 ;
        RECT 2325.830 2791.500 2374.450 2791.640 ;
        RECT 2325.830 2791.440 2326.150 2791.500 ;
        RECT 2374.130 2791.440 2374.450 2791.500 ;
        RECT 2387.930 2791.640 2388.250 2791.700 ;
        RECT 2391.610 2791.640 2391.930 2791.700 ;
        RECT 2435.770 2791.640 2436.090 2791.700 ;
        RECT 2387.930 2791.500 2436.090 2791.640 ;
        RECT 2387.930 2791.440 2388.250 2791.500 ;
        RECT 2391.610 2791.440 2391.930 2791.500 ;
        RECT 2435.770 2791.440 2436.090 2791.500 ;
        RECT 392.450 2791.300 392.770 2791.360 ;
        RECT 439.370 2791.300 439.690 2791.360 ;
        RECT 392.450 2791.160 439.690 2791.300 ;
        RECT 392.450 2791.100 392.770 2791.160 ;
        RECT 439.370 2791.100 439.690 2791.160 ;
        RECT 455.010 2791.300 455.330 2791.360 ;
        RECT 497.790 2791.300 498.110 2791.360 ;
        RECT 542.870 2791.300 543.190 2791.360 ;
        RECT 455.010 2791.160 543.190 2791.300 ;
        RECT 455.010 2791.100 455.330 2791.160 ;
        RECT 497.790 2791.100 498.110 2791.160 ;
        RECT 542.870 2791.100 543.190 2791.160 ;
        RECT 806.910 2791.300 807.230 2791.360 ;
        RECT 986.770 2791.300 987.090 2791.360 ;
        RECT 806.910 2791.160 987.090 2791.300 ;
        RECT 806.910 2791.100 807.230 2791.160 ;
        RECT 986.770 2791.100 987.090 2791.160 ;
        RECT 1083.370 2791.300 1083.690 2791.360 ;
        RECT 1087.970 2791.300 1088.290 2791.360 ;
        RECT 1131.670 2791.300 1131.990 2791.360 ;
        RECT 1083.370 2791.160 1131.990 2791.300 ;
        RECT 1083.370 2791.100 1083.690 2791.160 ;
        RECT 1087.970 2791.100 1088.290 2791.160 ;
        RECT 1131.670 2791.100 1131.990 2791.160 ;
        RECT 1138.570 2791.300 1138.890 2791.360 ;
        RECT 1186.870 2791.300 1187.190 2791.360 ;
        RECT 1138.570 2791.160 1187.190 2791.300 ;
        RECT 1138.570 2791.100 1138.890 2791.160 ;
        RECT 1186.870 2791.100 1187.190 2791.160 ;
        RECT 1459.190 2791.300 1459.510 2791.360 ;
        RECT 1649.170 2791.300 1649.490 2791.360 ;
        RECT 1459.190 2791.160 1649.490 2791.300 ;
        RECT 1459.190 2791.100 1459.510 2791.160 ;
        RECT 1649.170 2791.100 1649.490 2791.160 ;
        RECT 1670.330 2791.300 1670.650 2791.360 ;
        RECT 1718.630 2791.300 1718.950 2791.360 ;
        RECT 1670.330 2791.160 1718.950 2791.300 ;
        RECT 1670.330 2791.100 1670.650 2791.160 ;
        RECT 1718.630 2791.100 1718.950 2791.160 ;
        RECT 1731.510 2791.300 1731.830 2791.360 ;
        RECT 1773.370 2791.300 1773.690 2791.360 ;
        RECT 1731.510 2791.160 1773.690 2791.300 ;
        RECT 1731.510 2791.100 1731.830 2791.160 ;
        RECT 1773.370 2791.100 1773.690 2791.160 ;
        RECT 1797.750 2791.300 1798.070 2791.360 ;
        RECT 2290.870 2791.300 2291.190 2791.360 ;
        RECT 1797.750 2791.160 2291.190 2791.300 ;
        RECT 1797.750 2791.100 1798.070 2791.160 ;
        RECT 2290.870 2791.100 2291.190 2791.160 ;
        RECT 2335.490 2791.300 2335.810 2791.360 ;
        RECT 2442.670 2791.300 2442.990 2791.360 ;
        RECT 2335.490 2791.160 2442.990 2791.300 ;
        RECT 2335.490 2791.100 2335.810 2791.160 ;
        RECT 2442.670 2791.100 2442.990 2791.160 ;
        RECT 2218.190 2790.960 2218.510 2791.020 ;
        RECT 2297.770 2790.960 2298.090 2791.020 ;
        RECT 2218.190 2790.820 2298.090 2790.960 ;
        RECT 2218.190 2790.760 2218.510 2790.820 ;
        RECT 2297.770 2790.760 2298.090 2790.820 ;
        RECT 2328.590 2790.960 2328.910 2791.020 ;
        RECT 2435.770 2790.960 2436.090 2791.020 ;
        RECT 2328.590 2790.820 2436.090 2790.960 ;
        RECT 2328.590 2790.760 2328.910 2790.820 ;
        RECT 2435.770 2790.760 2436.090 2790.820 ;
        RECT 641.310 2790.620 641.630 2790.680 ;
        RECT 979.870 2790.620 980.190 2790.680 ;
        RECT 641.310 2790.480 980.190 2790.620 ;
        RECT 641.310 2790.420 641.630 2790.480 ;
        RECT 979.870 2790.420 980.190 2790.480 ;
        RECT 1024.490 2790.620 1024.810 2790.680 ;
        RECT 1069.570 2790.620 1069.890 2790.680 ;
        RECT 1024.490 2790.480 1069.890 2790.620 ;
        RECT 1024.490 2790.420 1024.810 2790.480 ;
        RECT 1069.570 2790.420 1069.890 2790.480 ;
        RECT 1452.290 2790.620 1452.610 2790.680 ;
        RECT 1656.070 2790.620 1656.390 2790.680 ;
        RECT 1452.290 2790.480 1656.390 2790.620 ;
        RECT 1452.290 2790.420 1452.610 2790.480 ;
        RECT 1656.070 2790.420 1656.390 2790.480 ;
        RECT 1748.990 2790.620 1749.310 2790.680 ;
        RECT 2263.270 2790.620 2263.590 2790.680 ;
        RECT 1748.990 2790.480 2263.590 2790.620 ;
        RECT 1748.990 2790.420 1749.310 2790.480 ;
        RECT 2263.270 2790.420 2263.590 2790.480 ;
        RECT 2273.390 2790.620 2273.710 2790.680 ;
        RECT 2321.230 2790.620 2321.550 2790.680 ;
        RECT 2273.390 2790.480 2321.550 2790.620 ;
        RECT 2273.390 2790.420 2273.710 2790.480 ;
        RECT 2321.230 2790.420 2321.550 2790.480 ;
        RECT 2321.690 2790.620 2322.010 2790.680 ;
        RECT 2428.870 2790.620 2429.190 2790.680 ;
        RECT 2321.690 2790.480 2429.190 2790.620 ;
        RECT 2321.690 2790.420 2322.010 2790.480 ;
        RECT 2428.870 2790.420 2429.190 2790.480 ;
        RECT 403.490 2790.280 403.810 2790.340 ;
        RECT 414.070 2790.280 414.390 2790.340 ;
        RECT 403.490 2790.140 414.390 2790.280 ;
        RECT 403.490 2790.080 403.810 2790.140 ;
        RECT 414.070 2790.080 414.390 2790.140 ;
        RECT 503.770 2790.280 504.090 2790.340 ;
        RECT 509.290 2790.280 509.610 2790.340 ;
        RECT 993.670 2790.280 993.990 2790.340 ;
        RECT 503.770 2790.140 993.990 2790.280 ;
        RECT 503.770 2790.080 504.090 2790.140 ;
        RECT 509.290 2790.080 509.610 2790.140 ;
        RECT 993.670 2790.080 993.990 2790.140 ;
        RECT 1031.390 2790.280 1031.710 2790.340 ;
        RECT 1076.470 2790.280 1076.790 2790.340 ;
        RECT 1031.390 2790.140 1076.790 2790.280 ;
        RECT 1031.390 2790.080 1031.710 2790.140 ;
        RECT 1076.470 2790.080 1076.790 2790.140 ;
        RECT 1610.990 2790.280 1611.310 2790.340 ;
        RECT 1642.270 2790.280 1642.590 2790.340 ;
        RECT 1610.990 2790.140 1642.590 2790.280 ;
        RECT 1610.990 2790.080 1611.310 2790.140 ;
        RECT 1642.270 2790.080 1642.590 2790.140 ;
        RECT 1645.490 2790.280 1645.810 2790.340 ;
        RECT 1686.890 2790.280 1687.210 2790.340 ;
        RECT 1645.490 2790.140 1687.210 2790.280 ;
        RECT 1645.490 2790.080 1645.810 2790.140 ;
        RECT 1686.890 2790.080 1687.210 2790.140 ;
        RECT 1762.790 2790.280 1763.110 2790.340 ;
        RECT 2380.570 2790.280 2380.890 2790.340 ;
        RECT 1762.790 2790.140 2380.890 2790.280 ;
        RECT 1762.790 2790.080 1763.110 2790.140 ;
        RECT 2380.570 2790.080 2380.890 2790.140 ;
        RECT 501.470 2789.940 501.790 2790.000 ;
        RECT 986.770 2789.940 987.090 2790.000 ;
        RECT 501.470 2789.800 987.090 2789.940 ;
        RECT 501.470 2789.740 501.790 2789.800 ;
        RECT 986.770 2789.740 987.090 2789.800 ;
        RECT 1046.110 2789.940 1046.430 2790.000 ;
        RECT 1083.370 2789.940 1083.690 2790.000 ;
        RECT 1046.110 2789.800 1083.690 2789.940 ;
        RECT 1046.110 2789.740 1046.430 2789.800 ;
        RECT 1083.370 2789.740 1083.690 2789.800 ;
        RECT 1638.590 2789.940 1638.910 2790.000 ;
        RECT 1683.210 2789.940 1683.530 2790.000 ;
        RECT 1638.590 2789.800 1683.530 2789.940 ;
        RECT 1638.590 2789.740 1638.910 2789.800 ;
        RECT 1683.210 2789.740 1683.530 2789.800 ;
        RECT 1763.250 2789.940 1763.570 2790.000 ;
        RECT 2387.470 2789.940 2387.790 2790.000 ;
        RECT 1763.250 2789.800 2387.790 2789.940 ;
        RECT 1763.250 2789.740 1763.570 2789.800 ;
        RECT 2387.470 2789.740 2387.790 2789.800 ;
        RECT 358.410 2789.600 358.730 2789.660 ;
        RECT 393.370 2789.600 393.690 2789.660 ;
        RECT 358.410 2789.460 393.690 2789.600 ;
        RECT 358.410 2789.400 358.730 2789.460 ;
        RECT 393.370 2789.400 393.690 2789.460 ;
        RECT 1010.690 2789.600 1011.010 2789.660 ;
        RECT 1055.770 2789.600 1056.090 2789.660 ;
        RECT 1010.690 2789.460 1056.090 2789.600 ;
        RECT 1010.690 2789.400 1011.010 2789.460 ;
        RECT 1055.770 2789.400 1056.090 2789.460 ;
        RECT 1611.450 2789.600 1611.770 2789.660 ;
        RECT 1656.530 2789.600 1656.850 2789.660 ;
        RECT 1611.450 2789.460 1656.850 2789.600 ;
        RECT 1611.450 2789.400 1611.770 2789.460 ;
        RECT 1656.530 2789.400 1656.850 2789.460 ;
        RECT 1763.710 2789.600 1764.030 2789.660 ;
        RECT 2394.370 2789.600 2394.690 2789.660 ;
        RECT 1763.710 2789.460 2394.690 2789.600 ;
        RECT 1763.710 2789.400 1764.030 2789.460 ;
        RECT 2394.370 2789.400 2394.690 2789.460 ;
        RECT 351.510 2789.260 351.830 2789.320 ;
        RECT 386.470 2789.260 386.790 2789.320 ;
        RECT 351.510 2789.120 386.790 2789.260 ;
        RECT 351.510 2789.060 351.830 2789.120 ;
        RECT 386.470 2789.060 386.790 2789.120 ;
        RECT 467.890 2789.260 468.210 2789.320 ;
        RECT 513.430 2789.260 513.750 2789.320 ;
        RECT 1007.470 2789.260 1007.790 2789.320 ;
        RECT 467.890 2789.120 1007.790 2789.260 ;
        RECT 467.890 2789.060 468.210 2789.120 ;
        RECT 513.430 2789.060 513.750 2789.120 ;
        RECT 1007.470 2789.060 1007.790 2789.120 ;
        RECT 1017.590 2789.260 1017.910 2789.320 ;
        RECT 1062.670 2789.260 1062.990 2789.320 ;
        RECT 1017.590 2789.120 1062.990 2789.260 ;
        RECT 1017.590 2789.060 1017.910 2789.120 ;
        RECT 1062.670 2789.060 1062.990 2789.120 ;
        RECT 1514.390 2789.260 1514.710 2789.320 ;
        RECT 1614.670 2789.260 1614.990 2789.320 ;
        RECT 1514.390 2789.120 1614.990 2789.260 ;
        RECT 1514.390 2789.060 1514.710 2789.120 ;
        RECT 1614.670 2789.060 1614.990 2789.120 ;
        RECT 1618.350 2789.260 1618.670 2789.320 ;
        RECT 1663.430 2789.260 1663.750 2789.320 ;
        RECT 1618.350 2789.120 1663.750 2789.260 ;
        RECT 1618.350 2789.060 1618.670 2789.120 ;
        RECT 1663.430 2789.060 1663.750 2789.120 ;
        RECT 1769.690 2789.260 1770.010 2789.320 ;
        RECT 2402.650 2789.260 2402.970 2789.320 ;
        RECT 1769.690 2789.120 2402.970 2789.260 ;
        RECT 1769.690 2789.060 1770.010 2789.120 ;
        RECT 2402.650 2789.060 2402.970 2789.120 ;
        RECT 330.810 2788.920 331.130 2788.980 ;
        RECT 372.670 2788.920 372.990 2788.980 ;
        RECT 330.810 2788.780 372.990 2788.920 ;
        RECT 330.810 2788.720 331.130 2788.780 ;
        RECT 372.670 2788.720 372.990 2788.780 ;
        RECT 530.450 2788.920 530.770 2788.980 ;
        RECT 1028.170 2788.920 1028.490 2788.980 ;
        RECT 530.450 2788.780 1028.490 2788.920 ;
        RECT 530.450 2788.720 530.770 2788.780 ;
        RECT 1028.170 2788.720 1028.490 2788.780 ;
        RECT 1438.950 2788.920 1439.270 2788.980 ;
        RECT 1587.070 2788.920 1587.390 2788.980 ;
        RECT 1438.950 2788.780 1587.390 2788.920 ;
        RECT 1438.950 2788.720 1439.270 2788.780 ;
        RECT 1587.070 2788.720 1587.390 2788.780 ;
        RECT 1624.790 2788.920 1625.110 2788.980 ;
        RECT 1670.330 2788.920 1670.650 2788.980 ;
        RECT 1624.790 2788.780 1670.650 2788.920 ;
        RECT 1624.790 2788.720 1625.110 2788.780 ;
        RECT 1670.330 2788.720 1670.650 2788.780 ;
        RECT 1783.490 2788.920 1783.810 2788.980 ;
        RECT 2415.070 2788.920 2415.390 2788.980 ;
        RECT 1783.490 2788.780 2415.390 2788.920 ;
        RECT 1783.490 2788.720 1783.810 2788.780 ;
        RECT 2415.070 2788.720 2415.390 2788.780 ;
        RECT 337.250 2788.580 337.570 2788.640 ;
        RECT 379.570 2788.580 379.890 2788.640 ;
        RECT 337.250 2788.440 379.890 2788.580 ;
        RECT 337.250 2788.380 337.570 2788.440 ;
        RECT 379.570 2788.380 379.890 2788.440 ;
        RECT 537.350 2788.580 537.670 2788.640 ;
        RECT 1035.070 2788.580 1035.390 2788.640 ;
        RECT 537.350 2788.440 1035.390 2788.580 ;
        RECT 537.350 2788.380 537.670 2788.440 ;
        RECT 1035.070 2788.380 1035.390 2788.440 ;
        RECT 1038.290 2788.580 1038.610 2788.640 ;
        RECT 1083.830 2788.580 1084.150 2788.640 ;
        RECT 1038.290 2788.440 1084.150 2788.580 ;
        RECT 1038.290 2788.380 1038.610 2788.440 ;
        RECT 1083.830 2788.380 1084.150 2788.440 ;
        RECT 1432.050 2788.580 1432.370 2788.640 ;
        RECT 1600.870 2788.580 1601.190 2788.640 ;
        RECT 1432.050 2788.440 1601.190 2788.580 ;
        RECT 1432.050 2788.380 1432.370 2788.440 ;
        RECT 1600.870 2788.380 1601.190 2788.440 ;
        RECT 1631.690 2788.580 1632.010 2788.640 ;
        RECT 1677.230 2788.580 1677.550 2788.640 ;
        RECT 1631.690 2788.440 1677.550 2788.580 ;
        RECT 1631.690 2788.380 1632.010 2788.440 ;
        RECT 1677.230 2788.380 1677.550 2788.440 ;
        RECT 1770.150 2788.580 1770.470 2788.640 ;
        RECT 2408.170 2788.580 2408.490 2788.640 ;
        RECT 1770.150 2788.440 2408.490 2788.580 ;
        RECT 1770.150 2788.380 1770.470 2788.440 ;
        RECT 2408.170 2788.380 2408.490 2788.440 ;
        RECT 317.010 2788.240 317.330 2788.300 ;
        RECT 365.770 2788.240 366.090 2788.300 ;
        RECT 317.010 2788.100 366.090 2788.240 ;
        RECT 317.010 2788.040 317.330 2788.100 ;
        RECT 365.770 2788.040 366.090 2788.100 ;
        RECT 523.550 2788.240 523.870 2788.300 ;
        RECT 1014.370 2788.240 1014.690 2788.300 ;
        RECT 523.550 2788.100 1014.690 2788.240 ;
        RECT 523.550 2788.040 523.870 2788.100 ;
        RECT 1014.370 2788.040 1014.690 2788.100 ;
        RECT 1045.190 2788.240 1045.510 2788.300 ;
        RECT 1090.270 2788.240 1090.590 2788.300 ;
        RECT 1045.190 2788.100 1090.590 2788.240 ;
        RECT 1045.190 2788.040 1045.510 2788.100 ;
        RECT 1090.270 2788.040 1090.590 2788.100 ;
        RECT 1646.410 2788.240 1646.730 2788.300 ;
        RECT 1694.710 2788.240 1695.030 2788.300 ;
        RECT 1646.410 2788.100 1695.030 2788.240 ;
        RECT 1646.410 2788.040 1646.730 2788.100 ;
        RECT 1694.710 2788.040 1695.030 2788.100 ;
        RECT 1790.390 2788.240 1790.710 2788.300 ;
        RECT 2270.170 2788.240 2270.490 2788.300 ;
        RECT 1790.390 2788.100 2270.490 2788.240 ;
        RECT 1790.390 2788.040 1790.710 2788.100 ;
        RECT 2270.170 2788.040 2270.490 2788.100 ;
        RECT 2280.290 2788.240 2280.610 2788.300 ;
        RECT 2325.830 2788.240 2326.150 2788.300 ;
        RECT 2280.290 2788.100 2326.150 2788.240 ;
        RECT 2280.290 2788.040 2280.610 2788.100 ;
        RECT 2325.830 2788.040 2326.150 2788.100 ;
        RECT 2342.850 2788.240 2343.170 2788.300 ;
        RECT 2387.930 2788.240 2388.250 2788.300 ;
        RECT 2342.850 2788.100 2388.250 2788.240 ;
        RECT 2342.850 2788.040 2343.170 2788.100 ;
        RECT 2387.930 2788.040 2388.250 2788.100 ;
        RECT 310.110 2787.900 310.430 2787.960 ;
        RECT 358.870 2787.900 359.190 2787.960 ;
        RECT 310.110 2787.760 359.190 2787.900 ;
        RECT 310.110 2787.700 310.430 2787.760 ;
        RECT 358.870 2787.700 359.190 2787.760 ;
        RECT 372.210 2787.900 372.530 2787.960 ;
        RECT 393.370 2787.900 393.690 2787.960 ;
        RECT 372.210 2787.760 393.690 2787.900 ;
        RECT 372.210 2787.700 372.530 2787.760 ;
        RECT 393.370 2787.700 393.690 2787.760 ;
        RECT 1052.090 2787.900 1052.410 2787.960 ;
        RECT 1100.390 2787.900 1100.710 2787.960 ;
        RECT 1139.030 2787.900 1139.350 2787.960 ;
        RECT 1052.090 2787.760 1139.350 2787.900 ;
        RECT 1052.090 2787.700 1052.410 2787.760 ;
        RECT 1100.390 2787.700 1100.710 2787.760 ;
        RECT 1139.030 2787.700 1139.350 2787.760 ;
        RECT 1652.390 2787.900 1652.710 2787.960 ;
        RECT 1699.310 2787.900 1699.630 2787.960 ;
        RECT 1652.390 2787.760 1699.630 2787.900 ;
        RECT 1652.390 2787.700 1652.710 2787.760 ;
        RECT 1699.310 2787.700 1699.630 2787.760 ;
        RECT 2252.690 2787.900 2253.010 2787.960 ;
        RECT 2256.830 2787.900 2257.150 2787.960 ;
        RECT 2252.690 2787.760 2257.150 2787.900 ;
        RECT 2252.690 2787.700 2253.010 2787.760 ;
        RECT 2256.830 2787.700 2257.150 2787.760 ;
        RECT 2287.190 2787.900 2287.510 2787.960 ;
        RECT 2332.730 2787.900 2333.050 2787.960 ;
        RECT 2373.210 2787.900 2373.530 2787.960 ;
        RECT 2287.190 2787.760 2373.530 2787.900 ;
        RECT 2287.190 2787.700 2287.510 2787.760 ;
        RECT 2332.730 2787.700 2333.050 2787.760 ;
        RECT 2373.210 2787.700 2373.530 2787.760 ;
        RECT 2374.130 2787.900 2374.450 2787.960 ;
        RECT 2415.070 2787.900 2415.390 2787.960 ;
        RECT 2374.130 2787.760 2415.390 2787.900 ;
        RECT 2374.130 2787.700 2374.450 2787.760 ;
        RECT 2415.070 2787.700 2415.390 2787.760 ;
        RECT 283.890 2718.540 284.210 2718.600 ;
        RECT 730.090 2718.540 730.410 2718.600 ;
        RECT 283.890 2718.400 730.410 2718.540 ;
        RECT 283.890 2718.340 284.210 2718.400 ;
        RECT 730.090 2718.340 730.410 2718.400 ;
        RECT 1034.610 2718.540 1034.930 2718.600 ;
        RECT 1103.610 2718.540 1103.930 2718.600 ;
        RECT 1034.610 2718.400 1103.930 2718.540 ;
        RECT 1034.610 2718.340 1034.930 2718.400 ;
        RECT 1103.610 2718.340 1103.930 2718.400 ;
        RECT 1145.010 2718.540 1145.330 2718.600 ;
        RECT 1300.950 2718.540 1301.270 2718.600 ;
        RECT 1145.010 2718.400 1301.270 2718.540 ;
        RECT 1145.010 2718.340 1145.330 2718.400 ;
        RECT 1300.950 2718.340 1301.270 2718.400 ;
        RECT 284.350 2718.200 284.670 2718.260 ;
        RECT 740.670 2718.200 740.990 2718.260 ;
        RECT 284.350 2718.060 740.990 2718.200 ;
        RECT 284.350 2718.000 284.670 2718.060 ;
        RECT 740.670 2718.000 740.990 2718.060 ;
        RECT 1027.710 2718.200 1028.030 2718.260 ;
        RECT 1093.490 2718.200 1093.810 2718.260 ;
        RECT 1027.710 2718.060 1093.810 2718.200 ;
        RECT 1027.710 2718.000 1028.030 2718.060 ;
        RECT 1093.490 2718.000 1093.810 2718.060 ;
        RECT 1138.110 2718.200 1138.430 2718.260 ;
        RECT 1290.370 2718.200 1290.690 2718.260 ;
        RECT 1138.110 2718.060 1290.690 2718.200 ;
        RECT 1138.110 2718.000 1138.430 2718.060 ;
        RECT 1290.370 2718.000 1290.690 2718.060 ;
        RECT 305.050 2717.860 305.370 2717.920 ;
        RECT 310.110 2717.860 310.430 2717.920 ;
        RECT 750.790 2717.860 751.110 2717.920 ;
        RECT 305.050 2717.720 310.430 2717.860 ;
        RECT 305.050 2717.660 305.370 2717.720 ;
        RECT 310.110 2717.660 310.430 2717.720 ;
        RECT 310.660 2717.720 751.110 2717.860 ;
        RECT 284.810 2717.520 285.130 2717.580 ;
        RECT 310.660 2717.520 310.800 2717.720 ;
        RECT 750.790 2717.660 751.110 2717.720 ;
        RECT 823.470 2717.860 823.790 2717.920 ;
        RECT 827.610 2717.860 827.930 2717.920 ;
        RECT 823.470 2717.720 827.930 2717.860 ;
        RECT 823.470 2717.660 823.790 2717.720 ;
        RECT 827.610 2717.660 827.930 2717.720 ;
        RECT 886.030 2717.860 886.350 2717.920 ;
        RECT 889.710 2717.860 890.030 2717.920 ;
        RECT 886.030 2717.720 890.030 2717.860 ;
        RECT 886.030 2717.660 886.350 2717.720 ;
        RECT 889.710 2717.660 890.030 2717.720 ;
        RECT 1041.510 2717.860 1041.830 2717.920 ;
        RECT 1114.190 2717.860 1114.510 2717.920 ;
        RECT 1041.510 2717.720 1114.510 2717.860 ;
        RECT 1041.510 2717.660 1041.830 2717.720 ;
        RECT 1114.190 2717.660 1114.510 2717.720 ;
        RECT 1158.810 2717.860 1159.130 2717.920 ;
        RECT 1321.650 2717.860 1321.970 2717.920 ;
        RECT 1158.810 2717.720 1321.970 2717.860 ;
        RECT 1158.810 2717.660 1159.130 2717.720 ;
        RECT 1321.650 2717.660 1321.970 2717.720 ;
        RECT 761.370 2717.520 761.690 2717.580 ;
        RECT 284.810 2717.380 310.800 2717.520 ;
        RECT 311.120 2717.380 761.690 2717.520 ;
        RECT 284.810 2717.320 285.130 2717.380 ;
        RECT 285.270 2717.180 285.590 2717.240 ;
        RECT 311.120 2717.180 311.260 2717.380 ;
        RECT 761.370 2717.320 761.690 2717.380 ;
        RECT 802.770 2717.520 803.090 2717.580 ;
        RECT 806.910 2717.520 807.230 2717.580 ;
        RECT 802.770 2717.380 807.230 2717.520 ;
        RECT 802.770 2717.320 803.090 2717.380 ;
        RECT 806.910 2717.320 807.230 2717.380 ;
        RECT 968.830 2717.520 969.150 2717.580 ;
        RECT 1045.190 2717.520 1045.510 2717.580 ;
        RECT 968.830 2717.380 1045.510 2717.520 ;
        RECT 968.830 2717.320 969.150 2717.380 ;
        RECT 1045.190 2717.320 1045.510 2717.380 ;
        RECT 1048.410 2717.520 1048.730 2717.580 ;
        RECT 1124.310 2717.520 1124.630 2717.580 ;
        RECT 1048.410 2717.380 1124.630 2717.520 ;
        RECT 1048.410 2717.320 1048.730 2717.380 ;
        RECT 1124.310 2717.320 1124.630 2717.380 ;
        RECT 1151.910 2717.520 1152.230 2717.580 ;
        RECT 1311.070 2717.520 1311.390 2717.580 ;
        RECT 1151.910 2717.380 1311.390 2717.520 ;
        RECT 1151.910 2717.320 1152.230 2717.380 ;
        RECT 1311.070 2717.320 1311.390 2717.380 ;
        RECT 771.950 2717.180 772.270 2717.240 ;
        RECT 285.270 2717.040 311.260 2717.180 ;
        RECT 311.580 2717.040 772.270 2717.180 ;
        RECT 285.270 2716.980 285.590 2717.040 ;
        RECT 285.730 2716.840 286.050 2716.900 ;
        RECT 311.580 2716.840 311.720 2717.040 ;
        RECT 771.950 2716.980 772.270 2717.040 ;
        RECT 979.410 2717.180 979.730 2717.240 ;
        RECT 1052.090 2717.180 1052.410 2717.240 ;
        RECT 979.410 2717.040 1052.410 2717.180 ;
        RECT 979.410 2716.980 979.730 2717.040 ;
        RECT 1052.090 2716.980 1052.410 2717.040 ;
        RECT 1054.850 2717.180 1055.170 2717.240 ;
        RECT 1134.890 2717.180 1135.210 2717.240 ;
        RECT 1054.850 2717.040 1135.210 2717.180 ;
        RECT 1054.850 2716.980 1055.170 2717.040 ;
        RECT 1134.890 2716.980 1135.210 2717.040 ;
        RECT 1165.250 2717.180 1165.570 2717.240 ;
        RECT 1332.230 2717.180 1332.550 2717.240 ;
        RECT 1165.250 2717.040 1332.550 2717.180 ;
        RECT 1165.250 2716.980 1165.570 2717.040 ;
        RECT 1332.230 2716.980 1332.550 2717.040 ;
        RECT 782.070 2716.840 782.390 2716.900 ;
        RECT 285.730 2716.700 311.720 2716.840 ;
        RECT 312.040 2716.700 782.390 2716.840 ;
        RECT 285.730 2716.640 286.050 2716.700 ;
        RECT 286.190 2716.500 286.510 2716.560 ;
        RECT 312.040 2716.500 312.180 2716.700 ;
        RECT 782.070 2716.640 782.390 2716.700 ;
        RECT 948.130 2716.840 948.450 2716.900 ;
        RECT 1038.290 2716.840 1038.610 2716.900 ;
        RECT 948.130 2716.700 1038.610 2716.840 ;
        RECT 948.130 2716.640 948.450 2716.700 ;
        RECT 1038.290 2716.640 1038.610 2716.700 ;
        RECT 1062.210 2716.840 1062.530 2716.900 ;
        RECT 1155.590 2716.840 1155.910 2716.900 ;
        RECT 1062.210 2716.700 1155.910 2716.840 ;
        RECT 1062.210 2716.640 1062.530 2716.700 ;
        RECT 1155.590 2716.640 1155.910 2716.700 ;
        RECT 1165.710 2716.840 1166.030 2716.900 ;
        RECT 1342.350 2716.840 1342.670 2716.900 ;
        RECT 1165.710 2716.700 1342.670 2716.840 ;
        RECT 1165.710 2716.640 1166.030 2716.700 ;
        RECT 1342.350 2716.640 1342.670 2716.700 ;
        RECT 286.190 2716.360 312.180 2716.500 ;
        RECT 325.750 2716.500 326.070 2716.560 ;
        RECT 330.810 2716.500 331.130 2716.560 ;
        RECT 325.750 2716.360 331.130 2716.500 ;
        RECT 286.190 2716.300 286.510 2716.360 ;
        RECT 325.750 2716.300 326.070 2716.360 ;
        RECT 330.810 2716.300 331.130 2716.360 ;
        RECT 367.150 2716.500 367.470 2716.560 ;
        RECT 372.210 2716.500 372.530 2716.560 ;
        RECT 367.150 2716.360 372.530 2716.500 ;
        RECT 367.150 2716.300 367.470 2716.360 ;
        RECT 372.210 2716.300 372.530 2716.360 ;
        RECT 387.850 2716.500 388.170 2716.560 ;
        RECT 396.590 2716.500 396.910 2716.560 ;
        RECT 387.850 2716.360 396.910 2716.500 ;
        RECT 387.850 2716.300 388.170 2716.360 ;
        RECT 396.590 2716.300 396.910 2716.360 ;
        RECT 398.430 2716.500 398.750 2716.560 ;
        RECT 403.490 2716.500 403.810 2716.560 ;
        RECT 398.430 2716.360 403.810 2716.500 ;
        RECT 398.430 2716.300 398.750 2716.360 ;
        RECT 403.490 2716.300 403.810 2716.360 ;
        RECT 403.950 2716.500 404.270 2716.560 ;
        RECT 844.170 2716.500 844.490 2716.560 ;
        RECT 403.950 2716.360 844.490 2716.500 ;
        RECT 403.950 2716.300 404.270 2716.360 ;
        RECT 844.170 2716.300 844.490 2716.360 ;
        RECT 958.710 2716.500 959.030 2716.560 ;
        RECT 1046.110 2716.500 1046.430 2716.560 ;
        RECT 958.710 2716.360 1046.430 2716.500 ;
        RECT 958.710 2716.300 959.030 2716.360 ;
        RECT 1046.110 2716.300 1046.430 2716.360 ;
        RECT 1055.310 2716.500 1055.630 2716.560 ;
        RECT 1145.470 2716.500 1145.790 2716.560 ;
        RECT 1055.310 2716.360 1145.790 2716.500 ;
        RECT 1055.310 2716.300 1055.630 2716.360 ;
        RECT 1145.470 2716.300 1145.790 2716.360 ;
        RECT 1172.610 2716.500 1172.930 2716.560 ;
        RECT 1352.930 2716.500 1353.250 2716.560 ;
        RECT 1172.610 2716.360 1353.250 2716.500 ;
        RECT 1172.610 2716.300 1172.930 2716.360 ;
        RECT 1352.930 2716.300 1353.250 2716.360 ;
        RECT 350.590 2716.160 350.910 2716.220 ;
        RECT 854.750 2716.160 855.070 2716.220 ;
        RECT 350.590 2716.020 855.070 2716.160 ;
        RECT 350.590 2715.960 350.910 2716.020 ;
        RECT 854.750 2715.960 855.070 2716.020 ;
        RECT 937.550 2716.160 937.870 2716.220 ;
        RECT 1031.390 2716.160 1031.710 2716.220 ;
        RECT 937.550 2716.020 1031.710 2716.160 ;
        RECT 937.550 2715.960 937.870 2716.020 ;
        RECT 1031.390 2715.960 1031.710 2716.020 ;
        RECT 1069.110 2716.160 1069.430 2716.220 ;
        RECT 1166.170 2716.160 1166.490 2716.220 ;
        RECT 1069.110 2716.020 1166.490 2716.160 ;
        RECT 1069.110 2715.960 1069.430 2716.020 ;
        RECT 1166.170 2715.960 1166.490 2716.020 ;
        RECT 1179.510 2716.160 1179.830 2716.220 ;
        RECT 1363.050 2716.160 1363.370 2716.220 ;
        RECT 1179.510 2716.020 1363.370 2716.160 ;
        RECT 1179.510 2715.960 1179.830 2716.020 ;
        RECT 1363.050 2715.960 1363.370 2716.020 ;
        RECT 351.050 2715.820 351.370 2715.880 ;
        RECT 865.330 2715.820 865.650 2715.880 ;
        RECT 351.050 2715.680 865.650 2715.820 ;
        RECT 351.050 2715.620 351.370 2715.680 ;
        RECT 865.330 2715.620 865.650 2715.680 ;
        RECT 927.430 2715.820 927.750 2715.880 ;
        RECT 1024.490 2715.820 1024.810 2715.880 ;
        RECT 927.430 2715.680 1024.810 2715.820 ;
        RECT 927.430 2715.620 927.750 2715.680 ;
        RECT 1024.490 2715.620 1024.810 2715.680 ;
        RECT 1082.910 2715.820 1083.230 2715.880 ;
        RECT 1186.870 2715.820 1187.190 2715.880 ;
        RECT 1082.910 2715.680 1187.190 2715.820 ;
        RECT 1082.910 2715.620 1083.230 2715.680 ;
        RECT 1186.870 2715.620 1187.190 2715.680 ;
        RECT 1193.310 2715.820 1193.630 2715.880 ;
        RECT 1383.750 2715.820 1384.070 2715.880 ;
        RECT 1193.310 2715.680 1384.070 2715.820 ;
        RECT 1193.310 2715.620 1193.630 2715.680 ;
        RECT 1383.750 2715.620 1384.070 2715.680 ;
        RECT 357.950 2715.480 358.270 2715.540 ;
        RECT 875.450 2715.480 875.770 2715.540 ;
        RECT 357.950 2715.340 875.770 2715.480 ;
        RECT 357.950 2715.280 358.270 2715.340 ;
        RECT 875.450 2715.280 875.770 2715.340 ;
        RECT 916.850 2715.480 917.170 2715.540 ;
        RECT 1017.590 2715.480 1017.910 2715.540 ;
        RECT 916.850 2715.340 1017.910 2715.480 ;
        RECT 916.850 2715.280 917.170 2715.340 ;
        RECT 1017.590 2715.280 1017.910 2715.340 ;
        RECT 1076.010 2715.480 1076.330 2715.540 ;
        RECT 1176.290 2715.480 1176.610 2715.540 ;
        RECT 1076.010 2715.340 1176.610 2715.480 ;
        RECT 1076.010 2715.280 1076.330 2715.340 ;
        RECT 1176.290 2715.280 1176.610 2715.340 ;
        RECT 1186.410 2715.480 1186.730 2715.540 ;
        RECT 1373.630 2715.480 1373.950 2715.540 ;
        RECT 1186.410 2715.340 1373.950 2715.480 ;
        RECT 1186.410 2715.280 1186.730 2715.340 ;
        RECT 1373.630 2715.280 1373.950 2715.340 ;
        RECT 283.430 2715.140 283.750 2715.200 ;
        RECT 896.150 2715.140 896.470 2715.200 ;
        RECT 283.430 2715.000 896.470 2715.140 ;
        RECT 283.430 2714.940 283.750 2715.000 ;
        RECT 896.150 2714.940 896.470 2715.000 ;
        RECT 906.730 2715.140 907.050 2715.200 ;
        RECT 1010.690 2715.140 1011.010 2715.200 ;
        RECT 906.730 2715.000 1011.010 2715.140 ;
        RECT 906.730 2714.940 907.050 2715.000 ;
        RECT 1010.690 2714.940 1011.010 2715.000 ;
        RECT 1013.910 2715.140 1014.230 2715.200 ;
        RECT 1072.790 2715.140 1073.110 2715.200 ;
        RECT 1013.910 2715.000 1073.110 2715.140 ;
        RECT 1013.910 2714.940 1014.230 2715.000 ;
        RECT 1072.790 2714.940 1073.110 2715.000 ;
        RECT 1089.810 2715.140 1090.130 2715.200 ;
        RECT 1196.990 2715.140 1197.310 2715.200 ;
        RECT 1089.810 2715.000 1197.310 2715.140 ;
        RECT 1089.810 2714.940 1090.130 2715.000 ;
        RECT 1196.990 2714.940 1197.310 2715.000 ;
        RECT 1200.210 2715.140 1200.530 2715.200 ;
        RECT 1394.330 2715.140 1394.650 2715.200 ;
        RECT 1200.210 2715.000 1394.650 2715.140 ;
        RECT 1200.210 2714.940 1200.530 2715.000 ;
        RECT 1394.330 2714.940 1394.650 2715.000 ;
        RECT 337.710 2714.800 338.030 2714.860 ;
        RECT 719.970 2714.800 720.290 2714.860 ;
        RECT 337.710 2714.660 720.290 2714.800 ;
        RECT 337.710 2714.600 338.030 2714.660 ;
        RECT 719.970 2714.600 720.290 2714.660 ;
        RECT 1020.810 2714.800 1021.130 2714.860 ;
        RECT 1082.910 2714.800 1083.230 2714.860 ;
        RECT 1020.810 2714.660 1083.230 2714.800 ;
        RECT 1020.810 2714.600 1021.130 2714.660 ;
        RECT 1082.910 2714.600 1083.230 2714.660 ;
        RECT 1131.210 2714.800 1131.530 2714.860 ;
        RECT 1280.250 2714.800 1280.570 2714.860 ;
        RECT 1131.210 2714.660 1280.570 2714.800 ;
        RECT 1131.210 2714.600 1131.530 2714.660 ;
        RECT 1280.250 2714.600 1280.570 2714.660 ;
        RECT 344.610 2714.460 344.930 2714.520 ;
        RECT 403.950 2714.460 404.270 2714.520 ;
        RECT 344.610 2714.320 404.270 2714.460 ;
        RECT 344.610 2714.260 344.930 2714.320 ;
        RECT 403.950 2714.260 404.270 2714.320 ;
        RECT 455.010 2714.460 455.330 2714.520 ;
        RECT 460.530 2714.460 460.850 2714.520 ;
        RECT 455.010 2714.320 460.850 2714.460 ;
        RECT 455.010 2714.260 455.330 2714.320 ;
        RECT 460.530 2714.260 460.850 2714.320 ;
        RECT 461.910 2714.460 462.230 2714.520 ;
        RECT 470.650 2714.460 470.970 2714.520 ;
        RECT 461.910 2714.320 470.970 2714.460 ;
        RECT 461.910 2714.260 462.230 2714.320 ;
        RECT 470.650 2714.260 470.970 2714.320 ;
        RECT 503.310 2714.460 503.630 2714.520 ;
        RECT 543.330 2714.460 543.650 2714.520 ;
        RECT 503.310 2714.320 543.650 2714.460 ;
        RECT 503.310 2714.260 503.630 2714.320 ;
        RECT 543.330 2714.260 543.650 2714.320 ;
        RECT 544.710 2714.460 545.030 2714.520 ;
        RECT 616.010 2714.460 616.330 2714.520 ;
        RECT 544.710 2714.320 616.330 2714.460 ;
        RECT 544.710 2714.260 545.030 2714.320 ;
        RECT 616.010 2714.260 616.330 2714.320 ;
        RECT 636.710 2714.460 637.030 2714.520 ;
        RECT 641.310 2714.460 641.630 2714.520 ;
        RECT 636.710 2714.320 641.630 2714.460 ;
        RECT 636.710 2714.260 637.030 2714.320 ;
        RECT 641.310 2714.260 641.630 2714.320 ;
        RECT 647.290 2714.460 647.610 2714.520 ;
        RECT 942.150 2714.460 942.470 2714.520 ;
        RECT 647.290 2714.320 942.470 2714.460 ;
        RECT 647.290 2714.260 647.610 2714.320 ;
        RECT 942.150 2714.260 942.470 2714.320 ;
        RECT 1130.750 2714.460 1131.070 2714.520 ;
        RECT 1269.670 2714.460 1269.990 2714.520 ;
        RECT 1130.750 2714.320 1269.990 2714.460 ;
        RECT 1130.750 2714.260 1131.070 2714.320 ;
        RECT 1269.670 2714.260 1269.990 2714.320 ;
        RECT 468.350 2714.120 468.670 2714.180 ;
        RECT 481.230 2714.120 481.550 2714.180 ;
        RECT 468.350 2713.980 481.550 2714.120 ;
        RECT 468.350 2713.920 468.670 2713.980 ;
        RECT 481.230 2713.920 481.550 2713.980 ;
        RECT 496.410 2714.120 496.730 2714.180 ;
        RECT 533.210 2714.120 533.530 2714.180 ;
        RECT 496.410 2713.980 533.530 2714.120 ;
        RECT 496.410 2713.920 496.730 2713.980 ;
        RECT 533.210 2713.920 533.530 2713.980 ;
        RECT 551.610 2714.120 551.930 2714.180 ;
        RECT 626.590 2714.120 626.910 2714.180 ;
        RECT 551.610 2713.980 626.910 2714.120 ;
        RECT 551.610 2713.920 551.930 2713.980 ;
        RECT 626.590 2713.920 626.910 2713.980 ;
        RECT 657.410 2714.120 657.730 2714.180 ;
        RECT 941.690 2714.120 942.010 2714.180 ;
        RECT 657.410 2713.980 942.010 2714.120 ;
        RECT 657.410 2713.920 657.730 2713.980 ;
        RECT 941.690 2713.920 942.010 2713.980 ;
        RECT 1117.410 2714.120 1117.730 2714.180 ;
        RECT 1248.970 2714.120 1249.290 2714.180 ;
        RECT 1117.410 2713.980 1249.290 2714.120 ;
        RECT 1117.410 2713.920 1117.730 2713.980 ;
        RECT 1248.970 2713.920 1249.290 2713.980 ;
        RECT 468.810 2713.780 469.130 2713.840 ;
        RECT 491.810 2713.780 492.130 2713.840 ;
        RECT 468.810 2713.640 492.130 2713.780 ;
        RECT 468.810 2713.580 469.130 2713.640 ;
        RECT 491.810 2713.580 492.130 2713.640 ;
        RECT 537.810 2713.780 538.130 2713.840 ;
        RECT 605.890 2713.780 606.210 2713.840 ;
        RECT 537.810 2713.640 606.210 2713.780 ;
        RECT 537.810 2713.580 538.130 2713.640 ;
        RECT 605.890 2713.580 606.210 2713.640 ;
        RECT 699.270 2713.780 699.590 2713.840 ;
        RECT 703.410 2713.780 703.730 2713.840 ;
        RECT 699.270 2713.640 703.730 2713.780 ;
        RECT 699.270 2713.580 699.590 2713.640 ;
        RECT 703.410 2713.580 703.730 2713.640 ;
        RECT 703.870 2713.780 704.190 2713.840 ;
        RECT 796.790 2713.780 797.110 2713.840 ;
        RECT 703.870 2713.640 797.110 2713.780 ;
        RECT 703.870 2713.580 704.190 2713.640 ;
        RECT 796.790 2713.580 797.110 2713.640 ;
        RECT 1123.390 2713.780 1123.710 2713.840 ;
        RECT 1259.550 2713.780 1259.870 2713.840 ;
        RECT 1123.390 2713.640 1259.870 2713.780 ;
        RECT 1123.390 2713.580 1123.710 2713.640 ;
        RECT 1259.550 2713.580 1259.870 2713.640 ;
        RECT 346.450 2713.440 346.770 2713.500 ;
        RECT 351.510 2713.440 351.830 2713.500 ;
        RECT 346.450 2713.300 351.830 2713.440 ;
        RECT 346.450 2713.240 346.770 2713.300 ;
        RECT 351.510 2713.240 351.830 2713.300 ;
        RECT 482.610 2713.440 482.930 2713.500 ;
        RECT 512.510 2713.440 512.830 2713.500 ;
        RECT 522.630 2713.440 522.950 2713.500 ;
        RECT 482.610 2713.300 512.830 2713.440 ;
        RECT 482.610 2713.240 482.930 2713.300 ;
        RECT 512.510 2713.240 512.830 2713.300 ;
        RECT 513.060 2713.300 522.950 2713.440 ;
        RECT 419.130 2713.100 419.450 2713.160 ;
        RECT 428.330 2713.100 428.650 2713.160 ;
        RECT 419.130 2712.960 428.650 2713.100 ;
        RECT 419.130 2712.900 419.450 2712.960 ;
        RECT 428.330 2712.900 428.650 2712.960 ;
        RECT 489.510 2713.100 489.830 2713.160 ;
        RECT 513.060 2713.100 513.200 2713.300 ;
        RECT 522.630 2713.240 522.950 2713.300 ;
        RECT 530.910 2713.440 531.230 2713.500 ;
        RECT 595.310 2713.440 595.630 2713.500 ;
        RECT 530.910 2713.300 595.630 2713.440 ;
        RECT 530.910 2713.240 531.230 2713.300 ;
        RECT 595.310 2713.240 595.630 2713.300 ;
        RECT 678.570 2713.440 678.890 2713.500 ;
        RECT 803.690 2713.440 804.010 2713.500 ;
        RECT 678.570 2713.300 804.010 2713.440 ;
        RECT 678.570 2713.240 678.890 2713.300 ;
        RECT 803.690 2713.240 804.010 2713.300 ;
        RECT 1102.690 2713.440 1103.010 2713.500 ;
        RECT 1228.270 2713.440 1228.590 2713.500 ;
        RECT 1102.690 2713.300 1228.590 2713.440 ;
        RECT 1102.690 2713.240 1103.010 2713.300 ;
        RECT 1228.270 2713.240 1228.590 2713.300 ;
        RECT 489.510 2712.960 513.200 2713.100 ;
        RECT 517.110 2713.100 517.430 2713.160 ;
        RECT 574.610 2713.100 574.930 2713.160 ;
        RECT 517.110 2712.960 574.930 2713.100 ;
        RECT 489.510 2712.900 489.830 2712.960 ;
        RECT 517.110 2712.900 517.430 2712.960 ;
        RECT 574.610 2712.900 574.930 2712.960 ;
        RECT 1110.510 2713.100 1110.830 2713.160 ;
        RECT 1238.850 2713.100 1239.170 2713.160 ;
        RECT 1110.510 2712.960 1239.170 2713.100 ;
        RECT 1110.510 2712.900 1110.830 2712.960 ;
        RECT 1238.850 2712.900 1239.170 2712.960 ;
        RECT 408.550 2712.760 408.870 2712.820 ;
        RECT 420.970 2712.760 421.290 2712.820 ;
        RECT 408.550 2712.620 421.290 2712.760 ;
        RECT 408.550 2712.560 408.870 2712.620 ;
        RECT 420.970 2712.560 421.290 2712.620 ;
        RECT 524.010 2712.760 524.330 2712.820 ;
        RECT 585.190 2712.760 585.510 2712.820 ;
        RECT 524.010 2712.620 585.510 2712.760 ;
        RECT 524.010 2712.560 524.330 2712.620 ;
        RECT 585.190 2712.560 585.510 2712.620 ;
        RECT 667.990 2712.760 668.310 2712.820 ;
        RECT 703.870 2712.760 704.190 2712.820 ;
        RECT 667.990 2712.620 704.190 2712.760 ;
        RECT 667.990 2712.560 668.310 2712.620 ;
        RECT 703.870 2712.560 704.190 2712.620 ;
        RECT 1089.350 2712.760 1089.670 2712.820 ;
        RECT 1207.570 2712.760 1207.890 2712.820 ;
        RECT 1089.350 2712.620 1207.890 2712.760 ;
        RECT 1089.350 2712.560 1089.670 2712.620 ;
        RECT 1207.570 2712.560 1207.890 2712.620 ;
        RECT 475.710 2712.420 476.030 2712.480 ;
        RECT 501.930 2712.420 502.250 2712.480 ;
        RECT 475.710 2712.280 502.250 2712.420 ;
        RECT 475.710 2712.220 476.030 2712.280 ;
        RECT 501.930 2712.220 502.250 2712.280 ;
        RECT 509.750 2712.420 510.070 2712.480 ;
        RECT 564.030 2712.420 564.350 2712.480 ;
        RECT 509.750 2712.280 564.350 2712.420 ;
        RECT 509.750 2712.220 510.070 2712.280 ;
        RECT 564.030 2712.220 564.350 2712.280 ;
        RECT 1096.710 2712.420 1097.030 2712.480 ;
        RECT 1217.690 2712.420 1218.010 2712.480 ;
        RECT 1096.710 2712.280 1218.010 2712.420 ;
        RECT 1096.710 2712.220 1097.030 2712.280 ;
        RECT 1217.690 2712.220 1218.010 2712.280 ;
        RECT 510.210 2712.080 510.530 2712.140 ;
        RECT 553.910 2712.080 554.230 2712.140 ;
        RECT 510.210 2711.940 554.230 2712.080 ;
        RECT 510.210 2711.880 510.530 2711.940 ;
        RECT 553.910 2711.880 554.230 2711.940 ;
        RECT 1055.770 2704.940 1056.090 2705.000 ;
        RECT 1057.150 2704.940 1057.470 2705.000 ;
        RECT 1055.770 2704.800 1057.470 2704.940 ;
        RECT 1055.770 2704.740 1056.090 2704.800 ;
        RECT 1057.150 2704.740 1057.470 2704.800 ;
      LAYER met1 ;
        RECT 305.130 1504.460 1394.730 2689.280 ;
      LAYER met1 ;
        RECT 1414.110 2683.860 1414.430 2683.920 ;
        RECT 2335.490 2683.860 2335.810 2683.920 ;
        RECT 1414.110 2683.720 2335.810 2683.860 ;
        RECT 1414.110 2683.660 1414.430 2683.720 ;
        RECT 2335.490 2683.660 2335.810 2683.720 ;
        RECT 1414.110 2677.060 1414.430 2677.120 ;
        RECT 2328.590 2677.060 2328.910 2677.120 ;
        RECT 1414.110 2676.920 2328.910 2677.060 ;
        RECT 1414.110 2676.860 1414.430 2676.920 ;
        RECT 2328.590 2676.860 2328.910 2676.920 ;
        RECT 1414.110 2663.460 1414.430 2663.520 ;
        RECT 2321.690 2663.460 2322.010 2663.520 ;
        RECT 1414.110 2663.320 2322.010 2663.460 ;
        RECT 1414.110 2663.260 1414.430 2663.320 ;
        RECT 2321.690 2663.260 2322.010 2663.320 ;
        RECT 1414.110 2656.320 1414.430 2656.380 ;
        RECT 1783.950 2656.320 1784.270 2656.380 ;
        RECT 1414.110 2656.180 1784.270 2656.320 ;
        RECT 1414.110 2656.120 1414.430 2656.180 ;
        RECT 1783.950 2656.120 1784.270 2656.180 ;
        RECT 1414.110 2642.720 1414.430 2642.780 ;
        RECT 1783.490 2642.720 1783.810 2642.780 ;
        RECT 1414.110 2642.580 1783.810 2642.720 ;
        RECT 1414.110 2642.520 1414.430 2642.580 ;
        RECT 1783.490 2642.520 1783.810 2642.580 ;
        RECT 1414.110 2628.780 1414.430 2628.840 ;
        RECT 1776.590 2628.780 1776.910 2628.840 ;
        RECT 1414.110 2628.640 1776.910 2628.780 ;
        RECT 1414.110 2628.580 1414.430 2628.640 ;
        RECT 1776.590 2628.580 1776.910 2628.640 ;
        RECT 1414.110 2621.980 1414.430 2622.040 ;
        RECT 1770.150 2621.980 1770.470 2622.040 ;
        RECT 1414.110 2621.840 1770.470 2621.980 ;
        RECT 1414.110 2621.780 1414.430 2621.840 ;
        RECT 1770.150 2621.780 1770.470 2621.840 ;
        RECT 1414.110 2608.040 1414.430 2608.100 ;
        RECT 1769.690 2608.040 1770.010 2608.100 ;
        RECT 1414.110 2607.900 1770.010 2608.040 ;
        RECT 1414.110 2607.840 1414.430 2607.900 ;
        RECT 1769.690 2607.840 1770.010 2607.900 ;
        RECT 1414.110 2601.240 1414.430 2601.300 ;
        RECT 1763.710 2601.240 1764.030 2601.300 ;
        RECT 1414.110 2601.100 1764.030 2601.240 ;
        RECT 1414.110 2601.040 1414.430 2601.100 ;
        RECT 1763.710 2601.040 1764.030 2601.100 ;
        RECT 1409.510 2587.300 1409.830 2587.360 ;
        RECT 1763.250 2587.300 1763.570 2587.360 ;
        RECT 1409.510 2587.160 1763.570 2587.300 ;
        RECT 1409.510 2587.100 1409.830 2587.160 ;
        RECT 1763.250 2587.100 1763.570 2587.160 ;
        RECT 1414.110 2573.700 1414.430 2573.760 ;
        RECT 1762.790 2573.700 1763.110 2573.760 ;
        RECT 1414.110 2573.560 1763.110 2573.700 ;
        RECT 1414.110 2573.500 1414.430 2573.560 ;
        RECT 1762.790 2573.500 1763.110 2573.560 ;
        RECT 1410.430 2566.560 1410.750 2566.620 ;
        RECT 2381.030 2566.560 2381.350 2566.620 ;
        RECT 1410.430 2566.420 2381.350 2566.560 ;
        RECT 1410.430 2566.360 1410.750 2566.420 ;
        RECT 2381.030 2566.360 2381.350 2566.420 ;
        RECT 1414.110 2552.960 1414.430 2553.020 ;
        RECT 2373.670 2552.960 2373.990 2553.020 ;
        RECT 1414.110 2552.820 2373.990 2552.960 ;
        RECT 1414.110 2552.760 1414.430 2552.820 ;
        RECT 2373.670 2552.760 2373.990 2552.820 ;
        RECT 1411.350 2546.160 1411.670 2546.220 ;
        RECT 2366.770 2546.160 2367.090 2546.220 ;
        RECT 1411.350 2546.020 2367.090 2546.160 ;
        RECT 1411.350 2545.960 1411.670 2546.020 ;
        RECT 2366.770 2545.960 2367.090 2546.020 ;
        RECT 1409.510 2532.220 1409.830 2532.280 ;
        RECT 2359.870 2532.220 2360.190 2532.280 ;
        RECT 1409.510 2532.080 2360.190 2532.220 ;
        RECT 1409.510 2532.020 1409.830 2532.080 ;
        RECT 2359.870 2532.020 2360.190 2532.080 ;
        RECT 1414.110 2518.280 1414.430 2518.340 ;
        RECT 2352.970 2518.280 2353.290 2518.340 ;
        RECT 1414.110 2518.140 2353.290 2518.280 ;
        RECT 1414.110 2518.080 1414.430 2518.140 ;
        RECT 2352.970 2518.080 2353.290 2518.140 ;
        RECT 1410.430 2511.480 1410.750 2511.540 ;
        RECT 2346.070 2511.480 2346.390 2511.540 ;
        RECT 1410.430 2511.340 2346.390 2511.480 ;
        RECT 1410.430 2511.280 1410.750 2511.340 ;
        RECT 2346.070 2511.280 2346.390 2511.340 ;
        RECT 1414.110 2497.540 1414.430 2497.600 ;
        RECT 2339.630 2497.540 2339.950 2497.600 ;
        RECT 1414.110 2497.400 2339.950 2497.540 ;
        RECT 1414.110 2497.340 1414.430 2497.400 ;
        RECT 2339.630 2497.340 2339.950 2497.400 ;
        RECT 1411.350 2490.740 1411.670 2490.800 ;
        RECT 2339.170 2490.740 2339.490 2490.800 ;
        RECT 1411.350 2490.600 2339.490 2490.740 ;
        RECT 1411.350 2490.540 1411.670 2490.600 ;
        RECT 2339.170 2490.540 2339.490 2490.600 ;
        RECT 1409.510 2477.140 1409.830 2477.200 ;
        RECT 2332.270 2477.140 2332.590 2477.200 ;
        RECT 1409.510 2477.000 2332.590 2477.140 ;
        RECT 1409.510 2476.940 1409.830 2477.000 ;
        RECT 2332.270 2476.940 2332.590 2477.000 ;
        RECT 1412.270 2470.000 1412.590 2470.060 ;
        RECT 2325.370 2470.000 2325.690 2470.060 ;
        RECT 1412.270 2469.860 2325.690 2470.000 ;
        RECT 1412.270 2469.800 1412.590 2469.860 ;
        RECT 2325.370 2469.800 2325.690 2469.860 ;
        RECT 1410.430 2456.400 1410.750 2456.460 ;
        RECT 2318.470 2456.400 2318.790 2456.460 ;
        RECT 1410.430 2456.260 2318.790 2456.400 ;
        RECT 1410.430 2456.200 1410.750 2456.260 ;
        RECT 2318.470 2456.200 2318.790 2456.260 ;
        RECT 1414.110 2442.460 1414.430 2442.520 ;
        RECT 2311.570 2442.460 2311.890 2442.520 ;
        RECT 1414.110 2442.320 2311.890 2442.460 ;
        RECT 1414.110 2442.260 1414.430 2442.320 ;
        RECT 2311.570 2442.260 2311.890 2442.320 ;
        RECT 1414.110 2435.660 1414.430 2435.720 ;
        RECT 2305.130 2435.660 2305.450 2435.720 ;
        RECT 1414.110 2435.520 2305.450 2435.660 ;
        RECT 1414.110 2435.460 1414.430 2435.520 ;
        RECT 2305.130 2435.460 2305.450 2435.520 ;
        RECT 1414.110 2421.720 1414.430 2421.780 ;
        RECT 2304.670 2421.720 2304.990 2421.780 ;
        RECT 1414.110 2421.580 2304.990 2421.720 ;
        RECT 1414.110 2421.520 1414.430 2421.580 ;
        RECT 2304.670 2421.520 2304.990 2421.580 ;
        RECT 1412.270 2414.920 1412.590 2414.980 ;
        RECT 2218.190 2414.920 2218.510 2414.980 ;
        RECT 1412.270 2414.780 2218.510 2414.920 ;
        RECT 1412.270 2414.720 1412.590 2414.780 ;
        RECT 2218.190 2414.720 2218.510 2414.780 ;
        RECT 1410.430 2400.980 1410.750 2401.040 ;
        RECT 1797.750 2400.980 1798.070 2401.040 ;
        RECT 1410.430 2400.840 1798.070 2400.980 ;
        RECT 1410.430 2400.780 1410.750 2400.840 ;
        RECT 1797.750 2400.780 1798.070 2400.840 ;
        RECT 1414.110 2387.380 1414.430 2387.440 ;
        RECT 1797.290 2387.380 1797.610 2387.440 ;
        RECT 1414.110 2387.240 1797.610 2387.380 ;
        RECT 1414.110 2387.180 1414.430 2387.240 ;
        RECT 1797.290 2387.180 1797.610 2387.240 ;
        RECT 1412.730 2380.240 1413.050 2380.300 ;
        RECT 1790.850 2380.240 1791.170 2380.300 ;
        RECT 1412.730 2380.100 1791.170 2380.240 ;
        RECT 1412.730 2380.040 1413.050 2380.100 ;
        RECT 1790.850 2380.040 1791.170 2380.100 ;
        RECT 1410.430 2366.640 1410.750 2366.700 ;
        RECT 1790.390 2366.640 1790.710 2366.700 ;
        RECT 1410.430 2366.500 1790.710 2366.640 ;
        RECT 1410.430 2366.440 1410.750 2366.500 ;
        RECT 1790.390 2366.440 1790.710 2366.500 ;
        RECT 1412.270 2359.840 1412.590 2359.900 ;
        RECT 1748.990 2359.840 1749.310 2359.900 ;
        RECT 1412.270 2359.700 1749.310 2359.840 ;
        RECT 1412.270 2359.640 1412.590 2359.700 ;
        RECT 1748.990 2359.640 1749.310 2359.700 ;
        RECT 1410.430 2345.900 1410.750 2345.960 ;
        RECT 2263.730 2345.900 2264.050 2345.960 ;
        RECT 1410.430 2345.760 2264.050 2345.900 ;
        RECT 1410.430 2345.700 1410.750 2345.760 ;
        RECT 2263.730 2345.700 2264.050 2345.760 ;
        RECT 1414.110 2331.960 1414.430 2332.020 ;
        RECT 1652.390 2331.960 1652.710 2332.020 ;
        RECT 1414.110 2331.820 1652.710 2331.960 ;
        RECT 1414.110 2331.760 1414.430 2331.820 ;
        RECT 1652.390 2331.760 1652.710 2331.820 ;
        RECT 1411.350 2325.160 1411.670 2325.220 ;
        RECT 1646.410 2325.160 1646.730 2325.220 ;
        RECT 1411.350 2325.020 1646.730 2325.160 ;
        RECT 1411.350 2324.960 1411.670 2325.020 ;
        RECT 1646.410 2324.960 1646.730 2325.020 ;
        RECT 1414.110 2311.560 1414.430 2311.620 ;
        RECT 1645.490 2311.560 1645.810 2311.620 ;
        RECT 1414.110 2311.420 1645.810 2311.560 ;
        RECT 1414.110 2311.360 1414.430 2311.420 ;
        RECT 1645.490 2311.360 1645.810 2311.420 ;
        RECT 1412.270 2304.420 1412.590 2304.480 ;
        RECT 1638.590 2304.420 1638.910 2304.480 ;
        RECT 1412.270 2304.280 1638.910 2304.420 ;
        RECT 1412.270 2304.220 1412.590 2304.280 ;
        RECT 1638.590 2304.220 1638.910 2304.280 ;
        RECT 1410.430 2290.820 1410.750 2290.880 ;
        RECT 1631.690 2290.820 1632.010 2290.880 ;
        RECT 1410.430 2290.680 1632.010 2290.820 ;
        RECT 1410.430 2290.620 1410.750 2290.680 ;
        RECT 1631.690 2290.620 1632.010 2290.680 ;
        RECT 1414.110 2276.880 1414.430 2276.940 ;
        RECT 1624.790 2276.880 1625.110 2276.940 ;
        RECT 1414.110 2276.740 1625.110 2276.880 ;
        RECT 1414.110 2276.680 1414.430 2276.740 ;
        RECT 1624.790 2276.680 1625.110 2276.740 ;
        RECT 1414.110 2270.080 1414.430 2270.140 ;
        RECT 1618.350 2270.080 1618.670 2270.140 ;
        RECT 1414.110 2269.940 1618.670 2270.080 ;
        RECT 1414.110 2269.880 1414.430 2269.940 ;
        RECT 1618.350 2269.880 1618.670 2269.940 ;
        RECT 1414.110 2256.140 1414.430 2256.200 ;
        RECT 1611.450 2256.140 1611.770 2256.200 ;
        RECT 1414.110 2256.000 1611.770 2256.140 ;
        RECT 1414.110 2255.940 1414.430 2256.000 ;
        RECT 1611.450 2255.940 1611.770 2256.000 ;
        RECT 1412.270 2249.340 1412.590 2249.400 ;
        RECT 2301.910 2249.340 2302.230 2249.400 ;
        RECT 1412.270 2249.200 2302.230 2249.340 ;
        RECT 1412.270 2249.140 1412.590 2249.200 ;
        RECT 2301.910 2249.140 2302.230 2249.200 ;
        RECT 1414.110 2235.400 1414.430 2235.460 ;
        RECT 2300.990 2235.400 2301.310 2235.460 ;
        RECT 1414.110 2235.260 2301.310 2235.400 ;
        RECT 1414.110 2235.200 1414.430 2235.260 ;
        RECT 2300.990 2235.200 2301.310 2235.260 ;
        RECT 1414.110 2221.800 1414.430 2221.860 ;
        RECT 2294.090 2221.800 2294.410 2221.860 ;
        RECT 1414.110 2221.660 2294.410 2221.800 ;
        RECT 1414.110 2221.600 1414.430 2221.660 ;
        RECT 2294.090 2221.600 2294.410 2221.660 ;
        RECT 1414.110 2214.660 1414.430 2214.720 ;
        RECT 2287.190 2214.660 2287.510 2214.720 ;
        RECT 1414.110 2214.520 2287.510 2214.660 ;
        RECT 1414.110 2214.460 1414.430 2214.520 ;
        RECT 2287.190 2214.460 2287.510 2214.520 ;
        RECT 1414.110 2201.060 1414.430 2201.120 ;
        RECT 2280.290 2201.060 2280.610 2201.120 ;
        RECT 1414.110 2200.920 2280.610 2201.060 ;
        RECT 1414.110 2200.860 1414.430 2200.920 ;
        RECT 2280.290 2200.860 2280.610 2200.920 ;
        RECT 1412.270 2194.260 1412.590 2194.320 ;
        RECT 2273.390 2194.260 2273.710 2194.320 ;
        RECT 1412.270 2194.120 2273.710 2194.260 ;
        RECT 1412.270 2194.060 1412.590 2194.120 ;
        RECT 2273.390 2194.060 2273.710 2194.120 ;
        RECT 1414.110 2180.320 1414.430 2180.380 ;
        RECT 2267.410 2180.320 2267.730 2180.380 ;
        RECT 1414.110 2180.180 2267.730 2180.320 ;
        RECT 1414.110 2180.120 1414.430 2180.180 ;
        RECT 2267.410 2180.120 2267.730 2180.180 ;
        RECT 1414.110 2166.380 1414.430 2166.440 ;
        RECT 2266.490 2166.380 2266.810 2166.440 ;
        RECT 1414.110 2166.240 2266.810 2166.380 ;
        RECT 1414.110 2166.180 1414.430 2166.240 ;
        RECT 2266.490 2166.180 2266.810 2166.240 ;
        RECT 1414.110 2159.580 1414.430 2159.640 ;
        RECT 1459.650 2159.580 1459.970 2159.640 ;
        RECT 1414.110 2159.440 1459.970 2159.580 ;
        RECT 1414.110 2159.380 1414.430 2159.440 ;
        RECT 1459.650 2159.380 1459.970 2159.440 ;
        RECT 1414.110 2145.640 1414.430 2145.700 ;
        RECT 1452.750 2145.640 1453.070 2145.700 ;
        RECT 1414.110 2145.500 1453.070 2145.640 ;
        RECT 1414.110 2145.440 1414.430 2145.500 ;
        RECT 1452.750 2145.440 1453.070 2145.500 ;
        RECT 1414.110 2133.060 1414.430 2133.120 ;
        RECT 1438.490 2133.060 1438.810 2133.120 ;
        RECT 1414.110 2132.920 1438.810 2133.060 ;
        RECT 1414.110 2132.860 1414.430 2132.920 ;
        RECT 1438.490 2132.860 1438.810 2132.920 ;
        RECT 1412.270 2125.240 1412.590 2125.300 ;
        RECT 1431.590 2125.240 1431.910 2125.300 ;
        RECT 1412.270 2125.100 1431.910 2125.240 ;
        RECT 1412.270 2125.040 1412.590 2125.100 ;
        RECT 1431.590 2125.040 1431.910 2125.100 ;
        RECT 1410.430 2111.300 1410.750 2111.360 ;
        RECT 1424.690 2111.300 1425.010 2111.360 ;
        RECT 1410.430 2111.160 1425.010 2111.300 ;
        RECT 1410.430 2111.100 1410.750 2111.160 ;
        RECT 1424.690 2111.100 1425.010 2111.160 ;
        RECT 1408.590 2104.160 1408.910 2104.220 ;
        RECT 1417.790 2104.160 1418.110 2104.220 ;
        RECT 1408.590 2104.020 1418.110 2104.160 ;
        RECT 1408.590 2103.960 1408.910 2104.020 ;
        RECT 1417.790 2103.960 1418.110 2104.020 ;
        RECT 1414.110 2090.560 1414.430 2090.620 ;
        RECT 1472.990 2090.560 1473.310 2090.620 ;
        RECT 1414.110 2090.420 1473.310 2090.560 ;
        RECT 1414.110 2090.360 1414.430 2090.420 ;
        RECT 1472.990 2090.360 1473.310 2090.420 ;
        RECT 1414.110 2083.760 1414.430 2083.820 ;
        RECT 1580.170 2083.760 1580.490 2083.820 ;
        RECT 1414.110 2083.620 1580.490 2083.760 ;
        RECT 1414.110 2083.560 1414.430 2083.620 ;
        RECT 1580.170 2083.560 1580.490 2083.620 ;
        RECT 1409.510 2069.820 1409.830 2069.880 ;
        RECT 1997.390 2069.820 1997.710 2069.880 ;
        RECT 1409.510 2069.680 1997.710 2069.820 ;
        RECT 1409.510 2069.620 1409.830 2069.680 ;
        RECT 1997.390 2069.620 1997.710 2069.680 ;
        RECT 1414.110 2056.220 1414.430 2056.280 ;
        RECT 1990.490 2056.220 1990.810 2056.280 ;
        RECT 1414.110 2056.080 1990.810 2056.220 ;
        RECT 1414.110 2056.020 1414.430 2056.080 ;
        RECT 1990.490 2056.020 1990.810 2056.080 ;
        RECT 1410.430 2049.080 1410.750 2049.140 ;
        RECT 1976.690 2049.080 1977.010 2049.140 ;
        RECT 1410.430 2048.940 1977.010 2049.080 ;
        RECT 1410.430 2048.880 1410.750 2048.940 ;
        RECT 1976.690 2048.880 1977.010 2048.940 ;
        RECT 1414.110 2035.480 1414.430 2035.540 ;
        RECT 1969.790 2035.480 1970.110 2035.540 ;
        RECT 1414.110 2035.340 1970.110 2035.480 ;
        RECT 1414.110 2035.280 1414.430 2035.340 ;
        RECT 1969.790 2035.280 1970.110 2035.340 ;
        RECT 1414.110 2028.340 1414.430 2028.400 ;
        RECT 1962.890 2028.340 1963.210 2028.400 ;
        RECT 1414.110 2028.200 1963.210 2028.340 ;
        RECT 1414.110 2028.140 1414.430 2028.200 ;
        RECT 1962.890 2028.140 1963.210 2028.200 ;
        RECT 1409.510 2014.740 1409.830 2014.800 ;
        RECT 1955.990 2014.740 1956.310 2014.800 ;
        RECT 1409.510 2014.600 1956.310 2014.740 ;
        RECT 1409.510 2014.540 1409.830 2014.600 ;
        RECT 1955.990 2014.540 1956.310 2014.600 ;
        RECT 1414.110 2000.800 1414.430 2000.860 ;
        RECT 1942.190 2000.800 1942.510 2000.860 ;
        RECT 1414.110 2000.660 1942.510 2000.800 ;
        RECT 1414.110 2000.600 1414.430 2000.660 ;
        RECT 1942.190 2000.600 1942.510 2000.660 ;
        RECT 1410.430 1994.000 1410.750 1994.060 ;
        RECT 2228.770 1994.000 2229.090 1994.060 ;
        RECT 1410.430 1993.860 2229.090 1994.000 ;
        RECT 1410.430 1993.800 1410.750 1993.860 ;
        RECT 2228.770 1993.800 2229.090 1993.860 ;
        RECT 1410.430 1979.380 1410.750 1979.440 ;
        RECT 1425.150 1979.380 1425.470 1979.440 ;
        RECT 1410.430 1979.240 1425.470 1979.380 ;
        RECT 1410.430 1979.180 1410.750 1979.240 ;
        RECT 1425.150 1979.180 1425.470 1979.240 ;
        RECT 1411.350 1973.260 1411.670 1973.320 ;
        RECT 2011.190 1973.260 2011.510 1973.320 ;
        RECT 1411.350 1973.120 2011.510 1973.260 ;
        RECT 1411.350 1973.060 1411.670 1973.120 ;
        RECT 2011.190 1973.060 2011.510 1973.120 ;
        RECT 1409.510 1959.660 1409.830 1959.720 ;
        RECT 1601.330 1959.660 1601.650 1959.720 ;
        RECT 1409.510 1959.520 1601.650 1959.660 ;
        RECT 1409.510 1959.460 1409.830 1959.520 ;
        RECT 1601.330 1959.460 1601.650 1959.520 ;
        RECT 1412.270 1949.120 1412.590 1949.180 ;
        RECT 1432.050 1949.120 1432.370 1949.180 ;
        RECT 1412.270 1948.980 1432.370 1949.120 ;
        RECT 1412.270 1948.920 1412.590 1948.980 ;
        RECT 1432.050 1948.920 1432.370 1948.980 ;
        RECT 1410.430 1938.920 1410.750 1938.980 ;
        RECT 1593.970 1938.920 1594.290 1938.980 ;
        RECT 1410.430 1938.780 1594.290 1938.920 ;
        RECT 1410.430 1938.720 1410.750 1938.780 ;
        RECT 1593.970 1938.720 1594.290 1938.780 ;
        RECT 1414.110 1923.280 1414.430 1923.340 ;
        RECT 1438.950 1923.280 1439.270 1923.340 ;
        RECT 1414.110 1923.140 1439.270 1923.280 ;
        RECT 1414.110 1923.080 1414.430 1923.140 ;
        RECT 1438.950 1923.080 1439.270 1923.140 ;
        RECT 1414.110 1918.180 1414.430 1918.240 ;
        RECT 2252.690 1918.180 2253.010 1918.240 ;
        RECT 1414.110 1918.040 2253.010 1918.180 ;
        RECT 1414.110 1917.980 1414.430 1918.040 ;
        RECT 2252.690 1917.980 2253.010 1918.040 ;
        RECT 1414.110 1904.240 1414.430 1904.300 ;
        RECT 2245.790 1904.240 2246.110 1904.300 ;
        RECT 1414.110 1904.100 2246.110 1904.240 ;
        RECT 1414.110 1904.040 1414.430 1904.100 ;
        RECT 2245.790 1904.040 2246.110 1904.100 ;
        RECT 1412.270 1897.440 1412.590 1897.500 ;
        RECT 2238.890 1897.440 2239.210 1897.500 ;
        RECT 1412.270 1897.300 2239.210 1897.440 ;
        RECT 1412.270 1897.240 1412.590 1897.300 ;
        RECT 2238.890 1897.240 2239.210 1897.300 ;
        RECT 1410.430 1883.500 1410.750 1883.560 ;
        RECT 2231.990 1883.500 2232.310 1883.560 ;
        RECT 1410.430 1883.360 2232.310 1883.500 ;
        RECT 1410.430 1883.300 1410.750 1883.360 ;
        RECT 2231.990 1883.300 2232.310 1883.360 ;
        RECT 1414.110 1869.900 1414.430 1869.960 ;
        RECT 1794.070 1869.900 1794.390 1869.960 ;
        RECT 1414.110 1869.760 1794.390 1869.900 ;
        RECT 1414.110 1869.700 1414.430 1869.760 ;
        RECT 1794.070 1869.700 1794.390 1869.760 ;
        RECT 1412.730 1862.760 1413.050 1862.820 ;
        RECT 1787.170 1862.760 1787.490 1862.820 ;
        RECT 1412.730 1862.620 1787.490 1862.760 ;
        RECT 1412.730 1862.560 1413.050 1862.620 ;
        RECT 1787.170 1862.560 1787.490 1862.620 ;
        RECT 1414.110 1849.160 1414.430 1849.220 ;
        RECT 1780.270 1849.160 1780.590 1849.220 ;
        RECT 1414.110 1849.020 1780.590 1849.160 ;
        RECT 1414.110 1848.960 1414.430 1849.020 ;
        RECT 1780.270 1848.960 1780.590 1849.020 ;
        RECT 1412.270 1842.360 1412.590 1842.420 ;
        RECT 1773.830 1842.360 1774.150 1842.420 ;
        RECT 1412.270 1842.220 1774.150 1842.360 ;
        RECT 1412.270 1842.160 1412.590 1842.220 ;
        RECT 1773.830 1842.160 1774.150 1842.220 ;
        RECT 1410.430 1828.420 1410.750 1828.480 ;
        RECT 1766.470 1828.420 1766.790 1828.480 ;
        RECT 1410.430 1828.280 1766.790 1828.420 ;
        RECT 1410.430 1828.220 1410.750 1828.280 ;
        RECT 1766.470 1828.220 1766.790 1828.280 ;
        RECT 1414.110 1814.480 1414.430 1814.540 ;
        RECT 1760.030 1814.480 1760.350 1814.540 ;
        RECT 1414.110 1814.340 1760.350 1814.480 ;
        RECT 1414.110 1814.280 1414.430 1814.340 ;
        RECT 1760.030 1814.280 1760.350 1814.340 ;
        RECT 1412.730 1807.680 1413.050 1807.740 ;
        RECT 1760.950 1807.680 1761.270 1807.740 ;
        RECT 1412.730 1807.540 1761.270 1807.680 ;
        RECT 1412.730 1807.480 1413.050 1807.540 ;
        RECT 1760.950 1807.480 1761.270 1807.540 ;
        RECT 1414.110 1793.740 1414.430 1793.800 ;
        RECT 1752.670 1793.740 1752.990 1793.800 ;
        RECT 1414.110 1793.600 1752.990 1793.740 ;
        RECT 1414.110 1793.540 1414.430 1793.600 ;
        RECT 1752.670 1793.540 1752.990 1793.600 ;
        RECT 1412.270 1786.940 1412.590 1787.000 ;
        RECT 1745.770 1786.940 1746.090 1787.000 ;
        RECT 1412.270 1786.800 1746.090 1786.940 ;
        RECT 1412.270 1786.740 1412.590 1786.800 ;
        RECT 1745.770 1786.740 1746.090 1786.800 ;
        RECT 1410.430 1773.340 1410.750 1773.400 ;
        RECT 1738.870 1773.340 1739.190 1773.400 ;
        RECT 1410.430 1773.200 1739.190 1773.340 ;
        RECT 1410.430 1773.140 1410.750 1773.200 ;
        RECT 1738.870 1773.140 1739.190 1773.200 ;
        RECT 1414.110 1759.400 1414.430 1759.460 ;
        RECT 1731.970 1759.400 1732.290 1759.460 ;
        RECT 1414.110 1759.260 1732.290 1759.400 ;
        RECT 1414.110 1759.200 1414.430 1759.260 ;
        RECT 1731.970 1759.200 1732.290 1759.260 ;
        RECT 1412.730 1752.600 1413.050 1752.660 ;
        RECT 1725.070 1752.600 1725.390 1752.660 ;
        RECT 1412.730 1752.460 1725.390 1752.600 ;
        RECT 1412.730 1752.400 1413.050 1752.460 ;
        RECT 1725.070 1752.400 1725.390 1752.460 ;
        RECT 1414.110 1738.660 1414.430 1738.720 ;
        RECT 1718.630 1738.660 1718.950 1738.720 ;
        RECT 1414.110 1738.520 1718.950 1738.660 ;
        RECT 1414.110 1738.460 1414.430 1738.520 ;
        RECT 1718.630 1738.460 1718.950 1738.520 ;
        RECT 1412.270 1731.860 1412.590 1731.920 ;
        RECT 1718.170 1731.860 1718.490 1731.920 ;
        RECT 1412.270 1731.720 1718.490 1731.860 ;
        RECT 1412.270 1731.660 1412.590 1731.720 ;
        RECT 1718.170 1731.660 1718.490 1731.720 ;
        RECT 1414.110 1717.920 1414.430 1717.980 ;
        RECT 1711.270 1717.920 1711.590 1717.980 ;
        RECT 1414.110 1717.780 1711.590 1717.920 ;
        RECT 1414.110 1717.720 1414.430 1717.780 ;
        RECT 1711.270 1717.720 1711.590 1717.780 ;
        RECT 1414.110 1704.320 1414.430 1704.380 ;
        RECT 1704.370 1704.320 1704.690 1704.380 ;
        RECT 1414.110 1704.180 1704.690 1704.320 ;
        RECT 1414.110 1704.120 1414.430 1704.180 ;
        RECT 1704.370 1704.120 1704.690 1704.180 ;
        RECT 1414.110 1697.180 1414.430 1697.240 ;
        RECT 1697.470 1697.180 1697.790 1697.240 ;
        RECT 1414.110 1697.040 1697.790 1697.180 ;
        RECT 1414.110 1696.980 1414.430 1697.040 ;
        RECT 1697.470 1696.980 1697.790 1697.040 ;
        RECT 1414.110 1683.580 1414.430 1683.640 ;
        RECT 1690.570 1683.580 1690.890 1683.640 ;
        RECT 1414.110 1683.440 1690.890 1683.580 ;
        RECT 1414.110 1683.380 1414.430 1683.440 ;
        RECT 1690.570 1683.380 1690.890 1683.440 ;
        RECT 1411.810 1676.440 1412.130 1676.500 ;
        RECT 1684.130 1676.440 1684.450 1676.500 ;
        RECT 1411.810 1676.300 1684.450 1676.440 ;
        RECT 1411.810 1676.240 1412.130 1676.300 ;
        RECT 1684.130 1676.240 1684.450 1676.300 ;
        RECT 1414.110 1662.840 1414.430 1662.900 ;
        RECT 1683.670 1662.840 1683.990 1662.900 ;
        RECT 1414.110 1662.700 1683.990 1662.840 ;
        RECT 1414.110 1662.640 1414.430 1662.700 ;
        RECT 1683.670 1662.640 1683.990 1662.700 ;
        RECT 1414.110 1648.900 1414.430 1648.960 ;
        RECT 1676.770 1648.900 1677.090 1648.960 ;
        RECT 1414.110 1648.760 1677.090 1648.900 ;
        RECT 1414.110 1648.700 1414.430 1648.760 ;
        RECT 1676.770 1648.700 1677.090 1648.760 ;
        RECT 1414.110 1642.100 1414.430 1642.160 ;
        RECT 1669.870 1642.100 1670.190 1642.160 ;
        RECT 1414.110 1641.960 1670.190 1642.100 ;
        RECT 1414.110 1641.900 1414.430 1641.960 ;
        RECT 1669.870 1641.900 1670.190 1641.960 ;
        RECT 1414.110 1628.160 1414.430 1628.220 ;
        RECT 1662.970 1628.160 1663.290 1628.220 ;
        RECT 1414.110 1628.020 1663.290 1628.160 ;
        RECT 1414.110 1627.960 1414.430 1628.020 ;
        RECT 1662.970 1627.960 1663.290 1628.020 ;
        RECT 1411.810 1621.360 1412.130 1621.420 ;
        RECT 1452.290 1621.360 1452.610 1621.420 ;
        RECT 1411.810 1621.220 1452.610 1621.360 ;
        RECT 1411.810 1621.160 1412.130 1621.220 ;
        RECT 1452.290 1621.160 1452.610 1621.220 ;
        RECT 1414.110 1607.760 1414.430 1607.820 ;
        RECT 1649.630 1607.760 1649.950 1607.820 ;
        RECT 1414.110 1607.620 1649.950 1607.760 ;
        RECT 1414.110 1607.560 1414.430 1607.620 ;
        RECT 1649.630 1607.560 1649.950 1607.620 ;
        RECT 1414.110 1593.820 1414.430 1593.880 ;
        RECT 1459.190 1593.820 1459.510 1593.880 ;
        RECT 1414.110 1593.680 1459.510 1593.820 ;
        RECT 1414.110 1593.620 1414.430 1593.680 ;
        RECT 1459.190 1593.620 1459.510 1593.680 ;
        RECT 1414.110 1587.020 1414.430 1587.080 ;
        RECT 1610.990 1587.020 1611.310 1587.080 ;
        RECT 1414.110 1586.880 1611.310 1587.020 ;
        RECT 1414.110 1586.820 1414.430 1586.880 ;
        RECT 1610.990 1586.820 1611.310 1586.880 ;
        RECT 1414.110 1573.080 1414.430 1573.140 ;
        RECT 1635.370 1573.080 1635.690 1573.140 ;
        RECT 1414.110 1572.940 1635.690 1573.080 ;
        RECT 1414.110 1572.880 1414.430 1572.940 ;
        RECT 1635.370 1572.880 1635.690 1572.940 ;
        RECT 1411.810 1566.280 1412.130 1566.340 ;
        RECT 1628.470 1566.280 1628.790 1566.340 ;
        RECT 1411.810 1566.140 1628.790 1566.280 ;
        RECT 1411.810 1566.080 1412.130 1566.140 ;
        RECT 1628.470 1566.080 1628.790 1566.140 ;
        RECT 1409.510 1552.340 1409.830 1552.400 ;
        RECT 1617.890 1552.340 1618.210 1552.400 ;
        RECT 1409.510 1552.200 1618.210 1552.340 ;
        RECT 1409.510 1552.140 1409.830 1552.200 ;
        RECT 1617.890 1552.140 1618.210 1552.200 ;
        RECT 1414.110 1538.740 1414.430 1538.800 ;
        RECT 1514.390 1538.740 1514.710 1538.800 ;
        RECT 1414.110 1538.600 1514.710 1538.740 ;
        RECT 1414.110 1538.540 1414.430 1538.600 ;
        RECT 1514.390 1538.540 1514.710 1538.600 ;
        RECT 1410.430 1531.600 1410.750 1531.660 ;
        RECT 1607.770 1531.600 1608.090 1531.660 ;
        RECT 1410.430 1531.460 1608.090 1531.600 ;
        RECT 1410.430 1531.400 1410.750 1531.460 ;
        RECT 1607.770 1531.400 1608.090 1531.460 ;
      LAYER via ;
        RECT 2539.300 3266.760 2539.560 3267.020 ;
        RECT 2566.900 3266.760 2567.160 3267.020 ;
        RECT 2566.900 3264.040 2567.160 3264.300 ;
        RECT 2594.500 3264.040 2594.760 3264.300 ;
        RECT 646.400 3263.700 646.660 3263.960 ;
        RECT 668.020 3263.700 668.280 3263.960 ;
        RECT 697.920 3263.700 698.180 3263.960 ;
        RECT 1295.920 3263.700 1296.180 3263.960 ;
        RECT 1318.920 3263.700 1319.180 3263.960 ;
        RECT 1345.600 3263.700 1345.860 3263.960 ;
        RECT 1892.540 3263.700 1892.800 3263.960 ;
        RECT 1917.380 3263.700 1917.640 3263.960 ;
        RECT 1946.820 3263.700 1947.080 3263.960 ;
        RECT 2539.300 3263.700 2539.560 3263.960 ;
        RECT 697.000 3251.800 697.260 3252.060 ;
        RECT 1331.800 3251.800 1332.060 3252.060 ;
        RECT 1410.000 3251.800 1410.260 3252.060 ;
        RECT 1945.900 3251.800 1946.160 3252.060 ;
        RECT 2582.080 3251.800 2582.340 3252.060 ;
        RECT 710.340 3229.360 710.600 3229.620 ;
        RECT 938.500 3229.360 938.760 3229.620 ;
        RECT 703.440 3222.220 703.700 3222.480 ;
        RECT 938.500 3222.220 938.760 3222.480 ;
        RECT 689.640 3215.420 689.900 3215.680 ;
        RECT 938.500 3215.420 938.760 3215.680 ;
        RECT 803.720 3208.620 803.980 3208.880 ;
        RECT 938.500 3208.620 938.760 3208.880 ;
        RECT 796.820 3201.480 797.080 3201.740 ;
        RECT 938.500 3201.480 938.760 3201.740 ;
        RECT 889.740 2898.200 890.000 2898.460 ;
        RECT 938.500 2898.200 938.760 2898.460 ;
        RECT 1331.800 3250.100 1332.060 3250.360 ;
        RECT 1407.700 3250.100 1407.960 3250.360 ;
        RECT 1410.000 3250.100 1410.260 3250.360 ;
        RECT 1459.680 3229.360 1459.940 3229.620 ;
        RECT 1536.960 3229.360 1537.220 3229.620 ;
        RECT 1452.780 3222.220 1453.040 3222.480 ;
        RECT 1535.580 3222.220 1535.840 3222.480 ;
        RECT 1438.520 3215.420 1438.780 3215.680 ;
        RECT 1535.580 3215.420 1535.840 3215.680 ;
        RECT 1431.620 3208.620 1431.880 3208.880 ;
        RECT 1538.340 3208.620 1538.600 3208.880 ;
        RECT 1424.720 3201.480 1424.980 3201.740 ;
        RECT 1538.340 3201.480 1538.600 3201.740 ;
        RECT 1417.820 3194.680 1418.080 3194.940 ;
        RECT 1533.280 3194.680 1533.540 3194.940 ;
        RECT 1473.020 3187.880 1473.280 3188.140 ;
        RECT 1497.860 3187.880 1498.120 3188.140 ;
        RECT 1350.200 2901.260 1350.460 2901.520 ;
        RECT 1408.160 2901.260 1408.420 2901.520 ;
        RECT 1425.180 2898.200 1425.440 2898.460 ;
        RECT 1534.660 2898.200 1534.920 2898.460 ;
        RECT 1410.920 2891.060 1411.180 2891.320 ;
        RECT 1531.900 2891.060 1532.160 2891.320 ;
        RECT 1408.620 2808.100 1408.880 2808.360 ;
        RECT 1410.920 2808.100 1411.180 2808.360 ;
        RECT 1997.420 3229.360 1997.680 3229.620 ;
        RECT 2187.400 3229.360 2187.660 3229.620 ;
        RECT 1990.520 3222.220 1990.780 3222.480 ;
        RECT 2187.400 3222.220 2187.660 3222.480 ;
        RECT 1976.720 3215.420 1976.980 3215.680 ;
        RECT 2187.400 3215.420 2187.660 3215.680 ;
        RECT 1969.820 3208.620 1970.080 3208.880 ;
        RECT 2187.400 3208.620 2187.660 3208.880 ;
        RECT 1962.920 3201.480 1963.180 3201.740 ;
        RECT 2187.400 3201.480 2187.660 3201.740 ;
        RECT 1956.020 3194.680 1956.280 3194.940 ;
        RECT 2187.400 3194.680 2187.660 3194.940 ;
        RECT 1942.220 3187.880 1942.480 3188.140 ;
        RECT 2187.400 3187.880 2187.660 3188.140 ;
        RECT 2011.220 2898.200 2011.480 2898.460 ;
        RECT 2187.400 2898.200 2187.660 2898.460 ;
        RECT 298.180 2804.360 298.440 2804.620 ;
        RECT 944.940 2804.360 945.200 2804.620 ;
        RECT 1408.620 2804.360 1408.880 2804.620 ;
        RECT 1531.440 2804.360 1531.700 2804.620 ;
        RECT 2190.620 2804.360 2190.880 2804.620 ;
        RECT 396.620 2794.160 396.880 2794.420 ;
        RECT 407.200 2794.160 407.460 2794.420 ;
        RECT 407.660 2794.160 407.920 2794.420 ;
        RECT 434.340 2794.160 434.600 2794.420 ;
        RECT 403.520 2793.820 403.780 2794.080 ;
        RECT 450.440 2794.160 450.700 2794.420 ;
        RECT 455.040 2794.160 455.300 2794.420 ;
        RECT 1677.260 2794.160 1677.520 2794.420 ;
        RECT 1721.420 2794.160 1721.680 2794.420 ;
        RECT 1776.620 2794.160 1776.880 2794.420 ;
        RECT 2415.100 2794.160 2415.360 2794.420 ;
        RECT 439.400 2793.820 439.660 2794.080 ;
        RECT 483.100 2793.820 483.360 2794.080 ;
        RECT 1117.900 2793.820 1118.160 2794.080 ;
        RECT 1159.760 2793.820 1160.020 2794.080 ;
        RECT 1718.660 2793.820 1718.920 2794.080 ;
        RECT 1759.600 2793.820 1759.860 2794.080 ;
        RECT 2294.120 2793.820 2294.380 2794.080 ;
        RECT 2340.120 2793.820 2340.380 2794.080 ;
        RECT 2385.660 2793.820 2385.920 2794.080 ;
        RECT 2428.900 2793.820 2429.160 2794.080 ;
        RECT 397.540 2793.480 397.800 2793.740 ;
        RECT 444.920 2793.480 445.180 2793.740 ;
        RECT 386.960 2793.140 387.220 2793.400 ;
        RECT 407.660 2793.140 407.920 2793.400 ;
        RECT 408.120 2793.140 408.380 2793.400 ;
        RECT 456.880 2793.140 457.140 2793.400 ;
        RECT 501.500 2793.480 501.760 2793.740 ;
        RECT 1083.860 2793.480 1084.120 2793.740 ;
        RECT 1128.940 2793.480 1129.200 2793.740 ;
        RECT 1131.700 2793.480 1131.960 2793.740 ;
        RECT 1135.840 2793.480 1136.100 2793.740 ;
        RECT 1180.000 2793.480 1180.260 2793.740 ;
        RECT 1721.420 2793.480 1721.680 2793.740 ;
        RECT 1766.500 2793.480 1766.760 2793.740 ;
        RECT 2303.320 2793.480 2303.580 2793.740 ;
        RECT 2342.880 2793.480 2343.140 2793.740 ;
        RECT 2377.840 2793.480 2378.100 2793.740 ;
        RECT 2422.000 2793.480 2422.260 2793.740 ;
        RECT 476.660 2793.140 476.920 2793.400 ;
        RECT 526.800 2793.140 527.060 2793.400 ;
        RECT 530.480 2793.140 530.740 2793.400 ;
        RECT 1076.500 2793.140 1076.760 2793.400 ;
        RECT 1122.040 2793.140 1122.300 2793.400 ;
        RECT 1166.200 2793.140 1166.460 2793.400 ;
        RECT 1694.740 2793.140 1695.000 2793.400 ;
        RECT 1741.660 2793.140 1741.920 2793.400 ;
        RECT 1787.200 2793.140 1787.460 2793.400 ;
        RECT 378.680 2792.800 378.940 2793.060 ;
        RECT 421.460 2792.800 421.720 2793.060 ;
        RECT 467.920 2792.800 468.180 2793.060 ;
        RECT 542.900 2792.800 543.160 2793.060 ;
        RECT 1056.720 2792.800 1056.980 2793.060 ;
        RECT 1062.700 2792.800 1062.960 2793.060 ;
        RECT 1065.920 2792.800 1066.180 2793.060 ;
        RECT 1111.460 2792.800 1111.720 2793.060 ;
        RECT 1159.300 2792.800 1159.560 2793.060 ;
        RECT 1683.240 2792.800 1683.500 2793.060 ;
        RECT 1731.540 2792.800 1731.800 2793.060 ;
        RECT 1734.760 2792.800 1735.020 2793.060 ;
        RECT 1780.300 2792.800 1780.560 2793.060 ;
        RECT 1783.980 2792.800 1784.240 2793.060 ;
        RECT 2422.460 2793.140 2422.720 2793.400 ;
        RECT 2267.440 2792.800 2267.700 2793.060 ;
        RECT 2314.820 2792.800 2315.080 2793.060 ;
        RECT 2318.040 2792.800 2318.300 2793.060 ;
        RECT 2321.720 2792.800 2321.980 2793.060 ;
        RECT 2367.720 2792.800 2367.980 2793.060 ;
        RECT 2415.100 2792.800 2415.360 2793.060 ;
        RECT 362.120 2792.460 362.380 2792.720 ;
        RECT 408.120 2792.460 408.380 2792.720 ;
        RECT 434.340 2792.460 434.600 2792.720 ;
        RECT 476.660 2792.460 476.920 2792.720 ;
        RECT 483.100 2792.460 483.360 2792.720 ;
        RECT 531.400 2792.460 531.660 2792.720 ;
        RECT 537.380 2792.460 537.640 2792.720 ;
        RECT 539.220 2792.460 539.480 2792.720 ;
        RECT 1048.900 2792.460 1049.160 2792.720 ;
        RECT 1055.800 2792.460 1056.060 2792.720 ;
        RECT 1059.480 2792.460 1059.740 2792.720 ;
        RECT 1105.480 2792.460 1105.740 2792.720 ;
        RECT 1152.400 2792.460 1152.660 2792.720 ;
        RECT 1686.920 2792.460 1687.180 2792.720 ;
        RECT 2301.940 2792.460 2302.200 2792.720 ;
        RECT 2304.240 2792.460 2304.500 2792.720 ;
        RECT 2350.240 2792.460 2350.500 2792.720 ;
        RECT 2397.160 2792.460 2397.420 2792.720 ;
        RECT 2442.700 2792.460 2442.960 2792.720 ;
        RECT 380.060 2792.120 380.320 2792.380 ;
        RECT 426.980 2792.120 427.240 2792.380 ;
        RECT 472.980 2792.120 473.240 2792.380 ;
        RECT 519.900 2792.120 520.160 2792.380 ;
        RECT 523.580 2792.120 523.840 2792.380 ;
        RECT 834.540 2792.120 834.800 2792.380 ;
        RECT 1007.500 2792.120 1007.760 2792.380 ;
        RECT 1656.560 2792.120 1656.820 2792.380 ;
        RECT 1658.860 2792.120 1659.120 2792.380 ;
        RECT 1704.860 2792.120 1705.120 2792.380 ;
        RECT 1752.700 2792.120 1752.960 2792.380 ;
        RECT 2266.520 2792.120 2266.780 2792.380 ;
        RECT 2308.840 2792.120 2309.100 2792.380 ;
        RECT 2356.220 2792.120 2356.480 2792.380 ;
        RECT 2402.220 2792.120 2402.480 2792.380 ;
        RECT 368.560 2791.780 368.820 2792.040 ;
        RECT 414.560 2791.780 414.820 2792.040 ;
        RECT 462.400 2791.780 462.660 2792.040 ;
        RECT 503.800 2791.780 504.060 2792.040 ;
        RECT 827.640 2791.780 827.900 2792.040 ;
        RECT 1001.060 2791.780 1001.320 2792.040 ;
        RECT 1090.300 2791.780 1090.560 2792.040 ;
        RECT 1094.440 2791.780 1094.700 2792.040 ;
        RECT 1138.600 2791.780 1138.860 2792.040 ;
        RECT 1139.060 2791.780 1139.320 2792.040 ;
        RECT 1147.340 2791.780 1147.600 2792.040 ;
        RECT 1193.800 2791.780 1194.060 2792.040 ;
        RECT 1663.460 2791.780 1663.720 2792.040 ;
        RECT 1712.680 2791.780 1712.940 2792.040 ;
        RECT 1739.820 2791.780 1740.080 2792.040 ;
        RECT 1790.880 2791.780 1791.140 2792.040 ;
        RECT 2277.100 2791.780 2277.360 2792.040 ;
        RECT 2318.040 2791.780 2318.300 2792.040 ;
        RECT 2361.280 2791.780 2361.540 2792.040 ;
        RECT 2408.200 2791.780 2408.460 2792.040 ;
        RECT 379.140 2791.440 379.400 2791.700 ;
        RECT 400.300 2791.440 400.560 2791.700 ;
        RECT 444.920 2791.440 445.180 2791.700 ;
        RECT 491.380 2791.440 491.640 2791.700 ;
        RECT 539.220 2791.440 539.480 2791.700 ;
        RECT 813.840 2791.440 814.100 2791.700 ;
        RECT 993.700 2791.440 993.960 2791.700 ;
        RECT 1069.600 2791.440 1069.860 2791.700 ;
        RECT 1117.900 2791.440 1118.160 2791.700 ;
        RECT 1128.940 2791.440 1129.200 2791.700 ;
        RECT 1173.100 2791.440 1173.360 2791.700 ;
        RECT 1699.340 2791.440 1699.600 2791.700 ;
        RECT 1747.640 2791.440 1747.900 2791.700 ;
        RECT 1788.580 2791.440 1788.840 2791.700 ;
        RECT 1797.320 2791.440 1797.580 2791.700 ;
        RECT 2284.000 2791.440 2284.260 2791.700 ;
        RECT 2325.860 2791.440 2326.120 2791.700 ;
        RECT 2374.160 2791.440 2374.420 2791.700 ;
        RECT 2387.960 2791.440 2388.220 2791.700 ;
        RECT 2391.640 2791.440 2391.900 2791.700 ;
        RECT 2435.800 2791.440 2436.060 2791.700 ;
        RECT 392.480 2791.100 392.740 2791.360 ;
        RECT 439.400 2791.100 439.660 2791.360 ;
        RECT 455.040 2791.100 455.300 2791.360 ;
        RECT 497.820 2791.100 498.080 2791.360 ;
        RECT 542.900 2791.100 543.160 2791.360 ;
        RECT 806.940 2791.100 807.200 2791.360 ;
        RECT 986.800 2791.100 987.060 2791.360 ;
        RECT 1083.400 2791.100 1083.660 2791.360 ;
        RECT 1088.000 2791.100 1088.260 2791.360 ;
        RECT 1131.700 2791.100 1131.960 2791.360 ;
        RECT 1138.600 2791.100 1138.860 2791.360 ;
        RECT 1186.900 2791.100 1187.160 2791.360 ;
        RECT 1459.220 2791.100 1459.480 2791.360 ;
        RECT 1649.200 2791.100 1649.460 2791.360 ;
        RECT 1670.360 2791.100 1670.620 2791.360 ;
        RECT 1718.660 2791.100 1718.920 2791.360 ;
        RECT 1731.540 2791.100 1731.800 2791.360 ;
        RECT 1773.400 2791.100 1773.660 2791.360 ;
        RECT 1797.780 2791.100 1798.040 2791.360 ;
        RECT 2290.900 2791.100 2291.160 2791.360 ;
        RECT 2335.520 2791.100 2335.780 2791.360 ;
        RECT 2442.700 2791.100 2442.960 2791.360 ;
        RECT 2218.220 2790.760 2218.480 2791.020 ;
        RECT 2297.800 2790.760 2298.060 2791.020 ;
        RECT 2328.620 2790.760 2328.880 2791.020 ;
        RECT 2435.800 2790.760 2436.060 2791.020 ;
        RECT 641.340 2790.420 641.600 2790.680 ;
        RECT 979.900 2790.420 980.160 2790.680 ;
        RECT 1024.520 2790.420 1024.780 2790.680 ;
        RECT 1069.600 2790.420 1069.860 2790.680 ;
        RECT 1452.320 2790.420 1452.580 2790.680 ;
        RECT 1656.100 2790.420 1656.360 2790.680 ;
        RECT 1749.020 2790.420 1749.280 2790.680 ;
        RECT 2263.300 2790.420 2263.560 2790.680 ;
        RECT 2273.420 2790.420 2273.680 2790.680 ;
        RECT 2321.260 2790.420 2321.520 2790.680 ;
        RECT 2321.720 2790.420 2321.980 2790.680 ;
        RECT 2428.900 2790.420 2429.160 2790.680 ;
        RECT 403.520 2790.080 403.780 2790.340 ;
        RECT 414.100 2790.080 414.360 2790.340 ;
        RECT 503.800 2790.080 504.060 2790.340 ;
        RECT 509.320 2790.080 509.580 2790.340 ;
        RECT 993.700 2790.080 993.960 2790.340 ;
        RECT 1031.420 2790.080 1031.680 2790.340 ;
        RECT 1076.500 2790.080 1076.760 2790.340 ;
        RECT 1611.020 2790.080 1611.280 2790.340 ;
        RECT 1642.300 2790.080 1642.560 2790.340 ;
        RECT 1645.520 2790.080 1645.780 2790.340 ;
        RECT 1686.920 2790.080 1687.180 2790.340 ;
        RECT 1762.820 2790.080 1763.080 2790.340 ;
        RECT 2380.600 2790.080 2380.860 2790.340 ;
        RECT 501.500 2789.740 501.760 2790.000 ;
        RECT 986.800 2789.740 987.060 2790.000 ;
        RECT 1046.140 2789.740 1046.400 2790.000 ;
        RECT 1083.400 2789.740 1083.660 2790.000 ;
        RECT 1638.620 2789.740 1638.880 2790.000 ;
        RECT 1683.240 2789.740 1683.500 2790.000 ;
        RECT 1763.280 2789.740 1763.540 2790.000 ;
        RECT 2387.500 2789.740 2387.760 2790.000 ;
        RECT 358.440 2789.400 358.700 2789.660 ;
        RECT 393.400 2789.400 393.660 2789.660 ;
        RECT 1010.720 2789.400 1010.980 2789.660 ;
        RECT 1055.800 2789.400 1056.060 2789.660 ;
        RECT 1611.480 2789.400 1611.740 2789.660 ;
        RECT 1656.560 2789.400 1656.820 2789.660 ;
        RECT 1763.740 2789.400 1764.000 2789.660 ;
        RECT 2394.400 2789.400 2394.660 2789.660 ;
        RECT 351.540 2789.060 351.800 2789.320 ;
        RECT 386.500 2789.060 386.760 2789.320 ;
        RECT 467.920 2789.060 468.180 2789.320 ;
        RECT 513.460 2789.060 513.720 2789.320 ;
        RECT 1007.500 2789.060 1007.760 2789.320 ;
        RECT 1017.620 2789.060 1017.880 2789.320 ;
        RECT 1062.700 2789.060 1062.960 2789.320 ;
        RECT 1514.420 2789.060 1514.680 2789.320 ;
        RECT 1614.700 2789.060 1614.960 2789.320 ;
        RECT 1618.380 2789.060 1618.640 2789.320 ;
        RECT 1663.460 2789.060 1663.720 2789.320 ;
        RECT 1769.720 2789.060 1769.980 2789.320 ;
        RECT 2402.680 2789.060 2402.940 2789.320 ;
        RECT 330.840 2788.720 331.100 2788.980 ;
        RECT 372.700 2788.720 372.960 2788.980 ;
        RECT 530.480 2788.720 530.740 2788.980 ;
        RECT 1028.200 2788.720 1028.460 2788.980 ;
        RECT 1438.980 2788.720 1439.240 2788.980 ;
        RECT 1587.100 2788.720 1587.360 2788.980 ;
        RECT 1624.820 2788.720 1625.080 2788.980 ;
        RECT 1670.360 2788.720 1670.620 2788.980 ;
        RECT 1783.520 2788.720 1783.780 2788.980 ;
        RECT 2415.100 2788.720 2415.360 2788.980 ;
        RECT 337.280 2788.380 337.540 2788.640 ;
        RECT 379.600 2788.380 379.860 2788.640 ;
        RECT 537.380 2788.380 537.640 2788.640 ;
        RECT 1035.100 2788.380 1035.360 2788.640 ;
        RECT 1038.320 2788.380 1038.580 2788.640 ;
        RECT 1083.860 2788.380 1084.120 2788.640 ;
        RECT 1432.080 2788.380 1432.340 2788.640 ;
        RECT 1600.900 2788.380 1601.160 2788.640 ;
        RECT 1631.720 2788.380 1631.980 2788.640 ;
        RECT 1677.260 2788.380 1677.520 2788.640 ;
        RECT 1770.180 2788.380 1770.440 2788.640 ;
        RECT 2408.200 2788.380 2408.460 2788.640 ;
        RECT 317.040 2788.040 317.300 2788.300 ;
        RECT 365.800 2788.040 366.060 2788.300 ;
        RECT 523.580 2788.040 523.840 2788.300 ;
        RECT 1014.400 2788.040 1014.660 2788.300 ;
        RECT 1045.220 2788.040 1045.480 2788.300 ;
        RECT 1090.300 2788.040 1090.560 2788.300 ;
        RECT 1646.440 2788.040 1646.700 2788.300 ;
        RECT 1694.740 2788.040 1695.000 2788.300 ;
        RECT 1790.420 2788.040 1790.680 2788.300 ;
        RECT 2270.200 2788.040 2270.460 2788.300 ;
        RECT 2280.320 2788.040 2280.580 2788.300 ;
        RECT 2325.860 2788.040 2326.120 2788.300 ;
        RECT 2342.880 2788.040 2343.140 2788.300 ;
        RECT 2387.960 2788.040 2388.220 2788.300 ;
        RECT 310.140 2787.700 310.400 2787.960 ;
        RECT 358.900 2787.700 359.160 2787.960 ;
        RECT 372.240 2787.700 372.500 2787.960 ;
        RECT 393.400 2787.700 393.660 2787.960 ;
        RECT 1052.120 2787.700 1052.380 2787.960 ;
        RECT 1100.420 2787.700 1100.680 2787.960 ;
        RECT 1139.060 2787.700 1139.320 2787.960 ;
        RECT 1652.420 2787.700 1652.680 2787.960 ;
        RECT 1699.340 2787.700 1699.600 2787.960 ;
        RECT 2252.720 2787.700 2252.980 2787.960 ;
        RECT 2256.860 2787.700 2257.120 2787.960 ;
        RECT 2287.220 2787.700 2287.480 2787.960 ;
        RECT 2332.760 2787.700 2333.020 2787.960 ;
        RECT 2373.240 2787.700 2373.500 2787.960 ;
        RECT 2374.160 2787.700 2374.420 2787.960 ;
        RECT 2415.100 2787.700 2415.360 2787.960 ;
        RECT 283.920 2718.340 284.180 2718.600 ;
        RECT 730.120 2718.340 730.380 2718.600 ;
        RECT 1034.640 2718.340 1034.900 2718.600 ;
        RECT 1103.640 2718.340 1103.900 2718.600 ;
        RECT 1145.040 2718.340 1145.300 2718.600 ;
        RECT 1300.980 2718.340 1301.240 2718.600 ;
        RECT 284.380 2718.000 284.640 2718.260 ;
        RECT 740.700 2718.000 740.960 2718.260 ;
        RECT 1027.740 2718.000 1028.000 2718.260 ;
        RECT 1093.520 2718.000 1093.780 2718.260 ;
        RECT 1138.140 2718.000 1138.400 2718.260 ;
        RECT 1290.400 2718.000 1290.660 2718.260 ;
        RECT 305.080 2717.660 305.340 2717.920 ;
        RECT 310.140 2717.660 310.400 2717.920 ;
        RECT 284.840 2717.320 285.100 2717.580 ;
        RECT 750.820 2717.660 751.080 2717.920 ;
        RECT 823.500 2717.660 823.760 2717.920 ;
        RECT 827.640 2717.660 827.900 2717.920 ;
        RECT 886.060 2717.660 886.320 2717.920 ;
        RECT 889.740 2717.660 890.000 2717.920 ;
        RECT 1041.540 2717.660 1041.800 2717.920 ;
        RECT 1114.220 2717.660 1114.480 2717.920 ;
        RECT 1158.840 2717.660 1159.100 2717.920 ;
        RECT 1321.680 2717.660 1321.940 2717.920 ;
        RECT 285.300 2716.980 285.560 2717.240 ;
        RECT 761.400 2717.320 761.660 2717.580 ;
        RECT 802.800 2717.320 803.060 2717.580 ;
        RECT 806.940 2717.320 807.200 2717.580 ;
        RECT 968.860 2717.320 969.120 2717.580 ;
        RECT 1045.220 2717.320 1045.480 2717.580 ;
        RECT 1048.440 2717.320 1048.700 2717.580 ;
        RECT 1124.340 2717.320 1124.600 2717.580 ;
        RECT 1151.940 2717.320 1152.200 2717.580 ;
        RECT 1311.100 2717.320 1311.360 2717.580 ;
        RECT 285.760 2716.640 286.020 2716.900 ;
        RECT 771.980 2716.980 772.240 2717.240 ;
        RECT 979.440 2716.980 979.700 2717.240 ;
        RECT 1052.120 2716.980 1052.380 2717.240 ;
        RECT 1054.880 2716.980 1055.140 2717.240 ;
        RECT 1134.920 2716.980 1135.180 2717.240 ;
        RECT 1165.280 2716.980 1165.540 2717.240 ;
        RECT 1332.260 2716.980 1332.520 2717.240 ;
        RECT 286.220 2716.300 286.480 2716.560 ;
        RECT 782.100 2716.640 782.360 2716.900 ;
        RECT 948.160 2716.640 948.420 2716.900 ;
        RECT 1038.320 2716.640 1038.580 2716.900 ;
        RECT 1062.240 2716.640 1062.500 2716.900 ;
        RECT 1155.620 2716.640 1155.880 2716.900 ;
        RECT 1165.740 2716.640 1166.000 2716.900 ;
        RECT 1342.380 2716.640 1342.640 2716.900 ;
        RECT 325.780 2716.300 326.040 2716.560 ;
        RECT 330.840 2716.300 331.100 2716.560 ;
        RECT 367.180 2716.300 367.440 2716.560 ;
        RECT 372.240 2716.300 372.500 2716.560 ;
        RECT 387.880 2716.300 388.140 2716.560 ;
        RECT 396.620 2716.300 396.880 2716.560 ;
        RECT 398.460 2716.300 398.720 2716.560 ;
        RECT 403.520 2716.300 403.780 2716.560 ;
        RECT 403.980 2716.300 404.240 2716.560 ;
        RECT 844.200 2716.300 844.460 2716.560 ;
        RECT 958.740 2716.300 959.000 2716.560 ;
        RECT 1046.140 2716.300 1046.400 2716.560 ;
        RECT 1055.340 2716.300 1055.600 2716.560 ;
        RECT 1145.500 2716.300 1145.760 2716.560 ;
        RECT 1172.640 2716.300 1172.900 2716.560 ;
        RECT 1352.960 2716.300 1353.220 2716.560 ;
        RECT 350.620 2715.960 350.880 2716.220 ;
        RECT 854.780 2715.960 855.040 2716.220 ;
        RECT 937.580 2715.960 937.840 2716.220 ;
        RECT 1031.420 2715.960 1031.680 2716.220 ;
        RECT 1069.140 2715.960 1069.400 2716.220 ;
        RECT 1166.200 2715.960 1166.460 2716.220 ;
        RECT 1179.540 2715.960 1179.800 2716.220 ;
        RECT 1363.080 2715.960 1363.340 2716.220 ;
        RECT 351.080 2715.620 351.340 2715.880 ;
        RECT 865.360 2715.620 865.620 2715.880 ;
        RECT 927.460 2715.620 927.720 2715.880 ;
        RECT 1024.520 2715.620 1024.780 2715.880 ;
        RECT 1082.940 2715.620 1083.200 2715.880 ;
        RECT 1186.900 2715.620 1187.160 2715.880 ;
        RECT 1193.340 2715.620 1193.600 2715.880 ;
        RECT 1383.780 2715.620 1384.040 2715.880 ;
        RECT 357.980 2715.280 358.240 2715.540 ;
        RECT 875.480 2715.280 875.740 2715.540 ;
        RECT 916.880 2715.280 917.140 2715.540 ;
        RECT 1017.620 2715.280 1017.880 2715.540 ;
        RECT 1076.040 2715.280 1076.300 2715.540 ;
        RECT 1176.320 2715.280 1176.580 2715.540 ;
        RECT 1186.440 2715.280 1186.700 2715.540 ;
        RECT 1373.660 2715.280 1373.920 2715.540 ;
        RECT 283.460 2714.940 283.720 2715.200 ;
        RECT 896.180 2714.940 896.440 2715.200 ;
        RECT 906.760 2714.940 907.020 2715.200 ;
        RECT 1010.720 2714.940 1010.980 2715.200 ;
        RECT 1013.940 2714.940 1014.200 2715.200 ;
        RECT 1072.820 2714.940 1073.080 2715.200 ;
        RECT 1089.840 2714.940 1090.100 2715.200 ;
        RECT 1197.020 2714.940 1197.280 2715.200 ;
        RECT 1200.240 2714.940 1200.500 2715.200 ;
        RECT 1394.360 2714.940 1394.620 2715.200 ;
        RECT 337.740 2714.600 338.000 2714.860 ;
        RECT 720.000 2714.600 720.260 2714.860 ;
        RECT 1020.840 2714.600 1021.100 2714.860 ;
        RECT 1082.940 2714.600 1083.200 2714.860 ;
        RECT 1131.240 2714.600 1131.500 2714.860 ;
        RECT 1280.280 2714.600 1280.540 2714.860 ;
        RECT 344.640 2714.260 344.900 2714.520 ;
        RECT 403.980 2714.260 404.240 2714.520 ;
        RECT 455.040 2714.260 455.300 2714.520 ;
        RECT 460.560 2714.260 460.820 2714.520 ;
        RECT 461.940 2714.260 462.200 2714.520 ;
        RECT 470.680 2714.260 470.940 2714.520 ;
        RECT 503.340 2714.260 503.600 2714.520 ;
        RECT 543.360 2714.260 543.620 2714.520 ;
        RECT 544.740 2714.260 545.000 2714.520 ;
        RECT 616.040 2714.260 616.300 2714.520 ;
        RECT 636.740 2714.260 637.000 2714.520 ;
        RECT 641.340 2714.260 641.600 2714.520 ;
        RECT 647.320 2714.260 647.580 2714.520 ;
        RECT 942.180 2714.260 942.440 2714.520 ;
        RECT 1130.780 2714.260 1131.040 2714.520 ;
        RECT 1269.700 2714.260 1269.960 2714.520 ;
        RECT 468.380 2713.920 468.640 2714.180 ;
        RECT 481.260 2713.920 481.520 2714.180 ;
        RECT 496.440 2713.920 496.700 2714.180 ;
        RECT 533.240 2713.920 533.500 2714.180 ;
        RECT 551.640 2713.920 551.900 2714.180 ;
        RECT 626.620 2713.920 626.880 2714.180 ;
        RECT 657.440 2713.920 657.700 2714.180 ;
        RECT 941.720 2713.920 941.980 2714.180 ;
        RECT 1117.440 2713.920 1117.700 2714.180 ;
        RECT 1249.000 2713.920 1249.260 2714.180 ;
        RECT 468.840 2713.580 469.100 2713.840 ;
        RECT 491.840 2713.580 492.100 2713.840 ;
        RECT 537.840 2713.580 538.100 2713.840 ;
        RECT 605.920 2713.580 606.180 2713.840 ;
        RECT 699.300 2713.580 699.560 2713.840 ;
        RECT 703.440 2713.580 703.700 2713.840 ;
        RECT 703.900 2713.580 704.160 2713.840 ;
        RECT 796.820 2713.580 797.080 2713.840 ;
        RECT 1123.420 2713.580 1123.680 2713.840 ;
        RECT 1259.580 2713.580 1259.840 2713.840 ;
        RECT 346.480 2713.240 346.740 2713.500 ;
        RECT 351.540 2713.240 351.800 2713.500 ;
        RECT 482.640 2713.240 482.900 2713.500 ;
        RECT 512.540 2713.240 512.800 2713.500 ;
        RECT 419.160 2712.900 419.420 2713.160 ;
        RECT 428.360 2712.900 428.620 2713.160 ;
        RECT 489.540 2712.900 489.800 2713.160 ;
        RECT 522.660 2713.240 522.920 2713.500 ;
        RECT 530.940 2713.240 531.200 2713.500 ;
        RECT 595.340 2713.240 595.600 2713.500 ;
        RECT 678.600 2713.240 678.860 2713.500 ;
        RECT 803.720 2713.240 803.980 2713.500 ;
        RECT 1102.720 2713.240 1102.980 2713.500 ;
        RECT 1228.300 2713.240 1228.560 2713.500 ;
        RECT 517.140 2712.900 517.400 2713.160 ;
        RECT 574.640 2712.900 574.900 2713.160 ;
        RECT 1110.540 2712.900 1110.800 2713.160 ;
        RECT 1238.880 2712.900 1239.140 2713.160 ;
        RECT 408.580 2712.560 408.840 2712.820 ;
        RECT 421.000 2712.560 421.260 2712.820 ;
        RECT 524.040 2712.560 524.300 2712.820 ;
        RECT 585.220 2712.560 585.480 2712.820 ;
        RECT 668.020 2712.560 668.280 2712.820 ;
        RECT 703.900 2712.560 704.160 2712.820 ;
        RECT 1089.380 2712.560 1089.640 2712.820 ;
        RECT 1207.600 2712.560 1207.860 2712.820 ;
        RECT 475.740 2712.220 476.000 2712.480 ;
        RECT 501.960 2712.220 502.220 2712.480 ;
        RECT 509.780 2712.220 510.040 2712.480 ;
        RECT 564.060 2712.220 564.320 2712.480 ;
        RECT 1096.740 2712.220 1097.000 2712.480 ;
        RECT 1217.720 2712.220 1217.980 2712.480 ;
        RECT 510.240 2711.880 510.500 2712.140 ;
        RECT 553.940 2711.880 554.200 2712.140 ;
        RECT 1055.800 2704.740 1056.060 2705.000 ;
        RECT 1057.180 2704.740 1057.440 2705.000 ;
        RECT 1414.140 2683.660 1414.400 2683.920 ;
        RECT 2335.520 2683.660 2335.780 2683.920 ;
        RECT 1414.140 2676.860 1414.400 2677.120 ;
        RECT 2328.620 2676.860 2328.880 2677.120 ;
        RECT 1414.140 2663.260 1414.400 2663.520 ;
        RECT 2321.720 2663.260 2321.980 2663.520 ;
        RECT 1414.140 2656.120 1414.400 2656.380 ;
        RECT 1783.980 2656.120 1784.240 2656.380 ;
        RECT 1414.140 2642.520 1414.400 2642.780 ;
        RECT 1783.520 2642.520 1783.780 2642.780 ;
        RECT 1414.140 2628.580 1414.400 2628.840 ;
        RECT 1776.620 2628.580 1776.880 2628.840 ;
        RECT 1414.140 2621.780 1414.400 2622.040 ;
        RECT 1770.180 2621.780 1770.440 2622.040 ;
        RECT 1414.140 2607.840 1414.400 2608.100 ;
        RECT 1769.720 2607.840 1769.980 2608.100 ;
        RECT 1414.140 2601.040 1414.400 2601.300 ;
        RECT 1763.740 2601.040 1764.000 2601.300 ;
        RECT 1409.540 2587.100 1409.800 2587.360 ;
        RECT 1763.280 2587.100 1763.540 2587.360 ;
        RECT 1414.140 2573.500 1414.400 2573.760 ;
        RECT 1762.820 2573.500 1763.080 2573.760 ;
        RECT 1410.460 2566.360 1410.720 2566.620 ;
        RECT 2381.060 2566.360 2381.320 2566.620 ;
        RECT 1414.140 2552.760 1414.400 2553.020 ;
        RECT 2373.700 2552.760 2373.960 2553.020 ;
        RECT 1411.380 2545.960 1411.640 2546.220 ;
        RECT 2366.800 2545.960 2367.060 2546.220 ;
        RECT 1409.540 2532.020 1409.800 2532.280 ;
        RECT 2359.900 2532.020 2360.160 2532.280 ;
        RECT 1414.140 2518.080 1414.400 2518.340 ;
        RECT 2353.000 2518.080 2353.260 2518.340 ;
        RECT 1410.460 2511.280 1410.720 2511.540 ;
        RECT 2346.100 2511.280 2346.360 2511.540 ;
        RECT 1414.140 2497.340 1414.400 2497.600 ;
        RECT 2339.660 2497.340 2339.920 2497.600 ;
        RECT 1411.380 2490.540 1411.640 2490.800 ;
        RECT 2339.200 2490.540 2339.460 2490.800 ;
        RECT 1409.540 2476.940 1409.800 2477.200 ;
        RECT 2332.300 2476.940 2332.560 2477.200 ;
        RECT 1412.300 2469.800 1412.560 2470.060 ;
        RECT 2325.400 2469.800 2325.660 2470.060 ;
        RECT 1410.460 2456.200 1410.720 2456.460 ;
        RECT 2318.500 2456.200 2318.760 2456.460 ;
        RECT 1414.140 2442.260 1414.400 2442.520 ;
        RECT 2311.600 2442.260 2311.860 2442.520 ;
        RECT 1414.140 2435.460 1414.400 2435.720 ;
        RECT 2305.160 2435.460 2305.420 2435.720 ;
        RECT 1414.140 2421.520 1414.400 2421.780 ;
        RECT 2304.700 2421.520 2304.960 2421.780 ;
        RECT 1412.300 2414.720 1412.560 2414.980 ;
        RECT 2218.220 2414.720 2218.480 2414.980 ;
        RECT 1410.460 2400.780 1410.720 2401.040 ;
        RECT 1797.780 2400.780 1798.040 2401.040 ;
        RECT 1414.140 2387.180 1414.400 2387.440 ;
        RECT 1797.320 2387.180 1797.580 2387.440 ;
        RECT 1412.760 2380.040 1413.020 2380.300 ;
        RECT 1790.880 2380.040 1791.140 2380.300 ;
        RECT 1410.460 2366.440 1410.720 2366.700 ;
        RECT 1790.420 2366.440 1790.680 2366.700 ;
        RECT 1412.300 2359.640 1412.560 2359.900 ;
        RECT 1749.020 2359.640 1749.280 2359.900 ;
        RECT 1410.460 2345.700 1410.720 2345.960 ;
        RECT 2263.760 2345.700 2264.020 2345.960 ;
        RECT 1414.140 2331.760 1414.400 2332.020 ;
        RECT 1652.420 2331.760 1652.680 2332.020 ;
        RECT 1411.380 2324.960 1411.640 2325.220 ;
        RECT 1646.440 2324.960 1646.700 2325.220 ;
        RECT 1414.140 2311.360 1414.400 2311.620 ;
        RECT 1645.520 2311.360 1645.780 2311.620 ;
        RECT 1412.300 2304.220 1412.560 2304.480 ;
        RECT 1638.620 2304.220 1638.880 2304.480 ;
        RECT 1410.460 2290.620 1410.720 2290.880 ;
        RECT 1631.720 2290.620 1631.980 2290.880 ;
        RECT 1414.140 2276.680 1414.400 2276.940 ;
        RECT 1624.820 2276.680 1625.080 2276.940 ;
        RECT 1414.140 2269.880 1414.400 2270.140 ;
        RECT 1618.380 2269.880 1618.640 2270.140 ;
        RECT 1414.140 2255.940 1414.400 2256.200 ;
        RECT 1611.480 2255.940 1611.740 2256.200 ;
        RECT 1412.300 2249.140 1412.560 2249.400 ;
        RECT 2301.940 2249.140 2302.200 2249.400 ;
        RECT 1414.140 2235.200 1414.400 2235.460 ;
        RECT 2301.020 2235.200 2301.280 2235.460 ;
        RECT 1414.140 2221.600 1414.400 2221.860 ;
        RECT 2294.120 2221.600 2294.380 2221.860 ;
        RECT 1414.140 2214.460 1414.400 2214.720 ;
        RECT 2287.220 2214.460 2287.480 2214.720 ;
        RECT 1414.140 2200.860 1414.400 2201.120 ;
        RECT 2280.320 2200.860 2280.580 2201.120 ;
        RECT 1412.300 2194.060 1412.560 2194.320 ;
        RECT 2273.420 2194.060 2273.680 2194.320 ;
        RECT 1414.140 2180.120 1414.400 2180.380 ;
        RECT 2267.440 2180.120 2267.700 2180.380 ;
        RECT 1414.140 2166.180 1414.400 2166.440 ;
        RECT 2266.520 2166.180 2266.780 2166.440 ;
        RECT 1414.140 2159.380 1414.400 2159.640 ;
        RECT 1459.680 2159.380 1459.940 2159.640 ;
        RECT 1414.140 2145.440 1414.400 2145.700 ;
        RECT 1452.780 2145.440 1453.040 2145.700 ;
        RECT 1414.140 2132.860 1414.400 2133.120 ;
        RECT 1438.520 2132.860 1438.780 2133.120 ;
        RECT 1412.300 2125.040 1412.560 2125.300 ;
        RECT 1431.620 2125.040 1431.880 2125.300 ;
        RECT 1410.460 2111.100 1410.720 2111.360 ;
        RECT 1424.720 2111.100 1424.980 2111.360 ;
        RECT 1408.620 2103.960 1408.880 2104.220 ;
        RECT 1417.820 2103.960 1418.080 2104.220 ;
        RECT 1414.140 2090.360 1414.400 2090.620 ;
        RECT 1473.020 2090.360 1473.280 2090.620 ;
        RECT 1414.140 2083.560 1414.400 2083.820 ;
        RECT 1580.200 2083.560 1580.460 2083.820 ;
        RECT 1409.540 2069.620 1409.800 2069.880 ;
        RECT 1997.420 2069.620 1997.680 2069.880 ;
        RECT 1414.140 2056.020 1414.400 2056.280 ;
        RECT 1990.520 2056.020 1990.780 2056.280 ;
        RECT 1410.460 2048.880 1410.720 2049.140 ;
        RECT 1976.720 2048.880 1976.980 2049.140 ;
        RECT 1414.140 2035.280 1414.400 2035.540 ;
        RECT 1969.820 2035.280 1970.080 2035.540 ;
        RECT 1414.140 2028.140 1414.400 2028.400 ;
        RECT 1962.920 2028.140 1963.180 2028.400 ;
        RECT 1409.540 2014.540 1409.800 2014.800 ;
        RECT 1956.020 2014.540 1956.280 2014.800 ;
        RECT 1414.140 2000.600 1414.400 2000.860 ;
        RECT 1942.220 2000.600 1942.480 2000.860 ;
        RECT 1410.460 1993.800 1410.720 1994.060 ;
        RECT 2228.800 1993.800 2229.060 1994.060 ;
        RECT 1410.460 1979.180 1410.720 1979.440 ;
        RECT 1425.180 1979.180 1425.440 1979.440 ;
        RECT 1411.380 1973.060 1411.640 1973.320 ;
        RECT 2011.220 1973.060 2011.480 1973.320 ;
        RECT 1409.540 1959.460 1409.800 1959.720 ;
        RECT 1601.360 1959.460 1601.620 1959.720 ;
        RECT 1412.300 1948.920 1412.560 1949.180 ;
        RECT 1432.080 1948.920 1432.340 1949.180 ;
        RECT 1410.460 1938.720 1410.720 1938.980 ;
        RECT 1594.000 1938.720 1594.260 1938.980 ;
        RECT 1414.140 1923.080 1414.400 1923.340 ;
        RECT 1438.980 1923.080 1439.240 1923.340 ;
        RECT 1414.140 1917.980 1414.400 1918.240 ;
        RECT 2252.720 1917.980 2252.980 1918.240 ;
        RECT 1414.140 1904.040 1414.400 1904.300 ;
        RECT 2245.820 1904.040 2246.080 1904.300 ;
        RECT 1412.300 1897.240 1412.560 1897.500 ;
        RECT 2238.920 1897.240 2239.180 1897.500 ;
        RECT 1410.460 1883.300 1410.720 1883.560 ;
        RECT 2232.020 1883.300 2232.280 1883.560 ;
        RECT 1414.140 1869.700 1414.400 1869.960 ;
        RECT 1794.100 1869.700 1794.360 1869.960 ;
        RECT 1412.760 1862.560 1413.020 1862.820 ;
        RECT 1787.200 1862.560 1787.460 1862.820 ;
        RECT 1414.140 1848.960 1414.400 1849.220 ;
        RECT 1780.300 1848.960 1780.560 1849.220 ;
        RECT 1412.300 1842.160 1412.560 1842.420 ;
        RECT 1773.860 1842.160 1774.120 1842.420 ;
        RECT 1410.460 1828.220 1410.720 1828.480 ;
        RECT 1766.500 1828.220 1766.760 1828.480 ;
        RECT 1414.140 1814.280 1414.400 1814.540 ;
        RECT 1760.060 1814.280 1760.320 1814.540 ;
        RECT 1412.760 1807.480 1413.020 1807.740 ;
        RECT 1760.980 1807.480 1761.240 1807.740 ;
        RECT 1414.140 1793.540 1414.400 1793.800 ;
        RECT 1752.700 1793.540 1752.960 1793.800 ;
        RECT 1412.300 1786.740 1412.560 1787.000 ;
        RECT 1745.800 1786.740 1746.060 1787.000 ;
        RECT 1410.460 1773.140 1410.720 1773.400 ;
        RECT 1738.900 1773.140 1739.160 1773.400 ;
        RECT 1414.140 1759.200 1414.400 1759.460 ;
        RECT 1732.000 1759.200 1732.260 1759.460 ;
        RECT 1412.760 1752.400 1413.020 1752.660 ;
        RECT 1725.100 1752.400 1725.360 1752.660 ;
        RECT 1414.140 1738.460 1414.400 1738.720 ;
        RECT 1718.660 1738.460 1718.920 1738.720 ;
        RECT 1412.300 1731.660 1412.560 1731.920 ;
        RECT 1718.200 1731.660 1718.460 1731.920 ;
        RECT 1414.140 1717.720 1414.400 1717.980 ;
        RECT 1711.300 1717.720 1711.560 1717.980 ;
        RECT 1414.140 1704.120 1414.400 1704.380 ;
        RECT 1704.400 1704.120 1704.660 1704.380 ;
        RECT 1414.140 1696.980 1414.400 1697.240 ;
        RECT 1697.500 1696.980 1697.760 1697.240 ;
        RECT 1414.140 1683.380 1414.400 1683.640 ;
        RECT 1690.600 1683.380 1690.860 1683.640 ;
        RECT 1411.840 1676.240 1412.100 1676.500 ;
        RECT 1684.160 1676.240 1684.420 1676.500 ;
        RECT 1414.140 1662.640 1414.400 1662.900 ;
        RECT 1683.700 1662.640 1683.960 1662.900 ;
        RECT 1414.140 1648.700 1414.400 1648.960 ;
        RECT 1676.800 1648.700 1677.060 1648.960 ;
        RECT 1414.140 1641.900 1414.400 1642.160 ;
        RECT 1669.900 1641.900 1670.160 1642.160 ;
        RECT 1414.140 1627.960 1414.400 1628.220 ;
        RECT 1663.000 1627.960 1663.260 1628.220 ;
        RECT 1411.840 1621.160 1412.100 1621.420 ;
        RECT 1452.320 1621.160 1452.580 1621.420 ;
        RECT 1414.140 1607.560 1414.400 1607.820 ;
        RECT 1649.660 1607.560 1649.920 1607.820 ;
        RECT 1414.140 1593.620 1414.400 1593.880 ;
        RECT 1459.220 1593.620 1459.480 1593.880 ;
        RECT 1414.140 1586.820 1414.400 1587.080 ;
        RECT 1611.020 1586.820 1611.280 1587.080 ;
        RECT 1414.140 1572.880 1414.400 1573.140 ;
        RECT 1635.400 1572.880 1635.660 1573.140 ;
        RECT 1411.840 1566.080 1412.100 1566.340 ;
        RECT 1628.500 1566.080 1628.760 1566.340 ;
        RECT 1409.540 1552.140 1409.800 1552.400 ;
        RECT 1617.920 1552.140 1618.180 1552.400 ;
        RECT 1414.140 1538.540 1414.400 1538.800 ;
        RECT 1514.420 1538.540 1514.680 1538.800 ;
        RECT 1410.460 1531.400 1410.720 1531.660 ;
        RECT 1607.800 1531.400 1608.060 1531.660 ;
      LAYER met2 ;
        RECT 2539.300 3266.730 2539.560 3267.050 ;
        RECT 2566.900 3266.730 2567.160 3267.050 ;
        RECT 2539.360 3264.525 2539.500 3266.730 ;
        RECT 2566.960 3264.525 2567.100 3266.730 ;
        RECT 646.390 3264.155 646.670 3264.525 ;
        RECT 668.010 3264.155 668.290 3264.525 ;
        RECT 1295.910 3264.155 1296.190 3264.525 ;
        RECT 1318.910 3264.155 1319.190 3264.525 ;
        RECT 1892.530 3264.155 1892.810 3264.525 ;
        RECT 1917.370 3264.155 1917.650 3264.525 ;
        RECT 2539.290 3264.155 2539.570 3264.525 ;
        RECT 2566.890 3264.155 2567.170 3264.525 ;
        RECT 646.460 3263.990 646.600 3264.155 ;
        RECT 668.080 3263.990 668.220 3264.155 ;
        RECT 1295.980 3263.990 1296.120 3264.155 ;
        RECT 1318.980 3263.990 1319.120 3264.155 ;
        RECT 1892.600 3263.990 1892.740 3264.155 ;
        RECT 1917.440 3263.990 1917.580 3264.155 ;
        RECT 2539.360 3263.990 2539.500 3264.155 ;
        RECT 2566.900 3264.010 2567.160 3264.155 ;
        RECT 2594.500 3264.010 2594.760 3264.330 ;
        RECT 646.400 3263.670 646.660 3263.990 ;
        RECT 668.020 3263.670 668.280 3263.990 ;
        RECT 697.920 3263.670 698.180 3263.990 ;
        RECT 1295.920 3263.670 1296.180 3263.990 ;
        RECT 1318.920 3263.670 1319.180 3263.990 ;
        RECT 1345.600 3263.670 1345.860 3263.990 ;
        RECT 1892.540 3263.670 1892.800 3263.990 ;
        RECT 1917.380 3263.670 1917.640 3263.990 ;
        RECT 1946.820 3263.670 1947.080 3263.990 ;
        RECT 2539.300 3263.670 2539.560 3263.990 ;
        RECT 2566.960 3263.855 2567.100 3264.010 ;
        RECT 697.000 3251.770 697.260 3252.090 ;
        RECT 282.990 3230.155 283.270 3230.525 ;
        RECT 283.060 2715.085 283.200 3230.155 ;
        RECT 286.210 3224.715 286.490 3225.085 ;
        RECT 285.750 3215.875 286.030 3216.245 ;
        RECT 285.290 3209.755 285.570 3210.125 ;
        RECT 284.830 3201.595 285.110 3201.965 ;
        RECT 284.370 3196.155 284.650 3196.525 ;
        RECT 283.910 3187.995 284.190 3188.365 ;
        RECT 283.450 2898.315 283.730 2898.685 ;
        RECT 283.520 2715.230 283.660 2898.315 ;
        RECT 283.980 2718.630 284.120 3187.995 ;
        RECT 283.920 2718.310 284.180 2718.630 ;
        RECT 284.440 2718.290 284.580 3196.155 ;
        RECT 284.380 2717.970 284.640 2718.290 ;
        RECT 284.900 2717.610 285.040 3201.595 ;
        RECT 284.840 2717.290 285.100 2717.610 ;
        RECT 285.360 2717.270 285.500 3209.755 ;
        RECT 285.300 2716.950 285.560 2717.270 ;
        RECT 285.820 2716.930 285.960 3215.875 ;
        RECT 285.760 2716.610 286.020 2716.930 ;
        RECT 286.280 2716.590 286.420 3224.715 ;
        RECT 298.170 2892.590 298.450 2892.960 ;
        RECT 298.240 2804.650 298.380 2892.590 ;
      LAYER met2 ;
        RECT 305.000 2805.000 681.480 3251.235 ;
      LAYER met2 ;
        RECT 697.060 3249.565 697.200 3251.770 ;
        RECT 696.990 3249.195 697.270 3249.565 ;
        RECT 697.980 3248.770 698.120 3263.670 ;
        RECT 1331.800 3251.770 1332.060 3252.090 ;
        RECT 697.060 3248.630 698.120 3248.770 ;
        RECT 689.640 3215.390 689.900 3215.710 ;
        RECT 298.180 2804.330 298.440 2804.650 ;
        RECT 337.730 2794.275 338.010 2794.645 ;
        RECT 350.610 2794.275 350.890 2794.645 ;
        RECT 362.110 2794.275 362.390 2794.645 ;
        RECT 368.550 2794.275 368.830 2794.645 ;
        RECT 378.670 2794.275 378.950 2794.645 ;
        RECT 380.050 2794.275 380.330 2794.645 ;
        RECT 386.950 2794.275 387.230 2794.645 ;
        RECT 392.470 2794.275 392.750 2794.645 ;
        RECT 330.840 2788.690 331.100 2789.010 ;
        RECT 317.040 2788.010 317.300 2788.330 ;
        RECT 310.140 2787.670 310.400 2787.990 ;
        RECT 310.200 2717.950 310.340 2787.670 ;
        RECT 305.080 2717.630 305.340 2717.950 ;
        RECT 310.140 2717.630 310.400 2717.950 ;
        RECT 286.220 2716.270 286.480 2716.590 ;
        RECT 282.990 2714.715 283.270 2715.085 ;
        RECT 283.460 2714.910 283.720 2715.230 ;
        RECT 305.140 2700.000 305.280 2717.630 ;
        RECT 317.100 2700.010 317.240 2788.010 ;
        RECT 330.900 2716.590 331.040 2788.690 ;
        RECT 337.280 2788.350 337.540 2788.670 ;
        RECT 325.780 2716.270 326.040 2716.590 ;
        RECT 330.840 2716.270 331.100 2716.590 ;
        RECT 315.330 2700.000 317.240 2700.010 ;
        RECT 305.140 2699.940 305.430 2700.000 ;
        RECT 305.150 2696.000 305.430 2699.940 ;
        RECT 315.270 2699.870 317.240 2700.000 ;
        RECT 325.840 2700.000 325.980 2716.270 ;
        RECT 337.340 2700.010 337.480 2788.350 ;
        RECT 337.800 2714.890 337.940 2794.275 ;
        RECT 344.630 2790.195 344.910 2790.565 ;
        RECT 337.740 2714.570 338.000 2714.890 ;
        RECT 344.700 2714.550 344.840 2790.195 ;
        RECT 350.680 2716.250 350.820 2794.275 ;
        RECT 351.070 2793.595 351.350 2793.965 ;
        RECT 350.620 2715.930 350.880 2716.250 ;
        RECT 351.140 2715.910 351.280 2793.595 ;
        RECT 362.180 2792.750 362.320 2794.275 ;
        RECT 362.120 2792.430 362.380 2792.750 ;
        RECT 368.620 2792.070 368.760 2794.275 ;
        RECT 378.740 2793.090 378.880 2794.275 ;
        RECT 378.680 2792.770 378.940 2793.090 ;
        RECT 380.120 2792.410 380.260 2794.275 ;
        RECT 387.020 2793.430 387.160 2794.275 ;
        RECT 386.960 2793.110 387.220 2793.430 ;
        RECT 380.060 2792.090 380.320 2792.410 ;
        RECT 368.560 2791.750 368.820 2792.070 ;
        RECT 379.140 2791.410 379.400 2791.730 ;
        RECT 386.490 2791.555 386.770 2791.925 ;
        RECT 365.790 2790.875 366.070 2791.245 ;
        RECT 358.440 2789.370 358.700 2789.690 ;
        RECT 351.540 2789.030 351.800 2789.350 ;
        RECT 351.080 2715.590 351.340 2715.910 ;
        RECT 344.640 2714.230 344.900 2714.550 ;
        RECT 351.600 2713.530 351.740 2789.030 ;
        RECT 357.970 2787.475 358.250 2787.845 ;
        RECT 358.040 2715.570 358.180 2787.475 ;
        RECT 357.980 2715.250 358.240 2715.570 ;
        RECT 346.480 2713.210 346.740 2713.530 ;
        RECT 351.540 2713.210 351.800 2713.530 ;
        RECT 336.030 2700.000 337.480 2700.010 ;
        RECT 325.840 2699.940 326.130 2700.000 ;
        RECT 315.270 2696.000 315.550 2699.870 ;
        RECT 325.850 2696.000 326.130 2699.940 ;
        RECT 335.970 2699.870 337.480 2700.000 ;
        RECT 346.540 2700.000 346.680 2713.210 ;
        RECT 358.500 2700.010 358.640 2789.370 ;
        RECT 358.890 2788.155 359.170 2788.525 ;
        RECT 365.860 2788.330 366.000 2790.875 ;
        RECT 372.690 2788.835 372.970 2789.205 ;
        RECT 372.700 2788.690 372.960 2788.835 ;
        RECT 358.960 2787.990 359.100 2788.155 ;
        RECT 365.800 2788.010 366.060 2788.330 ;
        RECT 358.900 2787.670 359.160 2787.990 ;
        RECT 372.240 2787.670 372.500 2787.990 ;
        RECT 372.300 2716.590 372.440 2787.670 ;
        RECT 367.180 2716.270 367.440 2716.590 ;
        RECT 372.240 2716.270 372.500 2716.590 ;
        RECT 356.730 2700.000 358.640 2700.010 ;
        RECT 346.540 2699.940 346.830 2700.000 ;
        RECT 335.970 2696.000 336.250 2699.870 ;
        RECT 346.550 2696.000 346.830 2699.940 ;
        RECT 356.670 2699.870 358.640 2700.000 ;
        RECT 367.240 2700.000 367.380 2716.270 ;
        RECT 379.200 2700.010 379.340 2791.410 ;
        RECT 386.560 2789.350 386.700 2791.555 ;
        RECT 392.540 2791.390 392.680 2794.275 ;
        RECT 396.620 2794.130 396.880 2794.450 ;
        RECT 397.530 2794.275 397.810 2794.645 ;
        RECT 403.510 2794.275 403.790 2794.645 ;
        RECT 407.190 2794.275 407.470 2794.645 ;
        RECT 392.480 2791.070 392.740 2791.390 ;
        RECT 393.390 2789.515 393.670 2789.885 ;
        RECT 393.400 2789.370 393.660 2789.515 ;
        RECT 379.590 2788.835 379.870 2789.205 ;
        RECT 386.500 2789.030 386.760 2789.350 ;
        RECT 379.660 2788.670 379.800 2788.835 ;
        RECT 379.600 2788.350 379.860 2788.670 ;
        RECT 393.390 2788.155 393.670 2788.525 ;
        RECT 393.460 2787.990 393.600 2788.155 ;
        RECT 393.400 2787.670 393.660 2787.990 ;
        RECT 396.680 2716.590 396.820 2794.130 ;
        RECT 397.600 2793.770 397.740 2794.275 ;
        RECT 403.580 2794.110 403.720 2794.275 ;
        RECT 407.200 2794.130 407.460 2794.275 ;
        RECT 407.660 2794.130 407.920 2794.450 ;
        RECT 414.550 2794.275 414.830 2794.645 ;
        RECT 420.990 2794.275 421.270 2794.645 ;
        RECT 426.970 2794.275 427.250 2794.645 ;
        RECT 428.350 2794.275 428.630 2794.645 ;
        RECT 431.110 2794.275 431.390 2794.645 ;
        RECT 397.540 2793.450 397.800 2793.770 ;
        RECT 400.290 2793.595 400.570 2793.965 ;
        RECT 403.520 2793.790 403.780 2794.110 ;
        RECT 400.360 2791.730 400.500 2793.595 ;
        RECT 407.720 2793.430 407.860 2794.130 ;
        RECT 408.110 2793.595 408.390 2793.965 ;
        RECT 408.180 2793.430 408.320 2793.595 ;
        RECT 407.660 2793.110 407.920 2793.430 ;
        RECT 408.120 2793.110 408.380 2793.430 ;
        RECT 408.180 2792.750 408.320 2793.110 ;
        RECT 408.120 2792.430 408.380 2792.750 ;
        RECT 414.620 2792.070 414.760 2794.275 ;
        RECT 400.300 2791.410 400.560 2791.730 ;
        RECT 414.090 2791.555 414.370 2791.925 ;
        RECT 414.560 2791.750 414.820 2792.070 ;
        RECT 414.160 2790.370 414.300 2791.555 ;
        RECT 403.520 2790.050 403.780 2790.370 ;
        RECT 414.100 2790.050 414.360 2790.370 ;
        RECT 403.580 2716.590 403.720 2790.050 ;
        RECT 387.880 2716.270 388.140 2716.590 ;
        RECT 396.620 2716.270 396.880 2716.590 ;
        RECT 398.460 2716.270 398.720 2716.590 ;
        RECT 403.520 2716.270 403.780 2716.590 ;
        RECT 403.980 2716.270 404.240 2716.590 ;
        RECT 377.430 2700.000 379.340 2700.010 ;
        RECT 367.240 2699.940 367.530 2700.000 ;
        RECT 356.670 2696.000 356.950 2699.870 ;
        RECT 367.250 2696.000 367.530 2699.940 ;
        RECT 377.370 2699.870 379.340 2700.000 ;
        RECT 387.940 2700.000 388.080 2716.270 ;
        RECT 398.520 2700.000 398.660 2716.270 ;
        RECT 404.040 2714.550 404.180 2716.270 ;
        RECT 403.980 2714.230 404.240 2714.550 ;
        RECT 419.160 2712.870 419.420 2713.190 ;
        RECT 408.580 2712.530 408.840 2712.850 ;
        RECT 408.640 2700.000 408.780 2712.530 ;
        RECT 419.220 2700.000 419.360 2712.870 ;
        RECT 421.060 2712.850 421.200 2794.275 ;
        RECT 421.450 2793.595 421.730 2793.965 ;
        RECT 421.520 2793.090 421.660 2793.595 ;
        RECT 421.460 2792.770 421.720 2793.090 ;
        RECT 427.040 2792.410 427.180 2794.275 ;
        RECT 426.980 2792.090 427.240 2792.410 ;
        RECT 428.420 2713.190 428.560 2794.275 ;
        RECT 428.360 2712.870 428.620 2713.190 ;
        RECT 421.000 2712.530 421.260 2712.850 ;
        RECT 431.180 2700.010 431.320 2794.275 ;
        RECT 434.340 2794.130 434.600 2794.450 ;
        RECT 438.010 2794.275 438.290 2794.645 ;
        RECT 444.910 2794.275 445.190 2794.645 ;
        RECT 448.130 2794.275 448.410 2794.645 ;
        RECT 450.430 2794.275 450.710 2794.645 ;
        RECT 434.400 2793.965 434.540 2794.130 ;
        RECT 434.330 2793.595 434.610 2793.965 ;
        RECT 434.400 2792.750 434.540 2793.595 ;
        RECT 434.340 2792.430 434.600 2792.750 ;
        RECT 429.410 2700.000 431.320 2700.010 ;
        RECT 387.940 2699.940 388.230 2700.000 ;
        RECT 398.520 2699.940 398.810 2700.000 ;
        RECT 408.640 2699.940 408.930 2700.000 ;
        RECT 419.220 2699.940 419.510 2700.000 ;
        RECT 377.370 2696.000 377.650 2699.870 ;
        RECT 387.950 2696.000 388.230 2699.940 ;
        RECT 398.530 2696.000 398.810 2699.940 ;
        RECT 408.650 2696.000 408.930 2699.940 ;
        RECT 419.230 2696.000 419.510 2699.940 ;
        RECT 429.350 2699.870 431.320 2700.000 ;
        RECT 438.080 2700.010 438.220 2794.275 ;
        RECT 439.400 2793.965 439.660 2794.110 ;
        RECT 439.390 2793.595 439.670 2793.965 ;
        RECT 444.980 2793.770 445.120 2794.275 ;
        RECT 439.460 2791.390 439.600 2793.595 ;
        RECT 444.920 2793.450 445.180 2793.770 ;
        RECT 444.980 2791.730 445.120 2793.450 ;
        RECT 444.920 2791.410 445.180 2791.730 ;
        RECT 439.400 2791.070 439.660 2791.390 ;
        RECT 448.200 2712.250 448.340 2794.275 ;
        RECT 450.440 2794.130 450.700 2794.275 ;
        RECT 455.040 2794.130 455.300 2794.450 ;
        RECT 456.870 2794.275 457.150 2794.645 ;
        RECT 462.390 2794.275 462.670 2794.645 ;
        RECT 467.910 2794.275 468.190 2794.645 ;
        RECT 472.970 2794.275 473.250 2794.645 ;
        RECT 476.650 2794.275 476.930 2794.645 ;
        RECT 483.090 2794.275 483.370 2794.645 ;
        RECT 491.370 2794.275 491.650 2794.645 ;
        RECT 497.810 2794.275 498.090 2794.645 ;
        RECT 503.330 2794.275 503.610 2794.645 ;
        RECT 509.770 2794.275 510.050 2794.645 ;
        RECT 513.450 2794.275 513.730 2794.645 ;
        RECT 517.130 2794.275 517.410 2794.645 ;
        RECT 519.890 2794.275 520.170 2794.645 ;
        RECT 524.030 2794.275 524.310 2794.645 ;
        RECT 526.790 2794.275 527.070 2794.645 ;
        RECT 530.930 2794.275 531.210 2794.645 ;
        RECT 537.830 2794.275 538.110 2794.645 ;
        RECT 539.210 2794.275 539.490 2794.645 ;
        RECT 544.730 2794.275 545.010 2794.645 ;
        RECT 551.630 2794.275 551.910 2794.645 ;
        RECT 455.100 2791.390 455.240 2794.130 ;
        RECT 456.940 2793.430 457.080 2794.275 ;
        RECT 456.880 2793.110 457.140 2793.430 ;
        RECT 462.460 2792.070 462.600 2794.275 ;
        RECT 467.980 2793.090 468.120 2794.275 ;
        RECT 467.920 2792.770 468.180 2793.090 ;
        RECT 462.400 2791.750 462.660 2792.070 ;
        RECT 455.040 2791.070 455.300 2791.390 ;
        RECT 467.980 2789.350 468.120 2792.770 ;
        RECT 473.040 2792.410 473.180 2794.275 ;
        RECT 476.720 2793.430 476.860 2794.275 ;
        RECT 483.160 2794.110 483.300 2794.275 ;
        RECT 483.100 2793.790 483.360 2794.110 ;
        RECT 476.660 2793.110 476.920 2793.430 ;
        RECT 476.720 2792.750 476.860 2793.110 ;
        RECT 483.160 2792.750 483.300 2793.790 ;
        RECT 476.660 2792.430 476.920 2792.750 ;
        RECT 483.100 2792.430 483.360 2792.750 ;
        RECT 472.980 2792.090 473.240 2792.410 ;
        RECT 491.440 2791.730 491.580 2794.275 ;
        RECT 491.380 2791.410 491.640 2791.730 ;
        RECT 497.880 2791.390 498.020 2794.275 ;
        RECT 501.490 2793.595 501.770 2793.965 ;
        RECT 501.500 2793.450 501.760 2793.595 ;
        RECT 497.820 2791.070 498.080 2791.390 ;
        RECT 501.560 2790.030 501.700 2793.450 ;
        RECT 501.500 2789.710 501.760 2790.030 ;
        RECT 467.920 2789.030 468.180 2789.350 ;
        RECT 468.370 2788.155 468.650 2788.525 ;
        RECT 455.030 2787.475 455.310 2787.845 ;
        RECT 461.930 2787.475 462.210 2787.845 ;
        RECT 455.100 2714.550 455.240 2787.475 ;
        RECT 462.000 2714.550 462.140 2787.475 ;
        RECT 455.040 2714.230 455.300 2714.550 ;
        RECT 460.560 2714.230 460.820 2714.550 ;
        RECT 461.940 2714.230 462.200 2714.550 ;
        RECT 448.200 2712.110 448.800 2712.250 ;
        RECT 448.660 2700.010 448.800 2712.110 ;
        RECT 438.080 2700.000 439.990 2700.010 ;
        RECT 448.660 2700.000 450.110 2700.010 ;
        RECT 460.620 2700.000 460.760 2714.230 ;
        RECT 468.440 2714.210 468.580 2788.155 ;
        RECT 468.830 2787.475 469.110 2787.845 ;
        RECT 475.730 2787.475 476.010 2787.845 ;
        RECT 482.630 2787.475 482.910 2787.845 ;
        RECT 489.530 2787.475 489.810 2787.845 ;
        RECT 496.430 2787.475 496.710 2787.845 ;
        RECT 468.380 2713.890 468.640 2714.210 ;
        RECT 468.900 2713.870 469.040 2787.475 ;
        RECT 470.680 2714.230 470.940 2714.550 ;
        RECT 468.840 2713.550 469.100 2713.870 ;
        RECT 470.740 2700.000 470.880 2714.230 ;
        RECT 475.800 2712.510 475.940 2787.475 ;
        RECT 481.260 2713.890 481.520 2714.210 ;
        RECT 475.740 2712.190 476.000 2712.510 ;
        RECT 481.320 2700.000 481.460 2713.890 ;
        RECT 482.700 2713.530 482.840 2787.475 ;
        RECT 482.640 2713.210 482.900 2713.530 ;
        RECT 489.600 2713.190 489.740 2787.475 ;
        RECT 496.500 2714.210 496.640 2787.475 ;
        RECT 503.400 2714.550 503.540 2794.275 ;
        RECT 509.310 2792.915 509.590 2793.285 ;
        RECT 503.800 2791.750 504.060 2792.070 ;
        RECT 503.860 2790.370 504.000 2791.750 ;
        RECT 509.380 2790.370 509.520 2792.915 ;
        RECT 503.800 2790.050 504.060 2790.370 ;
        RECT 509.320 2790.050 509.580 2790.370 ;
        RECT 503.340 2714.230 503.600 2714.550 ;
        RECT 496.440 2713.890 496.700 2714.210 ;
        RECT 491.840 2713.550 492.100 2713.870 ;
        RECT 489.540 2712.870 489.800 2713.190 ;
        RECT 491.900 2700.000 492.040 2713.550 ;
        RECT 509.840 2712.510 509.980 2794.275 ;
        RECT 510.230 2793.595 510.510 2793.965 ;
        RECT 501.960 2712.190 502.220 2712.510 ;
        RECT 509.780 2712.190 510.040 2712.510 ;
        RECT 502.020 2700.000 502.160 2712.190 ;
        RECT 510.300 2712.170 510.440 2793.595 ;
        RECT 513.520 2789.350 513.660 2794.275 ;
        RECT 513.460 2789.030 513.720 2789.350 ;
        RECT 512.540 2713.210 512.800 2713.530 ;
        RECT 510.240 2711.850 510.500 2712.170 ;
        RECT 512.600 2700.000 512.740 2713.210 ;
        RECT 517.200 2713.190 517.340 2794.275 ;
        RECT 519.960 2792.410 520.100 2794.275 ;
        RECT 519.900 2792.090 520.160 2792.410 ;
        RECT 523.580 2792.090 523.840 2792.410 ;
        RECT 523.640 2788.330 523.780 2792.090 ;
        RECT 523.580 2788.010 523.840 2788.330 ;
        RECT 522.660 2713.210 522.920 2713.530 ;
        RECT 517.140 2712.870 517.400 2713.190 ;
        RECT 522.720 2700.000 522.860 2713.210 ;
        RECT 524.100 2712.850 524.240 2794.275 ;
        RECT 526.860 2793.430 527.000 2794.275 ;
        RECT 526.800 2793.110 527.060 2793.430 ;
        RECT 530.480 2793.110 530.740 2793.430 ;
        RECT 530.540 2789.010 530.680 2793.110 ;
        RECT 530.480 2788.690 530.740 2789.010 ;
        RECT 531.000 2713.530 531.140 2794.275 ;
        RECT 531.390 2793.595 531.670 2793.965 ;
        RECT 531.460 2792.750 531.600 2793.595 ;
        RECT 531.400 2792.430 531.660 2792.750 ;
        RECT 537.380 2792.430 537.640 2792.750 ;
        RECT 537.440 2788.670 537.580 2792.430 ;
        RECT 537.380 2788.350 537.640 2788.670 ;
        RECT 533.240 2713.890 533.500 2714.210 ;
        RECT 530.940 2713.210 531.200 2713.530 ;
        RECT 524.040 2712.530 524.300 2712.850 ;
        RECT 533.300 2700.000 533.440 2713.890 ;
        RECT 537.900 2713.870 538.040 2794.275 ;
        RECT 539.280 2792.750 539.420 2794.275 ;
        RECT 542.890 2793.595 543.170 2793.965 ;
        RECT 542.960 2793.090 543.100 2793.595 ;
        RECT 542.900 2792.770 543.160 2793.090 ;
        RECT 539.220 2792.430 539.480 2792.750 ;
        RECT 539.280 2791.730 539.420 2792.430 ;
        RECT 539.220 2791.410 539.480 2791.730 ;
        RECT 542.960 2791.390 543.100 2792.770 ;
        RECT 542.900 2791.070 543.160 2791.390 ;
        RECT 544.800 2714.550 544.940 2794.275 ;
        RECT 543.360 2714.230 543.620 2714.550 ;
        RECT 544.740 2714.230 545.000 2714.550 ;
        RECT 537.840 2713.550 538.100 2713.870 ;
        RECT 543.420 2700.000 543.560 2714.230 ;
        RECT 551.700 2714.210 551.840 2794.275 ;
        RECT 641.340 2790.390 641.600 2790.710 ;
        RECT 641.400 2714.550 641.540 2790.390 ;
        RECT 616.040 2714.230 616.300 2714.550 ;
        RECT 636.740 2714.230 637.000 2714.550 ;
        RECT 641.340 2714.230 641.600 2714.550 ;
        RECT 647.320 2714.230 647.580 2714.550 ;
        RECT 551.640 2713.890 551.900 2714.210 ;
        RECT 605.920 2713.550 606.180 2713.870 ;
        RECT 595.340 2713.210 595.600 2713.530 ;
        RECT 574.640 2712.870 574.900 2713.190 ;
        RECT 564.060 2712.190 564.320 2712.510 ;
        RECT 553.940 2711.850 554.200 2712.170 ;
        RECT 554.000 2700.000 554.140 2711.850 ;
        RECT 564.120 2700.000 564.260 2712.190 ;
        RECT 574.700 2700.000 574.840 2712.870 ;
        RECT 585.220 2712.530 585.480 2712.850 ;
        RECT 585.280 2700.000 585.420 2712.530 ;
        RECT 595.400 2700.000 595.540 2713.210 ;
        RECT 605.980 2700.000 606.120 2713.550 ;
        RECT 616.100 2700.000 616.240 2714.230 ;
        RECT 626.620 2713.890 626.880 2714.210 ;
        RECT 626.680 2700.000 626.820 2713.890 ;
        RECT 636.800 2700.000 636.940 2714.230 ;
        RECT 647.380 2700.000 647.520 2714.230 ;
        RECT 657.440 2713.890 657.700 2714.210 ;
        RECT 657.500 2700.000 657.640 2713.890 ;
        RECT 678.600 2713.210 678.860 2713.530 ;
        RECT 668.020 2712.530 668.280 2712.850 ;
        RECT 668.080 2700.000 668.220 2712.530 ;
        RECT 678.660 2700.000 678.800 2713.210 ;
        RECT 689.700 2700.010 689.840 3215.390 ;
        RECT 697.060 2948.325 697.200 3248.630 ;
        RECT 938.490 3230.835 938.770 3231.205 ;
        RECT 938.560 3229.650 938.700 3230.835 ;
        RECT 710.340 3229.330 710.600 3229.650 ;
        RECT 938.500 3229.330 938.760 3229.650 ;
        RECT 703.440 3222.190 703.700 3222.510 ;
        RECT 696.990 2947.955 697.270 2948.325 ;
        RECT 703.500 2713.870 703.640 3222.190 ;
        RECT 699.300 2713.550 699.560 2713.870 ;
        RECT 703.440 2713.550 703.700 2713.870 ;
        RECT 703.900 2713.550 704.160 2713.870 ;
        RECT 688.850 2700.000 689.840 2700.010 ;
        RECT 438.080 2699.870 440.210 2700.000 ;
        RECT 448.660 2699.870 450.330 2700.000 ;
        RECT 460.620 2699.940 460.910 2700.000 ;
        RECT 470.740 2699.940 471.030 2700.000 ;
        RECT 481.320 2699.940 481.610 2700.000 ;
        RECT 491.900 2699.940 492.190 2700.000 ;
        RECT 502.020 2699.940 502.310 2700.000 ;
        RECT 512.600 2699.940 512.890 2700.000 ;
        RECT 522.720 2699.940 523.010 2700.000 ;
        RECT 533.300 2699.940 533.590 2700.000 ;
        RECT 543.420 2699.940 543.710 2700.000 ;
        RECT 554.000 2699.940 554.290 2700.000 ;
        RECT 564.120 2699.940 564.410 2700.000 ;
        RECT 574.700 2699.940 574.990 2700.000 ;
        RECT 585.280 2699.940 585.570 2700.000 ;
        RECT 595.400 2699.940 595.690 2700.000 ;
        RECT 605.980 2699.940 606.270 2700.000 ;
        RECT 616.100 2699.940 616.390 2700.000 ;
        RECT 626.680 2699.940 626.970 2700.000 ;
        RECT 636.800 2699.940 637.090 2700.000 ;
        RECT 647.380 2699.940 647.670 2700.000 ;
        RECT 657.500 2699.940 657.790 2700.000 ;
        RECT 668.080 2699.940 668.370 2700.000 ;
        RECT 678.660 2699.940 678.950 2700.000 ;
        RECT 429.350 2696.000 429.630 2699.870 ;
        RECT 439.930 2696.000 440.210 2699.870 ;
        RECT 450.050 2696.000 450.330 2699.870 ;
        RECT 460.630 2696.000 460.910 2699.940 ;
        RECT 470.750 2696.000 471.030 2699.940 ;
        RECT 481.330 2696.000 481.610 2699.940 ;
        RECT 491.910 2696.000 492.190 2699.940 ;
        RECT 502.030 2696.000 502.310 2699.940 ;
        RECT 512.610 2696.000 512.890 2699.940 ;
        RECT 522.730 2696.000 523.010 2699.940 ;
        RECT 533.310 2696.000 533.590 2699.940 ;
        RECT 543.430 2696.000 543.710 2699.940 ;
        RECT 554.010 2696.000 554.290 2699.940 ;
        RECT 564.130 2696.000 564.410 2699.940 ;
        RECT 574.710 2696.000 574.990 2699.940 ;
        RECT 585.290 2696.000 585.570 2699.940 ;
        RECT 595.410 2696.000 595.690 2699.940 ;
        RECT 605.990 2696.000 606.270 2699.940 ;
        RECT 616.110 2696.000 616.390 2699.940 ;
        RECT 626.690 2696.000 626.970 2699.940 ;
        RECT 636.810 2696.000 637.090 2699.940 ;
        RECT 647.390 2696.000 647.670 2699.940 ;
        RECT 657.510 2696.000 657.790 2699.940 ;
        RECT 668.090 2696.000 668.370 2699.940 ;
        RECT 678.670 2696.000 678.950 2699.940 ;
        RECT 688.790 2699.870 689.840 2700.000 ;
        RECT 699.360 2700.000 699.500 2713.550 ;
        RECT 703.960 2712.850 704.100 2713.550 ;
        RECT 703.900 2712.530 704.160 2712.850 ;
        RECT 710.400 2700.010 710.540 3229.330 ;
        RECT 938.490 3224.035 938.770 3224.405 ;
        RECT 938.560 3222.510 938.700 3224.035 ;
        RECT 938.500 3222.190 938.760 3222.510 ;
        RECT 938.490 3215.875 938.770 3216.245 ;
        RECT 938.560 3215.710 938.700 3215.875 ;
        RECT 938.500 3215.390 938.760 3215.710 ;
        RECT 938.490 3209.755 938.770 3210.125 ;
        RECT 938.560 3208.910 938.700 3209.755 ;
        RECT 803.720 3208.590 803.980 3208.910 ;
        RECT 938.500 3208.590 938.760 3208.910 ;
        RECT 796.820 3201.450 797.080 3201.770 ;
        RECT 730.120 2718.310 730.380 2718.630 ;
        RECT 720.000 2714.570 720.260 2714.890 ;
        RECT 709.550 2700.000 710.540 2700.010 ;
        RECT 699.360 2699.940 699.650 2700.000 ;
        RECT 688.790 2696.000 689.070 2699.870 ;
        RECT 699.370 2696.000 699.650 2699.940 ;
        RECT 709.490 2699.870 710.540 2700.000 ;
        RECT 720.060 2700.000 720.200 2714.570 ;
        RECT 730.180 2700.000 730.320 2718.310 ;
        RECT 740.700 2717.970 740.960 2718.290 ;
        RECT 740.760 2700.000 740.900 2717.970 ;
        RECT 750.820 2717.630 751.080 2717.950 ;
        RECT 750.880 2700.000 751.020 2717.630 ;
        RECT 761.400 2717.290 761.660 2717.610 ;
        RECT 761.460 2700.000 761.600 2717.290 ;
        RECT 771.980 2716.950 772.240 2717.270 ;
        RECT 772.040 2700.000 772.180 2716.950 ;
        RECT 782.100 2716.610 782.360 2716.930 ;
        RECT 782.160 2700.000 782.300 2716.610 ;
        RECT 792.670 2714.715 792.950 2715.085 ;
        RECT 792.740 2700.000 792.880 2714.715 ;
        RECT 796.880 2713.870 797.020 3201.450 ;
        RECT 802.800 2717.290 803.060 2717.610 ;
        RECT 796.820 2713.550 797.080 2713.870 ;
        RECT 802.860 2700.000 803.000 2717.290 ;
        RECT 803.780 2713.530 803.920 3208.590 ;
        RECT 938.490 3201.595 938.770 3201.965 ;
        RECT 938.500 3201.450 938.760 3201.595 ;
        RECT 941.710 3196.155 941.990 3196.525 ;
        RECT 889.740 2898.170 890.000 2898.490 ;
        RECT 938.490 2898.315 938.770 2898.685 ;
        RECT 938.500 2898.170 938.760 2898.315 ;
        RECT 834.540 2792.090 834.800 2792.410 ;
        RECT 827.640 2791.750 827.900 2792.070 ;
        RECT 813.840 2791.410 814.100 2791.730 ;
        RECT 806.940 2791.070 807.200 2791.390 ;
        RECT 807.000 2717.610 807.140 2791.070 ;
        RECT 806.940 2717.290 807.200 2717.610 ;
        RECT 803.720 2713.210 803.980 2713.530 ;
        RECT 813.900 2700.010 814.040 2791.410 ;
        RECT 827.700 2717.950 827.840 2791.750 ;
        RECT 823.500 2717.630 823.760 2717.950 ;
        RECT 827.640 2717.630 827.900 2717.950 ;
        RECT 813.510 2700.000 814.040 2700.010 ;
        RECT 720.060 2699.940 720.350 2700.000 ;
        RECT 730.180 2699.940 730.470 2700.000 ;
        RECT 740.760 2699.940 741.050 2700.000 ;
        RECT 750.880 2699.940 751.170 2700.000 ;
        RECT 761.460 2699.940 761.750 2700.000 ;
        RECT 772.040 2699.940 772.330 2700.000 ;
        RECT 782.160 2699.940 782.450 2700.000 ;
        RECT 792.740 2699.940 793.030 2700.000 ;
        RECT 802.860 2699.940 803.150 2700.000 ;
        RECT 709.490 2696.000 709.770 2699.870 ;
        RECT 720.070 2696.000 720.350 2699.940 ;
        RECT 730.190 2696.000 730.470 2699.940 ;
        RECT 740.770 2696.000 741.050 2699.940 ;
        RECT 750.890 2696.000 751.170 2699.940 ;
        RECT 761.470 2696.000 761.750 2699.940 ;
        RECT 772.050 2696.000 772.330 2699.940 ;
        RECT 782.170 2696.000 782.450 2699.940 ;
        RECT 792.750 2696.000 793.030 2699.940 ;
        RECT 802.870 2696.000 803.150 2699.940 ;
        RECT 813.450 2699.870 814.040 2700.000 ;
        RECT 823.560 2700.000 823.700 2717.630 ;
        RECT 834.600 2700.010 834.740 2792.090 ;
        RECT 889.800 2717.950 889.940 2898.170 ;
        RECT 886.060 2717.630 886.320 2717.950 ;
        RECT 889.740 2717.630 890.000 2717.950 ;
        RECT 844.200 2716.270 844.460 2716.590 ;
        RECT 834.210 2700.000 834.740 2700.010 ;
        RECT 823.560 2699.940 823.850 2700.000 ;
        RECT 813.450 2696.000 813.730 2699.870 ;
        RECT 823.570 2696.000 823.850 2699.940 ;
        RECT 834.150 2699.870 834.740 2700.000 ;
        RECT 844.260 2700.000 844.400 2716.270 ;
        RECT 854.780 2715.930 855.040 2716.250 ;
        RECT 854.840 2700.000 854.980 2715.930 ;
        RECT 865.360 2715.590 865.620 2715.910 ;
        RECT 865.420 2700.000 865.560 2715.590 ;
        RECT 875.480 2715.250 875.740 2715.570 ;
        RECT 875.540 2700.000 875.680 2715.250 ;
        RECT 886.120 2700.000 886.260 2717.630 ;
        RECT 937.580 2715.930 937.840 2716.250 ;
        RECT 927.460 2715.590 927.720 2715.910 ;
        RECT 916.880 2715.250 917.140 2715.570 ;
        RECT 896.180 2714.910 896.440 2715.230 ;
        RECT 906.760 2714.910 907.020 2715.230 ;
        RECT 896.240 2700.000 896.380 2714.910 ;
        RECT 906.820 2700.000 906.960 2714.910 ;
        RECT 916.940 2700.000 917.080 2715.250 ;
        RECT 927.520 2700.000 927.660 2715.590 ;
        RECT 937.640 2700.000 937.780 2715.930 ;
        RECT 941.780 2714.210 941.920 3196.155 ;
        RECT 942.170 3187.995 942.450 3188.365 ;
        RECT 942.240 2714.550 942.380 3187.995 ;
        RECT 944.930 2891.515 945.210 2891.885 ;
        RECT 945.000 2804.650 945.140 2891.515 ;
      LAYER met2 ;
        RECT 955.000 2805.000 1331.480 3251.235 ;
      LAYER met2 ;
        RECT 1331.860 3250.390 1332.000 3251.770 ;
        RECT 1331.800 3250.070 1332.060 3250.390 ;
        RECT 1331.860 3249.450 1332.000 3250.070 ;
        RECT 1332.250 3249.450 1332.530 3249.565 ;
        RECT 1331.860 3249.310 1332.530 3249.450 ;
        RECT 1332.250 3249.195 1332.530 3249.310 ;
        RECT 1345.660 2946.965 1345.800 3263.670 ;
        RECT 1410.000 3251.770 1410.260 3252.090 ;
        RECT 1945.900 3251.770 1946.160 3252.090 ;
        RECT 1410.060 3250.390 1410.200 3251.770 ;
        RECT 1407.700 3250.070 1407.960 3250.390 ;
        RECT 1410.000 3250.070 1410.260 3250.390 ;
        RECT 1345.590 2946.595 1345.870 2946.965 ;
        RECT 1345.660 2938.805 1345.800 2946.595 ;
        RECT 1345.590 2938.435 1345.870 2938.805 ;
        RECT 1350.190 2904.435 1350.470 2904.805 ;
        RECT 1350.260 2901.550 1350.400 2904.435 ;
        RECT 1350.200 2901.230 1350.460 2901.550 ;
        RECT 944.940 2804.330 945.200 2804.650 ;
        RECT 1055.330 2799.715 1055.610 2800.085 ;
        RECT 1052.110 2799.035 1052.390 2799.405 ;
        RECT 1013.930 2794.275 1014.210 2794.645 ;
        RECT 1020.830 2794.275 1021.110 2794.645 ;
        RECT 1027.730 2794.275 1028.010 2794.645 ;
        RECT 979.890 2793.595 980.170 2793.965 ;
        RECT 1007.490 2793.595 1007.770 2793.965 ;
        RECT 1010.710 2793.595 1010.990 2793.965 ;
        RECT 979.960 2790.710 980.100 2793.595 ;
        RECT 986.790 2792.915 987.070 2793.285 ;
        RECT 986.860 2791.390 987.000 2792.915 ;
        RECT 993.690 2792.235 993.970 2792.605 ;
        RECT 1001.050 2792.235 1001.330 2792.605 ;
        RECT 1007.560 2792.410 1007.700 2793.595 ;
        RECT 993.760 2791.730 993.900 2792.235 ;
        RECT 1001.120 2792.070 1001.260 2792.235 ;
        RECT 1007.500 2792.090 1007.760 2792.410 ;
        RECT 1001.060 2791.750 1001.320 2792.070 ;
        RECT 993.700 2791.410 993.960 2791.730 ;
        RECT 986.800 2791.070 987.060 2791.390 ;
        RECT 979.900 2790.390 980.160 2790.710 ;
        RECT 993.700 2790.050 993.960 2790.370 ;
        RECT 986.800 2789.710 987.060 2790.030 ;
        RECT 968.860 2717.290 969.120 2717.610 ;
        RECT 948.160 2716.610 948.420 2716.930 ;
        RECT 942.180 2714.230 942.440 2714.550 ;
        RECT 941.720 2713.890 941.980 2714.210 ;
        RECT 948.220 2700.000 948.360 2716.610 ;
        RECT 958.740 2716.270 959.000 2716.590 ;
        RECT 958.800 2700.000 958.940 2716.270 ;
        RECT 968.920 2700.000 969.060 2717.290 ;
        RECT 979.440 2716.950 979.700 2717.270 ;
        RECT 979.500 2700.000 979.640 2716.950 ;
        RECT 844.260 2699.940 844.550 2700.000 ;
        RECT 854.840 2699.940 855.130 2700.000 ;
        RECT 865.420 2699.940 865.710 2700.000 ;
        RECT 875.540 2699.940 875.830 2700.000 ;
        RECT 886.120 2699.940 886.410 2700.000 ;
        RECT 896.240 2699.940 896.530 2700.000 ;
        RECT 906.820 2699.940 907.110 2700.000 ;
        RECT 916.940 2699.940 917.230 2700.000 ;
        RECT 927.520 2699.940 927.810 2700.000 ;
        RECT 937.640 2699.940 937.930 2700.000 ;
        RECT 948.220 2699.940 948.510 2700.000 ;
        RECT 958.800 2699.940 959.090 2700.000 ;
        RECT 968.920 2699.940 969.210 2700.000 ;
        RECT 979.500 2699.940 979.790 2700.000 ;
        RECT 834.150 2696.000 834.430 2699.870 ;
        RECT 844.270 2696.000 844.550 2699.940 ;
        RECT 854.850 2696.000 855.130 2699.940 ;
        RECT 865.430 2696.000 865.710 2699.940 ;
        RECT 875.550 2696.000 875.830 2699.940 ;
        RECT 886.130 2696.000 886.410 2699.940 ;
        RECT 896.250 2696.000 896.530 2699.940 ;
        RECT 906.830 2696.000 907.110 2699.940 ;
        RECT 916.950 2696.000 917.230 2699.940 ;
        RECT 927.530 2696.000 927.810 2699.940 ;
        RECT 937.650 2696.000 937.930 2699.940 ;
        RECT 948.230 2696.000 948.510 2699.940 ;
        RECT 958.810 2696.000 959.090 2699.940 ;
        RECT 968.930 2696.000 969.210 2699.940 ;
        RECT 979.510 2696.000 979.790 2699.940 ;
        RECT 986.860 2699.330 987.000 2789.710 ;
        RECT 989.630 2699.330 989.910 2700.000 ;
        RECT 986.860 2699.190 989.910 2699.330 ;
        RECT 993.760 2699.330 993.900 2790.050 ;
        RECT 1010.780 2789.690 1010.920 2793.595 ;
        RECT 1010.720 2789.370 1010.980 2789.690 ;
        RECT 1007.500 2789.030 1007.760 2789.350 ;
        RECT 1000.210 2699.330 1000.490 2700.000 ;
        RECT 993.760 2699.190 1000.490 2699.330 ;
        RECT 1007.560 2699.330 1007.700 2789.030 ;
        RECT 1010.780 2715.230 1010.920 2789.370 ;
        RECT 1014.000 2715.230 1014.140 2794.275 ;
        RECT 1017.610 2792.915 1017.890 2793.285 ;
        RECT 1017.680 2789.350 1017.820 2792.915 ;
        RECT 1017.620 2789.030 1017.880 2789.350 ;
        RECT 1014.400 2788.010 1014.660 2788.330 ;
        RECT 1010.720 2714.910 1010.980 2715.230 ;
        RECT 1013.940 2714.910 1014.200 2715.230 ;
        RECT 1014.460 2700.690 1014.600 2788.010 ;
        RECT 1017.680 2715.570 1017.820 2789.030 ;
        RECT 1017.620 2715.250 1017.880 2715.570 ;
        RECT 1020.900 2714.890 1021.040 2794.275 ;
        RECT 1024.510 2793.595 1024.790 2793.965 ;
        RECT 1024.580 2790.710 1024.720 2793.595 ;
        RECT 1024.520 2790.390 1024.780 2790.710 ;
        RECT 1024.580 2715.910 1024.720 2790.390 ;
        RECT 1027.800 2718.290 1027.940 2794.275 ;
        RECT 1045.210 2792.915 1045.490 2793.285 ;
        RECT 1031.410 2790.195 1031.690 2790.565 ;
        RECT 1031.420 2790.050 1031.680 2790.195 ;
        RECT 1028.200 2788.690 1028.460 2789.010 ;
        RECT 1027.740 2717.970 1028.000 2718.290 ;
        RECT 1024.520 2715.590 1024.780 2715.910 ;
        RECT 1020.840 2714.570 1021.100 2714.890 ;
        RECT 1014.460 2700.550 1019.200 2700.690 ;
        RECT 1019.060 2700.010 1019.200 2700.550 ;
        RECT 1019.060 2700.000 1020.970 2700.010 ;
        RECT 1010.330 2699.330 1010.610 2700.000 ;
        RECT 1019.060 2699.870 1021.190 2700.000 ;
        RECT 1007.560 2699.190 1010.610 2699.330 ;
        RECT 989.630 2696.000 989.910 2699.190 ;
        RECT 1000.210 2696.000 1000.490 2699.190 ;
        RECT 1010.330 2696.000 1010.610 2699.190 ;
        RECT 1020.910 2696.000 1021.190 2699.870 ;
        RECT 1028.260 2699.330 1028.400 2788.690 ;
        RECT 1031.480 2716.250 1031.620 2790.050 ;
        RECT 1038.380 2788.670 1038.520 2788.825 ;
        RECT 1035.100 2788.350 1035.360 2788.670 ;
        RECT 1038.320 2788.525 1038.580 2788.670 ;
        RECT 1034.630 2787.475 1034.910 2787.845 ;
        RECT 1034.700 2718.630 1034.840 2787.475 ;
        RECT 1034.640 2718.310 1034.900 2718.630 ;
        RECT 1031.420 2715.930 1031.680 2716.250 ;
        RECT 1035.160 2700.690 1035.300 2788.350 ;
        RECT 1038.310 2788.155 1038.590 2788.525 ;
        RECT 1045.280 2788.330 1045.420 2792.915 ;
        RECT 1048.900 2792.430 1049.160 2792.750 ;
        RECT 1046.140 2789.710 1046.400 2790.030 ;
        RECT 1046.200 2788.525 1046.340 2789.710 ;
        RECT 1038.380 2716.930 1038.520 2788.155 ;
        RECT 1045.220 2788.010 1045.480 2788.330 ;
        RECT 1046.130 2788.155 1046.410 2788.525 ;
        RECT 1041.530 2787.475 1041.810 2787.845 ;
        RECT 1041.600 2717.950 1041.740 2787.475 ;
        RECT 1041.540 2717.630 1041.800 2717.950 ;
        RECT 1045.280 2717.610 1045.420 2788.010 ;
        RECT 1045.220 2717.290 1045.480 2717.610 ;
        RECT 1038.320 2716.610 1038.580 2716.930 ;
        RECT 1046.200 2716.590 1046.340 2788.155 ;
        RECT 1048.430 2787.475 1048.710 2787.845 ;
        RECT 1048.500 2717.610 1048.640 2787.475 ;
        RECT 1048.440 2717.290 1048.700 2717.610 ;
        RECT 1046.140 2716.270 1046.400 2716.590 ;
        RECT 1035.160 2700.550 1039.440 2700.690 ;
        RECT 1039.300 2700.010 1039.440 2700.550 ;
        RECT 1039.300 2700.000 1041.670 2700.010 ;
        RECT 1031.030 2699.330 1031.310 2700.000 ;
        RECT 1039.300 2699.870 1041.890 2700.000 ;
        RECT 1028.260 2699.190 1031.310 2699.330 ;
        RECT 1031.030 2696.000 1031.310 2699.190 ;
        RECT 1041.610 2696.000 1041.890 2699.870 ;
        RECT 1048.960 2699.330 1049.100 2792.430 ;
        RECT 1052.180 2787.990 1052.320 2799.035 ;
        RECT 1054.870 2788.155 1055.150 2788.525 ;
        RECT 1052.120 2787.670 1052.380 2787.990 ;
        RECT 1052.180 2717.270 1052.320 2787.670 ;
        RECT 1054.940 2717.270 1055.080 2788.155 ;
        RECT 1052.120 2716.950 1052.380 2717.270 ;
        RECT 1054.880 2716.950 1055.140 2717.270 ;
        RECT 1055.400 2716.590 1055.540 2799.715 ;
        RECT 1059.470 2794.275 1059.750 2794.645 ;
        RECT 1065.910 2794.275 1066.190 2794.645 ;
        RECT 1069.590 2794.275 1069.870 2794.645 ;
        RECT 1082.930 2794.275 1083.210 2794.645 ;
        RECT 1087.990 2794.275 1088.270 2794.645 ;
        RECT 1089.370 2794.275 1089.650 2794.645 ;
        RECT 1094.430 2794.275 1094.710 2794.645 ;
        RECT 1096.730 2794.275 1097.010 2794.645 ;
        RECT 1100.410 2794.275 1100.690 2794.645 ;
        RECT 1103.630 2794.275 1103.910 2794.645 ;
        RECT 1105.470 2794.275 1105.750 2794.645 ;
        RECT 1110.530 2794.275 1110.810 2794.645 ;
        RECT 1111.450 2794.275 1111.730 2794.645 ;
        RECT 1117.430 2794.275 1117.710 2794.645 ;
        RECT 1124.330 2794.275 1124.610 2794.645 ;
        RECT 1128.930 2794.275 1129.210 2794.645 ;
        RECT 1131.230 2794.275 1131.510 2794.645 ;
        RECT 1135.830 2794.275 1136.110 2794.645 ;
        RECT 1138.130 2794.275 1138.410 2794.645 ;
        RECT 1145.030 2794.275 1145.310 2794.645 ;
        RECT 1147.330 2794.275 1147.610 2794.645 ;
        RECT 1151.930 2794.275 1152.210 2794.645 ;
        RECT 1158.830 2794.275 1159.110 2794.645 ;
        RECT 1159.750 2794.275 1160.030 2794.645 ;
        RECT 1165.730 2794.275 1166.010 2794.645 ;
        RECT 1172.630 2794.275 1172.910 2794.645 ;
        RECT 1179.530 2794.275 1179.810 2794.645 ;
        RECT 1186.430 2794.275 1186.710 2794.645 ;
        RECT 1200.230 2794.275 1200.510 2794.645 ;
        RECT 1056.720 2792.770 1056.980 2793.090 ;
        RECT 1055.800 2792.430 1056.060 2792.750 ;
        RECT 1055.860 2789.690 1056.000 2792.430 ;
        RECT 1055.800 2789.370 1056.060 2789.690 ;
        RECT 1056.780 2766.650 1056.920 2792.770 ;
        RECT 1059.540 2792.750 1059.680 2794.275 ;
        RECT 1065.980 2793.090 1066.120 2794.275 ;
        RECT 1062.700 2792.770 1062.960 2793.090 ;
        RECT 1065.920 2792.770 1066.180 2793.090 ;
        RECT 1059.480 2792.430 1059.740 2792.750 ;
        RECT 1062.760 2789.350 1062.900 2792.770 ;
        RECT 1069.660 2791.730 1069.800 2794.275 ;
        RECT 1076.490 2793.595 1076.770 2793.965 ;
        RECT 1076.560 2793.430 1076.700 2793.595 ;
        RECT 1076.500 2793.110 1076.760 2793.430 ;
        RECT 1069.600 2791.410 1069.860 2791.730 ;
        RECT 1069.660 2790.710 1069.800 2791.410 ;
        RECT 1069.600 2790.390 1069.860 2790.710 ;
        RECT 1076.560 2790.370 1076.700 2793.110 ;
        RECT 1076.500 2790.050 1076.760 2790.370 ;
        RECT 1062.700 2789.030 1062.960 2789.350 ;
        RECT 1062.230 2787.475 1062.510 2787.845 ;
        RECT 1069.130 2787.475 1069.410 2787.845 ;
        RECT 1076.030 2787.475 1076.310 2787.845 ;
        RECT 1056.320 2766.510 1056.920 2766.650 ;
        RECT 1056.320 2753.165 1056.460 2766.510 ;
        RECT 1056.250 2752.795 1056.530 2753.165 ;
        RECT 1057.170 2752.795 1057.450 2753.165 ;
        RECT 1055.340 2716.270 1055.600 2716.590 ;
        RECT 1057.240 2705.030 1057.380 2752.795 ;
        RECT 1062.300 2716.930 1062.440 2787.475 ;
        RECT 1062.240 2716.610 1062.500 2716.930 ;
        RECT 1069.200 2716.250 1069.340 2787.475 ;
        RECT 1069.140 2715.930 1069.400 2716.250 ;
        RECT 1076.100 2715.570 1076.240 2787.475 ;
        RECT 1083.000 2715.910 1083.140 2794.275 ;
        RECT 1083.850 2793.595 1084.130 2793.965 ;
        RECT 1083.860 2793.450 1084.120 2793.595 ;
        RECT 1083.400 2791.070 1083.660 2791.390 ;
        RECT 1083.460 2790.030 1083.600 2791.070 ;
        RECT 1083.400 2789.710 1083.660 2790.030 ;
        RECT 1083.920 2788.670 1084.060 2793.450 ;
        RECT 1088.060 2791.390 1088.200 2794.275 ;
        RECT 1088.000 2791.070 1088.260 2791.390 ;
        RECT 1083.860 2788.350 1084.120 2788.670 ;
        RECT 1082.940 2715.590 1083.200 2715.910 ;
        RECT 1076.040 2715.250 1076.300 2715.570 ;
        RECT 1072.820 2714.910 1073.080 2715.230 ;
        RECT 1055.800 2704.710 1056.060 2705.030 ;
        RECT 1057.180 2704.710 1057.440 2705.030 ;
        RECT 1055.860 2700.690 1056.000 2704.710 ;
        RECT 1055.860 2700.550 1060.140 2700.690 ;
        RECT 1052.190 2699.330 1052.470 2700.000 ;
        RECT 1048.960 2699.190 1052.470 2699.330 ;
        RECT 1060.000 2699.330 1060.140 2700.550 ;
        RECT 1072.880 2700.000 1073.020 2714.910 ;
        RECT 1082.940 2714.570 1083.200 2714.890 ;
        RECT 1083.000 2700.000 1083.140 2714.570 ;
        RECT 1089.440 2712.850 1089.580 2794.275 ;
        RECT 1089.830 2793.595 1090.110 2793.965 ;
        RECT 1089.900 2715.230 1090.040 2793.595 ;
        RECT 1094.500 2792.070 1094.640 2794.275 ;
        RECT 1090.300 2791.750 1090.560 2792.070 ;
        RECT 1094.440 2791.750 1094.700 2792.070 ;
        RECT 1090.360 2788.330 1090.500 2791.750 ;
        RECT 1090.300 2788.010 1090.560 2788.330 ;
        RECT 1093.520 2717.970 1093.780 2718.290 ;
        RECT 1089.840 2714.910 1090.100 2715.230 ;
        RECT 1089.380 2712.530 1089.640 2712.850 ;
        RECT 1093.580 2700.000 1093.720 2717.970 ;
        RECT 1096.800 2712.510 1096.940 2794.275 ;
        RECT 1100.480 2787.990 1100.620 2794.275 ;
        RECT 1100.420 2787.670 1100.680 2787.990 ;
        RECT 1103.700 2726.530 1103.840 2794.275 ;
        RECT 1105.540 2792.750 1105.680 2794.275 ;
        RECT 1105.480 2792.430 1105.740 2792.750 ;
        RECT 1102.780 2726.390 1103.840 2726.530 ;
        RECT 1102.780 2713.530 1102.920 2726.390 ;
        RECT 1103.640 2718.310 1103.900 2718.630 ;
        RECT 1102.720 2713.210 1102.980 2713.530 ;
        RECT 1096.740 2712.190 1097.000 2712.510 ;
        RECT 1103.700 2700.000 1103.840 2718.310 ;
        RECT 1110.600 2713.190 1110.740 2794.275 ;
        RECT 1111.520 2793.090 1111.660 2794.275 ;
        RECT 1111.460 2792.770 1111.720 2793.090 ;
        RECT 1114.220 2717.630 1114.480 2717.950 ;
        RECT 1110.540 2712.870 1110.800 2713.190 ;
        RECT 1114.280 2700.000 1114.420 2717.630 ;
        RECT 1117.500 2714.210 1117.640 2794.275 ;
        RECT 1117.960 2794.110 1118.100 2794.265 ;
        RECT 1117.900 2793.965 1118.160 2794.110 ;
        RECT 1117.890 2793.595 1118.170 2793.965 ;
        RECT 1122.030 2793.595 1122.310 2793.965 ;
        RECT 1117.960 2791.730 1118.100 2793.595 ;
        RECT 1122.100 2793.430 1122.240 2793.595 ;
        RECT 1122.040 2793.110 1122.300 2793.430 ;
        RECT 1117.900 2791.410 1118.160 2791.730 ;
        RECT 1124.400 2726.530 1124.540 2794.275 ;
        RECT 1129.000 2793.770 1129.140 2794.275 ;
        RECT 1128.940 2793.450 1129.200 2793.770 ;
        RECT 1130.770 2793.595 1131.050 2793.965 ;
        RECT 1129.000 2791.730 1129.140 2793.450 ;
        RECT 1128.940 2791.410 1129.200 2791.730 ;
        RECT 1123.480 2726.390 1124.540 2726.530 ;
        RECT 1117.440 2713.890 1117.700 2714.210 ;
        RECT 1123.480 2713.870 1123.620 2726.390 ;
        RECT 1124.340 2717.290 1124.600 2717.610 ;
        RECT 1123.420 2713.550 1123.680 2713.870 ;
        RECT 1124.400 2700.000 1124.540 2717.290 ;
        RECT 1130.840 2714.550 1130.980 2793.595 ;
        RECT 1131.300 2714.890 1131.440 2794.275 ;
        RECT 1135.900 2793.770 1136.040 2794.275 ;
        RECT 1131.700 2793.450 1131.960 2793.770 ;
        RECT 1135.840 2793.450 1136.100 2793.770 ;
        RECT 1131.760 2791.390 1131.900 2793.450 ;
        RECT 1131.700 2791.070 1131.960 2791.390 ;
        RECT 1138.200 2718.290 1138.340 2794.275 ;
        RECT 1138.590 2793.595 1138.870 2793.965 ;
        RECT 1138.660 2792.070 1138.800 2793.595 ;
        RECT 1138.600 2791.750 1138.860 2792.070 ;
        RECT 1139.060 2791.750 1139.320 2792.070 ;
        RECT 1138.660 2791.390 1138.800 2791.750 ;
        RECT 1138.600 2791.070 1138.860 2791.390 ;
        RECT 1139.120 2787.990 1139.260 2791.750 ;
        RECT 1139.060 2787.670 1139.320 2787.990 ;
        RECT 1145.100 2718.630 1145.240 2794.275 ;
        RECT 1147.400 2792.070 1147.540 2794.275 ;
        RECT 1147.340 2791.750 1147.600 2792.070 ;
        RECT 1145.040 2718.310 1145.300 2718.630 ;
        RECT 1138.140 2717.970 1138.400 2718.290 ;
        RECT 1152.000 2717.610 1152.140 2794.275 ;
        RECT 1152.390 2792.915 1152.670 2793.285 ;
        RECT 1152.460 2792.750 1152.600 2792.915 ;
        RECT 1152.400 2792.430 1152.660 2792.750 ;
        RECT 1158.900 2717.950 1159.040 2794.275 ;
        RECT 1159.820 2794.110 1159.960 2794.275 ;
        RECT 1159.760 2793.790 1160.020 2794.110 ;
        RECT 1165.270 2793.595 1165.550 2793.965 ;
        RECT 1159.290 2792.915 1159.570 2793.285 ;
        RECT 1159.300 2792.770 1159.560 2792.915 ;
        RECT 1158.840 2717.630 1159.100 2717.950 ;
        RECT 1151.940 2717.290 1152.200 2717.610 ;
        RECT 1165.340 2717.270 1165.480 2793.595 ;
        RECT 1134.920 2716.950 1135.180 2717.270 ;
        RECT 1165.280 2716.950 1165.540 2717.270 ;
        RECT 1131.240 2714.570 1131.500 2714.890 ;
        RECT 1130.780 2714.230 1131.040 2714.550 ;
        RECT 1134.980 2700.000 1135.120 2716.950 ;
        RECT 1165.800 2716.930 1165.940 2794.275 ;
        RECT 1166.190 2793.595 1166.470 2793.965 ;
        RECT 1166.260 2793.430 1166.400 2793.595 ;
        RECT 1166.200 2793.110 1166.460 2793.430 ;
        RECT 1155.620 2716.610 1155.880 2716.930 ;
        RECT 1165.740 2716.610 1166.000 2716.930 ;
        RECT 1145.500 2716.270 1145.760 2716.590 ;
        RECT 1145.560 2700.000 1145.700 2716.270 ;
        RECT 1155.680 2700.000 1155.820 2716.610 ;
        RECT 1172.700 2716.590 1172.840 2794.275 ;
        RECT 1173.090 2792.915 1173.370 2793.285 ;
        RECT 1173.160 2791.730 1173.300 2792.915 ;
        RECT 1173.100 2791.410 1173.360 2791.730 ;
        RECT 1172.640 2716.270 1172.900 2716.590 ;
        RECT 1179.600 2716.250 1179.740 2794.275 ;
        RECT 1179.990 2793.595 1180.270 2793.965 ;
        RECT 1180.000 2793.450 1180.260 2793.595 ;
        RECT 1166.200 2715.930 1166.460 2716.250 ;
        RECT 1179.540 2715.930 1179.800 2716.250 ;
        RECT 1166.260 2700.000 1166.400 2715.930 ;
        RECT 1186.500 2715.570 1186.640 2794.275 ;
        RECT 1186.890 2792.235 1187.170 2792.605 ;
        RECT 1193.790 2792.235 1194.070 2792.605 ;
        RECT 1186.960 2791.390 1187.100 2792.235 ;
        RECT 1193.860 2792.070 1194.000 2792.235 ;
        RECT 1193.800 2791.750 1194.060 2792.070 ;
        RECT 1186.900 2791.070 1187.160 2791.390 ;
        RECT 1193.330 2790.195 1193.610 2790.565 ;
        RECT 1193.400 2715.910 1193.540 2790.195 ;
        RECT 1186.900 2715.590 1187.160 2715.910 ;
        RECT 1193.340 2715.590 1193.600 2715.910 ;
        RECT 1176.320 2715.250 1176.580 2715.570 ;
        RECT 1186.440 2715.250 1186.700 2715.570 ;
        RECT 1176.380 2700.000 1176.520 2715.250 ;
        RECT 1186.960 2700.000 1187.100 2715.590 ;
        RECT 1200.300 2715.230 1200.440 2794.275 ;
        RECT 1300.980 2718.310 1301.240 2718.630 ;
        RECT 1290.400 2717.970 1290.660 2718.290 ;
        RECT 1197.020 2714.910 1197.280 2715.230 ;
        RECT 1200.240 2714.910 1200.500 2715.230 ;
        RECT 1197.080 2700.000 1197.220 2714.910 ;
        RECT 1280.280 2714.570 1280.540 2714.890 ;
        RECT 1269.700 2714.230 1269.960 2714.550 ;
        RECT 1249.000 2713.890 1249.260 2714.210 ;
        RECT 1228.300 2713.210 1228.560 2713.530 ;
        RECT 1207.600 2712.530 1207.860 2712.850 ;
        RECT 1207.660 2700.000 1207.800 2712.530 ;
        RECT 1217.720 2712.190 1217.980 2712.510 ;
        RECT 1217.780 2700.000 1217.920 2712.190 ;
        RECT 1228.360 2700.000 1228.500 2713.210 ;
        RECT 1238.880 2712.870 1239.140 2713.190 ;
        RECT 1238.940 2700.000 1239.080 2712.870 ;
        RECT 1249.060 2700.000 1249.200 2713.890 ;
        RECT 1259.580 2713.550 1259.840 2713.870 ;
        RECT 1259.640 2700.000 1259.780 2713.550 ;
        RECT 1269.760 2700.000 1269.900 2714.230 ;
        RECT 1280.340 2700.000 1280.480 2714.570 ;
        RECT 1290.460 2700.000 1290.600 2717.970 ;
        RECT 1301.040 2700.000 1301.180 2718.310 ;
        RECT 1321.680 2717.630 1321.940 2717.950 ;
        RECT 1311.100 2717.290 1311.360 2717.610 ;
        RECT 1311.160 2700.000 1311.300 2717.290 ;
        RECT 1321.740 2700.000 1321.880 2717.630 ;
        RECT 1332.260 2716.950 1332.520 2717.270 ;
        RECT 1332.320 2700.000 1332.460 2716.950 ;
        RECT 1342.380 2716.610 1342.640 2716.930 ;
        RECT 1342.440 2700.000 1342.580 2716.610 ;
        RECT 1352.960 2716.270 1353.220 2716.590 ;
        RECT 1353.020 2700.000 1353.160 2716.270 ;
        RECT 1363.080 2715.930 1363.340 2716.250 ;
        RECT 1363.140 2700.000 1363.280 2715.930 ;
        RECT 1383.780 2715.590 1384.040 2715.910 ;
        RECT 1373.660 2715.250 1373.920 2715.570 ;
        RECT 1373.720 2700.000 1373.860 2715.250 ;
        RECT 1383.840 2700.000 1383.980 2715.590 ;
        RECT 1394.360 2714.910 1394.620 2715.230 ;
        RECT 1394.420 2700.000 1394.560 2714.910 ;
        RECT 1062.310 2699.330 1062.590 2700.000 ;
        RECT 1072.880 2699.940 1073.170 2700.000 ;
        RECT 1083.000 2699.940 1083.290 2700.000 ;
        RECT 1093.580 2699.940 1093.870 2700.000 ;
        RECT 1103.700 2699.940 1103.990 2700.000 ;
        RECT 1114.280 2699.940 1114.570 2700.000 ;
        RECT 1124.400 2699.940 1124.690 2700.000 ;
        RECT 1134.980 2699.940 1135.270 2700.000 ;
        RECT 1145.560 2699.940 1145.850 2700.000 ;
        RECT 1155.680 2699.940 1155.970 2700.000 ;
        RECT 1166.260 2699.940 1166.550 2700.000 ;
        RECT 1176.380 2699.940 1176.670 2700.000 ;
        RECT 1186.960 2699.940 1187.250 2700.000 ;
        RECT 1197.080 2699.940 1197.370 2700.000 ;
        RECT 1207.660 2699.940 1207.950 2700.000 ;
        RECT 1217.780 2699.940 1218.070 2700.000 ;
        RECT 1228.360 2699.940 1228.650 2700.000 ;
        RECT 1238.940 2699.940 1239.230 2700.000 ;
        RECT 1249.060 2699.940 1249.350 2700.000 ;
        RECT 1259.640 2699.940 1259.930 2700.000 ;
        RECT 1269.760 2699.940 1270.050 2700.000 ;
        RECT 1280.340 2699.940 1280.630 2700.000 ;
        RECT 1290.460 2699.940 1290.750 2700.000 ;
        RECT 1301.040 2699.940 1301.330 2700.000 ;
        RECT 1311.160 2699.940 1311.450 2700.000 ;
        RECT 1321.740 2699.940 1322.030 2700.000 ;
        RECT 1332.320 2699.940 1332.610 2700.000 ;
        RECT 1342.440 2699.940 1342.730 2700.000 ;
        RECT 1353.020 2699.940 1353.310 2700.000 ;
        RECT 1363.140 2699.940 1363.430 2700.000 ;
        RECT 1373.720 2699.940 1374.010 2700.000 ;
        RECT 1383.840 2699.940 1384.130 2700.000 ;
        RECT 1394.420 2699.940 1394.710 2700.000 ;
        RECT 1060.000 2699.190 1062.590 2699.330 ;
        RECT 1052.190 2696.000 1052.470 2699.190 ;
        RECT 1062.310 2696.000 1062.590 2699.190 ;
        RECT 1072.890 2696.000 1073.170 2699.940 ;
        RECT 1083.010 2696.000 1083.290 2699.940 ;
        RECT 1093.590 2696.000 1093.870 2699.940 ;
        RECT 1103.710 2696.000 1103.990 2699.940 ;
        RECT 1114.290 2696.000 1114.570 2699.940 ;
        RECT 1124.410 2696.000 1124.690 2699.940 ;
        RECT 1134.990 2696.000 1135.270 2699.940 ;
        RECT 1145.570 2696.000 1145.850 2699.940 ;
        RECT 1155.690 2696.000 1155.970 2699.940 ;
        RECT 1166.270 2696.000 1166.550 2699.940 ;
        RECT 1176.390 2696.000 1176.670 2699.940 ;
        RECT 1186.970 2696.000 1187.250 2699.940 ;
        RECT 1197.090 2696.000 1197.370 2699.940 ;
        RECT 1207.670 2696.000 1207.950 2699.940 ;
        RECT 1217.790 2696.000 1218.070 2699.940 ;
        RECT 1228.370 2696.000 1228.650 2699.940 ;
        RECT 1238.950 2696.000 1239.230 2699.940 ;
        RECT 1249.070 2696.000 1249.350 2699.940 ;
        RECT 1259.650 2696.000 1259.930 2699.940 ;
        RECT 1269.770 2696.000 1270.050 2699.940 ;
        RECT 1280.350 2696.000 1280.630 2699.940 ;
        RECT 1290.470 2696.000 1290.750 2699.940 ;
        RECT 1301.050 2696.000 1301.330 2699.940 ;
        RECT 1311.170 2696.000 1311.450 2699.940 ;
        RECT 1321.750 2696.000 1322.030 2699.940 ;
        RECT 1332.330 2696.000 1332.610 2699.940 ;
        RECT 1342.450 2696.000 1342.730 2699.940 ;
        RECT 1353.030 2696.000 1353.310 2699.940 ;
        RECT 1363.150 2696.000 1363.430 2699.940 ;
        RECT 1373.730 2696.000 1374.010 2699.940 ;
        RECT 1383.850 2696.000 1384.130 2699.940 ;
        RECT 1394.430 2696.000 1394.710 2699.940 ;
      LAYER met2 ;
        RECT 304.760 2695.720 304.870 2696.000 ;
        RECT 305.710 2695.720 314.990 2696.000 ;
        RECT 315.830 2695.720 325.570 2696.000 ;
        RECT 326.410 2695.720 335.690 2696.000 ;
        RECT 336.530 2695.720 346.270 2696.000 ;
        RECT 347.110 2695.720 356.390 2696.000 ;
        RECT 357.230 2695.720 366.970 2696.000 ;
        RECT 367.810 2695.720 377.090 2696.000 ;
        RECT 377.930 2695.720 387.670 2696.000 ;
        RECT 388.510 2695.720 398.250 2696.000 ;
        RECT 399.090 2695.720 408.370 2696.000 ;
        RECT 409.210 2695.720 418.950 2696.000 ;
        RECT 419.790 2695.720 429.070 2696.000 ;
        RECT 429.910 2695.720 439.650 2696.000 ;
        RECT 440.490 2695.720 449.770 2696.000 ;
        RECT 450.610 2695.720 460.350 2696.000 ;
        RECT 461.190 2695.720 470.470 2696.000 ;
        RECT 471.310 2695.720 481.050 2696.000 ;
        RECT 481.890 2695.720 491.630 2696.000 ;
        RECT 492.470 2695.720 501.750 2696.000 ;
        RECT 502.590 2695.720 512.330 2696.000 ;
        RECT 513.170 2695.720 522.450 2696.000 ;
        RECT 523.290 2695.720 533.030 2696.000 ;
        RECT 533.870 2695.720 543.150 2696.000 ;
        RECT 543.990 2695.720 553.730 2696.000 ;
        RECT 554.570 2695.720 563.850 2696.000 ;
        RECT 564.690 2695.720 574.430 2696.000 ;
        RECT 575.270 2695.720 585.010 2696.000 ;
        RECT 585.850 2695.720 595.130 2696.000 ;
        RECT 595.970 2695.720 605.710 2696.000 ;
        RECT 606.550 2695.720 615.830 2696.000 ;
        RECT 616.670 2695.720 626.410 2696.000 ;
        RECT 627.250 2695.720 636.530 2696.000 ;
        RECT 637.370 2695.720 647.110 2696.000 ;
        RECT 647.950 2695.720 657.230 2696.000 ;
        RECT 658.070 2695.720 667.810 2696.000 ;
        RECT 668.650 2695.720 678.390 2696.000 ;
        RECT 679.230 2695.720 688.510 2696.000 ;
        RECT 689.350 2695.720 699.090 2696.000 ;
        RECT 699.930 2695.720 709.210 2696.000 ;
        RECT 710.050 2695.720 719.790 2696.000 ;
        RECT 720.630 2695.720 729.910 2696.000 ;
        RECT 730.750 2695.720 740.490 2696.000 ;
        RECT 741.330 2695.720 750.610 2696.000 ;
        RECT 751.450 2695.720 761.190 2696.000 ;
        RECT 762.030 2695.720 771.770 2696.000 ;
        RECT 772.610 2695.720 781.890 2696.000 ;
        RECT 782.730 2695.720 792.470 2696.000 ;
        RECT 793.310 2695.720 802.590 2696.000 ;
        RECT 803.430 2695.720 813.170 2696.000 ;
        RECT 814.010 2695.720 823.290 2696.000 ;
        RECT 824.130 2695.720 833.870 2696.000 ;
        RECT 834.710 2695.720 843.990 2696.000 ;
        RECT 844.830 2695.720 854.570 2696.000 ;
        RECT 855.410 2695.720 865.150 2696.000 ;
        RECT 865.990 2695.720 875.270 2696.000 ;
        RECT 876.110 2695.720 885.850 2696.000 ;
        RECT 886.690 2695.720 895.970 2696.000 ;
        RECT 896.810 2695.720 906.550 2696.000 ;
        RECT 907.390 2695.720 916.670 2696.000 ;
        RECT 917.510 2695.720 927.250 2696.000 ;
        RECT 928.090 2695.720 937.370 2696.000 ;
        RECT 938.210 2695.720 947.950 2696.000 ;
        RECT 948.790 2695.720 958.530 2696.000 ;
        RECT 959.370 2695.720 968.650 2696.000 ;
        RECT 969.490 2695.720 979.230 2696.000 ;
        RECT 980.070 2695.720 989.350 2696.000 ;
        RECT 990.190 2695.720 999.930 2696.000 ;
        RECT 1000.770 2695.720 1010.050 2696.000 ;
        RECT 1010.890 2695.720 1020.630 2696.000 ;
        RECT 1021.470 2695.720 1030.750 2696.000 ;
        RECT 1031.590 2695.720 1041.330 2696.000 ;
        RECT 1042.170 2695.720 1051.910 2696.000 ;
        RECT 1052.750 2695.720 1062.030 2696.000 ;
        RECT 1062.870 2695.720 1072.610 2696.000 ;
        RECT 1073.450 2695.720 1082.730 2696.000 ;
        RECT 1083.570 2695.720 1093.310 2696.000 ;
        RECT 1094.150 2695.720 1103.430 2696.000 ;
        RECT 1104.270 2695.720 1114.010 2696.000 ;
        RECT 1114.850 2695.720 1124.130 2696.000 ;
        RECT 1124.970 2695.720 1134.710 2696.000 ;
        RECT 1135.550 2695.720 1145.290 2696.000 ;
        RECT 1146.130 2695.720 1155.410 2696.000 ;
        RECT 1156.250 2695.720 1165.990 2696.000 ;
        RECT 1166.830 2695.720 1176.110 2696.000 ;
        RECT 1176.950 2695.720 1186.690 2696.000 ;
        RECT 1187.530 2695.720 1196.810 2696.000 ;
        RECT 1197.650 2695.720 1207.390 2696.000 ;
        RECT 1208.230 2695.720 1217.510 2696.000 ;
        RECT 1218.350 2695.720 1228.090 2696.000 ;
        RECT 1228.930 2695.720 1238.670 2696.000 ;
        RECT 1239.510 2695.720 1248.790 2696.000 ;
        RECT 1249.630 2695.720 1259.370 2696.000 ;
        RECT 1260.210 2695.720 1269.490 2696.000 ;
        RECT 1270.330 2695.720 1280.070 2696.000 ;
        RECT 1280.910 2695.720 1290.190 2696.000 ;
        RECT 1291.030 2695.720 1300.770 2696.000 ;
        RECT 1301.610 2695.720 1310.890 2696.000 ;
        RECT 1311.730 2695.720 1321.470 2696.000 ;
        RECT 1322.310 2695.720 1332.050 2696.000 ;
        RECT 1332.890 2695.720 1342.170 2696.000 ;
        RECT 1343.010 2695.720 1352.750 2696.000 ;
        RECT 1353.590 2695.720 1362.870 2696.000 ;
        RECT 1363.710 2695.720 1373.450 2696.000 ;
        RECT 1374.290 2695.720 1383.570 2696.000 ;
        RECT 1384.410 2695.720 1394.150 2696.000 ;
        RECT 1394.990 2695.720 1395.630 2696.000 ;
        RECT 304.760 1504.280 1395.630 2695.720 ;
      LAYER met2 ;
        RECT 1407.760 1516.925 1407.900 3250.070 ;
        RECT 1536.950 3230.155 1537.230 3230.525 ;
        RECT 1537.020 3229.650 1537.160 3230.155 ;
        RECT 1459.680 3229.330 1459.940 3229.650 ;
        RECT 1536.960 3229.330 1537.220 3229.650 ;
        RECT 1452.780 3222.190 1453.040 3222.510 ;
        RECT 1438.520 3215.390 1438.780 3215.710 ;
        RECT 1431.620 3208.590 1431.880 3208.910 ;
        RECT 1424.720 3201.450 1424.980 3201.770 ;
        RECT 1417.820 3194.650 1418.080 3194.970 ;
        RECT 1408.160 2901.230 1408.420 2901.550 ;
        RECT 1407.690 1516.555 1407.970 1516.925 ;
        RECT 1408.220 1506.045 1408.360 2901.230 ;
        RECT 1410.920 2891.030 1411.180 2891.350 ;
        RECT 1410.980 2808.390 1411.120 2891.030 ;
        RECT 1408.620 2808.070 1408.880 2808.390 ;
        RECT 1410.920 2808.070 1411.180 2808.390 ;
        RECT 1408.680 2804.650 1408.820 2808.070 ;
        RECT 1408.620 2804.330 1408.880 2804.650 ;
        RECT 1408.680 2694.685 1408.820 2804.330 ;
        RECT 1408.610 2694.315 1408.890 2694.685 ;
        RECT 1414.140 2683.805 1414.400 2683.950 ;
        RECT 1414.130 2683.435 1414.410 2683.805 ;
        RECT 1414.140 2676.830 1414.400 2677.150 ;
        RECT 1414.200 2672.925 1414.340 2676.830 ;
        RECT 1414.130 2672.555 1414.410 2672.925 ;
        RECT 1414.140 2663.230 1414.400 2663.550 ;
        RECT 1414.200 2662.045 1414.340 2663.230 ;
        RECT 1414.130 2661.675 1414.410 2662.045 ;
        RECT 1414.140 2656.090 1414.400 2656.410 ;
        RECT 1414.200 2651.165 1414.340 2656.090 ;
        RECT 1414.130 2650.795 1414.410 2651.165 ;
        RECT 1414.140 2642.490 1414.400 2642.810 ;
        RECT 1414.200 2639.605 1414.340 2642.490 ;
        RECT 1414.130 2639.235 1414.410 2639.605 ;
        RECT 1414.140 2628.725 1414.400 2628.870 ;
        RECT 1414.130 2628.355 1414.410 2628.725 ;
        RECT 1414.140 2621.750 1414.400 2622.070 ;
        RECT 1414.200 2617.845 1414.340 2621.750 ;
        RECT 1414.130 2617.475 1414.410 2617.845 ;
        RECT 1414.140 2607.810 1414.400 2608.130 ;
        RECT 1414.200 2606.965 1414.340 2607.810 ;
        RECT 1414.130 2606.595 1414.410 2606.965 ;
        RECT 1414.140 2601.010 1414.400 2601.330 ;
        RECT 1414.200 2596.085 1414.340 2601.010 ;
        RECT 1414.130 2595.715 1414.410 2596.085 ;
        RECT 1409.540 2587.070 1409.800 2587.390 ;
        RECT 1409.600 2584.525 1409.740 2587.070 ;
        RECT 1409.530 2584.155 1409.810 2584.525 ;
        RECT 1414.140 2573.645 1414.400 2573.790 ;
        RECT 1414.130 2573.275 1414.410 2573.645 ;
        RECT 1410.460 2566.330 1410.720 2566.650 ;
        RECT 1410.520 2562.765 1410.660 2566.330 ;
        RECT 1410.450 2562.395 1410.730 2562.765 ;
        RECT 1414.140 2552.730 1414.400 2553.050 ;
        RECT 1414.200 2551.885 1414.340 2552.730 ;
        RECT 1414.130 2551.515 1414.410 2551.885 ;
        RECT 1411.380 2545.930 1411.640 2546.250 ;
        RECT 1411.440 2541.005 1411.580 2545.930 ;
        RECT 1411.370 2540.635 1411.650 2541.005 ;
        RECT 1409.540 2531.990 1409.800 2532.310 ;
        RECT 1409.600 2529.445 1409.740 2531.990 ;
        RECT 1409.530 2529.075 1409.810 2529.445 ;
        RECT 1414.130 2518.195 1414.410 2518.565 ;
        RECT 1414.140 2518.050 1414.400 2518.195 ;
        RECT 1410.460 2511.250 1410.720 2511.570 ;
        RECT 1410.520 2507.685 1410.660 2511.250 ;
        RECT 1410.450 2507.315 1410.730 2507.685 ;
        RECT 1414.140 2497.310 1414.400 2497.630 ;
        RECT 1414.200 2496.805 1414.340 2497.310 ;
        RECT 1414.130 2496.435 1414.410 2496.805 ;
        RECT 1411.380 2490.510 1411.640 2490.830 ;
        RECT 1411.440 2485.925 1411.580 2490.510 ;
        RECT 1411.370 2485.555 1411.650 2485.925 ;
        RECT 1409.540 2476.910 1409.800 2477.230 ;
        RECT 1409.600 2474.365 1409.740 2476.910 ;
        RECT 1409.530 2473.995 1409.810 2474.365 ;
        RECT 1412.300 2469.770 1412.560 2470.090 ;
        RECT 1412.360 2463.485 1412.500 2469.770 ;
        RECT 1412.290 2463.115 1412.570 2463.485 ;
        RECT 1410.460 2456.170 1410.720 2456.490 ;
        RECT 1410.520 2452.605 1410.660 2456.170 ;
        RECT 1410.450 2452.235 1410.730 2452.605 ;
        RECT 1414.140 2442.230 1414.400 2442.550 ;
        RECT 1414.200 2441.725 1414.340 2442.230 ;
        RECT 1414.130 2441.355 1414.410 2441.725 ;
        RECT 1414.140 2435.430 1414.400 2435.750 ;
        RECT 1414.200 2430.845 1414.340 2435.430 ;
        RECT 1414.130 2430.475 1414.410 2430.845 ;
        RECT 1414.140 2421.490 1414.400 2421.810 ;
        RECT 1414.200 2419.285 1414.340 2421.490 ;
        RECT 1414.130 2418.915 1414.410 2419.285 ;
        RECT 1412.300 2414.690 1412.560 2415.010 ;
        RECT 1412.360 2408.405 1412.500 2414.690 ;
        RECT 1412.290 2408.035 1412.570 2408.405 ;
        RECT 1410.460 2400.750 1410.720 2401.070 ;
        RECT 1410.520 2397.525 1410.660 2400.750 ;
        RECT 1410.450 2397.155 1410.730 2397.525 ;
        RECT 1414.140 2387.150 1414.400 2387.470 ;
        RECT 1414.200 2386.645 1414.340 2387.150 ;
        RECT 1414.130 2386.275 1414.410 2386.645 ;
        RECT 1412.760 2380.010 1413.020 2380.330 ;
        RECT 1412.820 2375.765 1412.960 2380.010 ;
        RECT 1412.750 2375.395 1413.030 2375.765 ;
        RECT 1410.460 2366.410 1410.720 2366.730 ;
        RECT 1410.520 2364.885 1410.660 2366.410 ;
        RECT 1410.450 2364.515 1410.730 2364.885 ;
        RECT 1412.300 2359.610 1412.560 2359.930 ;
        RECT 1412.360 2353.325 1412.500 2359.610 ;
        RECT 1412.290 2352.955 1412.570 2353.325 ;
        RECT 1410.460 2345.670 1410.720 2345.990 ;
        RECT 1410.520 2342.445 1410.660 2345.670 ;
        RECT 1410.450 2342.075 1410.730 2342.445 ;
        RECT 1414.140 2331.730 1414.400 2332.050 ;
        RECT 1414.200 2331.565 1414.340 2331.730 ;
        RECT 1414.130 2331.195 1414.410 2331.565 ;
        RECT 1411.380 2324.930 1411.640 2325.250 ;
        RECT 1411.440 2320.685 1411.580 2324.930 ;
        RECT 1411.370 2320.315 1411.650 2320.685 ;
        RECT 1414.140 2311.330 1414.400 2311.650 ;
        RECT 1414.200 2309.805 1414.340 2311.330 ;
        RECT 1414.130 2309.435 1414.410 2309.805 ;
        RECT 1412.300 2304.190 1412.560 2304.510 ;
        RECT 1412.360 2298.245 1412.500 2304.190 ;
        RECT 1412.290 2297.875 1412.570 2298.245 ;
        RECT 1410.460 2290.590 1410.720 2290.910 ;
        RECT 1410.520 2287.365 1410.660 2290.590 ;
        RECT 1410.450 2286.995 1410.730 2287.365 ;
        RECT 1414.140 2276.650 1414.400 2276.970 ;
        RECT 1414.200 2276.485 1414.340 2276.650 ;
        RECT 1414.130 2276.115 1414.410 2276.485 ;
        RECT 1414.140 2269.850 1414.400 2270.170 ;
        RECT 1414.200 2265.605 1414.340 2269.850 ;
        RECT 1414.130 2265.235 1414.410 2265.605 ;
        RECT 1414.140 2255.910 1414.400 2256.230 ;
        RECT 1414.200 2254.725 1414.340 2255.910 ;
        RECT 1414.130 2254.355 1414.410 2254.725 ;
        RECT 1412.300 2249.110 1412.560 2249.430 ;
        RECT 1412.360 2243.165 1412.500 2249.110 ;
        RECT 1412.290 2242.795 1412.570 2243.165 ;
        RECT 1414.140 2235.170 1414.400 2235.490 ;
        RECT 1414.200 2232.285 1414.340 2235.170 ;
        RECT 1414.130 2231.915 1414.410 2232.285 ;
        RECT 1414.140 2221.570 1414.400 2221.890 ;
        RECT 1414.200 2221.405 1414.340 2221.570 ;
        RECT 1414.130 2221.035 1414.410 2221.405 ;
        RECT 1414.140 2214.430 1414.400 2214.750 ;
        RECT 1414.200 2210.525 1414.340 2214.430 ;
        RECT 1414.130 2210.155 1414.410 2210.525 ;
        RECT 1414.140 2200.830 1414.400 2201.150 ;
        RECT 1414.200 2199.645 1414.340 2200.830 ;
        RECT 1414.130 2199.275 1414.410 2199.645 ;
        RECT 1412.300 2194.030 1412.560 2194.350 ;
        RECT 1412.360 2188.085 1412.500 2194.030 ;
        RECT 1412.290 2187.715 1412.570 2188.085 ;
        RECT 1414.140 2180.090 1414.400 2180.410 ;
        RECT 1414.200 2177.205 1414.340 2180.090 ;
        RECT 1414.130 2176.835 1414.410 2177.205 ;
        RECT 1414.140 2166.325 1414.400 2166.470 ;
        RECT 1414.130 2165.955 1414.410 2166.325 ;
        RECT 1414.140 2159.350 1414.400 2159.670 ;
        RECT 1414.200 2155.445 1414.340 2159.350 ;
        RECT 1414.130 2155.075 1414.410 2155.445 ;
        RECT 1414.140 2145.410 1414.400 2145.730 ;
        RECT 1414.200 2144.565 1414.340 2145.410 ;
        RECT 1414.130 2144.195 1414.410 2144.565 ;
        RECT 1414.140 2133.005 1414.400 2133.150 ;
        RECT 1414.130 2132.635 1414.410 2133.005 ;
        RECT 1412.300 2125.010 1412.560 2125.330 ;
        RECT 1412.360 2122.125 1412.500 2125.010 ;
        RECT 1412.290 2121.755 1412.570 2122.125 ;
        RECT 1410.460 2111.245 1410.720 2111.390 ;
        RECT 1410.450 2110.875 1410.730 2111.245 ;
        RECT 1417.880 2104.250 1418.020 3194.650 ;
        RECT 1424.780 2111.390 1424.920 3201.450 ;
        RECT 1425.180 2898.170 1425.440 2898.490 ;
        RECT 1424.720 2111.070 1424.980 2111.390 ;
        RECT 1408.620 2103.930 1408.880 2104.250 ;
        RECT 1417.820 2103.930 1418.080 2104.250 ;
        RECT 1408.680 2100.365 1408.820 2103.930 ;
        RECT 1408.610 2099.995 1408.890 2100.365 ;
        RECT 1414.140 2090.330 1414.400 2090.650 ;
        RECT 1414.200 2089.485 1414.340 2090.330 ;
        RECT 1414.130 2089.115 1414.410 2089.485 ;
        RECT 1414.140 2083.530 1414.400 2083.850 ;
        RECT 1414.200 2078.605 1414.340 2083.530 ;
        RECT 1414.130 2078.235 1414.410 2078.605 ;
        RECT 1409.540 2069.590 1409.800 2069.910 ;
        RECT 1409.600 2067.045 1409.740 2069.590 ;
        RECT 1409.530 2066.675 1409.810 2067.045 ;
        RECT 1414.140 2056.165 1414.400 2056.310 ;
        RECT 1414.130 2055.795 1414.410 2056.165 ;
        RECT 1410.460 2048.850 1410.720 2049.170 ;
        RECT 1410.520 2045.285 1410.660 2048.850 ;
        RECT 1410.450 2044.915 1410.730 2045.285 ;
        RECT 1414.140 2035.250 1414.400 2035.570 ;
        RECT 1414.200 2034.405 1414.340 2035.250 ;
        RECT 1414.130 2034.035 1414.410 2034.405 ;
        RECT 1414.140 2028.110 1414.400 2028.430 ;
        RECT 1414.200 2023.525 1414.340 2028.110 ;
        RECT 1414.130 2023.155 1414.410 2023.525 ;
        RECT 1409.540 2014.510 1409.800 2014.830 ;
        RECT 1409.600 2011.965 1409.740 2014.510 ;
        RECT 1409.530 2011.595 1409.810 2011.965 ;
        RECT 1414.130 2000.715 1414.410 2001.085 ;
        RECT 1414.140 2000.570 1414.400 2000.715 ;
        RECT 1410.460 1993.770 1410.720 1994.090 ;
        RECT 1410.520 1990.205 1410.660 1993.770 ;
        RECT 1410.450 1989.835 1410.730 1990.205 ;
        RECT 1425.240 1979.470 1425.380 2898.170 ;
        RECT 1431.680 2125.330 1431.820 3208.590 ;
        RECT 1432.080 2788.350 1432.340 2788.670 ;
        RECT 1431.620 2125.010 1431.880 2125.330 ;
        RECT 1410.460 1979.325 1410.720 1979.470 ;
        RECT 1410.450 1978.955 1410.730 1979.325 ;
        RECT 1425.180 1979.150 1425.440 1979.470 ;
        RECT 1411.380 1973.030 1411.640 1973.350 ;
        RECT 1411.440 1968.445 1411.580 1973.030 ;
        RECT 1411.370 1968.075 1411.650 1968.445 ;
        RECT 1409.540 1959.430 1409.800 1959.750 ;
        RECT 1409.600 1956.885 1409.740 1959.430 ;
        RECT 1409.530 1956.515 1409.810 1956.885 ;
        RECT 1432.140 1949.210 1432.280 2788.350 ;
        RECT 1438.580 2133.150 1438.720 3215.390 ;
        RECT 1452.320 2790.390 1452.580 2790.710 ;
        RECT 1438.980 2788.690 1439.240 2789.010 ;
        RECT 1438.520 2132.830 1438.780 2133.150 ;
        RECT 1412.300 1948.890 1412.560 1949.210 ;
        RECT 1432.080 1948.890 1432.340 1949.210 ;
        RECT 1412.360 1946.005 1412.500 1948.890 ;
        RECT 1412.290 1945.635 1412.570 1946.005 ;
        RECT 1410.460 1938.690 1410.720 1939.010 ;
        RECT 1410.520 1935.125 1410.660 1938.690 ;
        RECT 1410.450 1934.755 1410.730 1935.125 ;
        RECT 1414.130 1923.875 1414.410 1924.245 ;
        RECT 1414.200 1923.370 1414.340 1923.875 ;
        RECT 1439.040 1923.370 1439.180 2788.690 ;
        RECT 1414.140 1923.050 1414.400 1923.370 ;
        RECT 1438.980 1923.050 1439.240 1923.370 ;
        RECT 1414.140 1917.950 1414.400 1918.270 ;
        RECT 1414.200 1913.365 1414.340 1917.950 ;
        RECT 1414.130 1912.995 1414.410 1913.365 ;
        RECT 1414.140 1904.010 1414.400 1904.330 ;
        RECT 1414.200 1901.805 1414.340 1904.010 ;
        RECT 1414.130 1901.435 1414.410 1901.805 ;
        RECT 1412.300 1897.210 1412.560 1897.530 ;
        RECT 1412.360 1890.925 1412.500 1897.210 ;
        RECT 1412.290 1890.555 1412.570 1890.925 ;
        RECT 1410.460 1883.270 1410.720 1883.590 ;
        RECT 1410.520 1880.045 1410.660 1883.270 ;
        RECT 1410.450 1879.675 1410.730 1880.045 ;
        RECT 1414.140 1869.670 1414.400 1869.990 ;
        RECT 1414.200 1869.165 1414.340 1869.670 ;
        RECT 1414.130 1868.795 1414.410 1869.165 ;
        RECT 1412.760 1862.530 1413.020 1862.850 ;
        RECT 1412.820 1858.285 1412.960 1862.530 ;
        RECT 1412.750 1857.915 1413.030 1858.285 ;
        RECT 1414.140 1848.930 1414.400 1849.250 ;
        RECT 1414.200 1846.725 1414.340 1848.930 ;
        RECT 1414.130 1846.355 1414.410 1846.725 ;
        RECT 1412.300 1842.130 1412.560 1842.450 ;
        RECT 1412.360 1835.845 1412.500 1842.130 ;
        RECT 1412.290 1835.475 1412.570 1835.845 ;
        RECT 1410.460 1828.190 1410.720 1828.510 ;
        RECT 1410.520 1824.965 1410.660 1828.190 ;
        RECT 1410.450 1824.595 1410.730 1824.965 ;
        RECT 1414.140 1814.250 1414.400 1814.570 ;
        RECT 1414.200 1814.085 1414.340 1814.250 ;
        RECT 1414.130 1813.715 1414.410 1814.085 ;
        RECT 1412.760 1807.450 1413.020 1807.770 ;
        RECT 1412.820 1803.205 1412.960 1807.450 ;
        RECT 1412.750 1802.835 1413.030 1803.205 ;
        RECT 1414.140 1793.510 1414.400 1793.830 ;
        RECT 1414.200 1792.325 1414.340 1793.510 ;
        RECT 1414.130 1791.955 1414.410 1792.325 ;
        RECT 1412.300 1786.710 1412.560 1787.030 ;
        RECT 1412.360 1780.765 1412.500 1786.710 ;
        RECT 1412.290 1780.395 1412.570 1780.765 ;
        RECT 1410.460 1773.110 1410.720 1773.430 ;
        RECT 1410.520 1769.885 1410.660 1773.110 ;
        RECT 1410.450 1769.515 1410.730 1769.885 ;
        RECT 1414.140 1759.170 1414.400 1759.490 ;
        RECT 1414.200 1759.005 1414.340 1759.170 ;
        RECT 1414.130 1758.635 1414.410 1759.005 ;
        RECT 1412.760 1752.370 1413.020 1752.690 ;
        RECT 1412.820 1748.125 1412.960 1752.370 ;
        RECT 1412.750 1747.755 1413.030 1748.125 ;
        RECT 1414.140 1738.430 1414.400 1738.750 ;
        RECT 1414.200 1737.245 1414.340 1738.430 ;
        RECT 1414.130 1736.875 1414.410 1737.245 ;
        RECT 1412.300 1731.630 1412.560 1731.950 ;
        RECT 1412.360 1725.685 1412.500 1731.630 ;
        RECT 1412.290 1725.315 1412.570 1725.685 ;
        RECT 1414.140 1717.690 1414.400 1718.010 ;
        RECT 1414.200 1714.805 1414.340 1717.690 ;
        RECT 1414.130 1714.435 1414.410 1714.805 ;
        RECT 1414.140 1704.090 1414.400 1704.410 ;
        RECT 1414.200 1703.925 1414.340 1704.090 ;
        RECT 1414.130 1703.555 1414.410 1703.925 ;
        RECT 1414.140 1696.950 1414.400 1697.270 ;
        RECT 1414.200 1693.045 1414.340 1696.950 ;
        RECT 1414.130 1692.675 1414.410 1693.045 ;
        RECT 1414.140 1683.350 1414.400 1683.670 ;
        RECT 1414.200 1682.165 1414.340 1683.350 ;
        RECT 1414.130 1681.795 1414.410 1682.165 ;
        RECT 1411.840 1676.210 1412.100 1676.530 ;
        RECT 1411.900 1670.605 1412.040 1676.210 ;
        RECT 1411.830 1670.235 1412.110 1670.605 ;
        RECT 1414.140 1662.610 1414.400 1662.930 ;
        RECT 1414.200 1659.725 1414.340 1662.610 ;
        RECT 1414.130 1659.355 1414.410 1659.725 ;
        RECT 1414.140 1648.845 1414.400 1648.990 ;
        RECT 1414.130 1648.475 1414.410 1648.845 ;
        RECT 1414.140 1641.870 1414.400 1642.190 ;
        RECT 1414.200 1637.965 1414.340 1641.870 ;
        RECT 1414.130 1637.595 1414.410 1637.965 ;
        RECT 1414.140 1627.930 1414.400 1628.250 ;
        RECT 1414.200 1627.085 1414.340 1627.930 ;
        RECT 1414.130 1626.715 1414.410 1627.085 ;
        RECT 1452.380 1621.450 1452.520 2790.390 ;
        RECT 1452.840 2145.730 1452.980 3222.190 ;
        RECT 1459.220 2791.070 1459.480 2791.390 ;
        RECT 1452.780 2145.410 1453.040 2145.730 ;
        RECT 1411.840 1621.130 1412.100 1621.450 ;
        RECT 1452.320 1621.130 1452.580 1621.450 ;
        RECT 1411.900 1615.525 1412.040 1621.130 ;
        RECT 1411.830 1615.155 1412.110 1615.525 ;
        RECT 1414.140 1607.530 1414.400 1607.850 ;
        RECT 1414.200 1604.645 1414.340 1607.530 ;
        RECT 1414.130 1604.275 1414.410 1604.645 ;
        RECT 1459.280 1593.910 1459.420 2791.070 ;
        RECT 1459.740 2159.670 1459.880 3229.330 ;
        RECT 1535.570 3224.715 1535.850 3225.085 ;
        RECT 1535.640 3222.510 1535.780 3224.715 ;
        RECT 1535.580 3222.190 1535.840 3222.510 ;
        RECT 1535.570 3217.235 1535.850 3217.605 ;
        RECT 1535.640 3215.710 1535.780 3217.235 ;
        RECT 1535.580 3215.390 1535.840 3215.710 ;
        RECT 1538.330 3210.435 1538.610 3210.805 ;
        RECT 1538.400 3208.910 1538.540 3210.435 ;
        RECT 1538.340 3208.590 1538.600 3208.910 ;
        RECT 1538.330 3202.275 1538.610 3202.645 ;
        RECT 1538.400 3201.770 1538.540 3202.275 ;
        RECT 1538.340 3201.450 1538.600 3201.770 ;
        RECT 1533.270 3196.835 1533.550 3197.205 ;
        RECT 1533.340 3194.970 1533.480 3196.835 ;
        RECT 1533.280 3194.650 1533.540 3194.970 ;
        RECT 1497.850 3189.355 1498.130 3189.725 ;
        RECT 1497.920 3188.170 1498.060 3189.355 ;
        RECT 1473.020 3187.850 1473.280 3188.170 ;
        RECT 1497.860 3187.850 1498.120 3188.170 ;
        RECT 1459.680 2159.350 1459.940 2159.670 ;
        RECT 1473.080 2090.650 1473.220 3187.850 ;
        RECT 1534.650 2899.675 1534.930 2900.045 ;
        RECT 1534.720 2898.490 1534.860 2899.675 ;
        RECT 1534.660 2898.170 1534.920 2898.490 ;
        RECT 1531.890 2891.515 1532.170 2891.885 ;
        RECT 1531.960 2891.350 1532.100 2891.515 ;
        RECT 1531.900 2891.090 1532.160 2891.350 ;
        RECT 1531.500 2891.030 1532.160 2891.090 ;
        RECT 1531.500 2890.950 1532.100 2891.030 ;
        RECT 1531.500 2804.650 1531.640 2890.950 ;
        RECT 1531.960 2890.705 1532.100 2890.950 ;
      LAYER met2 ;
        RECT 1555.000 2805.000 1931.480 3251.235 ;
      LAYER met2 ;
        RECT 1945.960 3249.565 1946.100 3251.770 ;
        RECT 1945.890 3249.195 1946.170 3249.565 ;
        RECT 1946.880 3248.770 1947.020 3263.670 ;
        RECT 2582.080 3251.770 2582.340 3252.090 ;
        RECT 1945.960 3248.630 1947.020 3248.770 ;
        RECT 1942.220 3187.850 1942.480 3188.170 ;
        RECT 1531.440 2804.330 1531.700 2804.650 ;
        RECT 1739.810 2796.315 1740.090 2796.685 ;
        RECT 1788.570 2796.315 1788.850 2796.685 ;
        RECT 1580.190 2794.275 1580.470 2794.645 ;
        RECT 1593.990 2794.275 1594.270 2794.645 ;
        RECT 1601.350 2794.275 1601.630 2794.645 ;
        RECT 1607.790 2794.275 1608.070 2794.645 ;
        RECT 1617.910 2794.275 1618.190 2794.645 ;
        RECT 1628.490 2794.275 1628.770 2794.645 ;
        RECT 1635.390 2794.275 1635.670 2794.645 ;
        RECT 1649.650 2794.275 1649.930 2794.645 ;
        RECT 1658.850 2794.275 1659.130 2794.645 ;
        RECT 1662.990 2794.275 1663.270 2794.645 ;
        RECT 1669.890 2794.275 1670.170 2794.645 ;
        RECT 1676.790 2794.275 1677.070 2794.645 ;
        RECT 1514.420 2789.030 1514.680 2789.350 ;
        RECT 1473.020 2090.330 1473.280 2090.650 ;
        RECT 1414.140 1593.765 1414.400 1593.910 ;
        RECT 1414.130 1593.395 1414.410 1593.765 ;
        RECT 1459.220 1593.590 1459.480 1593.910 ;
        RECT 1414.140 1586.790 1414.400 1587.110 ;
        RECT 1414.200 1582.885 1414.340 1586.790 ;
        RECT 1414.130 1582.515 1414.410 1582.885 ;
        RECT 1414.140 1572.850 1414.400 1573.170 ;
        RECT 1414.200 1572.005 1414.340 1572.850 ;
        RECT 1414.130 1571.635 1414.410 1572.005 ;
        RECT 1411.840 1566.050 1412.100 1566.370 ;
        RECT 1411.900 1560.445 1412.040 1566.050 ;
        RECT 1411.830 1560.075 1412.110 1560.445 ;
        RECT 1409.540 1552.110 1409.800 1552.430 ;
        RECT 1409.600 1549.565 1409.740 1552.110 ;
        RECT 1409.530 1549.195 1409.810 1549.565 ;
        RECT 1514.480 1538.830 1514.620 2789.030 ;
        RECT 1580.260 2083.850 1580.400 2794.275 ;
        RECT 1587.090 2792.235 1587.370 2792.605 ;
        RECT 1587.160 2789.010 1587.300 2792.235 ;
        RECT 1587.100 2788.690 1587.360 2789.010 ;
        RECT 1580.200 2083.530 1580.460 2083.850 ;
        RECT 1594.060 1939.010 1594.200 2794.275 ;
        RECT 1600.890 2788.835 1601.170 2789.205 ;
        RECT 1600.960 2788.670 1601.100 2788.835 ;
        RECT 1600.900 2788.350 1601.160 2788.670 ;
        RECT 1601.420 1959.750 1601.560 2794.275 ;
        RECT 1601.360 1959.430 1601.620 1959.750 ;
        RECT 1594.000 1938.690 1594.260 1939.010 ;
        RECT 1414.140 1538.685 1414.400 1538.830 ;
        RECT 1414.130 1538.315 1414.410 1538.685 ;
        RECT 1514.420 1538.510 1514.680 1538.830 ;
        RECT 1607.860 1531.690 1608.000 2794.275 ;
        RECT 1611.470 2793.595 1611.750 2793.965 ;
        RECT 1611.020 2790.050 1611.280 2790.370 ;
        RECT 1611.080 1587.110 1611.220 2790.050 ;
        RECT 1611.540 2789.690 1611.680 2793.595 ;
        RECT 1611.480 2789.370 1611.740 2789.690 ;
        RECT 1614.690 2789.515 1614.970 2789.885 ;
        RECT 1611.540 2256.230 1611.680 2789.370 ;
        RECT 1614.760 2789.350 1614.900 2789.515 ;
        RECT 1614.700 2789.030 1614.960 2789.350 ;
        RECT 1611.480 2255.910 1611.740 2256.230 ;
        RECT 1611.020 1586.790 1611.280 1587.110 ;
        RECT 1617.980 1552.430 1618.120 2794.275 ;
        RECT 1618.370 2792.915 1618.650 2793.285 ;
        RECT 1624.810 2792.915 1625.090 2793.285 ;
        RECT 1618.440 2789.350 1618.580 2792.915 ;
        RECT 1618.380 2789.030 1618.640 2789.350 ;
        RECT 1618.440 2270.170 1618.580 2789.030 ;
        RECT 1624.880 2789.010 1625.020 2792.915 ;
        RECT 1624.820 2788.690 1625.080 2789.010 ;
        RECT 1624.880 2276.970 1625.020 2788.690 ;
        RECT 1624.820 2276.650 1625.080 2276.970 ;
        RECT 1618.380 2269.850 1618.640 2270.170 ;
        RECT 1628.560 1566.370 1628.700 2794.275 ;
        RECT 1631.710 2792.915 1631.990 2793.285 ;
        RECT 1631.780 2788.670 1631.920 2792.915 ;
        RECT 1631.720 2788.350 1631.980 2788.670 ;
        RECT 1631.780 2290.910 1631.920 2788.350 ;
        RECT 1631.720 2290.590 1631.980 2290.910 ;
        RECT 1635.460 1573.170 1635.600 2794.275 ;
        RECT 1638.610 2793.595 1638.890 2793.965 ;
        RECT 1645.510 2793.595 1645.790 2793.965 ;
        RECT 1638.680 2790.030 1638.820 2793.595 ;
        RECT 1642.290 2790.875 1642.570 2791.245 ;
        RECT 1642.360 2790.370 1642.500 2790.875 ;
        RECT 1645.580 2790.370 1645.720 2793.595 ;
        RECT 1646.430 2792.915 1646.710 2793.285 ;
        RECT 1642.300 2790.050 1642.560 2790.370 ;
        RECT 1645.520 2790.050 1645.780 2790.370 ;
        RECT 1638.620 2789.710 1638.880 2790.030 ;
        RECT 1638.680 2304.510 1638.820 2789.710 ;
        RECT 1645.580 2311.650 1645.720 2790.050 ;
        RECT 1646.500 2788.330 1646.640 2792.915 ;
        RECT 1649.190 2791.555 1649.470 2791.925 ;
        RECT 1649.260 2791.390 1649.400 2791.555 ;
        RECT 1649.200 2791.070 1649.460 2791.390 ;
        RECT 1646.440 2788.010 1646.700 2788.330 ;
        RECT 1646.500 2325.250 1646.640 2788.010 ;
        RECT 1646.440 2324.930 1646.700 2325.250 ;
        RECT 1645.520 2311.330 1645.780 2311.650 ;
        RECT 1638.620 2304.190 1638.880 2304.510 ;
        RECT 1649.720 1607.850 1649.860 2794.275 ;
        RECT 1652.410 2792.915 1652.690 2793.285 ;
        RECT 1652.480 2787.990 1652.620 2792.915 ;
        RECT 1658.920 2792.410 1659.060 2794.275 ;
        RECT 1656.560 2792.090 1656.820 2792.410 ;
        RECT 1658.860 2792.090 1659.120 2792.410 ;
        RECT 1656.090 2790.875 1656.370 2791.245 ;
        RECT 1656.160 2790.710 1656.300 2790.875 ;
        RECT 1656.100 2790.390 1656.360 2790.710 ;
        RECT 1656.620 2789.690 1656.760 2792.090 ;
        RECT 1656.560 2789.370 1656.820 2789.690 ;
        RECT 1652.420 2787.670 1652.680 2787.990 ;
        RECT 1652.480 2332.050 1652.620 2787.670 ;
        RECT 1652.420 2331.730 1652.680 2332.050 ;
        RECT 1663.060 1628.250 1663.200 2794.275 ;
        RECT 1663.450 2793.595 1663.730 2793.965 ;
        RECT 1663.520 2792.070 1663.660 2793.595 ;
        RECT 1663.460 2791.750 1663.720 2792.070 ;
        RECT 1663.520 2789.350 1663.660 2791.750 ;
        RECT 1663.460 2789.030 1663.720 2789.350 ;
        RECT 1669.960 1642.190 1670.100 2794.275 ;
        RECT 1670.350 2793.595 1670.630 2793.965 ;
        RECT 1670.420 2791.390 1670.560 2793.595 ;
        RECT 1670.360 2791.070 1670.620 2791.390 ;
        RECT 1670.420 2789.010 1670.560 2791.070 ;
        RECT 1670.360 2788.690 1670.620 2789.010 ;
        RECT 1676.860 1648.990 1677.000 2794.275 ;
        RECT 1677.260 2794.130 1677.520 2794.450 ;
        RECT 1683.690 2794.275 1683.970 2794.645 ;
        RECT 1686.910 2794.275 1687.190 2794.645 ;
        RECT 1690.590 2794.275 1690.870 2794.645 ;
        RECT 1697.490 2794.275 1697.770 2794.645 ;
        RECT 1704.390 2794.275 1704.670 2794.645 ;
        RECT 1711.290 2794.275 1711.570 2794.645 ;
        RECT 1718.190 2794.275 1718.470 2794.645 ;
        RECT 1721.410 2794.275 1721.690 2794.645 ;
        RECT 1725.090 2794.275 1725.370 2794.645 ;
        RECT 1731.990 2794.275 1732.270 2794.645 ;
        RECT 1738.890 2794.275 1739.170 2794.645 ;
        RECT 1677.320 2793.965 1677.460 2794.130 ;
        RECT 1677.250 2793.595 1677.530 2793.965 ;
        RECT 1683.230 2793.595 1683.510 2793.965 ;
        RECT 1677.320 2788.670 1677.460 2793.595 ;
        RECT 1683.300 2793.090 1683.440 2793.595 ;
        RECT 1683.240 2792.770 1683.500 2793.090 ;
        RECT 1683.300 2790.030 1683.440 2792.770 ;
        RECT 1683.240 2789.710 1683.500 2790.030 ;
        RECT 1677.260 2788.350 1677.520 2788.670 ;
        RECT 1683.760 1662.930 1683.900 2794.275 ;
        RECT 1686.980 2792.750 1687.120 2794.275 ;
        RECT 1684.150 2792.235 1684.430 2792.605 ;
        RECT 1686.920 2792.430 1687.180 2792.750 ;
        RECT 1684.220 1676.530 1684.360 2792.235 ;
        RECT 1686.980 2790.370 1687.120 2792.430 ;
        RECT 1686.920 2790.050 1687.180 2790.370 ;
        RECT 1690.660 1683.670 1690.800 2794.275 ;
        RECT 1694.730 2793.595 1695.010 2793.965 ;
        RECT 1694.800 2793.430 1694.940 2793.595 ;
        RECT 1694.740 2793.110 1695.000 2793.430 ;
        RECT 1694.800 2788.330 1694.940 2793.110 ;
        RECT 1694.740 2788.010 1695.000 2788.330 ;
        RECT 1697.560 1697.270 1697.700 2794.275 ;
        RECT 1699.330 2793.595 1699.610 2793.965 ;
        RECT 1699.400 2791.730 1699.540 2793.595 ;
        RECT 1699.340 2791.410 1699.600 2791.730 ;
        RECT 1699.400 2787.990 1699.540 2791.410 ;
        RECT 1699.340 2787.670 1699.600 2787.990 ;
        RECT 1704.460 1704.410 1704.600 2794.275 ;
        RECT 1704.850 2793.595 1705.130 2793.965 ;
        RECT 1704.920 2792.410 1705.060 2793.595 ;
        RECT 1704.860 2792.090 1705.120 2792.410 ;
        RECT 1711.360 1718.010 1711.500 2794.275 ;
        RECT 1712.670 2793.595 1712.950 2793.965 ;
        RECT 1712.740 2792.070 1712.880 2793.595 ;
        RECT 1712.680 2791.750 1712.940 2792.070 ;
        RECT 1718.260 1731.950 1718.400 2794.275 ;
        RECT 1721.420 2794.130 1721.680 2794.275 ;
        RECT 1718.660 2793.965 1718.920 2794.110 ;
        RECT 1718.650 2793.595 1718.930 2793.965 ;
        RECT 1721.480 2793.770 1721.620 2794.130 ;
        RECT 1718.720 2791.390 1718.860 2793.595 ;
        RECT 1721.420 2793.450 1721.680 2793.770 ;
        RECT 1718.660 2791.070 1718.920 2791.390 ;
        RECT 1718.650 2788.155 1718.930 2788.525 ;
        RECT 1718.720 1738.750 1718.860 2788.155 ;
        RECT 1725.160 1752.690 1725.300 2794.275 ;
        RECT 1731.530 2793.595 1731.810 2793.965 ;
        RECT 1731.600 2793.090 1731.740 2793.595 ;
        RECT 1731.540 2792.770 1731.800 2793.090 ;
        RECT 1731.600 2791.390 1731.740 2792.770 ;
        RECT 1731.540 2791.070 1731.800 2791.390 ;
        RECT 1732.060 1759.490 1732.200 2794.275 ;
        RECT 1734.750 2793.595 1735.030 2793.965 ;
        RECT 1734.820 2793.090 1734.960 2793.595 ;
        RECT 1734.760 2792.770 1735.020 2793.090 ;
        RECT 1738.960 1773.430 1739.100 2794.275 ;
        RECT 1739.880 2792.070 1740.020 2796.315 ;
        RECT 1745.790 2794.275 1746.070 2794.645 ;
        RECT 1759.590 2794.275 1759.870 2794.645 ;
        RECT 1741.650 2793.595 1741.930 2793.965 ;
        RECT 1741.720 2793.430 1741.860 2793.595 ;
        RECT 1741.660 2793.110 1741.920 2793.430 ;
        RECT 1739.820 2791.750 1740.080 2792.070 ;
        RECT 1745.860 1787.030 1746.000 2794.275 ;
        RECT 1759.660 2794.110 1759.800 2794.275 ;
        RECT 1776.620 2794.130 1776.880 2794.450 ;
        RECT 1747.630 2793.595 1747.910 2793.965 ;
        RECT 1759.600 2793.790 1759.860 2794.110 ;
        RECT 1766.490 2793.595 1766.770 2793.965 ;
        RECT 1747.700 2791.730 1747.840 2793.595 ;
        RECT 1766.500 2793.450 1766.760 2793.595 ;
        RECT 1752.690 2792.235 1752.970 2792.605 ;
        RECT 1752.700 2792.090 1752.960 2792.235 ;
        RECT 1747.640 2791.410 1747.900 2791.730 ;
        RECT 1773.390 2791.555 1773.670 2791.925 ;
        RECT 1773.460 2791.390 1773.600 2791.555 ;
        RECT 1773.400 2791.070 1773.660 2791.390 ;
        RECT 1749.020 2790.390 1749.280 2790.710 ;
        RECT 1749.080 2359.930 1749.220 2790.390 ;
        RECT 1762.820 2790.050 1763.080 2790.370 ;
        RECT 1760.050 2788.155 1760.330 2788.525 ;
        RECT 1752.690 2787.475 1752.970 2787.845 ;
        RECT 1749.020 2359.610 1749.280 2359.930 ;
        RECT 1752.760 1793.830 1752.900 2787.475 ;
        RECT 1760.120 1814.570 1760.260 2788.155 ;
        RECT 1760.970 2777.275 1761.250 2777.645 ;
        RECT 1760.060 1814.250 1760.320 1814.570 ;
        RECT 1761.040 1807.770 1761.180 2777.275 ;
        RECT 1762.880 2573.790 1763.020 2790.050 ;
        RECT 1763.280 2789.710 1763.540 2790.030 ;
        RECT 1763.340 2587.390 1763.480 2789.710 ;
        RECT 1763.740 2789.370 1764.000 2789.690 ;
        RECT 1763.800 2601.330 1763.940 2789.370 ;
        RECT 1769.720 2789.030 1769.980 2789.350 ;
        RECT 1766.490 2787.475 1766.770 2787.845 ;
        RECT 1763.740 2601.010 1764.000 2601.330 ;
        RECT 1763.280 2587.070 1763.540 2587.390 ;
        RECT 1762.820 2573.470 1763.080 2573.790 ;
        RECT 1766.560 1828.510 1766.700 2787.475 ;
        RECT 1769.780 2608.130 1769.920 2789.030 ;
        RECT 1770.180 2788.350 1770.440 2788.670 ;
        RECT 1770.240 2622.070 1770.380 2788.350 ;
        RECT 1773.850 2787.475 1774.130 2787.845 ;
        RECT 1770.180 2621.750 1770.440 2622.070 ;
        RECT 1769.720 2607.810 1769.980 2608.130 ;
        RECT 1773.920 1842.450 1774.060 2787.475 ;
        RECT 1776.680 2628.870 1776.820 2794.130 ;
        RECT 1787.190 2793.595 1787.470 2793.965 ;
        RECT 1787.260 2793.430 1787.400 2793.595 ;
        RECT 1780.290 2792.915 1780.570 2793.285 ;
        RECT 1787.200 2793.110 1787.460 2793.430 ;
        RECT 1780.300 2792.770 1780.560 2792.915 ;
        RECT 1783.980 2792.770 1784.240 2793.090 ;
        RECT 1783.520 2788.690 1783.780 2789.010 ;
        RECT 1780.290 2787.475 1780.570 2787.845 ;
        RECT 1776.620 2628.550 1776.880 2628.870 ;
        RECT 1780.360 1849.250 1780.500 2787.475 ;
        RECT 1783.580 2642.810 1783.720 2788.690 ;
        RECT 1784.040 2656.410 1784.180 2792.770 ;
        RECT 1788.640 2791.730 1788.780 2796.315 ;
        RECT 1790.880 2791.750 1791.140 2792.070 ;
        RECT 1788.580 2791.410 1788.840 2791.730 ;
        RECT 1790.420 2788.010 1790.680 2788.330 ;
        RECT 1787.190 2787.475 1787.470 2787.845 ;
        RECT 1783.980 2656.090 1784.240 2656.410 ;
        RECT 1783.520 2642.490 1783.780 2642.810 ;
        RECT 1787.260 1862.850 1787.400 2787.475 ;
        RECT 1790.480 2366.730 1790.620 2788.010 ;
        RECT 1790.940 2380.330 1791.080 2791.750 ;
        RECT 1797.320 2791.410 1797.580 2791.730 ;
        RECT 1794.090 2777.275 1794.370 2777.645 ;
        RECT 1790.880 2380.010 1791.140 2380.330 ;
        RECT 1790.420 2366.410 1790.680 2366.730 ;
        RECT 1794.160 1869.990 1794.300 2777.275 ;
        RECT 1797.380 2387.470 1797.520 2791.410 ;
        RECT 1797.780 2791.070 1798.040 2791.390 ;
        RECT 1797.840 2401.070 1797.980 2791.070 ;
        RECT 1797.780 2400.750 1798.040 2401.070 ;
        RECT 1797.320 2387.150 1797.580 2387.470 ;
        RECT 1942.280 2000.890 1942.420 3187.850 ;
        RECT 1945.960 2948.325 1946.100 3248.630 ;
        RECT 2187.390 3230.835 2187.670 3231.205 ;
        RECT 2187.460 3229.650 2187.600 3230.835 ;
        RECT 1997.420 3229.330 1997.680 3229.650 ;
        RECT 2187.400 3229.330 2187.660 3229.650 ;
        RECT 1990.520 3222.190 1990.780 3222.510 ;
        RECT 1976.720 3215.390 1976.980 3215.710 ;
        RECT 1969.820 3208.590 1970.080 3208.910 ;
        RECT 1962.920 3201.450 1963.180 3201.770 ;
        RECT 1956.020 3194.650 1956.280 3194.970 ;
        RECT 1945.890 2947.955 1946.170 2948.325 ;
        RECT 1956.080 2014.830 1956.220 3194.650 ;
        RECT 1962.980 2028.430 1963.120 3201.450 ;
        RECT 1969.880 2035.570 1970.020 3208.590 ;
        RECT 1976.780 2049.170 1976.920 3215.390 ;
        RECT 1990.580 2056.310 1990.720 3222.190 ;
        RECT 1997.480 2069.910 1997.620 3229.330 ;
        RECT 2187.390 3224.035 2187.670 3224.405 ;
        RECT 2187.460 3222.510 2187.600 3224.035 ;
        RECT 2187.400 3222.190 2187.660 3222.510 ;
        RECT 2187.390 3215.875 2187.670 3216.245 ;
        RECT 2187.460 3215.710 2187.600 3215.875 ;
        RECT 2187.400 3215.390 2187.660 3215.710 ;
        RECT 2187.390 3209.755 2187.670 3210.125 ;
        RECT 2187.460 3208.910 2187.600 3209.755 ;
        RECT 2187.400 3208.590 2187.660 3208.910 ;
        RECT 2187.390 3201.595 2187.670 3201.965 ;
        RECT 2187.400 3201.450 2187.660 3201.595 ;
        RECT 2187.390 3196.155 2187.670 3196.525 ;
        RECT 2187.460 3194.970 2187.600 3196.155 ;
        RECT 2187.400 3194.650 2187.660 3194.970 ;
        RECT 2187.390 3187.995 2187.670 3188.365 ;
        RECT 2187.400 3187.850 2187.660 3187.995 ;
        RECT 2011.220 2898.170 2011.480 2898.490 ;
        RECT 2187.390 2898.315 2187.670 2898.685 ;
        RECT 2187.400 2898.170 2187.660 2898.315 ;
        RECT 1997.420 2069.590 1997.680 2069.910 ;
        RECT 1990.520 2055.990 1990.780 2056.310 ;
        RECT 1976.720 2048.850 1976.980 2049.170 ;
        RECT 1969.820 2035.250 1970.080 2035.570 ;
        RECT 1962.920 2028.110 1963.180 2028.430 ;
        RECT 1956.020 2014.510 1956.280 2014.830 ;
        RECT 1942.220 2000.570 1942.480 2000.890 ;
        RECT 2011.280 1973.350 2011.420 2898.170 ;
        RECT 2190.610 2891.515 2190.890 2891.885 ;
        RECT 2190.680 2804.650 2190.820 2891.515 ;
      LAYER met2 ;
        RECT 2205.000 2805.000 2581.480 3251.235 ;
      LAYER met2 ;
        RECT 2582.140 3249.565 2582.280 3251.770 ;
        RECT 2582.070 3249.195 2582.350 3249.565 ;
        RECT 2594.560 2946.965 2594.700 3264.010 ;
        RECT 2594.490 2946.595 2594.770 2946.965 ;
        RECT 2594.560 2938.805 2594.700 2946.595 ;
        RECT 2594.490 2938.435 2594.770 2938.805 ;
        RECT 2190.620 2804.330 2190.880 2804.650 ;
        RECT 2228.790 2794.275 2229.070 2794.645 ;
        RECT 2232.010 2794.275 2232.290 2794.645 ;
        RECT 2238.910 2794.275 2239.190 2794.645 ;
        RECT 2245.810 2794.275 2246.090 2794.645 ;
        RECT 2263.750 2794.275 2264.030 2794.645 ;
        RECT 2267.430 2794.275 2267.710 2794.645 ;
        RECT 2273.410 2794.275 2273.690 2794.645 ;
        RECT 2294.110 2794.275 2294.390 2794.645 ;
        RECT 2304.690 2794.275 2304.970 2794.645 ;
        RECT 2308.830 2794.275 2309.110 2794.645 ;
        RECT 2311.590 2794.275 2311.870 2794.645 ;
        RECT 2318.490 2794.275 2318.770 2794.645 ;
        RECT 2325.390 2794.275 2325.670 2794.645 ;
        RECT 2332.290 2794.275 2332.570 2794.645 ;
        RECT 2339.190 2794.275 2339.470 2794.645 ;
        RECT 2342.870 2794.275 2343.150 2794.645 ;
        RECT 2346.090 2794.275 2346.370 2794.645 ;
        RECT 2352.990 2794.275 2353.270 2794.645 ;
        RECT 2359.890 2794.275 2360.170 2794.645 ;
        RECT 2366.790 2794.275 2367.070 2794.645 ;
        RECT 2373.690 2794.275 2373.970 2794.645 ;
        RECT 2381.050 2794.275 2381.330 2794.645 ;
        RECT 2385.650 2794.275 2385.930 2794.645 ;
        RECT 2391.630 2794.275 2391.910 2794.645 ;
        RECT 2397.150 2794.275 2397.430 2794.645 ;
        RECT 2402.670 2794.275 2402.950 2794.645 ;
        RECT 2415.090 2794.275 2415.370 2794.645 ;
        RECT 2422.450 2794.275 2422.730 2794.645 ;
        RECT 2428.890 2794.275 2429.170 2794.645 ;
        RECT 2218.220 2790.730 2218.480 2791.050 ;
        RECT 2218.280 2415.010 2218.420 2790.730 ;
        RECT 2218.220 2414.690 2218.480 2415.010 ;
        RECT 2228.860 1994.090 2229.000 2794.275 ;
        RECT 2228.800 1993.770 2229.060 1994.090 ;
        RECT 2011.220 1973.030 2011.480 1973.350 ;
        RECT 2232.080 1883.590 2232.220 2794.275 ;
        RECT 2238.980 1897.530 2239.120 2794.275 ;
        RECT 2245.880 1904.330 2246.020 2794.275 ;
        RECT 2263.290 2790.875 2263.570 2791.245 ;
        RECT 2263.360 2790.710 2263.500 2790.875 ;
        RECT 2263.300 2790.390 2263.560 2790.710 ;
        RECT 2256.850 2788.155 2257.130 2788.525 ;
        RECT 2256.920 2787.990 2257.060 2788.155 ;
        RECT 2252.720 2787.670 2252.980 2787.990 ;
        RECT 2256.860 2787.670 2257.120 2787.990 ;
        RECT 2252.780 1918.270 2252.920 2787.670 ;
        RECT 2263.820 2345.990 2263.960 2794.275 ;
        RECT 2266.510 2793.595 2266.790 2793.965 ;
        RECT 2266.580 2792.410 2266.720 2793.595 ;
        RECT 2267.500 2793.090 2267.640 2794.275 ;
        RECT 2267.440 2792.770 2267.700 2793.090 ;
        RECT 2266.520 2792.090 2266.780 2792.410 ;
        RECT 2263.760 2345.670 2264.020 2345.990 ;
        RECT 2266.580 2166.470 2266.720 2792.090 ;
        RECT 2267.500 2180.410 2267.640 2792.770 ;
        RECT 2270.190 2791.555 2270.470 2791.925 ;
        RECT 2270.260 2788.330 2270.400 2791.555 ;
        RECT 2273.480 2790.710 2273.620 2794.275 ;
        RECT 2294.180 2794.110 2294.320 2794.275 ;
        RECT 2294.120 2793.790 2294.380 2794.110 ;
        RECT 2280.310 2792.915 2280.590 2793.285 ;
        RECT 2287.210 2792.915 2287.490 2793.285 ;
        RECT 2277.090 2792.235 2277.370 2792.605 ;
        RECT 2277.160 2792.070 2277.300 2792.235 ;
        RECT 2277.100 2791.750 2277.360 2792.070 ;
        RECT 2273.420 2790.390 2273.680 2790.710 ;
        RECT 2270.200 2788.010 2270.460 2788.330 ;
        RECT 2273.480 2194.350 2273.620 2790.390 ;
        RECT 2280.380 2788.330 2280.520 2792.915 ;
        RECT 2283.990 2791.555 2284.270 2791.925 ;
        RECT 2284.000 2791.410 2284.260 2791.555 ;
        RECT 2280.320 2788.010 2280.580 2788.330 ;
        RECT 2280.380 2201.150 2280.520 2788.010 ;
        RECT 2287.280 2787.990 2287.420 2792.915 ;
        RECT 2290.890 2791.555 2291.170 2791.925 ;
        RECT 2290.960 2791.390 2291.100 2791.555 ;
        RECT 2290.900 2791.070 2291.160 2791.390 ;
        RECT 2287.220 2787.670 2287.480 2787.990 ;
        RECT 2287.280 2214.750 2287.420 2787.670 ;
        RECT 2294.180 2221.890 2294.320 2793.790 ;
        RECT 2301.010 2793.595 2301.290 2793.965 ;
        RECT 2303.310 2793.595 2303.590 2793.965 ;
        RECT 2297.790 2790.875 2298.070 2791.245 ;
        RECT 2297.800 2790.730 2298.060 2790.875 ;
        RECT 2301.080 2235.490 2301.220 2793.595 ;
        RECT 2303.320 2793.450 2303.580 2793.595 ;
        RECT 2304.230 2792.915 2304.510 2793.285 ;
        RECT 2304.300 2792.750 2304.440 2792.915 ;
        RECT 2301.940 2792.430 2302.200 2792.750 ;
        RECT 2304.240 2792.430 2304.500 2792.750 ;
        RECT 2302.000 2249.430 2302.140 2792.430 ;
        RECT 2304.760 2421.810 2304.900 2794.275 ;
        RECT 2305.150 2793.595 2305.430 2793.965 ;
        RECT 2305.220 2435.750 2305.360 2793.595 ;
        RECT 2308.900 2792.410 2309.040 2794.275 ;
        RECT 2308.840 2792.090 2309.100 2792.410 ;
        RECT 2311.660 2442.550 2311.800 2794.275 ;
        RECT 2314.810 2793.595 2315.090 2793.965 ;
        RECT 2314.880 2793.090 2315.020 2793.595 ;
        RECT 2314.820 2792.770 2315.080 2793.090 ;
        RECT 2318.040 2792.770 2318.300 2793.090 ;
        RECT 2318.100 2792.070 2318.240 2792.770 ;
        RECT 2318.040 2791.750 2318.300 2792.070 ;
        RECT 2318.560 2456.490 2318.700 2794.275 ;
        RECT 2321.710 2793.595 2321.990 2793.965 ;
        RECT 2321.780 2793.090 2321.920 2793.595 ;
        RECT 2321.720 2792.770 2321.980 2793.090 ;
        RECT 2321.780 2791.130 2321.920 2792.770 ;
        RECT 2321.320 2790.990 2321.920 2791.130 ;
        RECT 2321.320 2790.710 2321.460 2790.990 ;
        RECT 2321.260 2790.390 2321.520 2790.710 ;
        RECT 2321.720 2790.390 2321.980 2790.710 ;
        RECT 2321.780 2663.550 2321.920 2790.390 ;
        RECT 2321.720 2663.230 2321.980 2663.550 ;
        RECT 2325.460 2470.090 2325.600 2794.275 ;
        RECT 2325.850 2793.595 2326.130 2793.965 ;
        RECT 2325.920 2791.730 2326.060 2793.595 ;
        RECT 2325.860 2791.410 2326.120 2791.730 ;
        RECT 2325.920 2788.330 2326.060 2791.410 ;
        RECT 2328.620 2790.730 2328.880 2791.050 ;
        RECT 2325.860 2788.010 2326.120 2788.330 ;
        RECT 2328.680 2677.150 2328.820 2790.730 ;
        RECT 2328.620 2676.830 2328.880 2677.150 ;
        RECT 2332.360 2477.230 2332.500 2794.275 ;
        RECT 2332.750 2792.915 2333.030 2793.285 ;
        RECT 2332.820 2787.990 2332.960 2792.915 ;
        RECT 2335.520 2791.070 2335.780 2791.390 ;
        RECT 2332.760 2787.670 2333.020 2787.990 ;
        RECT 2335.580 2683.950 2335.720 2791.070 ;
        RECT 2335.520 2683.630 2335.780 2683.950 ;
        RECT 2339.260 2490.830 2339.400 2794.275 ;
        RECT 2339.650 2793.595 2339.930 2793.965 ;
        RECT 2340.120 2793.790 2340.380 2794.110 ;
        RECT 2339.720 2497.630 2339.860 2793.595 ;
        RECT 2340.180 2793.285 2340.320 2793.790 ;
        RECT 2342.940 2793.770 2343.080 2794.275 ;
        RECT 2342.880 2793.450 2343.140 2793.770 ;
        RECT 2340.110 2792.915 2340.390 2793.285 ;
        RECT 2342.940 2788.330 2343.080 2793.450 ;
        RECT 2342.880 2788.010 2343.140 2788.330 ;
        RECT 2346.160 2511.570 2346.300 2794.275 ;
        RECT 2350.230 2793.595 2350.510 2793.965 ;
        RECT 2350.300 2792.750 2350.440 2793.595 ;
        RECT 2350.240 2792.430 2350.500 2792.750 ;
        RECT 2353.060 2518.370 2353.200 2794.275 ;
        RECT 2356.210 2793.595 2356.490 2793.965 ;
        RECT 2356.280 2792.410 2356.420 2793.595 ;
        RECT 2356.220 2792.090 2356.480 2792.410 ;
        RECT 2359.960 2532.310 2360.100 2794.275 ;
        RECT 2361.270 2793.595 2361.550 2793.965 ;
        RECT 2361.340 2792.070 2361.480 2793.595 ;
        RECT 2361.280 2791.750 2361.540 2792.070 ;
        RECT 2366.860 2546.250 2367.000 2794.275 ;
        RECT 2367.710 2793.595 2367.990 2793.965 ;
        RECT 2367.780 2793.090 2367.920 2793.595 ;
        RECT 2367.720 2792.770 2367.980 2793.090 ;
        RECT 2373.230 2788.155 2373.510 2788.525 ;
        RECT 2373.300 2787.990 2373.440 2788.155 ;
        RECT 2373.240 2787.670 2373.500 2787.990 ;
        RECT 2373.760 2553.050 2373.900 2794.275 ;
        RECT 2374.150 2793.595 2374.430 2793.965 ;
        RECT 2377.830 2793.595 2378.110 2793.965 ;
        RECT 2374.220 2791.730 2374.360 2793.595 ;
        RECT 2377.840 2793.450 2378.100 2793.595 ;
        RECT 2374.160 2791.410 2374.420 2791.730 ;
        RECT 2374.220 2787.990 2374.360 2791.410 ;
        RECT 2380.590 2790.195 2380.870 2790.565 ;
        RECT 2380.600 2790.050 2380.860 2790.195 ;
        RECT 2374.160 2787.670 2374.420 2787.990 ;
        RECT 2381.120 2566.650 2381.260 2794.275 ;
        RECT 2385.720 2794.110 2385.860 2794.275 ;
        RECT 2385.660 2793.790 2385.920 2794.110 ;
        RECT 2391.700 2791.730 2391.840 2794.275 ;
        RECT 2397.220 2792.750 2397.360 2794.275 ;
        RECT 2402.210 2793.595 2402.490 2793.965 ;
        RECT 2397.160 2792.430 2397.420 2792.750 ;
        RECT 2402.280 2792.410 2402.420 2793.595 ;
        RECT 2402.220 2792.090 2402.480 2792.410 ;
        RECT 2387.960 2791.410 2388.220 2791.730 ;
        RECT 2391.640 2791.410 2391.900 2791.730 ;
        RECT 2387.490 2790.195 2387.770 2790.565 ;
        RECT 2387.560 2790.030 2387.700 2790.195 ;
        RECT 2387.500 2789.710 2387.760 2790.030 ;
        RECT 2388.020 2788.330 2388.160 2791.410 ;
        RECT 2394.390 2789.515 2394.670 2789.885 ;
        RECT 2394.400 2789.370 2394.660 2789.515 ;
        RECT 2402.740 2789.350 2402.880 2794.275 ;
        RECT 2415.100 2794.130 2415.360 2794.275 ;
        RECT 2421.990 2793.595 2422.270 2793.965 ;
        RECT 2422.000 2793.450 2422.260 2793.595 ;
        RECT 2422.520 2793.430 2422.660 2794.275 ;
        RECT 2428.960 2794.110 2429.100 2794.275 ;
        RECT 2428.900 2793.790 2429.160 2794.110 ;
        RECT 2415.090 2792.915 2415.370 2793.285 ;
        RECT 2422.460 2793.110 2422.720 2793.430 ;
        RECT 2442.690 2792.915 2442.970 2793.285 ;
        RECT 2415.100 2792.770 2415.360 2792.915 ;
        RECT 2442.760 2792.750 2442.900 2792.915 ;
        RECT 2408.190 2792.235 2408.470 2792.605 ;
        RECT 2435.790 2792.235 2436.070 2792.605 ;
        RECT 2442.700 2792.430 2442.960 2792.750 ;
        RECT 2408.260 2792.070 2408.400 2792.235 ;
        RECT 2408.200 2791.750 2408.460 2792.070 ;
        RECT 2435.860 2791.730 2436.000 2792.235 ;
        RECT 2435.800 2791.410 2436.060 2791.730 ;
        RECT 2442.690 2791.555 2442.970 2791.925 ;
        RECT 2442.760 2791.390 2442.900 2791.555 ;
        RECT 2415.090 2790.875 2415.370 2791.245 ;
        RECT 2428.890 2790.875 2429.170 2791.245 ;
        RECT 2435.790 2790.875 2436.070 2791.245 ;
        RECT 2442.700 2791.070 2442.960 2791.390 ;
        RECT 2402.680 2789.030 2402.940 2789.350 ;
        RECT 2408.190 2788.835 2408.470 2789.205 ;
        RECT 2415.160 2789.010 2415.300 2790.875 ;
        RECT 2428.960 2790.710 2429.100 2790.875 ;
        RECT 2435.800 2790.730 2436.060 2790.875 ;
        RECT 2428.900 2790.390 2429.160 2790.710 ;
        RECT 2408.260 2788.670 2408.400 2788.835 ;
        RECT 2415.100 2788.690 2415.360 2789.010 ;
        RECT 2408.200 2788.350 2408.460 2788.670 ;
        RECT 2387.960 2788.010 2388.220 2788.330 ;
        RECT 2415.090 2788.155 2415.370 2788.525 ;
        RECT 2415.160 2787.990 2415.300 2788.155 ;
        RECT 2415.100 2787.670 2415.360 2787.990 ;
        RECT 2381.060 2566.330 2381.320 2566.650 ;
        RECT 2373.700 2552.730 2373.960 2553.050 ;
        RECT 2366.800 2545.930 2367.060 2546.250 ;
        RECT 2359.900 2531.990 2360.160 2532.310 ;
        RECT 2353.000 2518.050 2353.260 2518.370 ;
        RECT 2346.100 2511.250 2346.360 2511.570 ;
        RECT 2339.660 2497.310 2339.920 2497.630 ;
        RECT 2339.200 2490.510 2339.460 2490.830 ;
        RECT 2332.300 2476.910 2332.560 2477.230 ;
        RECT 2325.400 2469.770 2325.660 2470.090 ;
        RECT 2318.500 2456.170 2318.760 2456.490 ;
        RECT 2311.600 2442.230 2311.860 2442.550 ;
        RECT 2305.160 2435.430 2305.420 2435.750 ;
        RECT 2304.700 2421.490 2304.960 2421.810 ;
        RECT 2301.940 2249.110 2302.200 2249.430 ;
        RECT 2301.020 2235.170 2301.280 2235.490 ;
        RECT 2294.120 2221.570 2294.380 2221.890 ;
        RECT 2287.220 2214.430 2287.480 2214.750 ;
        RECT 2280.320 2200.830 2280.580 2201.150 ;
        RECT 2273.420 2194.030 2273.680 2194.350 ;
        RECT 2267.440 2180.090 2267.700 2180.410 ;
        RECT 2266.520 2166.150 2266.780 2166.470 ;
        RECT 2252.720 1917.950 2252.980 1918.270 ;
        RECT 2245.820 1904.010 2246.080 1904.330 ;
        RECT 2238.920 1897.210 2239.180 1897.530 ;
        RECT 2232.020 1883.270 2232.280 1883.590 ;
        RECT 1794.100 1869.670 1794.360 1869.990 ;
        RECT 1787.200 1862.530 1787.460 1862.850 ;
        RECT 1780.300 1848.930 1780.560 1849.250 ;
        RECT 1773.860 1842.130 1774.120 1842.450 ;
        RECT 1766.500 1828.190 1766.760 1828.510 ;
        RECT 1760.980 1807.450 1761.240 1807.770 ;
        RECT 1752.700 1793.510 1752.960 1793.830 ;
        RECT 1745.800 1786.710 1746.060 1787.030 ;
        RECT 1738.900 1773.110 1739.160 1773.430 ;
        RECT 1732.000 1759.170 1732.260 1759.490 ;
        RECT 1725.100 1752.370 1725.360 1752.690 ;
        RECT 1718.660 1738.430 1718.920 1738.750 ;
        RECT 1718.200 1731.630 1718.460 1731.950 ;
        RECT 1711.300 1717.690 1711.560 1718.010 ;
        RECT 1704.400 1704.090 1704.660 1704.410 ;
        RECT 1697.500 1696.950 1697.760 1697.270 ;
        RECT 1690.600 1683.350 1690.860 1683.670 ;
        RECT 1684.160 1676.210 1684.420 1676.530 ;
        RECT 1683.700 1662.610 1683.960 1662.930 ;
        RECT 1676.800 1648.670 1677.060 1648.990 ;
        RECT 1669.900 1641.870 1670.160 1642.190 ;
        RECT 1663.000 1627.930 1663.260 1628.250 ;
        RECT 1649.660 1607.530 1649.920 1607.850 ;
        RECT 1635.400 1572.850 1635.660 1573.170 ;
        RECT 1628.500 1566.050 1628.760 1566.370 ;
        RECT 1617.920 1552.110 1618.180 1552.430 ;
        RECT 1410.460 1531.370 1410.720 1531.690 ;
        RECT 1607.800 1531.370 1608.060 1531.690 ;
        RECT 1410.520 1527.805 1410.660 1531.370 ;
        RECT 1410.450 1527.435 1410.730 1527.805 ;
        RECT 1408.150 1505.675 1408.430 1506.045 ;
      LAYER met2 ;
        RECT 305.250 1504.000 314.070 1504.280 ;
        RECT 314.910 1504.000 323.730 1504.280 ;
        RECT 324.570 1504.000 333.390 1504.280 ;
        RECT 334.230 1504.000 343.050 1504.280 ;
        RECT 343.890 1504.000 352.710 1504.280 ;
        RECT 353.550 1504.000 362.370 1504.280 ;
        RECT 363.210 1504.000 372.490 1504.280 ;
        RECT 373.330 1504.000 382.150 1504.280 ;
        RECT 382.990 1504.000 391.810 1504.280 ;
        RECT 392.650 1504.000 401.470 1504.280 ;
        RECT 402.310 1504.000 411.130 1504.280 ;
        RECT 411.970 1504.000 420.790 1504.280 ;
        RECT 421.630 1504.000 430.910 1504.280 ;
        RECT 431.750 1504.000 440.570 1504.280 ;
        RECT 441.410 1504.000 450.230 1504.280 ;
        RECT 451.070 1504.000 459.890 1504.280 ;
        RECT 460.730 1504.000 469.550 1504.280 ;
        RECT 470.390 1504.000 479.210 1504.280 ;
        RECT 480.050 1504.000 489.330 1504.280 ;
        RECT 490.170 1504.000 498.990 1504.280 ;
        RECT 499.830 1504.000 508.650 1504.280 ;
        RECT 509.490 1504.000 518.310 1504.280 ;
        RECT 519.150 1504.000 527.970 1504.280 ;
        RECT 528.810 1504.000 537.630 1504.280 ;
        RECT 538.470 1504.000 547.290 1504.280 ;
        RECT 548.130 1504.000 557.410 1504.280 ;
        RECT 558.250 1504.000 567.070 1504.280 ;
        RECT 567.910 1504.000 576.730 1504.280 ;
        RECT 577.570 1504.000 586.390 1504.280 ;
        RECT 587.230 1504.000 596.050 1504.280 ;
        RECT 596.890 1504.000 605.710 1504.280 ;
        RECT 606.550 1504.000 615.830 1504.280 ;
        RECT 616.670 1504.000 625.490 1504.280 ;
        RECT 626.330 1504.000 635.150 1504.280 ;
        RECT 635.990 1504.000 644.810 1504.280 ;
        RECT 645.650 1504.000 654.470 1504.280 ;
        RECT 655.310 1504.000 664.130 1504.280 ;
        RECT 664.970 1504.000 674.250 1504.280 ;
        RECT 675.090 1504.000 683.910 1504.280 ;
        RECT 684.750 1504.000 693.570 1504.280 ;
        RECT 694.410 1504.000 703.230 1504.280 ;
        RECT 704.070 1504.000 712.890 1504.280 ;
        RECT 713.730 1504.000 722.550 1504.280 ;
        RECT 723.390 1504.000 732.670 1504.280 ;
        RECT 733.510 1504.000 742.330 1504.280 ;
        RECT 743.170 1504.000 751.990 1504.280 ;
        RECT 752.830 1504.000 761.650 1504.280 ;
        RECT 762.490 1504.000 771.310 1504.280 ;
        RECT 772.150 1504.000 780.970 1504.280 ;
        RECT 781.810 1504.000 790.630 1504.280 ;
        RECT 791.470 1504.000 800.750 1504.280 ;
        RECT 801.590 1504.000 810.410 1504.280 ;
        RECT 811.250 1504.000 820.070 1504.280 ;
        RECT 820.910 1504.000 829.730 1504.280 ;
        RECT 830.570 1504.000 839.390 1504.280 ;
        RECT 840.230 1504.000 849.050 1504.280 ;
        RECT 849.890 1504.000 859.170 1504.280 ;
        RECT 860.010 1504.000 868.830 1504.280 ;
        RECT 869.670 1504.000 878.490 1504.280 ;
        RECT 879.330 1504.000 888.150 1504.280 ;
        RECT 888.990 1504.000 897.810 1504.280 ;
        RECT 898.650 1504.000 907.470 1504.280 ;
        RECT 908.310 1504.000 917.590 1504.280 ;
        RECT 918.430 1504.000 927.250 1504.280 ;
        RECT 928.090 1504.000 936.910 1504.280 ;
        RECT 937.750 1504.000 946.570 1504.280 ;
        RECT 947.410 1504.000 956.230 1504.280 ;
        RECT 957.070 1504.000 965.890 1504.280 ;
        RECT 966.730 1504.000 975.550 1504.280 ;
        RECT 976.390 1504.000 985.670 1504.280 ;
        RECT 986.510 1504.000 995.330 1504.280 ;
        RECT 996.170 1504.000 1004.990 1504.280 ;
        RECT 1005.830 1504.000 1014.650 1504.280 ;
        RECT 1015.490 1504.000 1024.310 1504.280 ;
        RECT 1025.150 1504.000 1033.970 1504.280 ;
        RECT 1034.810 1504.000 1044.090 1504.280 ;
        RECT 1044.930 1504.000 1053.750 1504.280 ;
        RECT 1054.590 1504.000 1063.410 1504.280 ;
        RECT 1064.250 1504.000 1073.070 1504.280 ;
        RECT 1073.910 1504.000 1082.730 1504.280 ;
        RECT 1083.570 1504.000 1092.390 1504.280 ;
        RECT 1093.230 1504.000 1102.510 1504.280 ;
        RECT 1103.350 1504.000 1112.170 1504.280 ;
        RECT 1113.010 1504.000 1121.830 1504.280 ;
        RECT 1122.670 1504.000 1131.490 1504.280 ;
        RECT 1132.330 1504.000 1141.150 1504.280 ;
        RECT 1141.990 1504.000 1150.810 1504.280 ;
        RECT 1151.650 1504.000 1160.930 1504.280 ;
        RECT 1161.770 1504.000 1170.590 1504.280 ;
        RECT 1171.430 1504.000 1180.250 1504.280 ;
        RECT 1181.090 1504.000 1189.910 1504.280 ;
        RECT 1190.750 1504.000 1199.570 1504.280 ;
        RECT 1200.410 1504.000 1209.230 1504.280 ;
        RECT 1210.070 1504.000 1218.890 1504.280 ;
        RECT 1219.730 1504.000 1229.010 1504.280 ;
        RECT 1229.850 1504.000 1238.670 1504.280 ;
        RECT 1239.510 1504.000 1248.330 1504.280 ;
        RECT 1249.170 1504.000 1257.990 1504.280 ;
        RECT 1258.830 1504.000 1267.650 1504.280 ;
        RECT 1268.490 1504.000 1277.310 1504.280 ;
        RECT 1278.150 1504.000 1287.430 1504.280 ;
        RECT 1288.270 1504.000 1297.090 1504.280 ;
        RECT 1297.930 1504.000 1306.750 1504.280 ;
        RECT 1307.590 1504.000 1316.410 1504.280 ;
        RECT 1317.250 1504.000 1326.070 1504.280 ;
        RECT 1326.910 1504.000 1335.730 1504.280 ;
        RECT 1336.570 1504.000 1345.850 1504.280 ;
        RECT 1346.690 1504.000 1355.510 1504.280 ;
        RECT 1356.350 1504.000 1365.170 1504.280 ;
        RECT 1366.010 1504.000 1374.830 1504.280 ;
        RECT 1375.670 1504.000 1384.490 1504.280 ;
        RECT 1385.330 1504.000 1394.150 1504.280 ;
        RECT 1394.990 1504.000 1395.630 1504.280 ;
      LAYER via2 ;
        RECT 646.390 3264.200 646.670 3264.480 ;
        RECT 668.010 3264.200 668.290 3264.480 ;
        RECT 1295.910 3264.200 1296.190 3264.480 ;
        RECT 1318.910 3264.200 1319.190 3264.480 ;
        RECT 1892.530 3264.200 1892.810 3264.480 ;
        RECT 1917.370 3264.200 1917.650 3264.480 ;
        RECT 2539.290 3264.200 2539.570 3264.480 ;
        RECT 2566.890 3264.200 2567.170 3264.480 ;
        RECT 282.990 3230.200 283.270 3230.480 ;
        RECT 286.210 3224.760 286.490 3225.040 ;
        RECT 285.750 3215.920 286.030 3216.200 ;
        RECT 285.290 3209.800 285.570 3210.080 ;
        RECT 284.830 3201.640 285.110 3201.920 ;
        RECT 284.370 3196.200 284.650 3196.480 ;
        RECT 283.910 3188.040 284.190 3188.320 ;
        RECT 283.450 2898.360 283.730 2898.640 ;
        RECT 298.170 2892.635 298.450 2892.915 ;
        RECT 696.990 3249.240 697.270 3249.520 ;
        RECT 337.730 2794.320 338.010 2794.600 ;
        RECT 350.610 2794.320 350.890 2794.600 ;
        RECT 362.110 2794.320 362.390 2794.600 ;
        RECT 368.550 2794.320 368.830 2794.600 ;
        RECT 378.670 2794.320 378.950 2794.600 ;
        RECT 380.050 2794.320 380.330 2794.600 ;
        RECT 386.950 2794.320 387.230 2794.600 ;
        RECT 392.470 2794.320 392.750 2794.600 ;
        RECT 282.990 2714.760 283.270 2715.040 ;
        RECT 344.630 2790.240 344.910 2790.520 ;
        RECT 351.070 2793.640 351.350 2793.920 ;
        RECT 386.490 2791.600 386.770 2791.880 ;
        RECT 365.790 2790.920 366.070 2791.200 ;
        RECT 357.970 2787.520 358.250 2787.800 ;
        RECT 358.890 2788.200 359.170 2788.480 ;
        RECT 372.690 2788.880 372.970 2789.160 ;
        RECT 397.530 2794.320 397.810 2794.600 ;
        RECT 403.510 2794.320 403.790 2794.600 ;
        RECT 407.190 2794.320 407.470 2794.600 ;
        RECT 393.390 2789.560 393.670 2789.840 ;
        RECT 379.590 2788.880 379.870 2789.160 ;
        RECT 393.390 2788.200 393.670 2788.480 ;
        RECT 414.550 2794.320 414.830 2794.600 ;
        RECT 420.990 2794.320 421.270 2794.600 ;
        RECT 426.970 2794.320 427.250 2794.600 ;
        RECT 428.350 2794.320 428.630 2794.600 ;
        RECT 431.110 2794.320 431.390 2794.600 ;
        RECT 400.290 2793.640 400.570 2793.920 ;
        RECT 408.110 2793.640 408.390 2793.920 ;
        RECT 414.090 2791.600 414.370 2791.880 ;
        RECT 421.450 2793.640 421.730 2793.920 ;
        RECT 438.010 2794.320 438.290 2794.600 ;
        RECT 444.910 2794.320 445.190 2794.600 ;
        RECT 448.130 2794.320 448.410 2794.600 ;
        RECT 450.430 2794.320 450.710 2794.600 ;
        RECT 434.330 2793.640 434.610 2793.920 ;
        RECT 439.390 2793.640 439.670 2793.920 ;
        RECT 456.870 2794.320 457.150 2794.600 ;
        RECT 462.390 2794.320 462.670 2794.600 ;
        RECT 467.910 2794.320 468.190 2794.600 ;
        RECT 472.970 2794.320 473.250 2794.600 ;
        RECT 476.650 2794.320 476.930 2794.600 ;
        RECT 483.090 2794.320 483.370 2794.600 ;
        RECT 491.370 2794.320 491.650 2794.600 ;
        RECT 497.810 2794.320 498.090 2794.600 ;
        RECT 503.330 2794.320 503.610 2794.600 ;
        RECT 509.770 2794.320 510.050 2794.600 ;
        RECT 513.450 2794.320 513.730 2794.600 ;
        RECT 517.130 2794.320 517.410 2794.600 ;
        RECT 519.890 2794.320 520.170 2794.600 ;
        RECT 524.030 2794.320 524.310 2794.600 ;
        RECT 526.790 2794.320 527.070 2794.600 ;
        RECT 530.930 2794.320 531.210 2794.600 ;
        RECT 537.830 2794.320 538.110 2794.600 ;
        RECT 539.210 2794.320 539.490 2794.600 ;
        RECT 544.730 2794.320 545.010 2794.600 ;
        RECT 551.630 2794.320 551.910 2794.600 ;
        RECT 501.490 2793.640 501.770 2793.920 ;
        RECT 468.370 2788.200 468.650 2788.480 ;
        RECT 455.030 2787.520 455.310 2787.800 ;
        RECT 461.930 2787.520 462.210 2787.800 ;
        RECT 468.830 2787.520 469.110 2787.800 ;
        RECT 475.730 2787.520 476.010 2787.800 ;
        RECT 482.630 2787.520 482.910 2787.800 ;
        RECT 489.530 2787.520 489.810 2787.800 ;
        RECT 496.430 2787.520 496.710 2787.800 ;
        RECT 509.310 2792.960 509.590 2793.240 ;
        RECT 510.230 2793.640 510.510 2793.920 ;
        RECT 531.390 2793.640 531.670 2793.920 ;
        RECT 542.890 2793.640 543.170 2793.920 ;
        RECT 938.490 3230.880 938.770 3231.160 ;
        RECT 696.990 2948.000 697.270 2948.280 ;
        RECT 938.490 3224.080 938.770 3224.360 ;
        RECT 938.490 3215.920 938.770 3216.200 ;
        RECT 938.490 3209.800 938.770 3210.080 ;
        RECT 792.670 2714.760 792.950 2715.040 ;
        RECT 938.490 3201.640 938.770 3201.920 ;
        RECT 941.710 3196.200 941.990 3196.480 ;
        RECT 938.490 2898.360 938.770 2898.640 ;
        RECT 942.170 3188.040 942.450 3188.320 ;
        RECT 944.930 2891.560 945.210 2891.840 ;
        RECT 1332.250 3249.240 1332.530 3249.520 ;
        RECT 1345.590 2946.640 1345.870 2946.920 ;
        RECT 1345.590 2938.480 1345.870 2938.760 ;
        RECT 1350.190 2904.480 1350.470 2904.760 ;
        RECT 1055.330 2799.760 1055.610 2800.040 ;
        RECT 1052.110 2799.080 1052.390 2799.360 ;
        RECT 1013.930 2794.320 1014.210 2794.600 ;
        RECT 1020.830 2794.320 1021.110 2794.600 ;
        RECT 1027.730 2794.320 1028.010 2794.600 ;
        RECT 979.890 2793.640 980.170 2793.920 ;
        RECT 1007.490 2793.640 1007.770 2793.920 ;
        RECT 1010.710 2793.640 1010.990 2793.920 ;
        RECT 986.790 2792.960 987.070 2793.240 ;
        RECT 993.690 2792.280 993.970 2792.560 ;
        RECT 1001.050 2792.280 1001.330 2792.560 ;
        RECT 1017.610 2792.960 1017.890 2793.240 ;
        RECT 1024.510 2793.640 1024.790 2793.920 ;
        RECT 1045.210 2792.960 1045.490 2793.240 ;
        RECT 1031.410 2790.240 1031.690 2790.520 ;
        RECT 1034.630 2787.520 1034.910 2787.800 ;
        RECT 1038.310 2788.200 1038.590 2788.480 ;
        RECT 1046.130 2788.200 1046.410 2788.480 ;
        RECT 1041.530 2787.520 1041.810 2787.800 ;
        RECT 1048.430 2787.520 1048.710 2787.800 ;
        RECT 1054.870 2788.200 1055.150 2788.480 ;
        RECT 1059.470 2794.320 1059.750 2794.600 ;
        RECT 1065.910 2794.320 1066.190 2794.600 ;
        RECT 1069.590 2794.320 1069.870 2794.600 ;
        RECT 1082.930 2794.320 1083.210 2794.600 ;
        RECT 1087.990 2794.320 1088.270 2794.600 ;
        RECT 1089.370 2794.320 1089.650 2794.600 ;
        RECT 1094.430 2794.320 1094.710 2794.600 ;
        RECT 1096.730 2794.320 1097.010 2794.600 ;
        RECT 1100.410 2794.320 1100.690 2794.600 ;
        RECT 1103.630 2794.320 1103.910 2794.600 ;
        RECT 1105.470 2794.320 1105.750 2794.600 ;
        RECT 1110.530 2794.320 1110.810 2794.600 ;
        RECT 1111.450 2794.320 1111.730 2794.600 ;
        RECT 1117.430 2794.320 1117.710 2794.600 ;
        RECT 1124.330 2794.320 1124.610 2794.600 ;
        RECT 1128.930 2794.320 1129.210 2794.600 ;
        RECT 1131.230 2794.320 1131.510 2794.600 ;
        RECT 1135.830 2794.320 1136.110 2794.600 ;
        RECT 1138.130 2794.320 1138.410 2794.600 ;
        RECT 1145.030 2794.320 1145.310 2794.600 ;
        RECT 1147.330 2794.320 1147.610 2794.600 ;
        RECT 1151.930 2794.320 1152.210 2794.600 ;
        RECT 1158.830 2794.320 1159.110 2794.600 ;
        RECT 1159.750 2794.320 1160.030 2794.600 ;
        RECT 1165.730 2794.320 1166.010 2794.600 ;
        RECT 1172.630 2794.320 1172.910 2794.600 ;
        RECT 1179.530 2794.320 1179.810 2794.600 ;
        RECT 1186.430 2794.320 1186.710 2794.600 ;
        RECT 1200.230 2794.320 1200.510 2794.600 ;
        RECT 1076.490 2793.640 1076.770 2793.920 ;
        RECT 1062.230 2787.520 1062.510 2787.800 ;
        RECT 1069.130 2787.520 1069.410 2787.800 ;
        RECT 1076.030 2787.520 1076.310 2787.800 ;
        RECT 1056.250 2752.840 1056.530 2753.120 ;
        RECT 1057.170 2752.840 1057.450 2753.120 ;
        RECT 1083.850 2793.640 1084.130 2793.920 ;
        RECT 1089.830 2793.640 1090.110 2793.920 ;
        RECT 1117.890 2793.640 1118.170 2793.920 ;
        RECT 1122.030 2793.640 1122.310 2793.920 ;
        RECT 1130.770 2793.640 1131.050 2793.920 ;
        RECT 1138.590 2793.640 1138.870 2793.920 ;
        RECT 1152.390 2792.960 1152.670 2793.240 ;
        RECT 1165.270 2793.640 1165.550 2793.920 ;
        RECT 1159.290 2792.960 1159.570 2793.240 ;
        RECT 1166.190 2793.640 1166.470 2793.920 ;
        RECT 1173.090 2792.960 1173.370 2793.240 ;
        RECT 1179.990 2793.640 1180.270 2793.920 ;
        RECT 1186.890 2792.280 1187.170 2792.560 ;
        RECT 1193.790 2792.280 1194.070 2792.560 ;
        RECT 1193.330 2790.240 1193.610 2790.520 ;
        RECT 1536.950 3230.200 1537.230 3230.480 ;
        RECT 1407.690 1516.600 1407.970 1516.880 ;
        RECT 1408.610 2694.360 1408.890 2694.640 ;
        RECT 1414.130 2683.480 1414.410 2683.760 ;
        RECT 1414.130 2672.600 1414.410 2672.880 ;
        RECT 1414.130 2661.720 1414.410 2662.000 ;
        RECT 1414.130 2650.840 1414.410 2651.120 ;
        RECT 1414.130 2639.280 1414.410 2639.560 ;
        RECT 1414.130 2628.400 1414.410 2628.680 ;
        RECT 1414.130 2617.520 1414.410 2617.800 ;
        RECT 1414.130 2606.640 1414.410 2606.920 ;
        RECT 1414.130 2595.760 1414.410 2596.040 ;
        RECT 1409.530 2584.200 1409.810 2584.480 ;
        RECT 1414.130 2573.320 1414.410 2573.600 ;
        RECT 1410.450 2562.440 1410.730 2562.720 ;
        RECT 1414.130 2551.560 1414.410 2551.840 ;
        RECT 1411.370 2540.680 1411.650 2540.960 ;
        RECT 1409.530 2529.120 1409.810 2529.400 ;
        RECT 1414.130 2518.240 1414.410 2518.520 ;
        RECT 1410.450 2507.360 1410.730 2507.640 ;
        RECT 1414.130 2496.480 1414.410 2496.760 ;
        RECT 1411.370 2485.600 1411.650 2485.880 ;
        RECT 1409.530 2474.040 1409.810 2474.320 ;
        RECT 1412.290 2463.160 1412.570 2463.440 ;
        RECT 1410.450 2452.280 1410.730 2452.560 ;
        RECT 1414.130 2441.400 1414.410 2441.680 ;
        RECT 1414.130 2430.520 1414.410 2430.800 ;
        RECT 1414.130 2418.960 1414.410 2419.240 ;
        RECT 1412.290 2408.080 1412.570 2408.360 ;
        RECT 1410.450 2397.200 1410.730 2397.480 ;
        RECT 1414.130 2386.320 1414.410 2386.600 ;
        RECT 1412.750 2375.440 1413.030 2375.720 ;
        RECT 1410.450 2364.560 1410.730 2364.840 ;
        RECT 1412.290 2353.000 1412.570 2353.280 ;
        RECT 1410.450 2342.120 1410.730 2342.400 ;
        RECT 1414.130 2331.240 1414.410 2331.520 ;
        RECT 1411.370 2320.360 1411.650 2320.640 ;
        RECT 1414.130 2309.480 1414.410 2309.760 ;
        RECT 1412.290 2297.920 1412.570 2298.200 ;
        RECT 1410.450 2287.040 1410.730 2287.320 ;
        RECT 1414.130 2276.160 1414.410 2276.440 ;
        RECT 1414.130 2265.280 1414.410 2265.560 ;
        RECT 1414.130 2254.400 1414.410 2254.680 ;
        RECT 1412.290 2242.840 1412.570 2243.120 ;
        RECT 1414.130 2231.960 1414.410 2232.240 ;
        RECT 1414.130 2221.080 1414.410 2221.360 ;
        RECT 1414.130 2210.200 1414.410 2210.480 ;
        RECT 1414.130 2199.320 1414.410 2199.600 ;
        RECT 1412.290 2187.760 1412.570 2188.040 ;
        RECT 1414.130 2176.880 1414.410 2177.160 ;
        RECT 1414.130 2166.000 1414.410 2166.280 ;
        RECT 1414.130 2155.120 1414.410 2155.400 ;
        RECT 1414.130 2144.240 1414.410 2144.520 ;
        RECT 1414.130 2132.680 1414.410 2132.960 ;
        RECT 1412.290 2121.800 1412.570 2122.080 ;
        RECT 1410.450 2110.920 1410.730 2111.200 ;
        RECT 1408.610 2100.040 1408.890 2100.320 ;
        RECT 1414.130 2089.160 1414.410 2089.440 ;
        RECT 1414.130 2078.280 1414.410 2078.560 ;
        RECT 1409.530 2066.720 1409.810 2067.000 ;
        RECT 1414.130 2055.840 1414.410 2056.120 ;
        RECT 1410.450 2044.960 1410.730 2045.240 ;
        RECT 1414.130 2034.080 1414.410 2034.360 ;
        RECT 1414.130 2023.200 1414.410 2023.480 ;
        RECT 1409.530 2011.640 1409.810 2011.920 ;
        RECT 1414.130 2000.760 1414.410 2001.040 ;
        RECT 1410.450 1989.880 1410.730 1990.160 ;
        RECT 1410.450 1979.000 1410.730 1979.280 ;
        RECT 1411.370 1968.120 1411.650 1968.400 ;
        RECT 1409.530 1956.560 1409.810 1956.840 ;
        RECT 1412.290 1945.680 1412.570 1945.960 ;
        RECT 1410.450 1934.800 1410.730 1935.080 ;
        RECT 1414.130 1923.920 1414.410 1924.200 ;
        RECT 1414.130 1913.040 1414.410 1913.320 ;
        RECT 1414.130 1901.480 1414.410 1901.760 ;
        RECT 1412.290 1890.600 1412.570 1890.880 ;
        RECT 1410.450 1879.720 1410.730 1880.000 ;
        RECT 1414.130 1868.840 1414.410 1869.120 ;
        RECT 1412.750 1857.960 1413.030 1858.240 ;
        RECT 1414.130 1846.400 1414.410 1846.680 ;
        RECT 1412.290 1835.520 1412.570 1835.800 ;
        RECT 1410.450 1824.640 1410.730 1824.920 ;
        RECT 1414.130 1813.760 1414.410 1814.040 ;
        RECT 1412.750 1802.880 1413.030 1803.160 ;
        RECT 1414.130 1792.000 1414.410 1792.280 ;
        RECT 1412.290 1780.440 1412.570 1780.720 ;
        RECT 1410.450 1769.560 1410.730 1769.840 ;
        RECT 1414.130 1758.680 1414.410 1758.960 ;
        RECT 1412.750 1747.800 1413.030 1748.080 ;
        RECT 1414.130 1736.920 1414.410 1737.200 ;
        RECT 1412.290 1725.360 1412.570 1725.640 ;
        RECT 1414.130 1714.480 1414.410 1714.760 ;
        RECT 1414.130 1703.600 1414.410 1703.880 ;
        RECT 1414.130 1692.720 1414.410 1693.000 ;
        RECT 1414.130 1681.840 1414.410 1682.120 ;
        RECT 1411.830 1670.280 1412.110 1670.560 ;
        RECT 1414.130 1659.400 1414.410 1659.680 ;
        RECT 1414.130 1648.520 1414.410 1648.800 ;
        RECT 1414.130 1637.640 1414.410 1637.920 ;
        RECT 1414.130 1626.760 1414.410 1627.040 ;
        RECT 1411.830 1615.200 1412.110 1615.480 ;
        RECT 1414.130 1604.320 1414.410 1604.600 ;
        RECT 1535.570 3224.760 1535.850 3225.040 ;
        RECT 1535.570 3217.280 1535.850 3217.560 ;
        RECT 1538.330 3210.480 1538.610 3210.760 ;
        RECT 1538.330 3202.320 1538.610 3202.600 ;
        RECT 1533.270 3196.880 1533.550 3197.160 ;
        RECT 1497.850 3189.400 1498.130 3189.680 ;
        RECT 1534.650 2899.720 1534.930 2900.000 ;
        RECT 1531.890 2891.560 1532.170 2891.840 ;
        RECT 1945.890 3249.240 1946.170 3249.520 ;
        RECT 1739.810 2796.360 1740.090 2796.640 ;
        RECT 1788.570 2796.360 1788.850 2796.640 ;
        RECT 1580.190 2794.320 1580.470 2794.600 ;
        RECT 1593.990 2794.320 1594.270 2794.600 ;
        RECT 1601.350 2794.320 1601.630 2794.600 ;
        RECT 1607.790 2794.320 1608.070 2794.600 ;
        RECT 1617.910 2794.320 1618.190 2794.600 ;
        RECT 1628.490 2794.320 1628.770 2794.600 ;
        RECT 1635.390 2794.320 1635.670 2794.600 ;
        RECT 1649.650 2794.320 1649.930 2794.600 ;
        RECT 1658.850 2794.320 1659.130 2794.600 ;
        RECT 1662.990 2794.320 1663.270 2794.600 ;
        RECT 1669.890 2794.320 1670.170 2794.600 ;
        RECT 1676.790 2794.320 1677.070 2794.600 ;
        RECT 1414.130 1593.440 1414.410 1593.720 ;
        RECT 1414.130 1582.560 1414.410 1582.840 ;
        RECT 1414.130 1571.680 1414.410 1571.960 ;
        RECT 1411.830 1560.120 1412.110 1560.400 ;
        RECT 1409.530 1549.240 1409.810 1549.520 ;
        RECT 1587.090 2792.280 1587.370 2792.560 ;
        RECT 1600.890 2788.880 1601.170 2789.160 ;
        RECT 1414.130 1538.360 1414.410 1538.640 ;
        RECT 1611.470 2793.640 1611.750 2793.920 ;
        RECT 1614.690 2789.560 1614.970 2789.840 ;
        RECT 1618.370 2792.960 1618.650 2793.240 ;
        RECT 1624.810 2792.960 1625.090 2793.240 ;
        RECT 1631.710 2792.960 1631.990 2793.240 ;
        RECT 1638.610 2793.640 1638.890 2793.920 ;
        RECT 1645.510 2793.640 1645.790 2793.920 ;
        RECT 1642.290 2790.920 1642.570 2791.200 ;
        RECT 1646.430 2792.960 1646.710 2793.240 ;
        RECT 1649.190 2791.600 1649.470 2791.880 ;
        RECT 1652.410 2792.960 1652.690 2793.240 ;
        RECT 1656.090 2790.920 1656.370 2791.200 ;
        RECT 1663.450 2793.640 1663.730 2793.920 ;
        RECT 1670.350 2793.640 1670.630 2793.920 ;
        RECT 1683.690 2794.320 1683.970 2794.600 ;
        RECT 1686.910 2794.320 1687.190 2794.600 ;
        RECT 1690.590 2794.320 1690.870 2794.600 ;
        RECT 1697.490 2794.320 1697.770 2794.600 ;
        RECT 1704.390 2794.320 1704.670 2794.600 ;
        RECT 1711.290 2794.320 1711.570 2794.600 ;
        RECT 1718.190 2794.320 1718.470 2794.600 ;
        RECT 1721.410 2794.320 1721.690 2794.600 ;
        RECT 1725.090 2794.320 1725.370 2794.600 ;
        RECT 1731.990 2794.320 1732.270 2794.600 ;
        RECT 1738.890 2794.320 1739.170 2794.600 ;
        RECT 1677.250 2793.640 1677.530 2793.920 ;
        RECT 1683.230 2793.640 1683.510 2793.920 ;
        RECT 1684.150 2792.280 1684.430 2792.560 ;
        RECT 1694.730 2793.640 1695.010 2793.920 ;
        RECT 1699.330 2793.640 1699.610 2793.920 ;
        RECT 1704.850 2793.640 1705.130 2793.920 ;
        RECT 1712.670 2793.640 1712.950 2793.920 ;
        RECT 1718.650 2793.640 1718.930 2793.920 ;
        RECT 1718.650 2788.200 1718.930 2788.480 ;
        RECT 1731.530 2793.640 1731.810 2793.920 ;
        RECT 1734.750 2793.640 1735.030 2793.920 ;
        RECT 1745.790 2794.320 1746.070 2794.600 ;
        RECT 1759.590 2794.320 1759.870 2794.600 ;
        RECT 1741.650 2793.640 1741.930 2793.920 ;
        RECT 1747.630 2793.640 1747.910 2793.920 ;
        RECT 1766.490 2793.640 1766.770 2793.920 ;
        RECT 1752.690 2792.280 1752.970 2792.560 ;
        RECT 1773.390 2791.600 1773.670 2791.880 ;
        RECT 1760.050 2788.200 1760.330 2788.480 ;
        RECT 1752.690 2787.520 1752.970 2787.800 ;
        RECT 1760.970 2777.320 1761.250 2777.600 ;
        RECT 1766.490 2787.520 1766.770 2787.800 ;
        RECT 1773.850 2787.520 1774.130 2787.800 ;
        RECT 1787.190 2793.640 1787.470 2793.920 ;
        RECT 1780.290 2792.960 1780.570 2793.240 ;
        RECT 1780.290 2787.520 1780.570 2787.800 ;
        RECT 1787.190 2787.520 1787.470 2787.800 ;
        RECT 1794.090 2777.320 1794.370 2777.600 ;
        RECT 2187.390 3230.880 2187.670 3231.160 ;
        RECT 1945.890 2948.000 1946.170 2948.280 ;
        RECT 2187.390 3224.080 2187.670 3224.360 ;
        RECT 2187.390 3215.920 2187.670 3216.200 ;
        RECT 2187.390 3209.800 2187.670 3210.080 ;
        RECT 2187.390 3201.640 2187.670 3201.920 ;
        RECT 2187.390 3196.200 2187.670 3196.480 ;
        RECT 2187.390 3188.040 2187.670 3188.320 ;
        RECT 2187.390 2898.360 2187.670 2898.640 ;
        RECT 2190.610 2891.560 2190.890 2891.840 ;
        RECT 2582.070 3249.240 2582.350 3249.520 ;
        RECT 2594.490 2946.640 2594.770 2946.920 ;
        RECT 2594.490 2938.480 2594.770 2938.760 ;
        RECT 2228.790 2794.320 2229.070 2794.600 ;
        RECT 2232.010 2794.320 2232.290 2794.600 ;
        RECT 2238.910 2794.320 2239.190 2794.600 ;
        RECT 2245.810 2794.320 2246.090 2794.600 ;
        RECT 2263.750 2794.320 2264.030 2794.600 ;
        RECT 2267.430 2794.320 2267.710 2794.600 ;
        RECT 2273.410 2794.320 2273.690 2794.600 ;
        RECT 2294.110 2794.320 2294.390 2794.600 ;
        RECT 2304.690 2794.320 2304.970 2794.600 ;
        RECT 2308.830 2794.320 2309.110 2794.600 ;
        RECT 2311.590 2794.320 2311.870 2794.600 ;
        RECT 2318.490 2794.320 2318.770 2794.600 ;
        RECT 2325.390 2794.320 2325.670 2794.600 ;
        RECT 2332.290 2794.320 2332.570 2794.600 ;
        RECT 2339.190 2794.320 2339.470 2794.600 ;
        RECT 2342.870 2794.320 2343.150 2794.600 ;
        RECT 2346.090 2794.320 2346.370 2794.600 ;
        RECT 2352.990 2794.320 2353.270 2794.600 ;
        RECT 2359.890 2794.320 2360.170 2794.600 ;
        RECT 2366.790 2794.320 2367.070 2794.600 ;
        RECT 2373.690 2794.320 2373.970 2794.600 ;
        RECT 2381.050 2794.320 2381.330 2794.600 ;
        RECT 2385.650 2794.320 2385.930 2794.600 ;
        RECT 2391.630 2794.320 2391.910 2794.600 ;
        RECT 2397.150 2794.320 2397.430 2794.600 ;
        RECT 2402.670 2794.320 2402.950 2794.600 ;
        RECT 2415.090 2794.320 2415.370 2794.600 ;
        RECT 2422.450 2794.320 2422.730 2794.600 ;
        RECT 2428.890 2794.320 2429.170 2794.600 ;
        RECT 2263.290 2790.920 2263.570 2791.200 ;
        RECT 2256.850 2788.200 2257.130 2788.480 ;
        RECT 2266.510 2793.640 2266.790 2793.920 ;
        RECT 2270.190 2791.600 2270.470 2791.880 ;
        RECT 2280.310 2792.960 2280.590 2793.240 ;
        RECT 2287.210 2792.960 2287.490 2793.240 ;
        RECT 2277.090 2792.280 2277.370 2792.560 ;
        RECT 2283.990 2791.600 2284.270 2791.880 ;
        RECT 2290.890 2791.600 2291.170 2791.880 ;
        RECT 2301.010 2793.640 2301.290 2793.920 ;
        RECT 2303.310 2793.640 2303.590 2793.920 ;
        RECT 2297.790 2790.920 2298.070 2791.200 ;
        RECT 2304.230 2792.960 2304.510 2793.240 ;
        RECT 2305.150 2793.640 2305.430 2793.920 ;
        RECT 2314.810 2793.640 2315.090 2793.920 ;
        RECT 2321.710 2793.640 2321.990 2793.920 ;
        RECT 2325.850 2793.640 2326.130 2793.920 ;
        RECT 2332.750 2792.960 2333.030 2793.240 ;
        RECT 2339.650 2793.640 2339.930 2793.920 ;
        RECT 2340.110 2792.960 2340.390 2793.240 ;
        RECT 2350.230 2793.640 2350.510 2793.920 ;
        RECT 2356.210 2793.640 2356.490 2793.920 ;
        RECT 2361.270 2793.640 2361.550 2793.920 ;
        RECT 2367.710 2793.640 2367.990 2793.920 ;
        RECT 2373.230 2788.200 2373.510 2788.480 ;
        RECT 2374.150 2793.640 2374.430 2793.920 ;
        RECT 2377.830 2793.640 2378.110 2793.920 ;
        RECT 2380.590 2790.240 2380.870 2790.520 ;
        RECT 2402.210 2793.640 2402.490 2793.920 ;
        RECT 2387.490 2790.240 2387.770 2790.520 ;
        RECT 2394.390 2789.560 2394.670 2789.840 ;
        RECT 2421.990 2793.640 2422.270 2793.920 ;
        RECT 2415.090 2792.960 2415.370 2793.240 ;
        RECT 2442.690 2792.960 2442.970 2793.240 ;
        RECT 2408.190 2792.280 2408.470 2792.560 ;
        RECT 2435.790 2792.280 2436.070 2792.560 ;
        RECT 2442.690 2791.600 2442.970 2791.880 ;
        RECT 2415.090 2790.920 2415.370 2791.200 ;
        RECT 2428.890 2790.920 2429.170 2791.200 ;
        RECT 2435.790 2790.920 2436.070 2791.200 ;
        RECT 2408.190 2788.880 2408.470 2789.160 ;
        RECT 2415.090 2788.200 2415.370 2788.480 ;
        RECT 1410.450 1527.480 1410.730 1527.760 ;
        RECT 1408.150 1505.720 1408.430 1506.000 ;
      LAYER met3 ;
        RECT 646.365 3264.500 646.695 3264.505 ;
        RECT 646.110 3264.490 646.695 3264.500 ;
        RECT 645.910 3264.190 646.695 3264.490 ;
        RECT 646.110 3264.180 646.695 3264.190 ;
        RECT 646.365 3264.175 646.695 3264.180 ;
        RECT 667.985 3264.500 668.315 3264.505 ;
        RECT 1295.885 3264.500 1296.215 3264.505 ;
        RECT 1318.885 3264.500 1319.215 3264.505 ;
        RECT 667.985 3264.490 668.570 3264.500 ;
        RECT 1295.630 3264.490 1296.215 3264.500 ;
        RECT 1318.630 3264.490 1319.215 3264.500 ;
        RECT 667.985 3264.190 668.770 3264.490 ;
        RECT 1295.430 3264.190 1296.215 3264.490 ;
        RECT 1318.430 3264.190 1319.215 3264.490 ;
        RECT 667.985 3264.180 668.570 3264.190 ;
        RECT 1295.630 3264.180 1296.215 3264.190 ;
        RECT 1318.630 3264.180 1319.215 3264.190 ;
        RECT 667.985 3264.175 668.315 3264.180 ;
        RECT 1295.885 3264.175 1296.215 3264.180 ;
        RECT 1318.885 3264.175 1319.215 3264.180 ;
        RECT 1892.505 3264.500 1892.835 3264.505 ;
        RECT 1917.345 3264.500 1917.675 3264.505 ;
        RECT 2539.265 3264.500 2539.595 3264.505 ;
        RECT 2566.865 3264.500 2567.195 3264.505 ;
        RECT 1892.505 3264.490 1893.090 3264.500 ;
        RECT 1917.345 3264.490 1917.930 3264.500 ;
        RECT 2539.265 3264.490 2539.850 3264.500 ;
        RECT 2566.865 3264.490 2567.450 3264.500 ;
        RECT 1892.505 3264.190 1893.290 3264.490 ;
        RECT 1917.345 3264.190 1918.130 3264.490 ;
        RECT 2539.265 3264.190 2540.050 3264.490 ;
        RECT 2566.865 3264.190 2567.650 3264.490 ;
        RECT 1892.505 3264.180 1893.090 3264.190 ;
        RECT 1917.345 3264.180 1917.930 3264.190 ;
        RECT 2539.265 3264.180 2539.850 3264.190 ;
        RECT 2566.865 3264.180 2567.450 3264.190 ;
        RECT 1892.505 3264.175 1892.835 3264.180 ;
        RECT 1917.345 3264.175 1917.675 3264.180 ;
        RECT 2539.265 3264.175 2539.595 3264.180 ;
        RECT 2566.865 3264.175 2567.195 3264.180 ;
        RECT 659.280 3251.235 661.020 3252.140 ;
        RECT 1309.280 3251.235 1311.020 3252.140 ;
        RECT 1909.280 3251.235 1911.020 3252.140 ;
        RECT 2559.280 3251.235 2561.020 3252.140 ;
        RECT 300.000 3232.785 304.600 3233.085 ;
        RECT 282.965 3230.490 283.295 3230.505 ;
        RECT 300.230 3230.490 300.530 3232.785 ;
        RECT 282.965 3230.190 300.530 3230.490 ;
        RECT 282.965 3230.175 283.295 3230.190 ;
        RECT 300.000 3227.145 304.600 3227.445 ;
        RECT 286.185 3225.050 286.515 3225.065 ;
        RECT 300.230 3225.050 300.530 3227.145 ;
        RECT 286.185 3224.750 300.530 3225.050 ;
        RECT 286.185 3224.735 286.515 3224.750 ;
        RECT 300.000 3218.645 304.600 3218.945 ;
        RECT 285.725 3216.210 286.055 3216.225 ;
        RECT 300.230 3216.210 300.530 3218.645 ;
        RECT 285.725 3215.910 300.530 3216.210 ;
        RECT 285.725 3215.895 286.055 3215.910 ;
        RECT 300.000 3213.005 304.600 3213.305 ;
        RECT 285.265 3210.090 285.595 3210.105 ;
        RECT 300.230 3210.090 300.530 3213.005 ;
        RECT 285.265 3209.790 300.530 3210.090 ;
        RECT 285.265 3209.775 285.595 3209.790 ;
        RECT 300.000 3204.505 304.600 3204.805 ;
        RECT 284.805 3201.930 285.135 3201.945 ;
        RECT 300.230 3201.930 300.530 3204.505 ;
        RECT 284.805 3201.630 300.530 3201.930 ;
        RECT 284.805 3201.615 285.135 3201.630 ;
        RECT 300.000 3198.865 304.600 3199.165 ;
        RECT 284.345 3196.490 284.675 3196.505 ;
        RECT 300.230 3196.490 300.530 3198.865 ;
        RECT 284.345 3196.190 300.530 3196.490 ;
        RECT 284.345 3196.175 284.675 3196.190 ;
        RECT 300.000 3190.365 304.600 3190.665 ;
        RECT 283.885 3188.330 284.215 3188.345 ;
        RECT 300.230 3188.330 300.530 3190.365 ;
        RECT 283.885 3188.030 300.530 3188.330 ;
        RECT 283.885 3188.015 284.215 3188.030 ;
        RECT 300.000 2901.125 304.600 2901.425 ;
        RECT 283.425 2898.650 283.755 2898.665 ;
        RECT 300.230 2898.650 300.530 2901.125 ;
        RECT 283.425 2898.350 300.530 2898.650 ;
        RECT 283.425 2898.335 283.755 2898.350 ;
        RECT 298.145 2892.925 298.475 2892.940 ;
        RECT 298.145 2892.625 304.600 2892.925 ;
        RECT 298.145 2892.610 298.475 2892.625 ;
      LAYER met3 ;
        RECT 305.000 2805.000 681.480 3251.235 ;
      LAYER met3 ;
        RECT 696.965 3249.530 697.295 3249.545 ;
        RECT 685.710 3249.230 697.295 3249.530 ;
        RECT 685.710 3248.565 686.010 3249.230 ;
        RECT 696.965 3249.215 697.295 3249.230 ;
        RECT 681.880 3248.265 686.480 3248.565 ;
        RECT 950.000 3232.785 954.600 3233.085 ;
        RECT 938.465 3231.170 938.795 3231.185 ;
        RECT 950.670 3231.170 950.970 3232.785 ;
        RECT 938.465 3230.870 950.970 3231.170 ;
        RECT 938.465 3230.855 938.795 3230.870 ;
        RECT 950.000 3227.145 954.600 3227.445 ;
        RECT 938.465 3224.370 938.795 3224.385 ;
        RECT 950.670 3224.370 950.970 3227.145 ;
        RECT 938.465 3224.070 950.970 3224.370 ;
        RECT 938.465 3224.055 938.795 3224.070 ;
        RECT 950.000 3218.645 954.600 3218.945 ;
        RECT 938.465 3216.210 938.795 3216.225 ;
        RECT 950.670 3216.210 950.970 3218.645 ;
        RECT 938.465 3215.910 950.970 3216.210 ;
        RECT 938.465 3215.895 938.795 3215.910 ;
        RECT 950.000 3213.005 954.600 3213.305 ;
        RECT 938.465 3210.090 938.795 3210.105 ;
        RECT 950.670 3210.090 950.970 3213.005 ;
        RECT 938.465 3209.790 950.970 3210.090 ;
        RECT 938.465 3209.775 938.795 3209.790 ;
        RECT 950.000 3204.505 954.600 3204.805 ;
        RECT 938.465 3201.930 938.795 3201.945 ;
        RECT 950.670 3201.930 950.970 3204.505 ;
        RECT 938.465 3201.630 950.970 3201.930 ;
        RECT 938.465 3201.615 938.795 3201.630 ;
        RECT 950.000 3198.865 954.600 3199.165 ;
        RECT 941.685 3196.490 942.015 3196.505 ;
        RECT 950.670 3196.490 950.970 3198.865 ;
        RECT 941.685 3196.190 950.970 3196.490 ;
        RECT 941.685 3196.175 942.015 3196.190 ;
        RECT 950.000 3190.365 954.600 3190.665 ;
        RECT 942.145 3188.330 942.475 3188.345 ;
        RECT 950.670 3188.330 950.970 3190.365 ;
        RECT 942.145 3188.030 950.970 3188.330 ;
        RECT 942.145 3188.015 942.475 3188.030 ;
        RECT 696.965 2948.290 697.295 2948.305 ;
        RECT 684.790 2947.990 697.295 2948.290 ;
        RECT 684.790 2947.210 685.090 2947.990 ;
        RECT 696.965 2947.975 697.295 2947.990 ;
        RECT 681.880 2946.910 686.480 2947.210 ;
        RECT 684.790 2938.710 685.090 2946.910 ;
        RECT 681.880 2938.410 686.480 2938.710 ;
        RECT 684.790 2933.070 685.090 2938.410 ;
        RECT 681.880 2932.770 686.480 2933.070 ;
        RECT 685.710 2924.570 686.010 2932.770 ;
        RECT 681.880 2924.270 686.480 2924.570 ;
        RECT 685.710 2918.930 686.010 2924.270 ;
        RECT 681.880 2918.630 686.480 2918.930 ;
        RECT 685.710 2910.430 686.010 2918.630 ;
        RECT 681.880 2910.130 686.480 2910.430 ;
        RECT 685.710 2904.790 686.010 2910.130 ;
        RECT 681.880 2904.490 686.480 2904.790 ;
        RECT 950.000 2901.125 954.600 2901.425 ;
        RECT 938.465 2898.650 938.795 2898.665 ;
        RECT 950.670 2898.650 950.970 2901.125 ;
        RECT 938.465 2898.350 950.970 2898.650 ;
        RECT 938.465 2898.335 938.795 2898.350 ;
        RECT 950.000 2892.625 954.600 2892.925 ;
        RECT 944.905 2891.850 945.235 2891.865 ;
        RECT 950.670 2891.850 950.970 2892.625 ;
        RECT 944.905 2891.550 950.970 2891.850 ;
        RECT 944.905 2891.535 945.235 2891.550 ;
      LAYER met3 ;
        RECT 955.000 2805.000 1331.480 3251.235 ;
      LAYER met3 ;
        RECT 1332.225 3249.530 1332.555 3249.545 ;
        RECT 1332.225 3249.215 1332.770 3249.530 ;
        RECT 1332.470 3248.565 1332.770 3249.215 ;
        RECT 1331.880 3248.265 1336.480 3248.565 ;
        RECT 1550.000 3232.785 1554.600 3233.085 ;
        RECT 1536.925 3230.490 1537.255 3230.505 ;
        RECT 1550.510 3230.490 1550.810 3232.785 ;
        RECT 1536.925 3230.190 1550.810 3230.490 ;
        RECT 1536.925 3230.175 1537.255 3230.190 ;
        RECT 1550.000 3227.145 1554.600 3227.445 ;
        RECT 1535.545 3225.050 1535.875 3225.065 ;
        RECT 1550.510 3225.050 1550.810 3227.145 ;
        RECT 1535.545 3224.750 1550.810 3225.050 ;
        RECT 1535.545 3224.735 1535.875 3224.750 ;
        RECT 1550.000 3218.645 1554.600 3218.945 ;
        RECT 1535.545 3217.570 1535.875 3217.585 ;
        RECT 1550.510 3217.570 1550.810 3218.645 ;
        RECT 1535.545 3217.270 1550.810 3217.570 ;
        RECT 1535.545 3217.255 1535.875 3217.270 ;
        RECT 1550.000 3213.005 1554.600 3213.305 ;
        RECT 1538.305 3210.770 1538.635 3210.785 ;
        RECT 1550.510 3210.770 1550.810 3213.005 ;
        RECT 1538.305 3210.470 1550.810 3210.770 ;
        RECT 1538.305 3210.455 1538.635 3210.470 ;
        RECT 1550.000 3204.505 1554.600 3204.805 ;
        RECT 1538.305 3202.610 1538.635 3202.625 ;
        RECT 1550.510 3202.610 1550.810 3204.505 ;
        RECT 1538.305 3202.310 1550.810 3202.610 ;
        RECT 1538.305 3202.295 1538.635 3202.310 ;
        RECT 1550.000 3198.865 1554.600 3199.165 ;
        RECT 1533.245 3197.170 1533.575 3197.185 ;
        RECT 1550.510 3197.170 1550.810 3198.865 ;
        RECT 1533.245 3196.870 1550.810 3197.170 ;
        RECT 1533.245 3196.855 1533.575 3196.870 ;
        RECT 1550.000 3190.365 1554.600 3190.665 ;
        RECT 1497.825 3189.690 1498.155 3189.705 ;
        RECT 1550.510 3189.690 1550.810 3190.365 ;
        RECT 1497.825 3189.390 1550.810 3189.690 ;
        RECT 1497.825 3189.375 1498.155 3189.390 ;
        RECT 1331.880 2946.930 1336.480 2947.210 ;
        RECT 1345.565 2946.930 1345.895 2946.945 ;
        RECT 1331.880 2946.910 1345.895 2946.930 ;
        RECT 1336.150 2946.630 1345.895 2946.910 ;
        RECT 1345.565 2946.615 1345.895 2946.630 ;
        RECT 1345.565 2938.770 1345.895 2938.785 ;
        RECT 1336.150 2938.710 1345.895 2938.770 ;
        RECT 1331.880 2938.470 1345.895 2938.710 ;
        RECT 1331.880 2938.410 1336.480 2938.470 ;
        RECT 1345.565 2938.455 1345.895 2938.470 ;
        RECT 1336.150 2933.070 1336.450 2938.410 ;
        RECT 1331.880 2932.770 1336.480 2933.070 ;
        RECT 1336.150 2924.570 1336.450 2932.770 ;
        RECT 1331.880 2924.270 1336.480 2924.570 ;
        RECT 1336.150 2918.930 1336.450 2924.270 ;
        RECT 1331.880 2918.630 1336.480 2918.930 ;
        RECT 1336.150 2910.430 1336.450 2918.630 ;
        RECT 1331.880 2910.130 1336.480 2910.430 ;
        RECT 1336.150 2904.790 1336.450 2910.130 ;
        RECT 1331.880 2904.770 1336.480 2904.790 ;
        RECT 1350.165 2904.770 1350.495 2904.785 ;
        RECT 1331.880 2904.490 1350.495 2904.770 ;
        RECT 1336.150 2904.470 1350.495 2904.490 ;
        RECT 1350.165 2904.455 1350.495 2904.470 ;
        RECT 1550.000 2901.125 1554.600 2901.425 ;
        RECT 1534.625 2900.010 1534.955 2900.025 ;
        RECT 1550.510 2900.010 1550.810 2901.125 ;
        RECT 1534.625 2899.710 1550.810 2900.010 ;
        RECT 1534.625 2899.695 1534.955 2899.710 ;
        RECT 1550.000 2892.625 1554.600 2892.925 ;
        RECT 1531.865 2891.850 1532.195 2891.865 ;
        RECT 1550.510 2891.850 1550.810 2892.625 ;
        RECT 1531.865 2891.550 1550.810 2891.850 ;
        RECT 1531.865 2891.535 1532.195 2891.550 ;
      LAYER met3 ;
        RECT 1555.000 2805.000 1931.480 3251.235 ;
      LAYER met3 ;
        RECT 1945.865 3249.530 1946.195 3249.545 ;
        RECT 1935.990 3249.230 1946.195 3249.530 ;
        RECT 1935.990 3248.565 1936.290 3249.230 ;
        RECT 1945.865 3249.215 1946.195 3249.230 ;
        RECT 1931.880 3248.265 1936.480 3248.565 ;
        RECT 2200.000 3232.785 2204.600 3233.085 ;
        RECT 2187.365 3231.170 2187.695 3231.185 ;
        RECT 2200.030 3231.170 2200.330 3232.785 ;
        RECT 2187.365 3230.870 2200.330 3231.170 ;
        RECT 2187.365 3230.855 2187.695 3230.870 ;
        RECT 2200.000 3227.145 2204.600 3227.445 ;
        RECT 2187.365 3224.370 2187.695 3224.385 ;
        RECT 2200.030 3224.370 2200.330 3227.145 ;
        RECT 2187.365 3224.070 2200.330 3224.370 ;
        RECT 2187.365 3224.055 2187.695 3224.070 ;
        RECT 2200.000 3218.645 2204.600 3218.945 ;
        RECT 2187.365 3216.210 2187.695 3216.225 ;
        RECT 2200.030 3216.210 2200.330 3218.645 ;
        RECT 2187.365 3215.910 2200.330 3216.210 ;
        RECT 2187.365 3215.895 2187.695 3215.910 ;
        RECT 2200.000 3213.005 2204.600 3213.305 ;
        RECT 2187.365 3210.090 2187.695 3210.105 ;
        RECT 2200.030 3210.090 2200.330 3213.005 ;
        RECT 2187.365 3209.790 2200.330 3210.090 ;
        RECT 2187.365 3209.775 2187.695 3209.790 ;
        RECT 2200.000 3204.505 2204.600 3204.805 ;
        RECT 2187.365 3201.930 2187.695 3201.945 ;
        RECT 2200.030 3201.930 2200.330 3204.505 ;
        RECT 2187.365 3201.630 2200.330 3201.930 ;
        RECT 2187.365 3201.615 2187.695 3201.630 ;
        RECT 2200.000 3198.865 2204.600 3199.165 ;
        RECT 2187.365 3196.490 2187.695 3196.505 ;
        RECT 2200.030 3196.490 2200.330 3198.865 ;
        RECT 2187.365 3196.190 2200.330 3196.490 ;
        RECT 2187.365 3196.175 2187.695 3196.190 ;
        RECT 2200.000 3190.365 2204.600 3190.665 ;
        RECT 2187.365 3188.330 2187.695 3188.345 ;
        RECT 2200.030 3188.330 2200.330 3190.365 ;
        RECT 2187.365 3188.030 2200.330 3188.330 ;
        RECT 2187.365 3188.015 2187.695 3188.030 ;
        RECT 1945.865 2948.290 1946.195 2948.305 ;
        RECT 1935.070 2947.990 1946.195 2948.290 ;
        RECT 1935.070 2947.210 1935.370 2947.990 ;
        RECT 1945.865 2947.975 1946.195 2947.990 ;
        RECT 1931.880 2946.910 1936.480 2947.210 ;
        RECT 1935.070 2938.710 1935.370 2946.910 ;
        RECT 1931.880 2938.410 1936.480 2938.710 ;
        RECT 1935.070 2933.070 1935.370 2938.410 ;
        RECT 1931.880 2932.770 1936.480 2933.070 ;
        RECT 1935.990 2924.570 1936.290 2932.770 ;
        RECT 1931.880 2924.270 1936.480 2924.570 ;
        RECT 1935.990 2918.930 1936.290 2924.270 ;
        RECT 1931.880 2918.630 1936.480 2918.930 ;
        RECT 1935.990 2910.430 1936.290 2918.630 ;
        RECT 1931.880 2910.130 1936.480 2910.430 ;
        RECT 1935.990 2904.790 1936.290 2910.130 ;
        RECT 1931.880 2904.490 1936.480 2904.790 ;
        RECT 2200.000 2901.125 2204.600 2901.425 ;
        RECT 2187.365 2898.650 2187.695 2898.665 ;
        RECT 2200.030 2898.650 2200.330 2901.125 ;
        RECT 2187.365 2898.350 2200.330 2898.650 ;
        RECT 2187.365 2898.335 2187.695 2898.350 ;
        RECT 2200.000 2892.625 2204.600 2892.925 ;
        RECT 2190.585 2891.850 2190.915 2891.865 ;
        RECT 2200.030 2891.850 2200.330 2892.625 ;
        RECT 2190.585 2891.550 2200.330 2891.850 ;
        RECT 2190.585 2891.535 2190.915 2891.550 ;
      LAYER met3 ;
        RECT 2205.000 2805.000 2581.480 3251.235 ;
      LAYER met3 ;
        RECT 2582.045 3249.530 2582.375 3249.545 ;
        RECT 2582.045 3249.230 2583.050 3249.530 ;
        RECT 2582.045 3249.215 2582.375 3249.230 ;
        RECT 2582.750 3248.565 2583.050 3249.230 ;
        RECT 2581.880 3248.265 2586.480 3248.565 ;
        RECT 2581.880 2946.930 2586.480 2947.210 ;
        RECT 2594.465 2946.930 2594.795 2946.945 ;
        RECT 2581.880 2946.910 2594.795 2946.930 ;
        RECT 2585.510 2946.630 2594.795 2946.910 ;
        RECT 2594.465 2946.615 2594.795 2946.630 ;
        RECT 2594.465 2938.770 2594.795 2938.785 ;
        RECT 2585.510 2938.710 2594.795 2938.770 ;
        RECT 2581.880 2938.470 2594.795 2938.710 ;
        RECT 2581.880 2938.410 2586.480 2938.470 ;
        RECT 2594.465 2938.455 2594.795 2938.470 ;
        RECT 2585.510 2933.070 2585.810 2938.410 ;
        RECT 2581.880 2932.770 2586.480 2933.070 ;
        RECT 2585.510 2924.570 2585.810 2932.770 ;
        RECT 2581.880 2924.270 2586.480 2924.570 ;
        RECT 2585.510 2918.930 2585.810 2924.270 ;
        RECT 2581.880 2918.630 2586.480 2918.930 ;
        RECT 2585.510 2910.430 2585.810 2918.630 ;
        RECT 2581.880 2910.130 2586.480 2910.430 ;
        RECT 2585.510 2904.790 2585.810 2910.130 ;
        RECT 2581.880 2904.490 2586.480 2904.790 ;
        RECT 1055.305 2800.060 1055.635 2800.065 ;
        RECT 1055.305 2800.050 1055.890 2800.060 ;
        RECT 1055.305 2799.750 1056.090 2800.050 ;
        RECT 1055.305 2799.740 1055.890 2799.750 ;
        RECT 1055.305 2799.735 1055.635 2799.740 ;
        RECT 1052.085 2799.370 1052.415 2799.385 ;
        RECT 1052.750 2799.370 1053.130 2799.380 ;
        RECT 1052.085 2799.070 1053.130 2799.370 ;
        RECT 1052.085 2799.055 1052.415 2799.070 ;
        RECT 1052.750 2799.060 1053.130 2799.070 ;
        RECT 1739.785 2796.650 1740.115 2796.665 ;
        RECT 1759.310 2796.650 1759.690 2796.660 ;
        RECT 1739.785 2796.350 1759.690 2796.650 ;
        RECT 1739.785 2796.335 1740.115 2796.350 ;
        RECT 1759.310 2796.340 1759.690 2796.350 ;
        RECT 1788.545 2796.650 1788.875 2796.665 ;
        RECT 1794.270 2796.650 1794.650 2796.660 ;
        RECT 1788.545 2796.350 1794.650 2796.650 ;
        RECT 1788.545 2796.335 1788.875 2796.350 ;
        RECT 1794.270 2796.340 1794.650 2796.350 ;
        RECT 336.990 2794.610 337.370 2794.620 ;
        RECT 337.705 2794.610 338.035 2794.625 ;
        RECT 336.990 2794.310 338.035 2794.610 ;
        RECT 336.990 2794.300 337.370 2794.310 ;
        RECT 337.705 2794.295 338.035 2794.310 ;
        RECT 348.950 2794.610 349.330 2794.620 ;
        RECT 350.585 2794.610 350.915 2794.625 ;
        RECT 362.085 2794.620 362.415 2794.625 ;
        RECT 368.525 2794.620 368.855 2794.625 ;
        RECT 361.830 2794.610 362.415 2794.620 ;
        RECT 368.270 2794.610 368.855 2794.620 ;
        RECT 348.950 2794.310 350.915 2794.610 ;
        RECT 361.630 2794.310 362.415 2794.610 ;
        RECT 368.070 2794.310 368.855 2794.610 ;
        RECT 348.950 2794.300 349.330 2794.310 ;
        RECT 350.585 2794.295 350.915 2794.310 ;
        RECT 361.830 2794.300 362.415 2794.310 ;
        RECT 368.270 2794.300 368.855 2794.310 ;
        RECT 374.710 2794.610 375.090 2794.620 ;
        RECT 378.645 2794.610 378.975 2794.625 ;
        RECT 374.710 2794.310 378.975 2794.610 ;
        RECT 374.710 2794.300 375.090 2794.310 ;
        RECT 362.085 2794.295 362.415 2794.300 ;
        RECT 368.525 2794.295 368.855 2794.300 ;
        RECT 378.645 2794.295 378.975 2794.310 ;
        RECT 379.310 2794.610 379.690 2794.620 ;
        RECT 380.025 2794.610 380.355 2794.625 ;
        RECT 386.925 2794.620 387.255 2794.625 ;
        RECT 392.445 2794.620 392.775 2794.625 ;
        RECT 386.670 2794.610 387.255 2794.620 ;
        RECT 392.190 2794.610 392.775 2794.620 ;
        RECT 379.310 2794.310 380.355 2794.610 ;
        RECT 386.470 2794.310 387.255 2794.610 ;
        RECT 391.990 2794.310 392.775 2794.610 ;
        RECT 379.310 2794.300 379.690 2794.310 ;
        RECT 380.025 2794.295 380.355 2794.310 ;
        RECT 386.670 2794.300 387.255 2794.310 ;
        RECT 392.190 2794.300 392.775 2794.310 ;
        RECT 396.790 2794.610 397.170 2794.620 ;
        RECT 397.505 2794.610 397.835 2794.625 ;
        RECT 403.485 2794.620 403.815 2794.625 ;
        RECT 403.230 2794.610 403.815 2794.620 ;
        RECT 396.790 2794.310 397.835 2794.610 ;
        RECT 403.030 2794.310 403.815 2794.610 ;
        RECT 396.790 2794.300 397.170 2794.310 ;
        RECT 386.925 2794.295 387.255 2794.300 ;
        RECT 392.445 2794.295 392.775 2794.300 ;
        RECT 397.505 2794.295 397.835 2794.310 ;
        RECT 403.230 2794.300 403.815 2794.310 ;
        RECT 403.485 2794.295 403.815 2794.300 ;
        RECT 407.165 2794.610 407.495 2794.625 ;
        RECT 414.525 2794.620 414.855 2794.625 ;
        RECT 410.590 2794.610 410.970 2794.620 ;
        RECT 414.270 2794.610 414.855 2794.620 ;
        RECT 407.165 2794.310 410.970 2794.610 ;
        RECT 414.070 2794.310 414.855 2794.610 ;
        RECT 407.165 2794.295 407.495 2794.310 ;
        RECT 410.590 2794.300 410.970 2794.310 ;
        RECT 414.270 2794.300 414.855 2794.310 ;
        RECT 414.525 2794.295 414.855 2794.300 ;
        RECT 420.965 2794.610 421.295 2794.625 ;
        RECT 426.945 2794.620 427.275 2794.625 ;
        RECT 428.325 2794.620 428.655 2794.625 ;
        RECT 423.470 2794.610 423.850 2794.620 ;
        RECT 420.965 2794.310 423.850 2794.610 ;
        RECT 420.965 2794.295 421.295 2794.310 ;
        RECT 423.470 2794.300 423.850 2794.310 ;
        RECT 426.945 2794.610 427.530 2794.620 ;
        RECT 428.070 2794.610 428.655 2794.620 ;
        RECT 431.085 2794.610 431.415 2794.625 ;
        RECT 433.590 2794.610 433.970 2794.620 ;
        RECT 426.945 2794.310 427.730 2794.610 ;
        RECT 428.070 2794.310 428.880 2794.610 ;
        RECT 431.085 2794.310 433.970 2794.610 ;
        RECT 426.945 2794.300 427.530 2794.310 ;
        RECT 428.070 2794.300 428.655 2794.310 ;
        RECT 426.945 2794.295 427.275 2794.300 ;
        RECT 428.325 2794.295 428.655 2794.300 ;
        RECT 431.085 2794.295 431.415 2794.310 ;
        RECT 433.590 2794.300 433.970 2794.310 ;
        RECT 437.985 2794.610 438.315 2794.625 ;
        RECT 444.885 2794.620 445.215 2794.625 ;
        RECT 440.950 2794.610 441.330 2794.620 ;
        RECT 444.630 2794.610 445.215 2794.620 ;
        RECT 437.985 2794.310 441.330 2794.610 ;
        RECT 444.430 2794.310 445.215 2794.610 ;
        RECT 437.985 2794.295 438.315 2794.310 ;
        RECT 440.950 2794.300 441.330 2794.310 ;
        RECT 444.630 2794.300 445.215 2794.310 ;
        RECT 445.550 2794.610 445.930 2794.620 ;
        RECT 448.105 2794.610 448.435 2794.625 ;
        RECT 450.405 2794.620 450.735 2794.625 ;
        RECT 456.845 2794.620 457.175 2794.625 ;
        RECT 462.365 2794.620 462.695 2794.625 ;
        RECT 467.885 2794.620 468.215 2794.625 ;
        RECT 450.150 2794.610 450.735 2794.620 ;
        RECT 456.590 2794.610 457.175 2794.620 ;
        RECT 462.110 2794.610 462.695 2794.620 ;
        RECT 467.630 2794.610 468.215 2794.620 ;
        RECT 445.550 2794.310 448.435 2794.610 ;
        RECT 449.950 2794.310 450.735 2794.610 ;
        RECT 456.390 2794.310 457.175 2794.610 ;
        RECT 461.910 2794.310 462.695 2794.610 ;
        RECT 467.430 2794.310 468.215 2794.610 ;
        RECT 445.550 2794.300 445.930 2794.310 ;
        RECT 444.885 2794.295 445.215 2794.300 ;
        RECT 448.105 2794.295 448.435 2794.310 ;
        RECT 450.150 2794.300 450.735 2794.310 ;
        RECT 456.590 2794.300 457.175 2794.310 ;
        RECT 462.110 2794.300 462.695 2794.310 ;
        RECT 467.630 2794.300 468.215 2794.310 ;
        RECT 450.405 2794.295 450.735 2794.300 ;
        RECT 456.845 2794.295 457.175 2794.300 ;
        RECT 462.365 2794.295 462.695 2794.300 ;
        RECT 467.885 2794.295 468.215 2794.300 ;
        RECT 472.945 2794.620 473.275 2794.625 ;
        RECT 476.625 2794.620 476.955 2794.625 ;
        RECT 483.065 2794.620 483.395 2794.625 ;
        RECT 491.345 2794.620 491.675 2794.625 ;
        RECT 497.785 2794.620 498.115 2794.625 ;
        RECT 472.945 2794.610 473.530 2794.620 ;
        RECT 476.625 2794.610 477.210 2794.620 ;
        RECT 483.065 2794.610 483.650 2794.620 ;
        RECT 491.345 2794.610 491.930 2794.620 ;
        RECT 497.785 2794.610 498.370 2794.620 ;
        RECT 500.750 2794.610 501.130 2794.620 ;
        RECT 503.305 2794.610 503.635 2794.625 ;
        RECT 509.745 2794.620 510.075 2794.625 ;
        RECT 513.425 2794.620 513.755 2794.625 ;
        RECT 509.745 2794.610 510.330 2794.620 ;
        RECT 472.945 2794.310 473.730 2794.610 ;
        RECT 476.625 2794.310 477.410 2794.610 ;
        RECT 483.065 2794.310 483.850 2794.610 ;
        RECT 491.345 2794.310 492.130 2794.610 ;
        RECT 497.785 2794.310 498.570 2794.610 ;
        RECT 500.750 2794.310 503.635 2794.610 ;
        RECT 509.520 2794.310 510.330 2794.610 ;
        RECT 472.945 2794.300 473.530 2794.310 ;
        RECT 476.625 2794.300 477.210 2794.310 ;
        RECT 483.065 2794.300 483.650 2794.310 ;
        RECT 491.345 2794.300 491.930 2794.310 ;
        RECT 497.785 2794.300 498.370 2794.310 ;
        RECT 500.750 2794.300 501.130 2794.310 ;
        RECT 472.945 2794.295 473.275 2794.300 ;
        RECT 476.625 2794.295 476.955 2794.300 ;
        RECT 483.065 2794.295 483.395 2794.300 ;
        RECT 491.345 2794.295 491.675 2794.300 ;
        RECT 497.785 2794.295 498.115 2794.300 ;
        RECT 503.305 2794.295 503.635 2794.310 ;
        RECT 509.745 2794.300 510.330 2794.310 ;
        RECT 513.425 2794.610 514.010 2794.620 ;
        RECT 516.390 2794.610 516.770 2794.620 ;
        RECT 517.105 2794.610 517.435 2794.625 ;
        RECT 513.425 2794.310 514.210 2794.610 ;
        RECT 516.390 2794.310 517.435 2794.610 ;
        RECT 513.425 2794.300 514.010 2794.310 ;
        RECT 516.390 2794.300 516.770 2794.310 ;
        RECT 509.745 2794.295 510.075 2794.300 ;
        RECT 513.425 2794.295 513.755 2794.300 ;
        RECT 517.105 2794.295 517.435 2794.310 ;
        RECT 519.865 2794.620 520.195 2794.625 ;
        RECT 524.005 2794.620 524.335 2794.625 ;
        RECT 526.765 2794.620 527.095 2794.625 ;
        RECT 519.865 2794.610 520.450 2794.620 ;
        RECT 523.750 2794.610 524.335 2794.620 ;
        RECT 526.510 2794.610 527.095 2794.620 ;
        RECT 519.865 2794.310 520.650 2794.610 ;
        RECT 523.750 2794.310 524.560 2794.610 ;
        RECT 526.310 2794.310 527.095 2794.610 ;
        RECT 519.865 2794.300 520.450 2794.310 ;
        RECT 523.750 2794.300 524.335 2794.310 ;
        RECT 526.510 2794.300 527.095 2794.310 ;
        RECT 530.190 2794.610 530.570 2794.620 ;
        RECT 530.905 2794.610 531.235 2794.625 ;
        RECT 530.190 2794.310 531.235 2794.610 ;
        RECT 530.190 2794.300 530.570 2794.310 ;
        RECT 519.865 2794.295 520.195 2794.300 ;
        RECT 524.005 2794.295 524.335 2794.300 ;
        RECT 526.765 2794.295 527.095 2794.300 ;
        RECT 530.905 2794.295 531.235 2794.310 ;
        RECT 535.710 2794.610 536.090 2794.620 ;
        RECT 537.805 2794.610 538.135 2794.625 ;
        RECT 535.710 2794.310 538.135 2794.610 ;
        RECT 535.710 2794.300 536.090 2794.310 ;
        RECT 537.805 2794.295 538.135 2794.310 ;
        RECT 538.470 2794.610 538.850 2794.620 ;
        RECT 539.185 2794.610 539.515 2794.625 ;
        RECT 538.470 2794.310 539.515 2794.610 ;
        RECT 538.470 2794.300 538.850 2794.310 ;
        RECT 539.185 2794.295 539.515 2794.310 ;
        RECT 542.150 2794.610 542.530 2794.620 ;
        RECT 544.705 2794.610 545.035 2794.625 ;
        RECT 542.150 2794.310 545.035 2794.610 ;
        RECT 542.150 2794.300 542.530 2794.310 ;
        RECT 544.705 2794.295 545.035 2794.310 ;
        RECT 547.670 2794.610 548.050 2794.620 ;
        RECT 551.605 2794.610 551.935 2794.625 ;
        RECT 547.670 2794.310 551.935 2794.610 ;
        RECT 547.670 2794.300 548.050 2794.310 ;
        RECT 551.605 2794.295 551.935 2794.310 ;
        RECT 1013.190 2794.610 1013.570 2794.620 ;
        RECT 1013.905 2794.610 1014.235 2794.625 ;
        RECT 1013.190 2794.310 1014.235 2794.610 ;
        RECT 1013.190 2794.300 1013.570 2794.310 ;
        RECT 1013.905 2794.295 1014.235 2794.310 ;
        RECT 1019.630 2794.610 1020.010 2794.620 ;
        RECT 1020.805 2794.610 1021.135 2794.625 ;
        RECT 1019.630 2794.310 1021.135 2794.610 ;
        RECT 1019.630 2794.300 1020.010 2794.310 ;
        RECT 1020.805 2794.295 1021.135 2794.310 ;
        RECT 1026.990 2794.610 1027.370 2794.620 ;
        RECT 1027.705 2794.610 1028.035 2794.625 ;
        RECT 1059.445 2794.620 1059.775 2794.625 ;
        RECT 1065.885 2794.620 1066.215 2794.625 ;
        RECT 1059.190 2794.610 1059.775 2794.620 ;
        RECT 1065.630 2794.610 1066.215 2794.620 ;
        RECT 1026.990 2794.310 1028.035 2794.610 ;
        RECT 1058.990 2794.310 1059.775 2794.610 ;
        RECT 1065.430 2794.310 1066.215 2794.610 ;
        RECT 1026.990 2794.300 1027.370 2794.310 ;
        RECT 1027.705 2794.295 1028.035 2794.310 ;
        RECT 1059.190 2794.300 1059.775 2794.310 ;
        RECT 1065.630 2794.300 1066.215 2794.310 ;
        RECT 1059.445 2794.295 1059.775 2794.300 ;
        RECT 1065.885 2794.295 1066.215 2794.300 ;
        RECT 1069.565 2794.610 1069.895 2794.625 ;
        RECT 1070.230 2794.610 1070.610 2794.620 ;
        RECT 1069.565 2794.310 1070.610 2794.610 ;
        RECT 1069.565 2794.295 1069.895 2794.310 ;
        RECT 1070.230 2794.300 1070.610 2794.310 ;
        RECT 1081.270 2794.610 1081.650 2794.620 ;
        RECT 1082.905 2794.610 1083.235 2794.625 ;
        RECT 1087.965 2794.620 1088.295 2794.625 ;
        RECT 1087.710 2794.610 1088.295 2794.620 ;
        RECT 1089.345 2794.620 1089.675 2794.625 ;
        RECT 1094.405 2794.620 1094.735 2794.625 ;
        RECT 1089.345 2794.610 1089.930 2794.620 ;
        RECT 1094.150 2794.610 1094.735 2794.620 ;
        RECT 1081.270 2794.310 1083.235 2794.610 ;
        RECT 1087.510 2794.310 1088.295 2794.610 ;
        RECT 1089.120 2794.310 1089.930 2794.610 ;
        RECT 1093.950 2794.310 1094.735 2794.610 ;
        RECT 1081.270 2794.300 1081.650 2794.310 ;
        RECT 1082.905 2794.295 1083.235 2794.310 ;
        RECT 1087.710 2794.300 1088.295 2794.310 ;
        RECT 1087.965 2794.295 1088.295 2794.300 ;
        RECT 1089.345 2794.300 1089.930 2794.310 ;
        RECT 1094.150 2794.300 1094.735 2794.310 ;
        RECT 1095.990 2794.610 1096.370 2794.620 ;
        RECT 1096.705 2794.610 1097.035 2794.625 ;
        RECT 1095.990 2794.310 1097.035 2794.610 ;
        RECT 1095.990 2794.300 1096.370 2794.310 ;
        RECT 1089.345 2794.295 1089.675 2794.300 ;
        RECT 1094.405 2794.295 1094.735 2794.300 ;
        RECT 1096.705 2794.295 1097.035 2794.310 ;
        RECT 1100.385 2794.620 1100.715 2794.625 ;
        RECT 1103.605 2794.620 1103.935 2794.625 ;
        RECT 1105.445 2794.620 1105.775 2794.625 ;
        RECT 1100.385 2794.610 1100.970 2794.620 ;
        RECT 1103.350 2794.610 1103.935 2794.620 ;
        RECT 1105.190 2794.610 1105.775 2794.620 ;
        RECT 1100.385 2794.310 1101.170 2794.610 ;
        RECT 1103.350 2794.310 1104.160 2794.610 ;
        RECT 1104.990 2794.310 1105.775 2794.610 ;
        RECT 1100.385 2794.300 1100.970 2794.310 ;
        RECT 1103.350 2794.300 1103.935 2794.310 ;
        RECT 1105.190 2794.300 1105.775 2794.310 ;
        RECT 1109.790 2794.610 1110.170 2794.620 ;
        RECT 1110.505 2794.610 1110.835 2794.625 ;
        RECT 1109.790 2794.310 1110.835 2794.610 ;
        RECT 1109.790 2794.300 1110.170 2794.310 ;
        RECT 1100.385 2794.295 1100.715 2794.300 ;
        RECT 1103.605 2794.295 1103.935 2794.300 ;
        RECT 1105.445 2794.295 1105.775 2794.300 ;
        RECT 1110.505 2794.295 1110.835 2794.310 ;
        RECT 1111.425 2794.620 1111.755 2794.625 ;
        RECT 1111.425 2794.610 1112.010 2794.620 ;
        RECT 1116.230 2794.610 1116.610 2794.620 ;
        RECT 1117.405 2794.610 1117.735 2794.625 ;
        RECT 1111.425 2794.310 1112.210 2794.610 ;
        RECT 1116.230 2794.310 1117.735 2794.610 ;
        RECT 1111.425 2794.300 1112.010 2794.310 ;
        RECT 1116.230 2794.300 1116.610 2794.310 ;
        RECT 1111.425 2794.295 1111.755 2794.300 ;
        RECT 1117.405 2794.295 1117.735 2794.310 ;
        RECT 1121.750 2794.610 1122.130 2794.620 ;
        RECT 1124.305 2794.610 1124.635 2794.625 ;
        RECT 1121.750 2794.310 1124.635 2794.610 ;
        RECT 1121.750 2794.300 1122.130 2794.310 ;
        RECT 1124.305 2794.295 1124.635 2794.310 ;
        RECT 1128.905 2794.620 1129.235 2794.625 ;
        RECT 1131.205 2794.620 1131.535 2794.625 ;
        RECT 1135.805 2794.620 1136.135 2794.625 ;
        RECT 1128.905 2794.610 1129.490 2794.620 ;
        RECT 1130.950 2794.610 1131.535 2794.620 ;
        RECT 1135.550 2794.610 1136.135 2794.620 ;
        RECT 1128.905 2794.310 1129.690 2794.610 ;
        RECT 1130.950 2794.310 1131.760 2794.610 ;
        RECT 1135.350 2794.310 1136.135 2794.610 ;
        RECT 1128.905 2794.300 1129.490 2794.310 ;
        RECT 1130.950 2794.300 1131.535 2794.310 ;
        RECT 1135.550 2794.300 1136.135 2794.310 ;
        RECT 1137.390 2794.610 1137.770 2794.620 ;
        RECT 1138.105 2794.610 1138.435 2794.625 ;
        RECT 1137.390 2794.310 1138.435 2794.610 ;
        RECT 1137.390 2794.300 1137.770 2794.310 ;
        RECT 1128.905 2794.295 1129.235 2794.300 ;
        RECT 1131.205 2794.295 1131.535 2794.300 ;
        RECT 1135.805 2794.295 1136.135 2794.300 ;
        RECT 1138.105 2794.295 1138.435 2794.310 ;
        RECT 1143.830 2794.610 1144.210 2794.620 ;
        RECT 1145.005 2794.610 1145.335 2794.625 ;
        RECT 1143.830 2794.310 1145.335 2794.610 ;
        RECT 1143.830 2794.300 1144.210 2794.310 ;
        RECT 1145.005 2794.295 1145.335 2794.310 ;
        RECT 1147.305 2794.620 1147.635 2794.625 ;
        RECT 1147.305 2794.610 1147.890 2794.620 ;
        RECT 1151.190 2794.610 1151.570 2794.620 ;
        RECT 1151.905 2794.610 1152.235 2794.625 ;
        RECT 1147.305 2794.310 1148.090 2794.610 ;
        RECT 1151.190 2794.310 1152.235 2794.610 ;
        RECT 1147.305 2794.300 1147.890 2794.310 ;
        RECT 1151.190 2794.300 1151.570 2794.310 ;
        RECT 1147.305 2794.295 1147.635 2794.300 ;
        RECT 1151.905 2794.295 1152.235 2794.310 ;
        RECT 1153.950 2794.610 1154.330 2794.620 ;
        RECT 1158.805 2794.610 1159.135 2794.625 ;
        RECT 1153.950 2794.310 1159.135 2794.610 ;
        RECT 1153.950 2794.300 1154.330 2794.310 ;
        RECT 1158.805 2794.295 1159.135 2794.310 ;
        RECT 1159.725 2794.610 1160.055 2794.625 ;
        RECT 1164.070 2794.610 1164.450 2794.620 ;
        RECT 1159.725 2794.310 1164.450 2794.610 ;
        RECT 1159.725 2794.295 1160.055 2794.310 ;
        RECT 1164.070 2794.300 1164.450 2794.310 ;
        RECT 1164.990 2794.610 1165.370 2794.620 ;
        RECT 1165.705 2794.610 1166.035 2794.625 ;
        RECT 1172.605 2794.620 1172.935 2794.625 ;
        RECT 1164.990 2794.310 1166.035 2794.610 ;
        RECT 1164.990 2794.300 1165.370 2794.310 ;
        RECT 1165.705 2794.295 1166.035 2794.310 ;
        RECT 1172.350 2794.610 1172.935 2794.620 ;
        RECT 1178.790 2794.610 1179.170 2794.620 ;
        RECT 1179.505 2794.610 1179.835 2794.625 ;
        RECT 1186.405 2794.620 1186.735 2794.625 ;
        RECT 1172.350 2794.310 1173.160 2794.610 ;
        RECT 1178.790 2794.310 1179.835 2794.610 ;
        RECT 1172.350 2794.300 1172.935 2794.310 ;
        RECT 1178.790 2794.300 1179.170 2794.310 ;
        RECT 1172.605 2794.295 1172.935 2794.300 ;
        RECT 1179.505 2794.295 1179.835 2794.310 ;
        RECT 1186.150 2794.610 1186.735 2794.620 ;
        RECT 1198.110 2794.610 1198.490 2794.620 ;
        RECT 1200.205 2794.610 1200.535 2794.625 ;
        RECT 1186.150 2794.310 1186.960 2794.610 ;
        RECT 1198.110 2794.310 1200.535 2794.610 ;
        RECT 1186.150 2794.300 1186.735 2794.310 ;
        RECT 1198.110 2794.300 1198.490 2794.310 ;
        RECT 1186.405 2794.295 1186.735 2794.300 ;
        RECT 1200.205 2794.295 1200.535 2794.310 ;
        RECT 1580.165 2794.610 1580.495 2794.625 ;
        RECT 1580.830 2794.610 1581.210 2794.620 ;
        RECT 1580.165 2794.310 1581.210 2794.610 ;
        RECT 1580.165 2794.295 1580.495 2794.310 ;
        RECT 1580.830 2794.300 1581.210 2794.310 ;
        RECT 1593.965 2794.610 1594.295 2794.625 ;
        RECT 1594.630 2794.610 1595.010 2794.620 ;
        RECT 1593.965 2794.310 1595.010 2794.610 ;
        RECT 1593.965 2794.295 1594.295 2794.310 ;
        RECT 1594.630 2794.300 1595.010 2794.310 ;
        RECT 1601.325 2794.610 1601.655 2794.625 ;
        RECT 1604.750 2794.610 1605.130 2794.620 ;
        RECT 1601.325 2794.310 1605.130 2794.610 ;
        RECT 1601.325 2794.295 1601.655 2794.310 ;
        RECT 1604.750 2794.300 1605.130 2794.310 ;
        RECT 1607.765 2794.610 1608.095 2794.625 ;
        RECT 1613.950 2794.610 1614.330 2794.620 ;
        RECT 1607.765 2794.310 1614.330 2794.610 ;
        RECT 1607.765 2794.295 1608.095 2794.310 ;
        RECT 1613.950 2794.300 1614.330 2794.310 ;
        RECT 1617.885 2794.610 1618.215 2794.625 ;
        RECT 1625.910 2794.610 1626.290 2794.620 ;
        RECT 1617.885 2794.310 1626.290 2794.610 ;
        RECT 1617.885 2794.295 1618.215 2794.310 ;
        RECT 1625.910 2794.300 1626.290 2794.310 ;
        RECT 1628.465 2794.610 1628.795 2794.625 ;
        RECT 1631.430 2794.610 1631.810 2794.620 ;
        RECT 1628.465 2794.310 1631.810 2794.610 ;
        RECT 1628.465 2794.295 1628.795 2794.310 ;
        RECT 1631.430 2794.300 1631.810 2794.310 ;
        RECT 1635.365 2794.610 1635.695 2794.625 ;
        RECT 1637.870 2794.610 1638.250 2794.620 ;
        RECT 1635.365 2794.310 1638.250 2794.610 ;
        RECT 1635.365 2794.295 1635.695 2794.310 ;
        RECT 1637.870 2794.300 1638.250 2794.310 ;
        RECT 1649.625 2794.610 1649.955 2794.625 ;
        RECT 1658.825 2794.620 1659.155 2794.625 ;
        RECT 1655.350 2794.610 1655.730 2794.620 ;
        RECT 1649.625 2794.310 1655.730 2794.610 ;
        RECT 1649.625 2794.295 1649.955 2794.310 ;
        RECT 1655.350 2794.300 1655.730 2794.310 ;
        RECT 1658.825 2794.610 1659.410 2794.620 ;
        RECT 1662.965 2794.610 1663.295 2794.625 ;
        RECT 1666.390 2794.610 1666.770 2794.620 ;
        RECT 1658.825 2794.310 1659.610 2794.610 ;
        RECT 1662.965 2794.310 1666.770 2794.610 ;
        RECT 1658.825 2794.300 1659.410 2794.310 ;
        RECT 1658.825 2794.295 1659.155 2794.300 ;
        RECT 1662.965 2794.295 1663.295 2794.310 ;
        RECT 1666.390 2794.300 1666.770 2794.310 ;
        RECT 1669.865 2794.610 1670.195 2794.625 ;
        RECT 1672.830 2794.610 1673.210 2794.620 ;
        RECT 1669.865 2794.310 1673.210 2794.610 ;
        RECT 1669.865 2794.295 1670.195 2794.310 ;
        RECT 1672.830 2794.300 1673.210 2794.310 ;
        RECT 1676.765 2794.610 1677.095 2794.625 ;
        RECT 1683.665 2794.620 1683.995 2794.625 ;
        RECT 1679.270 2794.610 1679.650 2794.620 ;
        RECT 1683.665 2794.610 1684.250 2794.620 ;
        RECT 1676.765 2794.310 1679.650 2794.610 ;
        RECT 1683.440 2794.310 1684.250 2794.610 ;
        RECT 1676.765 2794.295 1677.095 2794.310 ;
        RECT 1679.270 2794.300 1679.650 2794.310 ;
        RECT 1683.665 2794.300 1684.250 2794.310 ;
        RECT 1686.885 2794.610 1687.215 2794.625 ;
        RECT 1688.470 2794.610 1688.850 2794.620 ;
        RECT 1686.885 2794.310 1688.850 2794.610 ;
        RECT 1683.665 2794.295 1683.995 2794.300 ;
        RECT 1686.885 2794.295 1687.215 2794.310 ;
        RECT 1688.470 2794.300 1688.850 2794.310 ;
        RECT 1690.565 2794.610 1690.895 2794.625 ;
        RECT 1695.830 2794.610 1696.210 2794.620 ;
        RECT 1690.565 2794.310 1696.210 2794.610 ;
        RECT 1690.565 2794.295 1690.895 2794.310 ;
        RECT 1695.830 2794.300 1696.210 2794.310 ;
        RECT 1697.465 2794.610 1697.795 2794.625 ;
        RECT 1702.270 2794.610 1702.650 2794.620 ;
        RECT 1697.465 2794.310 1702.650 2794.610 ;
        RECT 1697.465 2794.295 1697.795 2794.310 ;
        RECT 1702.270 2794.300 1702.650 2794.310 ;
        RECT 1704.365 2794.610 1704.695 2794.625 ;
        RECT 1708.710 2794.610 1709.090 2794.620 ;
        RECT 1704.365 2794.310 1709.090 2794.610 ;
        RECT 1704.365 2794.295 1704.695 2794.310 ;
        RECT 1708.710 2794.300 1709.090 2794.310 ;
        RECT 1711.265 2794.610 1711.595 2794.625 ;
        RECT 1713.310 2794.610 1713.690 2794.620 ;
        RECT 1711.265 2794.310 1713.690 2794.610 ;
        RECT 1711.265 2794.295 1711.595 2794.310 ;
        RECT 1713.310 2794.300 1713.690 2794.310 ;
        RECT 1718.165 2794.610 1718.495 2794.625 ;
        RECT 1721.385 2794.620 1721.715 2794.625 ;
        RECT 1719.750 2794.610 1720.130 2794.620 ;
        RECT 1718.165 2794.310 1720.130 2794.610 ;
        RECT 1718.165 2794.295 1718.495 2794.310 ;
        RECT 1719.750 2794.300 1720.130 2794.310 ;
        RECT 1721.385 2794.610 1721.970 2794.620 ;
        RECT 1725.065 2794.610 1725.395 2794.625 ;
        RECT 1730.790 2794.610 1731.170 2794.620 ;
        RECT 1721.385 2794.310 1722.170 2794.610 ;
        RECT 1725.065 2794.310 1731.170 2794.610 ;
        RECT 1721.385 2794.300 1721.970 2794.310 ;
        RECT 1721.385 2794.295 1721.715 2794.300 ;
        RECT 1725.065 2794.295 1725.395 2794.310 ;
        RECT 1730.790 2794.300 1731.170 2794.310 ;
        RECT 1731.965 2794.610 1732.295 2794.625 ;
        RECT 1737.230 2794.610 1737.610 2794.620 ;
        RECT 1731.965 2794.310 1737.610 2794.610 ;
        RECT 1731.965 2794.295 1732.295 2794.310 ;
        RECT 1737.230 2794.300 1737.610 2794.310 ;
        RECT 1738.865 2794.610 1739.195 2794.625 ;
        RECT 1743.670 2794.610 1744.050 2794.620 ;
        RECT 1738.865 2794.310 1744.050 2794.610 ;
        RECT 1738.865 2794.295 1739.195 2794.310 ;
        RECT 1743.670 2794.300 1744.050 2794.310 ;
        RECT 1745.765 2794.610 1746.095 2794.625 ;
        RECT 1748.270 2794.610 1748.650 2794.620 ;
        RECT 1745.765 2794.310 1748.650 2794.610 ;
        RECT 1745.765 2794.295 1746.095 2794.310 ;
        RECT 1748.270 2794.300 1748.650 2794.310 ;
        RECT 1759.565 2794.610 1759.895 2794.625 ;
        RECT 1762.070 2794.610 1762.450 2794.620 ;
        RECT 1759.565 2794.310 1762.450 2794.610 ;
        RECT 1759.565 2794.295 1759.895 2794.310 ;
        RECT 1762.070 2794.300 1762.450 2794.310 ;
        RECT 2228.765 2794.610 2229.095 2794.625 ;
        RECT 2231.270 2794.610 2231.650 2794.620 ;
        RECT 2228.765 2794.310 2231.650 2794.610 ;
        RECT 2228.765 2794.295 2229.095 2794.310 ;
        RECT 2231.270 2794.300 2231.650 2794.310 ;
        RECT 2231.985 2794.610 2232.315 2794.625 ;
        RECT 2236.790 2794.610 2237.170 2794.620 ;
        RECT 2231.985 2794.310 2237.170 2794.610 ;
        RECT 2231.985 2794.295 2232.315 2794.310 ;
        RECT 2236.790 2794.300 2237.170 2794.310 ;
        RECT 2238.885 2794.610 2239.215 2794.625 ;
        RECT 2242.310 2794.610 2242.690 2794.620 ;
        RECT 2238.885 2794.310 2242.690 2794.610 ;
        RECT 2238.885 2794.295 2239.215 2794.310 ;
        RECT 2242.310 2794.300 2242.690 2794.310 ;
        RECT 2245.785 2794.610 2246.115 2794.625 ;
        RECT 2249.670 2794.610 2250.050 2794.620 ;
        RECT 2245.785 2794.310 2250.050 2794.610 ;
        RECT 2245.785 2794.295 2246.115 2794.310 ;
        RECT 2249.670 2794.300 2250.050 2794.310 ;
        RECT 2263.725 2794.610 2264.055 2794.625 ;
        RECT 2264.390 2794.610 2264.770 2794.620 ;
        RECT 2263.725 2794.310 2264.770 2794.610 ;
        RECT 2263.725 2794.295 2264.055 2794.310 ;
        RECT 2264.390 2794.300 2264.770 2794.310 ;
        RECT 2267.405 2794.610 2267.735 2794.625 ;
        RECT 2273.385 2794.620 2273.715 2794.625 ;
        RECT 2268.070 2794.610 2268.450 2794.620 ;
        RECT 2267.405 2794.310 2268.450 2794.610 ;
        RECT 2267.405 2794.295 2267.735 2794.310 ;
        RECT 2268.070 2794.300 2268.450 2794.310 ;
        RECT 2273.385 2794.610 2273.970 2794.620 ;
        RECT 2291.990 2794.610 2292.370 2794.620 ;
        RECT 2294.085 2794.610 2294.415 2794.625 ;
        RECT 2273.385 2794.310 2274.170 2794.610 ;
        RECT 2291.990 2794.310 2294.415 2794.610 ;
        RECT 2273.385 2794.300 2273.970 2794.310 ;
        RECT 2291.990 2794.300 2292.370 2794.310 ;
        RECT 2273.385 2794.295 2273.715 2794.300 ;
        RECT 2294.085 2794.295 2294.415 2794.310 ;
        RECT 2304.665 2794.620 2304.995 2794.625 ;
        RECT 2308.805 2794.620 2309.135 2794.625 ;
        RECT 2304.665 2794.610 2305.250 2794.620 ;
        RECT 2308.550 2794.610 2309.135 2794.620 ;
        RECT 2304.665 2794.310 2305.450 2794.610 ;
        RECT 2308.350 2794.310 2309.135 2794.610 ;
        RECT 2304.665 2794.300 2305.250 2794.310 ;
        RECT 2308.550 2794.300 2309.135 2794.310 ;
        RECT 2304.665 2794.295 2304.995 2794.300 ;
        RECT 2308.805 2794.295 2309.135 2794.300 ;
        RECT 2311.565 2794.610 2311.895 2794.625 ;
        RECT 2316.830 2794.610 2317.210 2794.620 ;
        RECT 2311.565 2794.310 2317.210 2794.610 ;
        RECT 2311.565 2794.295 2311.895 2794.310 ;
        RECT 2316.830 2794.300 2317.210 2794.310 ;
        RECT 2318.465 2794.610 2318.795 2794.625 ;
        RECT 2322.350 2794.610 2322.730 2794.620 ;
        RECT 2318.465 2794.310 2322.730 2794.610 ;
        RECT 2318.465 2794.295 2318.795 2794.310 ;
        RECT 2322.350 2794.300 2322.730 2794.310 ;
        RECT 2325.365 2794.610 2325.695 2794.625 ;
        RECT 2328.790 2794.610 2329.170 2794.620 ;
        RECT 2325.365 2794.310 2329.170 2794.610 ;
        RECT 2325.365 2794.295 2325.695 2794.310 ;
        RECT 2328.790 2794.300 2329.170 2794.310 ;
        RECT 2332.265 2794.610 2332.595 2794.625 ;
        RECT 2334.310 2794.610 2334.690 2794.620 ;
        RECT 2332.265 2794.310 2334.690 2794.610 ;
        RECT 2332.265 2794.295 2332.595 2794.310 ;
        RECT 2334.310 2794.300 2334.690 2794.310 ;
        RECT 2339.165 2794.610 2339.495 2794.625 ;
        RECT 2339.830 2794.610 2340.210 2794.620 ;
        RECT 2339.165 2794.310 2340.210 2794.610 ;
        RECT 2339.165 2794.295 2339.495 2794.310 ;
        RECT 2339.830 2794.300 2340.210 2794.310 ;
        RECT 2342.845 2794.610 2343.175 2794.625 ;
        RECT 2343.510 2794.610 2343.890 2794.620 ;
        RECT 2342.845 2794.310 2343.890 2794.610 ;
        RECT 2342.845 2794.295 2343.175 2794.310 ;
        RECT 2343.510 2794.300 2343.890 2794.310 ;
        RECT 2346.065 2794.610 2346.395 2794.625 ;
        RECT 2351.790 2794.610 2352.170 2794.620 ;
        RECT 2346.065 2794.310 2352.170 2794.610 ;
        RECT 2346.065 2794.295 2346.395 2794.310 ;
        RECT 2351.790 2794.300 2352.170 2794.310 ;
        RECT 2352.965 2794.610 2353.295 2794.625 ;
        RECT 2357.310 2794.610 2357.690 2794.620 ;
        RECT 2352.965 2794.310 2357.690 2794.610 ;
        RECT 2352.965 2794.295 2353.295 2794.310 ;
        RECT 2357.310 2794.300 2357.690 2794.310 ;
        RECT 2359.865 2794.610 2360.195 2794.625 ;
        RECT 2363.750 2794.610 2364.130 2794.620 ;
        RECT 2359.865 2794.310 2364.130 2794.610 ;
        RECT 2359.865 2794.295 2360.195 2794.310 ;
        RECT 2363.750 2794.300 2364.130 2794.310 ;
        RECT 2366.765 2794.610 2367.095 2794.625 ;
        RECT 2370.190 2794.610 2370.570 2794.620 ;
        RECT 2366.765 2794.310 2370.570 2794.610 ;
        RECT 2366.765 2794.295 2367.095 2794.310 ;
        RECT 2370.190 2794.300 2370.570 2794.310 ;
        RECT 2373.665 2794.610 2373.995 2794.625 ;
        RECT 2381.025 2794.620 2381.355 2794.625 ;
        RECT 2385.625 2794.620 2385.955 2794.625 ;
        RECT 2391.605 2794.620 2391.935 2794.625 ;
        RECT 2397.125 2794.620 2397.455 2794.625 ;
        RECT 2374.790 2794.610 2375.170 2794.620 ;
        RECT 2381.025 2794.610 2381.610 2794.620 ;
        RECT 2373.665 2794.310 2375.170 2794.610 ;
        RECT 2380.800 2794.310 2381.610 2794.610 ;
        RECT 2373.665 2794.295 2373.995 2794.310 ;
        RECT 2374.790 2794.300 2375.170 2794.310 ;
        RECT 2381.025 2794.300 2381.610 2794.310 ;
        RECT 2385.625 2794.610 2386.210 2794.620 ;
        RECT 2391.350 2794.610 2391.935 2794.620 ;
        RECT 2396.870 2794.610 2397.455 2794.620 ;
        RECT 2385.625 2794.310 2386.410 2794.610 ;
        RECT 2391.150 2794.310 2391.935 2794.610 ;
        RECT 2396.670 2794.310 2397.455 2794.610 ;
        RECT 2385.625 2794.300 2386.210 2794.310 ;
        RECT 2391.350 2794.300 2391.935 2794.310 ;
        RECT 2396.870 2794.300 2397.455 2794.310 ;
        RECT 2381.025 2794.295 2381.355 2794.300 ;
        RECT 2385.625 2794.295 2385.955 2794.300 ;
        RECT 2391.605 2794.295 2391.935 2794.300 ;
        RECT 2397.125 2794.295 2397.455 2794.300 ;
        RECT 2402.645 2794.610 2402.975 2794.625 ;
        RECT 2404.230 2794.610 2404.610 2794.620 ;
        RECT 2402.645 2794.310 2404.610 2794.610 ;
        RECT 2402.645 2794.295 2402.975 2794.310 ;
        RECT 2404.230 2794.300 2404.610 2794.310 ;
        RECT 2415.065 2794.610 2415.395 2794.625 ;
        RECT 2417.110 2794.610 2417.490 2794.620 ;
        RECT 2415.065 2794.310 2417.490 2794.610 ;
        RECT 2415.065 2794.295 2415.395 2794.310 ;
        RECT 2417.110 2794.300 2417.490 2794.310 ;
        RECT 2422.425 2794.610 2422.755 2794.625 ;
        RECT 2428.150 2794.610 2428.530 2794.620 ;
        RECT 2422.425 2794.310 2428.530 2794.610 ;
        RECT 2422.425 2794.295 2422.755 2794.310 ;
        RECT 2428.150 2794.300 2428.530 2794.310 ;
        RECT 2428.865 2794.610 2429.195 2794.625 ;
        RECT 2429.990 2794.610 2430.370 2794.620 ;
        RECT 2428.865 2794.310 2430.370 2794.610 ;
        RECT 2428.865 2794.295 2429.195 2794.310 ;
        RECT 2429.990 2794.300 2430.370 2794.310 ;
        RECT 351.045 2793.940 351.375 2793.945 ;
        RECT 350.790 2793.930 351.375 2793.940 ;
        RECT 400.265 2793.930 400.595 2793.945 ;
        RECT 405.070 2793.930 405.450 2793.940 ;
        RECT 350.790 2793.630 351.600 2793.930 ;
        RECT 400.265 2793.630 405.450 2793.930 ;
        RECT 350.790 2793.620 351.375 2793.630 ;
        RECT 351.045 2793.615 351.375 2793.620 ;
        RECT 400.265 2793.615 400.595 2793.630 ;
        RECT 405.070 2793.620 405.450 2793.630 ;
        RECT 408.085 2793.930 408.415 2793.945 ;
        RECT 408.750 2793.930 409.130 2793.940 ;
        RECT 408.085 2793.630 409.130 2793.930 ;
        RECT 408.085 2793.615 408.415 2793.630 ;
        RECT 408.750 2793.620 409.130 2793.630 ;
        RECT 420.710 2793.930 421.090 2793.940 ;
        RECT 421.425 2793.930 421.755 2793.945 ;
        RECT 420.710 2793.630 421.755 2793.930 ;
        RECT 420.710 2793.620 421.090 2793.630 ;
        RECT 421.425 2793.615 421.755 2793.630 ;
        RECT 431.750 2793.930 432.130 2793.940 ;
        RECT 434.305 2793.930 434.635 2793.945 ;
        RECT 439.365 2793.940 439.695 2793.945 ;
        RECT 439.110 2793.930 439.695 2793.940 ;
        RECT 431.750 2793.630 434.635 2793.930 ;
        RECT 438.910 2793.630 439.695 2793.930 ;
        RECT 431.750 2793.620 432.130 2793.630 ;
        RECT 434.305 2793.615 434.635 2793.630 ;
        RECT 439.110 2793.620 439.695 2793.630 ;
        RECT 439.365 2793.615 439.695 2793.620 ;
        RECT 501.465 2793.940 501.795 2793.945 ;
        RECT 501.465 2793.930 502.050 2793.940 ;
        RECT 507.190 2793.930 507.570 2793.940 ;
        RECT 510.205 2793.930 510.535 2793.945 ;
        RECT 531.365 2793.940 531.695 2793.945 ;
        RECT 531.110 2793.930 531.695 2793.940 ;
        RECT 501.465 2793.630 502.250 2793.930 ;
        RECT 507.190 2793.630 510.535 2793.930 ;
        RECT 530.910 2793.630 531.695 2793.930 ;
        RECT 501.465 2793.620 502.050 2793.630 ;
        RECT 507.190 2793.620 507.570 2793.630 ;
        RECT 501.465 2793.615 501.795 2793.620 ;
        RECT 510.205 2793.615 510.535 2793.630 ;
        RECT 531.110 2793.620 531.695 2793.630 ;
        RECT 531.365 2793.615 531.695 2793.620 ;
        RECT 542.865 2793.940 543.195 2793.945 ;
        RECT 542.865 2793.930 543.450 2793.940 ;
        RECT 979.865 2793.930 980.195 2793.945 ;
        RECT 980.990 2793.930 981.370 2793.940 ;
        RECT 542.865 2793.630 543.650 2793.930 ;
        RECT 979.865 2793.630 981.370 2793.930 ;
        RECT 542.865 2793.620 543.450 2793.630 ;
        RECT 542.865 2793.615 543.195 2793.620 ;
        RECT 979.865 2793.615 980.195 2793.630 ;
        RECT 980.990 2793.620 981.370 2793.630 ;
        RECT 1007.465 2793.930 1007.795 2793.945 ;
        RECT 1008.590 2793.930 1008.970 2793.940 ;
        RECT 1007.465 2793.630 1008.970 2793.930 ;
        RECT 1007.465 2793.615 1007.795 2793.630 ;
        RECT 1008.590 2793.620 1008.970 2793.630 ;
        RECT 1010.685 2793.930 1011.015 2793.945 ;
        RECT 1024.485 2793.940 1024.815 2793.945 ;
        RECT 1012.270 2793.930 1012.650 2793.940 ;
        RECT 1024.230 2793.930 1024.815 2793.940 ;
        RECT 1010.685 2793.630 1012.650 2793.930 ;
        RECT 1024.030 2793.630 1024.815 2793.930 ;
        RECT 1010.685 2793.615 1011.015 2793.630 ;
        RECT 1012.270 2793.620 1012.650 2793.630 ;
        RECT 1024.230 2793.620 1024.815 2793.630 ;
        RECT 1024.485 2793.615 1024.815 2793.620 ;
        RECT 1076.465 2793.940 1076.795 2793.945 ;
        RECT 1076.465 2793.930 1077.050 2793.940 ;
        RECT 1083.110 2793.930 1083.490 2793.940 ;
        RECT 1083.825 2793.930 1084.155 2793.945 ;
        RECT 1076.465 2793.630 1077.250 2793.930 ;
        RECT 1083.110 2793.630 1084.155 2793.930 ;
        RECT 1076.465 2793.620 1077.050 2793.630 ;
        RECT 1083.110 2793.620 1083.490 2793.630 ;
        RECT 1076.465 2793.615 1076.795 2793.620 ;
        RECT 1083.825 2793.615 1084.155 2793.630 ;
        RECT 1086.790 2793.930 1087.170 2793.940 ;
        RECT 1089.805 2793.930 1090.135 2793.945 ;
        RECT 1086.790 2793.630 1090.135 2793.930 ;
        RECT 1086.790 2793.620 1087.170 2793.630 ;
        RECT 1089.805 2793.615 1090.135 2793.630 ;
        RECT 1117.865 2793.940 1118.195 2793.945 ;
        RECT 1117.865 2793.930 1118.450 2793.940 ;
        RECT 1122.005 2793.930 1122.335 2793.945 ;
        RECT 1122.670 2793.930 1123.050 2793.940 ;
        RECT 1117.865 2793.630 1118.650 2793.930 ;
        RECT 1122.005 2793.630 1123.050 2793.930 ;
        RECT 1117.865 2793.620 1118.450 2793.630 ;
        RECT 1117.865 2793.615 1118.195 2793.620 ;
        RECT 1122.005 2793.615 1122.335 2793.630 ;
        RECT 1122.670 2793.620 1123.050 2793.630 ;
        RECT 1128.190 2793.930 1128.570 2793.940 ;
        RECT 1130.745 2793.930 1131.075 2793.945 ;
        RECT 1128.190 2793.630 1131.075 2793.930 ;
        RECT 1128.190 2793.620 1128.570 2793.630 ;
        RECT 1130.745 2793.615 1131.075 2793.630 ;
        RECT 1138.565 2793.930 1138.895 2793.945 ;
        RECT 1139.230 2793.930 1139.610 2793.940 ;
        RECT 1138.565 2793.630 1139.610 2793.930 ;
        RECT 1138.565 2793.615 1138.895 2793.630 ;
        RECT 1139.230 2793.620 1139.610 2793.630 ;
        RECT 1163.150 2793.930 1163.530 2793.940 ;
        RECT 1165.245 2793.930 1165.575 2793.945 ;
        RECT 1163.150 2793.630 1165.575 2793.930 ;
        RECT 1163.150 2793.620 1163.530 2793.630 ;
        RECT 1165.245 2793.615 1165.575 2793.630 ;
        RECT 1166.165 2793.930 1166.495 2793.945 ;
        RECT 1167.750 2793.930 1168.130 2793.940 ;
        RECT 1166.165 2793.630 1168.130 2793.930 ;
        RECT 1166.165 2793.615 1166.495 2793.630 ;
        RECT 1167.750 2793.620 1168.130 2793.630 ;
        RECT 1179.965 2793.930 1180.295 2793.945 ;
        RECT 1180.630 2793.930 1181.010 2793.940 ;
        RECT 1179.965 2793.630 1181.010 2793.930 ;
        RECT 1179.965 2793.615 1180.295 2793.630 ;
        RECT 1180.630 2793.620 1181.010 2793.630 ;
        RECT 1611.445 2793.930 1611.775 2793.945 ;
        RECT 1612.110 2793.930 1612.490 2793.940 ;
        RECT 1611.445 2793.630 1612.490 2793.930 ;
        RECT 1611.445 2793.615 1611.775 2793.630 ;
        RECT 1612.110 2793.620 1612.490 2793.630 ;
        RECT 1635.110 2793.930 1635.490 2793.940 ;
        RECT 1638.585 2793.930 1638.915 2793.945 ;
        RECT 1635.110 2793.630 1638.915 2793.930 ;
        RECT 1635.110 2793.620 1635.490 2793.630 ;
        RECT 1638.585 2793.615 1638.915 2793.630 ;
        RECT 1642.470 2793.930 1642.850 2793.940 ;
        RECT 1645.485 2793.930 1645.815 2793.945 ;
        RECT 1642.470 2793.630 1645.815 2793.930 ;
        RECT 1642.470 2793.620 1642.850 2793.630 ;
        RECT 1645.485 2793.615 1645.815 2793.630 ;
        RECT 1663.425 2793.940 1663.755 2793.945 ;
        RECT 1670.325 2793.940 1670.655 2793.945 ;
        RECT 1663.425 2793.930 1664.010 2793.940 ;
        RECT 1670.070 2793.930 1670.655 2793.940 ;
        RECT 1663.425 2793.630 1664.210 2793.930 ;
        RECT 1669.870 2793.630 1670.655 2793.930 ;
        RECT 1663.425 2793.620 1664.010 2793.630 ;
        RECT 1670.070 2793.620 1670.655 2793.630 ;
        RECT 1663.425 2793.615 1663.755 2793.620 ;
        RECT 1670.325 2793.615 1670.655 2793.620 ;
        RECT 1677.225 2793.940 1677.555 2793.945 ;
        RECT 1683.205 2793.940 1683.535 2793.945 ;
        RECT 1677.225 2793.930 1677.810 2793.940 ;
        RECT 1682.950 2793.930 1683.535 2793.940 ;
        RECT 1677.225 2793.630 1678.010 2793.930 ;
        RECT 1682.750 2793.630 1683.535 2793.930 ;
        RECT 1677.225 2793.620 1677.810 2793.630 ;
        RECT 1682.950 2793.620 1683.535 2793.630 ;
        RECT 1677.225 2793.615 1677.555 2793.620 ;
        RECT 1683.205 2793.615 1683.535 2793.620 ;
        RECT 1694.705 2793.940 1695.035 2793.945 ;
        RECT 1699.305 2793.940 1699.635 2793.945 ;
        RECT 1704.825 2793.940 1705.155 2793.945 ;
        RECT 1712.645 2793.940 1712.975 2793.945 ;
        RECT 1694.705 2793.930 1695.290 2793.940 ;
        RECT 1699.305 2793.930 1699.890 2793.940 ;
        RECT 1704.825 2793.930 1705.410 2793.940 ;
        RECT 1712.390 2793.930 1712.975 2793.940 ;
        RECT 1694.705 2793.630 1695.490 2793.930 ;
        RECT 1699.305 2793.630 1700.090 2793.930 ;
        RECT 1704.825 2793.630 1705.610 2793.930 ;
        RECT 1712.190 2793.630 1712.975 2793.930 ;
        RECT 1694.705 2793.620 1695.290 2793.630 ;
        RECT 1699.305 2793.620 1699.890 2793.630 ;
        RECT 1704.825 2793.620 1705.410 2793.630 ;
        RECT 1712.390 2793.620 1712.975 2793.630 ;
        RECT 1717.910 2793.930 1718.290 2793.940 ;
        RECT 1718.625 2793.930 1718.955 2793.945 ;
        RECT 1717.910 2793.630 1718.955 2793.930 ;
        RECT 1717.910 2793.620 1718.290 2793.630 ;
        RECT 1694.705 2793.615 1695.035 2793.620 ;
        RECT 1699.305 2793.615 1699.635 2793.620 ;
        RECT 1704.825 2793.615 1705.155 2793.620 ;
        RECT 1712.645 2793.615 1712.975 2793.620 ;
        RECT 1718.625 2793.615 1718.955 2793.630 ;
        RECT 1729.870 2793.930 1730.250 2793.940 ;
        RECT 1731.505 2793.930 1731.835 2793.945 ;
        RECT 1734.725 2793.940 1735.055 2793.945 ;
        RECT 1734.470 2793.930 1735.055 2793.940 ;
        RECT 1729.870 2793.630 1731.835 2793.930 ;
        RECT 1734.270 2793.630 1735.055 2793.930 ;
        RECT 1729.870 2793.620 1730.250 2793.630 ;
        RECT 1731.505 2793.615 1731.835 2793.630 ;
        RECT 1734.470 2793.620 1735.055 2793.630 ;
        RECT 1740.910 2793.930 1741.290 2793.940 ;
        RECT 1741.625 2793.930 1741.955 2793.945 ;
        RECT 1747.605 2793.940 1747.935 2793.945 ;
        RECT 1747.350 2793.930 1747.935 2793.940 ;
        RECT 1740.910 2793.630 1741.955 2793.930 ;
        RECT 1747.150 2793.630 1747.935 2793.930 ;
        RECT 1740.910 2793.620 1741.290 2793.630 ;
        RECT 1734.725 2793.615 1735.055 2793.620 ;
        RECT 1741.625 2793.615 1741.955 2793.630 ;
        RECT 1747.350 2793.620 1747.935 2793.630 ;
        RECT 1747.605 2793.615 1747.935 2793.620 ;
        RECT 1766.465 2793.930 1766.795 2793.945 ;
        RECT 1767.590 2793.930 1767.970 2793.940 ;
        RECT 1766.465 2793.630 1767.970 2793.930 ;
        RECT 1766.465 2793.615 1766.795 2793.630 ;
        RECT 1767.590 2793.620 1767.970 2793.630 ;
        RECT 1787.165 2793.930 1787.495 2793.945 ;
        RECT 1787.830 2793.930 1788.210 2793.940 ;
        RECT 1787.165 2793.630 1788.210 2793.930 ;
        RECT 1787.165 2793.615 1787.495 2793.630 ;
        RECT 1787.830 2793.620 1788.210 2793.630 ;
        RECT 2263.470 2793.930 2263.850 2793.940 ;
        RECT 2266.485 2793.930 2266.815 2793.945 ;
        RECT 2263.470 2793.630 2266.815 2793.930 ;
        RECT 2263.470 2793.620 2263.850 2793.630 ;
        RECT 2266.485 2793.615 2266.815 2793.630 ;
        RECT 2297.510 2793.930 2297.890 2793.940 ;
        RECT 2300.985 2793.930 2301.315 2793.945 ;
        RECT 2303.285 2793.930 2303.615 2793.945 ;
        RECT 2297.510 2793.630 2303.615 2793.930 ;
        RECT 2297.510 2793.620 2297.890 2793.630 ;
        RECT 2300.985 2793.615 2301.315 2793.630 ;
        RECT 2303.285 2793.615 2303.615 2793.630 ;
        RECT 2305.125 2793.930 2305.455 2793.945 ;
        RECT 2314.785 2793.940 2315.115 2793.945 ;
        RECT 2321.685 2793.940 2322.015 2793.945 ;
        RECT 2310.390 2793.930 2310.770 2793.940 ;
        RECT 2305.125 2793.630 2310.770 2793.930 ;
        RECT 2305.125 2793.615 2305.455 2793.630 ;
        RECT 2310.390 2793.620 2310.770 2793.630 ;
        RECT 2314.785 2793.930 2315.370 2793.940 ;
        RECT 2321.430 2793.930 2322.015 2793.940 ;
        RECT 2314.785 2793.630 2315.570 2793.930 ;
        RECT 2321.230 2793.630 2322.015 2793.930 ;
        RECT 2314.785 2793.620 2315.370 2793.630 ;
        RECT 2321.430 2793.620 2322.015 2793.630 ;
        RECT 2314.785 2793.615 2315.115 2793.620 ;
        RECT 2321.685 2793.615 2322.015 2793.620 ;
        RECT 2325.825 2793.940 2326.155 2793.945 ;
        RECT 2325.825 2793.930 2326.410 2793.940 ;
        RECT 2339.625 2793.930 2339.955 2793.945 ;
        RECT 2350.205 2793.940 2350.535 2793.945 ;
        RECT 2345.350 2793.930 2345.730 2793.940 ;
        RECT 2349.950 2793.930 2350.535 2793.940 ;
        RECT 2325.825 2793.630 2326.610 2793.930 ;
        RECT 2339.625 2793.630 2345.730 2793.930 ;
        RECT 2349.750 2793.630 2350.535 2793.930 ;
        RECT 2325.825 2793.620 2326.410 2793.630 ;
        RECT 2325.825 2793.615 2326.155 2793.620 ;
        RECT 2339.625 2793.615 2339.955 2793.630 ;
        RECT 2345.350 2793.620 2345.730 2793.630 ;
        RECT 2349.950 2793.620 2350.535 2793.630 ;
        RECT 2350.205 2793.615 2350.535 2793.620 ;
        RECT 2356.185 2793.940 2356.515 2793.945 ;
        RECT 2361.245 2793.940 2361.575 2793.945 ;
        RECT 2367.685 2793.940 2368.015 2793.945 ;
        RECT 2374.125 2793.940 2374.455 2793.945 ;
        RECT 2377.805 2793.940 2378.135 2793.945 ;
        RECT 2356.185 2793.930 2356.770 2793.940 ;
        RECT 2360.990 2793.930 2361.575 2793.940 ;
        RECT 2367.430 2793.930 2368.015 2793.940 ;
        RECT 2373.870 2793.930 2374.455 2793.940 ;
        RECT 2356.185 2793.630 2356.970 2793.930 ;
        RECT 2360.790 2793.630 2361.575 2793.930 ;
        RECT 2367.230 2793.630 2368.015 2793.930 ;
        RECT 2373.670 2793.630 2374.455 2793.930 ;
        RECT 2356.185 2793.620 2356.770 2793.630 ;
        RECT 2360.990 2793.620 2361.575 2793.630 ;
        RECT 2367.430 2793.620 2368.015 2793.630 ;
        RECT 2373.870 2793.620 2374.455 2793.630 ;
        RECT 2377.550 2793.930 2378.135 2793.940 ;
        RECT 2402.185 2793.940 2402.515 2793.945 ;
        RECT 2402.185 2793.930 2402.770 2793.940 ;
        RECT 2377.550 2793.630 2378.360 2793.930 ;
        RECT 2401.960 2793.630 2402.770 2793.930 ;
        RECT 2377.550 2793.620 2378.135 2793.630 ;
        RECT 2356.185 2793.615 2356.515 2793.620 ;
        RECT 2361.245 2793.615 2361.575 2793.620 ;
        RECT 2367.685 2793.615 2368.015 2793.620 ;
        RECT 2374.125 2793.615 2374.455 2793.620 ;
        RECT 2377.805 2793.615 2378.135 2793.620 ;
        RECT 2402.185 2793.620 2402.770 2793.630 ;
        RECT 2421.965 2793.930 2422.295 2793.945 ;
        RECT 2423.550 2793.930 2423.930 2793.940 ;
        RECT 2421.965 2793.630 2423.930 2793.930 ;
        RECT 2402.185 2793.615 2402.515 2793.620 ;
        RECT 2421.965 2793.615 2422.295 2793.630 ;
        RECT 2423.550 2793.620 2423.930 2793.630 ;
        RECT 509.285 2793.260 509.615 2793.265 ;
        RECT 509.030 2793.250 509.615 2793.260 ;
        RECT 508.830 2792.950 509.615 2793.250 ;
        RECT 509.030 2792.940 509.615 2792.950 ;
        RECT 509.285 2792.935 509.615 2792.940 ;
        RECT 986.765 2793.250 987.095 2793.265 ;
        RECT 987.430 2793.250 987.810 2793.260 ;
        RECT 986.765 2792.950 987.810 2793.250 ;
        RECT 986.765 2792.935 987.095 2792.950 ;
        RECT 987.430 2792.940 987.810 2792.950 ;
        RECT 1017.585 2793.250 1017.915 2793.265 ;
        RECT 1018.710 2793.250 1019.090 2793.260 ;
        RECT 1017.585 2792.950 1019.090 2793.250 ;
        RECT 1017.585 2792.935 1017.915 2792.950 ;
        RECT 1018.710 2792.940 1019.090 2792.950 ;
        RECT 1045.185 2793.250 1045.515 2793.265 ;
        RECT 1048.150 2793.250 1048.530 2793.260 ;
        RECT 1045.185 2792.950 1048.530 2793.250 ;
        RECT 1045.185 2792.935 1045.515 2792.950 ;
        RECT 1048.150 2792.940 1048.530 2792.950 ;
        RECT 1152.365 2793.250 1152.695 2793.265 ;
        RECT 1159.265 2793.260 1159.595 2793.265 ;
        RECT 1173.065 2793.260 1173.395 2793.265 ;
        RECT 1153.030 2793.250 1153.410 2793.260 ;
        RECT 1159.265 2793.250 1159.850 2793.260 ;
        RECT 1173.065 2793.250 1173.650 2793.260 ;
        RECT 1152.365 2792.950 1153.410 2793.250 ;
        RECT 1159.040 2792.950 1159.850 2793.250 ;
        RECT 1172.840 2792.950 1173.650 2793.250 ;
        RECT 1152.365 2792.935 1152.695 2792.950 ;
        RECT 1153.030 2792.940 1153.410 2792.950 ;
        RECT 1159.265 2792.940 1159.850 2792.950 ;
        RECT 1173.065 2792.940 1173.650 2792.950 ;
        RECT 1617.630 2793.250 1618.010 2793.260 ;
        RECT 1618.345 2793.250 1618.675 2793.265 ;
        RECT 1617.630 2792.950 1618.675 2793.250 ;
        RECT 1617.630 2792.940 1618.010 2792.950 ;
        RECT 1159.265 2792.935 1159.595 2792.940 ;
        RECT 1173.065 2792.935 1173.395 2792.940 ;
        RECT 1618.345 2792.935 1618.675 2792.950 ;
        RECT 1624.070 2793.250 1624.450 2793.260 ;
        RECT 1624.785 2793.250 1625.115 2793.265 ;
        RECT 1624.070 2792.950 1625.115 2793.250 ;
        RECT 1624.070 2792.940 1624.450 2792.950 ;
        RECT 1624.785 2792.935 1625.115 2792.950 ;
        RECT 1630.510 2793.250 1630.890 2793.260 ;
        RECT 1631.685 2793.250 1632.015 2793.265 ;
        RECT 1630.510 2792.950 1632.015 2793.250 ;
        RECT 1630.510 2792.940 1630.890 2792.950 ;
        RECT 1631.685 2792.935 1632.015 2792.950 ;
        RECT 1646.405 2793.250 1646.735 2793.265 ;
        RECT 1652.385 2793.260 1652.715 2793.265 ;
        RECT 1780.265 2793.260 1780.595 2793.265 ;
        RECT 2280.285 2793.260 2280.615 2793.265 ;
        RECT 1647.990 2793.250 1648.370 2793.260 ;
        RECT 1646.405 2792.950 1648.370 2793.250 ;
        RECT 1646.405 2792.935 1646.735 2792.950 ;
        RECT 1647.990 2792.940 1648.370 2792.950 ;
        RECT 1652.385 2793.250 1652.970 2793.260 ;
        RECT 1780.265 2793.250 1780.850 2793.260 ;
        RECT 2280.030 2793.250 2280.615 2793.260 ;
        RECT 1652.385 2792.950 1653.170 2793.250 ;
        RECT 1780.040 2792.950 1780.850 2793.250 ;
        RECT 2279.830 2792.950 2280.615 2793.250 ;
        RECT 1652.385 2792.940 1652.970 2792.950 ;
        RECT 1780.265 2792.940 1780.850 2792.950 ;
        RECT 2280.030 2792.940 2280.615 2792.950 ;
        RECT 2286.470 2793.250 2286.850 2793.260 ;
        RECT 2287.185 2793.250 2287.515 2793.265 ;
        RECT 2304.205 2793.260 2304.535 2793.265 ;
        RECT 2332.725 2793.260 2333.055 2793.265 ;
        RECT 2303.950 2793.250 2304.535 2793.260 ;
        RECT 2332.470 2793.250 2333.055 2793.260 ;
        RECT 2286.470 2792.950 2287.515 2793.250 ;
        RECT 2303.750 2792.950 2304.535 2793.250 ;
        RECT 2332.270 2792.950 2333.055 2793.250 ;
        RECT 2286.470 2792.940 2286.850 2792.950 ;
        RECT 1652.385 2792.935 1652.715 2792.940 ;
        RECT 1780.265 2792.935 1780.595 2792.940 ;
        RECT 2280.285 2792.935 2280.615 2792.940 ;
        RECT 2287.185 2792.935 2287.515 2792.950 ;
        RECT 2303.950 2792.940 2304.535 2792.950 ;
        RECT 2332.470 2792.940 2333.055 2792.950 ;
        RECT 2338.910 2793.250 2339.290 2793.260 ;
        RECT 2340.085 2793.250 2340.415 2793.265 ;
        RECT 2415.065 2793.260 2415.395 2793.265 ;
        RECT 2442.665 2793.260 2442.995 2793.265 ;
        RECT 2415.065 2793.250 2415.650 2793.260 ;
        RECT 2442.665 2793.250 2443.250 2793.260 ;
        RECT 2338.910 2792.950 2340.415 2793.250 ;
        RECT 2414.840 2792.950 2415.650 2793.250 ;
        RECT 2442.440 2792.950 2443.250 2793.250 ;
        RECT 2338.910 2792.940 2339.290 2792.950 ;
        RECT 2304.205 2792.935 2304.535 2792.940 ;
        RECT 2332.725 2792.935 2333.055 2792.940 ;
        RECT 2340.085 2792.935 2340.415 2792.950 ;
        RECT 2415.065 2792.940 2415.650 2792.950 ;
        RECT 2442.665 2792.940 2443.250 2792.950 ;
        RECT 2415.065 2792.935 2415.395 2792.940 ;
        RECT 2442.665 2792.935 2442.995 2792.940 ;
        RECT 993.665 2792.580 993.995 2792.585 ;
        RECT 1001.025 2792.580 1001.355 2792.585 ;
        RECT 1186.865 2792.580 1187.195 2792.585 ;
        RECT 1193.765 2792.580 1194.095 2792.585 ;
        RECT 993.665 2792.570 994.250 2792.580 ;
        RECT 1001.025 2792.570 1001.610 2792.580 ;
        RECT 1186.865 2792.570 1187.450 2792.580 ;
        RECT 993.440 2792.270 994.250 2792.570 ;
        RECT 1000.800 2792.270 1001.610 2792.570 ;
        RECT 1186.640 2792.270 1187.450 2792.570 ;
        RECT 993.665 2792.260 994.250 2792.270 ;
        RECT 1001.025 2792.260 1001.610 2792.270 ;
        RECT 1186.865 2792.260 1187.450 2792.270 ;
        RECT 1193.510 2792.570 1194.095 2792.580 ;
        RECT 1587.065 2792.580 1587.395 2792.585 ;
        RECT 1587.065 2792.570 1587.650 2792.580 ;
        RECT 1193.510 2792.270 1194.320 2792.570 ;
        RECT 1586.840 2792.270 1587.650 2792.570 ;
        RECT 1193.510 2792.260 1194.095 2792.270 ;
        RECT 993.665 2792.255 993.995 2792.260 ;
        RECT 1001.025 2792.255 1001.355 2792.260 ;
        RECT 1186.865 2792.255 1187.195 2792.260 ;
        RECT 1193.765 2792.255 1194.095 2792.260 ;
        RECT 1587.065 2792.260 1587.650 2792.270 ;
        RECT 1684.125 2792.570 1684.455 2792.585 ;
        RECT 1752.665 2792.580 1752.995 2792.585 ;
        RECT 1689.390 2792.570 1689.770 2792.580 ;
        RECT 1684.125 2792.270 1689.770 2792.570 ;
        RECT 1587.065 2792.255 1587.395 2792.260 ;
        RECT 1684.125 2792.255 1684.455 2792.270 ;
        RECT 1689.390 2792.260 1689.770 2792.270 ;
        RECT 1752.665 2792.570 1753.250 2792.580 ;
        RECT 2277.065 2792.570 2277.395 2792.585 ;
        RECT 2408.165 2792.580 2408.495 2792.585 ;
        RECT 2282.790 2792.570 2283.170 2792.580 ;
        RECT 1752.665 2792.270 1753.450 2792.570 ;
        RECT 2277.065 2792.270 2283.170 2792.570 ;
        RECT 1752.665 2792.260 1753.250 2792.270 ;
        RECT 1752.665 2792.255 1752.995 2792.260 ;
        RECT 2277.065 2792.255 2277.395 2792.270 ;
        RECT 2282.790 2792.260 2283.170 2792.270 ;
        RECT 2407.910 2792.570 2408.495 2792.580 ;
        RECT 2435.765 2792.570 2436.095 2792.585 ;
        RECT 2436.430 2792.570 2436.810 2792.580 ;
        RECT 2407.910 2792.270 2408.720 2792.570 ;
        RECT 2435.765 2792.270 2436.810 2792.570 ;
        RECT 2407.910 2792.260 2408.495 2792.270 ;
        RECT 2408.165 2792.255 2408.495 2792.260 ;
        RECT 2435.765 2792.255 2436.095 2792.270 ;
        RECT 2436.430 2792.260 2436.810 2792.270 ;
        RECT 386.465 2791.890 386.795 2791.905 ;
        RECT 388.510 2791.890 388.890 2791.900 ;
        RECT 386.465 2791.590 388.890 2791.890 ;
        RECT 386.465 2791.575 386.795 2791.590 ;
        RECT 388.510 2791.580 388.890 2791.590 ;
        RECT 414.065 2791.890 414.395 2791.905 ;
        RECT 1649.165 2791.900 1649.495 2791.905 ;
        RECT 417.030 2791.890 417.410 2791.900 ;
        RECT 414.065 2791.590 417.410 2791.890 ;
        RECT 414.065 2791.575 414.395 2791.590 ;
        RECT 417.030 2791.580 417.410 2791.590 ;
        RECT 1648.910 2791.890 1649.495 2791.900 ;
        RECT 1773.365 2791.890 1773.695 2791.905 ;
        RECT 1774.030 2791.890 1774.410 2791.900 ;
        RECT 1648.910 2791.590 1649.720 2791.890 ;
        RECT 1773.365 2791.590 1774.410 2791.890 ;
        RECT 1648.910 2791.580 1649.495 2791.590 ;
        RECT 1649.165 2791.575 1649.495 2791.580 ;
        RECT 1773.365 2791.575 1773.695 2791.590 ;
        RECT 1774.030 2791.580 1774.410 2791.590 ;
        RECT 2270.165 2791.890 2270.495 2791.905 ;
        RECT 2276.350 2791.890 2276.730 2791.900 ;
        RECT 2270.165 2791.590 2276.730 2791.890 ;
        RECT 2270.165 2791.575 2270.495 2791.590 ;
        RECT 2276.350 2791.580 2276.730 2791.590 ;
        RECT 2283.965 2791.890 2284.295 2791.905 ;
        RECT 2287.390 2791.890 2287.770 2791.900 ;
        RECT 2283.965 2791.590 2287.770 2791.890 ;
        RECT 2283.965 2791.575 2284.295 2791.590 ;
        RECT 2287.390 2791.580 2287.770 2791.590 ;
        RECT 2290.865 2791.890 2291.195 2791.905 ;
        RECT 2293.830 2791.890 2294.210 2791.900 ;
        RECT 2290.865 2791.590 2294.210 2791.890 ;
        RECT 2290.865 2791.575 2291.195 2791.590 ;
        RECT 2293.830 2791.580 2294.210 2791.590 ;
        RECT 2442.665 2791.890 2442.995 2791.905 ;
        RECT 2445.630 2791.890 2446.010 2791.900 ;
        RECT 2442.665 2791.590 2446.010 2791.890 ;
        RECT 2442.665 2791.575 2442.995 2791.590 ;
        RECT 2445.630 2791.580 2446.010 2791.590 ;
        RECT 365.765 2791.210 366.095 2791.225 ;
        RECT 371.030 2791.210 371.410 2791.220 ;
        RECT 365.765 2790.910 371.410 2791.210 ;
        RECT 365.765 2790.895 366.095 2790.910 ;
        RECT 371.030 2790.900 371.410 2790.910 ;
        RECT 1642.265 2791.210 1642.595 2791.225 ;
        RECT 1644.310 2791.210 1644.690 2791.220 ;
        RECT 1642.265 2790.910 1644.690 2791.210 ;
        RECT 1642.265 2790.895 1642.595 2790.910 ;
        RECT 1644.310 2790.900 1644.690 2790.910 ;
        RECT 1656.065 2791.210 1656.395 2791.225 ;
        RECT 1661.790 2791.210 1662.170 2791.220 ;
        RECT 1656.065 2790.910 1662.170 2791.210 ;
        RECT 1656.065 2790.895 1656.395 2790.910 ;
        RECT 1661.790 2790.900 1662.170 2790.910 ;
        RECT 2263.265 2791.210 2263.595 2791.225 ;
        RECT 2268.990 2791.210 2269.370 2791.220 ;
        RECT 2263.265 2790.910 2269.370 2791.210 ;
        RECT 2263.265 2790.895 2263.595 2790.910 ;
        RECT 2268.990 2790.900 2269.370 2790.910 ;
        RECT 2297.765 2791.210 2298.095 2791.225 ;
        RECT 2299.350 2791.210 2299.730 2791.220 ;
        RECT 2297.765 2790.910 2299.730 2791.210 ;
        RECT 2297.765 2790.895 2298.095 2790.910 ;
        RECT 2299.350 2790.900 2299.730 2790.910 ;
        RECT 2415.065 2791.210 2415.395 2791.225 ;
        RECT 2420.790 2791.210 2421.170 2791.220 ;
        RECT 2415.065 2790.910 2421.170 2791.210 ;
        RECT 2415.065 2790.895 2415.395 2790.910 ;
        RECT 2420.790 2790.900 2421.170 2790.910 ;
        RECT 2428.865 2791.210 2429.195 2791.225 ;
        RECT 2434.590 2791.210 2434.970 2791.220 ;
        RECT 2428.865 2790.910 2434.970 2791.210 ;
        RECT 2428.865 2790.895 2429.195 2790.910 ;
        RECT 2434.590 2790.900 2434.970 2790.910 ;
        RECT 2435.765 2791.210 2436.095 2791.225 ;
        RECT 2439.190 2791.210 2439.570 2791.220 ;
        RECT 2435.765 2790.910 2439.570 2791.210 ;
        RECT 2435.765 2790.895 2436.095 2790.910 ;
        RECT 2439.190 2790.900 2439.570 2790.910 ;
        RECT 342.510 2790.530 342.890 2790.540 ;
        RECT 344.605 2790.530 344.935 2790.545 ;
        RECT 342.510 2790.230 344.935 2790.530 ;
        RECT 342.510 2790.220 342.890 2790.230 ;
        RECT 344.605 2790.215 344.935 2790.230 ;
        RECT 1030.670 2790.530 1031.050 2790.540 ;
        RECT 1031.385 2790.530 1031.715 2790.545 ;
        RECT 1030.670 2790.230 1031.715 2790.530 ;
        RECT 1030.670 2790.220 1031.050 2790.230 ;
        RECT 1031.385 2790.215 1031.715 2790.230 ;
        RECT 1191.670 2790.530 1192.050 2790.540 ;
        RECT 1193.305 2790.530 1193.635 2790.545 ;
        RECT 1191.670 2790.230 1193.635 2790.530 ;
        RECT 1191.670 2790.220 1192.050 2790.230 ;
        RECT 1193.305 2790.215 1193.635 2790.230 ;
        RECT 2380.565 2790.530 2380.895 2790.545 ;
        RECT 2386.750 2790.530 2387.130 2790.540 ;
        RECT 2380.565 2790.230 2387.130 2790.530 ;
        RECT 2380.565 2790.215 2380.895 2790.230 ;
        RECT 2386.750 2790.220 2387.130 2790.230 ;
        RECT 2387.465 2790.530 2387.795 2790.545 ;
        RECT 2392.270 2790.530 2392.650 2790.540 ;
        RECT 2387.465 2790.230 2392.650 2790.530 ;
        RECT 2387.465 2790.215 2387.795 2790.230 ;
        RECT 2392.270 2790.220 2392.650 2790.230 ;
        RECT 393.365 2789.860 393.695 2789.865 ;
        RECT 393.110 2789.850 393.695 2789.860 ;
        RECT 1614.665 2789.850 1614.995 2789.865 ;
        RECT 1620.390 2789.850 1620.770 2789.860 ;
        RECT 393.110 2789.550 393.920 2789.850 ;
        RECT 1614.665 2789.550 1620.770 2789.850 ;
        RECT 393.110 2789.540 393.695 2789.550 ;
        RECT 393.365 2789.535 393.695 2789.540 ;
        RECT 1614.665 2789.535 1614.995 2789.550 ;
        RECT 1620.390 2789.540 1620.770 2789.550 ;
        RECT 2394.365 2789.850 2394.695 2789.865 ;
        RECT 2398.710 2789.850 2399.090 2789.860 ;
        RECT 2394.365 2789.550 2399.090 2789.850 ;
        RECT 2394.365 2789.535 2394.695 2789.550 ;
        RECT 2398.710 2789.540 2399.090 2789.550 ;
        RECT 372.665 2789.170 372.995 2789.185 ;
        RECT 375.630 2789.170 376.010 2789.180 ;
        RECT 372.665 2788.870 376.010 2789.170 ;
        RECT 372.665 2788.855 372.995 2788.870 ;
        RECT 375.630 2788.860 376.010 2788.870 ;
        RECT 379.565 2789.170 379.895 2789.185 ;
        RECT 1600.865 2789.180 1601.195 2789.185 ;
        RECT 382.070 2789.170 382.450 2789.180 ;
        RECT 1600.865 2789.170 1601.450 2789.180 ;
        RECT 379.565 2788.870 382.450 2789.170 ;
        RECT 1600.640 2788.870 1601.450 2789.170 ;
        RECT 379.565 2788.855 379.895 2788.870 ;
        RECT 382.070 2788.860 382.450 2788.870 ;
        RECT 1600.865 2788.860 1601.450 2788.870 ;
        RECT 2408.165 2789.170 2408.495 2789.185 ;
        RECT 2410.670 2789.170 2411.050 2789.180 ;
        RECT 2408.165 2788.870 2411.050 2789.170 ;
        RECT 1600.865 2788.855 1601.195 2788.860 ;
        RECT 2408.165 2788.855 2408.495 2788.870 ;
        RECT 2410.670 2788.860 2411.050 2788.870 ;
        RECT 358.865 2788.490 359.195 2788.505 ;
        RECT 364.590 2788.490 364.970 2788.500 ;
        RECT 358.865 2788.190 364.970 2788.490 ;
        RECT 358.865 2788.175 359.195 2788.190 ;
        RECT 364.590 2788.180 364.970 2788.190 ;
        RECT 393.365 2788.490 393.695 2788.505 ;
        RECT 399.550 2788.490 399.930 2788.500 ;
        RECT 393.365 2788.190 399.930 2788.490 ;
        RECT 393.365 2788.175 393.695 2788.190 ;
        RECT 399.550 2788.180 399.930 2788.190 ;
        RECT 465.790 2788.490 466.170 2788.500 ;
        RECT 468.345 2788.490 468.675 2788.505 ;
        RECT 465.790 2788.190 468.675 2788.490 ;
        RECT 465.790 2788.180 466.170 2788.190 ;
        RECT 468.345 2788.175 468.675 2788.190 ;
        RECT 1035.270 2788.490 1035.650 2788.500 ;
        RECT 1038.285 2788.490 1038.615 2788.505 ;
        RECT 1035.270 2788.190 1038.615 2788.490 ;
        RECT 1035.270 2788.180 1035.650 2788.190 ;
        RECT 1038.285 2788.175 1038.615 2788.190 ;
        RECT 1041.710 2788.490 1042.090 2788.500 ;
        RECT 1046.105 2788.490 1046.435 2788.505 ;
        RECT 1041.710 2788.190 1046.435 2788.490 ;
        RECT 1041.710 2788.180 1042.090 2788.190 ;
        RECT 1046.105 2788.175 1046.435 2788.190 ;
        RECT 1051.830 2788.490 1052.210 2788.500 ;
        RECT 1054.845 2788.490 1055.175 2788.505 ;
        RECT 1051.830 2788.190 1055.175 2788.490 ;
        RECT 1051.830 2788.180 1052.210 2788.190 ;
        RECT 1054.845 2788.175 1055.175 2788.190 ;
        RECT 1718.625 2788.490 1718.955 2788.505 ;
        RECT 1724.350 2788.490 1724.730 2788.500 ;
        RECT 1718.625 2788.190 1724.730 2788.490 ;
        RECT 1718.625 2788.175 1718.955 2788.190 ;
        RECT 1724.350 2788.180 1724.730 2788.190 ;
        RECT 1760.025 2788.490 1760.355 2788.505 ;
        RECT 2256.825 2788.500 2257.155 2788.505 ;
        RECT 1765.750 2788.490 1766.130 2788.500 ;
        RECT 2256.825 2788.490 2257.410 2788.500 ;
        RECT 1760.025 2788.190 1766.130 2788.490 ;
        RECT 2256.600 2788.190 2257.410 2788.490 ;
        RECT 1760.025 2788.175 1760.355 2788.190 ;
        RECT 1765.750 2788.180 1766.130 2788.190 ;
        RECT 2256.825 2788.180 2257.410 2788.190 ;
        RECT 2373.205 2788.490 2373.535 2788.505 ;
        RECT 2377.550 2788.490 2377.930 2788.500 ;
        RECT 2373.205 2788.190 2377.930 2788.490 ;
        RECT 2256.825 2788.175 2257.155 2788.180 ;
        RECT 2373.205 2788.175 2373.535 2788.190 ;
        RECT 2377.550 2788.180 2377.930 2788.190 ;
        RECT 2415.065 2788.490 2415.395 2788.505 ;
        RECT 2418.030 2788.490 2418.410 2788.500 ;
        RECT 2415.065 2788.190 2418.410 2788.490 ;
        RECT 2415.065 2788.175 2415.395 2788.190 ;
        RECT 2418.030 2788.180 2418.410 2788.190 ;
        RECT 357.230 2787.810 357.610 2787.820 ;
        RECT 357.945 2787.810 358.275 2787.825 ;
        RECT 455.005 2787.820 455.335 2787.825 ;
        RECT 357.230 2787.510 358.275 2787.810 ;
        RECT 357.230 2787.500 357.610 2787.510 ;
        RECT 357.945 2787.495 358.275 2787.510 ;
        RECT 454.750 2787.810 455.335 2787.820 ;
        RECT 460.270 2787.810 460.650 2787.820 ;
        RECT 461.905 2787.810 462.235 2787.825 ;
        RECT 468.805 2787.820 469.135 2787.825 ;
        RECT 454.750 2787.510 455.560 2787.810 ;
        RECT 460.270 2787.510 462.235 2787.810 ;
        RECT 454.750 2787.500 455.335 2787.510 ;
        RECT 460.270 2787.500 460.650 2787.510 ;
        RECT 455.005 2787.495 455.335 2787.500 ;
        RECT 461.905 2787.495 462.235 2787.510 ;
        RECT 468.550 2787.810 469.135 2787.820 ;
        RECT 474.990 2787.810 475.370 2787.820 ;
        RECT 475.705 2787.810 476.035 2787.825 ;
        RECT 482.605 2787.820 482.935 2787.825 ;
        RECT 468.550 2787.510 469.360 2787.810 ;
        RECT 474.990 2787.510 476.035 2787.810 ;
        RECT 468.550 2787.500 469.135 2787.510 ;
        RECT 474.990 2787.500 475.370 2787.510 ;
        RECT 468.805 2787.495 469.135 2787.500 ;
        RECT 475.705 2787.495 476.035 2787.510 ;
        RECT 482.350 2787.810 482.935 2787.820 ;
        RECT 488.790 2787.810 489.170 2787.820 ;
        RECT 489.505 2787.810 489.835 2787.825 ;
        RECT 482.350 2787.510 483.160 2787.810 ;
        RECT 488.790 2787.510 489.835 2787.810 ;
        RECT 482.350 2787.500 482.935 2787.510 ;
        RECT 488.790 2787.500 489.170 2787.510 ;
        RECT 482.605 2787.495 482.935 2787.500 ;
        RECT 489.505 2787.495 489.835 2787.510 ;
        RECT 495.230 2787.810 495.610 2787.820 ;
        RECT 496.405 2787.810 496.735 2787.825 ;
        RECT 1034.605 2787.820 1034.935 2787.825 ;
        RECT 495.230 2787.510 496.735 2787.810 ;
        RECT 495.230 2787.500 495.610 2787.510 ;
        RECT 496.405 2787.495 496.735 2787.510 ;
        RECT 1034.350 2787.810 1034.935 2787.820 ;
        RECT 1039.870 2787.810 1040.250 2787.820 ;
        RECT 1041.505 2787.810 1041.835 2787.825 ;
        RECT 1034.350 2787.510 1035.160 2787.810 ;
        RECT 1039.870 2787.510 1041.835 2787.810 ;
        RECT 1034.350 2787.500 1034.935 2787.510 ;
        RECT 1039.870 2787.500 1040.250 2787.510 ;
        RECT 1034.605 2787.495 1034.935 2787.500 ;
        RECT 1041.505 2787.495 1041.835 2787.510 ;
        RECT 1046.310 2787.810 1046.690 2787.820 ;
        RECT 1048.405 2787.810 1048.735 2787.825 ;
        RECT 1062.205 2787.820 1062.535 2787.825 ;
        RECT 1046.310 2787.510 1048.735 2787.810 ;
        RECT 1046.310 2787.500 1046.690 2787.510 ;
        RECT 1048.405 2787.495 1048.735 2787.510 ;
        RECT 1061.950 2787.810 1062.535 2787.820 ;
        RECT 1067.470 2787.810 1067.850 2787.820 ;
        RECT 1069.105 2787.810 1069.435 2787.825 ;
        RECT 1061.950 2787.510 1062.760 2787.810 ;
        RECT 1067.470 2787.510 1069.435 2787.810 ;
        RECT 1061.950 2787.500 1062.535 2787.510 ;
        RECT 1067.470 2787.500 1067.850 2787.510 ;
        RECT 1062.205 2787.495 1062.535 2787.500 ;
        RECT 1069.105 2787.495 1069.435 2787.510 ;
        RECT 1073.910 2787.810 1074.290 2787.820 ;
        RECT 1076.005 2787.810 1076.335 2787.825 ;
        RECT 1073.910 2787.510 1076.335 2787.810 ;
        RECT 1073.910 2787.500 1074.290 2787.510 ;
        RECT 1076.005 2787.495 1076.335 2787.510 ;
        RECT 1752.665 2787.810 1752.995 2787.825 ;
        RECT 1754.710 2787.810 1755.090 2787.820 ;
        RECT 1752.665 2787.510 1755.090 2787.810 ;
        RECT 1752.665 2787.495 1752.995 2787.510 ;
        RECT 1754.710 2787.500 1755.090 2787.510 ;
        RECT 1766.465 2787.810 1766.795 2787.825 ;
        RECT 1772.190 2787.810 1772.570 2787.820 ;
        RECT 1766.465 2787.510 1772.570 2787.810 ;
        RECT 1766.465 2787.495 1766.795 2787.510 ;
        RECT 1772.190 2787.500 1772.570 2787.510 ;
        RECT 1773.825 2787.810 1774.155 2787.825 ;
        RECT 1777.710 2787.810 1778.090 2787.820 ;
        RECT 1773.825 2787.510 1778.090 2787.810 ;
        RECT 1773.825 2787.495 1774.155 2787.510 ;
        RECT 1777.710 2787.500 1778.090 2787.510 ;
        RECT 1780.265 2787.810 1780.595 2787.825 ;
        RECT 1783.230 2787.810 1783.610 2787.820 ;
        RECT 1780.265 2787.510 1783.610 2787.810 ;
        RECT 1780.265 2787.495 1780.595 2787.510 ;
        RECT 1783.230 2787.500 1783.610 2787.510 ;
        RECT 1787.165 2787.810 1787.495 2787.825 ;
        RECT 1789.670 2787.810 1790.050 2787.820 ;
        RECT 1787.165 2787.510 1790.050 2787.810 ;
        RECT 1787.165 2787.495 1787.495 2787.510 ;
        RECT 1789.670 2787.500 1790.050 2787.510 ;
        RECT 1760.945 2777.620 1761.275 2777.625 ;
        RECT 1760.945 2777.610 1761.530 2777.620 ;
        RECT 1760.720 2777.310 1761.530 2777.610 ;
        RECT 1760.945 2777.300 1761.530 2777.310 ;
        RECT 1794.065 2777.610 1794.395 2777.625 ;
        RECT 1796.110 2777.610 1796.490 2777.620 ;
        RECT 1794.065 2777.310 1796.490 2777.610 ;
        RECT 1760.945 2777.295 1761.275 2777.300 ;
        RECT 1794.065 2777.295 1794.395 2777.310 ;
        RECT 1796.110 2777.300 1796.490 2777.310 ;
        RECT 1056.225 2753.130 1056.555 2753.145 ;
        RECT 1057.145 2753.130 1057.475 2753.145 ;
        RECT 1056.225 2752.830 1057.475 2753.130 ;
        RECT 1056.225 2752.815 1056.555 2752.830 ;
        RECT 1057.145 2752.815 1057.475 2752.830 ;
        RECT 282.965 2715.050 283.295 2715.065 ;
        RECT 792.645 2715.050 792.975 2715.065 ;
        RECT 282.965 2714.750 792.975 2715.050 ;
        RECT 282.965 2714.735 283.295 2714.750 ;
        RECT 792.645 2714.735 792.975 2714.750 ;
        RECT 1396.000 2694.650 1400.000 2694.720 ;
        RECT 1408.585 2694.650 1408.915 2694.665 ;
      LAYER met3 ;
        RECT 304.400 2693.720 1395.600 2694.585 ;
      LAYER met3 ;
        RECT 1396.000 2694.350 1408.915 2694.650 ;
        RECT 1396.000 2694.120 1400.000 2694.350 ;
        RECT 1408.585 2694.335 1408.915 2694.350 ;
      LAYER met3 ;
        RECT 303.990 2684.920 1396.000 2693.720 ;
        RECT 304.400 2684.240 1396.000 2684.920 ;
        RECT 304.400 2683.520 1395.600 2684.240 ;
        RECT 303.990 2682.840 1395.600 2683.520 ;
      LAYER met3 ;
        RECT 1396.000 2683.770 1400.000 2683.840 ;
        RECT 1414.105 2683.770 1414.435 2683.785 ;
        RECT 1396.000 2683.470 1414.435 2683.770 ;
        RECT 1396.000 2683.240 1400.000 2683.470 ;
        RECT 1414.105 2683.455 1414.435 2683.470 ;
      LAYER met3 ;
        RECT 303.990 2674.040 1396.000 2682.840 ;
        RECT 304.400 2673.360 1396.000 2674.040 ;
        RECT 304.400 2672.640 1395.600 2673.360 ;
        RECT 303.990 2671.960 1395.600 2672.640 ;
      LAYER met3 ;
        RECT 1396.000 2672.890 1400.000 2672.960 ;
        RECT 1414.105 2672.890 1414.435 2672.905 ;
        RECT 1396.000 2672.590 1414.435 2672.890 ;
        RECT 1396.000 2672.360 1400.000 2672.590 ;
        RECT 1414.105 2672.575 1414.435 2672.590 ;
      LAYER met3 ;
        RECT 303.990 2663.840 1396.000 2671.960 ;
        RECT 304.400 2662.480 1396.000 2663.840 ;
        RECT 304.400 2662.440 1395.600 2662.480 ;
        RECT 303.990 2661.080 1395.600 2662.440 ;
      LAYER met3 ;
        RECT 1396.000 2662.010 1400.000 2662.080 ;
        RECT 1414.105 2662.010 1414.435 2662.025 ;
        RECT 1396.000 2661.710 1414.435 2662.010 ;
        RECT 1396.000 2661.480 1400.000 2661.710 ;
        RECT 1414.105 2661.695 1414.435 2661.710 ;
      LAYER met3 ;
        RECT 303.990 2652.960 1396.000 2661.080 ;
        RECT 304.400 2651.600 1396.000 2652.960 ;
        RECT 304.400 2651.560 1395.600 2651.600 ;
        RECT 303.990 2650.200 1395.600 2651.560 ;
      LAYER met3 ;
        RECT 1396.000 2651.130 1400.000 2651.200 ;
        RECT 1414.105 2651.130 1414.435 2651.145 ;
        RECT 1396.000 2650.830 1414.435 2651.130 ;
        RECT 1396.000 2650.600 1400.000 2650.830 ;
        RECT 1414.105 2650.815 1414.435 2650.830 ;
      LAYER met3 ;
        RECT 303.990 2642.760 1396.000 2650.200 ;
        RECT 304.400 2641.360 1396.000 2642.760 ;
        RECT 303.990 2640.040 1396.000 2641.360 ;
        RECT 303.990 2638.640 1395.600 2640.040 ;
      LAYER met3 ;
        RECT 1396.000 2639.570 1400.000 2639.640 ;
        RECT 1414.105 2639.570 1414.435 2639.585 ;
        RECT 1396.000 2639.270 1414.435 2639.570 ;
        RECT 1396.000 2639.040 1400.000 2639.270 ;
        RECT 1414.105 2639.255 1414.435 2639.270 ;
      LAYER met3 ;
        RECT 303.990 2631.880 1396.000 2638.640 ;
        RECT 304.400 2630.480 1396.000 2631.880 ;
        RECT 303.990 2629.160 1396.000 2630.480 ;
        RECT 303.990 2627.760 1395.600 2629.160 ;
      LAYER met3 ;
        RECT 1396.000 2628.690 1400.000 2628.760 ;
        RECT 1414.105 2628.690 1414.435 2628.705 ;
        RECT 1396.000 2628.390 1414.435 2628.690 ;
        RECT 1396.000 2628.160 1400.000 2628.390 ;
        RECT 1414.105 2628.375 1414.435 2628.390 ;
      LAYER met3 ;
        RECT 303.990 2621.680 1396.000 2627.760 ;
        RECT 304.400 2620.280 1396.000 2621.680 ;
        RECT 303.990 2618.280 1396.000 2620.280 ;
        RECT 303.990 2616.880 1395.600 2618.280 ;
      LAYER met3 ;
        RECT 1396.000 2617.810 1400.000 2617.880 ;
        RECT 1414.105 2617.810 1414.435 2617.825 ;
        RECT 1396.000 2617.510 1414.435 2617.810 ;
        RECT 1396.000 2617.280 1400.000 2617.510 ;
        RECT 1414.105 2617.495 1414.435 2617.510 ;
      LAYER met3 ;
        RECT 303.990 2610.800 1396.000 2616.880 ;
        RECT 304.400 2609.400 1396.000 2610.800 ;
        RECT 303.990 2607.400 1396.000 2609.400 ;
        RECT 303.990 2606.000 1395.600 2607.400 ;
      LAYER met3 ;
        RECT 1396.000 2606.930 1400.000 2607.000 ;
        RECT 1414.105 2606.930 1414.435 2606.945 ;
        RECT 1396.000 2606.630 1414.435 2606.930 ;
        RECT 1396.000 2606.400 1400.000 2606.630 ;
        RECT 1414.105 2606.615 1414.435 2606.630 ;
      LAYER met3 ;
        RECT 303.990 2600.600 1396.000 2606.000 ;
        RECT 304.400 2599.200 1396.000 2600.600 ;
        RECT 303.990 2596.520 1396.000 2599.200 ;
        RECT 303.990 2595.120 1395.600 2596.520 ;
      LAYER met3 ;
        RECT 1396.000 2596.050 1400.000 2596.120 ;
        RECT 1414.105 2596.050 1414.435 2596.065 ;
        RECT 1396.000 2595.750 1414.435 2596.050 ;
        RECT 1396.000 2595.520 1400.000 2595.750 ;
        RECT 1414.105 2595.735 1414.435 2595.750 ;
      LAYER met3 ;
        RECT 303.990 2589.720 1396.000 2595.120 ;
        RECT 304.400 2588.320 1396.000 2589.720 ;
        RECT 303.990 2584.960 1396.000 2588.320 ;
        RECT 303.990 2583.560 1395.600 2584.960 ;
      LAYER met3 ;
        RECT 1396.000 2584.490 1400.000 2584.560 ;
        RECT 1409.505 2584.490 1409.835 2584.505 ;
        RECT 1396.000 2584.190 1409.835 2584.490 ;
        RECT 1396.000 2583.960 1400.000 2584.190 ;
        RECT 1409.505 2584.175 1409.835 2584.190 ;
      LAYER met3 ;
        RECT 303.990 2579.520 1396.000 2583.560 ;
        RECT 304.400 2578.120 1396.000 2579.520 ;
        RECT 303.990 2574.080 1396.000 2578.120 ;
        RECT 303.990 2572.680 1395.600 2574.080 ;
      LAYER met3 ;
        RECT 1396.000 2573.610 1400.000 2573.680 ;
        RECT 1414.105 2573.610 1414.435 2573.625 ;
        RECT 1396.000 2573.310 1414.435 2573.610 ;
        RECT 1396.000 2573.080 1400.000 2573.310 ;
        RECT 1414.105 2573.295 1414.435 2573.310 ;
      LAYER met3 ;
        RECT 303.990 2568.640 1396.000 2572.680 ;
        RECT 304.400 2567.240 1396.000 2568.640 ;
        RECT 303.990 2563.200 1396.000 2567.240 ;
        RECT 303.990 2561.800 1395.600 2563.200 ;
      LAYER met3 ;
        RECT 1396.000 2562.730 1400.000 2562.800 ;
        RECT 1410.425 2562.730 1410.755 2562.745 ;
        RECT 1396.000 2562.430 1410.755 2562.730 ;
        RECT 1396.000 2562.200 1400.000 2562.430 ;
        RECT 1410.425 2562.415 1410.755 2562.430 ;
      LAYER met3 ;
        RECT 303.990 2558.440 1396.000 2561.800 ;
        RECT 304.400 2557.040 1396.000 2558.440 ;
        RECT 303.990 2552.320 1396.000 2557.040 ;
        RECT 303.990 2550.920 1395.600 2552.320 ;
      LAYER met3 ;
        RECT 1396.000 2551.850 1400.000 2551.920 ;
        RECT 1414.105 2551.850 1414.435 2551.865 ;
        RECT 1396.000 2551.550 1414.435 2551.850 ;
        RECT 1396.000 2551.320 1400.000 2551.550 ;
        RECT 1414.105 2551.535 1414.435 2551.550 ;
      LAYER met3 ;
        RECT 303.990 2547.560 1396.000 2550.920 ;
        RECT 304.400 2546.160 1396.000 2547.560 ;
        RECT 303.990 2541.440 1396.000 2546.160 ;
        RECT 303.990 2540.040 1395.600 2541.440 ;
      LAYER met3 ;
        RECT 1396.000 2540.970 1400.000 2541.040 ;
        RECT 1411.345 2540.970 1411.675 2540.985 ;
        RECT 1396.000 2540.670 1411.675 2540.970 ;
        RECT 1396.000 2540.440 1400.000 2540.670 ;
        RECT 1411.345 2540.655 1411.675 2540.670 ;
      LAYER met3 ;
        RECT 303.990 2537.360 1396.000 2540.040 ;
        RECT 304.400 2535.960 1396.000 2537.360 ;
        RECT 303.990 2529.880 1396.000 2535.960 ;
        RECT 303.990 2528.480 1395.600 2529.880 ;
      LAYER met3 ;
        RECT 1396.000 2529.410 1400.000 2529.480 ;
        RECT 1409.505 2529.410 1409.835 2529.425 ;
        RECT 1396.000 2529.110 1409.835 2529.410 ;
        RECT 1396.000 2528.880 1400.000 2529.110 ;
        RECT 1409.505 2529.095 1409.835 2529.110 ;
      LAYER met3 ;
        RECT 303.990 2526.480 1396.000 2528.480 ;
        RECT 304.400 2525.080 1396.000 2526.480 ;
        RECT 303.990 2519.000 1396.000 2525.080 ;
        RECT 303.990 2517.600 1395.600 2519.000 ;
      LAYER met3 ;
        RECT 1396.000 2518.530 1400.000 2518.600 ;
        RECT 1414.105 2518.530 1414.435 2518.545 ;
        RECT 1396.000 2518.230 1414.435 2518.530 ;
        RECT 1396.000 2518.000 1400.000 2518.230 ;
        RECT 1414.105 2518.215 1414.435 2518.230 ;
      LAYER met3 ;
        RECT 303.990 2516.280 1396.000 2517.600 ;
        RECT 304.400 2514.880 1396.000 2516.280 ;
        RECT 303.990 2508.120 1396.000 2514.880 ;
        RECT 303.990 2506.720 1395.600 2508.120 ;
      LAYER met3 ;
        RECT 1396.000 2507.650 1400.000 2507.720 ;
        RECT 1410.425 2507.650 1410.755 2507.665 ;
        RECT 1396.000 2507.350 1410.755 2507.650 ;
        RECT 1396.000 2507.120 1400.000 2507.350 ;
        RECT 1410.425 2507.335 1410.755 2507.350 ;
      LAYER met3 ;
        RECT 303.990 2505.400 1396.000 2506.720 ;
        RECT 304.400 2504.000 1396.000 2505.400 ;
        RECT 303.990 2497.240 1396.000 2504.000 ;
        RECT 303.990 2495.840 1395.600 2497.240 ;
      LAYER met3 ;
        RECT 1396.000 2496.770 1400.000 2496.840 ;
        RECT 1414.105 2496.770 1414.435 2496.785 ;
        RECT 1396.000 2496.470 1414.435 2496.770 ;
        RECT 1396.000 2496.240 1400.000 2496.470 ;
        RECT 1414.105 2496.455 1414.435 2496.470 ;
      LAYER met3 ;
        RECT 303.990 2495.200 1396.000 2495.840 ;
        RECT 304.400 2493.800 1396.000 2495.200 ;
        RECT 303.990 2486.360 1396.000 2493.800 ;
        RECT 303.990 2484.960 1395.600 2486.360 ;
      LAYER met3 ;
        RECT 1396.000 2485.890 1400.000 2485.960 ;
        RECT 1411.345 2485.890 1411.675 2485.905 ;
        RECT 1396.000 2485.590 1411.675 2485.890 ;
        RECT 1396.000 2485.360 1400.000 2485.590 ;
        RECT 1411.345 2485.575 1411.675 2485.590 ;
      LAYER met3 ;
        RECT 303.990 2484.320 1396.000 2484.960 ;
        RECT 304.400 2482.920 1396.000 2484.320 ;
        RECT 303.990 2474.800 1396.000 2482.920 ;
        RECT 303.990 2474.120 1395.600 2474.800 ;
        RECT 304.400 2473.400 1395.600 2474.120 ;
      LAYER met3 ;
        RECT 1396.000 2474.330 1400.000 2474.400 ;
        RECT 1409.505 2474.330 1409.835 2474.345 ;
        RECT 1396.000 2474.030 1409.835 2474.330 ;
        RECT 1396.000 2473.800 1400.000 2474.030 ;
        RECT 1409.505 2474.015 1409.835 2474.030 ;
      LAYER met3 ;
        RECT 304.400 2472.720 1396.000 2473.400 ;
        RECT 303.990 2463.920 1396.000 2472.720 ;
        RECT 303.990 2463.240 1395.600 2463.920 ;
        RECT 304.400 2462.520 1395.600 2463.240 ;
      LAYER met3 ;
        RECT 1396.000 2463.450 1400.000 2463.520 ;
        RECT 1412.265 2463.450 1412.595 2463.465 ;
        RECT 1396.000 2463.150 1412.595 2463.450 ;
        RECT 1396.000 2462.920 1400.000 2463.150 ;
        RECT 1412.265 2463.135 1412.595 2463.150 ;
      LAYER met3 ;
        RECT 304.400 2461.840 1396.000 2462.520 ;
        RECT 303.990 2453.040 1396.000 2461.840 ;
        RECT 304.400 2451.640 1395.600 2453.040 ;
      LAYER met3 ;
        RECT 1396.000 2452.570 1400.000 2452.640 ;
        RECT 1410.425 2452.570 1410.755 2452.585 ;
        RECT 1396.000 2452.270 1410.755 2452.570 ;
        RECT 1396.000 2452.040 1400.000 2452.270 ;
        RECT 1410.425 2452.255 1410.755 2452.270 ;
      LAYER met3 ;
        RECT 303.990 2442.160 1396.000 2451.640 ;
        RECT 304.400 2440.760 1395.600 2442.160 ;
      LAYER met3 ;
        RECT 1396.000 2441.690 1400.000 2441.760 ;
        RECT 1414.105 2441.690 1414.435 2441.705 ;
        RECT 1396.000 2441.390 1414.435 2441.690 ;
        RECT 1396.000 2441.160 1400.000 2441.390 ;
        RECT 1414.105 2441.375 1414.435 2441.390 ;
      LAYER met3 ;
        RECT 303.990 2431.960 1396.000 2440.760 ;
        RECT 304.400 2431.280 1396.000 2431.960 ;
        RECT 304.400 2430.560 1395.600 2431.280 ;
        RECT 303.990 2429.880 1395.600 2430.560 ;
      LAYER met3 ;
        RECT 1396.000 2430.810 1400.000 2430.880 ;
        RECT 1414.105 2430.810 1414.435 2430.825 ;
        RECT 1396.000 2430.510 1414.435 2430.810 ;
        RECT 1396.000 2430.280 1400.000 2430.510 ;
        RECT 1414.105 2430.495 1414.435 2430.510 ;
      LAYER met3 ;
        RECT 303.990 2421.080 1396.000 2429.880 ;
        RECT 304.400 2419.720 1396.000 2421.080 ;
        RECT 304.400 2419.680 1395.600 2419.720 ;
        RECT 303.990 2418.320 1395.600 2419.680 ;
      LAYER met3 ;
        RECT 1396.000 2419.250 1400.000 2419.320 ;
        RECT 1414.105 2419.250 1414.435 2419.265 ;
        RECT 1396.000 2418.950 1414.435 2419.250 ;
        RECT 1396.000 2418.720 1400.000 2418.950 ;
        RECT 1414.105 2418.935 1414.435 2418.950 ;
      LAYER met3 ;
        RECT 303.990 2410.880 1396.000 2418.320 ;
        RECT 304.400 2409.480 1396.000 2410.880 ;
        RECT 303.990 2408.840 1396.000 2409.480 ;
        RECT 303.990 2407.440 1395.600 2408.840 ;
      LAYER met3 ;
        RECT 1396.000 2408.370 1400.000 2408.440 ;
        RECT 1412.265 2408.370 1412.595 2408.385 ;
        RECT 1396.000 2408.070 1412.595 2408.370 ;
        RECT 1396.000 2407.840 1400.000 2408.070 ;
        RECT 1412.265 2408.055 1412.595 2408.070 ;
      LAYER met3 ;
        RECT 303.990 2400.680 1396.000 2407.440 ;
        RECT 304.400 2399.280 1396.000 2400.680 ;
        RECT 303.990 2397.960 1396.000 2399.280 ;
        RECT 303.990 2396.560 1395.600 2397.960 ;
      LAYER met3 ;
        RECT 1396.000 2397.490 1400.000 2397.560 ;
        RECT 1410.425 2397.490 1410.755 2397.505 ;
        RECT 1396.000 2397.190 1410.755 2397.490 ;
        RECT 1396.000 2396.960 1400.000 2397.190 ;
        RECT 1410.425 2397.175 1410.755 2397.190 ;
      LAYER met3 ;
        RECT 303.990 2389.800 1396.000 2396.560 ;
        RECT 304.400 2388.400 1396.000 2389.800 ;
        RECT 303.990 2387.080 1396.000 2388.400 ;
        RECT 303.990 2385.680 1395.600 2387.080 ;
      LAYER met3 ;
        RECT 1396.000 2386.610 1400.000 2386.680 ;
        RECT 1414.105 2386.610 1414.435 2386.625 ;
        RECT 1396.000 2386.310 1414.435 2386.610 ;
        RECT 1396.000 2386.080 1400.000 2386.310 ;
        RECT 1414.105 2386.295 1414.435 2386.310 ;
      LAYER met3 ;
        RECT 303.990 2379.600 1396.000 2385.680 ;
        RECT 304.400 2378.200 1396.000 2379.600 ;
        RECT 303.990 2376.200 1396.000 2378.200 ;
        RECT 303.990 2374.800 1395.600 2376.200 ;
      LAYER met3 ;
        RECT 1396.000 2375.730 1400.000 2375.800 ;
        RECT 1412.725 2375.730 1413.055 2375.745 ;
        RECT 1396.000 2375.430 1413.055 2375.730 ;
        RECT 1396.000 2375.200 1400.000 2375.430 ;
        RECT 1412.725 2375.415 1413.055 2375.430 ;
      LAYER met3 ;
        RECT 303.990 2368.720 1396.000 2374.800 ;
        RECT 304.400 2367.320 1396.000 2368.720 ;
        RECT 303.990 2365.320 1396.000 2367.320 ;
        RECT 303.990 2363.920 1395.600 2365.320 ;
      LAYER met3 ;
        RECT 1396.000 2364.850 1400.000 2364.920 ;
        RECT 1410.425 2364.850 1410.755 2364.865 ;
        RECT 1396.000 2364.550 1410.755 2364.850 ;
        RECT 1396.000 2364.320 1400.000 2364.550 ;
        RECT 1410.425 2364.535 1410.755 2364.550 ;
      LAYER met3 ;
        RECT 303.990 2358.520 1396.000 2363.920 ;
        RECT 304.400 2357.120 1396.000 2358.520 ;
        RECT 303.990 2353.760 1396.000 2357.120 ;
        RECT 303.990 2352.360 1395.600 2353.760 ;
      LAYER met3 ;
        RECT 1396.000 2353.290 1400.000 2353.360 ;
        RECT 1412.265 2353.290 1412.595 2353.305 ;
        RECT 1396.000 2352.990 1412.595 2353.290 ;
        RECT 1396.000 2352.760 1400.000 2352.990 ;
        RECT 1412.265 2352.975 1412.595 2352.990 ;
      LAYER met3 ;
        RECT 303.990 2347.640 1396.000 2352.360 ;
        RECT 304.400 2346.240 1396.000 2347.640 ;
        RECT 303.990 2342.880 1396.000 2346.240 ;
        RECT 303.990 2341.480 1395.600 2342.880 ;
      LAYER met3 ;
        RECT 1396.000 2342.410 1400.000 2342.480 ;
        RECT 1410.425 2342.410 1410.755 2342.425 ;
        RECT 1396.000 2342.110 1410.755 2342.410 ;
        RECT 1396.000 2341.880 1400.000 2342.110 ;
        RECT 1410.425 2342.095 1410.755 2342.110 ;
      LAYER met3 ;
        RECT 303.990 2337.440 1396.000 2341.480 ;
        RECT 304.400 2336.040 1396.000 2337.440 ;
        RECT 303.990 2332.000 1396.000 2336.040 ;
        RECT 303.990 2330.600 1395.600 2332.000 ;
      LAYER met3 ;
        RECT 1396.000 2331.530 1400.000 2331.600 ;
        RECT 1414.105 2331.530 1414.435 2331.545 ;
        RECT 1396.000 2331.230 1414.435 2331.530 ;
        RECT 1396.000 2331.000 1400.000 2331.230 ;
        RECT 1414.105 2331.215 1414.435 2331.230 ;
      LAYER met3 ;
        RECT 303.990 2326.560 1396.000 2330.600 ;
        RECT 304.400 2325.160 1396.000 2326.560 ;
        RECT 303.990 2321.120 1396.000 2325.160 ;
        RECT 303.990 2319.720 1395.600 2321.120 ;
      LAYER met3 ;
        RECT 1396.000 2320.650 1400.000 2320.720 ;
        RECT 1411.345 2320.650 1411.675 2320.665 ;
        RECT 1396.000 2320.350 1411.675 2320.650 ;
        RECT 1396.000 2320.120 1400.000 2320.350 ;
        RECT 1411.345 2320.335 1411.675 2320.350 ;
      LAYER met3 ;
        RECT 303.990 2316.360 1396.000 2319.720 ;
        RECT 304.400 2314.960 1396.000 2316.360 ;
        RECT 303.990 2310.240 1396.000 2314.960 ;
        RECT 303.990 2308.840 1395.600 2310.240 ;
      LAYER met3 ;
        RECT 1396.000 2309.770 1400.000 2309.840 ;
        RECT 1414.105 2309.770 1414.435 2309.785 ;
        RECT 1396.000 2309.470 1414.435 2309.770 ;
        RECT 1396.000 2309.240 1400.000 2309.470 ;
        RECT 1414.105 2309.455 1414.435 2309.470 ;
      LAYER met3 ;
        RECT 303.990 2305.480 1396.000 2308.840 ;
        RECT 304.400 2304.080 1396.000 2305.480 ;
        RECT 303.990 2298.680 1396.000 2304.080 ;
        RECT 303.990 2297.280 1395.600 2298.680 ;
      LAYER met3 ;
        RECT 1396.000 2298.210 1400.000 2298.280 ;
        RECT 1412.265 2298.210 1412.595 2298.225 ;
        RECT 1396.000 2297.910 1412.595 2298.210 ;
        RECT 1396.000 2297.680 1400.000 2297.910 ;
        RECT 1412.265 2297.895 1412.595 2297.910 ;
      LAYER met3 ;
        RECT 303.990 2295.280 1396.000 2297.280 ;
        RECT 304.400 2293.880 1396.000 2295.280 ;
        RECT 303.990 2287.800 1396.000 2293.880 ;
        RECT 303.990 2286.400 1395.600 2287.800 ;
      LAYER met3 ;
        RECT 1396.000 2287.330 1400.000 2287.400 ;
        RECT 1410.425 2287.330 1410.755 2287.345 ;
        RECT 1396.000 2287.030 1410.755 2287.330 ;
        RECT 1396.000 2286.800 1400.000 2287.030 ;
        RECT 1410.425 2287.015 1410.755 2287.030 ;
      LAYER met3 ;
        RECT 303.990 2284.400 1396.000 2286.400 ;
        RECT 304.400 2283.000 1396.000 2284.400 ;
        RECT 303.990 2276.920 1396.000 2283.000 ;
        RECT 303.990 2275.520 1395.600 2276.920 ;
      LAYER met3 ;
        RECT 1396.000 2276.450 1400.000 2276.520 ;
        RECT 1414.105 2276.450 1414.435 2276.465 ;
        RECT 1396.000 2276.150 1414.435 2276.450 ;
        RECT 1396.000 2275.920 1400.000 2276.150 ;
        RECT 1414.105 2276.135 1414.435 2276.150 ;
      LAYER met3 ;
        RECT 303.990 2274.200 1396.000 2275.520 ;
        RECT 304.400 2272.800 1396.000 2274.200 ;
        RECT 303.990 2266.040 1396.000 2272.800 ;
        RECT 303.990 2264.640 1395.600 2266.040 ;
      LAYER met3 ;
        RECT 1396.000 2265.570 1400.000 2265.640 ;
        RECT 1414.105 2265.570 1414.435 2265.585 ;
        RECT 1396.000 2265.270 1414.435 2265.570 ;
        RECT 1396.000 2265.040 1400.000 2265.270 ;
        RECT 1414.105 2265.255 1414.435 2265.270 ;
      LAYER met3 ;
        RECT 303.990 2263.320 1396.000 2264.640 ;
        RECT 304.400 2261.920 1396.000 2263.320 ;
        RECT 303.990 2255.160 1396.000 2261.920 ;
        RECT 303.990 2253.760 1395.600 2255.160 ;
      LAYER met3 ;
        RECT 1396.000 2254.690 1400.000 2254.760 ;
        RECT 1414.105 2254.690 1414.435 2254.705 ;
        RECT 1396.000 2254.390 1414.435 2254.690 ;
        RECT 1396.000 2254.160 1400.000 2254.390 ;
        RECT 1414.105 2254.375 1414.435 2254.390 ;
      LAYER met3 ;
        RECT 303.990 2253.120 1396.000 2253.760 ;
        RECT 304.400 2251.720 1396.000 2253.120 ;
        RECT 303.990 2243.600 1396.000 2251.720 ;
        RECT 303.990 2242.240 1395.600 2243.600 ;
      LAYER met3 ;
        RECT 1396.000 2243.130 1400.000 2243.200 ;
        RECT 1412.265 2243.130 1412.595 2243.145 ;
        RECT 1396.000 2242.830 1412.595 2243.130 ;
        RECT 1396.000 2242.600 1400.000 2242.830 ;
        RECT 1412.265 2242.815 1412.595 2242.830 ;
      LAYER met3 ;
        RECT 304.400 2242.200 1395.600 2242.240 ;
        RECT 304.400 2240.840 1396.000 2242.200 ;
        RECT 303.990 2232.720 1396.000 2240.840 ;
        RECT 303.990 2232.040 1395.600 2232.720 ;
        RECT 304.400 2231.320 1395.600 2232.040 ;
      LAYER met3 ;
        RECT 1396.000 2232.250 1400.000 2232.320 ;
        RECT 1414.105 2232.250 1414.435 2232.265 ;
        RECT 1396.000 2231.950 1414.435 2232.250 ;
        RECT 1396.000 2231.720 1400.000 2231.950 ;
        RECT 1414.105 2231.935 1414.435 2231.950 ;
      LAYER met3 ;
        RECT 304.400 2230.640 1396.000 2231.320 ;
        RECT 303.990 2221.840 1396.000 2230.640 ;
        RECT 303.990 2221.160 1395.600 2221.840 ;
        RECT 304.400 2220.440 1395.600 2221.160 ;
      LAYER met3 ;
        RECT 1396.000 2221.370 1400.000 2221.440 ;
        RECT 1414.105 2221.370 1414.435 2221.385 ;
        RECT 1396.000 2221.070 1414.435 2221.370 ;
        RECT 1396.000 2220.840 1400.000 2221.070 ;
        RECT 1414.105 2221.055 1414.435 2221.070 ;
      LAYER met3 ;
        RECT 304.400 2219.760 1396.000 2220.440 ;
        RECT 303.990 2210.960 1396.000 2219.760 ;
        RECT 304.400 2209.560 1395.600 2210.960 ;
      LAYER met3 ;
        RECT 1396.000 2210.490 1400.000 2210.560 ;
        RECT 1414.105 2210.490 1414.435 2210.505 ;
        RECT 1396.000 2210.190 1414.435 2210.490 ;
        RECT 1396.000 2209.960 1400.000 2210.190 ;
        RECT 1414.105 2210.175 1414.435 2210.190 ;
      LAYER met3 ;
        RECT 303.990 2200.080 1396.000 2209.560 ;
        RECT 304.400 2198.680 1395.600 2200.080 ;
      LAYER met3 ;
        RECT 1396.000 2199.610 1400.000 2199.680 ;
        RECT 1414.105 2199.610 1414.435 2199.625 ;
        RECT 1396.000 2199.310 1414.435 2199.610 ;
        RECT 1396.000 2199.080 1400.000 2199.310 ;
        RECT 1414.105 2199.295 1414.435 2199.310 ;
      LAYER met3 ;
        RECT 303.990 2189.880 1396.000 2198.680 ;
        RECT 304.400 2188.520 1396.000 2189.880 ;
        RECT 304.400 2188.480 1395.600 2188.520 ;
        RECT 303.990 2187.120 1395.600 2188.480 ;
      LAYER met3 ;
        RECT 1396.000 2188.050 1400.000 2188.120 ;
        RECT 1412.265 2188.050 1412.595 2188.065 ;
        RECT 1396.000 2187.750 1412.595 2188.050 ;
        RECT 1396.000 2187.520 1400.000 2187.750 ;
        RECT 1412.265 2187.735 1412.595 2187.750 ;
      LAYER met3 ;
        RECT 303.990 2179.000 1396.000 2187.120 ;
        RECT 304.400 2177.640 1396.000 2179.000 ;
        RECT 304.400 2177.600 1395.600 2177.640 ;
        RECT 303.990 2176.240 1395.600 2177.600 ;
      LAYER met3 ;
        RECT 1396.000 2177.170 1400.000 2177.240 ;
        RECT 1414.105 2177.170 1414.435 2177.185 ;
        RECT 1396.000 2176.870 1414.435 2177.170 ;
        RECT 1396.000 2176.640 1400.000 2176.870 ;
        RECT 1414.105 2176.855 1414.435 2176.870 ;
      LAYER met3 ;
        RECT 303.990 2168.800 1396.000 2176.240 ;
        RECT 304.400 2167.400 1396.000 2168.800 ;
        RECT 303.990 2166.760 1396.000 2167.400 ;
        RECT 303.990 2165.360 1395.600 2166.760 ;
      LAYER met3 ;
        RECT 1396.000 2166.290 1400.000 2166.360 ;
        RECT 1414.105 2166.290 1414.435 2166.305 ;
        RECT 1396.000 2165.990 1414.435 2166.290 ;
        RECT 1396.000 2165.760 1400.000 2165.990 ;
        RECT 1414.105 2165.975 1414.435 2165.990 ;
      LAYER met3 ;
        RECT 303.990 2157.920 1396.000 2165.360 ;
        RECT 304.400 2156.520 1396.000 2157.920 ;
        RECT 303.990 2155.880 1396.000 2156.520 ;
        RECT 303.990 2154.480 1395.600 2155.880 ;
      LAYER met3 ;
        RECT 1396.000 2155.410 1400.000 2155.480 ;
        RECT 1414.105 2155.410 1414.435 2155.425 ;
        RECT 1396.000 2155.110 1414.435 2155.410 ;
        RECT 1396.000 2154.880 1400.000 2155.110 ;
        RECT 1414.105 2155.095 1414.435 2155.110 ;
      LAYER met3 ;
        RECT 303.990 2147.720 1396.000 2154.480 ;
        RECT 304.400 2146.320 1396.000 2147.720 ;
        RECT 303.990 2145.000 1396.000 2146.320 ;
        RECT 303.990 2143.600 1395.600 2145.000 ;
      LAYER met3 ;
        RECT 1396.000 2144.530 1400.000 2144.600 ;
        RECT 1414.105 2144.530 1414.435 2144.545 ;
        RECT 1396.000 2144.230 1414.435 2144.530 ;
        RECT 1396.000 2144.000 1400.000 2144.230 ;
        RECT 1414.105 2144.215 1414.435 2144.230 ;
      LAYER met3 ;
        RECT 303.990 2136.840 1396.000 2143.600 ;
        RECT 304.400 2135.440 1396.000 2136.840 ;
        RECT 303.990 2133.440 1396.000 2135.440 ;
        RECT 303.990 2132.040 1395.600 2133.440 ;
      LAYER met3 ;
        RECT 1396.000 2132.970 1400.000 2133.040 ;
        RECT 1414.105 2132.970 1414.435 2132.985 ;
        RECT 1396.000 2132.670 1414.435 2132.970 ;
        RECT 1396.000 2132.440 1400.000 2132.670 ;
        RECT 1414.105 2132.655 1414.435 2132.670 ;
      LAYER met3 ;
        RECT 303.990 2126.640 1396.000 2132.040 ;
        RECT 304.400 2125.240 1396.000 2126.640 ;
        RECT 303.990 2122.560 1396.000 2125.240 ;
        RECT 303.990 2121.160 1395.600 2122.560 ;
      LAYER met3 ;
        RECT 1396.000 2122.090 1400.000 2122.160 ;
        RECT 1412.265 2122.090 1412.595 2122.105 ;
        RECT 1396.000 2121.790 1412.595 2122.090 ;
        RECT 1396.000 2121.560 1400.000 2121.790 ;
        RECT 1412.265 2121.775 1412.595 2121.790 ;
      LAYER met3 ;
        RECT 303.990 2115.760 1396.000 2121.160 ;
        RECT 304.400 2114.360 1396.000 2115.760 ;
        RECT 303.990 2111.680 1396.000 2114.360 ;
        RECT 303.990 2110.280 1395.600 2111.680 ;
      LAYER met3 ;
        RECT 1396.000 2111.210 1400.000 2111.280 ;
        RECT 1410.425 2111.210 1410.755 2111.225 ;
        RECT 1396.000 2110.910 1410.755 2111.210 ;
        RECT 1396.000 2110.680 1400.000 2110.910 ;
        RECT 1410.425 2110.895 1410.755 2110.910 ;
      LAYER met3 ;
        RECT 303.990 2105.560 1396.000 2110.280 ;
        RECT 304.400 2104.160 1396.000 2105.560 ;
        RECT 303.990 2100.800 1396.000 2104.160 ;
        RECT 303.990 2099.400 1395.600 2100.800 ;
      LAYER met3 ;
        RECT 1396.000 2100.330 1400.000 2100.400 ;
        RECT 1408.585 2100.330 1408.915 2100.345 ;
        RECT 1396.000 2100.030 1408.915 2100.330 ;
        RECT 1396.000 2099.800 1400.000 2100.030 ;
        RECT 1408.585 2100.015 1408.915 2100.030 ;
      LAYER met3 ;
        RECT 303.990 2095.360 1396.000 2099.400 ;
        RECT 304.400 2093.960 1396.000 2095.360 ;
        RECT 303.990 2089.920 1396.000 2093.960 ;
        RECT 303.990 2088.520 1395.600 2089.920 ;
      LAYER met3 ;
        RECT 1396.000 2089.450 1400.000 2089.520 ;
        RECT 1414.105 2089.450 1414.435 2089.465 ;
        RECT 1396.000 2089.150 1414.435 2089.450 ;
        RECT 1396.000 2088.920 1400.000 2089.150 ;
        RECT 1414.105 2089.135 1414.435 2089.150 ;
      LAYER met3 ;
        RECT 303.990 2084.480 1396.000 2088.520 ;
        RECT 304.400 2083.080 1396.000 2084.480 ;
        RECT 303.990 2079.040 1396.000 2083.080 ;
        RECT 303.990 2077.640 1395.600 2079.040 ;
      LAYER met3 ;
        RECT 1396.000 2078.570 1400.000 2078.640 ;
        RECT 1414.105 2078.570 1414.435 2078.585 ;
        RECT 1396.000 2078.270 1414.435 2078.570 ;
        RECT 1396.000 2078.040 1400.000 2078.270 ;
        RECT 1414.105 2078.255 1414.435 2078.270 ;
      LAYER met3 ;
        RECT 303.990 2074.280 1396.000 2077.640 ;
        RECT 304.400 2072.880 1396.000 2074.280 ;
        RECT 303.990 2067.480 1396.000 2072.880 ;
        RECT 303.990 2066.080 1395.600 2067.480 ;
      LAYER met3 ;
        RECT 1396.000 2067.010 1400.000 2067.080 ;
        RECT 1409.505 2067.010 1409.835 2067.025 ;
        RECT 1396.000 2066.710 1409.835 2067.010 ;
        RECT 1396.000 2066.480 1400.000 2066.710 ;
        RECT 1409.505 2066.695 1409.835 2066.710 ;
      LAYER met3 ;
        RECT 303.990 2063.400 1396.000 2066.080 ;
        RECT 304.400 2062.000 1396.000 2063.400 ;
        RECT 303.990 2056.600 1396.000 2062.000 ;
        RECT 303.990 2055.200 1395.600 2056.600 ;
      LAYER met3 ;
        RECT 1396.000 2056.130 1400.000 2056.200 ;
        RECT 1414.105 2056.130 1414.435 2056.145 ;
        RECT 1396.000 2055.830 1414.435 2056.130 ;
        RECT 1396.000 2055.600 1400.000 2055.830 ;
        RECT 1414.105 2055.815 1414.435 2055.830 ;
      LAYER met3 ;
        RECT 303.990 2053.200 1396.000 2055.200 ;
        RECT 304.400 2051.800 1396.000 2053.200 ;
        RECT 303.990 2045.720 1396.000 2051.800 ;
        RECT 303.990 2044.320 1395.600 2045.720 ;
      LAYER met3 ;
        RECT 1396.000 2045.250 1400.000 2045.320 ;
        RECT 1410.425 2045.250 1410.755 2045.265 ;
        RECT 1396.000 2044.950 1410.755 2045.250 ;
        RECT 1396.000 2044.720 1400.000 2044.950 ;
        RECT 1410.425 2044.935 1410.755 2044.950 ;
      LAYER met3 ;
        RECT 303.990 2042.320 1396.000 2044.320 ;
        RECT 304.400 2040.920 1396.000 2042.320 ;
        RECT 303.990 2034.840 1396.000 2040.920 ;
        RECT 303.990 2033.440 1395.600 2034.840 ;
      LAYER met3 ;
        RECT 1396.000 2034.370 1400.000 2034.440 ;
        RECT 1414.105 2034.370 1414.435 2034.385 ;
        RECT 1396.000 2034.070 1414.435 2034.370 ;
        RECT 1396.000 2033.840 1400.000 2034.070 ;
        RECT 1414.105 2034.055 1414.435 2034.070 ;
      LAYER met3 ;
        RECT 303.990 2032.120 1396.000 2033.440 ;
        RECT 304.400 2030.720 1396.000 2032.120 ;
        RECT 303.990 2023.960 1396.000 2030.720 ;
        RECT 303.990 2022.560 1395.600 2023.960 ;
      LAYER met3 ;
        RECT 1396.000 2023.490 1400.000 2023.560 ;
        RECT 1414.105 2023.490 1414.435 2023.505 ;
        RECT 1396.000 2023.190 1414.435 2023.490 ;
        RECT 1396.000 2022.960 1400.000 2023.190 ;
        RECT 1414.105 2023.175 1414.435 2023.190 ;
      LAYER met3 ;
        RECT 303.990 2021.240 1396.000 2022.560 ;
        RECT 304.400 2019.840 1396.000 2021.240 ;
        RECT 303.990 2012.400 1396.000 2019.840 ;
        RECT 303.990 2011.040 1395.600 2012.400 ;
      LAYER met3 ;
        RECT 1396.000 2011.930 1400.000 2012.000 ;
        RECT 1409.505 2011.930 1409.835 2011.945 ;
        RECT 1396.000 2011.630 1409.835 2011.930 ;
        RECT 1396.000 2011.400 1400.000 2011.630 ;
        RECT 1409.505 2011.615 1409.835 2011.630 ;
      LAYER met3 ;
        RECT 304.400 2011.000 1395.600 2011.040 ;
        RECT 304.400 2009.640 1396.000 2011.000 ;
        RECT 303.990 2001.520 1396.000 2009.640 ;
        RECT 303.990 2000.160 1395.600 2001.520 ;
      LAYER met3 ;
        RECT 1396.000 2001.050 1400.000 2001.120 ;
        RECT 1414.105 2001.050 1414.435 2001.065 ;
        RECT 1396.000 2000.750 1414.435 2001.050 ;
        RECT 1396.000 2000.520 1400.000 2000.750 ;
        RECT 1414.105 2000.735 1414.435 2000.750 ;
      LAYER met3 ;
        RECT 304.400 2000.120 1395.600 2000.160 ;
        RECT 304.400 1998.760 1396.000 2000.120 ;
        RECT 303.990 1990.640 1396.000 1998.760 ;
        RECT 303.990 1989.960 1395.600 1990.640 ;
        RECT 304.400 1989.240 1395.600 1989.960 ;
      LAYER met3 ;
        RECT 1396.000 1990.170 1400.000 1990.240 ;
        RECT 1410.425 1990.170 1410.755 1990.185 ;
        RECT 1396.000 1989.870 1410.755 1990.170 ;
        RECT 1396.000 1989.640 1400.000 1989.870 ;
        RECT 1410.425 1989.855 1410.755 1989.870 ;
      LAYER met3 ;
        RECT 304.400 1988.560 1396.000 1989.240 ;
        RECT 303.990 1979.760 1396.000 1988.560 ;
        RECT 303.990 1979.080 1395.600 1979.760 ;
        RECT 304.400 1978.360 1395.600 1979.080 ;
      LAYER met3 ;
        RECT 1396.000 1979.290 1400.000 1979.360 ;
        RECT 1410.425 1979.290 1410.755 1979.305 ;
        RECT 1396.000 1978.990 1410.755 1979.290 ;
        RECT 1396.000 1978.760 1400.000 1978.990 ;
        RECT 1410.425 1978.975 1410.755 1978.990 ;
      LAYER met3 ;
        RECT 304.400 1977.680 1396.000 1978.360 ;
        RECT 303.990 1968.880 1396.000 1977.680 ;
        RECT 304.400 1967.480 1395.600 1968.880 ;
      LAYER met3 ;
        RECT 1396.000 1968.410 1400.000 1968.480 ;
        RECT 1411.345 1968.410 1411.675 1968.425 ;
        RECT 1396.000 1968.110 1411.675 1968.410 ;
        RECT 1396.000 1967.880 1400.000 1968.110 ;
        RECT 1411.345 1968.095 1411.675 1968.110 ;
      LAYER met3 ;
        RECT 303.990 1958.000 1396.000 1967.480 ;
        RECT 304.400 1957.320 1396.000 1958.000 ;
        RECT 304.400 1956.600 1395.600 1957.320 ;
        RECT 303.990 1955.920 1395.600 1956.600 ;
      LAYER met3 ;
        RECT 1396.000 1956.850 1400.000 1956.920 ;
        RECT 1409.505 1956.850 1409.835 1956.865 ;
        RECT 1396.000 1956.550 1409.835 1956.850 ;
        RECT 1396.000 1956.320 1400.000 1956.550 ;
        RECT 1409.505 1956.535 1409.835 1956.550 ;
      LAYER met3 ;
        RECT 303.990 1947.800 1396.000 1955.920 ;
        RECT 304.400 1946.440 1396.000 1947.800 ;
        RECT 304.400 1946.400 1395.600 1946.440 ;
        RECT 303.990 1945.040 1395.600 1946.400 ;
      LAYER met3 ;
        RECT 1396.000 1945.970 1400.000 1946.040 ;
        RECT 1412.265 1945.970 1412.595 1945.985 ;
        RECT 1396.000 1945.670 1412.595 1945.970 ;
        RECT 1396.000 1945.440 1400.000 1945.670 ;
        RECT 1412.265 1945.655 1412.595 1945.670 ;
      LAYER met3 ;
        RECT 303.990 1936.920 1396.000 1945.040 ;
        RECT 304.400 1935.560 1396.000 1936.920 ;
        RECT 304.400 1935.520 1395.600 1935.560 ;
        RECT 303.990 1934.160 1395.600 1935.520 ;
      LAYER met3 ;
        RECT 1396.000 1935.090 1400.000 1935.160 ;
        RECT 1410.425 1935.090 1410.755 1935.105 ;
        RECT 1396.000 1934.790 1410.755 1935.090 ;
        RECT 1396.000 1934.560 1400.000 1934.790 ;
        RECT 1410.425 1934.775 1410.755 1934.790 ;
      LAYER met3 ;
        RECT 303.990 1926.720 1396.000 1934.160 ;
        RECT 304.400 1925.320 1396.000 1926.720 ;
        RECT 303.990 1924.680 1396.000 1925.320 ;
        RECT 303.990 1923.280 1395.600 1924.680 ;
      LAYER met3 ;
        RECT 1396.000 1924.210 1400.000 1924.280 ;
        RECT 1414.105 1924.210 1414.435 1924.225 ;
        RECT 1396.000 1923.910 1414.435 1924.210 ;
        RECT 1396.000 1923.680 1400.000 1923.910 ;
        RECT 1414.105 1923.895 1414.435 1923.910 ;
      LAYER met3 ;
        RECT 303.990 1915.840 1396.000 1923.280 ;
        RECT 304.400 1914.440 1396.000 1915.840 ;
        RECT 303.990 1913.800 1396.000 1914.440 ;
        RECT 303.990 1912.400 1395.600 1913.800 ;
      LAYER met3 ;
        RECT 1396.000 1913.330 1400.000 1913.400 ;
        RECT 1414.105 1913.330 1414.435 1913.345 ;
        RECT 1396.000 1913.030 1414.435 1913.330 ;
        RECT 1396.000 1912.800 1400.000 1913.030 ;
        RECT 1414.105 1913.015 1414.435 1913.030 ;
      LAYER met3 ;
        RECT 303.990 1905.640 1396.000 1912.400 ;
        RECT 304.400 1904.240 1396.000 1905.640 ;
        RECT 303.990 1902.240 1396.000 1904.240 ;
        RECT 303.990 1900.840 1395.600 1902.240 ;
      LAYER met3 ;
        RECT 1396.000 1901.770 1400.000 1901.840 ;
        RECT 1414.105 1901.770 1414.435 1901.785 ;
        RECT 1396.000 1901.470 1414.435 1901.770 ;
        RECT 1396.000 1901.240 1400.000 1901.470 ;
        RECT 1414.105 1901.455 1414.435 1901.470 ;
      LAYER met3 ;
        RECT 303.990 1894.760 1396.000 1900.840 ;
        RECT 304.400 1893.360 1396.000 1894.760 ;
        RECT 303.990 1891.360 1396.000 1893.360 ;
        RECT 303.990 1889.960 1395.600 1891.360 ;
      LAYER met3 ;
        RECT 1396.000 1890.890 1400.000 1890.960 ;
        RECT 1412.265 1890.890 1412.595 1890.905 ;
        RECT 1396.000 1890.590 1412.595 1890.890 ;
        RECT 1396.000 1890.360 1400.000 1890.590 ;
        RECT 1412.265 1890.575 1412.595 1890.590 ;
      LAYER met3 ;
        RECT 303.990 1884.560 1396.000 1889.960 ;
        RECT 304.400 1883.160 1396.000 1884.560 ;
        RECT 303.990 1880.480 1396.000 1883.160 ;
        RECT 303.990 1879.080 1395.600 1880.480 ;
      LAYER met3 ;
        RECT 1396.000 1880.010 1400.000 1880.080 ;
        RECT 1410.425 1880.010 1410.755 1880.025 ;
        RECT 1396.000 1879.710 1410.755 1880.010 ;
        RECT 1396.000 1879.480 1400.000 1879.710 ;
        RECT 1410.425 1879.695 1410.755 1879.710 ;
      LAYER met3 ;
        RECT 303.990 1873.680 1396.000 1879.080 ;
        RECT 304.400 1872.280 1396.000 1873.680 ;
        RECT 303.990 1869.600 1396.000 1872.280 ;
        RECT 303.990 1868.200 1395.600 1869.600 ;
      LAYER met3 ;
        RECT 1396.000 1869.130 1400.000 1869.200 ;
        RECT 1414.105 1869.130 1414.435 1869.145 ;
        RECT 1396.000 1868.830 1414.435 1869.130 ;
        RECT 1396.000 1868.600 1400.000 1868.830 ;
        RECT 1414.105 1868.815 1414.435 1868.830 ;
      LAYER met3 ;
        RECT 303.990 1863.480 1396.000 1868.200 ;
        RECT 304.400 1862.080 1396.000 1863.480 ;
        RECT 303.990 1858.720 1396.000 1862.080 ;
        RECT 303.990 1857.320 1395.600 1858.720 ;
      LAYER met3 ;
        RECT 1396.000 1858.250 1400.000 1858.320 ;
        RECT 1412.725 1858.250 1413.055 1858.265 ;
        RECT 1396.000 1857.950 1413.055 1858.250 ;
        RECT 1396.000 1857.720 1400.000 1857.950 ;
        RECT 1412.725 1857.935 1413.055 1857.950 ;
      LAYER met3 ;
        RECT 303.990 1852.600 1396.000 1857.320 ;
        RECT 304.400 1851.200 1396.000 1852.600 ;
        RECT 303.990 1847.160 1396.000 1851.200 ;
        RECT 303.990 1845.760 1395.600 1847.160 ;
      LAYER met3 ;
        RECT 1396.000 1846.690 1400.000 1846.760 ;
        RECT 1414.105 1846.690 1414.435 1846.705 ;
        RECT 1396.000 1846.390 1414.435 1846.690 ;
        RECT 1396.000 1846.160 1400.000 1846.390 ;
        RECT 1414.105 1846.375 1414.435 1846.390 ;
      LAYER met3 ;
        RECT 303.990 1842.400 1396.000 1845.760 ;
        RECT 304.400 1841.000 1396.000 1842.400 ;
        RECT 303.990 1836.280 1396.000 1841.000 ;
        RECT 303.990 1834.880 1395.600 1836.280 ;
      LAYER met3 ;
        RECT 1396.000 1835.810 1400.000 1835.880 ;
        RECT 1412.265 1835.810 1412.595 1835.825 ;
        RECT 1396.000 1835.510 1412.595 1835.810 ;
        RECT 1396.000 1835.280 1400.000 1835.510 ;
        RECT 1412.265 1835.495 1412.595 1835.510 ;
      LAYER met3 ;
        RECT 303.990 1831.520 1396.000 1834.880 ;
        RECT 304.400 1830.120 1396.000 1831.520 ;
        RECT 303.990 1825.400 1396.000 1830.120 ;
        RECT 303.990 1824.000 1395.600 1825.400 ;
      LAYER met3 ;
        RECT 1396.000 1824.930 1400.000 1825.000 ;
        RECT 1410.425 1824.930 1410.755 1824.945 ;
        RECT 1396.000 1824.630 1410.755 1824.930 ;
        RECT 1396.000 1824.400 1400.000 1824.630 ;
        RECT 1410.425 1824.615 1410.755 1824.630 ;
      LAYER met3 ;
        RECT 303.990 1821.320 1396.000 1824.000 ;
        RECT 304.400 1819.920 1396.000 1821.320 ;
        RECT 303.990 1814.520 1396.000 1819.920 ;
        RECT 303.990 1813.120 1395.600 1814.520 ;
      LAYER met3 ;
        RECT 1396.000 1814.050 1400.000 1814.120 ;
        RECT 1414.105 1814.050 1414.435 1814.065 ;
        RECT 1396.000 1813.750 1414.435 1814.050 ;
        RECT 1396.000 1813.520 1400.000 1813.750 ;
        RECT 1414.105 1813.735 1414.435 1813.750 ;
      LAYER met3 ;
        RECT 303.990 1810.440 1396.000 1813.120 ;
        RECT 304.400 1809.040 1396.000 1810.440 ;
        RECT 303.990 1803.640 1396.000 1809.040 ;
        RECT 303.990 1802.240 1395.600 1803.640 ;
      LAYER met3 ;
        RECT 1396.000 1803.170 1400.000 1803.240 ;
        RECT 1412.725 1803.170 1413.055 1803.185 ;
        RECT 1396.000 1802.870 1413.055 1803.170 ;
        RECT 1396.000 1802.640 1400.000 1802.870 ;
        RECT 1412.725 1802.855 1413.055 1802.870 ;
      LAYER met3 ;
        RECT 303.990 1800.240 1396.000 1802.240 ;
        RECT 304.400 1798.840 1396.000 1800.240 ;
        RECT 303.990 1792.760 1396.000 1798.840 ;
        RECT 303.990 1791.360 1395.600 1792.760 ;
      LAYER met3 ;
        RECT 1396.000 1792.290 1400.000 1792.360 ;
        RECT 1414.105 1792.290 1414.435 1792.305 ;
        RECT 1396.000 1791.990 1414.435 1792.290 ;
        RECT 1396.000 1791.760 1400.000 1791.990 ;
        RECT 1414.105 1791.975 1414.435 1791.990 ;
      LAYER met3 ;
        RECT 303.990 1790.040 1396.000 1791.360 ;
        RECT 304.400 1788.640 1396.000 1790.040 ;
        RECT 303.990 1781.200 1396.000 1788.640 ;
        RECT 303.990 1779.800 1395.600 1781.200 ;
      LAYER met3 ;
        RECT 1396.000 1780.730 1400.000 1780.800 ;
        RECT 1412.265 1780.730 1412.595 1780.745 ;
        RECT 1396.000 1780.430 1412.595 1780.730 ;
        RECT 1396.000 1780.200 1400.000 1780.430 ;
        RECT 1412.265 1780.415 1412.595 1780.430 ;
      LAYER met3 ;
        RECT 303.990 1779.160 1396.000 1779.800 ;
        RECT 304.400 1777.760 1396.000 1779.160 ;
        RECT 303.990 1770.320 1396.000 1777.760 ;
        RECT 303.990 1768.960 1395.600 1770.320 ;
      LAYER met3 ;
        RECT 1396.000 1769.850 1400.000 1769.920 ;
        RECT 1410.425 1769.850 1410.755 1769.865 ;
        RECT 1396.000 1769.550 1410.755 1769.850 ;
        RECT 1396.000 1769.320 1400.000 1769.550 ;
        RECT 1410.425 1769.535 1410.755 1769.550 ;
      LAYER met3 ;
        RECT 304.400 1768.920 1395.600 1768.960 ;
        RECT 304.400 1767.560 1396.000 1768.920 ;
        RECT 303.990 1759.440 1396.000 1767.560 ;
        RECT 303.990 1758.080 1395.600 1759.440 ;
      LAYER met3 ;
        RECT 1396.000 1758.970 1400.000 1759.040 ;
        RECT 1414.105 1758.970 1414.435 1758.985 ;
        RECT 1396.000 1758.670 1414.435 1758.970 ;
        RECT 1396.000 1758.440 1400.000 1758.670 ;
        RECT 1414.105 1758.655 1414.435 1758.670 ;
      LAYER met3 ;
        RECT 304.400 1758.040 1395.600 1758.080 ;
        RECT 304.400 1756.680 1396.000 1758.040 ;
        RECT 303.990 1748.560 1396.000 1756.680 ;
        RECT 303.990 1747.880 1395.600 1748.560 ;
        RECT 304.400 1747.160 1395.600 1747.880 ;
      LAYER met3 ;
        RECT 1396.000 1748.090 1400.000 1748.160 ;
        RECT 1412.725 1748.090 1413.055 1748.105 ;
        RECT 1396.000 1747.790 1413.055 1748.090 ;
        RECT 1396.000 1747.560 1400.000 1747.790 ;
        RECT 1412.725 1747.775 1413.055 1747.790 ;
      LAYER met3 ;
        RECT 304.400 1746.480 1396.000 1747.160 ;
        RECT 303.990 1737.680 1396.000 1746.480 ;
        RECT 303.990 1737.000 1395.600 1737.680 ;
        RECT 304.400 1736.280 1395.600 1737.000 ;
      LAYER met3 ;
        RECT 1396.000 1737.210 1400.000 1737.280 ;
        RECT 1414.105 1737.210 1414.435 1737.225 ;
        RECT 1396.000 1736.910 1414.435 1737.210 ;
        RECT 1396.000 1736.680 1400.000 1736.910 ;
        RECT 1414.105 1736.895 1414.435 1736.910 ;
      LAYER met3 ;
        RECT 304.400 1735.600 1396.000 1736.280 ;
        RECT 303.990 1726.800 1396.000 1735.600 ;
        RECT 304.400 1726.120 1396.000 1726.800 ;
        RECT 304.400 1725.400 1395.600 1726.120 ;
        RECT 303.990 1724.720 1395.600 1725.400 ;
      LAYER met3 ;
        RECT 1396.000 1725.650 1400.000 1725.720 ;
        RECT 1412.265 1725.650 1412.595 1725.665 ;
        RECT 1396.000 1725.350 1412.595 1725.650 ;
        RECT 1396.000 1725.120 1400.000 1725.350 ;
        RECT 1412.265 1725.335 1412.595 1725.350 ;
      LAYER met3 ;
        RECT 303.990 1715.920 1396.000 1724.720 ;
        RECT 304.400 1715.240 1396.000 1715.920 ;
        RECT 304.400 1714.520 1395.600 1715.240 ;
        RECT 303.990 1713.840 1395.600 1714.520 ;
      LAYER met3 ;
        RECT 1396.000 1714.770 1400.000 1714.840 ;
        RECT 1414.105 1714.770 1414.435 1714.785 ;
        RECT 1396.000 1714.470 1414.435 1714.770 ;
        RECT 1396.000 1714.240 1400.000 1714.470 ;
        RECT 1414.105 1714.455 1414.435 1714.470 ;
      LAYER met3 ;
        RECT 303.990 1705.720 1396.000 1713.840 ;
        RECT 304.400 1704.360 1396.000 1705.720 ;
        RECT 304.400 1704.320 1395.600 1704.360 ;
        RECT 303.990 1702.960 1395.600 1704.320 ;
      LAYER met3 ;
        RECT 1396.000 1703.890 1400.000 1703.960 ;
        RECT 1414.105 1703.890 1414.435 1703.905 ;
        RECT 1396.000 1703.590 1414.435 1703.890 ;
        RECT 1396.000 1703.360 1400.000 1703.590 ;
        RECT 1414.105 1703.575 1414.435 1703.590 ;
      LAYER met3 ;
        RECT 303.990 1694.840 1396.000 1702.960 ;
        RECT 304.400 1693.480 1396.000 1694.840 ;
        RECT 304.400 1693.440 1395.600 1693.480 ;
        RECT 303.990 1692.080 1395.600 1693.440 ;
      LAYER met3 ;
        RECT 1396.000 1693.010 1400.000 1693.080 ;
        RECT 1414.105 1693.010 1414.435 1693.025 ;
        RECT 1396.000 1692.710 1414.435 1693.010 ;
        RECT 1396.000 1692.480 1400.000 1692.710 ;
        RECT 1414.105 1692.695 1414.435 1692.710 ;
      LAYER met3 ;
        RECT 303.990 1684.640 1396.000 1692.080 ;
        RECT 304.400 1683.240 1396.000 1684.640 ;
        RECT 303.990 1682.600 1396.000 1683.240 ;
        RECT 303.990 1681.200 1395.600 1682.600 ;
      LAYER met3 ;
        RECT 1396.000 1682.130 1400.000 1682.200 ;
        RECT 1414.105 1682.130 1414.435 1682.145 ;
        RECT 1396.000 1681.830 1414.435 1682.130 ;
        RECT 1396.000 1681.600 1400.000 1681.830 ;
        RECT 1414.105 1681.815 1414.435 1681.830 ;
      LAYER met3 ;
        RECT 303.990 1673.760 1396.000 1681.200 ;
        RECT 304.400 1672.360 1396.000 1673.760 ;
        RECT 303.990 1671.040 1396.000 1672.360 ;
        RECT 303.990 1669.640 1395.600 1671.040 ;
      LAYER met3 ;
        RECT 1396.000 1670.570 1400.000 1670.640 ;
        RECT 1411.805 1670.570 1412.135 1670.585 ;
        RECT 1396.000 1670.270 1412.135 1670.570 ;
        RECT 1396.000 1670.040 1400.000 1670.270 ;
        RECT 1411.805 1670.255 1412.135 1670.270 ;
      LAYER met3 ;
        RECT 303.990 1663.560 1396.000 1669.640 ;
        RECT 304.400 1662.160 1396.000 1663.560 ;
        RECT 303.990 1660.160 1396.000 1662.160 ;
        RECT 303.990 1658.760 1395.600 1660.160 ;
      LAYER met3 ;
        RECT 1396.000 1659.690 1400.000 1659.760 ;
        RECT 1414.105 1659.690 1414.435 1659.705 ;
        RECT 1396.000 1659.390 1414.435 1659.690 ;
        RECT 1396.000 1659.160 1400.000 1659.390 ;
        RECT 1414.105 1659.375 1414.435 1659.390 ;
      LAYER met3 ;
        RECT 303.990 1652.680 1396.000 1658.760 ;
        RECT 304.400 1651.280 1396.000 1652.680 ;
        RECT 303.990 1649.280 1396.000 1651.280 ;
        RECT 303.990 1647.880 1395.600 1649.280 ;
      LAYER met3 ;
        RECT 1396.000 1648.810 1400.000 1648.880 ;
        RECT 1414.105 1648.810 1414.435 1648.825 ;
        RECT 1396.000 1648.510 1414.435 1648.810 ;
        RECT 1396.000 1648.280 1400.000 1648.510 ;
        RECT 1414.105 1648.495 1414.435 1648.510 ;
      LAYER met3 ;
        RECT 303.990 1642.480 1396.000 1647.880 ;
        RECT 304.400 1641.080 1396.000 1642.480 ;
        RECT 303.990 1638.400 1396.000 1641.080 ;
        RECT 303.990 1637.000 1395.600 1638.400 ;
      LAYER met3 ;
        RECT 1396.000 1637.930 1400.000 1638.000 ;
        RECT 1414.105 1637.930 1414.435 1637.945 ;
        RECT 1396.000 1637.630 1414.435 1637.930 ;
        RECT 1396.000 1637.400 1400.000 1637.630 ;
        RECT 1414.105 1637.615 1414.435 1637.630 ;
      LAYER met3 ;
        RECT 303.990 1631.600 1396.000 1637.000 ;
        RECT 304.400 1630.200 1396.000 1631.600 ;
        RECT 303.990 1627.520 1396.000 1630.200 ;
        RECT 303.990 1626.120 1395.600 1627.520 ;
      LAYER met3 ;
        RECT 1396.000 1627.050 1400.000 1627.120 ;
        RECT 1414.105 1627.050 1414.435 1627.065 ;
        RECT 1396.000 1626.750 1414.435 1627.050 ;
        RECT 1396.000 1626.520 1400.000 1626.750 ;
        RECT 1414.105 1626.735 1414.435 1626.750 ;
      LAYER met3 ;
        RECT 303.990 1621.400 1396.000 1626.120 ;
        RECT 304.400 1620.000 1396.000 1621.400 ;
        RECT 303.990 1615.960 1396.000 1620.000 ;
        RECT 303.990 1614.560 1395.600 1615.960 ;
      LAYER met3 ;
        RECT 1396.000 1615.490 1400.000 1615.560 ;
        RECT 1411.805 1615.490 1412.135 1615.505 ;
        RECT 1396.000 1615.190 1412.135 1615.490 ;
        RECT 1396.000 1614.960 1400.000 1615.190 ;
        RECT 1411.805 1615.175 1412.135 1615.190 ;
      LAYER met3 ;
        RECT 303.990 1610.520 1396.000 1614.560 ;
        RECT 304.400 1609.120 1396.000 1610.520 ;
        RECT 303.990 1605.080 1396.000 1609.120 ;
        RECT 303.990 1603.680 1395.600 1605.080 ;
      LAYER met3 ;
        RECT 1396.000 1604.610 1400.000 1604.680 ;
        RECT 1414.105 1604.610 1414.435 1604.625 ;
        RECT 1396.000 1604.310 1414.435 1604.610 ;
        RECT 1396.000 1604.080 1400.000 1604.310 ;
        RECT 1414.105 1604.295 1414.435 1604.310 ;
      LAYER met3 ;
        RECT 303.990 1600.320 1396.000 1603.680 ;
        RECT 304.400 1598.920 1396.000 1600.320 ;
        RECT 303.990 1594.200 1396.000 1598.920 ;
        RECT 303.990 1592.800 1395.600 1594.200 ;
      LAYER met3 ;
        RECT 1396.000 1593.730 1400.000 1593.800 ;
        RECT 1414.105 1593.730 1414.435 1593.745 ;
        RECT 1396.000 1593.430 1414.435 1593.730 ;
        RECT 1396.000 1593.200 1400.000 1593.430 ;
        RECT 1414.105 1593.415 1414.435 1593.430 ;
      LAYER met3 ;
        RECT 303.990 1589.440 1396.000 1592.800 ;
        RECT 304.400 1588.040 1396.000 1589.440 ;
        RECT 303.990 1583.320 1396.000 1588.040 ;
        RECT 303.990 1581.920 1395.600 1583.320 ;
      LAYER met3 ;
        RECT 1396.000 1582.850 1400.000 1582.920 ;
        RECT 1414.105 1582.850 1414.435 1582.865 ;
        RECT 1396.000 1582.550 1414.435 1582.850 ;
        RECT 1396.000 1582.320 1400.000 1582.550 ;
        RECT 1414.105 1582.535 1414.435 1582.550 ;
      LAYER met3 ;
        RECT 303.990 1579.240 1396.000 1581.920 ;
        RECT 304.400 1577.840 1396.000 1579.240 ;
        RECT 303.990 1572.440 1396.000 1577.840 ;
        RECT 303.990 1571.040 1395.600 1572.440 ;
      LAYER met3 ;
        RECT 1396.000 1571.970 1400.000 1572.040 ;
        RECT 1414.105 1571.970 1414.435 1571.985 ;
        RECT 1396.000 1571.670 1414.435 1571.970 ;
        RECT 1396.000 1571.440 1400.000 1571.670 ;
        RECT 1414.105 1571.655 1414.435 1571.670 ;
      LAYER met3 ;
        RECT 303.990 1568.360 1396.000 1571.040 ;
        RECT 304.400 1566.960 1396.000 1568.360 ;
        RECT 303.990 1560.880 1396.000 1566.960 ;
        RECT 303.990 1559.480 1395.600 1560.880 ;
      LAYER met3 ;
        RECT 1396.000 1560.410 1400.000 1560.480 ;
        RECT 1411.805 1560.410 1412.135 1560.425 ;
        RECT 1396.000 1560.110 1412.135 1560.410 ;
        RECT 1396.000 1559.880 1400.000 1560.110 ;
        RECT 1411.805 1560.095 1412.135 1560.110 ;
      LAYER met3 ;
        RECT 303.990 1558.160 1396.000 1559.480 ;
        RECT 304.400 1556.760 1396.000 1558.160 ;
        RECT 303.990 1550.000 1396.000 1556.760 ;
        RECT 303.990 1548.600 1395.600 1550.000 ;
      LAYER met3 ;
        RECT 1396.000 1549.530 1400.000 1549.600 ;
        RECT 1409.505 1549.530 1409.835 1549.545 ;
        RECT 1396.000 1549.230 1409.835 1549.530 ;
        RECT 1396.000 1549.000 1400.000 1549.230 ;
        RECT 1409.505 1549.215 1409.835 1549.230 ;
      LAYER met3 ;
        RECT 303.990 1547.280 1396.000 1548.600 ;
        RECT 304.400 1545.880 1396.000 1547.280 ;
        RECT 303.990 1539.120 1396.000 1545.880 ;
        RECT 303.990 1537.720 1395.600 1539.120 ;
      LAYER met3 ;
        RECT 1396.000 1538.650 1400.000 1538.720 ;
        RECT 1414.105 1538.650 1414.435 1538.665 ;
        RECT 1396.000 1538.350 1414.435 1538.650 ;
        RECT 1396.000 1538.120 1400.000 1538.350 ;
        RECT 1414.105 1538.335 1414.435 1538.350 ;
      LAYER met3 ;
        RECT 303.990 1537.080 1396.000 1537.720 ;
        RECT 304.400 1535.680 1396.000 1537.080 ;
        RECT 303.990 1528.240 1396.000 1535.680 ;
        RECT 303.990 1526.840 1395.600 1528.240 ;
      LAYER met3 ;
        RECT 1396.000 1527.770 1400.000 1527.840 ;
        RECT 1410.425 1527.770 1410.755 1527.785 ;
        RECT 1396.000 1527.470 1410.755 1527.770 ;
        RECT 1396.000 1527.240 1400.000 1527.470 ;
        RECT 1410.425 1527.455 1410.755 1527.470 ;
      LAYER met3 ;
        RECT 303.990 1526.200 1396.000 1526.840 ;
        RECT 304.400 1524.800 1396.000 1526.200 ;
        RECT 303.990 1517.360 1396.000 1524.800 ;
        RECT 303.990 1516.000 1395.600 1517.360 ;
      LAYER met3 ;
        RECT 1396.000 1516.890 1400.000 1516.960 ;
        RECT 1407.665 1516.890 1407.995 1516.905 ;
        RECT 1396.000 1516.590 1407.995 1516.890 ;
        RECT 1396.000 1516.360 1400.000 1516.590 ;
        RECT 1407.665 1516.575 1407.995 1516.590 ;
      LAYER met3 ;
        RECT 304.400 1515.960 1395.600 1516.000 ;
        RECT 304.400 1514.600 1396.000 1515.960 ;
        RECT 303.990 1506.480 1396.000 1514.600 ;
        RECT 303.990 1505.800 1395.600 1506.480 ;
        RECT 304.400 1505.080 1395.600 1505.800 ;
      LAYER met3 ;
        RECT 1396.000 1506.010 1400.000 1506.080 ;
        RECT 1408.125 1506.010 1408.455 1506.025 ;
        RECT 1396.000 1505.710 1408.455 1506.010 ;
        RECT 1396.000 1505.480 1400.000 1505.710 ;
        RECT 1408.125 1505.695 1408.455 1505.710 ;
      LAYER met3 ;
        RECT 304.400 1504.400 1396.000 1505.080 ;
        RECT 303.990 1504.255 1396.000 1504.400 ;
      LAYER via3 ;
        RECT 646.140 3264.180 646.460 3264.500 ;
        RECT 668.220 3264.180 668.540 3264.500 ;
        RECT 1295.660 3264.180 1295.980 3264.500 ;
        RECT 1318.660 3264.180 1318.980 3264.500 ;
        RECT 1892.740 3264.180 1893.060 3264.500 ;
        RECT 1917.580 3264.180 1917.900 3264.500 ;
        RECT 2539.500 3264.180 2539.820 3264.500 ;
        RECT 2567.100 3264.180 2567.420 3264.500 ;
        RECT 1055.540 2799.740 1055.860 2800.060 ;
        RECT 1052.780 2799.060 1053.100 2799.380 ;
        RECT 1759.340 2796.340 1759.660 2796.660 ;
        RECT 1794.300 2796.340 1794.620 2796.660 ;
        RECT 337.020 2794.300 337.340 2794.620 ;
        RECT 348.980 2794.300 349.300 2794.620 ;
        RECT 361.860 2794.300 362.180 2794.620 ;
        RECT 368.300 2794.300 368.620 2794.620 ;
        RECT 374.740 2794.300 375.060 2794.620 ;
        RECT 379.340 2794.300 379.660 2794.620 ;
        RECT 386.700 2794.300 387.020 2794.620 ;
        RECT 392.220 2794.300 392.540 2794.620 ;
        RECT 396.820 2794.300 397.140 2794.620 ;
        RECT 403.260 2794.300 403.580 2794.620 ;
        RECT 410.620 2794.300 410.940 2794.620 ;
        RECT 414.300 2794.300 414.620 2794.620 ;
        RECT 423.500 2794.300 423.820 2794.620 ;
        RECT 427.180 2794.300 427.500 2794.620 ;
        RECT 428.100 2794.300 428.420 2794.620 ;
        RECT 433.620 2794.300 433.940 2794.620 ;
        RECT 440.980 2794.300 441.300 2794.620 ;
        RECT 444.660 2794.300 444.980 2794.620 ;
        RECT 445.580 2794.300 445.900 2794.620 ;
        RECT 450.180 2794.300 450.500 2794.620 ;
        RECT 456.620 2794.300 456.940 2794.620 ;
        RECT 462.140 2794.300 462.460 2794.620 ;
        RECT 467.660 2794.300 467.980 2794.620 ;
        RECT 473.180 2794.300 473.500 2794.620 ;
        RECT 476.860 2794.300 477.180 2794.620 ;
        RECT 483.300 2794.300 483.620 2794.620 ;
        RECT 491.580 2794.300 491.900 2794.620 ;
        RECT 498.020 2794.300 498.340 2794.620 ;
        RECT 500.780 2794.300 501.100 2794.620 ;
        RECT 509.980 2794.300 510.300 2794.620 ;
        RECT 513.660 2794.300 513.980 2794.620 ;
        RECT 516.420 2794.300 516.740 2794.620 ;
        RECT 520.100 2794.300 520.420 2794.620 ;
        RECT 523.780 2794.300 524.100 2794.620 ;
        RECT 526.540 2794.300 526.860 2794.620 ;
        RECT 530.220 2794.300 530.540 2794.620 ;
        RECT 535.740 2794.300 536.060 2794.620 ;
        RECT 538.500 2794.300 538.820 2794.620 ;
        RECT 542.180 2794.300 542.500 2794.620 ;
        RECT 547.700 2794.300 548.020 2794.620 ;
        RECT 1013.220 2794.300 1013.540 2794.620 ;
        RECT 1019.660 2794.300 1019.980 2794.620 ;
        RECT 1027.020 2794.300 1027.340 2794.620 ;
        RECT 1059.220 2794.300 1059.540 2794.620 ;
        RECT 1065.660 2794.300 1065.980 2794.620 ;
        RECT 1070.260 2794.300 1070.580 2794.620 ;
        RECT 1081.300 2794.300 1081.620 2794.620 ;
        RECT 1087.740 2794.300 1088.060 2794.620 ;
        RECT 1089.580 2794.300 1089.900 2794.620 ;
        RECT 1094.180 2794.300 1094.500 2794.620 ;
        RECT 1096.020 2794.300 1096.340 2794.620 ;
        RECT 1100.620 2794.300 1100.940 2794.620 ;
        RECT 1103.380 2794.300 1103.700 2794.620 ;
        RECT 1105.220 2794.300 1105.540 2794.620 ;
        RECT 1109.820 2794.300 1110.140 2794.620 ;
        RECT 1111.660 2794.300 1111.980 2794.620 ;
        RECT 1116.260 2794.300 1116.580 2794.620 ;
        RECT 1121.780 2794.300 1122.100 2794.620 ;
        RECT 1129.140 2794.300 1129.460 2794.620 ;
        RECT 1130.980 2794.300 1131.300 2794.620 ;
        RECT 1135.580 2794.300 1135.900 2794.620 ;
        RECT 1137.420 2794.300 1137.740 2794.620 ;
        RECT 1143.860 2794.300 1144.180 2794.620 ;
        RECT 1147.540 2794.300 1147.860 2794.620 ;
        RECT 1151.220 2794.300 1151.540 2794.620 ;
        RECT 1153.980 2794.300 1154.300 2794.620 ;
        RECT 1164.100 2794.300 1164.420 2794.620 ;
        RECT 1165.020 2794.300 1165.340 2794.620 ;
        RECT 1172.380 2794.300 1172.700 2794.620 ;
        RECT 1178.820 2794.300 1179.140 2794.620 ;
        RECT 1186.180 2794.300 1186.500 2794.620 ;
        RECT 1198.140 2794.300 1198.460 2794.620 ;
        RECT 1580.860 2794.300 1581.180 2794.620 ;
        RECT 1594.660 2794.300 1594.980 2794.620 ;
        RECT 1604.780 2794.300 1605.100 2794.620 ;
        RECT 1613.980 2794.300 1614.300 2794.620 ;
        RECT 1625.940 2794.300 1626.260 2794.620 ;
        RECT 1631.460 2794.300 1631.780 2794.620 ;
        RECT 1637.900 2794.300 1638.220 2794.620 ;
        RECT 1655.380 2794.300 1655.700 2794.620 ;
        RECT 1659.060 2794.300 1659.380 2794.620 ;
        RECT 1666.420 2794.300 1666.740 2794.620 ;
        RECT 1672.860 2794.300 1673.180 2794.620 ;
        RECT 1679.300 2794.300 1679.620 2794.620 ;
        RECT 1683.900 2794.300 1684.220 2794.620 ;
        RECT 1688.500 2794.300 1688.820 2794.620 ;
        RECT 1695.860 2794.300 1696.180 2794.620 ;
        RECT 1702.300 2794.300 1702.620 2794.620 ;
        RECT 1708.740 2794.300 1709.060 2794.620 ;
        RECT 1713.340 2794.300 1713.660 2794.620 ;
        RECT 1719.780 2794.300 1720.100 2794.620 ;
        RECT 1721.620 2794.300 1721.940 2794.620 ;
        RECT 1730.820 2794.300 1731.140 2794.620 ;
        RECT 1737.260 2794.300 1737.580 2794.620 ;
        RECT 1743.700 2794.300 1744.020 2794.620 ;
        RECT 1748.300 2794.300 1748.620 2794.620 ;
        RECT 1762.100 2794.300 1762.420 2794.620 ;
        RECT 2231.300 2794.300 2231.620 2794.620 ;
        RECT 2236.820 2794.300 2237.140 2794.620 ;
        RECT 2242.340 2794.300 2242.660 2794.620 ;
        RECT 2249.700 2794.300 2250.020 2794.620 ;
        RECT 2264.420 2794.300 2264.740 2794.620 ;
        RECT 2268.100 2794.300 2268.420 2794.620 ;
        RECT 2273.620 2794.300 2273.940 2794.620 ;
        RECT 2292.020 2794.300 2292.340 2794.620 ;
        RECT 2304.900 2794.300 2305.220 2794.620 ;
        RECT 2308.580 2794.300 2308.900 2794.620 ;
        RECT 2316.860 2794.300 2317.180 2794.620 ;
        RECT 2322.380 2794.300 2322.700 2794.620 ;
        RECT 2328.820 2794.300 2329.140 2794.620 ;
        RECT 2334.340 2794.300 2334.660 2794.620 ;
        RECT 2339.860 2794.300 2340.180 2794.620 ;
        RECT 2343.540 2794.300 2343.860 2794.620 ;
        RECT 2351.820 2794.300 2352.140 2794.620 ;
        RECT 2357.340 2794.300 2357.660 2794.620 ;
        RECT 2363.780 2794.300 2364.100 2794.620 ;
        RECT 2370.220 2794.300 2370.540 2794.620 ;
        RECT 2374.820 2794.300 2375.140 2794.620 ;
        RECT 2381.260 2794.300 2381.580 2794.620 ;
        RECT 2385.860 2794.300 2386.180 2794.620 ;
        RECT 2391.380 2794.300 2391.700 2794.620 ;
        RECT 2396.900 2794.300 2397.220 2794.620 ;
        RECT 2404.260 2794.300 2404.580 2794.620 ;
        RECT 2417.140 2794.300 2417.460 2794.620 ;
        RECT 2428.180 2794.300 2428.500 2794.620 ;
        RECT 2430.020 2794.300 2430.340 2794.620 ;
        RECT 350.820 2793.620 351.140 2793.940 ;
        RECT 405.100 2793.620 405.420 2793.940 ;
        RECT 408.780 2793.620 409.100 2793.940 ;
        RECT 420.740 2793.620 421.060 2793.940 ;
        RECT 431.780 2793.620 432.100 2793.940 ;
        RECT 439.140 2793.620 439.460 2793.940 ;
        RECT 501.700 2793.620 502.020 2793.940 ;
        RECT 507.220 2793.620 507.540 2793.940 ;
        RECT 531.140 2793.620 531.460 2793.940 ;
        RECT 543.100 2793.620 543.420 2793.940 ;
        RECT 981.020 2793.620 981.340 2793.940 ;
        RECT 1008.620 2793.620 1008.940 2793.940 ;
        RECT 1012.300 2793.620 1012.620 2793.940 ;
        RECT 1024.260 2793.620 1024.580 2793.940 ;
        RECT 1076.700 2793.620 1077.020 2793.940 ;
        RECT 1083.140 2793.620 1083.460 2793.940 ;
        RECT 1086.820 2793.620 1087.140 2793.940 ;
        RECT 1118.100 2793.620 1118.420 2793.940 ;
        RECT 1122.700 2793.620 1123.020 2793.940 ;
        RECT 1128.220 2793.620 1128.540 2793.940 ;
        RECT 1139.260 2793.620 1139.580 2793.940 ;
        RECT 1163.180 2793.620 1163.500 2793.940 ;
        RECT 1167.780 2793.620 1168.100 2793.940 ;
        RECT 1180.660 2793.620 1180.980 2793.940 ;
        RECT 1612.140 2793.620 1612.460 2793.940 ;
        RECT 1635.140 2793.620 1635.460 2793.940 ;
        RECT 1642.500 2793.620 1642.820 2793.940 ;
        RECT 1663.660 2793.620 1663.980 2793.940 ;
        RECT 1670.100 2793.620 1670.420 2793.940 ;
        RECT 1677.460 2793.620 1677.780 2793.940 ;
        RECT 1682.980 2793.620 1683.300 2793.940 ;
        RECT 1694.940 2793.620 1695.260 2793.940 ;
        RECT 1699.540 2793.620 1699.860 2793.940 ;
        RECT 1705.060 2793.620 1705.380 2793.940 ;
        RECT 1712.420 2793.620 1712.740 2793.940 ;
        RECT 1717.940 2793.620 1718.260 2793.940 ;
        RECT 1729.900 2793.620 1730.220 2793.940 ;
        RECT 1734.500 2793.620 1734.820 2793.940 ;
        RECT 1740.940 2793.620 1741.260 2793.940 ;
        RECT 1747.380 2793.620 1747.700 2793.940 ;
        RECT 1767.620 2793.620 1767.940 2793.940 ;
        RECT 1787.860 2793.620 1788.180 2793.940 ;
        RECT 2263.500 2793.620 2263.820 2793.940 ;
        RECT 2297.540 2793.620 2297.860 2793.940 ;
        RECT 2310.420 2793.620 2310.740 2793.940 ;
        RECT 2315.020 2793.620 2315.340 2793.940 ;
        RECT 2321.460 2793.620 2321.780 2793.940 ;
        RECT 2326.060 2793.620 2326.380 2793.940 ;
        RECT 2345.380 2793.620 2345.700 2793.940 ;
        RECT 2349.980 2793.620 2350.300 2793.940 ;
        RECT 2356.420 2793.620 2356.740 2793.940 ;
        RECT 2361.020 2793.620 2361.340 2793.940 ;
        RECT 2367.460 2793.620 2367.780 2793.940 ;
        RECT 2373.900 2793.620 2374.220 2793.940 ;
        RECT 2377.580 2793.620 2377.900 2793.940 ;
        RECT 2402.420 2793.620 2402.740 2793.940 ;
        RECT 2423.580 2793.620 2423.900 2793.940 ;
        RECT 509.060 2792.940 509.380 2793.260 ;
        RECT 987.460 2792.940 987.780 2793.260 ;
        RECT 1018.740 2792.940 1019.060 2793.260 ;
        RECT 1048.180 2792.940 1048.500 2793.260 ;
        RECT 1153.060 2792.940 1153.380 2793.260 ;
        RECT 1159.500 2792.940 1159.820 2793.260 ;
        RECT 1173.300 2792.940 1173.620 2793.260 ;
        RECT 1617.660 2792.940 1617.980 2793.260 ;
        RECT 1624.100 2792.940 1624.420 2793.260 ;
        RECT 1630.540 2792.940 1630.860 2793.260 ;
        RECT 1648.020 2792.940 1648.340 2793.260 ;
        RECT 1652.620 2792.940 1652.940 2793.260 ;
        RECT 1780.500 2792.940 1780.820 2793.260 ;
        RECT 2280.060 2792.940 2280.380 2793.260 ;
        RECT 2286.500 2792.940 2286.820 2793.260 ;
        RECT 2303.980 2792.940 2304.300 2793.260 ;
        RECT 2332.500 2792.940 2332.820 2793.260 ;
        RECT 2338.940 2792.940 2339.260 2793.260 ;
        RECT 2415.300 2792.940 2415.620 2793.260 ;
        RECT 2442.900 2792.940 2443.220 2793.260 ;
        RECT 993.900 2792.260 994.220 2792.580 ;
        RECT 1001.260 2792.260 1001.580 2792.580 ;
        RECT 1187.100 2792.260 1187.420 2792.580 ;
        RECT 1193.540 2792.260 1193.860 2792.580 ;
        RECT 1587.300 2792.260 1587.620 2792.580 ;
        RECT 1689.420 2792.260 1689.740 2792.580 ;
        RECT 1752.900 2792.260 1753.220 2792.580 ;
        RECT 2282.820 2792.260 2283.140 2792.580 ;
        RECT 2407.940 2792.260 2408.260 2792.580 ;
        RECT 2436.460 2792.260 2436.780 2792.580 ;
        RECT 388.540 2791.580 388.860 2791.900 ;
        RECT 417.060 2791.580 417.380 2791.900 ;
        RECT 1648.940 2791.580 1649.260 2791.900 ;
        RECT 1774.060 2791.580 1774.380 2791.900 ;
        RECT 2276.380 2791.580 2276.700 2791.900 ;
        RECT 2287.420 2791.580 2287.740 2791.900 ;
        RECT 2293.860 2791.580 2294.180 2791.900 ;
        RECT 2445.660 2791.580 2445.980 2791.900 ;
        RECT 371.060 2790.900 371.380 2791.220 ;
        RECT 1644.340 2790.900 1644.660 2791.220 ;
        RECT 1661.820 2790.900 1662.140 2791.220 ;
        RECT 2269.020 2790.900 2269.340 2791.220 ;
        RECT 2299.380 2790.900 2299.700 2791.220 ;
        RECT 2420.820 2790.900 2421.140 2791.220 ;
        RECT 2434.620 2790.900 2434.940 2791.220 ;
        RECT 2439.220 2790.900 2439.540 2791.220 ;
        RECT 342.540 2790.220 342.860 2790.540 ;
        RECT 1030.700 2790.220 1031.020 2790.540 ;
        RECT 1191.700 2790.220 1192.020 2790.540 ;
        RECT 2386.780 2790.220 2387.100 2790.540 ;
        RECT 2392.300 2790.220 2392.620 2790.540 ;
        RECT 393.140 2789.540 393.460 2789.860 ;
        RECT 1620.420 2789.540 1620.740 2789.860 ;
        RECT 2398.740 2789.540 2399.060 2789.860 ;
        RECT 375.660 2788.860 375.980 2789.180 ;
        RECT 382.100 2788.860 382.420 2789.180 ;
        RECT 1601.100 2788.860 1601.420 2789.180 ;
        RECT 2410.700 2788.860 2411.020 2789.180 ;
        RECT 364.620 2788.180 364.940 2788.500 ;
        RECT 399.580 2788.180 399.900 2788.500 ;
        RECT 465.820 2788.180 466.140 2788.500 ;
        RECT 1035.300 2788.180 1035.620 2788.500 ;
        RECT 1041.740 2788.180 1042.060 2788.500 ;
        RECT 1051.860 2788.180 1052.180 2788.500 ;
        RECT 1724.380 2788.180 1724.700 2788.500 ;
        RECT 1765.780 2788.180 1766.100 2788.500 ;
        RECT 2257.060 2788.180 2257.380 2788.500 ;
        RECT 2377.580 2788.180 2377.900 2788.500 ;
        RECT 2418.060 2788.180 2418.380 2788.500 ;
        RECT 357.260 2787.500 357.580 2787.820 ;
        RECT 454.780 2787.500 455.100 2787.820 ;
        RECT 460.300 2787.500 460.620 2787.820 ;
        RECT 468.580 2787.500 468.900 2787.820 ;
        RECT 475.020 2787.500 475.340 2787.820 ;
        RECT 482.380 2787.500 482.700 2787.820 ;
        RECT 488.820 2787.500 489.140 2787.820 ;
        RECT 495.260 2787.500 495.580 2787.820 ;
        RECT 1034.380 2787.500 1034.700 2787.820 ;
        RECT 1039.900 2787.500 1040.220 2787.820 ;
        RECT 1046.340 2787.500 1046.660 2787.820 ;
        RECT 1061.980 2787.500 1062.300 2787.820 ;
        RECT 1067.500 2787.500 1067.820 2787.820 ;
        RECT 1073.940 2787.500 1074.260 2787.820 ;
        RECT 1754.740 2787.500 1755.060 2787.820 ;
        RECT 1772.220 2787.500 1772.540 2787.820 ;
        RECT 1777.740 2787.500 1778.060 2787.820 ;
        RECT 1783.260 2787.500 1783.580 2787.820 ;
        RECT 1789.700 2787.500 1790.020 2787.820 ;
        RECT 1761.180 2777.300 1761.500 2777.620 ;
        RECT 1796.140 2777.300 1796.460 2777.620 ;
      LAYER met4 ;
        RECT 646.135 3264.175 646.465 3264.505 ;
        RECT 668.215 3264.175 668.545 3264.505 ;
        RECT 1295.655 3264.175 1295.985 3264.505 ;
        RECT 1318.655 3264.175 1318.985 3264.505 ;
        RECT 1892.735 3264.175 1893.065 3264.505 ;
        RECT 1917.575 3264.175 1917.905 3264.505 ;
        RECT 2539.495 3264.175 2539.825 3264.505 ;
        RECT 2567.095 3264.175 2567.425 3264.505 ;
        RECT 394.025 3251.635 394.325 3256.235 ;
        RECT 400.265 3251.635 400.565 3256.235 ;
        RECT 406.505 3251.635 406.805 3256.235 ;
        RECT 412.745 3251.635 413.045 3256.235 ;
        RECT 418.985 3251.635 419.285 3256.235 ;
        RECT 425.225 3251.635 425.525 3256.235 ;
        RECT 431.465 3251.635 431.765 3256.235 ;
        RECT 437.705 3251.635 438.005 3256.235 ;
        RECT 443.945 3251.635 444.245 3256.235 ;
        RECT 450.185 3251.635 450.485 3256.235 ;
        RECT 456.425 3251.635 456.725 3256.235 ;
        RECT 462.665 3251.635 462.965 3256.235 ;
        RECT 468.905 3251.635 469.205 3256.235 ;
        RECT 475.145 3251.635 475.445 3256.235 ;
        RECT 481.385 3251.635 481.685 3256.235 ;
        RECT 487.625 3251.635 487.925 3256.235 ;
        RECT 493.865 3251.635 494.165 3256.235 ;
        RECT 500.105 3251.635 500.405 3256.235 ;
        RECT 506.345 3251.635 506.645 3256.235 ;
        RECT 512.585 3251.635 512.885 3256.235 ;
        RECT 518.825 3251.635 519.125 3256.235 ;
        RECT 525.065 3251.635 525.365 3256.235 ;
        RECT 531.305 3251.635 531.605 3256.235 ;
        RECT 537.545 3251.635 537.845 3256.235 ;
        RECT 543.785 3251.635 544.085 3256.235 ;
        RECT 550.025 3251.635 550.325 3256.235 ;
        RECT 556.265 3251.635 556.565 3256.235 ;
        RECT 562.505 3251.635 562.805 3256.235 ;
        RECT 568.745 3251.635 569.045 3256.235 ;
        RECT 574.985 3251.635 575.285 3256.235 ;
        RECT 581.225 3251.635 581.525 3256.235 ;
        RECT 587.465 3251.635 587.765 3256.235 ;
        RECT 642.890 3255.650 643.190 3256.235 ;
        RECT 646.150 3255.650 646.450 3264.175 ;
        RECT 668.230 3259.050 668.530 3264.175 ;
        RECT 642.890 3255.350 646.450 3255.650 ;
        RECT 667.865 3258.750 668.530 3259.050 ;
        RECT 642.890 3251.635 643.190 3255.350 ;
        RECT 667.865 3251.635 668.165 3258.750 ;
        RECT 1044.025 3251.635 1044.325 3256.235 ;
        RECT 1050.265 3251.635 1050.565 3256.235 ;
        RECT 1056.505 3251.635 1056.805 3256.235 ;
        RECT 1062.745 3251.635 1063.045 3256.235 ;
        RECT 1068.985 3251.635 1069.285 3256.235 ;
        RECT 1075.225 3251.635 1075.525 3256.235 ;
        RECT 1081.465 3251.635 1081.765 3256.235 ;
        RECT 1087.705 3251.635 1088.005 3256.235 ;
        RECT 1093.945 3251.635 1094.245 3256.235 ;
        RECT 1100.185 3251.635 1100.485 3256.235 ;
        RECT 1106.425 3251.635 1106.725 3256.235 ;
        RECT 1112.665 3251.635 1112.965 3256.235 ;
        RECT 1118.905 3251.635 1119.205 3256.235 ;
        RECT 1125.145 3251.635 1125.445 3256.235 ;
        RECT 1131.385 3251.635 1131.685 3256.235 ;
        RECT 1137.625 3251.635 1137.925 3256.235 ;
        RECT 1143.865 3251.635 1144.165 3256.235 ;
        RECT 1150.105 3251.635 1150.405 3256.235 ;
        RECT 1156.345 3251.635 1156.645 3256.235 ;
        RECT 1162.585 3251.635 1162.885 3256.235 ;
        RECT 1168.825 3251.635 1169.125 3256.235 ;
        RECT 1175.065 3251.635 1175.365 3256.235 ;
        RECT 1181.305 3251.635 1181.605 3256.235 ;
        RECT 1187.545 3251.635 1187.845 3256.235 ;
        RECT 1193.785 3251.635 1194.085 3256.235 ;
        RECT 1200.025 3251.635 1200.325 3256.235 ;
        RECT 1206.265 3251.635 1206.565 3256.235 ;
        RECT 1212.505 3251.635 1212.805 3256.235 ;
        RECT 1218.745 3251.635 1219.045 3256.235 ;
        RECT 1224.985 3251.635 1225.285 3256.235 ;
        RECT 1231.225 3251.635 1231.525 3256.235 ;
        RECT 1237.465 3251.635 1237.765 3256.235 ;
        RECT 1292.890 3255.650 1293.190 3256.235 ;
        RECT 1295.670 3255.650 1295.970 3264.175 ;
        RECT 1292.890 3255.350 1295.970 3255.650 ;
        RECT 1317.865 3255.650 1318.165 3256.235 ;
        RECT 1318.670 3255.650 1318.970 3264.175 ;
        RECT 1892.750 3256.235 1893.050 3264.175 ;
        RECT 1917.590 3256.235 1917.890 3264.175 ;
        RECT 1317.865 3255.350 1318.970 3255.650 ;
        RECT 1292.890 3251.635 1293.190 3255.350 ;
        RECT 1317.865 3251.635 1318.165 3255.350 ;
        RECT 1644.025 3251.635 1644.325 3256.235 ;
        RECT 1650.265 3251.635 1650.565 3256.235 ;
        RECT 1656.505 3251.635 1656.805 3256.235 ;
        RECT 1662.745 3251.635 1663.045 3256.235 ;
        RECT 1668.985 3251.635 1669.285 3256.235 ;
        RECT 1675.225 3251.635 1675.525 3256.235 ;
        RECT 1681.465 3251.635 1681.765 3256.235 ;
        RECT 1687.705 3251.635 1688.005 3256.235 ;
        RECT 1693.945 3251.635 1694.245 3256.235 ;
        RECT 1700.185 3251.635 1700.485 3256.235 ;
        RECT 1706.425 3251.635 1706.725 3256.235 ;
        RECT 1712.665 3251.635 1712.965 3256.235 ;
        RECT 1718.905 3251.635 1719.205 3256.235 ;
        RECT 1725.145 3251.635 1725.445 3256.235 ;
        RECT 1731.385 3251.635 1731.685 3256.235 ;
        RECT 1737.625 3251.635 1737.925 3256.235 ;
        RECT 1743.865 3251.635 1744.165 3256.235 ;
        RECT 1750.105 3251.635 1750.405 3256.235 ;
        RECT 1756.345 3251.635 1756.645 3256.235 ;
        RECT 1762.585 3251.635 1762.885 3256.235 ;
        RECT 1768.825 3251.635 1769.125 3256.235 ;
        RECT 1775.065 3251.635 1775.365 3256.235 ;
        RECT 1781.305 3251.635 1781.605 3256.235 ;
        RECT 1787.545 3251.635 1787.845 3256.235 ;
        RECT 1793.785 3251.635 1794.085 3256.235 ;
        RECT 1800.025 3251.635 1800.325 3256.235 ;
        RECT 1806.265 3251.635 1806.565 3256.235 ;
        RECT 1812.505 3251.635 1812.805 3256.235 ;
        RECT 1818.745 3251.635 1819.045 3256.235 ;
        RECT 1824.985 3251.635 1825.285 3256.235 ;
        RECT 1831.225 3251.635 1831.525 3256.235 ;
        RECT 1837.465 3251.635 1837.765 3256.235 ;
        RECT 1892.750 3255.350 1893.190 3256.235 ;
        RECT 1917.590 3255.350 1918.165 3256.235 ;
        RECT 1892.890 3251.635 1893.190 3255.350 ;
        RECT 1917.865 3251.635 1918.165 3255.350 ;
        RECT 2294.025 3251.635 2294.325 3256.235 ;
        RECT 2300.265 3251.635 2300.565 3256.235 ;
        RECT 2306.505 3251.635 2306.805 3256.235 ;
        RECT 2312.745 3251.635 2313.045 3256.235 ;
        RECT 2318.985 3251.635 2319.285 3256.235 ;
        RECT 2325.225 3251.635 2325.525 3256.235 ;
        RECT 2331.465 3251.635 2331.765 3256.235 ;
        RECT 2337.705 3251.635 2338.005 3256.235 ;
        RECT 2343.945 3251.635 2344.245 3256.235 ;
        RECT 2350.185 3251.635 2350.485 3256.235 ;
        RECT 2356.425 3251.635 2356.725 3256.235 ;
        RECT 2362.665 3251.635 2362.965 3256.235 ;
        RECT 2368.905 3251.635 2369.205 3256.235 ;
        RECT 2375.145 3251.635 2375.445 3256.235 ;
        RECT 2381.385 3251.635 2381.685 3256.235 ;
        RECT 2387.625 3251.635 2387.925 3256.235 ;
        RECT 2393.865 3251.635 2394.165 3256.235 ;
        RECT 2400.105 3251.635 2400.405 3256.235 ;
        RECT 2406.345 3251.635 2406.645 3256.235 ;
        RECT 2412.585 3251.635 2412.885 3256.235 ;
        RECT 2418.825 3251.635 2419.125 3256.235 ;
        RECT 2425.065 3251.635 2425.365 3256.235 ;
        RECT 2431.305 3251.635 2431.605 3256.235 ;
        RECT 2437.545 3251.635 2437.845 3256.235 ;
        RECT 2443.785 3251.635 2444.085 3256.235 ;
        RECT 2450.025 3251.635 2450.325 3256.235 ;
        RECT 2456.265 3251.635 2456.565 3256.235 ;
        RECT 2462.505 3251.635 2462.805 3256.235 ;
        RECT 2468.745 3251.635 2469.045 3256.235 ;
        RECT 2474.985 3251.635 2475.285 3256.235 ;
        RECT 2481.225 3251.635 2481.525 3256.235 ;
        RECT 2487.465 3251.635 2487.765 3256.235 ;
        RECT 2539.510 3255.650 2539.810 3264.175 ;
        RECT 2542.890 3255.650 2543.190 3256.235 ;
        RECT 2539.510 3255.350 2543.190 3255.650 ;
        RECT 2567.110 3255.650 2567.410 3264.175 ;
        RECT 2567.865 3255.650 2568.165 3256.235 ;
        RECT 2567.110 3255.350 2568.165 3255.650 ;
        RECT 2542.890 3251.635 2543.190 3255.350 ;
        RECT 2567.865 3251.635 2568.165 3255.350 ;
      LAYER met4 ;
        RECT 305.000 2805.000 681.480 3251.235 ;
        RECT 955.000 2805.000 1331.480 3251.235 ;
        RECT 1555.000 2805.000 1931.480 3251.235 ;
        RECT 2205.000 2805.000 2581.480 3251.235 ;
      LAYER met4 ;
        RECT 334.010 2801.750 334.310 2804.600 ;
        RECT 339.850 2801.750 340.150 2804.600 ;
        RECT 345.690 2801.750 345.990 2804.600 ;
        RECT 351.530 2801.750 351.830 2804.600 ;
        RECT 357.370 2801.750 357.670 2804.600 ;
        RECT 363.210 2802.450 363.510 2804.600 ;
        RECT 334.010 2801.450 337.330 2801.750 ;
        RECT 334.010 2800.000 334.310 2801.450 ;
        RECT 337.030 2794.625 337.330 2801.450 ;
        RECT 339.850 2801.450 342.850 2801.750 ;
        RECT 339.850 2800.000 340.150 2801.450 ;
        RECT 337.015 2794.295 337.345 2794.625 ;
        RECT 342.550 2790.545 342.850 2801.450 ;
        RECT 345.690 2801.450 349.290 2801.750 ;
        RECT 345.690 2800.000 345.990 2801.450 ;
        RECT 348.990 2794.625 349.290 2801.450 ;
        RECT 350.830 2801.450 351.830 2801.750 ;
        RECT 348.975 2794.295 349.305 2794.625 ;
        RECT 350.830 2793.945 351.130 2801.450 ;
        RECT 351.530 2800.000 351.830 2801.450 ;
        RECT 357.270 2800.000 357.670 2801.750 ;
        RECT 361.870 2802.150 363.510 2802.450 ;
        RECT 350.815 2793.615 351.145 2793.945 ;
        RECT 342.535 2790.215 342.865 2790.545 ;
        RECT 357.270 2787.825 357.570 2800.000 ;
        RECT 361.870 2794.625 362.170 2802.150 ;
        RECT 363.210 2800.000 363.510 2802.150 ;
        RECT 363.830 2801.750 364.130 2804.600 ;
        RECT 369.050 2801.750 369.350 2804.600 ;
        RECT 363.830 2801.450 364.930 2801.750 ;
        RECT 363.830 2800.000 364.130 2801.450 ;
        RECT 361.855 2794.295 362.185 2794.625 ;
        RECT 364.630 2788.505 364.930 2801.450 ;
        RECT 368.310 2801.450 369.350 2801.750 ;
        RECT 368.310 2794.625 368.610 2801.450 ;
        RECT 369.050 2800.000 369.350 2801.450 ;
        RECT 369.670 2802.450 369.970 2804.600 ;
        RECT 369.670 2802.150 371.370 2802.450 ;
        RECT 369.670 2800.000 369.970 2802.150 ;
        RECT 368.295 2794.295 368.625 2794.625 ;
        RECT 371.070 2791.225 371.370 2802.150 ;
        RECT 374.890 2801.750 375.190 2804.600 ;
        RECT 374.750 2800.000 375.190 2801.750 ;
        RECT 375.510 2801.750 375.810 2804.600 ;
        RECT 380.730 2802.450 381.030 2804.600 ;
        RECT 379.350 2802.150 381.030 2802.450 ;
        RECT 375.510 2800.000 375.970 2801.750 ;
        RECT 374.750 2794.625 375.050 2800.000 ;
        RECT 374.735 2794.295 375.065 2794.625 ;
        RECT 371.055 2790.895 371.385 2791.225 ;
        RECT 375.670 2789.185 375.970 2800.000 ;
        RECT 379.350 2794.625 379.650 2802.150 ;
        RECT 380.730 2800.000 381.030 2802.150 ;
        RECT 381.350 2801.750 381.650 2804.600 ;
        RECT 381.350 2801.450 382.410 2801.750 ;
        RECT 381.350 2800.000 381.650 2801.450 ;
        RECT 379.335 2794.295 379.665 2794.625 ;
        RECT 382.110 2789.185 382.410 2801.450 ;
        RECT 386.570 2796.650 386.870 2804.600 ;
        RECT 387.190 2802.450 387.490 2804.600 ;
        RECT 387.190 2802.150 388.850 2802.450 ;
        RECT 387.190 2800.000 387.490 2802.150 ;
        RECT 386.570 2796.350 387.010 2796.650 ;
        RECT 386.710 2794.625 387.010 2796.350 ;
        RECT 386.695 2794.295 387.025 2794.625 ;
        RECT 388.550 2791.905 388.850 2802.150 ;
        RECT 392.410 2801.750 392.710 2804.600 ;
        RECT 392.230 2800.000 392.710 2801.750 ;
        RECT 393.030 2801.750 393.330 2804.600 ;
        RECT 398.250 2802.450 398.550 2804.600 ;
        RECT 396.830 2802.150 398.550 2802.450 ;
        RECT 393.030 2800.000 393.450 2801.750 ;
        RECT 392.230 2794.625 392.530 2800.000 ;
        RECT 392.215 2794.295 392.545 2794.625 ;
        RECT 388.535 2791.575 388.865 2791.905 ;
        RECT 393.150 2789.865 393.450 2800.000 ;
        RECT 396.830 2794.625 397.130 2802.150 ;
        RECT 398.250 2800.000 398.550 2802.150 ;
        RECT 398.870 2801.750 399.170 2804.600 ;
        RECT 404.090 2801.750 404.390 2804.600 ;
        RECT 398.870 2801.450 399.890 2801.750 ;
        RECT 398.870 2800.000 399.170 2801.450 ;
        RECT 396.815 2794.295 397.145 2794.625 ;
        RECT 393.135 2789.535 393.465 2789.865 ;
        RECT 375.655 2788.855 375.985 2789.185 ;
        RECT 382.095 2788.855 382.425 2789.185 ;
        RECT 399.590 2788.505 399.890 2801.450 ;
        RECT 403.270 2801.450 404.390 2801.750 ;
        RECT 403.270 2794.625 403.570 2801.450 ;
        RECT 404.090 2800.000 404.390 2801.450 ;
        RECT 404.710 2800.050 405.010 2804.600 ;
        RECT 409.930 2801.750 410.230 2804.600 ;
        RECT 408.790 2801.450 410.230 2801.750 ;
        RECT 404.710 2799.750 405.410 2800.050 ;
        RECT 403.255 2794.295 403.585 2794.625 ;
        RECT 405.110 2793.945 405.410 2799.750 ;
        RECT 408.790 2793.945 409.090 2801.450 ;
        RECT 409.930 2800.000 410.230 2801.450 ;
        RECT 410.550 2801.750 410.850 2804.600 ;
        RECT 415.770 2802.450 416.070 2804.600 ;
        RECT 414.310 2802.150 416.070 2802.450 ;
        RECT 410.550 2800.000 410.930 2801.750 ;
        RECT 410.630 2794.625 410.930 2800.000 ;
        RECT 414.310 2794.625 414.610 2802.150 ;
        RECT 415.770 2800.000 416.070 2802.150 ;
        RECT 416.390 2801.750 416.690 2804.600 ;
        RECT 421.610 2801.750 421.910 2804.600 ;
        RECT 416.390 2801.450 417.370 2801.750 ;
        RECT 416.390 2800.000 416.690 2801.450 ;
        RECT 410.615 2794.295 410.945 2794.625 ;
        RECT 414.295 2794.295 414.625 2794.625 ;
        RECT 405.095 2793.615 405.425 2793.945 ;
        RECT 408.775 2793.615 409.105 2793.945 ;
        RECT 417.070 2791.905 417.370 2801.450 ;
        RECT 420.750 2801.450 421.910 2801.750 ;
        RECT 420.750 2793.945 421.050 2801.450 ;
        RECT 421.610 2800.000 421.910 2801.450 ;
        RECT 422.230 2802.450 422.530 2804.600 ;
        RECT 422.230 2802.150 423.810 2802.450 ;
        RECT 422.230 2800.000 422.530 2802.150 ;
        RECT 423.510 2794.625 423.810 2802.150 ;
        RECT 427.450 2801.750 427.750 2804.600 ;
        RECT 427.190 2800.000 427.750 2801.750 ;
        RECT 428.070 2801.750 428.370 2804.600 ;
        RECT 433.290 2802.450 433.590 2804.600 ;
        RECT 431.790 2802.150 433.590 2802.450 ;
        RECT 428.070 2800.000 428.410 2801.750 ;
        RECT 427.190 2794.625 427.490 2800.000 ;
        RECT 428.110 2794.625 428.410 2800.000 ;
        RECT 423.495 2794.295 423.825 2794.625 ;
        RECT 427.175 2794.295 427.505 2794.625 ;
        RECT 428.095 2794.295 428.425 2794.625 ;
        RECT 431.790 2793.945 432.090 2802.150 ;
        RECT 433.290 2800.000 433.590 2802.150 ;
        RECT 433.910 2796.650 434.210 2804.600 ;
        RECT 439.130 2800.050 439.430 2804.600 ;
        RECT 439.750 2802.450 440.050 2804.600 ;
        RECT 439.750 2802.150 441.290 2802.450 ;
        RECT 439.130 2799.750 439.450 2800.050 ;
        RECT 439.750 2800.000 440.050 2802.150 ;
        RECT 433.630 2796.350 434.210 2796.650 ;
        RECT 433.630 2794.625 433.930 2796.350 ;
        RECT 433.615 2794.295 433.945 2794.625 ;
        RECT 439.150 2793.945 439.450 2799.750 ;
        RECT 440.990 2794.625 441.290 2802.150 ;
        RECT 444.970 2801.750 445.270 2804.600 ;
        RECT 444.670 2800.000 445.270 2801.750 ;
        RECT 444.670 2794.625 444.970 2800.000 ;
        RECT 445.590 2794.625 445.890 2804.600 ;
        RECT 450.810 2801.750 451.110 2804.600 ;
        RECT 450.190 2801.450 451.110 2801.750 ;
        RECT 450.190 2794.625 450.490 2801.450 ;
        RECT 450.810 2800.000 451.110 2801.450 ;
        RECT 451.430 2801.750 451.730 2804.600 ;
        RECT 456.650 2801.750 456.950 2804.600 ;
        RECT 451.430 2801.450 455.090 2801.750 ;
        RECT 451.430 2800.000 451.730 2801.450 ;
        RECT 440.975 2794.295 441.305 2794.625 ;
        RECT 444.655 2794.295 444.985 2794.625 ;
        RECT 445.575 2794.295 445.905 2794.625 ;
        RECT 450.175 2794.295 450.505 2794.625 ;
        RECT 420.735 2793.615 421.065 2793.945 ;
        RECT 431.775 2793.615 432.105 2793.945 ;
        RECT 439.135 2793.615 439.465 2793.945 ;
        RECT 417.055 2791.575 417.385 2791.905 ;
        RECT 364.615 2788.175 364.945 2788.505 ;
        RECT 399.575 2788.175 399.905 2788.505 ;
        RECT 454.790 2787.825 455.090 2801.450 ;
        RECT 456.630 2800.000 456.950 2801.750 ;
        RECT 457.270 2801.750 457.570 2804.600 ;
        RECT 457.270 2801.450 460.610 2801.750 ;
        RECT 457.270 2800.000 457.570 2801.450 ;
        RECT 456.630 2794.625 456.930 2800.000 ;
        RECT 456.615 2794.295 456.945 2794.625 ;
        RECT 460.310 2787.825 460.610 2801.450 ;
        RECT 462.490 2800.050 462.790 2804.600 ;
        RECT 462.150 2799.750 462.790 2800.050 ;
        RECT 463.110 2801.750 463.410 2804.600 ;
        RECT 468.330 2801.750 468.630 2804.600 ;
        RECT 463.110 2801.450 466.130 2801.750 ;
        RECT 463.110 2800.000 463.410 2801.450 ;
        RECT 462.150 2794.625 462.450 2799.750 ;
        RECT 462.135 2794.295 462.465 2794.625 ;
        RECT 465.830 2788.505 466.130 2801.450 ;
        RECT 467.670 2801.450 468.630 2801.750 ;
        RECT 467.670 2794.625 467.970 2801.450 ;
        RECT 468.330 2800.000 468.630 2801.450 ;
        RECT 468.950 2796.650 469.250 2804.600 ;
        RECT 474.170 2801.750 474.470 2804.600 ;
        RECT 468.590 2796.350 469.250 2796.650 ;
        RECT 473.190 2801.450 474.470 2801.750 ;
        RECT 467.655 2794.295 467.985 2794.625 ;
        RECT 465.815 2788.175 466.145 2788.505 ;
        RECT 468.590 2787.825 468.890 2796.350 ;
        RECT 473.190 2794.625 473.490 2801.450 ;
        RECT 474.170 2800.000 474.470 2801.450 ;
        RECT 474.790 2801.750 475.090 2804.600 ;
        RECT 480.010 2801.750 480.310 2804.600 ;
        RECT 474.790 2800.000 475.330 2801.750 ;
        RECT 473.175 2794.295 473.505 2794.625 ;
        RECT 475.030 2787.825 475.330 2800.000 ;
        RECT 476.870 2801.450 480.310 2801.750 ;
        RECT 476.870 2794.625 477.170 2801.450 ;
        RECT 480.010 2800.000 480.310 2801.450 ;
        RECT 480.630 2801.750 480.930 2804.600 ;
        RECT 485.850 2801.750 486.150 2804.600 ;
        RECT 480.630 2801.450 482.690 2801.750 ;
        RECT 480.630 2800.000 480.930 2801.450 ;
        RECT 476.855 2794.295 477.185 2794.625 ;
        RECT 482.390 2787.825 482.690 2801.450 ;
        RECT 483.310 2801.450 486.150 2801.750 ;
        RECT 483.310 2794.625 483.610 2801.450 ;
        RECT 485.850 2800.000 486.150 2801.450 ;
        RECT 486.470 2801.750 486.770 2804.600 ;
        RECT 491.690 2801.750 491.990 2804.600 ;
        RECT 486.470 2801.450 489.130 2801.750 ;
        RECT 486.470 2800.000 486.770 2801.450 ;
        RECT 483.295 2794.295 483.625 2794.625 ;
        RECT 488.830 2787.825 489.130 2801.450 ;
        RECT 491.590 2800.000 491.990 2801.750 ;
        RECT 492.310 2801.750 492.610 2804.600 ;
        RECT 492.310 2801.450 495.570 2801.750 ;
        RECT 492.310 2800.000 492.610 2801.450 ;
        RECT 491.590 2794.625 491.890 2800.000 ;
        RECT 491.575 2794.295 491.905 2794.625 ;
        RECT 495.270 2787.825 495.570 2801.450 ;
        RECT 497.530 2796.650 497.830 2804.600 ;
        RECT 498.150 2801.750 498.450 2804.600 ;
        RECT 503.370 2801.750 503.670 2804.600 ;
        RECT 498.150 2801.450 501.090 2801.750 ;
        RECT 498.150 2800.000 498.450 2801.450 ;
        RECT 497.530 2796.350 498.330 2796.650 ;
        RECT 498.030 2794.625 498.330 2796.350 ;
        RECT 500.790 2794.625 501.090 2801.450 ;
        RECT 501.710 2801.450 503.670 2801.750 ;
        RECT 498.015 2794.295 498.345 2794.625 ;
        RECT 500.775 2794.295 501.105 2794.625 ;
        RECT 501.710 2793.945 502.010 2801.450 ;
        RECT 503.370 2800.000 503.670 2801.450 ;
        RECT 503.990 2801.750 504.290 2804.600 ;
        RECT 509.210 2801.750 509.510 2804.600 ;
        RECT 503.990 2801.450 507.530 2801.750 ;
        RECT 503.990 2800.000 504.290 2801.450 ;
        RECT 507.230 2793.945 507.530 2801.450 ;
        RECT 509.070 2800.000 509.510 2801.750 ;
        RECT 509.830 2801.750 510.130 2804.600 ;
        RECT 515.050 2802.450 515.350 2804.600 ;
        RECT 513.670 2802.150 515.350 2802.450 ;
        RECT 509.830 2800.000 510.290 2801.750 ;
        RECT 501.695 2793.615 502.025 2793.945 ;
        RECT 507.215 2793.615 507.545 2793.945 ;
        RECT 509.070 2793.265 509.370 2800.000 ;
        RECT 509.990 2794.625 510.290 2800.000 ;
        RECT 513.670 2794.625 513.970 2802.150 ;
        RECT 515.050 2800.000 515.350 2802.150 ;
        RECT 515.670 2801.750 515.970 2804.600 ;
        RECT 520.890 2801.750 521.190 2804.600 ;
        RECT 515.670 2801.450 516.730 2801.750 ;
        RECT 515.670 2800.000 515.970 2801.450 ;
        RECT 516.430 2794.625 516.730 2801.450 ;
        RECT 520.110 2801.450 521.190 2801.750 ;
        RECT 520.110 2794.625 520.410 2801.450 ;
        RECT 520.890 2800.000 521.190 2801.450 ;
        RECT 521.510 2801.750 521.810 2804.600 ;
        RECT 526.730 2801.750 527.030 2804.600 ;
        RECT 521.510 2801.450 524.090 2801.750 ;
        RECT 521.510 2800.000 521.810 2801.450 ;
        RECT 523.790 2794.625 524.090 2801.450 ;
        RECT 526.550 2800.000 527.030 2801.750 ;
        RECT 527.350 2801.750 527.650 2804.600 ;
        RECT 532.570 2802.450 532.870 2804.600 ;
        RECT 531.150 2802.150 532.870 2802.450 ;
        RECT 527.350 2801.450 530.530 2801.750 ;
        RECT 527.350 2800.000 527.650 2801.450 ;
        RECT 526.550 2794.625 526.850 2800.000 ;
        RECT 530.230 2794.625 530.530 2801.450 ;
        RECT 509.975 2794.295 510.305 2794.625 ;
        RECT 513.655 2794.295 513.985 2794.625 ;
        RECT 516.415 2794.295 516.745 2794.625 ;
        RECT 520.095 2794.295 520.425 2794.625 ;
        RECT 523.775 2794.295 524.105 2794.625 ;
        RECT 526.535 2794.295 526.865 2794.625 ;
        RECT 530.215 2794.295 530.545 2794.625 ;
        RECT 531.150 2793.945 531.450 2802.150 ;
        RECT 532.570 2800.000 532.870 2802.150 ;
        RECT 533.190 2801.750 533.490 2804.600 ;
        RECT 533.190 2801.450 536.050 2801.750 ;
        RECT 533.190 2800.000 533.490 2801.450 ;
        RECT 535.750 2794.625 536.050 2801.450 ;
        RECT 538.410 2796.650 538.710 2804.600 ;
        RECT 539.030 2801.750 539.330 2804.600 ;
        RECT 544.250 2801.750 544.550 2804.600 ;
        RECT 539.030 2801.450 542.490 2801.750 ;
        RECT 539.030 2800.000 539.330 2801.450 ;
        RECT 538.410 2796.350 538.810 2796.650 ;
        RECT 538.510 2794.625 538.810 2796.350 ;
        RECT 542.190 2794.625 542.490 2801.450 ;
        RECT 543.110 2801.450 544.550 2801.750 ;
        RECT 535.735 2794.295 536.065 2794.625 ;
        RECT 538.495 2794.295 538.825 2794.625 ;
        RECT 542.175 2794.295 542.505 2794.625 ;
        RECT 543.110 2793.945 543.410 2801.450 ;
        RECT 544.250 2800.000 544.550 2801.450 ;
        RECT 544.870 2801.750 545.170 2804.600 ;
        RECT 984.010 2801.750 984.310 2804.600 ;
        RECT 989.850 2801.750 990.150 2804.600 ;
        RECT 995.690 2801.750 995.990 2804.600 ;
        RECT 1001.530 2801.750 1001.830 2804.600 ;
        RECT 544.870 2801.450 548.010 2801.750 ;
        RECT 544.870 2800.000 545.170 2801.450 ;
        RECT 547.710 2794.625 548.010 2801.450 ;
        RECT 981.030 2801.450 984.310 2801.750 ;
        RECT 547.695 2794.295 548.025 2794.625 ;
        RECT 981.030 2793.945 981.330 2801.450 ;
        RECT 984.010 2800.000 984.310 2801.450 ;
        RECT 987.470 2801.450 990.150 2801.750 ;
        RECT 531.135 2793.615 531.465 2793.945 ;
        RECT 543.095 2793.615 543.425 2793.945 ;
        RECT 981.015 2793.615 981.345 2793.945 ;
        RECT 987.470 2793.265 987.770 2801.450 ;
        RECT 989.850 2800.000 990.150 2801.450 ;
        RECT 993.910 2801.450 995.990 2801.750 ;
        RECT 509.055 2792.935 509.385 2793.265 ;
        RECT 987.455 2792.935 987.785 2793.265 ;
        RECT 993.910 2792.585 994.210 2801.450 ;
        RECT 995.690 2800.000 995.990 2801.450 ;
        RECT 1001.270 2800.000 1001.830 2801.750 ;
        RECT 1007.370 2802.450 1007.670 2804.600 ;
        RECT 1007.370 2802.150 1008.930 2802.450 ;
        RECT 1007.370 2800.000 1007.670 2802.150 ;
        RECT 1001.270 2792.585 1001.570 2800.000 ;
        RECT 1008.630 2793.945 1008.930 2802.150 ;
        RECT 1013.210 2801.750 1013.510 2804.600 ;
        RECT 1012.310 2801.450 1013.510 2801.750 ;
        RECT 1012.310 2793.945 1012.610 2801.450 ;
        RECT 1013.210 2800.000 1013.510 2801.450 ;
        RECT 1013.830 2796.650 1014.130 2804.600 ;
        RECT 1019.050 2801.750 1019.350 2804.600 ;
        RECT 1013.230 2796.350 1014.130 2796.650 ;
        RECT 1018.750 2800.000 1019.350 2801.750 ;
        RECT 1013.230 2794.625 1013.530 2796.350 ;
        RECT 1013.215 2794.295 1013.545 2794.625 ;
        RECT 1008.615 2793.615 1008.945 2793.945 ;
        RECT 1012.295 2793.615 1012.625 2793.945 ;
        RECT 1018.750 2793.265 1019.050 2800.000 ;
        RECT 1019.670 2794.625 1019.970 2804.600 ;
        RECT 1024.890 2801.750 1025.190 2804.600 ;
        RECT 1024.270 2801.450 1025.190 2801.750 ;
        RECT 1019.655 2794.295 1019.985 2794.625 ;
        RECT 1024.270 2793.945 1024.570 2801.450 ;
        RECT 1024.890 2800.000 1025.190 2801.450 ;
        RECT 1025.510 2801.750 1025.810 2804.600 ;
        RECT 1030.730 2801.750 1031.030 2804.600 ;
        RECT 1025.510 2801.450 1027.330 2801.750 ;
        RECT 1025.510 2800.000 1025.810 2801.450 ;
        RECT 1027.030 2794.625 1027.330 2801.450 ;
        RECT 1030.710 2800.000 1031.030 2801.750 ;
        RECT 1031.350 2801.750 1031.650 2804.600 ;
        RECT 1036.570 2802.450 1036.870 2804.600 ;
        RECT 1035.310 2802.150 1036.870 2802.450 ;
        RECT 1031.350 2801.450 1034.690 2801.750 ;
        RECT 1031.350 2800.000 1031.650 2801.450 ;
        RECT 1027.015 2794.295 1027.345 2794.625 ;
        RECT 1024.255 2793.615 1024.585 2793.945 ;
        RECT 1018.735 2792.935 1019.065 2793.265 ;
        RECT 993.895 2792.255 994.225 2792.585 ;
        RECT 1001.255 2792.255 1001.585 2792.585 ;
        RECT 1030.710 2790.545 1031.010 2800.000 ;
        RECT 1030.695 2790.215 1031.025 2790.545 ;
        RECT 1034.390 2787.825 1034.690 2801.450 ;
        RECT 1035.310 2788.505 1035.610 2802.150 ;
        RECT 1036.570 2800.000 1036.870 2802.150 ;
        RECT 1037.190 2801.750 1037.490 2804.600 ;
        RECT 1042.410 2801.750 1042.710 2804.600 ;
        RECT 1037.190 2801.450 1040.210 2801.750 ;
        RECT 1037.190 2800.000 1037.490 2801.450 ;
        RECT 1035.295 2788.175 1035.625 2788.505 ;
        RECT 1039.910 2787.825 1040.210 2801.450 ;
        RECT 1041.750 2801.450 1042.710 2801.750 ;
        RECT 1041.750 2788.505 1042.050 2801.450 ;
        RECT 1042.410 2800.000 1042.710 2801.450 ;
        RECT 1043.030 2801.750 1043.330 2804.600 ;
        RECT 1048.250 2801.750 1048.550 2804.600 ;
        RECT 1043.030 2801.450 1046.650 2801.750 ;
        RECT 1043.030 2800.000 1043.330 2801.450 ;
        RECT 1041.735 2788.175 1042.065 2788.505 ;
        RECT 1046.350 2787.825 1046.650 2801.450 ;
        RECT 1048.190 2800.000 1048.550 2801.750 ;
        RECT 1048.870 2801.750 1049.170 2804.600 ;
        RECT 1054.090 2802.450 1054.390 2804.600 ;
        RECT 1052.790 2802.150 1054.390 2802.450 ;
        RECT 1048.870 2801.450 1052.170 2801.750 ;
        RECT 1048.870 2800.000 1049.170 2801.450 ;
        RECT 1048.190 2793.265 1048.490 2800.000 ;
        RECT 1048.175 2792.935 1048.505 2793.265 ;
        RECT 1051.870 2788.505 1052.170 2801.450 ;
        RECT 1052.790 2799.385 1053.090 2802.150 ;
        RECT 1054.090 2800.000 1054.390 2802.150 ;
        RECT 1054.710 2800.050 1055.010 2804.600 ;
        RECT 1059.930 2801.750 1060.230 2804.600 ;
        RECT 1059.230 2801.450 1060.230 2801.750 ;
        RECT 1055.535 2800.050 1055.865 2800.065 ;
        RECT 1054.710 2799.750 1055.865 2800.050 ;
        RECT 1055.535 2799.735 1055.865 2799.750 ;
        RECT 1052.775 2799.055 1053.105 2799.385 ;
        RECT 1059.230 2794.625 1059.530 2801.450 ;
        RECT 1059.930 2800.000 1060.230 2801.450 ;
        RECT 1060.550 2801.750 1060.850 2804.600 ;
        RECT 1065.770 2801.750 1066.070 2804.600 ;
        RECT 1060.550 2801.450 1062.290 2801.750 ;
        RECT 1060.550 2800.000 1060.850 2801.450 ;
        RECT 1059.215 2794.295 1059.545 2794.625 ;
        RECT 1051.855 2788.175 1052.185 2788.505 ;
        RECT 1061.990 2787.825 1062.290 2801.450 ;
        RECT 1065.670 2800.000 1066.070 2801.750 ;
        RECT 1066.390 2801.750 1066.690 2804.600 ;
        RECT 1071.610 2801.750 1071.910 2804.600 ;
        RECT 1066.390 2801.450 1067.810 2801.750 ;
        RECT 1066.390 2800.000 1066.690 2801.450 ;
        RECT 1065.670 2794.625 1065.970 2800.000 ;
        RECT 1065.655 2794.295 1065.985 2794.625 ;
        RECT 1067.510 2787.825 1067.810 2801.450 ;
        RECT 1070.270 2801.450 1071.910 2801.750 ;
        RECT 1070.270 2794.625 1070.570 2801.450 ;
        RECT 1071.610 2800.000 1071.910 2801.450 ;
        RECT 1072.230 2801.750 1072.530 2804.600 ;
        RECT 1077.450 2801.750 1077.750 2804.600 ;
        RECT 1072.230 2801.450 1074.250 2801.750 ;
        RECT 1072.230 2800.000 1072.530 2801.450 ;
        RECT 1070.255 2794.295 1070.585 2794.625 ;
        RECT 1073.950 2787.825 1074.250 2801.450 ;
        RECT 1076.710 2801.450 1077.750 2801.750 ;
        RECT 1076.710 2793.945 1077.010 2801.450 ;
        RECT 1077.450 2800.000 1077.750 2801.450 ;
        RECT 1078.070 2801.750 1078.370 2804.600 ;
        RECT 1083.290 2801.750 1083.590 2804.600 ;
        RECT 1078.070 2801.450 1081.610 2801.750 ;
        RECT 1078.070 2800.000 1078.370 2801.450 ;
        RECT 1081.310 2794.625 1081.610 2801.450 ;
        RECT 1083.150 2800.000 1083.590 2801.750 ;
        RECT 1083.910 2801.750 1084.210 2804.600 ;
        RECT 1089.130 2801.750 1089.430 2804.600 ;
        RECT 1083.910 2801.450 1087.130 2801.750 ;
        RECT 1083.910 2800.000 1084.210 2801.450 ;
        RECT 1081.295 2794.295 1081.625 2794.625 ;
        RECT 1083.150 2793.945 1083.450 2800.000 ;
        RECT 1086.830 2793.945 1087.130 2801.450 ;
        RECT 1087.750 2801.450 1089.430 2801.750 ;
        RECT 1087.750 2794.625 1088.050 2801.450 ;
        RECT 1089.130 2800.000 1089.430 2801.450 ;
        RECT 1089.750 2796.650 1090.050 2804.600 ;
        RECT 1094.970 2801.750 1095.270 2804.600 ;
        RECT 1089.590 2796.350 1090.050 2796.650 ;
        RECT 1094.190 2801.450 1095.270 2801.750 ;
        RECT 1089.590 2794.625 1089.890 2796.350 ;
        RECT 1094.190 2794.625 1094.490 2801.450 ;
        RECT 1094.970 2800.000 1095.270 2801.450 ;
        RECT 1095.590 2800.050 1095.890 2804.600 ;
        RECT 1100.810 2801.750 1101.110 2804.600 ;
        RECT 1095.590 2799.750 1096.330 2800.050 ;
        RECT 1096.030 2794.625 1096.330 2799.750 ;
        RECT 1100.630 2800.000 1101.110 2801.750 ;
        RECT 1101.430 2801.750 1101.730 2804.600 ;
        RECT 1106.650 2802.450 1106.950 2804.600 ;
        RECT 1105.230 2802.150 1106.950 2802.450 ;
        RECT 1101.430 2801.450 1103.690 2801.750 ;
        RECT 1101.430 2800.000 1101.730 2801.450 ;
        RECT 1100.630 2794.625 1100.930 2800.000 ;
        RECT 1103.390 2794.625 1103.690 2801.450 ;
        RECT 1105.230 2794.625 1105.530 2802.150 ;
        RECT 1106.650 2800.000 1106.950 2802.150 ;
        RECT 1107.270 2801.750 1107.570 2804.600 ;
        RECT 1112.490 2801.750 1112.790 2804.600 ;
        RECT 1107.270 2801.450 1110.130 2801.750 ;
        RECT 1107.270 2800.000 1107.570 2801.450 ;
        RECT 1109.830 2794.625 1110.130 2801.450 ;
        RECT 1111.670 2801.450 1112.790 2801.750 ;
        RECT 1111.670 2794.625 1111.970 2801.450 ;
        RECT 1112.490 2800.000 1112.790 2801.450 ;
        RECT 1113.110 2801.750 1113.410 2804.600 ;
        RECT 1118.330 2801.750 1118.630 2804.600 ;
        RECT 1113.110 2801.450 1116.570 2801.750 ;
        RECT 1113.110 2800.000 1113.410 2801.450 ;
        RECT 1116.270 2794.625 1116.570 2801.450 ;
        RECT 1118.110 2800.000 1118.630 2801.750 ;
        RECT 1118.950 2801.750 1119.250 2804.600 ;
        RECT 1124.170 2801.750 1124.470 2804.600 ;
        RECT 1118.950 2801.450 1122.090 2801.750 ;
        RECT 1118.950 2800.000 1119.250 2801.450 ;
        RECT 1087.735 2794.295 1088.065 2794.625 ;
        RECT 1089.575 2794.295 1089.905 2794.625 ;
        RECT 1094.175 2794.295 1094.505 2794.625 ;
        RECT 1096.015 2794.295 1096.345 2794.625 ;
        RECT 1100.615 2794.295 1100.945 2794.625 ;
        RECT 1103.375 2794.295 1103.705 2794.625 ;
        RECT 1105.215 2794.295 1105.545 2794.625 ;
        RECT 1109.815 2794.295 1110.145 2794.625 ;
        RECT 1111.655 2794.295 1111.985 2794.625 ;
        RECT 1116.255 2794.295 1116.585 2794.625 ;
        RECT 1118.110 2793.945 1118.410 2800.000 ;
        RECT 1121.790 2794.625 1122.090 2801.450 ;
        RECT 1122.710 2801.450 1124.470 2801.750 ;
        RECT 1121.775 2794.295 1122.105 2794.625 ;
        RECT 1122.710 2793.945 1123.010 2801.450 ;
        RECT 1124.170 2800.000 1124.470 2801.450 ;
        RECT 1124.790 2801.750 1125.090 2804.600 ;
        RECT 1130.010 2801.750 1130.310 2804.600 ;
        RECT 1124.790 2801.450 1128.530 2801.750 ;
        RECT 1124.790 2800.000 1125.090 2801.450 ;
        RECT 1128.230 2793.945 1128.530 2801.450 ;
        RECT 1129.150 2801.450 1130.310 2801.750 ;
        RECT 1129.150 2794.625 1129.450 2801.450 ;
        RECT 1130.010 2800.000 1130.310 2801.450 ;
        RECT 1130.630 2800.050 1130.930 2804.600 ;
        RECT 1135.850 2801.750 1136.150 2804.600 ;
        RECT 1130.630 2799.750 1131.290 2800.050 ;
        RECT 1130.990 2794.625 1131.290 2799.750 ;
        RECT 1135.590 2800.000 1136.150 2801.750 ;
        RECT 1136.470 2801.750 1136.770 2804.600 ;
        RECT 1141.690 2801.750 1141.990 2804.600 ;
        RECT 1136.470 2801.450 1137.730 2801.750 ;
        RECT 1136.470 2800.000 1136.770 2801.450 ;
        RECT 1135.590 2794.625 1135.890 2800.000 ;
        RECT 1137.430 2794.625 1137.730 2801.450 ;
        RECT 1139.270 2801.450 1141.990 2801.750 ;
        RECT 1129.135 2794.295 1129.465 2794.625 ;
        RECT 1130.975 2794.295 1131.305 2794.625 ;
        RECT 1135.575 2794.295 1135.905 2794.625 ;
        RECT 1137.415 2794.295 1137.745 2794.625 ;
        RECT 1139.270 2793.945 1139.570 2801.450 ;
        RECT 1141.690 2800.000 1141.990 2801.450 ;
        RECT 1142.310 2801.750 1142.610 2804.600 ;
        RECT 1142.310 2801.450 1144.170 2801.750 ;
        RECT 1142.310 2800.000 1142.610 2801.450 ;
        RECT 1143.870 2794.625 1144.170 2801.450 ;
        RECT 1147.530 2800.050 1147.830 2804.600 ;
        RECT 1148.150 2801.750 1148.450 2804.600 ;
        RECT 1153.370 2801.750 1153.670 2804.600 ;
        RECT 1148.150 2801.450 1151.530 2801.750 ;
        RECT 1147.530 2799.750 1147.850 2800.050 ;
        RECT 1148.150 2800.000 1148.450 2801.450 ;
        RECT 1147.550 2794.625 1147.850 2799.750 ;
        RECT 1151.230 2794.625 1151.530 2801.450 ;
        RECT 1153.070 2800.000 1153.670 2801.750 ;
        RECT 1143.855 2794.295 1144.185 2794.625 ;
        RECT 1147.535 2794.295 1147.865 2794.625 ;
        RECT 1151.215 2794.295 1151.545 2794.625 ;
        RECT 1076.695 2793.615 1077.025 2793.945 ;
        RECT 1083.135 2793.615 1083.465 2793.945 ;
        RECT 1086.815 2793.615 1087.145 2793.945 ;
        RECT 1118.095 2793.615 1118.425 2793.945 ;
        RECT 1122.695 2793.615 1123.025 2793.945 ;
        RECT 1128.215 2793.615 1128.545 2793.945 ;
        RECT 1139.255 2793.615 1139.585 2793.945 ;
        RECT 1153.070 2793.265 1153.370 2800.000 ;
        RECT 1153.990 2794.625 1154.290 2804.600 ;
        RECT 1159.210 2796.650 1159.510 2804.600 ;
        RECT 1159.830 2801.750 1160.130 2804.600 ;
        RECT 1165.050 2801.750 1165.350 2804.600 ;
        RECT 1159.830 2801.450 1163.490 2801.750 ;
        RECT 1159.830 2800.000 1160.130 2801.450 ;
        RECT 1159.210 2796.350 1159.810 2796.650 ;
        RECT 1153.975 2794.295 1154.305 2794.625 ;
        RECT 1159.510 2793.265 1159.810 2796.350 ;
        RECT 1163.190 2793.945 1163.490 2801.450 ;
        RECT 1164.110 2801.450 1165.350 2801.750 ;
        RECT 1164.110 2794.625 1164.410 2801.450 ;
        RECT 1165.050 2800.000 1165.350 2801.450 ;
        RECT 1165.670 2796.650 1165.970 2804.600 ;
        RECT 1170.890 2801.750 1171.190 2804.600 ;
        RECT 1165.030 2796.350 1165.970 2796.650 ;
        RECT 1167.790 2801.450 1171.190 2801.750 ;
        RECT 1165.030 2794.625 1165.330 2796.350 ;
        RECT 1164.095 2794.295 1164.425 2794.625 ;
        RECT 1165.015 2794.295 1165.345 2794.625 ;
        RECT 1167.790 2793.945 1168.090 2801.450 ;
        RECT 1170.890 2800.000 1171.190 2801.450 ;
        RECT 1171.510 2801.750 1171.810 2804.600 ;
        RECT 1176.730 2801.750 1177.030 2804.600 ;
        RECT 1171.510 2801.450 1172.690 2801.750 ;
        RECT 1171.510 2800.000 1171.810 2801.450 ;
        RECT 1172.390 2794.625 1172.690 2801.450 ;
        RECT 1173.310 2801.450 1177.030 2801.750 ;
        RECT 1172.375 2794.295 1172.705 2794.625 ;
        RECT 1163.175 2793.615 1163.505 2793.945 ;
        RECT 1167.775 2793.615 1168.105 2793.945 ;
        RECT 1173.310 2793.265 1173.610 2801.450 ;
        RECT 1176.730 2800.000 1177.030 2801.450 ;
        RECT 1177.350 2801.750 1177.650 2804.600 ;
        RECT 1182.570 2801.750 1182.870 2804.600 ;
        RECT 1177.350 2801.450 1179.130 2801.750 ;
        RECT 1177.350 2800.000 1177.650 2801.450 ;
        RECT 1178.830 2794.625 1179.130 2801.450 ;
        RECT 1180.670 2801.450 1182.870 2801.750 ;
        RECT 1178.815 2794.295 1179.145 2794.625 ;
        RECT 1180.670 2793.945 1180.970 2801.450 ;
        RECT 1182.570 2800.000 1182.870 2801.450 ;
        RECT 1183.190 2801.750 1183.490 2804.600 ;
        RECT 1188.410 2801.750 1188.710 2804.600 ;
        RECT 1183.190 2801.450 1186.490 2801.750 ;
        RECT 1183.190 2800.000 1183.490 2801.450 ;
        RECT 1186.190 2794.625 1186.490 2801.450 ;
        RECT 1187.110 2801.450 1188.710 2801.750 ;
        RECT 1186.175 2794.295 1186.505 2794.625 ;
        RECT 1180.655 2793.615 1180.985 2793.945 ;
        RECT 1153.055 2792.935 1153.385 2793.265 ;
        RECT 1159.495 2792.935 1159.825 2793.265 ;
        RECT 1173.295 2792.935 1173.625 2793.265 ;
        RECT 1187.110 2792.585 1187.410 2801.450 ;
        RECT 1188.410 2800.000 1188.710 2801.450 ;
        RECT 1189.030 2801.750 1189.330 2804.600 ;
        RECT 1194.250 2801.750 1194.550 2804.600 ;
        RECT 1189.030 2801.450 1192.010 2801.750 ;
        RECT 1189.030 2800.000 1189.330 2801.450 ;
        RECT 1187.095 2792.255 1187.425 2792.585 ;
        RECT 1191.710 2790.545 1192.010 2801.450 ;
        RECT 1193.550 2801.450 1194.550 2801.750 ;
        RECT 1193.550 2792.585 1193.850 2801.450 ;
        RECT 1194.250 2800.000 1194.550 2801.450 ;
        RECT 1194.870 2801.750 1195.170 2804.600 ;
        RECT 1584.010 2801.750 1584.310 2804.600 ;
        RECT 1589.850 2801.750 1590.150 2804.600 ;
        RECT 1595.690 2801.750 1595.990 2804.600 ;
        RECT 1194.870 2801.450 1198.450 2801.750 ;
        RECT 1194.870 2800.000 1195.170 2801.450 ;
        RECT 1198.150 2794.625 1198.450 2801.450 ;
        RECT 1580.870 2801.450 1584.310 2801.750 ;
        RECT 1580.870 2794.625 1581.170 2801.450 ;
        RECT 1584.010 2800.000 1584.310 2801.450 ;
        RECT 1587.310 2801.450 1590.150 2801.750 ;
        RECT 1198.135 2794.295 1198.465 2794.625 ;
        RECT 1580.855 2794.295 1581.185 2794.625 ;
        RECT 1587.310 2792.585 1587.610 2801.450 ;
        RECT 1589.850 2800.000 1590.150 2801.450 ;
        RECT 1594.670 2801.450 1595.990 2801.750 ;
        RECT 1594.670 2794.625 1594.970 2801.450 ;
        RECT 1595.690 2800.000 1595.990 2801.450 ;
        RECT 1601.530 2800.050 1601.830 2804.600 ;
        RECT 1607.370 2801.750 1607.670 2804.600 ;
        RECT 1613.210 2801.750 1613.510 2804.600 ;
        RECT 1601.110 2799.750 1601.830 2800.050 ;
        RECT 1604.790 2801.450 1607.670 2801.750 ;
        RECT 1594.655 2794.295 1594.985 2794.625 ;
        RECT 1193.535 2792.255 1193.865 2792.585 ;
        RECT 1587.295 2792.255 1587.625 2792.585 ;
        RECT 1191.695 2790.215 1192.025 2790.545 ;
        RECT 1601.110 2789.185 1601.410 2799.750 ;
        RECT 1604.790 2794.625 1605.090 2801.450 ;
        RECT 1607.370 2800.000 1607.670 2801.450 ;
        RECT 1612.150 2801.450 1613.510 2801.750 ;
        RECT 1604.775 2794.295 1605.105 2794.625 ;
        RECT 1612.150 2793.945 1612.450 2801.450 ;
        RECT 1613.210 2800.000 1613.510 2801.450 ;
        RECT 1613.830 2801.750 1614.130 2804.600 ;
        RECT 1619.050 2802.450 1619.350 2804.600 ;
        RECT 1617.670 2802.150 1619.350 2802.450 ;
        RECT 1613.830 2800.000 1614.290 2801.750 ;
        RECT 1613.990 2794.625 1614.290 2800.000 ;
        RECT 1613.975 2794.295 1614.305 2794.625 ;
        RECT 1612.135 2793.615 1612.465 2793.945 ;
        RECT 1617.670 2793.265 1617.970 2802.150 ;
        RECT 1619.050 2800.000 1619.350 2802.150 ;
        RECT 1619.670 2801.750 1619.970 2804.600 ;
        RECT 1624.890 2801.750 1625.190 2804.600 ;
        RECT 1619.670 2801.450 1620.730 2801.750 ;
        RECT 1619.670 2800.000 1619.970 2801.450 ;
        RECT 1617.655 2792.935 1617.985 2793.265 ;
        RECT 1620.430 2789.865 1620.730 2801.450 ;
        RECT 1624.110 2801.450 1625.190 2801.750 ;
        RECT 1624.110 2793.265 1624.410 2801.450 ;
        RECT 1624.890 2800.000 1625.190 2801.450 ;
        RECT 1625.510 2800.050 1625.810 2804.600 ;
        RECT 1630.730 2801.750 1631.030 2804.600 ;
        RECT 1625.510 2799.750 1626.250 2800.050 ;
        RECT 1625.950 2794.625 1626.250 2799.750 ;
        RECT 1630.550 2800.000 1631.030 2801.750 ;
        RECT 1631.350 2801.750 1631.650 2804.600 ;
        RECT 1636.570 2802.450 1636.870 2804.600 ;
        RECT 1635.150 2802.150 1636.870 2802.450 ;
        RECT 1631.350 2800.000 1631.770 2801.750 ;
        RECT 1625.935 2794.295 1626.265 2794.625 ;
        RECT 1630.550 2793.265 1630.850 2800.000 ;
        RECT 1631.470 2794.625 1631.770 2800.000 ;
        RECT 1631.455 2794.295 1631.785 2794.625 ;
        RECT 1635.150 2793.945 1635.450 2802.150 ;
        RECT 1636.570 2800.000 1636.870 2802.150 ;
        RECT 1637.190 2801.750 1637.490 2804.600 ;
        RECT 1637.190 2801.450 1638.210 2801.750 ;
        RECT 1637.190 2800.000 1637.490 2801.450 ;
        RECT 1637.910 2794.625 1638.210 2801.450 ;
        RECT 1642.410 2796.650 1642.710 2804.600 ;
        RECT 1643.030 2802.450 1643.330 2804.600 ;
        RECT 1643.030 2802.150 1644.650 2802.450 ;
        RECT 1643.030 2800.000 1643.330 2802.150 ;
        RECT 1642.410 2796.350 1642.810 2796.650 ;
        RECT 1637.895 2794.295 1638.225 2794.625 ;
        RECT 1642.510 2793.945 1642.810 2796.350 ;
        RECT 1635.135 2793.615 1635.465 2793.945 ;
        RECT 1642.495 2793.615 1642.825 2793.945 ;
        RECT 1624.095 2792.935 1624.425 2793.265 ;
        RECT 1630.535 2792.935 1630.865 2793.265 ;
        RECT 1644.350 2791.225 1644.650 2802.150 ;
        RECT 1648.250 2801.750 1648.550 2804.600 ;
        RECT 1648.030 2800.000 1648.550 2801.750 ;
        RECT 1648.870 2801.750 1649.170 2804.600 ;
        RECT 1654.090 2802.450 1654.390 2804.600 ;
        RECT 1652.630 2802.150 1654.390 2802.450 ;
        RECT 1648.870 2800.000 1649.250 2801.750 ;
        RECT 1648.030 2793.265 1648.330 2800.000 ;
        RECT 1648.015 2792.935 1648.345 2793.265 ;
        RECT 1648.950 2791.905 1649.250 2800.000 ;
        RECT 1652.630 2793.265 1652.930 2802.150 ;
        RECT 1654.090 2800.000 1654.390 2802.150 ;
        RECT 1654.710 2801.750 1655.010 2804.600 ;
        RECT 1659.930 2801.750 1660.230 2804.600 ;
        RECT 1654.710 2801.450 1655.690 2801.750 ;
        RECT 1654.710 2800.000 1655.010 2801.450 ;
        RECT 1655.390 2794.625 1655.690 2801.450 ;
        RECT 1659.070 2801.450 1660.230 2801.750 ;
        RECT 1659.070 2794.625 1659.370 2801.450 ;
        RECT 1659.930 2800.000 1660.230 2801.450 ;
        RECT 1660.550 2802.450 1660.850 2804.600 ;
        RECT 1660.550 2802.150 1662.130 2802.450 ;
        RECT 1660.550 2800.000 1660.850 2802.150 ;
        RECT 1655.375 2794.295 1655.705 2794.625 ;
        RECT 1659.055 2794.295 1659.385 2794.625 ;
        RECT 1652.615 2792.935 1652.945 2793.265 ;
        RECT 1648.935 2791.575 1649.265 2791.905 ;
        RECT 1661.830 2791.225 1662.130 2802.150 ;
        RECT 1665.770 2801.750 1666.070 2804.600 ;
        RECT 1663.670 2801.450 1666.070 2801.750 ;
        RECT 1663.670 2793.945 1663.970 2801.450 ;
        RECT 1665.770 2800.000 1666.070 2801.450 ;
        RECT 1666.390 2801.750 1666.690 2804.600 ;
        RECT 1671.610 2802.450 1671.910 2804.600 ;
        RECT 1670.110 2802.150 1671.910 2802.450 ;
        RECT 1666.390 2800.000 1666.730 2801.750 ;
        RECT 1666.430 2794.625 1666.730 2800.000 ;
        RECT 1666.415 2794.295 1666.745 2794.625 ;
        RECT 1670.110 2793.945 1670.410 2802.150 ;
        RECT 1671.610 2800.000 1671.910 2802.150 ;
        RECT 1672.230 2801.750 1672.530 2804.600 ;
        RECT 1672.230 2801.450 1673.170 2801.750 ;
        RECT 1672.230 2800.000 1672.530 2801.450 ;
        RECT 1672.870 2794.625 1673.170 2801.450 ;
        RECT 1677.450 2800.050 1677.750 2804.600 ;
        RECT 1678.070 2802.450 1678.370 2804.600 ;
        RECT 1678.070 2802.150 1679.610 2802.450 ;
        RECT 1677.450 2799.750 1677.770 2800.050 ;
        RECT 1678.070 2800.000 1678.370 2802.150 ;
        RECT 1672.855 2794.295 1673.185 2794.625 ;
        RECT 1677.470 2793.945 1677.770 2799.750 ;
        RECT 1679.310 2794.625 1679.610 2802.150 ;
        RECT 1683.290 2801.750 1683.590 2804.600 ;
        RECT 1682.990 2800.000 1683.590 2801.750 ;
        RECT 1679.295 2794.295 1679.625 2794.625 ;
        RECT 1682.990 2793.945 1683.290 2800.000 ;
        RECT 1683.910 2794.625 1684.210 2804.600 ;
        RECT 1689.130 2801.750 1689.430 2804.600 ;
        RECT 1688.510 2801.450 1689.430 2801.750 ;
        RECT 1688.510 2794.625 1688.810 2801.450 ;
        RECT 1689.130 2800.000 1689.430 2801.450 ;
        RECT 1689.750 2796.650 1690.050 2804.600 ;
        RECT 1694.970 2801.750 1695.270 2804.600 ;
        RECT 1689.430 2796.350 1690.050 2796.650 ;
        RECT 1694.950 2800.000 1695.270 2801.750 ;
        RECT 1695.590 2801.750 1695.890 2804.600 ;
        RECT 1700.810 2802.450 1701.110 2804.600 ;
        RECT 1699.550 2802.150 1701.110 2802.450 ;
        RECT 1695.590 2800.000 1696.170 2801.750 ;
        RECT 1683.895 2794.295 1684.225 2794.625 ;
        RECT 1688.495 2794.295 1688.825 2794.625 ;
        RECT 1663.655 2793.615 1663.985 2793.945 ;
        RECT 1670.095 2793.615 1670.425 2793.945 ;
        RECT 1677.455 2793.615 1677.785 2793.945 ;
        RECT 1682.975 2793.615 1683.305 2793.945 ;
        RECT 1689.430 2792.585 1689.730 2796.350 ;
        RECT 1694.950 2793.945 1695.250 2800.000 ;
        RECT 1695.870 2794.625 1696.170 2800.000 ;
        RECT 1695.855 2794.295 1696.185 2794.625 ;
        RECT 1699.550 2793.945 1699.850 2802.150 ;
        RECT 1700.810 2800.000 1701.110 2802.150 ;
        RECT 1701.430 2801.750 1701.730 2804.600 ;
        RECT 1706.650 2801.750 1706.950 2804.600 ;
        RECT 1701.430 2801.450 1702.610 2801.750 ;
        RECT 1701.430 2800.000 1701.730 2801.450 ;
        RECT 1702.310 2794.625 1702.610 2801.450 ;
        RECT 1705.070 2801.450 1706.950 2801.750 ;
        RECT 1702.295 2794.295 1702.625 2794.625 ;
        RECT 1705.070 2793.945 1705.370 2801.450 ;
        RECT 1706.650 2800.000 1706.950 2801.450 ;
        RECT 1707.270 2802.450 1707.570 2804.600 ;
        RECT 1707.270 2802.150 1709.050 2802.450 ;
        RECT 1707.270 2800.000 1707.570 2802.150 ;
        RECT 1708.750 2794.625 1709.050 2802.150 ;
        RECT 1712.490 2801.750 1712.790 2804.600 ;
        RECT 1712.430 2800.000 1712.790 2801.750 ;
        RECT 1713.110 2801.750 1713.410 2804.600 ;
        RECT 1713.110 2800.000 1713.650 2801.750 ;
        RECT 1718.330 2800.050 1718.630 2804.600 ;
        RECT 1708.735 2794.295 1709.065 2794.625 ;
        RECT 1712.430 2793.945 1712.730 2800.000 ;
        RECT 1713.350 2794.625 1713.650 2800.000 ;
        RECT 1717.950 2799.750 1718.630 2800.050 ;
        RECT 1718.950 2801.750 1719.250 2804.600 ;
        RECT 1724.170 2801.750 1724.470 2804.600 ;
        RECT 1718.950 2801.450 1720.090 2801.750 ;
        RECT 1718.950 2800.000 1719.250 2801.450 ;
        RECT 1713.335 2794.295 1713.665 2794.625 ;
        RECT 1717.950 2793.945 1718.250 2799.750 ;
        RECT 1719.790 2794.625 1720.090 2801.450 ;
        RECT 1721.630 2801.450 1724.470 2801.750 ;
        RECT 1721.630 2794.625 1721.930 2801.450 ;
        RECT 1724.170 2800.000 1724.470 2801.450 ;
        RECT 1724.790 2796.650 1725.090 2804.600 ;
        RECT 1730.010 2801.750 1730.310 2804.600 ;
        RECT 1724.390 2796.350 1725.090 2796.650 ;
        RECT 1729.910 2800.000 1730.310 2801.750 ;
        RECT 1730.630 2801.750 1730.930 2804.600 ;
        RECT 1735.850 2802.450 1736.150 2804.600 ;
        RECT 1734.510 2802.150 1736.150 2802.450 ;
        RECT 1730.630 2800.000 1731.130 2801.750 ;
        RECT 1719.775 2794.295 1720.105 2794.625 ;
        RECT 1721.615 2794.295 1721.945 2794.625 ;
        RECT 1694.935 2793.615 1695.265 2793.945 ;
        RECT 1699.535 2793.615 1699.865 2793.945 ;
        RECT 1705.055 2793.615 1705.385 2793.945 ;
        RECT 1712.415 2793.615 1712.745 2793.945 ;
        RECT 1717.935 2793.615 1718.265 2793.945 ;
        RECT 1689.415 2792.255 1689.745 2792.585 ;
        RECT 1644.335 2790.895 1644.665 2791.225 ;
        RECT 1661.815 2790.895 1662.145 2791.225 ;
        RECT 1620.415 2789.535 1620.745 2789.865 ;
        RECT 1601.095 2788.855 1601.425 2789.185 ;
        RECT 1724.390 2788.505 1724.690 2796.350 ;
        RECT 1729.910 2793.945 1730.210 2800.000 ;
        RECT 1730.830 2794.625 1731.130 2800.000 ;
        RECT 1730.815 2794.295 1731.145 2794.625 ;
        RECT 1734.510 2793.945 1734.810 2802.150 ;
        RECT 1735.850 2800.000 1736.150 2802.150 ;
        RECT 1736.470 2801.750 1736.770 2804.600 ;
        RECT 1741.690 2801.750 1741.990 2804.600 ;
        RECT 1736.470 2801.450 1737.570 2801.750 ;
        RECT 1736.470 2800.000 1736.770 2801.450 ;
        RECT 1737.270 2794.625 1737.570 2801.450 ;
        RECT 1740.950 2801.450 1741.990 2801.750 ;
        RECT 1737.255 2794.295 1737.585 2794.625 ;
        RECT 1740.950 2793.945 1741.250 2801.450 ;
        RECT 1741.690 2800.000 1741.990 2801.450 ;
        RECT 1742.310 2802.450 1742.610 2804.600 ;
        RECT 1742.310 2802.150 1744.010 2802.450 ;
        RECT 1742.310 2800.000 1742.610 2802.150 ;
        RECT 1743.710 2794.625 1744.010 2802.150 ;
        RECT 1747.530 2801.750 1747.830 2804.600 ;
        RECT 1747.390 2800.000 1747.830 2801.750 ;
        RECT 1748.150 2801.750 1748.450 2804.600 ;
        RECT 1748.150 2800.000 1748.610 2801.750 ;
        RECT 1753.370 2800.050 1753.670 2804.600 ;
        RECT 1743.695 2794.295 1744.025 2794.625 ;
        RECT 1747.390 2793.945 1747.690 2800.000 ;
        RECT 1748.310 2794.625 1748.610 2800.000 ;
        RECT 1752.910 2799.750 1753.670 2800.050 ;
        RECT 1753.990 2801.750 1754.290 2804.600 ;
        RECT 1753.990 2801.450 1755.050 2801.750 ;
        RECT 1753.990 2800.000 1754.290 2801.450 ;
        RECT 1748.295 2794.295 1748.625 2794.625 ;
        RECT 1729.895 2793.615 1730.225 2793.945 ;
        RECT 1734.495 2793.615 1734.825 2793.945 ;
        RECT 1740.935 2793.615 1741.265 2793.945 ;
        RECT 1747.375 2793.615 1747.705 2793.945 ;
        RECT 1752.910 2792.585 1753.210 2799.750 ;
        RECT 1752.895 2792.255 1753.225 2792.585 ;
        RECT 1724.375 2788.175 1724.705 2788.505 ;
        RECT 1754.750 2787.825 1755.050 2801.450 ;
        RECT 1759.210 2796.665 1759.510 2804.600 ;
        RECT 1759.830 2802.450 1760.130 2804.600 ;
        RECT 1759.830 2802.150 1761.490 2802.450 ;
        RECT 1759.830 2800.000 1760.130 2802.150 ;
        RECT 1759.210 2796.350 1759.665 2796.665 ;
        RECT 1759.335 2796.335 1759.665 2796.350 ;
        RECT 357.255 2787.495 357.585 2787.825 ;
        RECT 454.775 2787.495 455.105 2787.825 ;
        RECT 460.295 2787.495 460.625 2787.825 ;
        RECT 468.575 2787.495 468.905 2787.825 ;
        RECT 475.015 2787.495 475.345 2787.825 ;
        RECT 482.375 2787.495 482.705 2787.825 ;
        RECT 488.815 2787.495 489.145 2787.825 ;
        RECT 495.255 2787.495 495.585 2787.825 ;
        RECT 1034.375 2787.495 1034.705 2787.825 ;
        RECT 1039.895 2787.495 1040.225 2787.825 ;
        RECT 1046.335 2787.495 1046.665 2787.825 ;
        RECT 1061.975 2787.495 1062.305 2787.825 ;
        RECT 1067.495 2787.495 1067.825 2787.825 ;
        RECT 1073.935 2787.495 1074.265 2787.825 ;
        RECT 1754.735 2787.495 1755.065 2787.825 ;
        RECT 292.020 2715.000 295.020 2785.000 ;
        RECT 310.020 2715.000 313.020 2785.000 ;
        RECT 328.020 2715.000 331.020 2785.000 ;
        RECT 364.020 2715.000 367.020 2785.000 ;
        RECT 454.020 2715.000 457.020 2785.000 ;
        RECT 472.020 2715.000 475.020 2785.000 ;
        RECT 490.020 2715.000 493.020 2785.000 ;
        RECT 508.020 2715.000 511.020 2785.000 ;
        RECT 544.020 2715.000 547.020 2785.000 ;
        RECT 634.020 2715.000 637.020 2785.000 ;
        RECT 652.020 2715.000 655.020 2785.000 ;
        RECT 670.020 2715.000 673.020 2785.000 ;
        RECT 688.020 2715.000 691.020 2785.000 ;
        RECT 994.020 2715.000 997.020 2785.000 ;
        RECT 1012.020 2715.000 1015.020 2785.000 ;
        RECT 1030.020 2715.000 1033.020 2785.000 ;
        RECT 1048.020 2715.000 1051.020 2785.000 ;
        RECT 1084.020 2715.000 1087.020 2785.000 ;
        RECT 1174.020 2715.000 1177.020 2785.000 ;
        RECT 1192.020 2715.000 1195.020 2785.000 ;
        RECT 1210.020 2715.000 1213.020 2785.000 ;
        RECT 1228.020 2715.000 1231.020 2785.000 ;
        RECT 1264.020 2715.000 1267.020 2785.000 ;
        RECT 1761.190 2777.625 1761.490 2802.150 ;
        RECT 1765.050 2801.750 1765.350 2804.600 ;
        RECT 1762.110 2801.450 1765.350 2801.750 ;
        RECT 1762.110 2794.625 1762.410 2801.450 ;
        RECT 1765.050 2800.000 1765.350 2801.450 ;
        RECT 1765.670 2801.750 1765.970 2804.600 ;
        RECT 1770.890 2801.750 1771.190 2804.600 ;
        RECT 1765.670 2800.000 1766.090 2801.750 ;
        RECT 1762.095 2794.295 1762.425 2794.625 ;
        RECT 1765.790 2788.505 1766.090 2800.000 ;
        RECT 1767.630 2801.450 1771.190 2801.750 ;
        RECT 1767.630 2793.945 1767.930 2801.450 ;
        RECT 1770.890 2800.000 1771.190 2801.450 ;
        RECT 1771.510 2801.750 1771.810 2804.600 ;
        RECT 1776.730 2801.750 1777.030 2804.600 ;
        RECT 1771.510 2801.450 1772.530 2801.750 ;
        RECT 1771.510 2800.000 1771.810 2801.450 ;
        RECT 1767.615 2793.615 1767.945 2793.945 ;
        RECT 1765.775 2788.175 1766.105 2788.505 ;
        RECT 1772.230 2787.825 1772.530 2801.450 ;
        RECT 1774.070 2801.450 1777.030 2801.750 ;
        RECT 1774.070 2791.905 1774.370 2801.450 ;
        RECT 1776.730 2800.000 1777.030 2801.450 ;
        RECT 1777.350 2800.050 1777.650 2804.600 ;
        RECT 1782.570 2801.750 1782.870 2804.600 ;
        RECT 1780.510 2801.450 1782.870 2801.750 ;
        RECT 1777.350 2799.750 1778.050 2800.050 ;
        RECT 1774.055 2791.575 1774.385 2791.905 ;
        RECT 1777.750 2787.825 1778.050 2799.750 ;
        RECT 1780.510 2793.265 1780.810 2801.450 ;
        RECT 1782.570 2800.000 1782.870 2801.450 ;
        RECT 1783.190 2801.750 1783.490 2804.600 ;
        RECT 1783.190 2800.000 1783.570 2801.750 ;
        RECT 1788.410 2800.050 1788.710 2804.600 ;
        RECT 1780.495 2792.935 1780.825 2793.265 ;
        RECT 1783.270 2787.825 1783.570 2800.000 ;
        RECT 1787.870 2799.750 1788.710 2800.050 ;
        RECT 1789.030 2801.750 1789.330 2804.600 ;
        RECT 1789.030 2801.450 1790.010 2801.750 ;
        RECT 1789.030 2800.000 1789.330 2801.450 ;
        RECT 1787.870 2793.945 1788.170 2799.750 ;
        RECT 1787.855 2793.615 1788.185 2793.945 ;
        RECT 1789.710 2787.825 1790.010 2801.450 ;
        RECT 1794.250 2796.665 1794.550 2804.600 ;
        RECT 1794.870 2802.450 1795.170 2804.600 ;
        RECT 1794.870 2802.150 1796.450 2802.450 ;
        RECT 1794.870 2800.000 1795.170 2802.150 ;
        RECT 1794.250 2796.350 1794.625 2796.665 ;
        RECT 1794.295 2796.335 1794.625 2796.350 ;
        RECT 1772.215 2787.495 1772.545 2787.825 ;
        RECT 1777.735 2787.495 1778.065 2787.825 ;
        RECT 1783.255 2787.495 1783.585 2787.825 ;
        RECT 1789.695 2787.495 1790.025 2787.825 ;
        RECT 1796.150 2777.625 1796.450 2802.150 ;
        RECT 2234.010 2801.750 2234.310 2804.600 ;
        RECT 2239.850 2801.750 2240.150 2804.600 ;
        RECT 2245.690 2801.750 2245.990 2804.600 ;
        RECT 2251.530 2801.750 2251.830 2804.600 ;
        RECT 2257.370 2801.750 2257.670 2804.600 ;
        RECT 2231.310 2801.450 2234.310 2801.750 ;
        RECT 2231.310 2794.625 2231.610 2801.450 ;
        RECT 2234.010 2800.000 2234.310 2801.450 ;
        RECT 2236.830 2801.450 2240.150 2801.750 ;
        RECT 2236.830 2794.625 2237.130 2801.450 ;
        RECT 2239.850 2800.000 2240.150 2801.450 ;
        RECT 2242.350 2801.450 2245.990 2801.750 ;
        RECT 2242.350 2794.625 2242.650 2801.450 ;
        RECT 2245.690 2800.000 2245.990 2801.450 ;
        RECT 2249.710 2801.450 2251.830 2801.750 ;
        RECT 2249.710 2794.625 2250.010 2801.450 ;
        RECT 2251.530 2800.000 2251.830 2801.450 ;
        RECT 2257.070 2800.000 2257.670 2801.750 ;
        RECT 2231.295 2794.295 2231.625 2794.625 ;
        RECT 2236.815 2794.295 2237.145 2794.625 ;
        RECT 2242.335 2794.295 2242.665 2794.625 ;
        RECT 2249.695 2794.295 2250.025 2794.625 ;
        RECT 2257.070 2788.505 2257.370 2800.000 ;
        RECT 2263.210 2796.650 2263.510 2804.600 ;
        RECT 2263.830 2801.750 2264.130 2804.600 ;
        RECT 2269.050 2801.750 2269.350 2804.600 ;
        RECT 2263.830 2801.450 2264.730 2801.750 ;
        RECT 2263.830 2800.000 2264.130 2801.450 ;
        RECT 2263.210 2796.350 2263.810 2796.650 ;
        RECT 2263.510 2793.945 2263.810 2796.350 ;
        RECT 2264.430 2794.625 2264.730 2801.450 ;
        RECT 2268.110 2801.450 2269.350 2801.750 ;
        RECT 2268.110 2794.625 2268.410 2801.450 ;
        RECT 2269.050 2800.000 2269.350 2801.450 ;
        RECT 2269.670 2796.650 2269.970 2804.600 ;
        RECT 2274.890 2802.450 2275.190 2804.600 ;
        RECT 2269.030 2796.350 2269.970 2796.650 ;
        RECT 2273.630 2802.150 2275.190 2802.450 ;
        RECT 2264.415 2794.295 2264.745 2794.625 ;
        RECT 2268.095 2794.295 2268.425 2794.625 ;
        RECT 2263.495 2793.615 2263.825 2793.945 ;
        RECT 2269.030 2791.225 2269.330 2796.350 ;
        RECT 2273.630 2794.625 2273.930 2802.150 ;
        RECT 2274.890 2800.000 2275.190 2802.150 ;
        RECT 2275.510 2801.750 2275.810 2804.600 ;
        RECT 2280.730 2801.750 2281.030 2804.600 ;
        RECT 2275.510 2801.450 2276.690 2801.750 ;
        RECT 2275.510 2800.000 2275.810 2801.450 ;
        RECT 2273.615 2794.295 2273.945 2794.625 ;
        RECT 2276.390 2791.905 2276.690 2801.450 ;
        RECT 2280.070 2801.450 2281.030 2801.750 ;
        RECT 2280.070 2793.265 2280.370 2801.450 ;
        RECT 2280.730 2800.000 2281.030 2801.450 ;
        RECT 2281.350 2802.450 2281.650 2804.600 ;
        RECT 2281.350 2802.150 2283.130 2802.450 ;
        RECT 2281.350 2800.000 2281.650 2802.150 ;
        RECT 2280.055 2792.935 2280.385 2793.265 ;
        RECT 2282.830 2792.585 2283.130 2802.150 ;
        RECT 2286.570 2801.750 2286.870 2804.600 ;
        RECT 2286.510 2800.000 2286.870 2801.750 ;
        RECT 2287.190 2801.750 2287.490 2804.600 ;
        RECT 2287.190 2800.000 2287.730 2801.750 ;
        RECT 2292.410 2800.050 2292.710 2804.600 ;
        RECT 2286.510 2793.265 2286.810 2800.000 ;
        RECT 2286.495 2792.935 2286.825 2793.265 ;
        RECT 2282.815 2792.255 2283.145 2792.585 ;
        RECT 2287.430 2791.905 2287.730 2800.000 ;
        RECT 2292.030 2799.750 2292.710 2800.050 ;
        RECT 2293.030 2801.750 2293.330 2804.600 ;
        RECT 2298.250 2801.750 2298.550 2804.600 ;
        RECT 2293.030 2801.450 2294.170 2801.750 ;
        RECT 2293.030 2800.000 2293.330 2801.450 ;
        RECT 2292.030 2794.625 2292.330 2799.750 ;
        RECT 2292.015 2794.295 2292.345 2794.625 ;
        RECT 2293.870 2791.905 2294.170 2801.450 ;
        RECT 2297.550 2801.450 2298.550 2801.750 ;
        RECT 2297.550 2793.945 2297.850 2801.450 ;
        RECT 2298.250 2800.000 2298.550 2801.450 ;
        RECT 2298.870 2800.050 2299.170 2804.600 ;
        RECT 2304.090 2801.750 2304.390 2804.600 ;
        RECT 2298.870 2799.750 2299.690 2800.050 ;
        RECT 2297.535 2793.615 2297.865 2793.945 ;
        RECT 2276.375 2791.575 2276.705 2791.905 ;
        RECT 2287.415 2791.575 2287.745 2791.905 ;
        RECT 2293.855 2791.575 2294.185 2791.905 ;
        RECT 2299.390 2791.225 2299.690 2799.750 ;
        RECT 2303.990 2800.000 2304.390 2801.750 ;
        RECT 2304.710 2801.750 2305.010 2804.600 ;
        RECT 2309.930 2802.450 2310.230 2804.600 ;
        RECT 2308.590 2802.150 2310.230 2802.450 ;
        RECT 2304.710 2800.000 2305.210 2801.750 ;
        RECT 2303.990 2793.265 2304.290 2800.000 ;
        RECT 2304.910 2794.625 2305.210 2800.000 ;
        RECT 2308.590 2794.625 2308.890 2802.150 ;
        RECT 2309.930 2800.000 2310.230 2802.150 ;
        RECT 2310.550 2796.650 2310.850 2804.600 ;
        RECT 2315.770 2801.750 2316.070 2804.600 ;
        RECT 2310.430 2796.350 2310.850 2796.650 ;
        RECT 2315.030 2801.450 2316.070 2801.750 ;
        RECT 2304.895 2794.295 2305.225 2794.625 ;
        RECT 2308.575 2794.295 2308.905 2794.625 ;
        RECT 2310.430 2793.945 2310.730 2796.350 ;
        RECT 2315.030 2793.945 2315.330 2801.450 ;
        RECT 2315.770 2800.000 2316.070 2801.450 ;
        RECT 2316.390 2800.050 2316.690 2804.600 ;
        RECT 2321.610 2801.750 2321.910 2804.600 ;
        RECT 2316.390 2799.750 2317.170 2800.050 ;
        RECT 2316.870 2794.625 2317.170 2799.750 ;
        RECT 2321.470 2800.000 2321.910 2801.750 ;
        RECT 2322.230 2801.750 2322.530 2804.600 ;
        RECT 2327.450 2802.450 2327.750 2804.600 ;
        RECT 2326.070 2802.150 2327.750 2802.450 ;
        RECT 2322.230 2800.000 2322.690 2801.750 ;
        RECT 2316.855 2794.295 2317.185 2794.625 ;
        RECT 2321.470 2793.945 2321.770 2800.000 ;
        RECT 2322.390 2794.625 2322.690 2800.000 ;
        RECT 2322.375 2794.295 2322.705 2794.625 ;
        RECT 2326.070 2793.945 2326.370 2802.150 ;
        RECT 2327.450 2800.000 2327.750 2802.150 ;
        RECT 2328.070 2801.750 2328.370 2804.600 ;
        RECT 2333.290 2801.750 2333.590 2804.600 ;
        RECT 2328.070 2801.450 2329.130 2801.750 ;
        RECT 2328.070 2800.000 2328.370 2801.450 ;
        RECT 2328.830 2794.625 2329.130 2801.450 ;
        RECT 2332.510 2801.450 2333.590 2801.750 ;
        RECT 2328.815 2794.295 2329.145 2794.625 ;
        RECT 2310.415 2793.615 2310.745 2793.945 ;
        RECT 2315.015 2793.615 2315.345 2793.945 ;
        RECT 2321.455 2793.615 2321.785 2793.945 ;
        RECT 2326.055 2793.615 2326.385 2793.945 ;
        RECT 2332.510 2793.265 2332.810 2801.450 ;
        RECT 2333.290 2800.000 2333.590 2801.450 ;
        RECT 2333.910 2800.050 2334.210 2804.600 ;
        RECT 2339.130 2801.750 2339.430 2804.600 ;
        RECT 2333.910 2799.750 2334.650 2800.050 ;
        RECT 2334.350 2794.625 2334.650 2799.750 ;
        RECT 2338.950 2800.000 2339.430 2801.750 ;
        RECT 2339.750 2801.750 2340.050 2804.600 ;
        RECT 2344.970 2801.750 2345.270 2804.600 ;
        RECT 2339.750 2800.000 2340.170 2801.750 ;
        RECT 2334.335 2794.295 2334.665 2794.625 ;
        RECT 2338.950 2793.265 2339.250 2800.000 ;
        RECT 2339.870 2794.625 2340.170 2800.000 ;
        RECT 2343.550 2801.450 2345.270 2801.750 ;
        RECT 2343.550 2794.625 2343.850 2801.450 ;
        RECT 2344.970 2800.000 2345.270 2801.450 ;
        RECT 2345.590 2796.650 2345.890 2804.600 ;
        RECT 2350.810 2801.750 2351.110 2804.600 ;
        RECT 2345.390 2796.350 2345.890 2796.650 ;
        RECT 2349.990 2801.450 2351.110 2801.750 ;
        RECT 2339.855 2794.295 2340.185 2794.625 ;
        RECT 2343.535 2794.295 2343.865 2794.625 ;
        RECT 2345.390 2793.945 2345.690 2796.350 ;
        RECT 2349.990 2793.945 2350.290 2801.450 ;
        RECT 2350.810 2800.000 2351.110 2801.450 ;
        RECT 2351.430 2800.050 2351.730 2804.600 ;
        RECT 2356.650 2801.750 2356.950 2804.600 ;
        RECT 2351.430 2799.750 2352.130 2800.050 ;
        RECT 2351.830 2794.625 2352.130 2799.750 ;
        RECT 2356.430 2800.000 2356.950 2801.750 ;
        RECT 2357.270 2801.750 2357.570 2804.600 ;
        RECT 2362.490 2802.450 2362.790 2804.600 ;
        RECT 2361.030 2802.150 2362.790 2802.450 ;
        RECT 2357.270 2800.000 2357.650 2801.750 ;
        RECT 2351.815 2794.295 2352.145 2794.625 ;
        RECT 2356.430 2793.945 2356.730 2800.000 ;
        RECT 2357.350 2794.625 2357.650 2800.000 ;
        RECT 2357.335 2794.295 2357.665 2794.625 ;
        RECT 2361.030 2793.945 2361.330 2802.150 ;
        RECT 2362.490 2800.000 2362.790 2802.150 ;
        RECT 2363.110 2801.750 2363.410 2804.600 ;
        RECT 2368.330 2801.750 2368.630 2804.600 ;
        RECT 2363.110 2801.450 2364.090 2801.750 ;
        RECT 2363.110 2800.000 2363.410 2801.450 ;
        RECT 2363.790 2794.625 2364.090 2801.450 ;
        RECT 2367.470 2801.450 2368.630 2801.750 ;
        RECT 2363.775 2794.295 2364.105 2794.625 ;
        RECT 2367.470 2793.945 2367.770 2801.450 ;
        RECT 2368.330 2800.000 2368.630 2801.450 ;
        RECT 2368.950 2802.450 2369.250 2804.600 ;
        RECT 2368.950 2802.150 2370.530 2802.450 ;
        RECT 2368.950 2800.000 2369.250 2802.150 ;
        RECT 2370.230 2794.625 2370.530 2802.150 ;
        RECT 2374.170 2801.750 2374.470 2804.600 ;
        RECT 2373.910 2800.000 2374.470 2801.750 ;
        RECT 2374.790 2801.750 2375.090 2804.600 ;
        RECT 2380.010 2801.750 2380.310 2804.600 ;
        RECT 2374.790 2800.000 2375.130 2801.750 ;
        RECT 2370.215 2794.295 2370.545 2794.625 ;
        RECT 2373.910 2793.945 2374.210 2800.000 ;
        RECT 2374.830 2794.625 2375.130 2800.000 ;
        RECT 2377.590 2801.450 2380.310 2801.750 ;
        RECT 2374.815 2794.295 2375.145 2794.625 ;
        RECT 2377.590 2793.945 2377.890 2801.450 ;
        RECT 2380.010 2800.000 2380.310 2801.450 ;
        RECT 2380.630 2801.750 2380.930 2804.600 ;
        RECT 2380.630 2801.450 2381.570 2801.750 ;
        RECT 2380.630 2800.000 2380.930 2801.450 ;
        RECT 2381.270 2794.625 2381.570 2801.450 ;
        RECT 2385.850 2800.050 2386.150 2804.600 ;
        RECT 2386.470 2800.050 2386.770 2804.600 ;
        RECT 2391.690 2801.750 2391.990 2804.600 ;
        RECT 2385.850 2799.750 2386.170 2800.050 ;
        RECT 2386.470 2799.750 2387.090 2800.050 ;
        RECT 2385.870 2794.625 2386.170 2799.750 ;
        RECT 2381.255 2794.295 2381.585 2794.625 ;
        RECT 2385.855 2794.295 2386.185 2794.625 ;
        RECT 2345.375 2793.615 2345.705 2793.945 ;
        RECT 2349.975 2793.615 2350.305 2793.945 ;
        RECT 2356.415 2793.615 2356.745 2793.945 ;
        RECT 2361.015 2793.615 2361.345 2793.945 ;
        RECT 2367.455 2793.615 2367.785 2793.945 ;
        RECT 2373.895 2793.615 2374.225 2793.945 ;
        RECT 2377.575 2793.615 2377.905 2793.945 ;
        RECT 2303.975 2792.935 2304.305 2793.265 ;
        RECT 2332.495 2792.935 2332.825 2793.265 ;
        RECT 2338.935 2792.935 2339.265 2793.265 ;
        RECT 2269.015 2790.895 2269.345 2791.225 ;
        RECT 2299.375 2790.895 2299.705 2791.225 ;
        RECT 2377.590 2788.505 2377.890 2793.615 ;
        RECT 2386.790 2790.545 2387.090 2799.750 ;
        RECT 2391.390 2800.000 2391.990 2801.750 ;
        RECT 2391.390 2794.625 2391.690 2800.000 ;
        RECT 2391.375 2794.295 2391.705 2794.625 ;
        RECT 2392.310 2790.545 2392.610 2804.600 ;
        RECT 2397.530 2801.750 2397.830 2804.600 ;
        RECT 2396.910 2801.450 2397.830 2801.750 ;
        RECT 2396.910 2794.625 2397.210 2801.450 ;
        RECT 2397.530 2800.000 2397.830 2801.450 ;
        RECT 2398.150 2801.750 2398.450 2804.600 ;
        RECT 2403.370 2801.750 2403.670 2804.600 ;
        RECT 2398.150 2801.450 2399.050 2801.750 ;
        RECT 2398.150 2800.000 2398.450 2801.450 ;
        RECT 2396.895 2794.295 2397.225 2794.625 ;
        RECT 2386.775 2790.215 2387.105 2790.545 ;
        RECT 2392.295 2790.215 2392.625 2790.545 ;
        RECT 2398.750 2789.865 2399.050 2801.450 ;
        RECT 2402.430 2801.450 2403.670 2801.750 ;
        RECT 2402.430 2793.945 2402.730 2801.450 ;
        RECT 2403.370 2800.000 2403.670 2801.450 ;
        RECT 2403.990 2801.750 2404.290 2804.600 ;
        RECT 2409.210 2802.450 2409.510 2804.600 ;
        RECT 2407.950 2802.150 2409.510 2802.450 ;
        RECT 2403.990 2800.000 2404.570 2801.750 ;
        RECT 2404.270 2794.625 2404.570 2800.000 ;
        RECT 2404.255 2794.295 2404.585 2794.625 ;
        RECT 2402.415 2793.615 2402.745 2793.945 ;
        RECT 2407.950 2792.585 2408.250 2802.150 ;
        RECT 2409.210 2800.000 2409.510 2802.150 ;
        RECT 2409.830 2801.750 2410.130 2804.600 ;
        RECT 2409.830 2801.450 2411.010 2801.750 ;
        RECT 2409.830 2800.000 2410.130 2801.450 ;
        RECT 2407.935 2792.255 2408.265 2792.585 ;
        RECT 2398.735 2789.535 2399.065 2789.865 ;
        RECT 2410.710 2789.185 2411.010 2801.450 ;
        RECT 2415.050 2796.650 2415.350 2804.600 ;
        RECT 2415.670 2802.450 2415.970 2804.600 ;
        RECT 2415.670 2802.150 2417.450 2802.450 ;
        RECT 2415.670 2800.000 2415.970 2802.150 ;
        RECT 2415.050 2796.350 2415.610 2796.650 ;
        RECT 2415.310 2793.265 2415.610 2796.350 ;
        RECT 2417.150 2794.625 2417.450 2802.150 ;
        RECT 2420.890 2801.750 2421.190 2804.600 ;
        RECT 2418.070 2801.450 2421.190 2801.750 ;
        RECT 2417.135 2794.295 2417.465 2794.625 ;
        RECT 2415.295 2792.935 2415.625 2793.265 ;
        RECT 2410.695 2788.855 2411.025 2789.185 ;
        RECT 2418.070 2788.505 2418.370 2801.450 ;
        RECT 2420.890 2800.000 2421.190 2801.450 ;
        RECT 2421.510 2796.650 2421.810 2804.600 ;
        RECT 2426.730 2801.750 2427.030 2804.600 ;
        RECT 2420.830 2796.350 2421.810 2796.650 ;
        RECT 2423.590 2801.450 2427.030 2801.750 ;
        RECT 2420.830 2791.225 2421.130 2796.350 ;
        RECT 2423.590 2793.945 2423.890 2801.450 ;
        RECT 2426.730 2800.000 2427.030 2801.450 ;
        RECT 2427.350 2801.750 2427.650 2804.600 ;
        RECT 2432.570 2801.750 2432.870 2804.600 ;
        RECT 2427.350 2801.450 2428.490 2801.750 ;
        RECT 2427.350 2800.000 2427.650 2801.450 ;
        RECT 2428.190 2794.625 2428.490 2801.450 ;
        RECT 2430.030 2801.450 2432.870 2801.750 ;
        RECT 2430.030 2794.625 2430.330 2801.450 ;
        RECT 2432.570 2800.000 2432.870 2801.450 ;
        RECT 2433.190 2802.450 2433.490 2804.600 ;
        RECT 2433.190 2802.150 2434.930 2802.450 ;
        RECT 2433.190 2800.000 2433.490 2802.150 ;
        RECT 2428.175 2794.295 2428.505 2794.625 ;
        RECT 2430.015 2794.295 2430.345 2794.625 ;
        RECT 2423.575 2793.615 2423.905 2793.945 ;
        RECT 2434.630 2791.225 2434.930 2802.150 ;
        RECT 2438.410 2801.750 2438.710 2804.600 ;
        RECT 2436.470 2801.450 2438.710 2801.750 ;
        RECT 2436.470 2792.585 2436.770 2801.450 ;
        RECT 2438.410 2800.000 2438.710 2801.450 ;
        RECT 2439.030 2801.750 2439.330 2804.600 ;
        RECT 2444.250 2801.750 2444.550 2804.600 ;
        RECT 2439.030 2800.000 2439.530 2801.750 ;
        RECT 2436.455 2792.255 2436.785 2792.585 ;
        RECT 2439.230 2791.225 2439.530 2800.000 ;
        RECT 2442.910 2801.450 2444.550 2801.750 ;
        RECT 2442.910 2793.265 2443.210 2801.450 ;
        RECT 2444.250 2800.000 2444.550 2801.450 ;
        RECT 2444.870 2801.750 2445.170 2804.600 ;
        RECT 2444.870 2801.450 2445.970 2801.750 ;
        RECT 2444.870 2800.000 2445.170 2801.450 ;
        RECT 2442.895 2792.935 2443.225 2793.265 ;
        RECT 2445.670 2791.905 2445.970 2801.450 ;
        RECT 2445.655 2791.575 2445.985 2791.905 ;
        RECT 2420.815 2790.895 2421.145 2791.225 ;
        RECT 2434.615 2790.895 2434.945 2791.225 ;
        RECT 2439.215 2790.895 2439.545 2791.225 ;
        RECT 2257.055 2788.175 2257.385 2788.505 ;
        RECT 2377.575 2788.175 2377.905 2788.505 ;
        RECT 2418.055 2788.175 2418.385 2788.505 ;
        RECT 1761.175 2777.295 1761.505 2777.625 ;
        RECT 1796.135 2777.295 1796.465 2777.625 ;
      LAYER met4 ;
        RECT 314.095 1510.640 320.640 2688.880 ;
        RECT 323.040 1510.640 397.440 2688.880 ;
        RECT 399.840 1510.640 1388.065 2688.880 ;
  END
END user_project_wrapper
END LIBRARY

