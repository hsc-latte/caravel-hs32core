magic
tech sky130A
magscale 1 2
timestamp 1608421104
<< locali >>
rect 260849 652783 260883 653361
rect 318809 650675 318843 650777
rect 280169 650539 280203 650641
rect 193229 650335 193263 650505
rect 202797 650403 202831 650505
rect 212549 650335 212583 650505
rect 222117 650403 222151 650505
rect 231869 650335 231903 650505
rect 241437 650403 241471 650505
rect 251189 650335 251223 650505
rect 260757 650403 260791 650505
rect 289737 650471 289771 650641
rect 328377 650607 328411 650777
rect 338129 650675 338163 650777
rect 347697 650607 347731 650777
rect 357449 650675 357483 650777
rect 367017 650607 367051 650777
rect 434729 650675 434763 650777
rect 311851 650573 311909 650607
rect 331171 650573 331229 650607
rect 350491 650573 350549 650607
rect 369903 650573 369961 650607
rect 273211 650437 273269 650471
rect 292531 650437 292589 650471
rect 405749 650199 405783 650505
rect 425069 650335 425103 650641
rect 444297 650607 444331 650777
rect 454049 650675 454083 650777
rect 463617 650607 463651 650777
rect 473369 650675 473403 650777
rect 482937 650607 482971 650777
rect 492689 650675 492723 650777
rect 502257 650607 502291 650777
rect 447091 650573 447149 650607
rect 466411 650573 466469 650607
rect 485731 650573 485789 650607
rect 505143 650573 505201 650607
rect 101965 558705 102885 558739
rect 101965 558671 101999 558705
rect 93869 557923 93903 558433
rect 97273 557923 97307 558637
rect 97123 557889 97307 557923
rect 99757 557923 99791 558637
rect 99849 557923 99883 558569
rect 208593 557923 208627 558365
rect 222209 557923 222243 558093
rect 231777 557923 231811 558025
rect 325709 557855 325743 558365
rect 93995 557821 94915 557855
rect 94881 557719 94915 557821
rect 98285 557719 98319 557821
rect 106289 557515 106323 557821
rect 115857 557515 115891 557753
rect 125425 557515 125459 557821
rect 128311 557549 128369 557583
rect 125609 556903 125643 557481
rect 145481 542487 145515 543677
rect 152381 542419 152415 543541
rect 152473 542555 152507 543677
rect 216781 542963 216815 543201
rect 281641 413899 281675 421345
rect 282101 417639 282135 431545
rect 384589 413831 384623 414001
rect 373917 412743 373951 412981
rect 375941 412947 375975 413457
rect 377413 413015 377447 413185
rect 377505 412743 377539 413185
rect 378609 413151 378643 413389
rect 378885 413219 378919 413389
rect 378735 413185 378919 413219
rect 381369 413015 381403 413593
rect 377355 412709 377539 412743
rect 384221 412607 384255 412913
rect 384313 412743 384347 413321
rect 384405 412743 384439 413389
rect 384497 413151 384531 413797
rect 386521 413627 386555 413797
rect 384589 413083 384623 413389
rect 387901 412675 387935 412981
rect 387993 412675 388027 413593
rect 282193 386427 282227 395981
rect 282285 367183 282319 369869
rect 282101 357459 282135 366877
rect 282377 328491 282411 338045
rect 97767 318597 98101 318631
rect 131037 317543 131071 318733
rect 131313 4913 131865 4947
rect 130117 4811 130151 4845
rect 131313 4811 131347 4913
rect 130117 4777 130485 4811
rect 55229 4131 55263 4505
rect 64797 4131 64831 4505
rect 16589 3995 16623 4097
rect 35909 3451 35943 3553
rect 80069 3383 80103 4029
rect 84853 3927 84887 4097
rect 6837 2907 6871 3145
rect 55229 2703 55263 3349
rect 58541 2839 58575 3349
rect 64797 2975 64831 3349
rect 69673 3179 69707 3281
rect 91293 3247 91327 3893
rect 108313 3859 108347 4029
rect 95617 3723 95651 3825
rect 68327 3077 68477 3111
rect 63509 2941 63785 2975
rect 63509 2839 63543 2941
<< viali >>
rect 260849 653361 260883 653395
rect 260849 652749 260883 652783
rect 318809 650777 318843 650811
rect 280169 650641 280203 650675
rect 193229 650505 193263 650539
rect 202797 650505 202831 650539
rect 202797 650369 202831 650403
rect 212549 650505 212583 650539
rect 193229 650301 193263 650335
rect 222117 650505 222151 650539
rect 222117 650369 222151 650403
rect 231869 650505 231903 650539
rect 212549 650301 212583 650335
rect 241437 650505 241471 650539
rect 241437 650369 241471 650403
rect 251189 650505 251223 650539
rect 231869 650301 231903 650335
rect 260757 650505 260791 650539
rect 280169 650505 280203 650539
rect 289737 650641 289771 650675
rect 318809 650641 318843 650675
rect 328377 650777 328411 650811
rect 338129 650777 338163 650811
rect 338129 650641 338163 650675
rect 347697 650777 347731 650811
rect 357449 650777 357483 650811
rect 357449 650641 357483 650675
rect 367017 650777 367051 650811
rect 434729 650777 434763 650811
rect 425069 650641 425103 650675
rect 434729 650641 434763 650675
rect 444297 650777 444331 650811
rect 311817 650573 311851 650607
rect 311909 650573 311943 650607
rect 328377 650573 328411 650607
rect 331137 650573 331171 650607
rect 331229 650573 331263 650607
rect 347697 650573 347731 650607
rect 350457 650573 350491 650607
rect 350549 650573 350583 650607
rect 367017 650573 367051 650607
rect 369869 650573 369903 650607
rect 369961 650573 369995 650607
rect 405749 650505 405783 650539
rect 273177 650437 273211 650471
rect 273269 650437 273303 650471
rect 289737 650437 289771 650471
rect 292497 650437 292531 650471
rect 292589 650437 292623 650471
rect 260757 650369 260791 650403
rect 251189 650301 251223 650335
rect 454049 650777 454083 650811
rect 454049 650641 454083 650675
rect 463617 650777 463651 650811
rect 473369 650777 473403 650811
rect 473369 650641 473403 650675
rect 482937 650777 482971 650811
rect 492689 650777 492723 650811
rect 492689 650641 492723 650675
rect 502257 650777 502291 650811
rect 444297 650573 444331 650607
rect 447057 650573 447091 650607
rect 447149 650573 447183 650607
rect 463617 650573 463651 650607
rect 466377 650573 466411 650607
rect 466469 650573 466503 650607
rect 482937 650573 482971 650607
rect 485697 650573 485731 650607
rect 485789 650573 485823 650607
rect 502257 650573 502291 650607
rect 505109 650573 505143 650607
rect 505201 650573 505235 650607
rect 425069 650301 425103 650335
rect 405749 650165 405783 650199
rect 102885 558705 102919 558739
rect 97273 558637 97307 558671
rect 93869 558433 93903 558467
rect 93869 557889 93903 557923
rect 97089 557889 97123 557923
rect 99757 558637 99791 558671
rect 101965 558637 101999 558671
rect 99757 557889 99791 557923
rect 99849 558569 99883 558603
rect 99849 557889 99883 557923
rect 208593 558365 208627 558399
rect 325709 558365 325743 558399
rect 208593 557889 208627 557923
rect 222209 558093 222243 558127
rect 222209 557889 222243 557923
rect 231777 558025 231811 558059
rect 231777 557889 231811 557923
rect 93961 557821 93995 557855
rect 94881 557685 94915 557719
rect 98285 557821 98319 557855
rect 98285 557685 98319 557719
rect 106289 557821 106323 557855
rect 125425 557821 125459 557855
rect 325709 557821 325743 557855
rect 106289 557481 106323 557515
rect 115857 557753 115891 557787
rect 115857 557481 115891 557515
rect 128277 557549 128311 557583
rect 128369 557549 128403 557583
rect 125425 557481 125459 557515
rect 125609 557481 125643 557515
rect 125609 556869 125643 556903
rect 145481 543677 145515 543711
rect 152473 543677 152507 543711
rect 145481 542453 145515 542487
rect 152381 543541 152415 543575
rect 216781 543201 216815 543235
rect 216781 542929 216815 542963
rect 152473 542521 152507 542555
rect 152381 542385 152415 542419
rect 282101 431545 282135 431579
rect 281641 421345 281675 421379
rect 282101 417605 282135 417639
rect 281641 413865 281675 413899
rect 384589 414001 384623 414035
rect 384497 413797 384531 413831
rect 384589 413797 384623 413831
rect 386521 413797 386555 413831
rect 381369 413593 381403 413627
rect 375941 413457 375975 413491
rect 373917 412981 373951 413015
rect 378609 413389 378643 413423
rect 377413 413185 377447 413219
rect 377413 412981 377447 413015
rect 377505 413185 377539 413219
rect 375941 412913 375975 412947
rect 378885 413389 378919 413423
rect 378701 413185 378735 413219
rect 378609 413117 378643 413151
rect 384405 413389 384439 413423
rect 381369 412981 381403 413015
rect 384313 413321 384347 413355
rect 373917 412709 373951 412743
rect 377321 412709 377355 412743
rect 384221 412913 384255 412947
rect 384313 412709 384347 412743
rect 386521 413593 386555 413627
rect 387993 413593 388027 413627
rect 384497 413117 384531 413151
rect 384589 413389 384623 413423
rect 384589 413049 384623 413083
rect 384405 412709 384439 412743
rect 387901 412981 387935 413015
rect 387901 412641 387935 412675
rect 387993 412641 388027 412675
rect 384221 412573 384255 412607
rect 282193 395981 282227 396015
rect 282193 386393 282227 386427
rect 282285 369869 282319 369903
rect 282285 367149 282319 367183
rect 282101 366877 282135 366911
rect 282101 357425 282135 357459
rect 282377 338045 282411 338079
rect 282377 328457 282411 328491
rect 131037 318733 131071 318767
rect 97733 318597 97767 318631
rect 98101 318597 98135 318631
rect 131037 317509 131071 317543
rect 131865 4913 131899 4947
rect 130117 4845 130151 4879
rect 130485 4777 130519 4811
rect 131313 4777 131347 4811
rect 55229 4505 55263 4539
rect 16589 4097 16623 4131
rect 55229 4097 55263 4131
rect 64797 4505 64831 4539
rect 64797 4097 64831 4131
rect 84853 4097 84887 4131
rect 16589 3961 16623 3995
rect 80069 4029 80103 4063
rect 35909 3553 35943 3587
rect 35909 3417 35943 3451
rect 108313 4029 108347 4063
rect 84853 3893 84887 3927
rect 91293 3893 91327 3927
rect 55229 3349 55263 3383
rect 6837 3145 6871 3179
rect 6837 2873 6871 2907
rect 58541 3349 58575 3383
rect 64797 3349 64831 3383
rect 80069 3349 80103 3383
rect 69673 3281 69707 3315
rect 95617 3825 95651 3859
rect 108313 3825 108347 3859
rect 95617 3689 95651 3723
rect 91293 3213 91327 3247
rect 69673 3145 69707 3179
rect 68293 3077 68327 3111
rect 68477 3077 68511 3111
rect 58541 2805 58575 2839
rect 63785 2941 63819 2975
rect 64797 2941 64831 2975
rect 63509 2805 63543 2839
rect 55229 2669 55263 2703
<< metal1 >>
rect 260837 653395 260895 653401
rect 260837 653361 260849 653395
rect 260883 653392 260895 653395
rect 263594 653392 263600 653404
rect 260883 653364 263600 653392
rect 260883 653361 260895 653364
rect 260837 653355 260895 653361
rect 263594 653352 263600 653364
rect 263652 653392 263658 653404
rect 378134 653392 378140 653404
rect 263652 653364 378140 653392
rect 263652 653352 263658 653364
rect 378134 653352 378140 653364
rect 378192 653352 378198 653404
rect 383562 653352 383568 653404
rect 383620 653392 383626 653404
rect 508406 653392 508412 653404
rect 383620 653364 508412 653392
rect 383620 653352 383626 653364
rect 508406 653352 508412 653364
rect 508464 653352 508470 653404
rect 378134 652876 378140 652928
rect 378192 652916 378198 652928
rect 383562 652916 383568 652928
rect 378192 652888 383568 652916
rect 378192 652876 378198 652888
rect 383562 652876 383568 652888
rect 383620 652876 383626 652928
rect 139394 652848 139400 652860
rect 137664 652820 139400 652848
rect 135162 652740 135168 652792
rect 135220 652780 135226 652792
rect 137664 652780 137692 652820
rect 139394 652808 139400 652820
rect 139452 652848 139458 652860
rect 139452 652820 139716 652848
rect 139452 652808 139458 652820
rect 135220 652752 137692 652780
rect 139688 652780 139716 652820
rect 508406 652808 508412 652860
rect 508464 652848 508470 652860
rect 513374 652848 513380 652860
rect 508464 652820 513380 652848
rect 508464 652808 508470 652820
rect 513374 652808 513380 652820
rect 513432 652808 513438 652860
rect 258534 652780 258540 652792
rect 139688 652752 258540 652780
rect 135220 652740 135226 652752
rect 258534 652740 258540 652752
rect 258592 652780 258598 652792
rect 260837 652783 260895 652789
rect 260837 652780 260849 652783
rect 258592 652752 260849 652780
rect 258592 652740 258598 652752
rect 260837 652749 260849 652752
rect 260883 652749 260895 652783
rect 513392 652780 513420 652808
rect 518894 652780 518900 652792
rect 513392 652752 518900 652780
rect 260837 652743 260895 652749
rect 518894 652740 518900 652752
rect 518952 652740 518958 652792
rect 318797 650811 318855 650817
rect 318797 650777 318809 650811
rect 318843 650808 318855 650811
rect 328365 650811 328423 650817
rect 328365 650808 328377 650811
rect 318843 650780 328377 650808
rect 318843 650777 318855 650780
rect 318797 650771 318855 650777
rect 328365 650777 328377 650780
rect 328411 650777 328423 650811
rect 328365 650771 328423 650777
rect 338117 650811 338175 650817
rect 338117 650777 338129 650811
rect 338163 650808 338175 650811
rect 347685 650811 347743 650817
rect 347685 650808 347697 650811
rect 338163 650780 347697 650808
rect 338163 650777 338175 650780
rect 338117 650771 338175 650777
rect 347685 650777 347697 650780
rect 347731 650777 347743 650811
rect 347685 650771 347743 650777
rect 357437 650811 357495 650817
rect 357437 650777 357449 650811
rect 357483 650808 357495 650811
rect 367005 650811 367063 650817
rect 367005 650808 367017 650811
rect 357483 650780 367017 650808
rect 357483 650777 357495 650780
rect 357437 650771 357495 650777
rect 367005 650777 367017 650780
rect 367051 650777 367063 650811
rect 367005 650771 367063 650777
rect 434717 650811 434775 650817
rect 434717 650777 434729 650811
rect 434763 650808 434775 650811
rect 444285 650811 444343 650817
rect 444285 650808 444297 650811
rect 434763 650780 444297 650808
rect 434763 650777 434775 650780
rect 434717 650771 434775 650777
rect 444285 650777 444297 650780
rect 444331 650777 444343 650811
rect 444285 650771 444343 650777
rect 454037 650811 454095 650817
rect 454037 650777 454049 650811
rect 454083 650808 454095 650811
rect 463605 650811 463663 650817
rect 463605 650808 463617 650811
rect 454083 650780 463617 650808
rect 454083 650777 454095 650780
rect 454037 650771 454095 650777
rect 463605 650777 463617 650780
rect 463651 650777 463663 650811
rect 463605 650771 463663 650777
rect 473357 650811 473415 650817
rect 473357 650777 473369 650811
rect 473403 650808 473415 650811
rect 482925 650811 482983 650817
rect 482925 650808 482937 650811
rect 473403 650780 482937 650808
rect 473403 650777 473415 650780
rect 473357 650771 473415 650777
rect 482925 650777 482937 650780
rect 482971 650777 482983 650811
rect 482925 650771 482983 650777
rect 492677 650811 492735 650817
rect 492677 650777 492689 650811
rect 492723 650808 492735 650811
rect 502245 650811 502303 650817
rect 502245 650808 502257 650811
rect 492723 650780 502257 650808
rect 492723 650777 492735 650780
rect 492677 650771 492735 650777
rect 502245 650777 502257 650780
rect 502291 650777 502303 650811
rect 502245 650771 502303 650777
rect 280157 650675 280215 650681
rect 280157 650641 280169 650675
rect 280203 650672 280215 650675
rect 289725 650675 289783 650681
rect 289725 650672 289737 650675
rect 280203 650644 289737 650672
rect 280203 650641 280215 650644
rect 280157 650635 280215 650641
rect 289725 650641 289737 650644
rect 289771 650641 289783 650675
rect 318797 650675 318855 650681
rect 318797 650672 318809 650675
rect 289725 650635 289783 650641
rect 313108 650644 318809 650672
rect 311805 650607 311863 650613
rect 311805 650604 311817 650607
rect 302160 650576 311817 650604
rect 193217 650539 193275 650545
rect 193217 650505 193229 650539
rect 193263 650536 193275 650539
rect 202785 650539 202843 650545
rect 202785 650536 202797 650539
rect 193263 650508 202797 650536
rect 193263 650505 193275 650508
rect 193217 650499 193275 650505
rect 202785 650505 202797 650508
rect 202831 650505 202843 650539
rect 202785 650499 202843 650505
rect 212537 650539 212595 650545
rect 212537 650505 212549 650539
rect 212583 650536 212595 650539
rect 222105 650539 222163 650545
rect 222105 650536 222117 650539
rect 212583 650508 222117 650536
rect 212583 650505 212595 650508
rect 212537 650499 212595 650505
rect 222105 650505 222117 650508
rect 222151 650505 222163 650539
rect 222105 650499 222163 650505
rect 231857 650539 231915 650545
rect 231857 650505 231869 650539
rect 231903 650536 231915 650539
rect 241425 650539 241483 650545
rect 241425 650536 241437 650539
rect 231903 650508 241437 650536
rect 231903 650505 231915 650508
rect 231857 650499 231915 650505
rect 241425 650505 241437 650508
rect 241471 650505 241483 650539
rect 241425 650499 241483 650505
rect 251177 650539 251235 650545
rect 251177 650505 251189 650539
rect 251223 650536 251235 650539
rect 260745 650539 260803 650545
rect 260745 650536 260757 650539
rect 251223 650508 260757 650536
rect 251223 650505 251235 650508
rect 251177 650499 251235 650505
rect 260745 650505 260757 650508
rect 260791 650505 260803 650539
rect 280157 650539 280215 650545
rect 280157 650536 280169 650539
rect 260745 650499 260803 650505
rect 274468 650508 280169 650536
rect 266630 650468 266636 650480
rect 263520 650440 266636 650468
rect 202785 650403 202843 650409
rect 202785 650369 202797 650403
rect 202831 650369 202843 650403
rect 202785 650363 202843 650369
rect 222105 650403 222163 650409
rect 222105 650369 222117 650403
rect 222151 650369 222163 650403
rect 222105 650363 222163 650369
rect 241425 650403 241483 650409
rect 241425 650369 241437 650403
rect 241471 650369 241483 650403
rect 241425 650363 241483 650369
rect 260745 650403 260803 650409
rect 260745 650369 260757 650403
rect 260791 650400 260803 650403
rect 263520 650400 263548 650440
rect 266630 650428 266636 650440
rect 266688 650468 266694 650480
rect 273165 650471 273223 650477
rect 273165 650468 273177 650471
rect 266688 650440 273177 650468
rect 266688 650428 266694 650440
rect 273165 650437 273177 650440
rect 273211 650437 273223 650471
rect 273165 650431 273223 650437
rect 273257 650471 273315 650477
rect 273257 650437 273269 650471
rect 273303 650468 273315 650471
rect 274468 650468 274496 650508
rect 280157 650505 280169 650508
rect 280203 650505 280215 650539
rect 302160 650536 302188 650576
rect 311805 650573 311817 650576
rect 311851 650573 311863 650607
rect 311805 650567 311863 650573
rect 311897 650607 311955 650613
rect 311897 650573 311909 650607
rect 311943 650604 311955 650607
rect 313108 650604 313136 650644
rect 318797 650641 318809 650644
rect 318843 650641 318855 650675
rect 338117 650675 338175 650681
rect 338117 650672 338129 650675
rect 318797 650635 318855 650641
rect 332428 650644 338129 650672
rect 311943 650576 313136 650604
rect 328365 650607 328423 650613
rect 311943 650573 311955 650576
rect 311897 650567 311955 650573
rect 328365 650573 328377 650607
rect 328411 650604 328423 650607
rect 331125 650607 331183 650613
rect 331125 650604 331137 650607
rect 328411 650576 331137 650604
rect 328411 650573 328423 650576
rect 328365 650567 328423 650573
rect 331125 650573 331137 650576
rect 331171 650573 331183 650607
rect 331125 650567 331183 650573
rect 331217 650607 331275 650613
rect 331217 650573 331229 650607
rect 331263 650604 331275 650607
rect 332428 650604 332456 650644
rect 338117 650641 338129 650644
rect 338163 650641 338175 650675
rect 357437 650675 357495 650681
rect 357437 650672 357449 650675
rect 338117 650635 338175 650641
rect 351748 650644 357449 650672
rect 331263 650576 332456 650604
rect 347685 650607 347743 650613
rect 331263 650573 331275 650576
rect 331217 650567 331275 650573
rect 347685 650573 347697 650607
rect 347731 650604 347743 650607
rect 350445 650607 350503 650613
rect 350445 650604 350457 650607
rect 347731 650576 350457 650604
rect 347731 650573 347743 650576
rect 347685 650567 347743 650573
rect 350445 650573 350457 650576
rect 350491 650573 350503 650607
rect 350445 650567 350503 650573
rect 350537 650607 350595 650613
rect 350537 650573 350549 650607
rect 350583 650604 350595 650607
rect 351748 650604 351776 650644
rect 357437 650641 357449 650644
rect 357483 650641 357495 650675
rect 357437 650635 357495 650641
rect 425057 650675 425115 650681
rect 425057 650641 425069 650675
rect 425103 650672 425115 650675
rect 434717 650675 434775 650681
rect 434717 650672 434729 650675
rect 425103 650644 434729 650672
rect 425103 650641 425115 650644
rect 425057 650635 425115 650641
rect 434717 650641 434729 650644
rect 434763 650641 434775 650675
rect 454037 650675 454095 650681
rect 454037 650672 454049 650675
rect 434717 650635 434775 650641
rect 448348 650644 454049 650672
rect 350583 650576 351776 650604
rect 367005 650607 367063 650613
rect 350583 650573 350595 650576
rect 350537 650567 350595 650573
rect 367005 650573 367017 650607
rect 367051 650604 367063 650607
rect 369857 650607 369915 650613
rect 369857 650604 369869 650607
rect 367051 650576 369869 650604
rect 367051 650573 367063 650576
rect 367005 650567 367063 650573
rect 369857 650573 369869 650576
rect 369903 650573 369915 650607
rect 369857 650567 369915 650573
rect 369949 650607 370007 650613
rect 369949 650573 369961 650607
rect 369995 650604 370007 650607
rect 444285 650607 444343 650613
rect 369995 650576 376708 650604
rect 369995 650573 370007 650576
rect 369949 650567 370007 650573
rect 280157 650499 280215 650505
rect 293788 650508 302188 650536
rect 376680 650536 376708 650576
rect 444285 650573 444297 650607
rect 444331 650604 444343 650607
rect 447045 650607 447103 650613
rect 447045 650604 447057 650607
rect 444331 650576 447057 650604
rect 444331 650573 444343 650576
rect 444285 650567 444343 650573
rect 447045 650573 447057 650576
rect 447091 650573 447103 650607
rect 447045 650567 447103 650573
rect 447137 650607 447195 650613
rect 447137 650573 447149 650607
rect 447183 650604 447195 650607
rect 448348 650604 448376 650644
rect 454037 650641 454049 650644
rect 454083 650641 454095 650675
rect 473357 650675 473415 650681
rect 473357 650672 473369 650675
rect 454037 650635 454095 650641
rect 467668 650644 473369 650672
rect 447183 650576 448376 650604
rect 463605 650607 463663 650613
rect 447183 650573 447195 650576
rect 447137 650567 447195 650573
rect 463605 650573 463617 650607
rect 463651 650604 463663 650607
rect 466365 650607 466423 650613
rect 466365 650604 466377 650607
rect 463651 650576 466377 650604
rect 463651 650573 463663 650576
rect 463605 650567 463663 650573
rect 466365 650573 466377 650576
rect 466411 650573 466423 650607
rect 466365 650567 466423 650573
rect 466457 650607 466515 650613
rect 466457 650573 466469 650607
rect 466503 650604 466515 650607
rect 467668 650604 467696 650644
rect 473357 650641 473369 650644
rect 473403 650641 473415 650675
rect 492677 650675 492735 650681
rect 492677 650672 492689 650675
rect 473357 650635 473415 650641
rect 486988 650644 492689 650672
rect 466503 650576 467696 650604
rect 482925 650607 482983 650613
rect 466503 650573 466515 650576
rect 466457 650567 466515 650573
rect 482925 650573 482937 650607
rect 482971 650604 482983 650607
rect 485685 650607 485743 650613
rect 485685 650604 485697 650607
rect 482971 650576 485697 650604
rect 482971 650573 482983 650576
rect 482925 650567 482983 650573
rect 485685 650573 485697 650576
rect 485731 650573 485743 650607
rect 485685 650567 485743 650573
rect 485777 650607 485835 650613
rect 485777 650573 485789 650607
rect 485823 650604 485835 650607
rect 486988 650604 487016 650644
rect 492677 650641 492689 650644
rect 492723 650641 492735 650675
rect 492677 650635 492735 650641
rect 485823 650576 487016 650604
rect 502245 650607 502303 650613
rect 485823 650573 485835 650576
rect 485777 650567 485835 650573
rect 502245 650573 502257 650607
rect 502291 650604 502303 650607
rect 505097 650607 505155 650613
rect 505097 650604 505109 650607
rect 502291 650576 505109 650604
rect 502291 650573 502303 650576
rect 502245 650567 502303 650573
rect 505097 650573 505109 650576
rect 505143 650573 505155 650607
rect 505097 650567 505155 650573
rect 505189 650607 505247 650613
rect 505189 650573 505201 650607
rect 505235 650604 505247 650607
rect 505235 650576 511948 650604
rect 505235 650573 505247 650576
rect 505189 650567 505247 650573
rect 405737 650539 405795 650545
rect 376680 650508 379468 650536
rect 273303 650440 274496 650468
rect 289725 650471 289783 650477
rect 273303 650437 273315 650440
rect 273257 650431 273315 650437
rect 289725 650437 289737 650471
rect 289771 650468 289783 650471
rect 292485 650471 292543 650477
rect 292485 650468 292497 650471
rect 289771 650440 292497 650468
rect 289771 650437 289783 650440
rect 289725 650431 289783 650437
rect 292485 650437 292497 650440
rect 292531 650437 292543 650471
rect 292485 650431 292543 650437
rect 292577 650471 292635 650477
rect 292577 650437 292589 650471
rect 292623 650468 292635 650471
rect 293788 650468 293816 650508
rect 292623 650440 293816 650468
rect 379440 650468 379468 650508
rect 405737 650505 405749 650539
rect 405783 650536 405795 650539
rect 407758 650536 407764 650548
rect 405783 650508 407764 650536
rect 405783 650505 405795 650508
rect 405737 650499 405795 650505
rect 407758 650496 407764 650508
rect 407816 650536 407822 650548
rect 511920 650536 511948 650576
rect 407816 650508 416268 650536
rect 511920 650508 514708 650536
rect 407816 650496 407822 650508
rect 387150 650468 387156 650480
rect 379440 650440 387156 650468
rect 292623 650437 292635 650440
rect 292577 650431 292635 650437
rect 387150 650428 387156 650440
rect 387208 650428 387214 650480
rect 260791 650372 263548 650400
rect 260791 650369 260803 650372
rect 260745 650363 260803 650369
rect 193217 650335 193275 650341
rect 193217 650332 193229 650335
rect 144840 650304 154620 650332
rect 137646 650224 137652 650276
rect 137704 650264 137710 650276
rect 144840 650264 144868 650304
rect 137704 650236 144868 650264
rect 154592 650264 154620 650304
rect 164160 650304 173940 650332
rect 164160 650264 164188 650304
rect 154592 650236 164188 650264
rect 173912 650264 173940 650304
rect 183480 650304 193229 650332
rect 183480 650264 183508 650304
rect 193217 650301 193229 650304
rect 193263 650301 193275 650335
rect 202800 650332 202828 650363
rect 212537 650335 212595 650341
rect 212537 650332 212549 650335
rect 202800 650304 212549 650332
rect 193217 650295 193275 650301
rect 212537 650301 212549 650304
rect 212583 650301 212595 650335
rect 222120 650332 222148 650363
rect 231857 650335 231915 650341
rect 231857 650332 231869 650335
rect 222120 650304 231869 650332
rect 212537 650295 212595 650301
rect 231857 650301 231869 650304
rect 231903 650301 231915 650335
rect 241440 650332 241468 650363
rect 251177 650335 251235 650341
rect 251177 650332 251189 650335
rect 241440 650304 251189 650332
rect 231857 650295 231915 650301
rect 251177 650301 251189 650304
rect 251223 650301 251235 650335
rect 416240 650332 416268 650508
rect 514680 650468 514708 650508
rect 516410 650468 516416 650480
rect 514680 650440 516416 650468
rect 516410 650428 516416 650440
rect 516468 650428 516474 650480
rect 425057 650335 425115 650341
rect 425057 650332 425069 650335
rect 416240 650304 425069 650332
rect 251177 650295 251235 650301
rect 425057 650301 425069 650304
rect 425103 650301 425115 650335
rect 425057 650295 425115 650301
rect 173912 650236 183508 650264
rect 137704 650224 137710 650236
rect 389174 650156 389180 650208
rect 389232 650196 389238 650208
rect 405737 650199 405795 650205
rect 405737 650196 405749 650199
rect 389232 650168 405749 650196
rect 389232 650156 389238 650168
rect 405737 650165 405749 650168
rect 405783 650165 405795 650199
rect 405737 650159 405795 650165
rect 291838 645872 291844 645924
rect 291896 645912 291902 645924
rect 307386 645912 307392 645924
rect 291896 645884 307392 645912
rect 291896 645872 291902 645884
rect 307386 645872 307392 645884
rect 307444 645872 307450 645924
rect 290458 644444 290464 644496
rect 290516 644484 290522 644496
rect 307110 644484 307116 644496
rect 290516 644456 307116 644484
rect 290516 644444 290522 644456
rect 307110 644444 307116 644456
rect 307168 644444 307174 644496
rect 287698 643084 287704 643136
rect 287756 643124 287762 643136
rect 307110 643124 307116 643136
rect 287756 643096 307116 643124
rect 287756 643084 287762 643096
rect 307110 643084 307116 643096
rect 307168 643084 307174 643136
rect 286318 641724 286324 641776
rect 286376 641764 286382 641776
rect 307662 641764 307668 641776
rect 286376 641736 307668 641764
rect 286376 641724 286382 641736
rect 307662 641724 307668 641736
rect 307720 641724 307726 641776
rect 284938 640296 284944 640348
rect 284996 640336 285002 640348
rect 307662 640336 307668 640348
rect 284996 640308 307668 640336
rect 284996 640296 285002 640308
rect 307662 640296 307668 640308
rect 307720 640296 307726 640348
rect 291930 637576 291936 637628
rect 291988 637616 291994 637628
rect 306834 637616 306840 637628
rect 291988 637588 306840 637616
rect 291988 637576 291994 637588
rect 306834 637576 306840 637588
rect 306892 637576 306898 637628
rect 270402 580252 270408 580304
rect 270460 580292 270466 580304
rect 279142 580292 279148 580304
rect 270460 580264 279148 580292
rect 270460 580252 270466 580264
rect 279142 580252 279148 580264
rect 279200 580252 279206 580304
rect 302878 579640 302884 579692
rect 302936 579680 302942 579692
rect 307662 579680 307668 579692
rect 302936 579652 307668 579680
rect 302936 579640 302942 579652
rect 307662 579640 307668 579652
rect 307720 579640 307726 579692
rect 313826 558940 313832 558952
rect 313292 558912 313832 558940
rect 77386 558832 77392 558884
rect 77444 558872 77450 558884
rect 86310 558872 86316 558884
rect 77444 558844 86316 558872
rect 77444 558832 77450 558844
rect 86310 558832 86316 558844
rect 86368 558872 86374 558884
rect 86678 558872 86684 558884
rect 86368 558844 86684 558872
rect 86368 558832 86374 558844
rect 86678 558832 86684 558844
rect 86736 558832 86742 558884
rect 93762 558832 93768 558884
rect 93820 558872 93826 558884
rect 137278 558872 137284 558884
rect 93820 558844 137284 558872
rect 93820 558832 93826 558844
rect 137278 558832 137284 558844
rect 137336 558832 137342 558884
rect 194410 558832 194416 558884
rect 194468 558872 194474 558884
rect 313292 558872 313320 558912
rect 313826 558900 313832 558912
rect 313884 558940 313890 558952
rect 413922 558940 413928 558952
rect 313884 558912 413928 558940
rect 313884 558900 313890 558912
rect 413922 558900 413928 558912
rect 413980 558900 413986 558952
rect 194468 558844 313320 558872
rect 194468 558832 194474 558844
rect 347682 558832 347688 558884
rect 347740 558872 347746 558884
rect 356054 558872 356060 558884
rect 347740 558844 356060 558872
rect 347740 558832 347746 558844
rect 356054 558832 356060 558844
rect 356112 558832 356118 558884
rect 468018 558832 468024 558884
rect 468076 558872 468082 558884
rect 476574 558872 476580 558884
rect 468076 558844 476580 558872
rect 468076 558832 468082 558844
rect 476574 558832 476580 558844
rect 476632 558832 476638 558884
rect 66162 558764 66168 558816
rect 66220 558804 66226 558816
rect 200206 558804 200212 558816
rect 66220 558776 200212 558804
rect 66220 558764 66226 558776
rect 200206 558764 200212 558776
rect 200264 558764 200270 558816
rect 215294 558764 215300 558816
rect 215352 558804 215358 558816
rect 224494 558804 224500 558816
rect 215352 558776 224500 558804
rect 215352 558764 215358 558776
rect 224494 558764 224500 558776
rect 224552 558764 224558 558816
rect 286410 558764 286416 558816
rect 286468 558804 286474 558816
rect 453666 558804 453672 558816
rect 286468 558776 453672 558804
rect 286468 558764 286474 558776
rect 453666 558764 453672 558776
rect 453724 558804 453730 558816
rect 453724 558776 455368 558804
rect 453724 558764 453730 558776
rect 74994 558696 75000 558748
rect 75052 558736 75058 558748
rect 84194 558736 84200 558748
rect 75052 558708 84200 558736
rect 75052 558696 75058 558708
rect 84194 558696 84200 558708
rect 84252 558736 84258 558748
rect 93302 558736 93308 558748
rect 84252 558708 93308 558736
rect 84252 558696 84258 558708
rect 93302 558696 93308 558708
rect 93360 558736 93366 558748
rect 102778 558736 102784 558748
rect 93360 558708 102784 558736
rect 93360 558696 93366 558708
rect 102778 558696 102784 558708
rect 102836 558696 102842 558748
rect 102873 558739 102931 558745
rect 102873 558705 102885 558739
rect 102919 558736 102931 558739
rect 106274 558736 106280 558748
rect 102919 558708 106280 558736
rect 102919 558705 102931 558708
rect 102873 558699 102931 558705
rect 106274 558696 106280 558708
rect 106332 558696 106338 558748
rect 107286 558696 107292 558748
rect 107344 558736 107350 558748
rect 141418 558736 141424 558748
rect 107344 558708 141424 558736
rect 107344 558696 107350 558708
rect 141418 558696 141424 558708
rect 141476 558696 141482 558748
rect 218790 558696 218796 558748
rect 218848 558736 218854 558748
rect 227990 558736 227996 558748
rect 218848 558708 227996 558736
rect 218848 558696 218854 558708
rect 227990 558696 227996 558708
rect 228048 558736 228054 558748
rect 237374 558736 237380 558748
rect 228048 558708 237380 558736
rect 228048 558696 228054 558708
rect 237374 558696 237380 558708
rect 237432 558696 237438 558748
rect 286502 558696 286508 558748
rect 286560 558736 286566 558748
rect 454770 558736 454776 558748
rect 286560 558708 454776 558736
rect 286560 558696 286566 558708
rect 454770 558696 454776 558708
rect 454828 558696 454834 558748
rect 78490 558628 78496 558680
rect 78548 558668 78554 558680
rect 87874 558668 87880 558680
rect 78548 558640 87880 558668
rect 78548 558628 78554 558640
rect 87874 558628 87880 558640
rect 87932 558668 87938 558680
rect 97166 558668 97172 558680
rect 87932 558640 97172 558668
rect 87932 558628 87938 558640
rect 97166 558628 97172 558640
rect 97224 558628 97230 558680
rect 97261 558671 97319 558677
rect 97261 558637 97273 558671
rect 97307 558668 97319 558671
rect 99466 558668 99472 558680
rect 97307 558640 99472 558668
rect 97307 558637 97319 558640
rect 97261 558631 97319 558637
rect 99466 558628 99472 558640
rect 99524 558628 99530 558680
rect 99745 558671 99803 558677
rect 99745 558637 99757 558671
rect 99791 558668 99803 558671
rect 101953 558671 102011 558677
rect 101953 558668 101965 558671
rect 99791 558640 101965 558668
rect 99791 558637 99803 558640
rect 99745 558631 99803 558637
rect 101953 558637 101965 558640
rect 101999 558637 102011 558671
rect 101953 558631 102011 558637
rect 102042 558628 102048 558680
rect 102100 558668 102106 558680
rect 140038 558668 140044 558680
rect 102100 558640 140044 558668
rect 102100 558628 102106 558640
rect 140038 558628 140044 558640
rect 140096 558628 140102 558680
rect 222194 558628 222200 558680
rect 222252 558668 222258 558680
rect 231854 558668 231860 558680
rect 222252 558640 231860 558668
rect 222252 558628 222258 558640
rect 231854 558628 231860 558640
rect 231912 558628 231918 558680
rect 326338 558628 326344 558680
rect 326396 558668 326402 558680
rect 335446 558668 335452 558680
rect 326396 558640 335452 558668
rect 326396 558628 326402 558640
rect 335446 558628 335452 558640
rect 335504 558668 335510 558680
rect 344278 558668 344284 558680
rect 335504 558640 344284 558668
rect 335504 558628 335510 558640
rect 344278 558628 344284 558640
rect 344336 558668 344342 558680
rect 353294 558668 353300 558680
rect 344336 558640 353300 558668
rect 344336 558628 344342 558640
rect 353294 558628 353300 558640
rect 353352 558628 353358 558680
rect 75914 558560 75920 558612
rect 75972 558600 75978 558612
rect 85390 558600 85396 558612
rect 75972 558572 85396 558600
rect 75972 558560 75978 558572
rect 85390 558560 85396 558572
rect 85448 558560 85454 558612
rect 86678 558560 86684 558612
rect 86736 558600 86742 558612
rect 95694 558600 95700 558612
rect 86736 558572 95700 558600
rect 86736 558560 86742 558572
rect 95694 558560 95700 558572
rect 95752 558600 95758 558612
rect 99837 558603 99895 558609
rect 99837 558600 99849 558603
rect 95752 558572 99849 558600
rect 95752 558560 95758 558572
rect 99837 558569 99849 558572
rect 99883 558569 99895 558603
rect 104158 558600 104164 558612
rect 99837 558563 99895 558569
rect 99944 558572 104164 558600
rect 79410 558492 79416 558544
rect 79468 558532 79474 558544
rect 88886 558532 88892 558544
rect 79468 558504 88892 558532
rect 79468 558492 79474 558504
rect 88886 558492 88892 558504
rect 88944 558532 88950 558544
rect 98362 558532 98368 558544
rect 88944 558504 98368 558532
rect 88944 558492 88950 558504
rect 98362 558492 98368 558504
rect 98420 558492 98426 558544
rect 99944 558532 99972 558572
rect 104158 558560 104164 558572
rect 104216 558560 104222 558612
rect 108482 558560 108488 558612
rect 108540 558600 108546 558612
rect 148318 558600 148324 558612
rect 108540 558572 148324 558600
rect 108540 558560 108546 558572
rect 148318 558560 148324 558572
rect 148376 558560 148382 558612
rect 217502 558560 217508 558612
rect 217560 558600 217566 558612
rect 225874 558600 225880 558612
rect 217560 558572 225880 558600
rect 217560 558560 217566 558572
rect 225874 558560 225880 558572
rect 225932 558600 225938 558612
rect 234614 558600 234620 558612
rect 225932 558572 234620 558600
rect 225932 558560 225938 558572
rect 234614 558560 234620 558572
rect 234672 558560 234678 558612
rect 336090 558560 336096 558612
rect 336148 558600 336154 558612
rect 336642 558600 336648 558612
rect 336148 558572 336648 558600
rect 336148 558560 336154 558572
rect 336642 558560 336648 558572
rect 336700 558600 336706 558612
rect 346026 558600 346032 558612
rect 336700 558572 346032 558600
rect 336700 558560 336706 558572
rect 346026 558560 346032 558572
rect 346084 558600 346090 558612
rect 354674 558600 354680 558612
rect 346084 558572 354680 558600
rect 346084 558560 346090 558572
rect 354674 558560 354680 558572
rect 354732 558560 354738 558612
rect 455340 558600 455368 558776
rect 457438 558764 457444 558816
rect 457496 558804 457502 558816
rect 466546 558804 466552 558816
rect 457496 558776 466552 558804
rect 457496 558764 457502 558776
rect 466546 558764 466552 558776
rect 466604 558804 466610 558816
rect 475470 558804 475476 558816
rect 466604 558776 475476 558804
rect 466604 558764 466610 558776
rect 475470 558764 475476 558776
rect 475528 558804 475534 558816
rect 475528 558776 477724 558804
rect 475528 558764 475534 558776
rect 458818 558696 458824 558748
rect 458876 558736 458882 558748
rect 468018 558736 468024 558748
rect 458876 558708 468024 558736
rect 458876 558696 458882 558708
rect 468018 558696 468024 558708
rect 468076 558696 468082 558748
rect 468110 558696 468116 558748
rect 468168 558736 468174 558748
rect 468754 558736 468760 558748
rect 468168 558708 468760 558736
rect 468168 558696 468174 558708
rect 468754 558696 468760 558708
rect 468812 558736 468818 558748
rect 477586 558736 477592 558748
rect 468812 558708 477592 558736
rect 468812 558696 468818 558708
rect 477586 558696 477592 558708
rect 477644 558696 477650 558748
rect 456058 558628 456064 558680
rect 456116 558668 456122 558680
rect 465258 558668 465264 558680
rect 456116 558640 465264 558668
rect 456116 558628 456122 558640
rect 465258 558628 465264 558640
rect 465316 558668 465322 558680
rect 474826 558668 474832 558680
rect 465316 558640 474832 558668
rect 465316 558628 465322 558640
rect 474826 558628 474832 558640
rect 474884 558628 474890 558680
rect 477696 558668 477724 558776
rect 484394 558668 484400 558680
rect 477696 558640 484400 558668
rect 484394 558628 484400 558640
rect 484452 558628 484458 558680
rect 463050 558600 463056 558612
rect 455340 558572 463056 558600
rect 463050 558560 463056 558572
rect 463108 558600 463114 558612
rect 472158 558600 472164 558612
rect 463108 558572 472164 558600
rect 463108 558560 463114 558572
rect 472158 558560 472164 558572
rect 472216 558600 472222 558612
rect 481634 558600 481640 558612
rect 472216 558572 481640 558600
rect 472216 558560 472222 558572
rect 481634 558560 481640 558572
rect 481692 558560 481698 558612
rect 98472 558504 99972 558532
rect 80790 558424 80796 558476
rect 80848 558464 80854 558476
rect 89806 558464 89812 558476
rect 80848 558436 89812 558464
rect 80848 558424 80854 558436
rect 89806 558424 89812 558436
rect 89864 558464 89870 558476
rect 93857 558467 93915 558473
rect 93857 558464 93869 558467
rect 89864 558436 93869 558464
rect 89864 558424 89870 558436
rect 93857 558433 93869 558436
rect 93903 558433 93915 558467
rect 93857 558427 93915 558433
rect 94774 558424 94780 558476
rect 94832 558464 94838 558476
rect 98472 558464 98500 558504
rect 100018 558492 100024 558544
rect 100076 558532 100082 558544
rect 100076 558504 104296 558532
rect 100076 558492 100082 558504
rect 94832 558436 98500 558464
rect 104268 558464 104296 558504
rect 104802 558492 104808 558544
rect 104860 558532 104866 558544
rect 144178 558532 144184 558544
rect 104860 558504 144184 558532
rect 104860 558492 104866 558504
rect 144178 558492 144184 558504
rect 144236 558492 144242 558544
rect 208486 558492 208492 558544
rect 208544 558532 208550 558544
rect 217594 558532 217600 558544
rect 208544 558504 217600 558532
rect 208544 558492 208550 558504
rect 217594 558492 217600 558504
rect 217652 558532 217658 558544
rect 227162 558532 227168 558544
rect 217652 558504 227168 558532
rect 217652 558492 217658 558504
rect 227162 558492 227168 558504
rect 227220 558532 227226 558544
rect 235994 558532 236000 558544
rect 227220 558504 236000 558532
rect 227220 558492 227226 558504
rect 235994 558492 236000 558504
rect 236052 558492 236058 558544
rect 330478 558492 330484 558544
rect 330536 558532 330542 558544
rect 339862 558532 339868 558544
rect 330536 558504 339868 558532
rect 330536 558492 330542 558504
rect 339862 558492 339868 558504
rect 339920 558532 339926 558544
rect 349706 558532 349712 558544
rect 339920 558504 349712 558532
rect 339920 558492 339926 558504
rect 349706 558492 349712 558504
rect 349764 558532 349770 558544
rect 358170 558532 358176 558544
rect 349764 558504 358176 558532
rect 349764 558492 349770 558504
rect 358170 558492 358176 558504
rect 358228 558492 358234 558544
rect 453298 558492 453304 558544
rect 453356 558532 453362 558544
rect 461670 558532 461676 558544
rect 453356 558504 461676 558532
rect 453356 558492 453362 558504
rect 461670 558492 461676 558504
rect 461728 558532 461734 558544
rect 471330 558532 471336 558544
rect 461728 558504 471336 558532
rect 461728 558492 461734 558504
rect 471330 558492 471336 558504
rect 471388 558532 471394 558544
rect 480346 558532 480352 558544
rect 471388 558504 480352 558532
rect 471388 558492 471394 558504
rect 480346 558492 480352 558504
rect 480404 558492 480410 558544
rect 140130 558464 140136 558476
rect 104268 558436 140136 558464
rect 94832 558424 94838 558436
rect 140130 558424 140136 558436
rect 140188 558424 140194 558476
rect 213178 558424 213184 558476
rect 213236 558464 213242 558476
rect 222194 558464 222200 558476
rect 213236 558436 222200 558464
rect 213236 558424 213242 558436
rect 222194 558424 222200 558436
rect 222252 558424 222258 558476
rect 329282 558424 329288 558476
rect 329340 558464 329346 558476
rect 339034 558464 339040 558476
rect 329340 558436 339040 558464
rect 329340 558424 329346 558436
rect 339034 558424 339040 558436
rect 339092 558464 339098 558476
rect 348234 558464 348240 558476
rect 339092 558436 348240 558464
rect 339092 558424 339098 558436
rect 348234 558424 348240 558436
rect 348292 558464 348298 558476
rect 357434 558464 357440 558476
rect 348292 558436 357440 558464
rect 348292 558424 348298 558436
rect 357434 558424 357440 558436
rect 357492 558424 357498 558476
rect 413922 558424 413928 558476
rect 413980 558464 413986 558476
rect 443086 558464 443092 558476
rect 413980 558436 443092 558464
rect 413980 558424 413986 558436
rect 443086 558424 443092 558436
rect 443144 558424 443150 558476
rect 454770 558424 454776 558476
rect 454828 558464 454834 558476
rect 464246 558464 464252 558476
rect 454828 558436 464252 558464
rect 454828 558424 454834 558436
rect 464246 558424 464252 558436
rect 464304 558464 464310 558476
rect 473446 558464 473452 558476
rect 464304 558436 473452 558464
rect 464304 558424 464310 558436
rect 473446 558424 473452 558436
rect 473504 558464 473510 558476
rect 483014 558464 483020 558476
rect 473504 558436 483020 558464
rect 473504 558424 473510 558436
rect 483014 558424 483020 558436
rect 483072 558424 483078 558476
rect 73706 558356 73712 558408
rect 73764 558396 73770 558408
rect 82906 558396 82912 558408
rect 73764 558368 82912 558396
rect 73764 558356 73770 558368
rect 82906 558356 82912 558368
rect 82964 558396 82970 558408
rect 92474 558396 92480 558408
rect 82964 558368 92480 558396
rect 82964 558356 82970 558368
rect 92474 558356 92480 558368
rect 92532 558396 92538 558408
rect 93118 558396 93124 558408
rect 92532 558368 93124 558396
rect 92532 558356 92538 558368
rect 93118 558356 93124 558368
rect 93176 558356 93182 558408
rect 97810 558356 97816 558408
rect 97868 558396 97874 558408
rect 138658 558396 138664 558408
rect 97868 558368 138664 558396
rect 97868 558356 97874 558368
rect 138658 558356 138664 558368
rect 138716 558356 138722 558408
rect 208581 558399 208639 558405
rect 208581 558365 208593 558399
rect 208627 558396 208639 558399
rect 210602 558396 210608 558408
rect 208627 558368 210608 558396
rect 208627 558365 208639 558368
rect 208581 558359 208639 558365
rect 210602 558356 210608 558368
rect 210660 558396 210666 558408
rect 220078 558396 220084 558408
rect 210660 558368 220084 558396
rect 210660 558356 210666 558368
rect 220078 558356 220084 558368
rect 220136 558396 220142 558408
rect 229462 558396 229468 558408
rect 220136 558368 229468 558396
rect 220136 558356 220142 558368
rect 229462 558356 229468 558368
rect 229520 558396 229526 558408
rect 325697 558399 325755 558405
rect 229520 558368 233372 558396
rect 229520 558356 229526 558368
rect 81434 558288 81440 558340
rect 81492 558328 81498 558340
rect 81986 558328 81992 558340
rect 81492 558300 81992 558328
rect 81492 558288 81498 558300
rect 81986 558288 81992 558300
rect 82044 558328 82050 558340
rect 91094 558328 91100 558340
rect 82044 558300 91100 558328
rect 82044 558288 82050 558300
rect 91094 558288 91100 558300
rect 91152 558288 91158 558340
rect 92198 558288 92204 558340
rect 92256 558328 92262 558340
rect 137462 558328 137468 558340
rect 92256 558300 137468 558328
rect 92256 558288 92262 558300
rect 137462 558288 137468 558300
rect 137520 558288 137526 558340
rect 211154 558288 211160 558340
rect 211212 558328 211218 558340
rect 211798 558328 211804 558340
rect 211212 558300 211804 558328
rect 211212 558288 211218 558300
rect 211798 558288 211804 558300
rect 211856 558328 211862 558340
rect 221090 558328 221096 558340
rect 211856 558300 221096 558328
rect 211856 558288 211862 558300
rect 221090 558288 221096 558300
rect 221148 558328 221154 558340
rect 230474 558328 230480 558340
rect 221148 558300 230480 558328
rect 221148 558288 221154 558300
rect 230474 558288 230480 558300
rect 230532 558288 230538 558340
rect 74258 558220 74264 558272
rect 74316 558260 74322 558272
rect 137370 558260 137376 558272
rect 74316 558232 137376 558260
rect 74316 558220 74322 558232
rect 137370 558220 137376 558232
rect 137428 558220 137434 558272
rect 206922 558220 206928 558272
rect 206980 558260 206986 558272
rect 215294 558260 215300 558272
rect 206980 558232 215300 558260
rect 206980 558220 206986 558232
rect 215294 558220 215300 558232
rect 215352 558220 215358 558272
rect 224494 558220 224500 558272
rect 224552 558260 224558 558272
rect 233234 558260 233240 558272
rect 224552 558232 233240 558260
rect 224552 558220 224558 558232
rect 233234 558220 233240 558232
rect 233292 558220 233298 558272
rect 233344 558260 233372 558368
rect 325697 558365 325709 558399
rect 325743 558396 325755 558399
rect 334066 558396 334072 558408
rect 325743 558368 334072 558396
rect 325743 558365 325755 558368
rect 325697 558359 325755 558365
rect 334066 558356 334072 558368
rect 334124 558396 334130 558408
rect 335262 558396 335268 558408
rect 334124 558368 335268 558396
rect 334124 558356 334130 558368
rect 335262 558356 335268 558368
rect 335320 558356 335326 558408
rect 337562 558356 337568 558408
rect 337620 558396 337626 558408
rect 347682 558396 347688 558408
rect 337620 558368 347688 558396
rect 337620 558356 337626 558368
rect 347682 558356 347688 558368
rect 347740 558356 347746 558408
rect 352558 558356 352564 558408
rect 352616 558396 352622 558408
rect 476206 558396 476212 558408
rect 352616 558368 476212 558396
rect 352616 558356 352622 558368
rect 476206 558356 476212 558368
rect 476264 558356 476270 558408
rect 476574 558356 476580 558408
rect 476632 558396 476638 558408
rect 485774 558396 485780 558408
rect 476632 558368 485780 558396
rect 476632 558356 476638 558368
rect 485774 558356 485780 558368
rect 485832 558356 485838 558408
rect 333146 558328 333152 558340
rect 331416 558300 333152 558328
rect 238754 558260 238760 558272
rect 233344 558232 238760 558260
rect 238754 558220 238760 558232
rect 238812 558220 238818 558272
rect 72510 558152 72516 558204
rect 72568 558192 72574 558204
rect 81434 558192 81440 558204
rect 72568 558164 81440 558192
rect 72568 558152 72574 558164
rect 81434 558152 81440 558164
rect 81492 558152 81498 558204
rect 83826 558152 83832 558204
rect 83884 558192 83890 558204
rect 149698 558192 149704 558204
rect 83884 558164 149704 558192
rect 83884 558152 83890 558164
rect 149698 558152 149704 558164
rect 149756 558152 149762 558204
rect 203794 558152 203800 558204
rect 203852 558192 203858 558204
rect 213178 558192 213184 558204
rect 203852 558164 213184 558192
rect 203852 558152 203858 558164
rect 213178 558152 213184 558164
rect 213236 558152 213242 558204
rect 76834 558084 76840 558136
rect 76892 558124 76898 558136
rect 145558 558124 145564 558136
rect 76892 558096 145564 558124
rect 76892 558084 76898 558096
rect 145558 558084 145564 558096
rect 145616 558084 145622 558136
rect 215202 558084 215208 558136
rect 215260 558124 215266 558136
rect 222197 558127 222255 558133
rect 222197 558124 222209 558127
rect 215260 558096 222209 558124
rect 215260 558084 215266 558096
rect 222197 558093 222209 558096
rect 222243 558093 222255 558127
rect 222197 558087 222255 558093
rect 285122 558084 285128 558136
rect 285180 558124 285186 558136
rect 328454 558124 328460 558136
rect 285180 558096 328460 558124
rect 285180 558084 285186 558096
rect 328454 558084 328460 558096
rect 328512 558084 328518 558136
rect 81250 558016 81256 558068
rect 81308 558056 81314 558068
rect 152550 558056 152556 558068
rect 81308 558028 152556 558056
rect 81308 558016 81314 558028
rect 152550 558016 152556 558028
rect 152608 558016 152614 558068
rect 231765 558059 231823 558065
rect 231765 558025 231777 558059
rect 231811 558056 231823 558059
rect 231854 558056 231860 558068
rect 231811 558028 231860 558056
rect 231811 558025 231823 558028
rect 231765 558019 231823 558025
rect 231854 558016 231860 558028
rect 231912 558016 231918 558068
rect 312538 558016 312544 558068
rect 312596 558056 312602 558068
rect 322934 558056 322940 558068
rect 312596 558028 322940 558056
rect 312596 558016 312602 558028
rect 322934 558016 322940 558028
rect 322992 558016 322998 558068
rect 323578 558016 323584 558068
rect 323636 558056 323642 558068
rect 331416 558056 331444 558300
rect 333146 558288 333152 558300
rect 333204 558328 333210 558340
rect 342530 558328 342536 558340
rect 333204 558300 342536 558328
rect 333204 558288 333210 558300
rect 342530 558288 342536 558300
rect 342588 558328 342594 558340
rect 348418 558328 348424 558340
rect 342588 558300 348424 558328
rect 342588 558288 342594 558300
rect 348418 558288 348424 558300
rect 348476 558288 348482 558340
rect 352650 558288 352656 558340
rect 352708 558328 352714 558340
rect 477494 558328 477500 558340
rect 352708 558300 477500 558328
rect 352708 558288 352714 558300
rect 477494 558288 477500 558300
rect 477552 558288 477558 558340
rect 477586 558288 477592 558340
rect 477644 558328 477650 558340
rect 487154 558328 487160 558340
rect 477644 558300 487160 558328
rect 477644 558288 477650 558300
rect 487154 558288 487160 558300
rect 487212 558288 487218 558340
rect 331766 558260 331772 558272
rect 323636 558028 331444 558056
rect 331508 558232 331772 558260
rect 323636 558016 323642 558028
rect 79318 557948 79324 558000
rect 79376 557988 79382 558000
rect 152458 557988 152464 558000
rect 79376 557960 152464 557988
rect 79376 557948 79382 557960
rect 152458 557948 152464 557960
rect 152516 557948 152522 558000
rect 309778 557948 309784 558000
rect 309836 557988 309842 558000
rect 321554 557988 321560 558000
rect 309836 557960 321560 557988
rect 309836 557948 309842 557960
rect 321554 557948 321560 557960
rect 321612 557948 321618 558000
rect 322198 557948 322204 558000
rect 322256 557988 322262 558000
rect 331508 557988 331536 558232
rect 331766 558220 331772 558232
rect 331824 558260 331830 558272
rect 341242 558260 341248 558272
rect 331824 558232 341248 558260
rect 331824 558220 331830 558232
rect 341242 558220 341248 558232
rect 341300 558260 341306 558272
rect 350534 558260 350540 558272
rect 341300 558232 350540 558260
rect 341300 558220 341306 558232
rect 350534 558220 350540 558232
rect 350592 558220 350598 558272
rect 353938 558220 353944 558272
rect 353996 558260 354002 558272
rect 478874 558260 478880 558272
rect 353996 558232 478880 558260
rect 353996 558220 354002 558232
rect 478874 558220 478880 558232
rect 478932 558220 478938 558272
rect 478966 558220 478972 558272
rect 479024 558260 479030 558272
rect 488534 558260 488540 558272
rect 479024 558232 488540 558260
rect 479024 558220 479030 558232
rect 488534 558220 488540 558232
rect 488592 558220 488598 558272
rect 335262 558152 335268 558204
rect 335320 558192 335326 558204
rect 343634 558192 343640 558204
rect 335320 558164 343640 558192
rect 335320 558152 335326 558164
rect 343634 558152 343640 558164
rect 343692 558192 343698 558204
rect 352006 558192 352012 558204
rect 343692 558164 352012 558192
rect 343692 558152 343698 558164
rect 352006 558152 352012 558164
rect 352064 558152 352070 558204
rect 354030 558152 354036 558204
rect 354088 558192 354094 558204
rect 480346 558192 480352 558204
rect 354088 558164 480352 558192
rect 354088 558152 354094 558164
rect 480346 558152 480352 558164
rect 480404 558152 480410 558204
rect 356698 558084 356704 558136
rect 356756 558124 356762 558136
rect 483014 558124 483020 558136
rect 356756 558096 483020 558124
rect 356756 558084 356762 558096
rect 483014 558084 483020 558096
rect 483072 558084 483078 558136
rect 355318 558016 355324 558068
rect 355376 558056 355382 558068
rect 481634 558056 481640 558068
rect 355376 558028 481640 558056
rect 355376 558016 355382 558028
rect 481634 558016 481640 558028
rect 481692 558016 481698 558068
rect 322256 557960 331536 557988
rect 322256 557948 322262 557960
rect 356790 557948 356796 558000
rect 356848 557988 356854 558000
rect 484394 557988 484400 558000
rect 356848 557960 484400 557988
rect 356848 557948 356854 557960
rect 484394 557948 484400 557960
rect 484452 557948 484458 558000
rect 93857 557923 93915 557929
rect 93857 557889 93869 557923
rect 93903 557920 93915 557923
rect 97077 557923 97135 557929
rect 97077 557920 97089 557923
rect 93903 557892 97089 557920
rect 93903 557889 93915 557892
rect 93857 557883 93915 557889
rect 97077 557889 97089 557892
rect 97123 557889 97135 557923
rect 97077 557883 97135 557889
rect 97166 557880 97172 557932
rect 97224 557920 97230 557932
rect 99745 557923 99803 557929
rect 99745 557920 99757 557923
rect 97224 557892 99757 557920
rect 97224 557880 97230 557892
rect 99745 557889 99757 557892
rect 99791 557889 99803 557923
rect 99745 557883 99803 557889
rect 99837 557923 99895 557929
rect 99837 557889 99849 557923
rect 99883 557920 99895 557923
rect 105538 557920 105544 557932
rect 99883 557892 105544 557920
rect 99883 557889 99895 557892
rect 99837 557883 99895 557889
rect 105538 557880 105544 557892
rect 105596 557880 105602 557932
rect 129642 557880 129648 557932
rect 129700 557920 129706 557932
rect 208581 557923 208639 557929
rect 208581 557920 208593 557923
rect 129700 557892 208593 557920
rect 129700 557880 129706 557892
rect 208581 557889 208593 557892
rect 208627 557889 208639 557923
rect 208581 557883 208639 557889
rect 222197 557923 222255 557929
rect 222197 557889 222209 557923
rect 222243 557920 222255 557923
rect 223574 557920 223580 557932
rect 222243 557892 223580 557920
rect 222243 557889 222255 557892
rect 222197 557883 222255 557889
rect 223574 557880 223580 557892
rect 223632 557920 223638 557932
rect 231765 557923 231823 557929
rect 231765 557920 231777 557923
rect 223632 557892 231777 557920
rect 223632 557880 223638 557892
rect 231765 557889 231777 557892
rect 231811 557889 231823 557923
rect 231765 557883 231823 557889
rect 286594 557880 286600 557932
rect 286652 557920 286658 557932
rect 329834 557920 329840 557932
rect 286652 557892 329840 557920
rect 286652 557880 286658 557892
rect 329834 557880 329840 557892
rect 329892 557880 329898 557932
rect 355410 557880 355416 557932
rect 355468 557920 355474 557932
rect 483014 557920 483020 557932
rect 355468 557892 483020 557920
rect 355468 557880 355474 557892
rect 483014 557880 483020 557892
rect 483072 557880 483078 557932
rect 89162 557812 89168 557864
rect 89220 557852 89226 557864
rect 93949 557855 94007 557861
rect 93949 557852 93961 557855
rect 89220 557824 93961 557852
rect 89220 557812 89226 557824
rect 93949 557821 93961 557824
rect 93995 557821 94007 557855
rect 93949 557815 94007 557821
rect 98273 557855 98331 557861
rect 98273 557821 98285 557855
rect 98319 557852 98331 557855
rect 106277 557855 106335 557861
rect 106277 557852 106289 557855
rect 98319 557824 106289 557852
rect 98319 557821 98331 557824
rect 98273 557815 98331 557821
rect 106277 557821 106289 557824
rect 106323 557821 106335 557855
rect 125413 557855 125471 557861
rect 125413 557852 125425 557855
rect 106277 557815 106335 557821
rect 121288 557824 125425 557852
rect 93118 557744 93124 557796
rect 93176 557784 93182 557796
rect 100846 557784 100852 557796
rect 93176 557756 100852 557784
rect 93176 557744 93182 557756
rect 100846 557744 100852 557756
rect 100904 557744 100910 557796
rect 115845 557787 115903 557793
rect 115845 557753 115857 557787
rect 115891 557784 115903 557787
rect 121288 557784 121316 557824
rect 125413 557821 125425 557824
rect 125459 557821 125471 557855
rect 125413 557815 125471 557821
rect 125502 557812 125508 557864
rect 125560 557852 125566 557864
rect 208486 557852 208492 557864
rect 125560 557824 208492 557852
rect 125560 557812 125566 557824
rect 208486 557812 208492 557824
rect 208544 557812 208550 557864
rect 324958 557812 324964 557864
rect 325016 557852 325022 557864
rect 325697 557855 325755 557861
rect 325697 557852 325709 557855
rect 325016 557824 325709 557852
rect 325016 557812 325022 557824
rect 325697 557821 325709 557824
rect 325743 557821 325755 557855
rect 325697 557815 325755 557821
rect 358078 557812 358084 557864
rect 358136 557852 358142 557864
rect 485774 557852 485780 557864
rect 358136 557824 485780 557852
rect 358136 557812 358142 557824
rect 485774 557812 485780 557824
rect 485832 557812 485838 557864
rect 115891 557756 121316 557784
rect 115891 557753 115903 557756
rect 115845 557747 115903 557753
rect 121362 557744 121368 557796
rect 121420 557784 121426 557796
rect 206922 557784 206928 557796
rect 121420 557756 206928 557784
rect 121420 557744 121426 557756
rect 206922 557744 206928 557756
rect 206980 557744 206986 557796
rect 209038 557744 209044 557796
rect 209096 557784 209102 557796
rect 218790 557784 218796 557796
rect 209096 557756 218796 557784
rect 209096 557744 209102 557756
rect 218790 557744 218796 557756
rect 218848 557744 218854 557796
rect 287790 557744 287796 557796
rect 287848 557784 287854 557796
rect 331214 557784 331220 557796
rect 287848 557756 331220 557784
rect 287848 557744 287854 557756
rect 331214 557744 331220 557756
rect 331272 557744 331278 557796
rect 358170 557744 358176 557796
rect 358228 557784 358234 557796
rect 487154 557784 487160 557796
rect 358228 557756 487160 557784
rect 358228 557744 358234 557756
rect 487154 557744 487160 557756
rect 487212 557744 487218 557796
rect 85390 557676 85396 557728
rect 85448 557716 85454 557728
rect 94774 557716 94780 557728
rect 85448 557688 94780 557716
rect 85448 557676 85454 557688
rect 94774 557676 94780 557688
rect 94832 557676 94838 557728
rect 94869 557719 94927 557725
rect 94869 557685 94881 557719
rect 94915 557716 94927 557719
rect 98273 557719 98331 557725
rect 98273 557716 98285 557719
rect 94915 557688 98285 557716
rect 94915 557685 94927 557688
rect 94869 557679 94927 557685
rect 98273 557685 98285 557688
rect 98319 557685 98331 557719
rect 98273 557679 98331 557685
rect 98362 557676 98368 557728
rect 98420 557716 98426 557728
rect 108298 557716 108304 557728
rect 98420 557688 108304 557716
rect 98420 557676 98426 557688
rect 108298 557676 108304 557688
rect 108356 557676 108362 557728
rect 117222 557676 117228 557728
rect 117280 557716 117286 557728
rect 203794 557716 203800 557728
rect 117280 557688 203800 557716
rect 117280 557676 117286 557688
rect 203794 557676 203800 557688
rect 203852 557676 203858 557728
rect 204898 557676 204904 557728
rect 204956 557716 204962 557728
rect 214006 557716 214012 557728
rect 204956 557688 214012 557716
rect 204956 557676 204962 557688
rect 214006 557676 214012 557688
rect 214064 557716 214070 557728
rect 215202 557716 215208 557728
rect 214064 557688 215208 557716
rect 214064 557676 214070 557688
rect 215202 557676 215208 557688
rect 215260 557676 215266 557728
rect 285030 557676 285036 557728
rect 285088 557716 285094 557728
rect 449894 557716 449900 557728
rect 285088 557688 449900 557716
rect 285088 557676 285094 557688
rect 449894 557676 449900 557688
rect 449952 557676 449958 557728
rect 460382 557676 460388 557728
rect 460440 557716 460446 557728
rect 468110 557716 468116 557728
rect 460440 557688 468116 557716
rect 460440 557676 460446 557688
rect 468110 557676 468116 557688
rect 468168 557676 468174 557728
rect 474826 557676 474832 557728
rect 474884 557716 474890 557728
rect 483014 557716 483020 557728
rect 474884 557688 483020 557716
rect 474884 557676 474890 557688
rect 483014 557676 483020 557688
rect 483072 557676 483078 557728
rect 91094 557608 91100 557660
rect 91152 557648 91158 557660
rect 100018 557648 100024 557660
rect 91152 557620 100024 557648
rect 91152 557608 91158 557620
rect 100018 557608 100024 557620
rect 100076 557608 100082 557660
rect 100386 557608 100392 557660
rect 100444 557648 100450 557660
rect 108482 557648 108488 557660
rect 100444 557620 108488 557648
rect 100444 557608 100450 557620
rect 108482 557608 108488 557620
rect 108540 557608 108546 557660
rect 202138 557608 202144 557660
rect 202196 557648 202202 557660
rect 211154 557648 211160 557660
rect 202196 557620 211160 557648
rect 202196 557608 202202 557620
rect 211154 557608 211160 557620
rect 211212 557608 211218 557660
rect 315298 557608 315304 557660
rect 315356 557648 315362 557660
rect 324314 557648 324320 557660
rect 315356 557620 324320 557648
rect 315356 557608 315362 557620
rect 324314 557608 324320 557620
rect 324372 557608 324378 557660
rect 327718 557608 327724 557660
rect 327776 557648 327782 557660
rect 336090 557648 336096 557660
rect 327776 557620 336096 557648
rect 327776 557608 327782 557620
rect 336090 557608 336096 557620
rect 336148 557608 336154 557660
rect 460198 557608 460204 557660
rect 460256 557648 460262 557660
rect 460842 557648 460848 557660
rect 460256 557620 460848 557648
rect 460256 557608 460262 557620
rect 460842 557608 460848 557620
rect 460900 557648 460906 557660
rect 470042 557648 470048 557660
rect 460900 557620 470048 557648
rect 460900 557608 460906 557620
rect 470042 557608 470048 557620
rect 470100 557648 470106 557660
rect 478966 557648 478972 557660
rect 470100 557620 478972 557648
rect 470100 557608 470106 557620
rect 478966 557608 478972 557620
rect 479024 557608 479030 557660
rect 67450 557540 67456 557592
rect 67508 557580 67514 557592
rect 128265 557583 128323 557589
rect 128265 557580 128277 557583
rect 67508 557552 128277 557580
rect 67508 557540 67514 557552
rect 128265 557549 128277 557552
rect 128311 557549 128323 557583
rect 128265 557543 128323 557549
rect 128357 557583 128415 557589
rect 128357 557549 128369 557583
rect 128403 557580 128415 557583
rect 201494 557580 201500 557592
rect 128403 557552 201500 557580
rect 128403 557549 128415 557552
rect 128357 557543 128415 557549
rect 201494 557540 201500 557552
rect 201552 557540 201558 557592
rect 207658 557540 207664 557592
rect 207716 557580 207722 557592
rect 217502 557580 217508 557592
rect 207716 557552 217508 557580
rect 207716 557540 207722 557552
rect 217502 557540 217508 557552
rect 217560 557540 217566 557592
rect 308398 557540 308404 557592
rect 308456 557580 308462 557592
rect 316310 557580 316316 557592
rect 308456 557552 316316 557580
rect 308456 557540 308462 557552
rect 316310 557540 316316 557552
rect 316368 557540 316374 557592
rect 329098 557540 329104 557592
rect 329156 557580 329162 557592
rect 337562 557580 337568 557592
rect 329156 557552 337568 557580
rect 329156 557540 329162 557552
rect 337562 557540 337568 557552
rect 337620 557540 337626 557592
rect 464338 557540 464344 557592
rect 464396 557580 464402 557592
rect 488534 557580 488540 557592
rect 464396 557552 488540 557580
rect 464396 557540 464402 557552
rect 488534 557540 488540 557552
rect 488592 557540 488598 557592
rect 106277 557515 106335 557521
rect 106277 557481 106289 557515
rect 106323 557512 106335 557515
rect 115845 557515 115903 557521
rect 115845 557512 115857 557515
rect 106323 557484 115857 557512
rect 106323 557481 106335 557484
rect 106277 557475 106335 557481
rect 115845 557481 115857 557484
rect 115891 557481 115903 557515
rect 115845 557475 115903 557481
rect 125413 557515 125471 557521
rect 125413 557481 125425 557515
rect 125459 557512 125471 557515
rect 125597 557515 125655 557521
rect 125597 557512 125609 557515
rect 125459 557484 125609 557512
rect 125459 557481 125471 557484
rect 125413 557475 125471 557481
rect 125597 557481 125609 557484
rect 125643 557481 125655 557515
rect 125597 557475 125655 557481
rect 125597 556903 125655 556909
rect 125597 556869 125609 556903
rect 125643 556900 125655 556903
rect 131758 556900 131764 556912
rect 125643 556872 131764 556900
rect 125643 556869 125655 556872
rect 125597 556863 125655 556869
rect 131758 556860 131764 556872
rect 131816 556860 131822 556912
rect 96522 545028 96528 545080
rect 96580 545068 96586 545080
rect 189626 545068 189632 545080
rect 96580 545040 189632 545068
rect 96580 545028 96586 545040
rect 189626 545028 189632 545040
rect 189684 545028 189690 545080
rect 94130 544960 94136 545012
rect 94188 545000 94194 545012
rect 188430 545000 188436 545012
rect 94188 544972 188436 545000
rect 94188 544960 94194 544972
rect 188430 544960 188436 544972
rect 188488 544960 188494 545012
rect 102042 544892 102048 544944
rect 102100 544932 102106 544944
rect 197906 544932 197912 544944
rect 102100 544904 197912 544932
rect 102100 544892 102106 544904
rect 197906 544892 197912 544904
rect 197964 544892 197970 544944
rect 92106 544824 92112 544876
rect 92164 544864 92170 544876
rect 188522 544864 188528 544876
rect 92164 544836 188528 544864
rect 92164 544824 92170 544836
rect 188522 544824 188528 544836
rect 188580 544824 188586 544876
rect 89990 544756 89996 544808
rect 90048 544796 90054 544808
rect 188614 544796 188620 544808
rect 90048 544768 188620 544796
rect 90048 544756 90054 544768
rect 188614 544756 188620 544768
rect 188672 544756 188678 544808
rect 106182 544688 106188 544740
rect 106240 544728 106246 544740
rect 206186 544728 206192 544740
rect 106240 544700 206192 544728
rect 106240 544688 106246 544700
rect 206186 544688 206192 544700
rect 206244 544688 206250 544740
rect 87966 544620 87972 544672
rect 88024 544660 88030 544672
rect 188706 544660 188712 544672
rect 88024 544632 188712 544660
rect 88024 544620 88030 544632
rect 188706 544620 188712 544632
rect 188764 544620 188770 544672
rect 110322 544552 110328 544604
rect 110380 544592 110386 544604
rect 212442 544592 212448 544604
rect 110380 544564 212448 544592
rect 110380 544552 110386 544564
rect 212442 544552 212448 544564
rect 212500 544552 212506 544604
rect 85850 544484 85856 544536
rect 85908 544524 85914 544536
rect 188798 544524 188804 544536
rect 85908 544496 188804 544524
rect 85908 544484 85914 544496
rect 188798 544484 188804 544496
rect 188856 544484 188862 544536
rect 83826 544416 83832 544468
rect 83884 544456 83890 544468
rect 188890 544456 188896 544468
rect 83884 544428 188896 544456
rect 83884 544416 83890 544428
rect 188890 544416 188896 544428
rect 188948 544416 188954 544468
rect 81710 544348 81716 544400
rect 81768 544388 81774 544400
rect 195974 544388 195980 544400
rect 81768 544360 195980 544388
rect 81768 544348 81774 544360
rect 195974 544348 195980 544360
rect 196032 544348 196038 544400
rect 86770 544280 86776 544332
rect 86828 544320 86834 544332
rect 173066 544320 173072 544332
rect 86828 544292 173072 544320
rect 86828 544280 86834 544292
rect 173066 544280 173072 544292
rect 173124 544280 173130 544332
rect 88242 544212 88248 544264
rect 88300 544252 88306 544264
rect 175090 544252 175096 544264
rect 88300 544224 175096 544252
rect 88300 544212 88306 544224
rect 175090 544212 175096 544224
rect 175148 544212 175154 544264
rect 85482 544144 85488 544196
rect 85540 544184 85546 544196
rect 168834 544184 168840 544196
rect 85540 544156 168840 544184
rect 85540 544144 85546 544156
rect 168834 544144 168840 544156
rect 168892 544144 168898 544196
rect 86862 544076 86868 544128
rect 86920 544116 86926 544128
rect 170950 544116 170956 544128
rect 86920 544088 170956 544116
rect 86920 544076 86926 544088
rect 170950 544076 170956 544088
rect 171008 544076 171014 544128
rect 82722 544008 82728 544060
rect 82780 544048 82786 544060
rect 164694 544048 164700 544060
rect 82780 544020 164700 544048
rect 82780 544008 82786 544020
rect 164694 544008 164700 544020
rect 164752 544008 164758 544060
rect 73062 543940 73068 543992
rect 73120 543980 73126 543992
rect 148134 543980 148140 543992
rect 73120 543952 148140 543980
rect 73120 543940 73126 543952
rect 148134 543940 148140 543952
rect 148192 543940 148198 543992
rect 57882 543872 57888 543924
rect 57940 543912 57946 543924
rect 112806 543912 112812 543924
rect 57940 543884 112812 543912
rect 57940 543872 57946 543884
rect 112806 543872 112812 543884
rect 112864 543872 112870 543924
rect 57790 543804 57796 543856
rect 57848 543844 57854 543856
rect 110782 543844 110788 543856
rect 57848 543816 110788 543844
rect 57848 543804 57854 543816
rect 110782 543804 110788 543816
rect 110840 543804 110846 543856
rect 220722 543736 220728 543788
rect 220780 543736 220786 543788
rect 71682 543668 71688 543720
rect 71740 543708 71746 543720
rect 75454 543708 75460 543720
rect 71740 543680 75460 543708
rect 71740 543668 71746 543680
rect 75454 543668 75460 543680
rect 75512 543668 75518 543720
rect 75822 543668 75828 543720
rect 75880 543708 75886 543720
rect 145469 543711 145527 543717
rect 145469 543708 145481 543711
rect 75880 543680 145481 543708
rect 75880 543668 75886 543680
rect 145469 543677 145481 543680
rect 145515 543677 145527 543711
rect 145469 543671 145527 543677
rect 145558 543668 145564 543720
rect 145616 543708 145622 543720
rect 152461 543711 152519 543717
rect 152461 543708 152473 543711
rect 145616 543680 152473 543708
rect 145616 543668 145622 543680
rect 152461 543677 152473 543680
rect 152507 543677 152519 543711
rect 152461 543671 152519 543677
rect 152550 543668 152556 543720
rect 152608 543708 152614 543720
rect 162670 543708 162676 543720
rect 152608 543680 162676 543708
rect 152608 543668 152614 543680
rect 162670 543668 162676 543680
rect 162728 543668 162734 543720
rect 205542 543668 205548 543720
rect 205600 543708 205606 543720
rect 218698 543708 218704 543720
rect 205600 543680 218704 543708
rect 205600 543668 205606 543680
rect 218698 543668 218704 543680
rect 218756 543668 218762 543720
rect 220538 543668 220544 543720
rect 220596 543708 220602 543720
rect 220740 543708 220768 543736
rect 220596 543680 220768 543708
rect 220596 543668 220602 543680
rect 229002 543668 229008 543720
rect 229060 543708 229066 543720
rect 260190 543708 260196 543720
rect 229060 543680 260196 543708
rect 229060 543668 229066 543680
rect 260190 543668 260196 543680
rect 260248 543668 260254 543720
rect 70302 543600 70308 543652
rect 70360 543640 70366 543652
rect 73430 543640 73436 543652
rect 70360 543612 73436 543640
rect 70360 543600 70366 543612
rect 73430 543600 73436 543612
rect 73488 543600 73494 543652
rect 78582 543600 78588 543652
rect 78640 543640 78646 543652
rect 156414 543640 156420 543652
rect 78640 543612 156420 543640
rect 78640 543600 78646 543612
rect 156414 543600 156420 543612
rect 156472 543600 156478 543652
rect 206922 543600 206928 543652
rect 206980 543640 206986 543652
rect 220722 543640 220728 543652
rect 206980 543612 220728 543640
rect 206980 543600 206986 543612
rect 220722 543600 220728 543612
rect 220780 543600 220786 543652
rect 227622 543600 227628 543652
rect 227680 543640 227686 543652
rect 258074 543640 258080 543652
rect 227680 543612 258080 543640
rect 227680 543600 227686 543612
rect 258074 543600 258080 543612
rect 258132 543600 258138 543652
rect 61010 543532 61016 543584
rect 61068 543572 61074 543584
rect 62022 543572 62028 543584
rect 61068 543544 62028 543572
rect 61068 543532 61074 543544
rect 62022 543532 62028 543544
rect 62080 543532 62086 543584
rect 65150 543532 65156 543584
rect 65208 543572 65214 543584
rect 66162 543572 66168 543584
rect 65208 543544 66168 543572
rect 65208 543532 65214 543544
rect 66162 543532 66168 543544
rect 66220 543532 66226 543584
rect 70210 543532 70216 543584
rect 70268 543572 70274 543584
rect 71314 543572 71320 543584
rect 70268 543544 71320 543572
rect 70268 543532 70274 543544
rect 71314 543532 71320 543544
rect 71372 543532 71378 543584
rect 79870 543532 79876 543584
rect 79928 543572 79934 543584
rect 152369 543575 152427 543581
rect 152369 543572 152381 543575
rect 79928 543544 152381 543572
rect 79928 543532 79934 543544
rect 152369 543541 152381 543544
rect 152415 543541 152427 543575
rect 152369 543535 152427 543541
rect 152458 543532 152464 543584
rect 152516 543572 152522 543584
rect 158530 543572 158536 543584
rect 152516 543544 158536 543572
rect 152516 543532 152522 543544
rect 158530 543532 158536 543544
rect 158588 543532 158594 543584
rect 208302 543532 208308 543584
rect 208360 543572 208366 543584
rect 222838 543572 222844 543584
rect 208360 543544 222844 543572
rect 208360 543532 208366 543544
rect 222838 543532 222844 543544
rect 222896 543532 222902 543584
rect 230382 543532 230388 543584
rect 230440 543572 230446 543584
rect 262214 543572 262220 543584
rect 230440 543544 262220 543572
rect 230440 543532 230446 543544
rect 262214 543532 262220 543544
rect 262272 543532 262278 543584
rect 57422 543464 57428 543516
rect 57480 543504 57486 543516
rect 102502 543504 102508 543516
rect 57480 543476 102508 543504
rect 57480 543464 57486 543476
rect 102502 543464 102508 543476
rect 102560 543464 102566 543516
rect 127342 543464 127348 543516
rect 127400 543504 127406 543516
rect 209038 543504 209044 543516
rect 127400 543476 209044 543504
rect 127400 543464 127406 543476
rect 209038 543464 209044 543476
rect 209096 543464 209102 543516
rect 209682 543464 209688 543516
rect 209740 543504 209746 543516
rect 224862 543504 224868 543516
rect 209740 543476 224868 543504
rect 209740 543464 209746 543476
rect 224862 543464 224868 543476
rect 224920 543464 224926 543516
rect 231762 543464 231768 543516
rect 231820 543504 231826 543516
rect 264330 543504 264336 543516
rect 231820 543476 264336 543504
rect 231820 543464 231826 543476
rect 264330 543464 264336 543476
rect 264388 543464 264394 543516
rect 57514 543396 57520 543448
rect 57572 543436 57578 543448
rect 104526 543436 104532 543448
rect 57572 543408 104532 543436
rect 57572 543396 57578 543408
rect 104526 543396 104532 543408
rect 104584 543396 104590 543448
rect 123202 543396 123208 543448
rect 123260 543436 123266 543448
rect 207658 543436 207664 543448
rect 123260 543408 207664 543436
rect 123260 543396 123266 543408
rect 207658 543396 207664 543408
rect 207716 543396 207722 543448
rect 211062 543396 211068 543448
rect 211120 543436 211126 543448
rect 226978 543436 226984 543448
rect 211120 543408 226984 543436
rect 211120 543396 211126 543408
rect 226978 543396 226984 543408
rect 227036 543396 227042 543448
rect 233142 543396 233148 543448
rect 233200 543436 233206 543448
rect 266446 543436 266452 543448
rect 233200 543408 266452 543436
rect 233200 543396 233206 543408
rect 266446 543396 266452 543408
rect 266504 543396 266510 543448
rect 57606 543328 57612 543380
rect 57664 543368 57670 543380
rect 106642 543368 106648 543380
rect 57664 543340 106648 543368
rect 57664 543328 57670 543340
rect 106642 543328 106648 543340
rect 106700 543328 106706 543380
rect 119062 543328 119068 543380
rect 119120 543368 119126 543380
rect 204898 543368 204904 543380
rect 119120 543340 204904 543368
rect 119120 543328 119126 543340
rect 204898 543328 204904 543340
rect 204956 543328 204962 543380
rect 212350 543328 212356 543380
rect 212408 543368 212414 543380
rect 231118 543368 231124 543380
rect 212408 543340 231124 543368
rect 212408 543328 212414 543340
rect 231118 543328 231124 543340
rect 231176 543328 231182 543380
rect 233050 543328 233056 543380
rect 233108 543368 233114 543380
rect 268470 543368 268476 543380
rect 233108 543340 268476 543368
rect 233108 543328 233114 543340
rect 268470 543328 268476 543340
rect 268528 543328 268534 543380
rect 91002 543260 91008 543312
rect 91060 543300 91066 543312
rect 179230 543300 179236 543312
rect 91060 543272 179236 543300
rect 91060 543260 91066 543272
rect 179230 543260 179236 543272
rect 179288 543260 179294 543312
rect 215202 543260 215208 543312
rect 215260 543300 215266 543312
rect 235258 543300 235264 543312
rect 215260 543272 235264 543300
rect 215260 543260 215266 543272
rect 235258 543260 235264 543272
rect 235316 543260 235322 543312
rect 235902 543260 235908 543312
rect 235960 543300 235966 543312
rect 272610 543300 272616 543312
rect 235960 543272 272616 543300
rect 235960 543260 235966 543272
rect 272610 543260 272616 543272
rect 272668 543260 272674 543312
rect 57698 543192 57704 543244
rect 57756 543232 57762 543244
rect 108666 543232 108672 543244
rect 57756 543204 108672 543232
rect 57756 543192 57762 543204
rect 108666 543192 108672 543204
rect 108724 543192 108730 543244
rect 114922 543192 114928 543244
rect 114980 543232 114986 543244
rect 202138 543232 202144 543244
rect 114980 543204 202144 543232
rect 114980 543192 114986 543204
rect 202138 543192 202144 543204
rect 202196 543192 202202 543244
rect 216490 543192 216496 543244
rect 216548 543232 216554 543244
rect 216769 543235 216827 543241
rect 216548 543204 216720 543232
rect 216548 543192 216554 543204
rect 93670 543124 93676 543176
rect 93728 543164 93734 543176
rect 183370 543164 183376 543176
rect 93728 543136 183376 543164
rect 93728 543124 93734 543136
rect 183370 543124 183376 543136
rect 183428 543124 183434 543176
rect 204162 543124 204168 543176
rect 204220 543164 204226 543176
rect 216582 543164 216588 543176
rect 204220 543136 216588 543164
rect 204220 543124 204226 543136
rect 216582 543124 216588 543136
rect 216640 543124 216646 543176
rect 216692 543164 216720 543204
rect 216769 543201 216781 543235
rect 216815 543232 216827 543235
rect 229094 543232 229100 543244
rect 216815 543204 229100 543232
rect 216815 543201 216827 543204
rect 216769 543195 216827 543201
rect 229094 543192 229100 543204
rect 229152 543192 229158 543244
rect 234522 543192 234528 543244
rect 234580 543232 234586 543244
rect 270586 543232 270592 543244
rect 234580 543204 270592 543232
rect 234580 543192 234586 543204
rect 270586 543192 270592 543204
rect 270644 543192 270650 543244
rect 237374 543164 237380 543176
rect 216692 543136 237380 543164
rect 237374 543124 237380 543136
rect 237432 543124 237438 543176
rect 238662 543124 238668 543176
rect 238720 543164 238726 543176
rect 276750 543164 276756 543176
rect 238720 543136 276756 543164
rect 238720 543124 238726 543136
rect 276750 543124 276756 543136
rect 276808 543124 276814 543176
rect 57238 543056 57244 543108
rect 57296 543096 57302 543108
rect 79686 543096 79692 543108
rect 57296 543068 79692 543096
rect 57296 543056 57302 543068
rect 79686 543056 79692 543068
rect 79744 543056 79750 543108
rect 95050 543056 95056 543108
rect 95108 543096 95114 543108
rect 187510 543096 187516 543108
rect 95108 543068 187516 543096
rect 95108 543056 95114 543068
rect 187510 543056 187516 543068
rect 187568 543056 187574 543108
rect 213822 543056 213828 543108
rect 213880 543096 213886 543108
rect 233234 543096 233240 543108
rect 213880 543068 233240 543096
rect 213880 543056 213886 543068
rect 233234 543056 233240 543068
rect 233292 543056 233298 543108
rect 237282 543056 237288 543108
rect 237340 543096 237346 543108
rect 274726 543096 274732 543108
rect 237340 543068 274732 543096
rect 237340 543056 237346 543068
rect 274726 543056 274732 543068
rect 274784 543056 274790 543108
rect 67542 542988 67548 543040
rect 67600 543028 67606 543040
rect 98362 543028 98368 543040
rect 67600 543000 98368 543028
rect 67600 542988 67606 543000
rect 98362 542988 98368 543000
rect 98420 542988 98426 543040
rect 99282 542988 99288 543040
rect 99340 543028 99346 543040
rect 193766 543028 193772 543040
rect 99340 543000 193772 543028
rect 99340 542988 99346 543000
rect 193766 542988 193772 543000
rect 193824 542988 193830 543040
rect 202782 542988 202788 543040
rect 202840 543028 202846 543040
rect 214558 543028 214564 543040
rect 202840 543000 214564 543028
rect 202840 542988 202846 543000
rect 214558 542988 214564 543000
rect 214616 542988 214622 543040
rect 217962 542988 217968 543040
rect 218020 543028 218026 543040
rect 239398 543028 239404 543040
rect 218020 543000 239404 543028
rect 218020 542988 218026 543000
rect 239398 542988 239404 543000
rect 239456 542988 239462 543040
rect 240042 542988 240048 543040
rect 240100 543028 240106 543040
rect 278866 543028 278872 543040
rect 240100 543000 278872 543028
rect 240100 542988 240106 543000
rect 278866 542988 278872 543000
rect 278924 542988 278930 543040
rect 57330 542920 57336 542972
rect 57388 542960 57394 542972
rect 100386 542960 100392 542972
rect 57388 542932 100392 542960
rect 57388 542920 57394 542932
rect 100386 542920 100392 542932
rect 100444 542920 100450 542972
rect 108298 542920 108304 542972
rect 108356 542960 108362 542972
rect 143994 542960 144000 542972
rect 108356 542932 144000 542960
rect 108356 542920 108362 542932
rect 143994 542920 144000 542932
rect 144052 542920 144058 542972
rect 144178 542920 144184 542972
rect 144236 542960 144242 542972
rect 204162 542960 204168 542972
rect 144236 542932 204168 542960
rect 144236 542920 144242 542932
rect 204162 542920 204168 542932
rect 204220 542920 204226 542972
rect 210970 542920 210976 542972
rect 211028 542960 211034 542972
rect 216769 542963 216827 542969
rect 216769 542960 216781 542963
rect 211028 542932 216781 542960
rect 211028 542920 211034 542932
rect 216769 542929 216781 542932
rect 216815 542929 216827 542963
rect 216769 542923 216827 542929
rect 226150 542920 226156 542972
rect 226208 542960 226214 542972
rect 256050 542960 256056 542972
rect 226208 542932 256056 542960
rect 226208 542920 226214 542932
rect 256050 542920 256056 542932
rect 256108 542920 256114 542972
rect 105538 542852 105544 542904
rect 105596 542892 105602 542904
rect 139854 542892 139860 542904
rect 105596 542864 139860 542892
rect 105596 542852 105602 542864
rect 139854 542852 139860 542864
rect 139912 542852 139918 542904
rect 140130 542852 140136 542904
rect 140188 542892 140194 542904
rect 195882 542892 195888 542904
rect 140188 542864 195888 542892
rect 140188 542852 140194 542864
rect 195882 542852 195888 542864
rect 195940 542852 195946 542904
rect 226242 542852 226248 542904
rect 226300 542892 226306 542904
rect 253934 542892 253940 542904
rect 226300 542864 253940 542892
rect 226300 542852 226306 542864
rect 253934 542852 253940 542864
rect 253992 542852 253998 542904
rect 102778 542784 102784 542836
rect 102836 542824 102842 542836
rect 135714 542824 135720 542836
rect 102836 542796 135720 542824
rect 102836 542784 102842 542796
rect 135714 542784 135720 542796
rect 135772 542784 135778 542836
rect 137278 542784 137284 542836
rect 137336 542824 137342 542836
rect 137336 542796 137876 542824
rect 137336 542784 137342 542796
rect 104158 542716 104164 542768
rect 104216 542756 104222 542768
rect 137738 542756 137744 542768
rect 104216 542728 137744 542756
rect 104216 542716 104222 542728
rect 137738 542716 137744 542728
rect 137796 542716 137802 542768
rect 137848 542756 137876 542796
rect 138658 542784 138664 542836
rect 138716 542824 138722 542836
rect 191742 542824 191748 542836
rect 138716 542796 191748 542824
rect 138716 542784 138722 542796
rect 191742 542784 191748 542796
rect 191800 542784 191806 542836
rect 223482 542784 223488 542836
rect 223540 542824 223546 542836
rect 249794 542824 249800 542836
rect 223540 542796 249800 542824
rect 223540 542784 223546 542796
rect 249794 542784 249800 542796
rect 249852 542784 249858 542836
rect 185486 542756 185492 542768
rect 137848 542728 185492 542756
rect 185486 542716 185492 542728
rect 185544 542716 185550 542768
rect 224678 542716 224684 542768
rect 224736 542756 224742 542768
rect 251910 542756 251916 542768
rect 224736 542728 251916 542756
rect 224736 542716 224742 542728
rect 251910 542716 251916 542728
rect 251968 542716 251974 542768
rect 100018 542648 100024 542700
rect 100076 542688 100082 542700
rect 131482 542688 131488 542700
rect 100076 542660 131488 542688
rect 100076 542648 100082 542660
rect 131482 542648 131488 542660
rect 131540 542648 131546 542700
rect 131758 542648 131764 542700
rect 131816 542688 131822 542700
rect 177206 542688 177212 542700
rect 131816 542660 177212 542688
rect 131816 542648 131822 542660
rect 177206 542648 177212 542660
rect 177264 542648 177270 542700
rect 220538 542648 220544 542700
rect 220596 542688 220602 542700
rect 245654 542688 245660 542700
rect 220596 542660 245660 542688
rect 220596 542648 220602 542660
rect 245654 542648 245660 542660
rect 245712 542648 245718 542700
rect 101398 542580 101404 542632
rect 101456 542620 101462 542632
rect 133598 542620 133604 542632
rect 101456 542592 133604 542620
rect 101456 542580 101462 542592
rect 133598 542580 133604 542592
rect 133656 542580 133662 542632
rect 137462 542580 137468 542632
rect 137520 542620 137526 542632
rect 181346 542620 181352 542632
rect 137520 542592 181352 542620
rect 137520 542580 137526 542592
rect 181346 542580 181352 542592
rect 181404 542580 181410 542632
rect 222102 542580 222108 542632
rect 222160 542620 222166 542632
rect 247770 542620 247776 542632
rect 222160 542592 247776 542620
rect 222160 542580 222166 542592
rect 247770 542580 247776 542592
rect 247828 542580 247834 542632
rect 108482 542512 108488 542564
rect 108540 542552 108546 542564
rect 146018 542552 146024 542564
rect 108540 542524 146024 542552
rect 108540 542512 108546 542524
rect 146018 542512 146024 542524
rect 146076 542512 146082 542564
rect 152274 542552 152280 542564
rect 146956 542524 152280 542552
rect 106918 542444 106924 542496
rect 106976 542484 106982 542496
rect 141878 542484 141884 542496
rect 106976 542456 141884 542484
rect 106976 542444 106982 542456
rect 141878 542444 141884 542456
rect 141936 542444 141942 542496
rect 145469 542487 145527 542493
rect 145469 542453 145481 542487
rect 145515 542484 145527 542487
rect 146956 542484 146984 542524
rect 152274 542512 152280 542524
rect 152332 542512 152338 542564
rect 152461 542555 152519 542561
rect 152461 542521 152473 542555
rect 152507 542552 152519 542555
rect 154390 542552 154396 542564
rect 152507 542524 154396 542552
rect 152507 542521 152519 542524
rect 152461 542515 152519 542521
rect 154390 542512 154396 542524
rect 154448 542512 154454 542564
rect 166810 542552 166816 542564
rect 156616 542524 166816 542552
rect 145515 542456 146984 542484
rect 145515 542453 145527 542456
rect 145469 542447 145527 542453
rect 149698 542444 149704 542496
rect 149756 542484 149762 542496
rect 156616 542484 156644 542524
rect 166810 542512 166816 542524
rect 166868 542512 166874 542564
rect 217870 542512 217876 542564
rect 217928 542552 217934 542564
rect 241514 542552 241520 542564
rect 217928 542524 241520 542552
rect 217928 542512 217934 542524
rect 241514 542512 241520 542524
rect 241572 542512 241578 542564
rect 149756 542456 156644 542484
rect 149756 542444 149762 542456
rect 219342 542444 219348 542496
rect 219400 542484 219406 542496
rect 243538 542484 243544 542496
rect 219400 542456 243544 542484
rect 219400 542444 219406 542456
rect 243538 542444 243544 542456
rect 243596 542444 243602 542496
rect 137370 542376 137376 542428
rect 137428 542416 137434 542428
rect 150158 542416 150164 542428
rect 137428 542388 150164 542416
rect 137428 542376 137434 542388
rect 150158 542376 150164 542388
rect 150216 542376 150222 542428
rect 152369 542419 152427 542425
rect 152369 542385 152381 542419
rect 152415 542416 152427 542419
rect 160554 542416 160560 542428
rect 152415 542388 160560 542416
rect 152415 542385 152427 542388
rect 152369 542379 152427 542385
rect 160554 542376 160560 542388
rect 160612 542376 160618 542428
rect 282270 538296 282276 538348
rect 282328 538336 282334 538348
rect 367094 538336 367100 538348
rect 282328 538308 367100 538336
rect 282328 538296 282334 538308
rect 367094 538296 367100 538308
rect 367152 538296 367158 538348
rect 282822 538228 282828 538280
rect 282880 538268 282886 538280
rect 368474 538268 368480 538280
rect 282880 538240 368480 538268
rect 282880 538228 282886 538240
rect 368474 538228 368480 538240
rect 368532 538228 368538 538280
rect 282822 536800 282828 536852
rect 282880 536840 282886 536852
rect 369854 536840 369860 536852
rect 282880 536812 369860 536840
rect 282880 536800 282886 536812
rect 369854 536800 369860 536812
rect 369912 536800 369918 536852
rect 282822 535440 282828 535492
rect 282880 535480 282886 535492
rect 371234 535480 371240 535492
rect 282880 535452 371240 535480
rect 282880 535440 282886 535452
rect 371234 535440 371240 535452
rect 371292 535440 371298 535492
rect 281718 534148 281724 534200
rect 281776 534188 281782 534200
rect 372614 534188 372620 534200
rect 281776 534160 372620 534188
rect 281776 534148 281782 534160
rect 372614 534148 372620 534160
rect 372672 534148 372678 534200
rect 282086 534080 282092 534132
rect 282144 534120 282150 534132
rect 373994 534120 374000 534132
rect 282144 534092 374000 534120
rect 282144 534080 282150 534092
rect 373994 534080 374000 534092
rect 374052 534080 374058 534132
rect 282086 532720 282092 532772
rect 282144 532760 282150 532772
rect 375374 532760 375380 532772
rect 282144 532732 375380 532760
rect 282144 532720 282150 532732
rect 375374 532720 375380 532732
rect 375432 532720 375438 532772
rect 282270 531360 282276 531412
rect 282328 531400 282334 531412
rect 375466 531400 375472 531412
rect 282328 531372 375472 531400
rect 282328 531360 282334 531372
rect 375466 531360 375472 531372
rect 375524 531360 375530 531412
rect 282822 531292 282828 531344
rect 282880 531332 282886 531344
rect 376754 531332 376760 531344
rect 282880 531304 376760 531332
rect 282880 531292 282886 531304
rect 376754 531292 376760 531304
rect 376812 531292 376818 531344
rect 282822 529932 282828 529984
rect 282880 529972 282886 529984
rect 378226 529972 378232 529984
rect 282880 529944 378232 529972
rect 282880 529932 282886 529944
rect 378226 529932 378232 529944
rect 378284 529932 378290 529984
rect 282822 528572 282828 528624
rect 282880 528612 282886 528624
rect 379606 528612 379612 528624
rect 282880 528584 379612 528612
rect 282880 528572 282886 528584
rect 379606 528572 379612 528584
rect 379664 528572 379670 528624
rect 282822 527212 282828 527264
rect 282880 527252 282886 527264
rect 376018 527252 376024 527264
rect 282880 527224 376024 527252
rect 282880 527212 282886 527224
rect 376018 527212 376024 527224
rect 376076 527212 376082 527264
rect 282270 527144 282276 527196
rect 282328 527184 282334 527196
rect 380986 527184 380992 527196
rect 282328 527156 380992 527184
rect 282328 527144 282334 527156
rect 380986 527144 380992 527156
rect 381044 527144 381050 527196
rect 281902 525784 281908 525836
rect 281960 525824 281966 525836
rect 374638 525824 374644 525836
rect 281960 525796 374644 525824
rect 281960 525784 281966 525796
rect 374638 525784 374644 525796
rect 374696 525784 374702 525836
rect 282822 524424 282828 524476
rect 282880 524464 282886 524476
rect 371878 524464 371884 524476
rect 282880 524436 371884 524464
rect 282880 524424 282886 524436
rect 371878 524424 371884 524436
rect 371936 524424 371942 524476
rect 282822 523064 282828 523116
rect 282880 523104 282886 523116
rect 354122 523104 354128 523116
rect 282880 523076 354128 523104
rect 282880 523064 282886 523076
rect 354122 523064 354128 523076
rect 354180 523064 354186 523116
rect 282362 522996 282368 523048
rect 282420 523036 282426 523048
rect 367738 523036 367744 523048
rect 282420 523008 367744 523036
rect 282420 522996 282426 523008
rect 367738 522996 367744 523008
rect 367796 522996 367802 523048
rect 282822 521636 282828 521688
rect 282880 521676 282886 521688
rect 387886 521676 387892 521688
rect 282880 521648 387892 521676
rect 282880 521636 282886 521648
rect 387886 521636 387892 521648
rect 387944 521636 387950 521688
rect 282822 520276 282828 520328
rect 282880 520316 282886 520328
rect 390646 520316 390652 520328
rect 282880 520288 390652 520316
rect 282880 520276 282886 520288
rect 390646 520276 390652 520288
rect 390704 520276 390710 520328
rect 281718 519052 281724 519104
rect 281776 519092 281782 519104
rect 283742 519092 283748 519104
rect 281776 519064 283748 519092
rect 281776 519052 281782 519064
rect 283742 519052 283748 519064
rect 283800 519052 283806 519104
rect 282086 517488 282092 517540
rect 282144 517528 282150 517540
rect 392026 517528 392032 517540
rect 282144 517500 392032 517528
rect 282144 517488 282150 517500
rect 392026 517488 392032 517500
rect 392084 517488 392090 517540
rect 282270 516196 282276 516248
rect 282328 516236 282334 516248
rect 387058 516236 387064 516248
rect 282328 516208 387064 516236
rect 282328 516196 282334 516208
rect 387058 516196 387064 516208
rect 387116 516196 387122 516248
rect 282822 516128 282828 516180
rect 282880 516168 282886 516180
rect 419534 516168 419540 516180
rect 282880 516140 419540 516168
rect 282880 516128 282886 516140
rect 419534 516128 419540 516140
rect 419592 516128 419598 516180
rect 282822 514768 282828 514820
rect 282880 514808 282886 514820
rect 385678 514808 385684 514820
rect 282880 514780 385684 514808
rect 282880 514768 282886 514780
rect 385678 514768 385684 514780
rect 385736 514768 385742 514820
rect 282270 513340 282276 513392
rect 282328 513380 282334 513392
rect 419626 513380 419632 513392
rect 282328 513352 419632 513380
rect 282328 513340 282334 513352
rect 419626 513340 419632 513352
rect 419684 513340 419690 513392
rect 282730 512048 282736 512100
rect 282788 512088 282794 512100
rect 385770 512088 385776 512100
rect 282788 512060 385776 512088
rect 282788 512048 282794 512060
rect 385770 512048 385776 512060
rect 385828 512048 385834 512100
rect 282822 511980 282828 512032
rect 282880 512020 282886 512032
rect 419718 512020 419724 512032
rect 282880 511992 419724 512020
rect 282880 511980 282886 511992
rect 419718 511980 419724 511992
rect 419776 511980 419782 512032
rect 281718 510620 281724 510672
rect 281776 510660 281782 510672
rect 384298 510660 384304 510672
rect 281776 510632 384304 510660
rect 281776 510620 281782 510632
rect 384298 510620 384304 510632
rect 384356 510620 384362 510672
rect 282270 509260 282276 509312
rect 282328 509300 282334 509312
rect 419810 509300 419816 509312
rect 282328 509272 419816 509300
rect 282328 509260 282334 509272
rect 419810 509260 419816 509272
rect 419868 509260 419874 509312
rect 282546 507900 282552 507952
rect 282604 507940 282610 507952
rect 382918 507940 382924 507952
rect 282604 507912 382924 507940
rect 282604 507900 282610 507912
rect 382918 507900 382924 507912
rect 382976 507900 382982 507952
rect 282822 507832 282828 507884
rect 282880 507872 282886 507884
rect 419902 507872 419908 507884
rect 282880 507844 419908 507872
rect 282880 507832 282886 507844
rect 419902 507832 419908 507844
rect 419960 507832 419966 507884
rect 282086 506472 282092 506524
rect 282144 506512 282150 506524
rect 383010 506512 383016 506524
rect 282144 506484 383016 506512
rect 282144 506472 282150 506484
rect 383010 506472 383016 506484
rect 383068 506472 383074 506524
rect 282822 505180 282828 505232
rect 282880 505220 282886 505232
rect 383102 505220 383108 505232
rect 282880 505192 383108 505220
rect 282880 505180 282886 505192
rect 383102 505180 383108 505192
rect 383160 505180 383166 505232
rect 282730 505112 282736 505164
rect 282788 505152 282794 505164
rect 419994 505152 420000 505164
rect 282788 505124 420000 505152
rect 282788 505112 282794 505124
rect 419994 505112 420000 505124
rect 420052 505112 420058 505164
rect 282822 503684 282828 503736
rect 282880 503724 282886 503736
rect 420086 503724 420092 503736
rect 282880 503696 420092 503724
rect 282880 503684 282886 503696
rect 420086 503684 420092 503696
rect 420144 503684 420150 503736
rect 282822 502324 282828 502376
rect 282880 502364 282886 502376
rect 383194 502364 383200 502376
rect 282880 502336 383200 502364
rect 282880 502324 282886 502336
rect 383194 502324 383200 502336
rect 383252 502324 383258 502376
rect 282822 501032 282828 501084
rect 282880 501072 282886 501084
rect 378778 501072 378784 501084
rect 282880 501044 378784 501072
rect 282880 501032 282886 501044
rect 378778 501032 378784 501044
rect 378836 501032 378842 501084
rect 282270 500964 282276 501016
rect 282328 501004 282334 501016
rect 410518 501004 410524 501016
rect 282328 500976 410524 501004
rect 282328 500964 282334 500976
rect 410518 500964 410524 500976
rect 410576 500964 410582 501016
rect 282822 498176 282828 498228
rect 282880 498216 282886 498228
rect 283926 498216 283932 498228
rect 282880 498188 283932 498216
rect 282880 498176 282886 498188
rect 283926 498176 283932 498188
rect 283984 498176 283990 498228
rect 282822 496816 282828 496868
rect 282880 496856 282886 496868
rect 416314 496856 416320 496868
rect 282880 496828 416320 496856
rect 282880 496816 282886 496828
rect 416314 496816 416320 496828
rect 416372 496816 416378 496868
rect 281902 495456 281908 495508
rect 281960 495496 281966 495508
rect 498838 495496 498844 495508
rect 281960 495468 498844 495496
rect 281960 495456 281966 495468
rect 498838 495456 498844 495468
rect 498896 495456 498902 495508
rect 282822 494028 282828 494080
rect 282880 494068 282886 494080
rect 496078 494068 496084 494080
rect 282880 494040 496084 494068
rect 282880 494028 282886 494040
rect 496078 494028 496084 494040
rect 496136 494028 496142 494080
rect 282822 492736 282828 492788
rect 282880 492776 282886 492788
rect 491938 492776 491944 492788
rect 282880 492748 491944 492776
rect 282880 492736 282886 492748
rect 491938 492736 491944 492748
rect 491996 492736 492002 492788
rect 282362 492668 282368 492720
rect 282420 492708 282426 492720
rect 493318 492708 493324 492720
rect 282420 492680 493324 492708
rect 282420 492668 282426 492680
rect 493318 492668 493324 492680
rect 493376 492668 493382 492720
rect 282822 491308 282828 491360
rect 282880 491348 282886 491360
rect 489178 491348 489184 491360
rect 282880 491320 489184 491348
rect 282880 491308 282886 491320
rect 489178 491308 489184 491320
rect 489236 491308 489242 491360
rect 282822 489948 282828 490000
rect 282880 489988 282886 490000
rect 483658 489988 483664 490000
rect 282880 489960 483664 489988
rect 282880 489948 282886 489960
rect 483658 489948 483664 489960
rect 483716 489948 483722 490000
rect 282270 489880 282276 489932
rect 282328 489920 282334 489932
rect 485038 489920 485044 489932
rect 282328 489892 485044 489920
rect 282328 489880 282334 489892
rect 485038 489880 485044 489892
rect 485096 489880 485102 489932
rect 282270 488520 282276 488572
rect 282328 488560 282334 488572
rect 482278 488560 482284 488572
rect 282328 488532 482284 488560
rect 282328 488520 282334 488532
rect 482278 488520 482284 488532
rect 482336 488520 482342 488572
rect 282822 487160 282828 487212
rect 282880 487200 282886 487212
rect 480898 487200 480904 487212
rect 282880 487172 480904 487200
rect 282880 487160 282886 487172
rect 480898 487160 480904 487172
rect 480956 487160 480962 487212
rect 282822 485868 282828 485920
rect 282880 485908 282886 485920
rect 465718 485908 465724 485920
rect 282880 485880 465724 485908
rect 282880 485868 282886 485880
rect 465718 485868 465724 485880
rect 465776 485868 465782 485920
rect 282270 485800 282276 485852
rect 282328 485840 282334 485852
rect 467098 485840 467104 485852
rect 282328 485812 467104 485840
rect 282328 485800 282334 485812
rect 467098 485800 467104 485812
rect 467156 485800 467162 485852
rect 281718 484372 281724 484424
rect 281776 484412 281782 484424
rect 449158 484412 449164 484424
rect 281776 484384 449164 484412
rect 281776 484372 281782 484384
rect 449158 484372 449164 484384
rect 449216 484372 449222 484424
rect 282270 483012 282276 483064
rect 282328 483052 282334 483064
rect 446398 483052 446404 483064
rect 282328 483024 446404 483052
rect 282328 483012 282334 483024
rect 446398 483012 446404 483024
rect 446456 483012 446462 483064
rect 282822 481720 282828 481772
rect 282880 481760 282886 481772
rect 442258 481760 442264 481772
rect 282880 481732 442264 481760
rect 282880 481720 282886 481732
rect 442258 481720 442264 481732
rect 442316 481720 442322 481772
rect 282546 481652 282552 481704
rect 282604 481692 282610 481704
rect 445018 481692 445024 481704
rect 282604 481664 445024 481692
rect 282604 481652 282610 481664
rect 445018 481652 445024 481664
rect 445076 481652 445082 481704
rect 282086 480224 282092 480276
rect 282144 480264 282150 480276
rect 435358 480264 435364 480276
rect 282144 480236 435364 480264
rect 282144 480224 282150 480236
rect 435358 480224 435364 480236
rect 435416 480224 435422 480276
rect 282822 478932 282828 478984
rect 282880 478972 282886 478984
rect 431218 478972 431224 478984
rect 282880 478944 431224 478972
rect 282880 478932 282886 478944
rect 431218 478932 431224 478944
rect 431276 478932 431282 478984
rect 282730 478864 282736 478916
rect 282788 478904 282794 478916
rect 433978 478904 433984 478916
rect 282788 478876 433984 478904
rect 282788 478864 282794 478876
rect 433978 478864 433984 478876
rect 434036 478864 434042 478916
rect 282822 477504 282828 477556
rect 282880 477544 282886 477556
rect 429838 477544 429844 477556
rect 282880 477516 429844 477544
rect 282880 477504 282886 477516
rect 429838 477504 429844 477516
rect 429896 477504 429902 477556
rect 282086 476076 282092 476128
rect 282144 476116 282150 476128
rect 428458 476116 428464 476128
rect 282144 476088 428464 476116
rect 282144 476076 282150 476088
rect 428458 476076 428464 476088
rect 428516 476076 428522 476128
rect 282822 474784 282828 474836
rect 282880 474824 282886 474836
rect 424318 474824 424324 474836
rect 282880 474796 424324 474824
rect 282880 474784 282886 474796
rect 424318 474784 424324 474796
rect 424376 474784 424382 474836
rect 282270 474716 282276 474768
rect 282328 474756 282334 474768
rect 427078 474756 427084 474768
rect 282328 474728 427084 474756
rect 282328 474716 282334 474728
rect 427078 474716 427084 474728
rect 427136 474716 427142 474768
rect 281718 473356 281724 473408
rect 281776 473396 281782 473408
rect 416038 473396 416044 473408
rect 281776 473368 416044 473396
rect 281776 473356 281782 473368
rect 416038 473356 416044 473368
rect 416096 473356 416102 473408
rect 282086 471996 282092 472048
rect 282144 472036 282150 472048
rect 477586 472036 477592 472048
rect 282144 472008 477592 472036
rect 282144 471996 282150 472008
rect 477586 471996 477592 472008
rect 477644 471996 477650 472048
rect 282822 470636 282828 470688
rect 282880 470676 282886 470688
rect 409138 470676 409144 470688
rect 282880 470648 409144 470676
rect 282880 470636 282886 470648
rect 409138 470636 409144 470648
rect 409196 470636 409202 470688
rect 282730 470568 282736 470620
rect 282788 470608 282794 470620
rect 411898 470608 411904 470620
rect 282788 470580 411904 470608
rect 282788 470568 282794 470580
rect 411898 470568 411904 470580
rect 411956 470568 411962 470620
rect 281902 469208 281908 469260
rect 281960 469248 281966 469260
rect 474826 469248 474832 469260
rect 281960 469220 474832 469248
rect 281960 469208 281966 469220
rect 474826 469208 474832 469220
rect 474884 469208 474890 469260
rect 282822 467848 282828 467900
rect 282880 467888 282886 467900
rect 473446 467888 473452 467900
rect 282880 467860 473452 467888
rect 282880 467848 282886 467860
rect 473446 467848 473452 467860
rect 473504 467848 473510 467900
rect 282730 466488 282736 466540
rect 282788 466528 282794 466540
rect 406378 466528 406384 466540
rect 282788 466500 406384 466528
rect 282788 466488 282794 466500
rect 406378 466488 406384 466500
rect 406436 466488 406442 466540
rect 282822 466420 282828 466472
rect 282880 466460 282886 466472
rect 470686 466460 470692 466472
rect 282880 466432 470692 466460
rect 282880 466420 282886 466432
rect 470686 466420 470692 466432
rect 470744 466420 470750 466472
rect 282822 465060 282828 465112
rect 282880 465100 282886 465112
rect 447778 465100 447784 465112
rect 282880 465072 447784 465100
rect 282880 465060 282886 465072
rect 447778 465060 447784 465072
rect 447836 465060 447842 465112
rect 282730 463768 282736 463820
rect 282788 463808 282794 463820
rect 417418 463808 417424 463820
rect 282788 463780 417424 463808
rect 282788 463768 282794 463780
rect 417418 463768 417424 463780
rect 417476 463768 417482 463820
rect 282822 463700 282828 463752
rect 282880 463740 282886 463752
rect 526346 463740 526352 463752
rect 282880 463712 526352 463740
rect 282880 463700 282886 463712
rect 526346 463700 526352 463712
rect 526404 463700 526410 463752
rect 282822 462340 282828 462392
rect 282880 462380 282886 462392
rect 283650 462380 283656 462392
rect 282880 462352 283656 462380
rect 282880 462340 282886 462352
rect 283650 462340 283656 462352
rect 283708 462340 283714 462392
rect 282822 460912 282828 460964
rect 282880 460952 282886 460964
rect 368566 460952 368572 460964
rect 282880 460924 368572 460952
rect 282880 460912 282886 460924
rect 368566 460912 368572 460924
rect 368624 460912 368630 460964
rect 282730 459620 282736 459672
rect 282788 459660 282794 459672
rect 283834 459660 283840 459672
rect 282788 459632 283840 459660
rect 282788 459620 282794 459632
rect 283834 459620 283840 459632
rect 283892 459620 283898 459672
rect 282822 459552 282828 459604
rect 282880 459592 282886 459604
rect 369946 459592 369952 459604
rect 282880 459564 369952 459592
rect 282880 459552 282886 459564
rect 369946 459552 369952 459564
rect 370004 459552 370010 459604
rect 281718 458192 281724 458244
rect 281776 458232 281782 458244
rect 284018 458232 284024 458244
rect 281776 458204 284024 458232
rect 281776 458192 281782 458204
rect 284018 458192 284024 458204
rect 284076 458192 284082 458244
rect 282086 456764 282092 456816
rect 282144 456804 282150 456816
rect 284110 456804 284116 456816
rect 282144 456776 284116 456804
rect 282144 456764 282150 456776
rect 284110 456764 284116 456776
rect 284168 456764 284174 456816
rect 281626 455472 281632 455524
rect 281684 455512 281690 455524
rect 284202 455512 284208 455524
rect 281684 455484 284208 455512
rect 281684 455472 281690 455484
rect 284202 455472 284208 455484
rect 284260 455472 284266 455524
rect 282822 455404 282828 455456
rect 282880 455444 282886 455456
rect 375558 455444 375564 455456
rect 282880 455416 375564 455444
rect 282880 455404 282886 455416
rect 375558 455404 375564 455416
rect 375616 455404 375622 455456
rect 282178 440376 282184 440428
rect 282236 440416 282242 440428
rect 384390 440416 384396 440428
rect 282236 440388 384396 440416
rect 282236 440376 282242 440388
rect 384390 440376 384396 440388
rect 384448 440376 384454 440428
rect 281442 440240 281448 440292
rect 281500 440280 281506 440292
rect 387150 440280 387156 440292
rect 281500 440252 387156 440280
rect 281500 440240 281506 440252
rect 387150 440240 387156 440252
rect 387208 440240 387214 440292
rect 282178 438880 282184 438932
rect 282236 438920 282242 438932
rect 381538 438920 381544 438932
rect 282236 438892 381544 438920
rect 282236 438880 282242 438892
rect 381538 438880 381544 438892
rect 381596 438880 381602 438932
rect 282178 436608 282184 436620
rect 282104 436580 282184 436608
rect 282104 436132 282132 436580
rect 282178 436568 282184 436580
rect 282236 436568 282242 436620
rect 282178 436160 282184 436212
rect 282236 436200 282242 436212
rect 377398 436200 377404 436212
rect 282236 436172 377404 436200
rect 282236 436160 282242 436172
rect 377398 436160 377404 436172
rect 377456 436160 377462 436212
rect 380158 436132 380164 436144
rect 282104 436104 380164 436132
rect 380158 436092 380164 436104
rect 380216 436092 380222 436144
rect 282178 434732 282184 434784
rect 282236 434772 282242 434784
rect 374730 434772 374736 434784
rect 282236 434744 374736 434772
rect 282236 434732 282242 434744
rect 374730 434732 374736 434744
rect 374788 434732 374794 434784
rect 282178 433304 282184 433356
rect 282236 433344 282242 433356
rect 373258 433344 373264 433356
rect 282236 433316 373264 433344
rect 282236 433304 282242 433316
rect 373258 433304 373264 433316
rect 373316 433304 373322 433356
rect 282089 431579 282147 431585
rect 282089 431545 282101 431579
rect 282135 431576 282147 431579
rect 282270 431576 282276 431588
rect 282135 431548 282276 431576
rect 282135 431545 282147 431548
rect 282089 431539 282147 431545
rect 282270 431536 282276 431548
rect 282328 431536 282334 431588
rect 282270 430652 282276 430704
rect 282328 430692 282334 430704
rect 388438 430692 388444 430704
rect 282328 430664 388444 430692
rect 282328 430652 282334 430664
rect 388438 430652 388444 430664
rect 388496 430652 388502 430704
rect 282270 430516 282276 430568
rect 282328 430556 282334 430568
rect 464338 430556 464344 430568
rect 282328 430528 464344 430556
rect 282328 430516 282334 430528
rect 464338 430516 464344 430528
rect 464396 430516 464402 430568
rect 281442 429156 281448 429208
rect 281500 429196 281506 429208
rect 416774 429196 416780 429208
rect 281500 429168 416780 429196
rect 281500 429156 281506 429168
rect 416774 429156 416780 429168
rect 416832 429156 416838 429208
rect 282270 429088 282276 429140
rect 282328 429128 282334 429140
rect 358170 429128 358176 429140
rect 282328 429100 358176 429128
rect 282328 429088 282334 429100
rect 358170 429088 358176 429100
rect 358228 429088 358234 429140
rect 282270 427728 282276 427780
rect 282328 427768 282334 427780
rect 358078 427768 358084 427780
rect 282328 427740 358084 427768
rect 282328 427728 282334 427740
rect 358078 427728 358084 427740
rect 358136 427728 358142 427780
rect 356790 427700 356796 427712
rect 283116 427672 356796 427700
rect 283116 427360 283144 427672
rect 356790 427660 356796 427672
rect 356848 427660 356854 427712
rect 282196 427332 283144 427360
rect 282196 427224 282224 427332
rect 282270 427224 282276 427236
rect 282196 427196 282276 427224
rect 282270 427184 282276 427196
rect 282328 427184 282334 427236
rect 282270 426368 282276 426420
rect 282328 426408 282334 426420
rect 356698 426408 356704 426420
rect 282328 426380 356704 426408
rect 282328 426368 282334 426380
rect 356698 426368 356704 426380
rect 356756 426368 356762 426420
rect 282270 425008 282276 425060
rect 282328 425048 282334 425060
rect 355410 425048 355416 425060
rect 282328 425020 355416 425048
rect 282328 425008 282334 425020
rect 355410 425008 355416 425020
rect 355468 425008 355474 425060
rect 282270 423580 282276 423632
rect 282328 423620 282334 423632
rect 355318 423620 355324 423632
rect 282328 423592 355324 423620
rect 282328 423580 282334 423592
rect 355318 423580 355324 423592
rect 355376 423580 355382 423632
rect 354030 423552 354036 423564
rect 282196 423524 354036 423552
rect 282196 423280 282224 423524
rect 354030 423512 354036 423524
rect 354088 423512 354094 423564
rect 282270 423280 282276 423292
rect 282196 423252 282276 423280
rect 282270 423240 282276 423252
rect 282328 423240 282334 423292
rect 282270 422220 282276 422272
rect 282328 422260 282334 422272
rect 353938 422260 353944 422272
rect 282328 422232 353944 422260
rect 282328 422220 282334 422232
rect 353938 422220 353944 422232
rect 353996 422220 354002 422272
rect 281626 421376 281632 421388
rect 281587 421348 281632 421376
rect 281626 421336 281632 421348
rect 281684 421336 281690 421388
rect 281626 421200 281632 421252
rect 281684 421240 281690 421252
rect 282454 421240 282460 421252
rect 281684 421212 282460 421240
rect 281684 421200 281690 421212
rect 282454 421200 282460 421212
rect 282512 421200 282518 421252
rect 282454 420996 282460 421048
rect 282512 421036 282518 421048
rect 282822 421036 282828 421048
rect 282512 421008 282828 421036
rect 282512 420996 282518 421008
rect 282822 420996 282828 421008
rect 282880 420996 282886 421048
rect 282822 420860 282828 420912
rect 282880 420900 282886 420912
rect 352650 420900 352656 420912
rect 282880 420872 352656 420900
rect 282880 420860 282886 420872
rect 352650 420860 352656 420872
rect 352708 420860 352714 420912
rect 282546 419432 282552 419484
rect 282604 419472 282610 419484
rect 476114 419472 476120 419484
rect 282604 419444 476120 419472
rect 282604 419432 282610 419444
rect 476114 419432 476120 419444
rect 476172 419432 476178 419484
rect 282822 419364 282828 419416
rect 282880 419404 282886 419416
rect 352558 419404 352564 419416
rect 282880 419376 352564 419404
rect 282880 419364 282886 419376
rect 352558 419364 352564 419376
rect 352616 419364 352622 419416
rect 282822 418072 282828 418124
rect 282880 418112 282886 418124
rect 474734 418112 474740 418124
rect 282880 418084 474740 418112
rect 282880 418072 282886 418084
rect 474734 418072 474740 418084
rect 474792 418072 474798 418124
rect 282270 417732 282276 417784
rect 282328 417772 282334 417784
rect 282546 417772 282552 417784
rect 282328 417744 282552 417772
rect 282328 417732 282334 417744
rect 282546 417732 282552 417744
rect 282604 417732 282610 417784
rect 282089 417639 282147 417645
rect 282089 417605 282101 417639
rect 282135 417636 282147 417639
rect 282270 417636 282276 417648
rect 282135 417608 282276 417636
rect 282135 417605 282147 417608
rect 282089 417599 282147 417605
rect 282270 417596 282276 417608
rect 282328 417596 282334 417648
rect 282822 416712 282828 416764
rect 282880 416752 282886 416764
rect 473354 416752 473360 416764
rect 282880 416724 473360 416752
rect 282880 416712 282886 416724
rect 473354 416712 473360 416724
rect 473412 416712 473418 416764
rect 284570 416372 284576 416424
rect 284628 416412 284634 416424
rect 453298 416412 453304 416424
rect 284628 416384 453304 416412
rect 284628 416372 284634 416384
rect 453298 416372 453304 416384
rect 453356 416372 453362 416424
rect 286226 416304 286232 416356
rect 286284 416344 286290 416356
rect 455414 416344 455420 416356
rect 286284 416316 455420 416344
rect 286284 416304 286290 416316
rect 455414 416304 455420 416316
rect 455472 416304 455478 416356
rect 286134 416236 286140 416288
rect 286192 416276 286198 416288
rect 456794 416276 456800 416288
rect 286192 416248 456800 416276
rect 286192 416236 286198 416248
rect 456794 416236 456800 416248
rect 456852 416236 456858 416288
rect 283282 416168 283288 416220
rect 283340 416208 283346 416220
rect 458174 416208 458180 416220
rect 283340 416180 458180 416208
rect 283340 416168 283346 416180
rect 458174 416168 458180 416180
rect 458232 416168 458238 416220
rect 283190 416100 283196 416152
rect 283248 416140 283254 416152
rect 459554 416140 459560 416152
rect 283248 416112 459560 416140
rect 283248 416100 283254 416112
rect 459554 416100 459560 416112
rect 459612 416100 459618 416152
rect 283098 416032 283104 416084
rect 283156 416072 283162 416084
rect 461026 416072 461032 416084
rect 283156 416044 461032 416072
rect 283156 416032 283162 416044
rect 461026 416032 461032 416044
rect 461084 416032 461090 416084
rect 282270 415420 282276 415472
rect 282328 415460 282334 415472
rect 282914 415460 282920 415472
rect 282328 415432 282920 415460
rect 282328 415420 282334 415432
rect 282914 415420 282920 415432
rect 282972 415420 282978 415472
rect 282822 415352 282828 415404
rect 282880 415392 282886 415404
rect 471974 415392 471980 415404
rect 282880 415364 471980 415392
rect 282880 415352 282886 415364
rect 471974 415352 471980 415364
rect 472032 415352 472038 415404
rect 282270 415284 282276 415336
rect 282328 415324 282334 415336
rect 470594 415324 470600 415336
rect 282328 415296 470600 415324
rect 282328 415284 282334 415296
rect 470594 415284 470600 415296
rect 470652 415284 470658 415336
rect 285398 415216 285404 415268
rect 285456 415256 285462 415268
rect 438578 415256 438584 415268
rect 285456 415228 438584 415256
rect 285456 415216 285462 415228
rect 438578 415216 438584 415228
rect 438636 415216 438642 415268
rect 285306 415148 285312 415200
rect 285364 415188 285370 415200
rect 438670 415188 438676 415200
rect 285364 415160 438676 415188
rect 285364 415148 285370 415160
rect 438670 415148 438676 415160
rect 438728 415148 438734 415200
rect 284754 415080 284760 415132
rect 284812 415120 284818 415132
rect 438118 415120 438124 415132
rect 284812 415092 438124 415120
rect 284812 415080 284818 415092
rect 438118 415080 438124 415092
rect 438176 415080 438182 415132
rect 284846 415012 284852 415064
rect 284904 415052 284910 415064
rect 438302 415052 438308 415064
rect 284904 415024 438308 415052
rect 284904 415012 284910 415024
rect 438302 415012 438308 415024
rect 438360 415012 438366 415064
rect 284662 414944 284668 414996
rect 284720 414984 284726 414996
rect 438210 414984 438216 414996
rect 284720 414956 438216 414984
rect 284720 414944 284726 414956
rect 438210 414944 438216 414956
rect 438268 414944 438274 414996
rect 285214 414876 285220 414928
rect 285272 414916 285278 414928
rect 445754 414916 445760 414928
rect 285272 414888 445760 414916
rect 285272 414876 285278 414888
rect 445754 414876 445760 414888
rect 445812 414876 445818 414928
rect 292022 414808 292028 414860
rect 292080 414848 292086 414860
rect 452746 414848 452752 414860
rect 292080 414820 452752 414848
rect 292080 414808 292086 414820
rect 452746 414808 452752 414820
rect 452804 414808 452810 414860
rect 283006 414740 283012 414792
rect 283064 414780 283070 414792
rect 467926 414780 467932 414792
rect 283064 414752 467932 414780
rect 283064 414740 283070 414752
rect 467926 414740 467932 414752
rect 467984 414740 467990 414792
rect 282914 414672 282920 414724
rect 282972 414712 282978 414724
rect 469214 414712 469220 414724
rect 282972 414684 469220 414712
rect 282972 414672 282978 414684
rect 469214 414672 469220 414684
rect 469272 414672 469278 414724
rect 285490 414604 285496 414656
rect 285548 414644 285554 414656
rect 438486 414644 438492 414656
rect 285548 414616 438492 414644
rect 285548 414604 285554 414616
rect 438486 414604 438492 414616
rect 438544 414604 438550 414656
rect 285582 414536 285588 414588
rect 285640 414576 285646 414588
rect 438394 414576 438400 414588
rect 285640 414548 438400 414576
rect 285640 414536 285646 414548
rect 438394 414536 438400 414548
rect 438452 414536 438458 414588
rect 337378 414468 337384 414520
rect 337436 414508 337442 414520
rect 454034 414508 454040 414520
rect 337436 414480 454040 414508
rect 337436 414468 337442 414480
rect 454034 414468 454040 414480
rect 454092 414468 454098 414520
rect 284386 414400 284392 414452
rect 284444 414440 284450 414452
rect 343726 414440 343732 414452
rect 284444 414412 343732 414440
rect 284444 414400 284450 414412
rect 343726 414400 343732 414412
rect 343784 414400 343790 414452
rect 284478 414332 284484 414384
rect 284536 414372 284542 414384
rect 342254 414372 342260 414384
rect 284536 414344 342260 414372
rect 284536 414332 284542 414344
rect 342254 414332 342260 414344
rect 342312 414332 342318 414384
rect 383102 413992 383108 414044
rect 383160 414032 383166 414044
rect 384577 414035 384635 414041
rect 384577 414032 384589 414035
rect 383160 414004 384589 414032
rect 383160 413992 383166 414004
rect 384577 414001 384589 414004
rect 384623 414001 384635 414035
rect 384577 413995 384635 414001
rect 282178 413924 282184 413976
rect 282236 413964 282242 413976
rect 402974 413964 402980 413976
rect 282236 413936 402980 413964
rect 282236 413924 282242 413936
rect 402974 413924 402980 413936
rect 403032 413924 403038 413976
rect 447778 413924 447784 413976
rect 447836 413964 447842 413976
rect 469398 413964 469404 413976
rect 447836 413936 469404 413964
rect 447836 413924 447842 413936
rect 469398 413924 469404 413936
rect 469456 413924 469462 413976
rect 496078 413924 496084 413976
rect 496136 413964 496142 413976
rect 505094 413964 505100 413976
rect 496136 413936 505100 413964
rect 496136 413924 496142 413936
rect 505094 413924 505100 413936
rect 505152 413924 505158 413976
rect 281629 413899 281687 413905
rect 281629 413865 281641 413899
rect 281675 413896 281687 413899
rect 282270 413896 282276 413908
rect 281675 413868 282276 413896
rect 281675 413865 281687 413868
rect 281629 413859 281687 413865
rect 282270 413856 282276 413868
rect 282328 413856 282334 413908
rect 283466 413856 283472 413908
rect 283524 413896 283530 413908
rect 396074 413896 396080 413908
rect 283524 413868 396080 413896
rect 283524 413856 283530 413868
rect 396074 413856 396080 413868
rect 396132 413856 396138 413908
rect 409138 413856 409144 413908
rect 409196 413896 409202 413908
rect 476114 413896 476120 413908
rect 409196 413868 476120 413896
rect 409196 413856 409202 413868
rect 476114 413856 476120 413868
rect 476172 413856 476178 413908
rect 489178 413856 489184 413908
rect 489236 413896 489242 413908
rect 502518 413896 502524 413908
rect 489236 413868 502524 413896
rect 489236 413856 489242 413868
rect 502518 413856 502524 413868
rect 502576 413856 502582 413908
rect 281718 413788 281724 413840
rect 281776 413828 281782 413840
rect 384485 413831 384543 413837
rect 384485 413828 384497 413831
rect 281776 413800 384497 413828
rect 281776 413788 281782 413800
rect 384485 413797 384497 413800
rect 384531 413797 384543 413831
rect 384485 413791 384543 413797
rect 384577 413831 384635 413837
rect 384577 413797 384589 413831
rect 384623 413828 384635 413831
rect 386509 413831 386567 413837
rect 386509 413828 386521 413831
rect 384623 413800 386521 413828
rect 384623 413797 384635 413800
rect 384577 413791 384635 413797
rect 386509 413797 386521 413800
rect 386555 413797 386567 413831
rect 386509 413791 386567 413797
rect 387150 413788 387156 413840
rect 387208 413828 387214 413840
rect 391934 413828 391940 413840
rect 387208 413800 391940 413828
rect 387208 413788 387214 413800
rect 391934 413788 391940 413800
rect 391992 413788 391998 413840
rect 411898 413788 411904 413840
rect 411956 413828 411962 413840
rect 477494 413828 477500 413840
rect 411956 413800 477500 413828
rect 411956 413788 411962 413800
rect 477494 413788 477500 413800
rect 477552 413788 477558 413840
rect 483658 413788 483664 413840
rect 483716 413828 483722 413840
rect 499574 413828 499580 413840
rect 483716 413800 499580 413828
rect 483716 413788 483722 413800
rect 499574 413788 499580 413800
rect 499632 413788 499638 413840
rect 281902 413720 281908 413772
rect 281960 413760 281966 413772
rect 389266 413760 389272 413772
rect 281960 413732 389272 413760
rect 281960 413720 281966 413732
rect 389266 413720 389272 413732
rect 389324 413720 389330 413772
rect 406378 413720 406384 413772
rect 406436 413760 406442 413772
rect 471974 413760 471980 413772
rect 406436 413732 471980 413760
rect 406436 413720 406442 413732
rect 471974 413720 471980 413732
rect 472032 413720 472038 413772
rect 491938 413720 491944 413772
rect 491996 413760 492002 413772
rect 503714 413760 503720 413772
rect 491996 413732 503720 413760
rect 491996 413720 492002 413732
rect 503714 413720 503720 413732
rect 503772 413720 503778 413772
rect 281994 413652 282000 413704
rect 282052 413692 282058 413704
rect 389174 413692 389180 413704
rect 282052 413664 389180 413692
rect 282052 413652 282058 413664
rect 389174 413652 389180 413664
rect 389232 413652 389238 413704
rect 416038 413652 416044 413704
rect 416096 413692 416102 413704
rect 478874 413692 478880 413704
rect 416096 413664 478880 413692
rect 416096 413652 416102 413664
rect 478874 413652 478880 413664
rect 478932 413652 478938 413704
rect 482278 413652 482284 413704
rect 482336 413692 482342 413704
rect 498286 413692 498292 413704
rect 482336 413664 498292 413692
rect 482336 413652 482342 413664
rect 498286 413652 498292 413664
rect 498344 413652 498350 413704
rect 498838 413652 498844 413704
rect 498896 413692 498902 413704
rect 506474 413692 506480 413704
rect 498896 413664 506480 413692
rect 498896 413652 498902 413664
rect 506474 413652 506480 413664
rect 506532 413652 506538 413704
rect 281810 413584 281816 413636
rect 281868 413624 281874 413636
rect 381357 413627 381415 413633
rect 381357 413624 381369 413627
rect 281868 413596 381369 413624
rect 281868 413584 281874 413596
rect 381357 413593 381369 413596
rect 381403 413593 381415 413627
rect 386414 413624 386420 413636
rect 381357 413587 381415 413593
rect 381464 413596 386420 413624
rect 282086 413516 282092 413568
rect 282144 413556 282150 413568
rect 381464 413556 381492 413596
rect 386414 413584 386420 413596
rect 386472 413584 386478 413636
rect 386509 413627 386567 413633
rect 386509 413593 386521 413627
rect 386555 413624 386567 413627
rect 387981 413627 388039 413633
rect 387981 413624 387993 413627
rect 386555 413596 387993 413624
rect 386555 413593 386567 413596
rect 386509 413587 386567 413593
rect 387981 413593 387993 413596
rect 388027 413593 388039 413627
rect 387981 413587 388039 413593
rect 388530 413584 388536 413636
rect 388588 413624 388594 413636
rect 404354 413624 404360 413636
rect 388588 413596 404360 413624
rect 388588 413584 388594 413596
rect 404354 413584 404360 413596
rect 404412 413584 404418 413636
rect 413922 413584 413928 413636
rect 413980 413624 413986 413636
rect 420178 413624 420184 413636
rect 413980 413596 420184 413624
rect 413980 413584 413986 413596
rect 420178 413584 420184 413596
rect 420236 413584 420242 413636
rect 424318 413584 424324 413636
rect 424376 413624 424382 413636
rect 480438 413624 480444 413636
rect 424376 413596 480444 413624
rect 424376 413584 424382 413596
rect 480438 413584 480444 413596
rect 480496 413584 480502 413636
rect 480898 413584 480904 413636
rect 480956 413624 480962 413636
rect 496814 413624 496820 413636
rect 480956 413596 496820 413624
rect 480956 413584 480962 413596
rect 496814 413584 496820 413596
rect 496872 413584 496878 413636
rect 282144 413528 381492 413556
rect 282144 413516 282150 413528
rect 381538 413516 381544 413568
rect 381596 413556 381602 413568
rect 394694 413556 394700 413568
rect 381596 413528 394700 413556
rect 381596 413516 381602 413528
rect 394694 413516 394700 413528
rect 394752 413516 394758 413568
rect 431218 413516 431224 413568
rect 431276 413556 431282 413568
rect 485774 413556 485780 413568
rect 431276 413528 485780 413556
rect 431276 413516 431282 413528
rect 485774 413516 485780 413528
rect 485832 413516 485838 413568
rect 282730 413448 282736 413500
rect 282788 413488 282794 413500
rect 375929 413491 375987 413497
rect 375929 413488 375941 413491
rect 282788 413460 375941 413488
rect 282788 413448 282794 413460
rect 375929 413457 375941 413460
rect 375975 413457 375987 413491
rect 375929 413451 375987 413457
rect 376018 413448 376024 413500
rect 376076 413488 376082 413500
rect 382274 413488 382280 413500
rect 376076 413460 382280 413488
rect 376076 413448 376082 413460
rect 382274 413448 382280 413460
rect 382332 413448 382338 413500
rect 383194 413448 383200 413500
rect 383252 413488 383258 413500
rect 401594 413488 401600 413500
rect 383252 413460 401600 413488
rect 383252 413448 383258 413460
rect 401594 413448 401600 413460
rect 401652 413448 401658 413500
rect 428458 413448 428464 413500
rect 428516 413488 428522 413500
rect 483014 413488 483020 413500
rect 428516 413460 483020 413488
rect 428516 413448 428522 413460
rect 483014 413448 483020 413460
rect 483072 413448 483078 413500
rect 493318 413448 493324 413500
rect 493376 413488 493382 413500
rect 503990 413488 503996 413500
rect 493376 413460 503996 413488
rect 493376 413448 493382 413460
rect 503990 413448 503996 413460
rect 504048 413448 504054 413500
rect 282638 413380 282644 413432
rect 282696 413420 282702 413432
rect 378597 413423 378655 413429
rect 378597 413420 378609 413423
rect 282696 413392 378609 413420
rect 282696 413380 282702 413392
rect 378597 413389 378609 413392
rect 378643 413389 378655 413423
rect 378597 413383 378655 413389
rect 378873 413423 378931 413429
rect 378873 413389 378885 413423
rect 378919 413420 378931 413423
rect 384393 413423 384451 413429
rect 384393 413420 384405 413423
rect 378919 413392 384405 413420
rect 378919 413389 378931 413392
rect 378873 413383 378931 413389
rect 384393 413389 384405 413392
rect 384439 413389 384451 413423
rect 384393 413383 384451 413389
rect 384577 413423 384635 413429
rect 384577 413389 384589 413423
rect 384623 413420 384635 413423
rect 397454 413420 397460 413432
rect 384623 413392 397460 413420
rect 384623 413389 384635 413392
rect 384577 413383 384635 413389
rect 397454 413380 397460 413392
rect 397512 413380 397518 413432
rect 427078 413380 427084 413432
rect 427136 413420 427142 413432
rect 481634 413420 481640 413432
rect 427136 413392 481640 413420
rect 427136 413380 427142 413392
rect 481634 413380 481640 413392
rect 481692 413380 481698 413432
rect 485038 413380 485044 413432
rect 485096 413420 485102 413432
rect 501046 413420 501052 413432
rect 485096 413392 501052 413420
rect 485096 413380 485102 413392
rect 501046 413380 501052 413392
rect 501104 413380 501110 413432
rect 282362 413312 282368 413364
rect 282420 413352 282426 413364
rect 382182 413352 382188 413364
rect 282420 413324 382188 413352
rect 282420 413312 282426 413324
rect 382182 413312 382188 413324
rect 382240 413312 382246 413364
rect 384301 413355 384359 413361
rect 384301 413321 384313 413355
rect 384347 413352 384359 413355
rect 397546 413352 397552 413364
rect 384347 413324 397552 413352
rect 384347 413321 384359 413324
rect 384301 413315 384359 413321
rect 397546 413312 397552 413324
rect 397604 413312 397610 413364
rect 429838 413312 429844 413364
rect 429896 413352 429902 413364
rect 484394 413352 484400 413364
rect 429896 413324 484400 413352
rect 429896 413312 429902 413324
rect 484394 413312 484400 413324
rect 484452 413312 484458 413364
rect 282454 413244 282460 413296
rect 282512 413284 282518 413296
rect 382366 413284 382372 413296
rect 282512 413256 382372 413284
rect 282512 413244 282518 413256
rect 382366 413244 382372 413256
rect 382424 413244 382430 413296
rect 383010 413244 383016 413296
rect 383068 413284 383074 413296
rect 398834 413284 398840 413296
rect 383068 413256 398840 413284
rect 383068 413244 383074 413256
rect 398834 413244 398840 413256
rect 398892 413244 398898 413296
rect 435358 413244 435364 413296
rect 435416 413284 435422 413296
rect 488534 413284 488540 413296
rect 435416 413256 488540 413284
rect 435416 413244 435422 413256
rect 488534 413244 488540 413256
rect 488592 413244 488598 413296
rect 282546 413176 282552 413228
rect 282604 413216 282610 413228
rect 377401 413219 377459 413225
rect 377401 413216 377413 413219
rect 282604 413188 377413 413216
rect 282604 413176 282610 413188
rect 377401 413185 377413 413188
rect 377447 413185 377459 413219
rect 377401 413179 377459 413185
rect 377493 413219 377551 413225
rect 377493 413185 377505 413219
rect 377539 413216 377551 413219
rect 378689 413219 378747 413225
rect 378689 413216 378701 413219
rect 377539 413188 378701 413216
rect 377539 413185 377551 413188
rect 377493 413179 377551 413185
rect 378689 413185 378701 413188
rect 378735 413185 378747 413219
rect 378689 413179 378747 413185
rect 378778 413176 378784 413228
rect 378836 413216 378842 413228
rect 384298 413216 384304 413228
rect 378836 413188 384304 413216
rect 378836 413176 378842 413188
rect 384298 413176 384304 413188
rect 384356 413176 384362 413228
rect 384390 413176 384396 413228
rect 384448 413216 384454 413228
rect 393314 413216 393320 413228
rect 384448 413188 393320 413216
rect 384448 413176 384454 413188
rect 393314 413176 393320 413188
rect 393372 413176 393378 413228
rect 433978 413176 433984 413228
rect 434036 413216 434042 413228
rect 487154 413216 487160 413228
rect 434036 413188 487160 413216
rect 434036 413176 434042 413188
rect 487154 413176 487160 413188
rect 487212 413176 487218 413228
rect 282730 413108 282736 413160
rect 282788 413148 282794 413160
rect 378597 413151 378655 413157
rect 282788 413120 378272 413148
rect 282788 413108 282794 413120
rect 281626 413040 281632 413092
rect 281684 413080 281690 413092
rect 378134 413080 378140 413092
rect 281684 413052 378140 413080
rect 281684 413040 281690 413052
rect 378134 413040 378140 413052
rect 378192 413040 378198 413092
rect 378244 413080 378272 413120
rect 378597 413117 378609 413151
rect 378643 413148 378655 413151
rect 383654 413148 383660 413160
rect 378643 413120 383660 413148
rect 378643 413117 378655 413120
rect 378597 413111 378655 413117
rect 383654 413108 383660 413120
rect 383712 413108 383718 413160
rect 384485 413151 384543 413157
rect 384485 413117 384497 413151
rect 384531 413148 384543 413151
rect 390554 413148 390560 413160
rect 384531 413120 390560 413148
rect 384531 413117 384543 413120
rect 384485 413111 384543 413117
rect 390554 413108 390560 413120
rect 390612 413108 390618 413160
rect 417418 413108 417424 413160
rect 417476 413148 417482 413160
rect 468110 413148 468116 413160
rect 417476 413120 468116 413148
rect 417476 413108 417482 413120
rect 468110 413108 468116 413120
rect 468168 413108 468174 413160
rect 379606 413080 379612 413092
rect 378244 413052 379612 413080
rect 379606 413040 379612 413052
rect 379664 413040 379670 413092
rect 380158 413040 380164 413092
rect 380216 413080 380222 413092
rect 384577 413083 384635 413089
rect 384577 413080 384589 413083
rect 380216 413052 384589 413080
rect 380216 413040 380222 413052
rect 384577 413049 384589 413052
rect 384623 413049 384635 413083
rect 384577 413043 384635 413049
rect 385770 413040 385776 413092
rect 385828 413080 385834 413092
rect 396074 413080 396080 413092
rect 385828 413052 396080 413080
rect 385828 413040 385834 413052
rect 396074 413040 396080 413052
rect 396132 413040 396138 413092
rect 442258 413040 442264 413092
rect 442316 413080 442322 413092
rect 489914 413080 489920 413092
rect 442316 413052 489920 413080
rect 442316 413040 442322 413052
rect 489914 413040 489920 413052
rect 489972 413040 489978 413092
rect 282270 412972 282276 413024
rect 282328 413012 282334 413024
rect 287054 413012 287060 413024
rect 282328 412984 287060 413012
rect 282328 412972 282334 412984
rect 287054 412972 287060 412984
rect 287112 412972 287118 413024
rect 296622 412972 296628 413024
rect 296680 413012 296686 413024
rect 306374 413012 306380 413024
rect 296680 412984 306380 413012
rect 296680 412972 296686 412984
rect 306374 412972 306380 412984
rect 306432 412972 306438 413024
rect 315942 412972 315948 413024
rect 316000 413012 316006 413024
rect 331122 413012 331128 413024
rect 316000 412984 331128 413012
rect 316000 412972 316006 412984
rect 331122 412972 331128 412984
rect 331180 412972 331186 413024
rect 335262 412972 335268 413024
rect 335320 413012 335326 413024
rect 350442 413012 350448 413024
rect 335320 412984 350448 413012
rect 335320 412972 335326 412984
rect 350442 412972 350448 412984
rect 350500 412972 350506 413024
rect 354582 412972 354588 413024
rect 354640 413012 354646 413024
rect 364334 413012 364340 413024
rect 354640 412984 364340 413012
rect 354640 412972 354646 412984
rect 364334 412972 364340 412984
rect 364392 412972 364398 413024
rect 373905 413015 373963 413021
rect 373905 412981 373917 413015
rect 373951 413012 373963 413015
rect 376754 413012 376760 413024
rect 373951 412984 376760 413012
rect 373951 412981 373963 412984
rect 373905 412975 373963 412981
rect 376754 412972 376760 412984
rect 376812 412972 376818 413024
rect 377401 413015 377459 413021
rect 377401 412981 377413 413015
rect 377447 413012 377459 413015
rect 380894 413012 380900 413024
rect 377447 412984 380900 413012
rect 377447 412981 377459 412984
rect 377401 412975 377459 412981
rect 380894 412972 380900 412984
rect 380952 412972 380958 413024
rect 381357 413015 381415 413021
rect 381357 412981 381369 413015
rect 381403 413012 381415 413015
rect 387794 413012 387800 413024
rect 381403 412984 387800 413012
rect 381403 412981 381415 412984
rect 381357 412975 381415 412981
rect 387794 412972 387800 412984
rect 387852 412972 387858 413024
rect 387889 413015 387947 413021
rect 387889 412981 387901 413015
rect 387935 413012 387947 413015
rect 397454 413012 397460 413024
rect 387935 412984 397460 413012
rect 387935 412981 387947 412984
rect 387889 412975 387947 412981
rect 397454 412972 397460 412984
rect 397512 412972 397518 413024
rect 445018 412972 445024 413024
rect 445076 413012 445082 413024
rect 491294 413012 491300 413024
rect 445076 412984 491300 413012
rect 445076 412972 445082 412984
rect 491294 412972 491300 412984
rect 491352 412972 491358 413024
rect 284110 412904 284116 412956
rect 284168 412944 284174 412956
rect 373994 412944 374000 412956
rect 284168 412916 374000 412944
rect 284168 412904 284174 412916
rect 373994 412904 374000 412916
rect 374052 412904 374058 412956
rect 375929 412947 375987 412953
rect 375929 412913 375941 412947
rect 375975 412944 375987 412947
rect 375975 412916 382688 412944
rect 375975 412913 375987 412916
rect 375929 412907 375987 412913
rect 284202 412836 284208 412888
rect 284260 412876 284266 412888
rect 374178 412876 374184 412888
rect 284260 412848 374184 412876
rect 284260 412836 284266 412848
rect 374178 412836 374184 412848
rect 374236 412836 374242 412888
rect 374638 412836 374644 412888
rect 374696 412876 374702 412888
rect 382274 412876 382280 412888
rect 374696 412848 382280 412876
rect 374696 412836 374702 412848
rect 382274 412836 382280 412848
rect 382332 412836 382338 412888
rect 382660 412876 382688 412916
rect 382918 412904 382924 412956
rect 382976 412944 382982 412956
rect 384209 412947 384267 412953
rect 384209 412944 384221 412947
rect 382976 412916 384221 412944
rect 382976 412904 382982 412916
rect 384209 412913 384221 412916
rect 384255 412913 384267 412947
rect 384209 412907 384267 412913
rect 384298 412904 384304 412956
rect 384356 412944 384362 412956
rect 403158 412944 403164 412956
rect 384356 412916 403164 412944
rect 384356 412904 384362 412916
rect 403158 412904 403164 412916
rect 403216 412904 403222 412956
rect 446398 412904 446404 412956
rect 446456 412944 446462 412956
rect 491386 412944 491392 412956
rect 446456 412916 491392 412944
rect 446456 412904 446462 412916
rect 491386 412904 491392 412916
rect 491444 412904 491450 412956
rect 385034 412876 385040 412888
rect 382660 412848 385040 412876
rect 385034 412836 385040 412848
rect 385092 412836 385098 412888
rect 385678 412836 385684 412888
rect 385736 412876 385742 412888
rect 394694 412876 394700 412888
rect 385736 412848 394700 412876
rect 385736 412836 385742 412848
rect 394694 412836 394700 412848
rect 394752 412836 394758 412888
rect 449158 412836 449164 412888
rect 449216 412876 449222 412888
rect 492674 412876 492680 412888
rect 449216 412848 492680 412876
rect 449216 412836 449222 412848
rect 492674 412836 492680 412848
rect 492732 412836 492738 412888
rect 284018 412768 284024 412820
rect 284076 412808 284082 412820
rect 372614 412808 372620 412820
rect 284076 412780 372620 412808
rect 284076 412768 284082 412780
rect 372614 412768 372620 412780
rect 372672 412768 372678 412820
rect 373258 412768 373264 412820
rect 373316 412808 373322 412820
rect 400214 412808 400220 412820
rect 373316 412780 400220 412808
rect 373316 412768 373322 412780
rect 400214 412768 400220 412780
rect 400272 412768 400278 412820
rect 410518 412768 410524 412820
rect 410576 412808 410582 412820
rect 517514 412808 517520 412820
rect 410576 412780 517520 412808
rect 410576 412768 410582 412780
rect 517514 412768 517520 412780
rect 517572 412768 517578 412820
rect 283834 412700 283840 412752
rect 283892 412740 283898 412752
rect 371234 412740 371240 412752
rect 283892 412712 371240 412740
rect 283892 412700 283898 412712
rect 371234 412700 371240 412712
rect 371292 412700 371298 412752
rect 371326 412700 371332 412752
rect 371384 412740 371390 412752
rect 373905 412743 373963 412749
rect 373905 412740 373917 412743
rect 371384 412712 373917 412740
rect 371384 412700 371390 412712
rect 373905 412709 373917 412712
rect 373951 412709 373963 412743
rect 373905 412703 373963 412709
rect 374730 412700 374736 412752
rect 374788 412740 374794 412752
rect 377309 412743 377367 412749
rect 377309 412740 377321 412743
rect 374788 412712 377321 412740
rect 374788 412700 374794 412712
rect 377309 412709 377321 412712
rect 377355 412709 377367 412743
rect 377309 412703 377367 412709
rect 377398 412700 377404 412752
rect 377456 412740 377462 412752
rect 384301 412743 384359 412749
rect 384301 412740 384313 412743
rect 377456 412712 384313 412740
rect 377456 412700 377462 412712
rect 384301 412709 384313 412712
rect 384347 412709 384359 412743
rect 384301 412703 384359 412709
rect 384393 412743 384451 412749
rect 384393 412709 384405 412743
rect 384439 412740 384451 412743
rect 398834 412740 398840 412752
rect 384439 412712 398840 412740
rect 384439 412709 384451 412712
rect 384393 412703 384451 412709
rect 398834 412700 398840 412712
rect 398892 412700 398898 412752
rect 467098 412700 467104 412752
rect 467156 412740 467162 412752
rect 495710 412740 495716 412752
rect 467156 412712 495716 412740
rect 467156 412700 467162 412712
rect 495710 412700 495716 412712
rect 495768 412700 495774 412752
rect 283650 412632 283656 412684
rect 283708 412672 283714 412684
rect 367094 412672 367100 412684
rect 283708 412644 367100 412672
rect 283708 412632 283714 412644
rect 367094 412632 367100 412644
rect 367152 412632 367158 412684
rect 367738 412632 367744 412684
rect 367796 412672 367802 412684
rect 385034 412672 385040 412684
rect 367796 412644 385040 412672
rect 367796 412632 367802 412644
rect 385034 412632 385040 412644
rect 385092 412632 385098 412684
rect 387889 412675 387947 412681
rect 387889 412672 387901 412675
rect 385144 412644 387901 412672
rect 283926 412564 283932 412616
rect 283984 412604 283990 412616
rect 352098 412604 352104 412616
rect 283984 412576 352104 412604
rect 283984 412564 283990 412576
rect 352098 412564 352104 412576
rect 352156 412564 352162 412616
rect 384209 412607 384267 412613
rect 384209 412573 384221 412607
rect 384255 412604 384267 412607
rect 385144 412604 385172 412644
rect 387889 412641 387901 412644
rect 387935 412641 387947 412675
rect 387889 412635 387947 412641
rect 387981 412675 388039 412681
rect 387981 412641 387993 412675
rect 388027 412672 388039 412675
rect 400214 412672 400220 412684
rect 388027 412644 400220 412672
rect 388027 412641 388039 412644
rect 387981 412635 388039 412641
rect 400214 412632 400220 412644
rect 400272 412632 400278 412684
rect 465718 412632 465724 412684
rect 465776 412672 465782 412684
rect 494054 412672 494060 412684
rect 465776 412644 494060 412672
rect 465776 412632 465782 412644
rect 494054 412632 494060 412644
rect 494112 412632 494118 412684
rect 384255 412576 385172 412604
rect 384255 412573 384267 412576
rect 384209 412567 384267 412573
rect 283742 412496 283748 412548
rect 283800 412536 283806 412548
rect 352006 412536 352012 412548
rect 283800 412508 352012 412536
rect 283800 412496 283806 412508
rect 352006 412496 352012 412508
rect 352064 412496 352070 412548
rect 283834 412428 283840 412480
rect 283892 412468 283898 412480
rect 353294 412468 353300 412480
rect 283892 412440 353300 412468
rect 283892 412428 283898 412440
rect 353294 412428 353300 412440
rect 353352 412428 353358 412480
rect 284018 412360 284024 412412
rect 284076 412400 284082 412412
rect 354674 412400 354680 412412
rect 284076 412372 354680 412400
rect 284076 412360 284082 412372
rect 354674 412360 354680 412372
rect 354732 412360 354738 412412
rect 284110 412292 284116 412344
rect 284168 412332 284174 412344
rect 356146 412332 356152 412344
rect 284168 412304 356152 412332
rect 284168 412292 284174 412304
rect 356146 412292 356152 412304
rect 356204 412292 356210 412344
rect 283466 412224 283472 412276
rect 283524 412264 283530 412276
rect 357526 412264 357532 412276
rect 283524 412236 357532 412264
rect 283524 412224 283530 412236
rect 357526 412224 357532 412236
rect 357584 412224 357590 412276
rect 284202 412156 284208 412208
rect 284260 412196 284266 412208
rect 358906 412196 358912 412208
rect 284260 412168 358912 412196
rect 284260 412156 284266 412168
rect 358906 412156 358912 412168
rect 358964 412156 358970 412208
rect 343082 412088 343088 412140
rect 343140 412128 343146 412140
rect 467834 412128 467840 412140
rect 343140 412100 467840 412128
rect 343140 412088 343146 412100
rect 467834 412088 467840 412100
rect 467892 412088 467898 412140
rect 338022 412020 338028 412072
rect 338080 412060 338086 412072
rect 463694 412060 463700 412072
rect 338080 412032 463700 412060
rect 338080 412020 338086 412032
rect 463694 412020 463700 412032
rect 463752 412020 463758 412072
rect 283374 411952 283380 412004
rect 283432 411992 283438 412004
rect 452654 411992 452660 412004
rect 283432 411964 452660 411992
rect 283432 411952 283438 411964
rect 452654 411952 452660 411964
rect 452712 411952 452718 412004
rect 292574 411884 292580 411936
rect 292632 411924 292638 411936
rect 465074 411924 465080 411936
rect 292632 411896 465080 411924
rect 292632 411884 292638 411896
rect 465074 411884 465080 411896
rect 465132 411884 465138 411936
rect 283650 411816 283656 411868
rect 283708 411856 283714 411868
rect 350626 411856 350632 411868
rect 283708 411828 350632 411856
rect 283708 411816 283714 411828
rect 350626 411816 350632 411828
rect 350684 411816 350690 411868
rect 283558 411748 283564 411800
rect 283616 411788 283622 411800
rect 349154 411788 349160 411800
rect 283616 411760 349160 411788
rect 283616 411748 283622 411760
rect 349154 411748 349160 411760
rect 349212 411748 349218 411800
rect 286962 411680 286968 411732
rect 287020 411720 287026 411732
rect 347774 411720 347780 411732
rect 287020 411692 347780 411720
rect 287020 411680 287026 411692
rect 347774 411680 347780 411692
rect 347832 411680 347838 411732
rect 286870 411612 286876 411664
rect 286928 411652 286934 411664
rect 346394 411652 346400 411664
rect 286928 411624 346400 411652
rect 286928 411612 286934 411624
rect 346394 411612 346400 411624
rect 346452 411612 346458 411664
rect 286686 411544 286692 411596
rect 286744 411584 286750 411596
rect 345014 411584 345020 411596
rect 286744 411556 345020 411584
rect 286744 411544 286750 411556
rect 345014 411544 345020 411556
rect 345072 411544 345078 411596
rect 286778 411476 286784 411528
rect 286836 411516 286842 411528
rect 343634 411516 343640 411528
rect 286836 411488 343640 411516
rect 286836 411476 286842 411488
rect 343634 411476 343640 411488
rect 343692 411476 343698 411528
rect 338758 411272 338764 411324
rect 338816 411312 338822 411324
rect 405734 411312 405740 411324
rect 338816 411284 405740 411312
rect 338816 411272 338822 411284
rect 405734 411272 405740 411284
rect 405792 411272 405798 411324
rect 282730 411204 282736 411256
rect 282788 411244 282794 411256
rect 466454 411244 466460 411256
rect 282788 411216 466460 411244
rect 282788 411204 282794 411216
rect 466454 411204 466460 411216
rect 466512 411204 466518 411256
rect 282822 411136 282828 411188
rect 282880 411176 282886 411188
rect 343082 411176 343088 411188
rect 282880 411148 343088 411176
rect 282880 411136 282886 411148
rect 343082 411136 343088 411148
rect 343140 411136 343146 411188
rect 281626 411068 281632 411120
rect 281684 411108 281690 411120
rect 438762 411108 438768 411120
rect 281684 411080 438768 411108
rect 281684 411068 281690 411080
rect 438762 411068 438768 411080
rect 438820 411068 438826 411120
rect 281994 411000 282000 411052
rect 282052 411040 282058 411052
rect 451274 411040 451280 411052
rect 282052 411012 451280 411040
rect 282052 411000 282058 411012
rect 451274 411000 451280 411012
rect 451332 411000 451338 411052
rect 282178 410932 282184 410984
rect 282236 410972 282242 410984
rect 456058 410972 456064 410984
rect 282236 410944 456064 410972
rect 282236 410932 282242 410944
rect 456058 410932 456064 410944
rect 456116 410932 456122 410984
rect 282270 410864 282276 410916
rect 282328 410904 282334 410916
rect 457438 410904 457444 410916
rect 282328 410876 457444 410904
rect 282328 410864 282334 410876
rect 457438 410864 457444 410876
rect 457496 410864 457502 410916
rect 282638 410796 282644 410848
rect 282696 410836 282702 410848
rect 458818 410836 458824 410848
rect 282696 410808 458824 410836
rect 282696 410796 282702 410808
rect 458818 410796 458824 410808
rect 458876 410796 458882 410848
rect 282546 410728 282552 410780
rect 282604 410768 282610 410780
rect 460198 410768 460204 410780
rect 282604 410740 460204 410768
rect 282604 410728 282610 410740
rect 460198 410728 460204 410740
rect 460256 410728 460262 410780
rect 282454 410660 282460 410712
rect 282512 410700 282518 410712
rect 460382 410700 460388 410712
rect 282512 410672 460388 410700
rect 282512 410660 282518 410672
rect 460382 410660 460388 410672
rect 460440 410660 460446 410712
rect 282362 410592 282368 410644
rect 282420 410632 282426 410644
rect 460934 410632 460940 410644
rect 282420 410604 460940 410632
rect 282420 410592 282426 410604
rect 460934 410592 460940 410604
rect 460992 410592 460998 410644
rect 282822 410524 282828 410576
rect 282880 410564 282886 410576
rect 462314 410564 462320 410576
rect 282880 410536 462320 410564
rect 282880 410524 282886 410536
rect 462314 410524 462320 410536
rect 462372 410524 462378 410576
rect 284294 410456 284300 410508
rect 284352 410496 284358 410508
rect 340874 410496 340880 410508
rect 284352 410468 340880 410496
rect 284352 410456 284358 410468
rect 340874 410456 340880 410468
rect 340932 410456 340938 410508
rect 281718 409776 281724 409828
rect 281776 409816 281782 409828
rect 292574 409816 292580 409828
rect 281776 409788 292580 409816
rect 281776 409776 281782 409788
rect 292574 409776 292580 409788
rect 292632 409776 292638 409828
rect 281718 408416 281724 408468
rect 281776 408456 281782 408468
rect 338022 408456 338028 408468
rect 281776 408428 338028 408456
rect 281776 408416 281782 408428
rect 338022 408416 338028 408428
rect 338080 408416 338086 408468
rect 281626 403996 281632 404048
rect 281684 404036 281690 404048
rect 283282 404036 283288 404048
rect 281684 404008 283288 404036
rect 281684 403996 281690 404008
rect 283282 403996 283288 404008
rect 283340 403996 283346 404048
rect 282822 402228 282828 402280
rect 282880 402268 282886 402280
rect 286134 402268 286140 402280
rect 282880 402240 286140 402268
rect 282880 402228 282886 402240
rect 286134 402228 286140 402240
rect 286192 402228 286198 402280
rect 282822 401140 282828 401192
rect 282880 401180 282886 401192
rect 286226 401180 286232 401192
rect 282880 401152 286232 401180
rect 282880 401140 282886 401152
rect 286226 401140 286232 401152
rect 286284 401140 286290 401192
rect 282822 400120 282828 400172
rect 282880 400160 282886 400172
rect 337378 400160 337384 400172
rect 282880 400132 337384 400160
rect 282880 400120 282886 400132
rect 337378 400120 337384 400132
rect 337436 400120 337442 400172
rect 282270 400052 282276 400104
rect 282328 400092 282334 400104
rect 292022 400092 292028 400104
rect 282328 400064 292028 400092
rect 282328 400052 282334 400064
rect 292022 400052 292028 400064
rect 292080 400052 292086 400104
rect 281626 398148 281632 398200
rect 281684 398188 281690 398200
rect 283374 398188 283380 398200
rect 281684 398160 283380 398188
rect 281684 398148 281690 398160
rect 283374 398148 283380 398160
rect 283432 398148 283438 398200
rect 281626 397196 281632 397248
rect 281684 397236 281690 397248
rect 284202 397236 284208 397248
rect 281684 397208 284208 397236
rect 281684 397196 281690 397208
rect 284202 397196 284208 397208
rect 284260 397196 284266 397248
rect 281626 396448 281632 396500
rect 281684 396488 281690 396500
rect 283466 396488 283472 396500
rect 281684 396460 283472 396488
rect 281684 396448 281690 396460
rect 283466 396448 283472 396460
rect 283524 396448 283530 396500
rect 282178 396012 282184 396024
rect 282139 395984 282184 396012
rect 282178 395972 282184 395984
rect 282236 395972 282242 396024
rect 281626 395768 281632 395820
rect 281684 395808 281690 395820
rect 284110 395808 284116 395820
rect 281684 395780 284116 395808
rect 281684 395768 281690 395780
rect 284110 395768 284116 395780
rect 284168 395768 284174 395820
rect 281626 394340 281632 394392
rect 281684 394380 281690 394392
rect 284018 394380 284024 394392
rect 281684 394352 284024 394380
rect 281684 394340 281690 394352
rect 284018 394340 284024 394352
rect 284076 394340 284082 394392
rect 281626 393184 281632 393236
rect 281684 393224 281690 393236
rect 283834 393224 283840 393236
rect 281684 393196 283840 393224
rect 281684 393184 281690 393196
rect 283834 393184 283840 393196
rect 283892 393184 283898 393236
rect 281626 392028 281632 392080
rect 281684 392068 281690 392080
rect 283926 392068 283932 392080
rect 281684 392040 283932 392068
rect 281684 392028 281690 392040
rect 283926 392028 283932 392040
rect 283984 392028 283990 392080
rect 281626 391620 281632 391672
rect 281684 391660 281690 391672
rect 283742 391660 283748 391672
rect 281684 391632 283748 391660
rect 281684 391620 281690 391632
rect 283742 391620 283748 391632
rect 283800 391620 283806 391672
rect 281626 390124 281632 390176
rect 281684 390164 281690 390176
rect 283650 390164 283656 390176
rect 281684 390136 283656 390164
rect 281684 390124 281690 390136
rect 283650 390124 283656 390136
rect 283708 390124 283714 390176
rect 281626 389036 281632 389088
rect 281684 389076 281690 389088
rect 283558 389076 283564 389088
rect 281684 389048 283564 389076
rect 281684 389036 281690 389048
rect 283558 389036 283564 389048
rect 283616 389036 283622 389088
rect 281626 388288 281632 388340
rect 281684 388328 281690 388340
rect 286962 388328 286968 388340
rect 281684 388300 286968 388328
rect 281684 388288 281690 388300
rect 286962 388288 286968 388300
rect 287020 388288 287026 388340
rect 281626 387064 281632 387116
rect 281684 387104 281690 387116
rect 286870 387104 286876 387116
rect 281684 387076 286876 387104
rect 281684 387064 281690 387076
rect 286870 387064 286876 387076
rect 286928 387064 286934 387116
rect 282181 386427 282239 386433
rect 282181 386393 282193 386427
rect 282227 386424 282239 386427
rect 282270 386424 282276 386436
rect 282227 386396 282276 386424
rect 282227 386393 282239 386396
rect 282181 386387 282239 386393
rect 282270 386384 282276 386396
rect 282328 386384 282334 386436
rect 281626 386044 281632 386096
rect 281684 386084 281690 386096
rect 286686 386084 286692 386096
rect 281684 386056 286692 386084
rect 281684 386044 281690 386056
rect 286686 386044 286692 386056
rect 286744 386044 286750 386096
rect 281626 385228 281632 385280
rect 281684 385268 281690 385280
rect 286778 385268 286784 385280
rect 281684 385240 286784 385268
rect 281684 385228 281690 385240
rect 286778 385228 286784 385240
rect 286836 385228 286842 385280
rect 281626 384004 281632 384056
rect 281684 384044 281690 384056
rect 284386 384044 284392 384056
rect 281684 384016 284392 384044
rect 281684 384004 281690 384016
rect 284386 384004 284392 384016
rect 284444 384004 284450 384056
rect 281626 383256 281632 383308
rect 281684 383296 281690 383308
rect 284478 383296 284484 383308
rect 281684 383268 284484 383296
rect 281684 383256 281690 383268
rect 284478 383256 284484 383268
rect 284536 383256 284542 383308
rect 281810 382168 281816 382220
rect 281868 382208 281874 382220
rect 339494 382208 339500 382220
rect 281868 382180 339500 382208
rect 281868 382168 281874 382180
rect 339494 382168 339500 382180
rect 339552 382168 339558 382220
rect 281626 382100 281632 382152
rect 281684 382140 281690 382152
rect 284294 382140 284300 382152
rect 281684 382112 284300 382140
rect 281684 382100 281690 382112
rect 284294 382100 284300 382112
rect 284352 382100 284358 382152
rect 281626 380808 281632 380860
rect 281684 380848 281690 380860
rect 338114 380848 338120 380860
rect 281684 380820 338120 380848
rect 281684 380808 281690 380820
rect 338114 380808 338120 380820
rect 338172 380808 338178 380860
rect 281626 379448 281632 379500
rect 281684 379488 281690 379500
rect 336826 379488 336832 379500
rect 281684 379460 336832 379488
rect 281684 379448 281690 379460
rect 336826 379448 336832 379460
rect 336884 379448 336890 379500
rect 281626 378088 281632 378140
rect 281684 378128 281690 378140
rect 336734 378128 336740 378140
rect 281684 378100 336740 378128
rect 281684 378088 281690 378100
rect 336734 378088 336740 378100
rect 336792 378088 336798 378140
rect 281810 378020 281816 378072
rect 281868 378060 281874 378072
rect 335354 378060 335360 378072
rect 281868 378032 335360 378060
rect 281868 378020 281874 378032
rect 335354 378020 335360 378032
rect 335412 378020 335418 378072
rect 281626 376660 281632 376712
rect 281684 376700 281690 376712
rect 333974 376700 333980 376712
rect 281684 376672 333980 376700
rect 281684 376660 281690 376672
rect 333974 376660 333980 376672
rect 334032 376660 334038 376712
rect 281626 375300 281632 375352
rect 281684 375340 281690 375352
rect 332594 375340 332600 375352
rect 281684 375312 332600 375340
rect 281684 375300 281690 375312
rect 332594 375300 332600 375312
rect 332652 375300 332658 375352
rect 281810 373940 281816 373992
rect 281868 373980 281874 373992
rect 329926 373980 329932 373992
rect 281868 373952 329932 373980
rect 281868 373940 281874 373952
rect 329926 373940 329932 373952
rect 329984 373940 329990 373992
rect 281626 373124 281632 373176
rect 281684 373164 281690 373176
rect 287790 373164 287796 373176
rect 281684 373136 287796 373164
rect 281684 373124 281690 373136
rect 287790 373124 287796 373136
rect 287848 373124 287854 373176
rect 281626 371900 281632 371952
rect 281684 371940 281690 371952
rect 286594 371940 286600 371952
rect 281684 371912 286600 371940
rect 281684 371900 281690 371912
rect 286594 371900 286600 371912
rect 286652 371900 286658 371952
rect 281810 371152 281816 371204
rect 281868 371192 281874 371204
rect 327074 371192 327080 371204
rect 281868 371164 327080 371192
rect 281868 371152 281874 371164
rect 327074 371152 327080 371164
rect 327132 371152 327138 371204
rect 281626 370948 281632 371000
rect 281684 370988 281690 371000
rect 285122 370988 285128 371000
rect 281684 370960 285128 370988
rect 281684 370948 281690 370960
rect 285122 370948 285128 370960
rect 285180 370948 285186 371000
rect 282270 369900 282276 369912
rect 282231 369872 282276 369900
rect 282270 369860 282276 369872
rect 282328 369860 282334 369912
rect 281626 369792 281632 369844
rect 281684 369832 281690 369844
rect 325694 369832 325700 369844
rect 281684 369804 325700 369832
rect 281684 369792 281690 369804
rect 325694 369792 325700 369804
rect 325752 369792 325758 369844
rect 281626 368432 281632 368484
rect 281684 368472 281690 368484
rect 315298 368472 315304 368484
rect 281684 368444 315304 368472
rect 281684 368432 281690 368444
rect 315298 368432 315304 368444
rect 315356 368432 315362 368484
rect 282178 367140 282184 367192
rect 282236 367180 282242 367192
rect 282273 367183 282331 367189
rect 282273 367180 282285 367183
rect 282236 367152 282285 367180
rect 282236 367140 282242 367152
rect 282273 367149 282285 367152
rect 282319 367149 282331 367183
rect 282273 367143 282331 367149
rect 282086 367004 282092 367056
rect 282144 367004 282150 367056
rect 284478 367004 284484 367056
rect 284536 367044 284542 367056
rect 312538 367044 312544 367056
rect 284536 367016 312544 367044
rect 284536 367004 284542 367016
rect 312538 367004 312544 367016
rect 312596 367004 312602 367056
rect 282104 366917 282132 367004
rect 285122 366936 285128 366988
rect 285180 366976 285186 366988
rect 309778 366976 309784 366988
rect 285180 366948 309784 366976
rect 285180 366936 285186 366948
rect 309778 366936 309784 366948
rect 309836 366936 309842 366988
rect 282089 366911 282147 366917
rect 282089 366877 282101 366911
rect 282135 366877 282147 366911
rect 282089 366871 282147 366877
rect 281626 365644 281632 365696
rect 281684 365684 281690 365696
rect 330478 365684 330484 365696
rect 281684 365656 330484 365684
rect 281684 365644 281690 365656
rect 330478 365644 330484 365656
rect 330536 365644 330542 365696
rect 282270 364964 282276 365016
rect 282328 365004 282334 365016
rect 282730 365004 282736 365016
rect 282328 364976 282736 365004
rect 282328 364964 282334 364976
rect 282730 364964 282736 364976
rect 282788 364964 282794 365016
rect 281626 364284 281632 364336
rect 281684 364324 281690 364336
rect 329282 364324 329288 364336
rect 281684 364296 329288 364324
rect 281684 364284 281690 364296
rect 329282 364284 329288 364296
rect 329340 364284 329346 364336
rect 281626 362856 281632 362908
rect 281684 362896 281690 362908
rect 329098 362896 329104 362908
rect 281684 362868 329104 362896
rect 281684 362856 281690 362868
rect 329098 362856 329104 362868
rect 329156 362856 329162 362908
rect 281810 362788 281816 362840
rect 281868 362828 281874 362840
rect 327718 362828 327724 362840
rect 281868 362800 327724 362828
rect 281868 362788 281874 362800
rect 327718 362788 327724 362800
rect 327776 362788 327782 362840
rect 281626 361496 281632 361548
rect 281684 361536 281690 361548
rect 326338 361536 326344 361548
rect 281684 361508 326344 361536
rect 281684 361496 281690 361508
rect 326338 361496 326344 361508
rect 326396 361496 326402 361548
rect 281626 360136 281632 360188
rect 281684 360176 281690 360188
rect 324958 360176 324964 360188
rect 281684 360148 324964 360176
rect 281684 360136 281690 360148
rect 324958 360136 324964 360148
rect 325016 360136 325022 360188
rect 281810 360068 281816 360120
rect 281868 360108 281874 360120
rect 323578 360108 323584 360120
rect 281868 360080 323584 360108
rect 281868 360068 281874 360080
rect 323578 360068 323584 360080
rect 323636 360068 323642 360120
rect 281626 358708 281632 358760
rect 281684 358748 281690 358760
rect 322198 358748 322204 358760
rect 281684 358720 322204 358748
rect 281684 358708 281690 358720
rect 322198 358708 322204 358720
rect 322256 358708 322262 358760
rect 282089 357459 282147 357465
rect 282089 357425 282101 357459
rect 282135 357456 282147 357459
rect 282178 357456 282184 357468
rect 282135 357428 282184 357456
rect 282135 357425 282147 357428
rect 282089 357419 282147 357425
rect 282178 357416 282184 357428
rect 282236 357416 282242 357468
rect 281626 351772 281632 351824
rect 281684 351812 281690 351824
rect 286502 351812 286508 351824
rect 281684 351784 286508 351812
rect 281684 351772 281690 351784
rect 286502 351772 286508 351784
rect 286560 351772 286566 351824
rect 281626 350888 281632 350940
rect 281684 350928 281690 350940
rect 286410 350928 286416 350940
rect 281684 350900 286416 350928
rect 281684 350888 281690 350900
rect 286410 350888 286416 350900
rect 286468 350888 286474 350940
rect 281626 350276 281632 350328
rect 281684 350316 281690 350328
rect 284570 350316 284576 350328
rect 281684 350288 284576 350316
rect 281684 350276 281690 350288
rect 284570 350276 284576 350288
rect 284628 350276 284634 350328
rect 281626 349052 281632 349104
rect 281684 349092 281690 349104
rect 291838 349092 291844 349104
rect 281684 349064 291844 349092
rect 281684 349052 281690 349064
rect 291838 349052 291844 349064
rect 291896 349052 291902 349104
rect 281626 347692 281632 347744
rect 281684 347732 281690 347744
rect 290458 347732 290464 347744
rect 281684 347704 290464 347732
rect 281684 347692 281690 347704
rect 290458 347692 290464 347704
rect 290516 347692 290522 347744
rect 281626 346740 281632 346792
rect 281684 346780 281690 346792
rect 287698 346780 287704 346792
rect 281684 346752 287704 346780
rect 281684 346740 281690 346752
rect 287698 346740 287704 346752
rect 287756 346740 287762 346792
rect 281626 345652 281632 345704
rect 281684 345692 281690 345704
rect 286318 345692 286324 345704
rect 281684 345664 286324 345692
rect 281684 345652 281690 345664
rect 286318 345652 286324 345664
rect 286376 345652 286382 345704
rect 281626 344836 281632 344888
rect 281684 344876 281690 344888
rect 284938 344876 284944 344888
rect 281684 344848 284944 344876
rect 281684 344836 281690 344848
rect 284938 344836 284944 344848
rect 284996 344836 285002 344888
rect 281626 343544 281632 343596
rect 281684 343584 281690 343596
rect 307018 343584 307024 343596
rect 281684 343556 307024 343584
rect 281684 343544 281690 343556
rect 307018 343544 307024 343556
rect 307076 343544 307082 343596
rect 281810 343476 281816 343528
rect 281868 343516 281874 343528
rect 291930 343516 291936 343528
rect 281868 343488 291936 343516
rect 281868 343476 281874 343488
rect 291930 343476 291936 343488
rect 291988 343476 291994 343528
rect 281626 342184 281632 342236
rect 281684 342224 281690 342236
rect 308398 342224 308404 342236
rect 281684 342196 308404 342224
rect 281684 342184 281690 342196
rect 308398 342184 308404 342196
rect 308456 342184 308462 342236
rect 282270 340824 282276 340876
rect 282328 340864 282334 340876
rect 282454 340864 282460 340876
rect 282328 340836 282460 340864
rect 282328 340824 282334 340836
rect 282454 340824 282460 340836
rect 282512 340824 282518 340876
rect 281626 340756 281632 340808
rect 281684 340796 281690 340808
rect 284754 340796 284760 340808
rect 281684 340768 284760 340796
rect 281684 340756 281690 340768
rect 284754 340756 284760 340768
rect 284812 340756 284818 340808
rect 281718 340620 281724 340672
rect 281776 340660 281782 340672
rect 284662 340660 284668 340672
rect 281776 340632 284668 340660
rect 281776 340620 281782 340632
rect 284662 340620 284668 340632
rect 284720 340620 284726 340672
rect 281626 338784 281632 338836
rect 281684 338824 281690 338836
rect 284846 338824 284852 338836
rect 281684 338796 284852 338824
rect 281684 338784 281690 338796
rect 284846 338784 284852 338796
rect 284904 338784 284910 338836
rect 282365 338079 282423 338085
rect 282365 338045 282377 338079
rect 282411 338076 282423 338079
rect 282454 338076 282460 338088
rect 282411 338048 282460 338076
rect 282411 338045 282423 338048
rect 282365 338039 282423 338045
rect 282454 338036 282460 338048
rect 282512 338036 282518 338088
rect 281626 337900 281632 337952
rect 281684 337940 281690 337952
rect 285582 337940 285588 337952
rect 281684 337912 285588 337940
rect 281684 337900 281690 337912
rect 285582 337900 285588 337912
rect 285640 337900 285646 337952
rect 281718 336676 281724 336728
rect 281776 336716 281782 336728
rect 285398 336716 285404 336728
rect 281776 336688 285404 336716
rect 281776 336676 281782 336688
rect 285398 336676 285404 336688
rect 285456 336676 285462 336728
rect 281626 336540 281632 336592
rect 281684 336580 281690 336592
rect 285490 336580 285496 336592
rect 281684 336552 285496 336580
rect 281684 336540 281690 336552
rect 285490 336540 285496 336552
rect 285548 336540 285554 336592
rect 281626 334568 281632 334620
rect 281684 334608 281690 334620
rect 285306 334608 285312 334620
rect 281684 334580 285312 334608
rect 281684 334568 281690 334580
rect 285306 334568 285312 334580
rect 285364 334568 285370 334620
rect 281718 333888 281724 333940
rect 281776 333928 281782 333940
rect 302878 333928 302884 333940
rect 281776 333900 302884 333928
rect 281776 333888 281782 333900
rect 302878 333888 302884 333900
rect 302936 333888 302942 333940
rect 281626 333616 281632 333668
rect 281684 333656 281690 333668
rect 285214 333656 285220 333668
rect 281684 333628 285220 333656
rect 281684 333616 281690 333628
rect 285214 333616 285220 333628
rect 285272 333616 285278 333668
rect 281626 331168 281632 331220
rect 281684 331208 281690 331220
rect 320266 331208 320272 331220
rect 281684 331180 320272 331208
rect 281684 331168 281690 331180
rect 320266 331168 320272 331180
rect 320324 331168 320330 331220
rect 281534 329740 281540 329792
rect 281592 329780 281598 329792
rect 320174 329780 320180 329792
rect 281592 329752 320180 329780
rect 281592 329740 281598 329752
rect 320174 329740 320180 329752
rect 320232 329740 320238 329792
rect 281626 329672 281632 329724
rect 281684 329712 281690 329724
rect 318794 329712 318800 329724
rect 281684 329684 318800 329712
rect 281684 329672 281690 329684
rect 318794 329672 318800 329684
rect 318852 329672 318858 329724
rect 282362 328488 282368 328500
rect 282323 328460 282368 328488
rect 282362 328448 282368 328460
rect 282420 328448 282426 328500
rect 281534 328380 281540 328432
rect 281592 328420 281598 328432
rect 317414 328420 317420 328432
rect 281592 328392 317420 328420
rect 281592 328380 281598 328392
rect 317414 328380 317420 328392
rect 317472 328380 317478 328432
rect 281534 325524 281540 325576
rect 281592 325564 281598 325576
rect 285030 325564 285036 325576
rect 281592 325536 285036 325564
rect 281592 325524 281598 325536
rect 285030 325524 285036 325536
rect 285088 325524 285094 325576
rect 282822 321512 282828 321564
rect 282880 321552 282886 321564
rect 338758 321552 338764 321564
rect 282880 321524 338764 321552
rect 282880 321512 282886 321524
rect 338758 321512 338764 321524
rect 338816 321512 338822 321564
rect 44082 318724 44088 318776
rect 44140 318764 44146 318776
rect 130930 318764 130936 318776
rect 44140 318736 130936 318764
rect 44140 318724 44146 318736
rect 130930 318724 130936 318736
rect 130988 318724 130994 318776
rect 131025 318767 131083 318773
rect 131025 318733 131037 318767
rect 131071 318764 131083 318767
rect 132862 318764 132868 318776
rect 131071 318736 132868 318764
rect 131071 318733 131083 318736
rect 131025 318727 131083 318733
rect 132862 318724 132868 318736
rect 132920 318724 132926 318776
rect 133138 318724 133144 318776
rect 133196 318764 133202 318776
rect 249702 318764 249708 318776
rect 133196 318736 249708 318764
rect 133196 318724 133202 318736
rect 249702 318724 249708 318736
rect 249760 318724 249766 318776
rect 343634 318724 343640 318776
rect 343692 318764 343698 318776
rect 420178 318764 420184 318776
rect 343692 318736 420184 318764
rect 343692 318724 343698 318736
rect 420178 318724 420184 318736
rect 420236 318764 420242 318776
rect 453114 318764 453120 318776
rect 420236 318736 453120 318764
rect 420236 318724 420242 318736
rect 453114 318724 453120 318736
rect 453172 318724 453178 318776
rect 20622 318656 20628 318708
rect 20680 318696 20686 318708
rect 92014 318696 92020 318708
rect 20680 318668 92020 318696
rect 20680 318656 20686 318668
rect 92014 318656 92020 318668
rect 92072 318656 92078 318708
rect 92382 318656 92388 318708
rect 92440 318696 92446 318708
rect 210786 318696 210792 318708
rect 92440 318668 210792 318696
rect 92440 318656 92446 318668
rect 210786 318656 210792 318668
rect 210844 318656 210850 318708
rect 22002 318588 22008 318640
rect 22060 318628 22066 318640
rect 93946 318628 93952 318640
rect 22060 318600 93952 318628
rect 22060 318588 22066 318600
rect 93946 318588 93952 318600
rect 94004 318588 94010 318640
rect 96522 318588 96528 318640
rect 96580 318628 96586 318640
rect 97721 318631 97779 318637
rect 97721 318628 97733 318631
rect 96580 318600 97733 318628
rect 96580 318588 96586 318600
rect 97721 318597 97733 318600
rect 97767 318597 97779 318631
rect 97721 318591 97779 318597
rect 98089 318631 98147 318637
rect 98089 318597 98101 318631
rect 98135 318628 98147 318631
rect 216582 318628 216588 318640
rect 98135 318600 216588 318628
rect 98135 318597 98147 318600
rect 98089 318591 98147 318597
rect 216582 318588 216588 318600
rect 216640 318588 216646 318640
rect 23382 318520 23388 318572
rect 23440 318560 23446 318572
rect 97902 318560 97908 318572
rect 23440 318532 97908 318560
rect 23440 318520 23446 318532
rect 97902 318520 97908 318532
rect 97960 318520 97966 318572
rect 97994 318520 98000 318572
rect 98052 318560 98058 318572
rect 218514 318560 218520 318572
rect 98052 318532 218520 318560
rect 98052 318520 98058 318532
rect 218514 318520 218520 318532
rect 218572 318520 218578 318572
rect 30282 318452 30288 318504
rect 30340 318492 30346 318504
rect 107562 318492 107568 318504
rect 30340 318464 107568 318492
rect 30340 318452 30346 318464
rect 107562 318452 107568 318464
rect 107620 318452 107626 318504
rect 107654 318452 107660 318504
rect 107712 318492 107718 318504
rect 234154 318492 234160 318504
rect 107712 318464 234160 318492
rect 107712 318452 107718 318464
rect 234154 318452 234160 318464
rect 234212 318452 234218 318504
rect 28902 318384 28908 318436
rect 28960 318424 28966 318436
rect 105630 318424 105636 318436
rect 28960 318396 105636 318424
rect 28960 318384 28966 318396
rect 105630 318384 105636 318396
rect 105688 318384 105694 318436
rect 110322 318384 110328 318436
rect 110380 318424 110386 318436
rect 239950 318424 239956 318436
rect 110380 318396 239956 318424
rect 110380 318384 110386 318396
rect 239950 318384 239956 318396
rect 240008 318384 240014 318436
rect 31662 318316 31668 318368
rect 31720 318356 31726 318368
rect 111518 318356 111524 318368
rect 31720 318328 111524 318356
rect 31720 318316 31726 318328
rect 111518 318316 111524 318328
rect 111576 318316 111582 318368
rect 111702 318316 111708 318368
rect 111760 318356 111766 318368
rect 241882 318356 241888 318368
rect 111760 318328 241888 318356
rect 111760 318316 111766 318328
rect 241882 318316 241888 318328
rect 241940 318316 241946 318368
rect 42702 318248 42708 318300
rect 42760 318288 42766 318300
rect 128998 318288 129004 318300
rect 42760 318260 129004 318288
rect 42760 318248 42766 318260
rect 128998 318248 129004 318260
rect 129056 318248 129062 318300
rect 130378 318248 130384 318300
rect 130436 318288 130442 318300
rect 261386 318288 261392 318300
rect 130436 318260 261392 318288
rect 130436 318248 130442 318260
rect 261386 318248 261392 318260
rect 261444 318248 261450 318300
rect 35802 318180 35808 318232
rect 35860 318220 35866 318232
rect 117314 318220 117320 318232
rect 35860 318192 117320 318220
rect 35860 318180 35866 318192
rect 117314 318180 117320 318192
rect 117372 318180 117378 318232
rect 118602 318180 118608 318232
rect 118660 318220 118666 318232
rect 253566 318220 253572 318232
rect 118660 318192 253572 318220
rect 118660 318180 118666 318192
rect 253566 318180 253572 318192
rect 253624 318180 253630 318232
rect 39942 318112 39948 318164
rect 40000 318152 40006 318164
rect 125134 318152 125140 318164
rect 40000 318124 125140 318152
rect 40000 318112 40006 318124
rect 125134 318112 125140 318124
rect 125192 318112 125198 318164
rect 125502 318112 125508 318164
rect 125560 318152 125566 318164
rect 265250 318152 265256 318164
rect 125560 318124 265256 318152
rect 125560 318112 125566 318124
rect 265250 318112 265256 318124
rect 265308 318112 265314 318164
rect 61378 318044 61384 318096
rect 61436 318084 61442 318096
rect 343634 318084 343640 318096
rect 61436 318056 343640 318084
rect 61436 318044 61442 318056
rect 343634 318044 343640 318056
rect 343692 318044 343698 318096
rect 16482 317976 16488 318028
rect 16540 318016 16546 318028
rect 86218 318016 86224 318028
rect 16540 317988 86224 318016
rect 16540 317976 16546 317988
rect 86218 317976 86224 317988
rect 86276 317976 86282 318028
rect 90910 317976 90916 318028
rect 90968 318016 90974 318028
rect 206830 318016 206836 318028
rect 90968 317988 206836 318016
rect 90968 317976 90974 317988
rect 206830 317976 206836 317988
rect 206888 317976 206894 318028
rect 12342 317908 12348 317960
rect 12400 317948 12406 317960
rect 78398 317948 78404 317960
rect 12400 317920 78404 317948
rect 12400 317908 12406 317920
rect 78398 317908 78404 317920
rect 78456 317908 78462 317960
rect 79962 317908 79968 317960
rect 80020 317948 80026 317960
rect 189350 317948 189356 317960
rect 80020 317920 189356 317948
rect 80020 317908 80026 317920
rect 189350 317908 189356 317920
rect 189408 317908 189414 317960
rect 5442 317840 5448 317892
rect 5500 317880 5506 317892
rect 68646 317880 68652 317892
rect 5500 317852 68652 317880
rect 5500 317840 5506 317852
rect 68646 317840 68652 317852
rect 68704 317840 68710 317892
rect 72970 317840 72976 317892
rect 73028 317880 73034 317892
rect 177666 317880 177672 317892
rect 73028 317852 177672 317880
rect 73028 317840 73034 317852
rect 177666 317840 177672 317852
rect 177724 317840 177730 317892
rect 57882 317772 57888 317824
rect 57940 317812 57946 317824
rect 154298 317812 154304 317824
rect 57940 317784 154304 317812
rect 57940 317772 57946 317784
rect 154298 317772 154304 317784
rect 154356 317772 154362 317824
rect 53742 317704 53748 317756
rect 53800 317744 53806 317756
rect 146570 317744 146576 317756
rect 53800 317716 146576 317744
rect 53800 317704 53806 317716
rect 146570 317704 146576 317716
rect 146628 317704 146634 317756
rect 50982 317636 50988 317688
rect 51040 317676 51046 317688
rect 142614 317676 142620 317688
rect 51040 317648 142620 317676
rect 51040 317636 51046 317648
rect 142614 317636 142620 317648
rect 142672 317636 142678 317688
rect 48130 317568 48136 317620
rect 48188 317608 48194 317620
rect 136818 317608 136824 317620
rect 48188 317580 136824 317608
rect 48188 317568 48194 317580
rect 136818 317568 136824 317580
rect 136876 317568 136882 317620
rect 38470 317500 38476 317552
rect 38528 317540 38534 317552
rect 123202 317540 123208 317552
rect 38528 317512 123208 317540
rect 38528 317500 38534 317512
rect 123202 317500 123208 317512
rect 123260 317500 123266 317552
rect 123478 317500 123484 317552
rect 123536 317540 123542 317552
rect 131025 317543 131083 317549
rect 131025 317540 131037 317543
rect 123536 317512 131037 317540
rect 123536 317500 123542 317512
rect 131025 317509 131037 317512
rect 131071 317509 131083 317543
rect 131025 317503 131083 317509
rect 131758 317500 131764 317552
rect 131816 317540 131822 317552
rect 169846 317540 169852 317552
rect 131816 317512 169852 317540
rect 131816 317500 131822 317512
rect 169846 317500 169852 317512
rect 169904 317500 169910 317552
rect 33042 317432 33048 317484
rect 33100 317472 33106 317484
rect 113450 317472 113456 317484
rect 33100 317444 113456 317472
rect 33100 317432 33106 317444
rect 113450 317432 113456 317444
rect 113508 317432 113514 317484
rect 124858 317432 124864 317484
rect 124916 317472 124922 317484
rect 158162 317472 158168 317484
rect 124916 317444 158168 317472
rect 124916 317432 124922 317444
rect 158162 317432 158168 317444
rect 158220 317432 158226 317484
rect 49326 6128 49332 6180
rect 49384 6168 49390 6180
rect 139394 6168 139400 6180
rect 49384 6140 139400 6168
rect 49384 6128 49390 6140
rect 139394 6128 139400 6140
rect 139452 6128 139458 6180
rect 80238 5448 80244 5500
rect 80296 5488 80302 5500
rect 190454 5488 190460 5500
rect 80296 5460 190460 5488
rect 80296 5448 80302 5460
rect 190454 5448 190460 5460
rect 190512 5448 190518 5500
rect 83826 5380 83832 5432
rect 83884 5420 83890 5432
rect 195974 5420 195980 5432
rect 83884 5392 195980 5420
rect 83884 5380 83890 5392
rect 195974 5380 195980 5392
rect 196032 5380 196038 5432
rect 87322 5312 87328 5364
rect 87380 5352 87386 5364
rect 202874 5352 202880 5364
rect 87380 5324 202880 5352
rect 87380 5312 87386 5324
rect 202874 5312 202880 5324
rect 202932 5312 202938 5364
rect 91002 5244 91008 5296
rect 91060 5284 91066 5296
rect 208394 5284 208400 5296
rect 91060 5256 208400 5284
rect 91060 5244 91066 5256
rect 208394 5244 208400 5256
rect 208452 5244 208458 5296
rect 94498 5176 94504 5228
rect 94556 5216 94562 5228
rect 213914 5216 213920 5228
rect 94556 5188 213920 5216
rect 94556 5176 94562 5188
rect 213914 5176 213920 5188
rect 213972 5176 213978 5228
rect 98086 5108 98092 5160
rect 98144 5148 98150 5160
rect 219434 5148 219440 5160
rect 98144 5120 219440 5148
rect 98144 5108 98150 5120
rect 219434 5108 219440 5120
rect 219492 5108 219498 5160
rect 101582 5040 101588 5092
rect 101640 5080 101646 5092
rect 226334 5080 226340 5092
rect 101640 5052 226340 5080
rect 101640 5040 101646 5052
rect 226334 5040 226340 5052
rect 226392 5040 226398 5092
rect 105170 4972 105176 5024
rect 105228 5012 105234 5024
rect 231854 5012 231860 5024
rect 105228 4984 231860 5012
rect 105228 4972 105234 4984
rect 231854 4972 231860 4984
rect 231912 4972 231918 5024
rect 67174 4904 67180 4956
rect 67232 4944 67238 4956
rect 131758 4944 131764 4956
rect 67232 4916 131764 4944
rect 67232 4904 67238 4916
rect 131758 4904 131764 4916
rect 131816 4904 131822 4956
rect 131853 4947 131911 4953
rect 131853 4913 131865 4947
rect 131899 4944 131911 4947
rect 266354 4944 266360 4956
rect 131899 4916 266360 4944
rect 131899 4913 131911 4916
rect 131853 4907 131911 4913
rect 266354 4904 266360 4916
rect 266412 4904 266418 4956
rect 59998 4836 60004 4888
rect 60056 4876 60062 4888
rect 124858 4876 124864 4888
rect 60056 4848 124864 4876
rect 60056 4836 60062 4848
rect 124858 4836 124864 4848
rect 124916 4836 124922 4888
rect 126606 4836 126612 4888
rect 126664 4876 126670 4888
rect 130105 4879 130163 4885
rect 130105 4876 130117 4879
rect 126664 4848 130117 4876
rect 126664 4836 126670 4848
rect 130105 4845 130117 4848
rect 130151 4845 130163 4879
rect 130105 4839 130163 4845
rect 130194 4836 130200 4888
rect 130252 4876 130258 4888
rect 271874 4876 271880 4888
rect 130252 4848 271880 4876
rect 130252 4836 130258 4848
rect 271874 4836 271880 4848
rect 271932 4836 271938 4888
rect 37366 4768 37372 4820
rect 37424 4808 37430 4820
rect 120074 4808 120080 4820
rect 37424 4780 120080 4808
rect 37424 4768 37430 4780
rect 120074 4768 120080 4780
rect 120132 4768 120138 4820
rect 123018 4768 123024 4820
rect 123076 4808 123082 4820
rect 130378 4808 130384 4820
rect 123076 4780 130384 4808
rect 123076 4768 123082 4780
rect 130378 4768 130384 4780
rect 130436 4768 130442 4820
rect 130473 4811 130531 4817
rect 130473 4777 130485 4811
rect 130519 4808 130531 4811
rect 131301 4811 131359 4817
rect 131301 4808 131313 4811
rect 130519 4780 131313 4808
rect 130519 4777 130531 4780
rect 130473 4771 130531 4777
rect 131301 4777 131313 4780
rect 131347 4777 131359 4811
rect 131301 4771 131359 4777
rect 131390 4768 131396 4820
rect 131448 4808 131454 4820
rect 274634 4808 274640 4820
rect 131448 4780 274640 4808
rect 131448 4768 131454 4780
rect 274634 4768 274640 4780
rect 274692 4768 274698 4820
rect 76650 4700 76656 4752
rect 76708 4740 76714 4752
rect 184934 4740 184940 4752
rect 76708 4712 184940 4740
rect 76708 4700 76714 4712
rect 184934 4700 184940 4712
rect 184992 4700 184998 4752
rect 73062 4632 73068 4684
rect 73120 4672 73126 4684
rect 179414 4672 179420 4684
rect 73120 4644 179420 4672
rect 73120 4632 73126 4644
rect 179414 4632 179420 4644
rect 179472 4632 179478 4684
rect 69474 4564 69480 4616
rect 69532 4604 69538 4616
rect 172514 4604 172520 4616
rect 69532 4576 172520 4604
rect 69532 4564 69538 4576
rect 172514 4564 172520 4576
rect 172572 4564 172578 4616
rect 55217 4539 55275 4545
rect 55217 4505 55229 4539
rect 55263 4536 55275 4539
rect 64785 4539 64843 4545
rect 64785 4536 64797 4539
rect 55263 4508 64797 4536
rect 55263 4505 55275 4508
rect 55217 4499 55275 4505
rect 64785 4505 64797 4508
rect 64831 4505 64843 4539
rect 64785 4499 64843 4505
rect 65978 4496 65984 4548
rect 66036 4536 66042 4548
rect 166994 4536 167000 4548
rect 66036 4508 167000 4536
rect 66036 4496 66042 4508
rect 166994 4496 167000 4508
rect 167052 4496 167058 4548
rect 62390 4428 62396 4480
rect 62448 4468 62454 4480
rect 161474 4468 161480 4480
rect 62448 4440 161480 4468
rect 62448 4428 62454 4440
rect 161474 4428 161480 4440
rect 161532 4428 161538 4480
rect 58802 4360 58808 4412
rect 58860 4400 58866 4412
rect 155954 4400 155960 4412
rect 58860 4372 155960 4400
rect 58860 4360 58866 4372
rect 155954 4360 155960 4372
rect 156012 4360 156018 4412
rect 55214 4292 55220 4344
rect 55272 4332 55278 4344
rect 150434 4332 150440 4344
rect 55272 4304 150440 4332
rect 55272 4292 55278 4304
rect 150434 4292 150440 4304
rect 150492 4292 150498 4344
rect 51626 4224 51632 4276
rect 51684 4264 51690 4276
rect 143534 4264 143540 4276
rect 51684 4236 143540 4264
rect 51684 4224 51690 4236
rect 143534 4224 143540 4236
rect 143592 4224 143598 4276
rect 46934 4156 46940 4208
rect 46992 4196 46998 4208
rect 48130 4196 48136 4208
rect 46992 4168 48136 4196
rect 46992 4156 46998 4168
rect 48130 4156 48136 4168
rect 48188 4156 48194 4208
rect 48222 4156 48228 4208
rect 48280 4196 48286 4208
rect 138014 4196 138020 4208
rect 48280 4168 138020 4196
rect 48280 4156 48286 4168
rect 138014 4156 138020 4168
rect 138072 4156 138078 4208
rect 16577 4131 16635 4137
rect 16577 4097 16589 4131
rect 16623 4128 16635 4131
rect 55217 4131 55275 4137
rect 55217 4128 55229 4131
rect 16623 4100 55229 4128
rect 16623 4097 16635 4100
rect 16577 4091 16635 4097
rect 55217 4097 55229 4100
rect 55263 4097 55275 4131
rect 55217 4091 55275 4097
rect 64785 4131 64843 4137
rect 64785 4097 64797 4131
rect 64831 4128 64843 4131
rect 81342 4128 81348 4140
rect 64831 4100 81348 4128
rect 64831 4097 64843 4100
rect 64785 4091 64843 4097
rect 81342 4088 81348 4100
rect 81400 4088 81406 4140
rect 84841 4131 84899 4137
rect 84841 4097 84853 4131
rect 84887 4128 84899 4131
rect 89714 4128 89720 4140
rect 84887 4100 89720 4128
rect 84887 4097 84899 4100
rect 84841 4091 84899 4097
rect 89714 4088 89720 4100
rect 89772 4088 89778 4140
rect 93302 4088 93308 4140
rect 93360 4128 93366 4140
rect 212534 4128 212540 4140
rect 93360 4100 212540 4128
rect 93360 4088 93366 4100
rect 212534 4088 212540 4100
rect 212592 4088 212598 4140
rect 14826 4020 14832 4072
rect 14884 4060 14890 4072
rect 55306 4060 55312 4072
rect 14884 4032 55312 4060
rect 14884 4020 14890 4032
rect 55306 4020 55312 4032
rect 55364 4020 55370 4072
rect 64690 4020 64696 4072
rect 64748 4060 64754 4072
rect 80057 4063 80115 4069
rect 80057 4060 80069 4063
rect 64748 4032 80069 4060
rect 64748 4020 64754 4032
rect 80057 4029 80069 4032
rect 80103 4029 80115 4063
rect 80057 4023 80115 4029
rect 81434 4020 81440 4072
rect 81492 4060 81498 4072
rect 82630 4060 82636 4072
rect 81492 4032 82636 4060
rect 81492 4020 81498 4032
rect 82630 4020 82636 4032
rect 82688 4020 82694 4072
rect 108301 4063 108359 4069
rect 108301 4029 108313 4063
rect 108347 4060 108359 4063
rect 223574 4060 223580 4072
rect 108347 4032 223580 4060
rect 108347 4029 108359 4032
rect 108301 4023 108359 4029
rect 223574 4020 223580 4032
rect 223632 4020 223638 4072
rect 13630 3952 13636 4004
rect 13688 3992 13694 4004
rect 16577 3995 16635 4001
rect 16577 3992 16589 3995
rect 13688 3964 16589 3992
rect 13688 3952 13694 3964
rect 16577 3961 16589 3964
rect 16623 3961 16635 3995
rect 16577 3955 16635 3961
rect 17218 3952 17224 4004
rect 17276 3992 17282 4004
rect 86954 3992 86960 4004
rect 17276 3964 86960 3992
rect 17276 3952 17282 3964
rect 86954 3952 86960 3964
rect 87012 3952 87018 4004
rect 99282 3952 99288 4004
rect 99340 3992 99346 4004
rect 222194 3992 222200 4004
rect 99340 3964 222200 3992
rect 99340 3952 99346 3964
rect 222194 3952 222200 3964
rect 222252 3952 222258 4004
rect 18322 3884 18328 3936
rect 18380 3924 18386 3936
rect 84841 3927 84899 3933
rect 84841 3924 84853 3927
rect 18380 3896 84853 3924
rect 18380 3884 18386 3896
rect 84841 3893 84853 3896
rect 84887 3893 84899 3927
rect 84841 3887 84899 3893
rect 84930 3884 84936 3936
rect 84988 3924 84994 3936
rect 91281 3927 91339 3933
rect 91281 3924 91293 3927
rect 84988 3896 91293 3924
rect 84988 3884 84994 3896
rect 91281 3893 91293 3896
rect 91327 3893 91339 3927
rect 91281 3887 91339 3893
rect 102778 3884 102784 3936
rect 102836 3924 102842 3936
rect 227714 3924 227720 3936
rect 102836 3896 227720 3924
rect 102836 3884 102842 3896
rect 227714 3884 227720 3896
rect 227772 3884 227778 3936
rect 19518 3816 19524 3868
rect 19576 3856 19582 3868
rect 20622 3856 20628 3868
rect 19576 3828 20628 3856
rect 19576 3816 19582 3828
rect 20622 3816 20628 3828
rect 20680 3816 20686 3868
rect 20714 3816 20720 3868
rect 20772 3856 20778 3868
rect 22002 3856 22008 3868
rect 20772 3828 22008 3856
rect 20772 3816 20778 3828
rect 22002 3816 22008 3828
rect 22060 3816 22066 3868
rect 95234 3856 95240 3868
rect 22112 3828 95240 3856
rect 21910 3748 21916 3800
rect 21968 3788 21974 3800
rect 22112 3788 22140 3828
rect 95234 3816 95240 3828
rect 95292 3816 95298 3868
rect 95605 3859 95663 3865
rect 95605 3825 95617 3859
rect 95651 3856 95663 3859
rect 99374 3856 99380 3868
rect 95651 3828 99380 3856
rect 95651 3825 95663 3828
rect 95605 3819 95663 3825
rect 99374 3816 99380 3828
rect 99432 3816 99438 3868
rect 100478 3816 100484 3868
rect 100536 3856 100542 3868
rect 108301 3859 108359 3865
rect 108301 3856 108313 3859
rect 100536 3828 108313 3856
rect 100536 3816 100542 3828
rect 108301 3825 108313 3828
rect 108347 3825 108359 3859
rect 235994 3856 236000 3868
rect 108301 3819 108359 3825
rect 109880 3828 236000 3856
rect 21968 3760 22140 3788
rect 21968 3748 21974 3760
rect 25498 3748 25504 3800
rect 25556 3788 25562 3800
rect 100754 3788 100760 3800
rect 25556 3760 100760 3788
rect 25556 3748 25562 3760
rect 100754 3748 100760 3760
rect 100812 3748 100818 3800
rect 107470 3748 107476 3800
rect 107528 3788 107534 3800
rect 109880 3788 109908 3828
rect 235994 3816 236000 3828
rect 236052 3816 236058 3868
rect 107528 3760 109908 3788
rect 107528 3748 107534 3760
rect 114738 3748 114744 3800
rect 114796 3788 114802 3800
rect 247034 3788 247040 3800
rect 114796 3760 247040 3788
rect 114796 3748 114802 3760
rect 247034 3748 247040 3760
rect 247092 3748 247098 3800
rect 24302 3680 24308 3732
rect 24360 3720 24366 3732
rect 95605 3723 95663 3729
rect 95605 3720 95617 3723
rect 24360 3692 95617 3720
rect 24360 3680 24366 3692
rect 95605 3689 95617 3692
rect 95651 3689 95663 3723
rect 95605 3683 95663 3689
rect 95694 3680 95700 3732
rect 95752 3720 95758 3732
rect 96522 3720 96528 3732
rect 95752 3692 96528 3720
rect 95752 3680 95758 3692
rect 96522 3680 96528 3692
rect 96580 3680 96586 3732
rect 96890 3680 96896 3732
rect 96948 3720 96954 3732
rect 97902 3720 97908 3732
rect 96948 3692 97908 3720
rect 96948 3680 96954 3692
rect 97902 3680 97908 3692
rect 97960 3680 97966 3732
rect 113542 3680 113548 3732
rect 113600 3720 113606 3732
rect 245654 3720 245660 3732
rect 113600 3692 245660 3720
rect 113600 3680 113606 3692
rect 245654 3680 245660 3692
rect 245712 3680 245718 3732
rect 26694 3612 26700 3664
rect 26752 3652 26758 3664
rect 103514 3652 103520 3664
rect 26752 3624 103520 3652
rect 26752 3612 26758 3624
rect 103514 3612 103520 3624
rect 103572 3612 103578 3664
rect 109034 3652 109040 3664
rect 103900 3624 109040 3652
rect 34974 3544 34980 3596
rect 35032 3584 35038 3596
rect 35802 3584 35808 3596
rect 35032 3556 35808 3584
rect 35032 3544 35038 3556
rect 35802 3544 35808 3556
rect 35860 3544 35866 3596
rect 35897 3587 35955 3593
rect 35897 3553 35909 3587
rect 35943 3584 35955 3587
rect 103900 3584 103928 3624
rect 109034 3612 109040 3624
rect 109092 3612 109098 3664
rect 117130 3612 117136 3664
rect 117188 3652 117194 3664
rect 251174 3652 251180 3664
rect 117188 3624 251180 3652
rect 117188 3612 117194 3624
rect 251174 3612 251180 3624
rect 251232 3612 251238 3664
rect 35943 3556 103928 3584
rect 35943 3553 35955 3556
rect 35897 3547 35955 3553
rect 103974 3544 103980 3596
rect 104032 3584 104038 3596
rect 104802 3584 104808 3596
rect 104032 3556 104808 3584
rect 104032 3544 104038 3556
rect 104802 3544 104808 3556
rect 104860 3544 104866 3596
rect 106366 3544 106372 3596
rect 106424 3584 106430 3596
rect 107562 3584 107568 3596
rect 106424 3556 107568 3584
rect 106424 3544 106430 3556
rect 107562 3544 107568 3556
rect 107620 3544 107626 3596
rect 111150 3544 111156 3596
rect 111208 3584 111214 3596
rect 111702 3584 111708 3596
rect 111208 3556 111708 3584
rect 111208 3544 111214 3556
rect 111702 3544 111708 3556
rect 111760 3544 111766 3596
rect 119430 3544 119436 3596
rect 119488 3584 119494 3596
rect 255314 3584 255320 3596
rect 119488 3556 255320 3584
rect 119488 3544 119494 3556
rect 255314 3544 255320 3556
rect 255372 3544 255378 3596
rect 11238 3476 11244 3528
rect 11296 3516 11302 3528
rect 12342 3516 12348 3528
rect 11296 3488 12348 3516
rect 11296 3476 11302 3488
rect 12342 3476 12348 3488
rect 12400 3476 12406 3528
rect 16022 3476 16028 3528
rect 16080 3516 16086 3528
rect 16482 3516 16488 3528
rect 16080 3488 16488 3516
rect 16080 3476 16086 3488
rect 16482 3476 16488 3488
rect 16540 3476 16546 3528
rect 27890 3476 27896 3528
rect 27948 3516 27954 3528
rect 28902 3516 28908 3528
rect 27948 3488 28908 3516
rect 27948 3476 27954 3488
rect 28902 3476 28908 3488
rect 28960 3476 28966 3528
rect 29086 3476 29092 3528
rect 29144 3516 29150 3528
rect 30282 3516 30288 3528
rect 29144 3488 30288 3516
rect 29144 3476 29150 3488
rect 30282 3476 30288 3488
rect 30340 3476 30346 3528
rect 33870 3476 33876 3528
rect 33928 3516 33934 3528
rect 114554 3516 114560 3528
rect 33928 3488 114560 3516
rect 33928 3476 33934 3488
rect 114554 3476 114560 3488
rect 114612 3476 114618 3528
rect 120626 3476 120632 3528
rect 120684 3516 120690 3528
rect 256694 3516 256700 3528
rect 120684 3488 256700 3516
rect 120684 3476 120690 3488
rect 256694 3476 256700 3488
rect 256752 3476 256758 3528
rect 30190 3408 30196 3460
rect 30248 3448 30254 3460
rect 35897 3451 35955 3457
rect 35897 3448 35909 3451
rect 30248 3420 35909 3448
rect 30248 3408 30254 3420
rect 35897 3417 35909 3420
rect 35943 3417 35955 3451
rect 35897 3411 35955 3417
rect 36170 3408 36176 3460
rect 36228 3448 36234 3460
rect 118694 3448 118700 3460
rect 36228 3420 118700 3448
rect 36228 3408 36234 3420
rect 118694 3408 118700 3420
rect 118752 3408 118758 3460
rect 124214 3408 124220 3460
rect 124272 3448 124278 3460
rect 262214 3448 262220 3460
rect 124272 3420 262220 3448
rect 124272 3408 124278 3420
rect 262214 3408 262220 3420
rect 262272 3408 262278 3460
rect 12434 3340 12440 3392
rect 12492 3380 12498 3392
rect 55217 3383 55275 3389
rect 55217 3380 55229 3383
rect 12492 3352 55229 3380
rect 12492 3340 12498 3352
rect 55217 3349 55229 3352
rect 55263 3349 55275 3383
rect 55217 3343 55275 3349
rect 58529 3383 58587 3389
rect 58529 3349 58541 3383
rect 58575 3380 58587 3383
rect 63678 3380 63684 3392
rect 58575 3352 63684 3380
rect 58575 3349 58587 3352
rect 58529 3343 58587 3349
rect 63678 3340 63684 3352
rect 63736 3340 63742 3392
rect 64785 3383 64843 3389
rect 64785 3349 64797 3383
rect 64831 3380 64843 3383
rect 64831 3352 76972 3380
rect 64831 3349 64843 3352
rect 64785 3343 64843 3349
rect 10042 3272 10048 3324
rect 10100 3312 10106 3324
rect 69661 3315 69719 3321
rect 69661 3312 69673 3315
rect 10100 3284 69673 3312
rect 10100 3272 10106 3284
rect 69661 3281 69673 3284
rect 69707 3281 69719 3315
rect 69661 3275 69719 3281
rect 71866 3272 71872 3324
rect 71924 3312 71930 3324
rect 72970 3312 72976 3324
rect 71924 3284 72976 3312
rect 71924 3272 71930 3284
rect 72970 3272 72976 3284
rect 73028 3272 73034 3324
rect 74534 3312 74540 3324
rect 73080 3284 74540 3312
rect 8846 3204 8852 3256
rect 8904 3244 8910 3256
rect 73080 3244 73108 3284
rect 74534 3272 74540 3284
rect 74592 3272 74598 3324
rect 76944 3312 76972 3352
rect 79042 3340 79048 3392
rect 79100 3380 79106 3392
rect 79962 3380 79968 3392
rect 79100 3352 79968 3380
rect 79100 3340 79106 3352
rect 79962 3340 79968 3352
rect 80020 3340 80026 3392
rect 80057 3383 80115 3389
rect 80057 3349 80069 3383
rect 80103 3380 80115 3383
rect 84194 3380 84200 3392
rect 80103 3352 84200 3380
rect 80103 3349 80115 3352
rect 80057 3343 80115 3349
rect 84194 3340 84200 3352
rect 84252 3340 84258 3392
rect 89714 3340 89720 3392
rect 89772 3380 89778 3392
rect 90910 3380 90916 3392
rect 89772 3352 90916 3380
rect 89772 3340 89778 3352
rect 90910 3340 90916 3352
rect 90968 3340 90974 3392
rect 204254 3380 204260 3392
rect 91112 3352 204260 3380
rect 80146 3312 80152 3324
rect 76944 3284 80152 3312
rect 80146 3272 80152 3284
rect 80204 3272 80210 3324
rect 88518 3272 88524 3324
rect 88576 3312 88582 3324
rect 91112 3312 91140 3352
rect 204254 3340 204260 3352
rect 204312 3340 204318 3392
rect 200114 3312 200120 3324
rect 88576 3284 91140 3312
rect 91204 3284 200120 3312
rect 88576 3272 88582 3284
rect 8904 3216 73108 3244
rect 8904 3204 8910 3216
rect 86126 3204 86132 3256
rect 86184 3244 86190 3256
rect 91204 3244 91232 3284
rect 200114 3272 200120 3284
rect 200172 3272 200178 3324
rect 86184 3216 91232 3244
rect 91281 3247 91339 3253
rect 86184 3204 86190 3216
rect 91281 3213 91293 3247
rect 91327 3244 91339 3247
rect 198734 3244 198740 3256
rect 91327 3216 198740 3244
rect 91327 3213 91339 3216
rect 91281 3207 91339 3213
rect 198734 3204 198740 3216
rect 198792 3204 198798 3256
rect 1670 3136 1676 3188
rect 1728 3176 1734 3188
rect 6825 3179 6883 3185
rect 6825 3176 6837 3179
rect 1728 3148 6837 3176
rect 1728 3136 1734 3148
rect 6825 3145 6837 3148
rect 6871 3145 6883 3179
rect 6825 3139 6883 3145
rect 7650 3136 7656 3188
rect 7708 3176 7714 3188
rect 69661 3179 69719 3185
rect 7708 3148 68416 3176
rect 7708 3136 7714 3148
rect 6454 3068 6460 3120
rect 6512 3108 6518 3120
rect 68281 3111 68339 3117
rect 68281 3108 68293 3111
rect 6512 3080 68293 3108
rect 6512 3068 6518 3080
rect 68281 3077 68293 3080
rect 68327 3077 68339 3111
rect 68281 3071 68339 3077
rect 4062 3000 4068 3052
rect 4120 3040 4126 3052
rect 66346 3040 66352 3052
rect 4120 3012 66352 3040
rect 4120 3000 4126 3012
rect 66346 3000 66352 3012
rect 66404 3000 66410 3052
rect 68388 3040 68416 3148
rect 69661 3145 69673 3179
rect 69707 3176 69719 3179
rect 76006 3176 76012 3188
rect 69707 3148 76012 3176
rect 69707 3145 69719 3148
rect 69661 3139 69719 3145
rect 76006 3136 76012 3148
rect 76064 3136 76070 3188
rect 77846 3136 77852 3188
rect 77904 3176 77910 3188
rect 186314 3176 186320 3188
rect 77904 3148 186320 3176
rect 77904 3136 77910 3148
rect 186314 3136 186320 3148
rect 186372 3136 186378 3188
rect 68465 3111 68523 3117
rect 68465 3077 68477 3111
rect 68511 3108 68523 3111
rect 70394 3108 70400 3120
rect 68511 3080 70400 3108
rect 68511 3077 68523 3080
rect 68465 3071 68523 3077
rect 70394 3068 70400 3080
rect 70452 3068 70458 3120
rect 71958 3108 71964 3120
rect 70504 3080 71964 3108
rect 70504 3040 70532 3080
rect 71958 3068 71964 3080
rect 72016 3068 72022 3120
rect 75454 3068 75460 3120
rect 75512 3108 75518 3120
rect 183554 3108 183560 3120
rect 75512 3080 183560 3108
rect 75512 3068 75518 3080
rect 183554 3068 183560 3080
rect 183612 3068 183618 3120
rect 68388 3012 70532 3040
rect 70670 3000 70676 3052
rect 70728 3040 70734 3052
rect 175274 3040 175280 3052
rect 70728 3012 175280 3040
rect 70728 3000 70734 3012
rect 175274 3000 175280 3012
rect 175332 3000 175338 3052
rect 566 2932 572 2984
rect 624 2972 630 2984
rect 61378 2972 61384 2984
rect 624 2944 61384 2972
rect 624 2932 630 2944
rect 61378 2932 61384 2944
rect 61436 2932 61442 2984
rect 63773 2975 63831 2981
rect 63773 2941 63785 2975
rect 63819 2972 63831 2975
rect 64785 2975 64843 2981
rect 64785 2972 64797 2975
rect 63819 2944 64797 2972
rect 63819 2941 63831 2944
rect 63773 2935 63831 2941
rect 64785 2941 64797 2944
rect 64831 2941 64843 2975
rect 64785 2935 64843 2941
rect 68278 2932 68284 2984
rect 68336 2972 68342 2984
rect 171134 2972 171140 2984
rect 68336 2944 171140 2972
rect 68336 2932 68342 2944
rect 171134 2932 171140 2944
rect 171192 2932 171198 2984
rect 6825 2907 6883 2913
rect 6825 2873 6837 2907
rect 6871 2904 6883 2907
rect 6871 2876 58940 2904
rect 6871 2873 6883 2876
rect 6825 2867 6883 2873
rect 2866 2796 2872 2848
rect 2924 2836 2930 2848
rect 58529 2839 58587 2845
rect 58529 2836 58541 2839
rect 2924 2808 58541 2836
rect 2924 2796 2930 2808
rect 58529 2805 58541 2808
rect 58575 2805 58587 2839
rect 58912 2836 58940 2876
rect 61194 2864 61200 2916
rect 61252 2904 61258 2916
rect 160094 2904 160100 2916
rect 61252 2876 160100 2904
rect 61252 2864 61258 2876
rect 160094 2864 160100 2876
rect 160152 2864 160158 2916
rect 62206 2836 62212 2848
rect 58912 2808 62212 2836
rect 58529 2799 58587 2805
rect 62206 2796 62212 2808
rect 62264 2796 62270 2848
rect 63497 2839 63555 2845
rect 63497 2836 63509 2839
rect 62316 2808 63509 2836
rect 55217 2703 55275 2709
rect 55217 2669 55229 2703
rect 55263 2700 55275 2703
rect 62316 2700 62344 2808
rect 63497 2805 63509 2808
rect 63543 2805 63555 2839
rect 63497 2799 63555 2805
rect 63586 2796 63592 2848
rect 63644 2836 63650 2848
rect 162854 2836 162860 2848
rect 63644 2808 162860 2836
rect 63644 2796 63650 2808
rect 162854 2796 162860 2808
rect 162912 2796 162918 2848
rect 55263 2672 62344 2700
rect 55263 2669 55275 2672
rect 55217 2663 55275 2669
rect 5258 552 5264 604
rect 5316 592 5322 604
rect 5442 592 5448 604
rect 5316 564 5448 592
rect 5316 552 5322 564
rect 5442 552 5448 564
rect 5500 552 5506 604
rect 74258 552 74264 604
rect 74316 592 74322 604
rect 74442 592 74448 604
rect 74316 564 74448 592
rect 74316 552 74322 564
rect 74442 552 74448 564
rect 74500 552 74506 604
<< via1 >>
rect 263600 653352 263652 653404
rect 378140 653352 378192 653404
rect 383568 653352 383620 653404
rect 508412 653352 508464 653404
rect 378140 652876 378192 652928
rect 383568 652876 383620 652928
rect 135168 652740 135220 652792
rect 139400 652808 139452 652860
rect 508412 652808 508464 652860
rect 513380 652808 513432 652860
rect 258540 652740 258592 652792
rect 518900 652740 518952 652792
rect 266636 650428 266688 650480
rect 407764 650496 407816 650548
rect 387156 650428 387208 650480
rect 137652 650224 137704 650276
rect 516416 650428 516468 650480
rect 389180 650156 389232 650208
rect 291844 645872 291896 645924
rect 307392 645872 307444 645924
rect 290464 644444 290516 644496
rect 307116 644444 307168 644496
rect 287704 643084 287756 643136
rect 307116 643084 307168 643136
rect 286324 641724 286376 641776
rect 307668 641724 307720 641776
rect 284944 640296 284996 640348
rect 307668 640296 307720 640348
rect 291936 637576 291988 637628
rect 306840 637576 306892 637628
rect 270408 580252 270460 580304
rect 279148 580252 279200 580304
rect 302884 579640 302936 579692
rect 307668 579640 307720 579692
rect 77392 558832 77444 558884
rect 86316 558832 86368 558884
rect 86684 558832 86736 558884
rect 93768 558832 93820 558884
rect 137284 558832 137336 558884
rect 194416 558832 194468 558884
rect 313832 558900 313884 558952
rect 413928 558900 413980 558952
rect 347688 558832 347740 558884
rect 356060 558832 356112 558884
rect 468024 558832 468076 558884
rect 476580 558832 476632 558884
rect 66168 558764 66220 558816
rect 200212 558764 200264 558816
rect 215300 558764 215352 558816
rect 224500 558764 224552 558816
rect 286416 558764 286468 558816
rect 453672 558764 453724 558816
rect 75000 558696 75052 558748
rect 84200 558696 84252 558748
rect 93308 558696 93360 558748
rect 102784 558696 102836 558748
rect 106280 558696 106332 558748
rect 107292 558696 107344 558748
rect 141424 558696 141476 558748
rect 218796 558696 218848 558748
rect 227996 558696 228048 558748
rect 237380 558696 237432 558748
rect 286508 558696 286560 558748
rect 454776 558696 454828 558748
rect 78496 558628 78548 558680
rect 87880 558628 87932 558680
rect 97172 558628 97224 558680
rect 99472 558628 99524 558680
rect 102048 558628 102100 558680
rect 140044 558628 140096 558680
rect 222200 558628 222252 558680
rect 231860 558628 231912 558680
rect 326344 558628 326396 558680
rect 335452 558628 335504 558680
rect 344284 558628 344336 558680
rect 353300 558628 353352 558680
rect 75920 558560 75972 558612
rect 85396 558560 85448 558612
rect 86684 558560 86736 558612
rect 95700 558560 95752 558612
rect 79416 558492 79468 558544
rect 88892 558492 88944 558544
rect 98368 558492 98420 558544
rect 104164 558560 104216 558612
rect 108488 558560 108540 558612
rect 148324 558560 148376 558612
rect 217508 558560 217560 558612
rect 225880 558560 225932 558612
rect 234620 558560 234672 558612
rect 336096 558560 336148 558612
rect 336648 558560 336700 558612
rect 346032 558560 346084 558612
rect 354680 558560 354732 558612
rect 457444 558764 457496 558816
rect 466552 558764 466604 558816
rect 475476 558764 475528 558816
rect 458824 558696 458876 558748
rect 468024 558696 468076 558748
rect 468116 558696 468168 558748
rect 468760 558696 468812 558748
rect 477592 558696 477644 558748
rect 456064 558628 456116 558680
rect 465264 558628 465316 558680
rect 474832 558628 474884 558680
rect 484400 558628 484452 558680
rect 463056 558560 463108 558612
rect 472164 558560 472216 558612
rect 481640 558560 481692 558612
rect 80796 558424 80848 558476
rect 89812 558424 89864 558476
rect 94780 558424 94832 558476
rect 100024 558492 100076 558544
rect 104808 558492 104860 558544
rect 144184 558492 144236 558544
rect 208492 558492 208544 558544
rect 217600 558492 217652 558544
rect 227168 558492 227220 558544
rect 236000 558492 236052 558544
rect 330484 558492 330536 558544
rect 339868 558492 339920 558544
rect 349712 558492 349764 558544
rect 358176 558492 358228 558544
rect 453304 558492 453356 558544
rect 461676 558492 461728 558544
rect 471336 558492 471388 558544
rect 480352 558492 480404 558544
rect 140136 558424 140188 558476
rect 213184 558424 213236 558476
rect 222200 558424 222252 558476
rect 329288 558424 329340 558476
rect 339040 558424 339092 558476
rect 348240 558424 348292 558476
rect 357440 558424 357492 558476
rect 413928 558424 413980 558476
rect 443092 558424 443144 558476
rect 454776 558424 454828 558476
rect 464252 558424 464304 558476
rect 473452 558424 473504 558476
rect 483020 558424 483072 558476
rect 73712 558356 73764 558408
rect 82912 558356 82964 558408
rect 92480 558356 92532 558408
rect 93124 558356 93176 558408
rect 97816 558356 97868 558408
rect 138664 558356 138716 558408
rect 210608 558356 210660 558408
rect 220084 558356 220136 558408
rect 229468 558356 229520 558408
rect 81440 558288 81492 558340
rect 81992 558288 82044 558340
rect 91100 558288 91152 558340
rect 92204 558288 92256 558340
rect 137468 558288 137520 558340
rect 211160 558288 211212 558340
rect 211804 558288 211856 558340
rect 221096 558288 221148 558340
rect 230480 558288 230532 558340
rect 74264 558220 74316 558272
rect 137376 558220 137428 558272
rect 206928 558220 206980 558272
rect 215300 558220 215352 558272
rect 224500 558220 224552 558272
rect 233240 558220 233292 558272
rect 334072 558356 334124 558408
rect 335268 558356 335320 558408
rect 337568 558356 337620 558408
rect 347688 558356 347740 558408
rect 352564 558356 352616 558408
rect 476212 558356 476264 558408
rect 476580 558356 476632 558408
rect 485780 558356 485832 558408
rect 238760 558220 238812 558272
rect 72516 558152 72568 558204
rect 81440 558152 81492 558204
rect 83832 558152 83884 558204
rect 149704 558152 149756 558204
rect 203800 558152 203852 558204
rect 213184 558152 213236 558204
rect 76840 558084 76892 558136
rect 145564 558084 145616 558136
rect 215208 558084 215260 558136
rect 285128 558084 285180 558136
rect 328460 558084 328512 558136
rect 81256 558016 81308 558068
rect 152556 558016 152608 558068
rect 231860 558016 231912 558068
rect 312544 558016 312596 558068
rect 322940 558016 322992 558068
rect 323584 558016 323636 558068
rect 333152 558288 333204 558340
rect 342536 558288 342588 558340
rect 348424 558288 348476 558340
rect 352656 558288 352708 558340
rect 477500 558288 477552 558340
rect 477592 558288 477644 558340
rect 487160 558288 487212 558340
rect 79324 557948 79376 558000
rect 152464 557948 152516 558000
rect 309784 557948 309836 558000
rect 321560 557948 321612 558000
rect 322204 557948 322256 558000
rect 331772 558220 331824 558272
rect 341248 558220 341300 558272
rect 350540 558220 350592 558272
rect 353944 558220 353996 558272
rect 478880 558220 478932 558272
rect 478972 558220 479024 558272
rect 488540 558220 488592 558272
rect 335268 558152 335320 558204
rect 343640 558152 343692 558204
rect 352012 558152 352064 558204
rect 354036 558152 354088 558204
rect 480352 558152 480404 558204
rect 356704 558084 356756 558136
rect 483020 558084 483072 558136
rect 355324 558016 355376 558068
rect 481640 558016 481692 558068
rect 356796 557948 356848 558000
rect 484400 557948 484452 558000
rect 97172 557880 97224 557932
rect 105544 557880 105596 557932
rect 129648 557880 129700 557932
rect 223580 557880 223632 557932
rect 286600 557880 286652 557932
rect 329840 557880 329892 557932
rect 355416 557880 355468 557932
rect 483020 557880 483072 557932
rect 89168 557812 89220 557864
rect 93124 557744 93176 557796
rect 100852 557744 100904 557796
rect 125508 557812 125560 557864
rect 208492 557812 208544 557864
rect 324964 557812 325016 557864
rect 358084 557812 358136 557864
rect 485780 557812 485832 557864
rect 121368 557744 121420 557796
rect 206928 557744 206980 557796
rect 209044 557744 209096 557796
rect 218796 557744 218848 557796
rect 287796 557744 287848 557796
rect 331220 557744 331272 557796
rect 358176 557744 358228 557796
rect 487160 557744 487212 557796
rect 85396 557676 85448 557728
rect 94780 557676 94832 557728
rect 98368 557676 98420 557728
rect 108304 557676 108356 557728
rect 117228 557676 117280 557728
rect 203800 557676 203852 557728
rect 204904 557676 204956 557728
rect 214012 557676 214064 557728
rect 215208 557676 215260 557728
rect 285036 557676 285088 557728
rect 449900 557676 449952 557728
rect 460388 557676 460440 557728
rect 468116 557676 468168 557728
rect 474832 557676 474884 557728
rect 483020 557676 483072 557728
rect 91100 557608 91152 557660
rect 100024 557608 100076 557660
rect 100392 557608 100444 557660
rect 108488 557608 108540 557660
rect 202144 557608 202196 557660
rect 211160 557608 211212 557660
rect 315304 557608 315356 557660
rect 324320 557608 324372 557660
rect 327724 557608 327776 557660
rect 336096 557608 336148 557660
rect 460204 557608 460256 557660
rect 460848 557608 460900 557660
rect 470048 557608 470100 557660
rect 478972 557608 479024 557660
rect 67456 557540 67508 557592
rect 201500 557540 201552 557592
rect 207664 557540 207716 557592
rect 217508 557540 217560 557592
rect 308404 557540 308456 557592
rect 316316 557540 316368 557592
rect 329104 557540 329156 557592
rect 337568 557540 337620 557592
rect 464344 557540 464396 557592
rect 488540 557540 488592 557592
rect 131764 556860 131816 556912
rect 96528 545028 96580 545080
rect 189632 545028 189684 545080
rect 94136 544960 94188 545012
rect 188436 544960 188488 545012
rect 102048 544892 102100 544944
rect 197912 544892 197964 544944
rect 92112 544824 92164 544876
rect 188528 544824 188580 544876
rect 89996 544756 90048 544808
rect 188620 544756 188672 544808
rect 106188 544688 106240 544740
rect 206192 544688 206244 544740
rect 87972 544620 88024 544672
rect 188712 544620 188764 544672
rect 110328 544552 110380 544604
rect 212448 544552 212500 544604
rect 85856 544484 85908 544536
rect 188804 544484 188856 544536
rect 83832 544416 83884 544468
rect 188896 544416 188948 544468
rect 81716 544348 81768 544400
rect 195980 544348 196032 544400
rect 86776 544280 86828 544332
rect 173072 544280 173124 544332
rect 88248 544212 88300 544264
rect 175096 544212 175148 544264
rect 85488 544144 85540 544196
rect 168840 544144 168892 544196
rect 86868 544076 86920 544128
rect 170956 544076 171008 544128
rect 82728 544008 82780 544060
rect 164700 544008 164752 544060
rect 73068 543940 73120 543992
rect 148140 543940 148192 543992
rect 57888 543872 57940 543924
rect 112812 543872 112864 543924
rect 57796 543804 57848 543856
rect 110788 543804 110840 543856
rect 220728 543736 220780 543788
rect 71688 543668 71740 543720
rect 75460 543668 75512 543720
rect 75828 543668 75880 543720
rect 145564 543668 145616 543720
rect 152556 543668 152608 543720
rect 162676 543668 162728 543720
rect 205548 543668 205600 543720
rect 218704 543668 218756 543720
rect 220544 543668 220596 543720
rect 229008 543668 229060 543720
rect 260196 543668 260248 543720
rect 70308 543600 70360 543652
rect 73436 543600 73488 543652
rect 78588 543600 78640 543652
rect 156420 543600 156472 543652
rect 206928 543600 206980 543652
rect 220728 543600 220780 543652
rect 227628 543600 227680 543652
rect 258080 543600 258132 543652
rect 61016 543532 61068 543584
rect 62028 543532 62080 543584
rect 65156 543532 65208 543584
rect 66168 543532 66220 543584
rect 70216 543532 70268 543584
rect 71320 543532 71372 543584
rect 79876 543532 79928 543584
rect 152464 543532 152516 543584
rect 158536 543532 158588 543584
rect 208308 543532 208360 543584
rect 222844 543532 222896 543584
rect 230388 543532 230440 543584
rect 262220 543532 262272 543584
rect 57428 543464 57480 543516
rect 102508 543464 102560 543516
rect 127348 543464 127400 543516
rect 209044 543464 209096 543516
rect 209688 543464 209740 543516
rect 224868 543464 224920 543516
rect 231768 543464 231820 543516
rect 264336 543464 264388 543516
rect 57520 543396 57572 543448
rect 104532 543396 104584 543448
rect 123208 543396 123260 543448
rect 207664 543396 207716 543448
rect 211068 543396 211120 543448
rect 226984 543396 227036 543448
rect 233148 543396 233200 543448
rect 266452 543396 266504 543448
rect 57612 543328 57664 543380
rect 106648 543328 106700 543380
rect 119068 543328 119120 543380
rect 204904 543328 204956 543380
rect 212356 543328 212408 543380
rect 231124 543328 231176 543380
rect 233056 543328 233108 543380
rect 268476 543328 268528 543380
rect 91008 543260 91060 543312
rect 179236 543260 179288 543312
rect 215208 543260 215260 543312
rect 235264 543260 235316 543312
rect 235908 543260 235960 543312
rect 272616 543260 272668 543312
rect 57704 543192 57756 543244
rect 108672 543192 108724 543244
rect 114928 543192 114980 543244
rect 202144 543192 202196 543244
rect 216496 543192 216548 543244
rect 93676 543124 93728 543176
rect 183376 543124 183428 543176
rect 204168 543124 204220 543176
rect 216588 543124 216640 543176
rect 229100 543192 229152 543244
rect 234528 543192 234580 543244
rect 270592 543192 270644 543244
rect 237380 543124 237432 543176
rect 238668 543124 238720 543176
rect 276756 543124 276808 543176
rect 57244 543056 57296 543108
rect 79692 543056 79744 543108
rect 95056 543056 95108 543108
rect 187516 543056 187568 543108
rect 213828 543056 213880 543108
rect 233240 543056 233292 543108
rect 237288 543056 237340 543108
rect 274732 543056 274784 543108
rect 67548 542988 67600 543040
rect 98368 542988 98420 543040
rect 99288 542988 99340 543040
rect 193772 542988 193824 543040
rect 202788 542988 202840 543040
rect 214564 542988 214616 543040
rect 217968 542988 218020 543040
rect 239404 542988 239456 543040
rect 240048 542988 240100 543040
rect 278872 542988 278924 543040
rect 57336 542920 57388 542972
rect 100392 542920 100444 542972
rect 108304 542920 108356 542972
rect 144000 542920 144052 542972
rect 144184 542920 144236 542972
rect 204168 542920 204220 542972
rect 210976 542920 211028 542972
rect 226156 542920 226208 542972
rect 256056 542920 256108 542972
rect 105544 542852 105596 542904
rect 139860 542852 139912 542904
rect 140136 542852 140188 542904
rect 195888 542852 195940 542904
rect 226248 542852 226300 542904
rect 253940 542852 253992 542904
rect 102784 542784 102836 542836
rect 135720 542784 135772 542836
rect 137284 542784 137336 542836
rect 104164 542716 104216 542768
rect 137744 542716 137796 542768
rect 138664 542784 138716 542836
rect 191748 542784 191800 542836
rect 223488 542784 223540 542836
rect 249800 542784 249852 542836
rect 185492 542716 185544 542768
rect 224684 542716 224736 542768
rect 251916 542716 251968 542768
rect 100024 542648 100076 542700
rect 131488 542648 131540 542700
rect 131764 542648 131816 542700
rect 177212 542648 177264 542700
rect 220544 542648 220596 542700
rect 245660 542648 245712 542700
rect 101404 542580 101456 542632
rect 133604 542580 133656 542632
rect 137468 542580 137520 542632
rect 181352 542580 181404 542632
rect 222108 542580 222160 542632
rect 247776 542580 247828 542632
rect 108488 542512 108540 542564
rect 146024 542512 146076 542564
rect 106924 542444 106976 542496
rect 141884 542444 141936 542496
rect 152280 542512 152332 542564
rect 154396 542512 154448 542564
rect 149704 542444 149756 542496
rect 166816 542512 166868 542564
rect 217876 542512 217928 542564
rect 241520 542512 241572 542564
rect 219348 542444 219400 542496
rect 243544 542444 243596 542496
rect 137376 542376 137428 542428
rect 150164 542376 150216 542428
rect 160560 542376 160612 542428
rect 282276 538296 282328 538348
rect 367100 538296 367152 538348
rect 282828 538228 282880 538280
rect 368480 538228 368532 538280
rect 282828 536800 282880 536852
rect 369860 536800 369912 536852
rect 282828 535440 282880 535492
rect 371240 535440 371292 535492
rect 281724 534148 281776 534200
rect 372620 534148 372672 534200
rect 282092 534080 282144 534132
rect 374000 534080 374052 534132
rect 282092 532720 282144 532772
rect 375380 532720 375432 532772
rect 282276 531360 282328 531412
rect 375472 531360 375524 531412
rect 282828 531292 282880 531344
rect 376760 531292 376812 531344
rect 282828 529932 282880 529984
rect 378232 529932 378284 529984
rect 282828 528572 282880 528624
rect 379612 528572 379664 528624
rect 282828 527212 282880 527264
rect 376024 527212 376076 527264
rect 282276 527144 282328 527196
rect 380992 527144 381044 527196
rect 281908 525784 281960 525836
rect 374644 525784 374696 525836
rect 282828 524424 282880 524476
rect 371884 524424 371936 524476
rect 282828 523064 282880 523116
rect 354128 523064 354180 523116
rect 282368 522996 282420 523048
rect 367744 522996 367796 523048
rect 282828 521636 282880 521688
rect 387892 521636 387944 521688
rect 282828 520276 282880 520328
rect 390652 520276 390704 520328
rect 281724 519052 281776 519104
rect 283748 519052 283800 519104
rect 282092 517488 282144 517540
rect 392032 517488 392084 517540
rect 282276 516196 282328 516248
rect 387064 516196 387116 516248
rect 282828 516128 282880 516180
rect 419540 516128 419592 516180
rect 282828 514768 282880 514820
rect 385684 514768 385736 514820
rect 282276 513340 282328 513392
rect 419632 513340 419684 513392
rect 282736 512048 282788 512100
rect 385776 512048 385828 512100
rect 282828 511980 282880 512032
rect 419724 511980 419776 512032
rect 281724 510620 281776 510672
rect 384304 510620 384356 510672
rect 282276 509260 282328 509312
rect 419816 509260 419868 509312
rect 282552 507900 282604 507952
rect 382924 507900 382976 507952
rect 282828 507832 282880 507884
rect 419908 507832 419960 507884
rect 282092 506472 282144 506524
rect 383016 506472 383068 506524
rect 282828 505180 282880 505232
rect 383108 505180 383160 505232
rect 282736 505112 282788 505164
rect 420000 505112 420052 505164
rect 282828 503684 282880 503736
rect 420092 503684 420144 503736
rect 282828 502324 282880 502376
rect 383200 502324 383252 502376
rect 282828 501032 282880 501084
rect 378784 501032 378836 501084
rect 282276 500964 282328 501016
rect 410524 500964 410576 501016
rect 282828 498176 282880 498228
rect 283932 498176 283984 498228
rect 282828 496816 282880 496868
rect 416320 496816 416372 496868
rect 281908 495456 281960 495508
rect 498844 495456 498896 495508
rect 282828 494028 282880 494080
rect 496084 494028 496136 494080
rect 282828 492736 282880 492788
rect 491944 492736 491996 492788
rect 282368 492668 282420 492720
rect 493324 492668 493376 492720
rect 282828 491308 282880 491360
rect 489184 491308 489236 491360
rect 282828 489948 282880 490000
rect 483664 489948 483716 490000
rect 282276 489880 282328 489932
rect 485044 489880 485096 489932
rect 282276 488520 282328 488572
rect 482284 488520 482336 488572
rect 282828 487160 282880 487212
rect 480904 487160 480956 487212
rect 282828 485868 282880 485920
rect 465724 485868 465776 485920
rect 282276 485800 282328 485852
rect 467104 485800 467156 485852
rect 281724 484372 281776 484424
rect 449164 484372 449216 484424
rect 282276 483012 282328 483064
rect 446404 483012 446456 483064
rect 282828 481720 282880 481772
rect 442264 481720 442316 481772
rect 282552 481652 282604 481704
rect 445024 481652 445076 481704
rect 282092 480224 282144 480276
rect 435364 480224 435416 480276
rect 282828 478932 282880 478984
rect 431224 478932 431276 478984
rect 282736 478864 282788 478916
rect 433984 478864 434036 478916
rect 282828 477504 282880 477556
rect 429844 477504 429896 477556
rect 282092 476076 282144 476128
rect 428464 476076 428516 476128
rect 282828 474784 282880 474836
rect 424324 474784 424376 474836
rect 282276 474716 282328 474768
rect 427084 474716 427136 474768
rect 281724 473356 281776 473408
rect 416044 473356 416096 473408
rect 282092 471996 282144 472048
rect 477592 471996 477644 472048
rect 282828 470636 282880 470688
rect 409144 470636 409196 470688
rect 282736 470568 282788 470620
rect 411904 470568 411956 470620
rect 281908 469208 281960 469260
rect 474832 469208 474884 469260
rect 282828 467848 282880 467900
rect 473452 467848 473504 467900
rect 282736 466488 282788 466540
rect 406384 466488 406436 466540
rect 282828 466420 282880 466472
rect 470692 466420 470744 466472
rect 282828 465060 282880 465112
rect 447784 465060 447836 465112
rect 282736 463768 282788 463820
rect 417424 463768 417476 463820
rect 282828 463700 282880 463752
rect 526352 463700 526404 463752
rect 282828 462340 282880 462392
rect 283656 462340 283708 462392
rect 282828 460912 282880 460964
rect 368572 460912 368624 460964
rect 282736 459620 282788 459672
rect 283840 459620 283892 459672
rect 282828 459552 282880 459604
rect 369952 459552 370004 459604
rect 281724 458192 281776 458244
rect 284024 458192 284076 458244
rect 282092 456764 282144 456816
rect 284116 456764 284168 456816
rect 281632 455472 281684 455524
rect 284208 455472 284260 455524
rect 282828 455404 282880 455456
rect 375564 455404 375616 455456
rect 282184 440376 282236 440428
rect 384396 440376 384448 440428
rect 281448 440240 281500 440292
rect 387156 440240 387208 440292
rect 282184 438880 282236 438932
rect 381544 438880 381596 438932
rect 282184 436568 282236 436620
rect 282184 436160 282236 436212
rect 377404 436160 377456 436212
rect 380164 436092 380216 436144
rect 282184 434732 282236 434784
rect 374736 434732 374788 434784
rect 282184 433304 282236 433356
rect 373264 433304 373316 433356
rect 282276 431536 282328 431588
rect 282276 430652 282328 430704
rect 388444 430652 388496 430704
rect 282276 430516 282328 430568
rect 464344 430516 464396 430568
rect 281448 429156 281500 429208
rect 416780 429156 416832 429208
rect 282276 429088 282328 429140
rect 358176 429088 358228 429140
rect 282276 427728 282328 427780
rect 358084 427728 358136 427780
rect 356796 427660 356848 427712
rect 282276 427184 282328 427236
rect 282276 426368 282328 426420
rect 356704 426368 356756 426420
rect 282276 425008 282328 425060
rect 355416 425008 355468 425060
rect 282276 423580 282328 423632
rect 355324 423580 355376 423632
rect 354036 423512 354088 423564
rect 282276 423240 282328 423292
rect 282276 422220 282328 422272
rect 353944 422220 353996 422272
rect 281632 421379 281684 421388
rect 281632 421345 281641 421379
rect 281641 421345 281675 421379
rect 281675 421345 281684 421379
rect 281632 421336 281684 421345
rect 281632 421200 281684 421252
rect 282460 421200 282512 421252
rect 282460 420996 282512 421048
rect 282828 420996 282880 421048
rect 282828 420860 282880 420912
rect 352656 420860 352708 420912
rect 282552 419432 282604 419484
rect 476120 419432 476172 419484
rect 282828 419364 282880 419416
rect 352564 419364 352616 419416
rect 282828 418072 282880 418124
rect 474740 418072 474792 418124
rect 282276 417732 282328 417784
rect 282552 417732 282604 417784
rect 282276 417596 282328 417648
rect 282828 416712 282880 416764
rect 473360 416712 473412 416764
rect 284576 416372 284628 416424
rect 453304 416372 453356 416424
rect 286232 416304 286284 416356
rect 455420 416304 455472 416356
rect 286140 416236 286192 416288
rect 456800 416236 456852 416288
rect 283288 416168 283340 416220
rect 458180 416168 458232 416220
rect 283196 416100 283248 416152
rect 459560 416100 459612 416152
rect 283104 416032 283156 416084
rect 461032 416032 461084 416084
rect 282276 415420 282328 415472
rect 282920 415420 282972 415472
rect 282828 415352 282880 415404
rect 471980 415352 472032 415404
rect 282276 415284 282328 415336
rect 470600 415284 470652 415336
rect 285404 415216 285456 415268
rect 438584 415216 438636 415268
rect 285312 415148 285364 415200
rect 438676 415148 438728 415200
rect 284760 415080 284812 415132
rect 438124 415080 438176 415132
rect 284852 415012 284904 415064
rect 438308 415012 438360 415064
rect 284668 414944 284720 414996
rect 438216 414944 438268 414996
rect 285220 414876 285272 414928
rect 445760 414876 445812 414928
rect 292028 414808 292080 414860
rect 452752 414808 452804 414860
rect 283012 414740 283064 414792
rect 467932 414740 467984 414792
rect 282920 414672 282972 414724
rect 469220 414672 469272 414724
rect 285496 414604 285548 414656
rect 438492 414604 438544 414656
rect 285588 414536 285640 414588
rect 438400 414536 438452 414588
rect 337384 414468 337436 414520
rect 454040 414468 454092 414520
rect 284392 414400 284444 414452
rect 343732 414400 343784 414452
rect 284484 414332 284536 414384
rect 342260 414332 342312 414384
rect 383108 413992 383160 414044
rect 282184 413924 282236 413976
rect 402980 413924 403032 413976
rect 447784 413924 447836 413976
rect 469404 413924 469456 413976
rect 496084 413924 496136 413976
rect 505100 413924 505152 413976
rect 282276 413856 282328 413908
rect 283472 413856 283524 413908
rect 396080 413856 396132 413908
rect 409144 413856 409196 413908
rect 476120 413856 476172 413908
rect 489184 413856 489236 413908
rect 502524 413856 502576 413908
rect 281724 413788 281776 413840
rect 387156 413788 387208 413840
rect 391940 413788 391992 413840
rect 411904 413788 411956 413840
rect 477500 413788 477552 413840
rect 483664 413788 483716 413840
rect 499580 413788 499632 413840
rect 281908 413720 281960 413772
rect 389272 413720 389324 413772
rect 406384 413720 406436 413772
rect 471980 413720 472032 413772
rect 491944 413720 491996 413772
rect 503720 413720 503772 413772
rect 282000 413652 282052 413704
rect 389180 413652 389232 413704
rect 416044 413652 416096 413704
rect 478880 413652 478932 413704
rect 482284 413652 482336 413704
rect 498292 413652 498344 413704
rect 498844 413652 498896 413704
rect 506480 413652 506532 413704
rect 281816 413584 281868 413636
rect 282092 413516 282144 413568
rect 386420 413584 386472 413636
rect 388536 413584 388588 413636
rect 404360 413584 404412 413636
rect 413928 413584 413980 413636
rect 420184 413584 420236 413636
rect 424324 413584 424376 413636
rect 480444 413584 480496 413636
rect 480904 413584 480956 413636
rect 496820 413584 496872 413636
rect 381544 413516 381596 413568
rect 394700 413516 394752 413568
rect 431224 413516 431276 413568
rect 485780 413516 485832 413568
rect 282736 413448 282788 413500
rect 376024 413448 376076 413500
rect 382280 413448 382332 413500
rect 383200 413448 383252 413500
rect 401600 413448 401652 413500
rect 428464 413448 428516 413500
rect 483020 413448 483072 413500
rect 493324 413448 493376 413500
rect 503996 413448 504048 413500
rect 282644 413380 282696 413432
rect 397460 413380 397512 413432
rect 427084 413380 427136 413432
rect 481640 413380 481692 413432
rect 485044 413380 485096 413432
rect 501052 413380 501104 413432
rect 282368 413312 282420 413364
rect 382188 413312 382240 413364
rect 397552 413312 397604 413364
rect 429844 413312 429896 413364
rect 484400 413312 484452 413364
rect 282460 413244 282512 413296
rect 382372 413244 382424 413296
rect 383016 413244 383068 413296
rect 398840 413244 398892 413296
rect 435364 413244 435416 413296
rect 488540 413244 488592 413296
rect 282552 413176 282604 413228
rect 378784 413176 378836 413228
rect 384304 413176 384356 413228
rect 384396 413176 384448 413228
rect 393320 413176 393372 413228
rect 433984 413176 434036 413228
rect 487160 413176 487212 413228
rect 282736 413108 282788 413160
rect 281632 413040 281684 413092
rect 378140 413040 378192 413092
rect 383660 413108 383712 413160
rect 390560 413108 390612 413160
rect 417424 413108 417476 413160
rect 468116 413108 468168 413160
rect 379612 413040 379664 413092
rect 380164 413040 380216 413092
rect 385776 413040 385828 413092
rect 396080 413040 396132 413092
rect 442264 413040 442316 413092
rect 489920 413040 489972 413092
rect 282276 412972 282328 413024
rect 287060 412972 287112 413024
rect 296628 412972 296680 413024
rect 306380 412972 306432 413024
rect 315948 412972 316000 413024
rect 331128 412972 331180 413024
rect 335268 412972 335320 413024
rect 350448 412972 350500 413024
rect 354588 412972 354640 413024
rect 364340 412972 364392 413024
rect 376760 412972 376812 413024
rect 380900 412972 380952 413024
rect 387800 412972 387852 413024
rect 397460 412972 397512 413024
rect 445024 412972 445076 413024
rect 491300 412972 491352 413024
rect 284116 412904 284168 412956
rect 374000 412904 374052 412956
rect 284208 412836 284260 412888
rect 374184 412836 374236 412888
rect 374644 412836 374696 412888
rect 382280 412836 382332 412888
rect 382924 412904 382976 412956
rect 384304 412904 384356 412956
rect 403164 412904 403216 412956
rect 446404 412904 446456 412956
rect 491392 412904 491444 412956
rect 385040 412836 385092 412888
rect 385684 412836 385736 412888
rect 394700 412836 394752 412888
rect 449164 412836 449216 412888
rect 492680 412836 492732 412888
rect 284024 412768 284076 412820
rect 372620 412768 372672 412820
rect 373264 412768 373316 412820
rect 400220 412768 400272 412820
rect 410524 412768 410576 412820
rect 517520 412768 517572 412820
rect 283840 412700 283892 412752
rect 371240 412700 371292 412752
rect 371332 412700 371384 412752
rect 374736 412700 374788 412752
rect 377404 412700 377456 412752
rect 398840 412700 398892 412752
rect 467104 412700 467156 412752
rect 495716 412700 495768 412752
rect 283656 412632 283708 412684
rect 367100 412632 367152 412684
rect 367744 412632 367796 412684
rect 385040 412632 385092 412684
rect 283932 412564 283984 412616
rect 352104 412564 352156 412616
rect 400220 412632 400272 412684
rect 465724 412632 465776 412684
rect 494060 412632 494112 412684
rect 283748 412496 283800 412548
rect 352012 412496 352064 412548
rect 283840 412428 283892 412480
rect 353300 412428 353352 412480
rect 284024 412360 284076 412412
rect 354680 412360 354732 412412
rect 284116 412292 284168 412344
rect 356152 412292 356204 412344
rect 283472 412224 283524 412276
rect 357532 412224 357584 412276
rect 284208 412156 284260 412208
rect 358912 412156 358964 412208
rect 343088 412088 343140 412140
rect 467840 412088 467892 412140
rect 338028 412020 338080 412072
rect 463700 412020 463752 412072
rect 283380 411952 283432 412004
rect 452660 411952 452712 412004
rect 292580 411884 292632 411936
rect 465080 411884 465132 411936
rect 283656 411816 283708 411868
rect 350632 411816 350684 411868
rect 283564 411748 283616 411800
rect 349160 411748 349212 411800
rect 286968 411680 287020 411732
rect 347780 411680 347832 411732
rect 286876 411612 286928 411664
rect 346400 411612 346452 411664
rect 286692 411544 286744 411596
rect 345020 411544 345072 411596
rect 286784 411476 286836 411528
rect 343640 411476 343692 411528
rect 338764 411272 338816 411324
rect 405740 411272 405792 411324
rect 282736 411204 282788 411256
rect 466460 411204 466512 411256
rect 282828 411136 282880 411188
rect 343088 411136 343140 411188
rect 281632 411068 281684 411120
rect 438768 411068 438820 411120
rect 282000 411000 282052 411052
rect 451280 411000 451332 411052
rect 282184 410932 282236 410984
rect 456064 410932 456116 410984
rect 282276 410864 282328 410916
rect 457444 410864 457496 410916
rect 282644 410796 282696 410848
rect 458824 410796 458876 410848
rect 282552 410728 282604 410780
rect 460204 410728 460256 410780
rect 282460 410660 282512 410712
rect 460388 410660 460440 410712
rect 282368 410592 282420 410644
rect 460940 410592 460992 410644
rect 282828 410524 282880 410576
rect 462320 410524 462372 410576
rect 284300 410456 284352 410508
rect 340880 410456 340932 410508
rect 281724 409776 281776 409828
rect 292580 409776 292632 409828
rect 281724 408416 281776 408468
rect 338028 408416 338080 408468
rect 281632 403996 281684 404048
rect 283288 403996 283340 404048
rect 282828 402228 282880 402280
rect 286140 402228 286192 402280
rect 282828 401140 282880 401192
rect 286232 401140 286284 401192
rect 282828 400120 282880 400172
rect 337384 400120 337436 400172
rect 282276 400052 282328 400104
rect 292028 400052 292080 400104
rect 281632 398148 281684 398200
rect 283380 398148 283432 398200
rect 281632 397196 281684 397248
rect 284208 397196 284260 397248
rect 281632 396448 281684 396500
rect 283472 396448 283524 396500
rect 282184 396015 282236 396024
rect 282184 395981 282193 396015
rect 282193 395981 282227 396015
rect 282227 395981 282236 396015
rect 282184 395972 282236 395981
rect 281632 395768 281684 395820
rect 284116 395768 284168 395820
rect 281632 394340 281684 394392
rect 284024 394340 284076 394392
rect 281632 393184 281684 393236
rect 283840 393184 283892 393236
rect 281632 392028 281684 392080
rect 283932 392028 283984 392080
rect 281632 391620 281684 391672
rect 283748 391620 283800 391672
rect 281632 390124 281684 390176
rect 283656 390124 283708 390176
rect 281632 389036 281684 389088
rect 283564 389036 283616 389088
rect 281632 388288 281684 388340
rect 286968 388288 287020 388340
rect 281632 387064 281684 387116
rect 286876 387064 286928 387116
rect 282276 386384 282328 386436
rect 281632 386044 281684 386096
rect 286692 386044 286744 386096
rect 281632 385228 281684 385280
rect 286784 385228 286836 385280
rect 281632 384004 281684 384056
rect 284392 384004 284444 384056
rect 281632 383256 281684 383308
rect 284484 383256 284536 383308
rect 281816 382168 281868 382220
rect 339500 382168 339552 382220
rect 281632 382100 281684 382152
rect 284300 382100 284352 382152
rect 281632 380808 281684 380860
rect 338120 380808 338172 380860
rect 281632 379448 281684 379500
rect 336832 379448 336884 379500
rect 281632 378088 281684 378140
rect 336740 378088 336792 378140
rect 281816 378020 281868 378072
rect 335360 378020 335412 378072
rect 281632 376660 281684 376712
rect 333980 376660 334032 376712
rect 281632 375300 281684 375352
rect 332600 375300 332652 375352
rect 281816 373940 281868 373992
rect 329932 373940 329984 373992
rect 281632 373124 281684 373176
rect 287796 373124 287848 373176
rect 281632 371900 281684 371952
rect 286600 371900 286652 371952
rect 281816 371152 281868 371204
rect 327080 371152 327132 371204
rect 281632 370948 281684 371000
rect 285128 370948 285180 371000
rect 282276 369903 282328 369912
rect 282276 369869 282285 369903
rect 282285 369869 282319 369903
rect 282319 369869 282328 369903
rect 282276 369860 282328 369869
rect 281632 369792 281684 369844
rect 325700 369792 325752 369844
rect 281632 368432 281684 368484
rect 315304 368432 315356 368484
rect 282184 367140 282236 367192
rect 282092 367004 282144 367056
rect 284484 367004 284536 367056
rect 312544 367004 312596 367056
rect 285128 366936 285180 366988
rect 309784 366936 309836 366988
rect 281632 365644 281684 365696
rect 330484 365644 330536 365696
rect 282276 364964 282328 365016
rect 282736 364964 282788 365016
rect 281632 364284 281684 364336
rect 329288 364284 329340 364336
rect 281632 362856 281684 362908
rect 329104 362856 329156 362908
rect 281816 362788 281868 362840
rect 327724 362788 327776 362840
rect 281632 361496 281684 361548
rect 326344 361496 326396 361548
rect 281632 360136 281684 360188
rect 324964 360136 325016 360188
rect 281816 360068 281868 360120
rect 323584 360068 323636 360120
rect 281632 358708 281684 358760
rect 322204 358708 322256 358760
rect 282184 357416 282236 357468
rect 281632 351772 281684 351824
rect 286508 351772 286560 351824
rect 281632 350888 281684 350940
rect 286416 350888 286468 350940
rect 281632 350276 281684 350328
rect 284576 350276 284628 350328
rect 281632 349052 281684 349104
rect 291844 349052 291896 349104
rect 281632 347692 281684 347744
rect 290464 347692 290516 347744
rect 281632 346740 281684 346792
rect 287704 346740 287756 346792
rect 281632 345652 281684 345704
rect 286324 345652 286376 345704
rect 281632 344836 281684 344888
rect 284944 344836 284996 344888
rect 281632 343544 281684 343596
rect 307024 343544 307076 343596
rect 281816 343476 281868 343528
rect 291936 343476 291988 343528
rect 281632 342184 281684 342236
rect 308404 342184 308456 342236
rect 282276 340824 282328 340876
rect 282460 340824 282512 340876
rect 281632 340756 281684 340808
rect 284760 340756 284812 340808
rect 281724 340620 281776 340672
rect 284668 340620 284720 340672
rect 281632 338784 281684 338836
rect 284852 338784 284904 338836
rect 282460 338036 282512 338088
rect 281632 337900 281684 337952
rect 285588 337900 285640 337952
rect 281724 336676 281776 336728
rect 285404 336676 285456 336728
rect 281632 336540 281684 336592
rect 285496 336540 285548 336592
rect 281632 334568 281684 334620
rect 285312 334568 285364 334620
rect 281724 333888 281776 333940
rect 302884 333888 302936 333940
rect 281632 333616 281684 333668
rect 285220 333616 285272 333668
rect 281632 331168 281684 331220
rect 320272 331168 320324 331220
rect 281540 329740 281592 329792
rect 320180 329740 320232 329792
rect 281632 329672 281684 329724
rect 318800 329672 318852 329724
rect 282368 328491 282420 328500
rect 282368 328457 282377 328491
rect 282377 328457 282411 328491
rect 282411 328457 282420 328491
rect 282368 328448 282420 328457
rect 281540 328380 281592 328432
rect 317420 328380 317472 328432
rect 281540 325524 281592 325576
rect 285036 325524 285088 325576
rect 282828 321512 282880 321564
rect 338764 321512 338816 321564
rect 44088 318724 44140 318776
rect 130936 318724 130988 318776
rect 132868 318724 132920 318776
rect 133144 318724 133196 318776
rect 249708 318724 249760 318776
rect 343640 318724 343692 318776
rect 420184 318724 420236 318776
rect 453120 318724 453172 318776
rect 20628 318656 20680 318708
rect 92020 318656 92072 318708
rect 92388 318656 92440 318708
rect 210792 318656 210844 318708
rect 22008 318588 22060 318640
rect 93952 318588 94004 318640
rect 96528 318588 96580 318640
rect 216588 318588 216640 318640
rect 23388 318520 23440 318572
rect 97908 318520 97960 318572
rect 98000 318520 98052 318572
rect 218520 318520 218572 318572
rect 30288 318452 30340 318504
rect 107568 318452 107620 318504
rect 107660 318452 107712 318504
rect 234160 318452 234212 318504
rect 28908 318384 28960 318436
rect 105636 318384 105688 318436
rect 110328 318384 110380 318436
rect 239956 318384 240008 318436
rect 31668 318316 31720 318368
rect 111524 318316 111576 318368
rect 111708 318316 111760 318368
rect 241888 318316 241940 318368
rect 42708 318248 42760 318300
rect 129004 318248 129056 318300
rect 130384 318248 130436 318300
rect 261392 318248 261444 318300
rect 35808 318180 35860 318232
rect 117320 318180 117372 318232
rect 118608 318180 118660 318232
rect 253572 318180 253624 318232
rect 39948 318112 40000 318164
rect 125140 318112 125192 318164
rect 125508 318112 125560 318164
rect 265256 318112 265308 318164
rect 61384 318044 61436 318096
rect 343640 318044 343692 318096
rect 16488 317976 16540 318028
rect 86224 317976 86276 318028
rect 90916 317976 90968 318028
rect 206836 317976 206888 318028
rect 12348 317908 12400 317960
rect 78404 317908 78456 317960
rect 79968 317908 80020 317960
rect 189356 317908 189408 317960
rect 5448 317840 5500 317892
rect 68652 317840 68704 317892
rect 72976 317840 73028 317892
rect 177672 317840 177724 317892
rect 57888 317772 57940 317824
rect 154304 317772 154356 317824
rect 53748 317704 53800 317756
rect 146576 317704 146628 317756
rect 50988 317636 51040 317688
rect 142620 317636 142672 317688
rect 48136 317568 48188 317620
rect 136824 317568 136876 317620
rect 38476 317500 38528 317552
rect 123208 317500 123260 317552
rect 123484 317500 123536 317552
rect 131764 317500 131816 317552
rect 169852 317500 169904 317552
rect 33048 317432 33100 317484
rect 113456 317432 113508 317484
rect 124864 317432 124916 317484
rect 158168 317432 158220 317484
rect 49332 6128 49384 6180
rect 139400 6128 139452 6180
rect 80244 5448 80296 5500
rect 190460 5448 190512 5500
rect 83832 5380 83884 5432
rect 195980 5380 196032 5432
rect 87328 5312 87380 5364
rect 202880 5312 202932 5364
rect 91008 5244 91060 5296
rect 208400 5244 208452 5296
rect 94504 5176 94556 5228
rect 213920 5176 213972 5228
rect 98092 5108 98144 5160
rect 219440 5108 219492 5160
rect 101588 5040 101640 5092
rect 226340 5040 226392 5092
rect 105176 4972 105228 5024
rect 231860 4972 231912 5024
rect 67180 4904 67232 4956
rect 131764 4904 131816 4956
rect 266360 4904 266412 4956
rect 60004 4836 60056 4888
rect 124864 4836 124916 4888
rect 126612 4836 126664 4888
rect 130200 4836 130252 4888
rect 271880 4836 271932 4888
rect 37372 4768 37424 4820
rect 120080 4768 120132 4820
rect 123024 4768 123076 4820
rect 130384 4768 130436 4820
rect 131396 4768 131448 4820
rect 274640 4768 274692 4820
rect 76656 4700 76708 4752
rect 184940 4700 184992 4752
rect 73068 4632 73120 4684
rect 179420 4632 179472 4684
rect 69480 4564 69532 4616
rect 172520 4564 172572 4616
rect 65984 4496 66036 4548
rect 167000 4496 167052 4548
rect 62396 4428 62448 4480
rect 161480 4428 161532 4480
rect 58808 4360 58860 4412
rect 155960 4360 156012 4412
rect 55220 4292 55272 4344
rect 150440 4292 150492 4344
rect 51632 4224 51684 4276
rect 143540 4224 143592 4276
rect 46940 4156 46992 4208
rect 48136 4156 48188 4208
rect 48228 4156 48280 4208
rect 138020 4156 138072 4208
rect 81348 4088 81400 4140
rect 89720 4088 89772 4140
rect 93308 4088 93360 4140
rect 212540 4088 212592 4140
rect 14832 4020 14884 4072
rect 55312 4020 55364 4072
rect 64696 4020 64748 4072
rect 81440 4020 81492 4072
rect 82636 4020 82688 4072
rect 223580 4020 223632 4072
rect 13636 3952 13688 4004
rect 17224 3952 17276 4004
rect 86960 3952 87012 4004
rect 99288 3952 99340 4004
rect 222200 3952 222252 4004
rect 18328 3884 18380 3936
rect 84936 3884 84988 3936
rect 102784 3884 102836 3936
rect 227720 3884 227772 3936
rect 19524 3816 19576 3868
rect 20628 3816 20680 3868
rect 20720 3816 20772 3868
rect 22008 3816 22060 3868
rect 21916 3748 21968 3800
rect 95240 3816 95292 3868
rect 99380 3816 99432 3868
rect 100484 3816 100536 3868
rect 25504 3748 25556 3800
rect 100760 3748 100812 3800
rect 107476 3748 107528 3800
rect 236000 3816 236052 3868
rect 114744 3748 114796 3800
rect 247040 3748 247092 3800
rect 24308 3680 24360 3732
rect 95700 3680 95752 3732
rect 96528 3680 96580 3732
rect 96896 3680 96948 3732
rect 97908 3680 97960 3732
rect 113548 3680 113600 3732
rect 245660 3680 245712 3732
rect 26700 3612 26752 3664
rect 103520 3612 103572 3664
rect 34980 3544 35032 3596
rect 35808 3544 35860 3596
rect 109040 3612 109092 3664
rect 117136 3612 117188 3664
rect 251180 3612 251232 3664
rect 103980 3544 104032 3596
rect 104808 3544 104860 3596
rect 106372 3544 106424 3596
rect 107568 3544 107620 3596
rect 111156 3544 111208 3596
rect 111708 3544 111760 3596
rect 119436 3544 119488 3596
rect 255320 3544 255372 3596
rect 11244 3476 11296 3528
rect 12348 3476 12400 3528
rect 16028 3476 16080 3528
rect 16488 3476 16540 3528
rect 27896 3476 27948 3528
rect 28908 3476 28960 3528
rect 29092 3476 29144 3528
rect 30288 3476 30340 3528
rect 33876 3476 33928 3528
rect 114560 3476 114612 3528
rect 120632 3476 120684 3528
rect 256700 3476 256752 3528
rect 30196 3408 30248 3460
rect 36176 3408 36228 3460
rect 118700 3408 118752 3460
rect 124220 3408 124272 3460
rect 262220 3408 262272 3460
rect 12440 3340 12492 3392
rect 63684 3340 63736 3392
rect 10048 3272 10100 3324
rect 71872 3272 71924 3324
rect 72976 3272 73028 3324
rect 8852 3204 8904 3256
rect 74540 3272 74592 3324
rect 79048 3340 79100 3392
rect 79968 3340 80020 3392
rect 84200 3340 84252 3392
rect 89720 3340 89772 3392
rect 90916 3340 90968 3392
rect 80152 3272 80204 3324
rect 88524 3272 88576 3324
rect 204260 3340 204312 3392
rect 86132 3204 86184 3256
rect 200120 3272 200172 3324
rect 198740 3204 198792 3256
rect 1676 3136 1728 3188
rect 7656 3136 7708 3188
rect 6460 3068 6512 3120
rect 4068 3000 4120 3052
rect 66352 3000 66404 3052
rect 76012 3136 76064 3188
rect 77852 3136 77904 3188
rect 186320 3136 186372 3188
rect 70400 3068 70452 3120
rect 71964 3068 72016 3120
rect 75460 3068 75512 3120
rect 183560 3068 183612 3120
rect 70676 3000 70728 3052
rect 175280 3000 175332 3052
rect 572 2932 624 2984
rect 61384 2932 61436 2984
rect 68284 2932 68336 2984
rect 171140 2932 171192 2984
rect 2872 2796 2924 2848
rect 61200 2864 61252 2916
rect 160100 2864 160152 2916
rect 62212 2796 62264 2848
rect 63592 2796 63644 2848
rect 162860 2796 162912 2848
rect 5264 552 5316 604
rect 5448 552 5500 604
rect 74264 552 74316 604
rect 74448 552 74500 604
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 263600 653404 263652 653410
rect 263600 653346 263652 653352
rect 378140 653404 378192 653410
rect 378140 653346 378192 653352
rect 383568 653404 383620 653410
rect 383568 653346 383620 653352
rect 508412 653404 508464 653410
rect 508412 653346 508464 653352
rect 139400 652860 139452 652866
rect 139400 652802 139452 652808
rect 135168 652792 135220 652798
rect 135088 652752 135168 652780
rect 135088 651137 135116 652752
rect 135168 652734 135220 652740
rect 135074 651128 135130 651137
rect 135074 651063 135130 651072
rect 137652 650276 137704 650282
rect 137652 650218 137704 650224
rect 137664 649720 137692 650218
rect 137650 649711 137706 649720
rect 137650 649646 137706 649655
rect 57886 646096 57942 646105
rect 57886 646031 57942 646040
rect 57794 645008 57850 645017
rect 57794 644943 57850 644952
rect 57702 643240 57758 643249
rect 57702 643175 57758 643184
rect 57610 642016 57666 642025
rect 57610 641951 57666 641960
rect 57518 640384 57574 640393
rect 57518 640319 57574 640328
rect 57426 639296 57482 639305
rect 57426 639231 57482 639240
rect 57334 637664 57390 637673
rect 57334 637599 57390 637608
rect 57242 579728 57298 579737
rect 57242 579663 57298 579672
rect 57256 543114 57284 579663
rect 57244 543108 57296 543114
rect 57244 543050 57296 543056
rect 57348 542978 57376 637599
rect 57440 543522 57468 639231
rect 57428 543516 57480 543522
rect 57428 543458 57480 543464
rect 57532 543454 57560 640319
rect 57520 543448 57572 543454
rect 57520 543390 57572 543396
rect 57624 543386 57652 641951
rect 57612 543380 57664 543386
rect 57612 543322 57664 543328
rect 57716 543250 57744 643175
rect 57808 543862 57836 644943
rect 57900 543930 57928 646031
rect 139412 589665 139440 652802
rect 258540 652792 258592 652798
rect 258540 652734 258592 652740
rect 258552 651681 258580 652734
rect 263612 651681 263640 653346
rect 378152 652934 378180 653346
rect 383580 652934 383608 653346
rect 378140 652928 378192 652934
rect 378138 652896 378140 652905
rect 383568 652928 383620 652934
rect 378192 652896 378194 652905
rect 378138 652831 378194 652840
rect 383566 652896 383568 652905
rect 508424 652905 508452 653346
rect 383620 652896 383622 652905
rect 383566 652831 383622 652840
rect 508410 652896 508466 652905
rect 508410 652831 508412 652840
rect 383580 652805 383608 652831
rect 508464 652831 508466 652840
rect 513378 652896 513434 652905
rect 513378 652831 513380 652840
rect 508412 652802 508464 652808
rect 513432 652831 513434 652840
rect 513380 652802 513432 652808
rect 508424 652771 508452 652802
rect 518900 652792 518952 652798
rect 518900 652734 518952 652740
rect 258538 651672 258594 651681
rect 258538 651607 258594 651616
rect 263598 651672 263654 651681
rect 263598 651607 263654 651616
rect 407764 650548 407816 650554
rect 407764 650490 407816 650496
rect 266636 650480 266688 650486
rect 266636 650422 266688 650428
rect 387156 650480 387208 650486
rect 387156 650422 387208 650428
rect 266648 649913 266676 650422
rect 387168 649913 387196 650422
rect 389180 650208 389232 650214
rect 389180 650150 389232 650156
rect 389192 649913 389220 650150
rect 266634 649904 266690 649913
rect 266634 649839 266690 649848
rect 387154 649904 387210 649913
rect 387154 649839 387210 649848
rect 389178 649904 389234 649913
rect 389178 649839 389234 649848
rect 188342 646096 188398 646105
rect 188342 646031 188398 646040
rect 307390 646096 307446 646105
rect 307390 646031 307446 646040
rect 139398 589656 139454 589665
rect 139398 589591 139454 589600
rect 67546 558920 67602 558929
rect 67546 558855 67602 558864
rect 68926 558920 68982 558929
rect 68926 558855 68982 558864
rect 70306 558920 70362 558929
rect 70306 558855 70362 558864
rect 71686 558920 71742 558929
rect 71686 558855 71742 558864
rect 72514 558920 72570 558929
rect 72514 558855 72570 558864
rect 73066 558920 73122 558929
rect 73066 558855 73122 558864
rect 73710 558920 73766 558929
rect 73710 558855 73766 558864
rect 74262 558920 74318 558929
rect 74262 558855 74318 558864
rect 74998 558920 75054 558929
rect 74998 558855 75054 558864
rect 75826 558920 75882 558929
rect 75826 558855 75882 558864
rect 76838 558920 76894 558929
rect 76838 558855 76894 558864
rect 77390 558920 77446 558929
rect 77390 558855 77392 558864
rect 66168 558816 66220 558822
rect 66168 558758 66220 558764
rect 62026 558376 62082 558385
rect 62026 558311 62082 558320
rect 57888 543924 57940 543930
rect 57888 543866 57940 543872
rect 57796 543856 57848 543862
rect 57796 543798 57848 543804
rect 62040 543590 62068 558311
rect 63406 558240 63462 558249
rect 63406 558175 63462 558184
rect 61016 543584 61068 543590
rect 61016 543526 61068 543532
rect 62028 543584 62080 543590
rect 62028 543526 62080 543532
rect 57704 543244 57756 543250
rect 57704 543186 57756 543192
rect 57336 542972 57388 542978
rect 57336 542914 57388 542920
rect 61028 539988 61056 543526
rect 63420 540002 63448 558175
rect 66180 543590 66208 558758
rect 67456 557592 67508 557598
rect 67456 557534 67508 557540
rect 65156 543584 65208 543590
rect 65156 543526 65208 543532
rect 66168 543584 66220 543590
rect 66168 543526 66220 543532
rect 63066 539974 63448 540002
rect 65168 539988 65196 543526
rect 67468 540002 67496 557534
rect 67560 543046 67588 558855
rect 67548 543040 67600 543046
rect 67548 542982 67600 542988
rect 68940 542450 68968 558855
rect 70214 558648 70270 558657
rect 70214 558583 70270 558592
rect 70228 543590 70256 558583
rect 70320 543658 70348 558855
rect 71700 543726 71728 558855
rect 72528 558210 72556 558855
rect 72516 558204 72568 558210
rect 72516 558146 72568 558152
rect 73080 543998 73108 558855
rect 73724 558414 73752 558855
rect 73712 558408 73764 558414
rect 73712 558350 73764 558356
rect 74276 558278 74304 558855
rect 75012 558754 75040 558855
rect 75000 558748 75052 558754
rect 75000 558690 75052 558696
rect 74264 558272 74316 558278
rect 74264 558214 74316 558220
rect 73068 543992 73120 543998
rect 73068 543934 73120 543940
rect 75840 543726 75868 558855
rect 75918 558648 75974 558657
rect 75918 558583 75920 558592
rect 75972 558583 75974 558592
rect 75920 558554 75972 558560
rect 76852 558142 76880 558855
rect 77444 558855 77446 558864
rect 78586 558920 78642 558929
rect 78586 558855 78642 558864
rect 79322 558920 79378 558929
rect 79322 558855 79378 558864
rect 79874 558920 79930 558929
rect 79874 558855 79930 558864
rect 80794 558920 80850 558929
rect 80794 558855 80850 558864
rect 81254 558920 81310 558929
rect 81254 558855 81310 558864
rect 81990 558920 82046 558929
rect 81990 558855 82046 558864
rect 82910 558920 82966 558929
rect 82910 558855 82966 558864
rect 83830 558920 83886 558929
rect 83830 558855 83886 558864
rect 84198 558920 84254 558929
rect 84198 558855 84254 558864
rect 85486 558920 85542 558929
rect 85486 558855 85542 558864
rect 86314 558920 86370 558929
rect 86774 558920 86830 558929
rect 86314 558855 86316 558864
rect 77392 558826 77444 558832
rect 78496 558680 78548 558686
rect 78494 558648 78496 558657
rect 78548 558648 78550 558657
rect 78494 558583 78550 558592
rect 76840 558136 76892 558142
rect 76840 558078 76892 558084
rect 71688 543720 71740 543726
rect 71688 543662 71740 543668
rect 75460 543720 75512 543726
rect 75460 543662 75512 543668
rect 75828 543720 75880 543726
rect 75828 543662 75880 543668
rect 70308 543652 70360 543658
rect 70308 543594 70360 543600
rect 73436 543652 73488 543658
rect 73436 543594 73488 543600
rect 70216 543584 70268 543590
rect 70216 543526 70268 543532
rect 71320 543584 71372 543590
rect 71320 543526 71372 543532
rect 68940 542422 69060 542450
rect 67206 539974 67496 540002
rect 69032 540002 69060 542422
rect 69032 539974 69322 540002
rect 71332 539988 71360 543526
rect 73448 539988 73476 543594
rect 75472 539988 75500 543662
rect 78600 543658 78628 558855
rect 79336 558006 79364 558855
rect 79414 558648 79470 558657
rect 79414 558583 79470 558592
rect 79428 558550 79456 558583
rect 79416 558544 79468 558550
rect 79416 558486 79468 558492
rect 79324 558000 79376 558006
rect 79324 557942 79376 557948
rect 78588 543652 78640 543658
rect 78588 543594 78640 543600
rect 79888 543590 79916 558855
rect 80808 558482 80836 558855
rect 80796 558476 80848 558482
rect 80796 558418 80848 558424
rect 81268 558074 81296 558855
rect 82004 558346 82032 558855
rect 82924 558414 82952 558855
rect 82912 558408 82964 558414
rect 82912 558350 82964 558356
rect 81440 558340 81492 558346
rect 81440 558282 81492 558288
rect 81992 558340 82044 558346
rect 81992 558282 82044 558288
rect 81452 558210 81480 558282
rect 83844 558210 83872 558855
rect 84212 558754 84240 558855
rect 84200 558748 84252 558754
rect 84200 558690 84252 558696
rect 85394 558648 85450 558657
rect 85394 558583 85396 558592
rect 85448 558583 85450 558592
rect 85396 558554 85448 558560
rect 81440 558204 81492 558210
rect 81440 558146 81492 558152
rect 83832 558204 83884 558210
rect 83832 558146 83884 558152
rect 81256 558068 81308 558074
rect 81256 558010 81308 558016
rect 82726 557968 82782 557977
rect 82726 557903 82782 557912
rect 81716 544400 81768 544406
rect 81716 544342 81768 544348
rect 79876 543584 79928 543590
rect 79876 543526 79928 543532
rect 79692 543108 79744 543114
rect 79692 543050 79744 543056
rect 77574 543008 77630 543017
rect 77574 542943 77630 542952
rect 77588 539988 77616 542943
rect 79704 539988 79732 543050
rect 81728 539988 81756 544342
rect 82740 544066 82768 557903
rect 85408 557734 85436 558554
rect 85396 557728 85448 557734
rect 85396 557670 85448 557676
rect 83832 544468 83884 544474
rect 83832 544410 83884 544416
rect 82728 544060 82780 544066
rect 82728 544002 82780 544008
rect 83844 539988 83872 544410
rect 85500 544202 85528 558855
rect 86368 558855 86370 558864
rect 86684 558884 86736 558890
rect 86316 558826 86368 558832
rect 86774 558855 86830 558864
rect 87878 558920 87934 558929
rect 87878 558855 87934 558864
rect 88246 558920 88302 558929
rect 88246 558855 88302 558864
rect 88890 558920 88946 558929
rect 88890 558855 88946 558864
rect 89166 558920 89222 558929
rect 89166 558855 89222 558864
rect 89810 558920 89866 558929
rect 89810 558855 89866 558864
rect 91006 558920 91062 558929
rect 91006 558855 91062 558864
rect 92202 558920 92258 558929
rect 92202 558855 92258 558864
rect 92478 558920 92534 558929
rect 92478 558855 92534 558864
rect 93306 558920 93362 558929
rect 93306 558855 93362 558864
rect 93766 558920 93822 558929
rect 93766 558855 93768 558864
rect 86684 558826 86736 558832
rect 86696 558618 86724 558826
rect 86684 558612 86736 558618
rect 86684 558554 86736 558560
rect 85856 544536 85908 544542
rect 85856 544478 85908 544484
rect 85488 544196 85540 544202
rect 85488 544138 85540 544144
rect 85868 539988 85896 544478
rect 86788 544338 86816 558855
rect 87892 558686 87920 558855
rect 87880 558680 87932 558686
rect 86866 558648 86922 558657
rect 87880 558622 87932 558628
rect 86866 558583 86922 558592
rect 86776 544332 86828 544338
rect 86776 544274 86828 544280
rect 86880 544134 86908 558583
rect 87972 544672 88024 544678
rect 87972 544614 88024 544620
rect 86868 544128 86920 544134
rect 86868 544070 86920 544076
rect 87984 539988 88012 544614
rect 88260 544270 88288 558855
rect 88904 558550 88932 558855
rect 88892 558544 88944 558550
rect 88892 558486 88944 558492
rect 89180 557870 89208 558855
rect 89824 558482 89852 558855
rect 89812 558476 89864 558482
rect 89812 558418 89864 558424
rect 89168 557864 89220 557870
rect 89168 557806 89220 557812
rect 89996 544808 90048 544814
rect 89996 544750 90048 544756
rect 88248 544264 88300 544270
rect 88248 544206 88300 544212
rect 90008 539988 90036 544750
rect 91020 543318 91048 558855
rect 91098 558648 91154 558657
rect 91098 558583 91154 558592
rect 91112 558346 91140 558583
rect 92216 558346 92244 558855
rect 92492 558414 92520 558855
rect 93320 558754 93348 558855
rect 93820 558855 93822 558864
rect 95054 558920 95110 558929
rect 95054 558855 95110 558864
rect 95698 558920 95754 558929
rect 95698 558855 95754 558864
rect 96526 558920 96582 558929
rect 96526 558855 96582 558864
rect 97170 558920 97226 558929
rect 97170 558855 97226 558864
rect 97814 558920 97870 558929
rect 97814 558855 97870 558864
rect 98366 558920 98422 558929
rect 98366 558855 98422 558864
rect 99286 558920 99342 558929
rect 99286 558855 99342 558864
rect 100022 558920 100078 558929
rect 100022 558855 100078 558864
rect 102046 558920 102102 558929
rect 102046 558855 102102 558864
rect 104806 558920 104862 558929
rect 104806 558855 104862 558864
rect 107290 558920 107346 558929
rect 107290 558855 107346 558864
rect 108486 558920 108542 558929
rect 108486 558855 108542 558864
rect 137284 558884 137336 558890
rect 93768 558826 93820 558832
rect 93308 558748 93360 558754
rect 93308 558690 93360 558696
rect 93674 558648 93730 558657
rect 93674 558583 93730 558592
rect 94778 558648 94834 558657
rect 94778 558583 94834 558592
rect 92480 558408 92532 558414
rect 92480 558350 92532 558356
rect 93124 558408 93176 558414
rect 93124 558350 93176 558356
rect 91100 558340 91152 558346
rect 91100 558282 91152 558288
rect 92204 558340 92256 558346
rect 92204 558282 92256 558288
rect 91112 557666 91140 558282
rect 93136 557802 93164 558350
rect 93124 557796 93176 557802
rect 93124 557738 93176 557744
rect 91100 557660 91152 557666
rect 91100 557602 91152 557608
rect 92112 544876 92164 544882
rect 92112 544818 92164 544824
rect 91008 543312 91060 543318
rect 91008 543254 91060 543260
rect 92124 539988 92152 544818
rect 93688 543182 93716 558583
rect 94792 558482 94820 558583
rect 94780 558476 94832 558482
rect 94780 558418 94832 558424
rect 94792 557734 94820 558418
rect 94780 557728 94832 557734
rect 94780 557670 94832 557676
rect 94136 545012 94188 545018
rect 94136 544954 94188 544960
rect 93676 543176 93728 543182
rect 93676 543118 93728 543124
rect 94148 539988 94176 544954
rect 95068 543114 95096 558855
rect 95712 558618 95740 558855
rect 95700 558612 95752 558618
rect 95700 558554 95752 558560
rect 96540 545086 96568 558855
rect 97184 558686 97212 558855
rect 97172 558680 97224 558686
rect 97172 558622 97224 558628
rect 97184 557938 97212 558622
rect 97828 558414 97856 558855
rect 98380 558550 98408 558855
rect 98368 558544 98420 558550
rect 98368 558486 98420 558492
rect 97816 558408 97868 558414
rect 97816 558350 97868 558356
rect 97172 557932 97224 557938
rect 97172 557874 97224 557880
rect 98380 557734 98408 558486
rect 98368 557728 98420 557734
rect 98368 557670 98420 557676
rect 96528 545080 96580 545086
rect 96528 545022 96580 545028
rect 96250 543280 96306 543289
rect 96250 543215 96306 543224
rect 95056 543108 95108 543114
rect 95056 543050 95108 543056
rect 96264 539988 96292 543215
rect 99300 543046 99328 558855
rect 99472 558680 99524 558686
rect 99472 558622 99524 558628
rect 99484 558521 99512 558622
rect 100036 558550 100064 558855
rect 102060 558686 102088 558855
rect 102784 558748 102836 558754
rect 102784 558690 102836 558696
rect 102048 558680 102100 558686
rect 102048 558622 102100 558628
rect 100024 558544 100076 558550
rect 99470 558512 99526 558521
rect 100024 558486 100076 558492
rect 100390 558512 100446 558521
rect 99470 558447 99526 558456
rect 100390 558447 100446 558456
rect 100022 557696 100078 557705
rect 100404 557666 100432 558447
rect 100850 557832 100906 557841
rect 100850 557767 100852 557776
rect 100904 557767 100906 557776
rect 101402 557832 101458 557841
rect 101402 557767 101458 557776
rect 100852 557738 100904 557744
rect 100022 557631 100024 557640
rect 100076 557631 100078 557640
rect 100392 557660 100444 557666
rect 100024 557602 100076 557608
rect 100392 557602 100444 557608
rect 98368 543040 98420 543046
rect 98368 542982 98420 542988
rect 99288 543040 99340 543046
rect 99288 542982 99340 542988
rect 98380 539988 98408 542982
rect 100036 542706 100064 557602
rect 100392 542972 100444 542978
rect 100392 542914 100444 542920
rect 100024 542700 100076 542706
rect 100024 542642 100076 542648
rect 100404 539988 100432 542914
rect 101416 542638 101444 557767
rect 102796 557569 102824 558690
rect 104164 558612 104216 558618
rect 104164 558554 104216 558560
rect 104176 557569 104204 558554
rect 104820 558550 104848 558855
rect 107304 558754 107332 558855
rect 106280 558748 106332 558754
rect 106280 558690 106332 558696
rect 107292 558748 107344 558754
rect 107292 558690 107344 558696
rect 106292 558657 106320 558690
rect 106278 558648 106334 558657
rect 108500 558618 108528 558855
rect 137284 558826 137336 558832
rect 106278 558583 106334 558592
rect 108488 558612 108540 558618
rect 108488 558554 108540 558560
rect 104808 558544 104860 558550
rect 104808 558486 104860 558492
rect 108486 558512 108542 558521
rect 108486 558447 108542 558456
rect 110326 558512 110382 558521
rect 110326 558447 110382 558456
rect 108302 557968 108358 557977
rect 105544 557932 105596 557938
rect 108302 557903 108358 557912
rect 105544 557874 105596 557880
rect 105556 557569 105584 557874
rect 108316 557734 108344 557903
rect 108304 557728 108356 557734
rect 106922 557696 106978 557705
rect 108304 557670 108356 557676
rect 106922 557631 106978 557640
rect 102046 557560 102102 557569
rect 102046 557495 102102 557504
rect 102782 557560 102838 557569
rect 102782 557495 102838 557504
rect 103426 557560 103482 557569
rect 103426 557495 103482 557504
rect 104162 557560 104218 557569
rect 104162 557495 104218 557504
rect 105542 557560 105598 557569
rect 105542 557495 105598 557504
rect 106186 557560 106242 557569
rect 106186 557495 106242 557504
rect 102060 544950 102088 557495
rect 102048 544944 102100 544950
rect 102048 544886 102100 544892
rect 102508 543516 102560 543522
rect 102508 543458 102560 543464
rect 101404 542632 101456 542638
rect 101404 542574 101456 542580
rect 102520 539988 102548 543458
rect 102796 542842 102824 557495
rect 103440 543153 103468 557495
rect 103426 543144 103482 543153
rect 103426 543079 103482 543088
rect 102784 542836 102836 542842
rect 102784 542778 102836 542784
rect 104176 542774 104204 557495
rect 104532 543448 104584 543454
rect 104532 543390 104584 543396
rect 104164 542768 104216 542774
rect 104164 542710 104216 542716
rect 104544 539988 104572 543390
rect 105556 542910 105584 557495
rect 106200 544746 106228 557495
rect 106188 544740 106240 544746
rect 106188 544682 106240 544688
rect 106648 543380 106700 543386
rect 106648 543322 106700 543328
rect 105544 542904 105596 542910
rect 105544 542846 105596 542852
rect 106660 539988 106688 543322
rect 106936 542502 106964 557631
rect 108316 542978 108344 557670
rect 108500 557666 108528 558447
rect 108488 557660 108540 557666
rect 108488 557602 108540 557608
rect 108304 542972 108356 542978
rect 108304 542914 108356 542920
rect 108500 542570 108528 557602
rect 110340 544610 110368 558447
rect 129648 557932 129700 557938
rect 129648 557874 129700 557880
rect 125508 557864 125560 557870
rect 125508 557806 125560 557812
rect 121368 557796 121420 557802
rect 121368 557738 121420 557744
rect 117228 557728 117280 557734
rect 117228 557670 117280 557676
rect 110328 544604 110380 544610
rect 110328 544546 110380 544552
rect 112812 543924 112864 543930
rect 112812 543866 112864 543872
rect 110788 543856 110840 543862
rect 110788 543798 110840 543804
rect 108672 543244 108724 543250
rect 108672 543186 108724 543192
rect 108488 542564 108540 542570
rect 108488 542506 108540 542512
rect 106924 542496 106976 542502
rect 106924 542438 106976 542444
rect 108684 539988 108712 543186
rect 110800 539988 110828 543798
rect 112824 539988 112852 543866
rect 114928 543244 114980 543250
rect 114928 543186 114980 543192
rect 114940 539988 114968 543186
rect 117240 540002 117268 557670
rect 119068 543380 119120 543386
rect 119068 543322 119120 543328
rect 117070 539974 117268 540002
rect 119080 539988 119108 543322
rect 121380 540002 121408 557738
rect 123208 543448 123260 543454
rect 123208 543390 123260 543396
rect 121210 539974 121408 540002
rect 123220 539988 123248 543390
rect 125520 540002 125548 557806
rect 127348 543516 127400 543522
rect 127348 543458 127400 543464
rect 125350 539974 125548 540002
rect 127360 539988 127388 543458
rect 129660 540002 129688 557874
rect 131764 556912 131816 556918
rect 131764 556854 131816 556860
rect 131776 542706 131804 556854
rect 137296 542842 137324 558826
rect 141424 558748 141476 558754
rect 141424 558690 141476 558696
rect 140044 558680 140096 558686
rect 140044 558622 140096 558628
rect 138664 558408 138716 558414
rect 138664 558350 138716 558356
rect 137468 558340 137520 558346
rect 137468 558282 137520 558288
rect 137376 558272 137428 558278
rect 137376 558214 137428 558220
rect 135720 542836 135772 542842
rect 135720 542778 135772 542784
rect 137284 542836 137336 542842
rect 137284 542778 137336 542784
rect 131488 542700 131540 542706
rect 131488 542642 131540 542648
rect 131764 542700 131816 542706
rect 131764 542642 131816 542648
rect 129490 539974 129688 540002
rect 131500 539988 131528 542642
rect 133604 542632 133656 542638
rect 133604 542574 133656 542580
rect 133616 539988 133644 542574
rect 135732 539988 135760 542778
rect 137388 542434 137416 558214
rect 137480 542638 137508 558282
rect 138676 542842 138704 558350
rect 140056 543697 140084 558622
rect 140136 558476 140188 558482
rect 140136 558418 140188 558424
rect 140042 543688 140098 543697
rect 140042 543623 140098 543632
rect 140148 542910 140176 558418
rect 141436 543425 141464 558690
rect 148324 558612 148376 558618
rect 148324 558554 148376 558560
rect 144184 558544 144236 558550
rect 144184 558486 144236 558492
rect 141422 543416 141478 543425
rect 141422 543351 141478 543360
rect 144196 542978 144224 558486
rect 145564 558136 145616 558142
rect 145564 558078 145616 558084
rect 145576 543726 145604 558078
rect 148140 543992 148192 543998
rect 148140 543934 148192 543940
rect 145564 543720 145616 543726
rect 145564 543662 145616 543668
rect 144000 542972 144052 542978
rect 144000 542914 144052 542920
rect 144184 542972 144236 542978
rect 144184 542914 144236 542920
rect 139860 542904 139912 542910
rect 139860 542846 139912 542852
rect 140136 542904 140188 542910
rect 140136 542846 140188 542852
rect 138664 542836 138716 542842
rect 138664 542778 138716 542784
rect 137744 542768 137796 542774
rect 137744 542710 137796 542716
rect 137468 542632 137520 542638
rect 137468 542574 137520 542580
rect 137376 542428 137428 542434
rect 137376 542370 137428 542376
rect 137756 539988 137784 542710
rect 139872 539988 139900 542846
rect 141884 542496 141936 542502
rect 141884 542438 141936 542444
rect 141896 539988 141924 542438
rect 144012 539988 144040 542914
rect 146024 542564 146076 542570
rect 146024 542506 146076 542512
rect 146036 539988 146064 542506
rect 148152 539988 148180 543934
rect 148336 543561 148364 558554
rect 149704 558204 149756 558210
rect 149704 558146 149756 558152
rect 148322 543552 148378 543561
rect 148322 543487 148378 543496
rect 149716 542502 149744 558146
rect 152556 558068 152608 558074
rect 152556 558010 152608 558016
rect 152464 558000 152516 558006
rect 152464 557942 152516 557948
rect 152476 543590 152504 557942
rect 152568 543726 152596 558010
rect 173072 544332 173124 544338
rect 173072 544274 173124 544280
rect 168840 544196 168892 544202
rect 168840 544138 168892 544144
rect 164700 544060 164752 544066
rect 164700 544002 164752 544008
rect 152556 543720 152608 543726
rect 152556 543662 152608 543668
rect 162676 543720 162728 543726
rect 162676 543662 162728 543668
rect 156420 543652 156472 543658
rect 156420 543594 156472 543600
rect 152464 543584 152516 543590
rect 152464 543526 152516 543532
rect 152280 542564 152332 542570
rect 152280 542506 152332 542512
rect 154396 542564 154448 542570
rect 154396 542506 154448 542512
rect 149704 542496 149756 542502
rect 149704 542438 149756 542444
rect 150164 542428 150216 542434
rect 150164 542370 150216 542376
rect 150176 539988 150204 542370
rect 152292 539988 152320 542506
rect 154408 539988 154436 542506
rect 156432 539988 156460 543594
rect 158536 543584 158588 543590
rect 158536 543526 158588 543532
rect 158548 539988 158576 543526
rect 160560 542428 160612 542434
rect 160560 542370 160612 542376
rect 160572 539988 160600 542370
rect 162688 539988 162716 543662
rect 164712 539988 164740 544002
rect 166816 542564 166868 542570
rect 166816 542506 166868 542512
rect 166828 539988 166856 542506
rect 168852 539988 168880 544138
rect 170956 544128 171008 544134
rect 170956 544070 171008 544076
rect 170968 539988 170996 544070
rect 173084 539988 173112 544274
rect 175096 544264 175148 544270
rect 175096 544206 175148 544212
rect 175108 539988 175136 544206
rect 179236 543312 179288 543318
rect 188356 543289 188384 646031
rect 307404 645930 307432 646031
rect 291844 645924 291896 645930
rect 291844 645866 291896 645872
rect 307392 645924 307444 645930
rect 307392 645866 307444 645872
rect 188434 645008 188490 645017
rect 188434 644943 188490 644952
rect 188448 545018 188476 644943
rect 290464 644496 290516 644502
rect 290464 644438 290516 644444
rect 188526 643240 188582 643249
rect 188526 643175 188582 643184
rect 188436 545012 188488 545018
rect 188436 544954 188488 544960
rect 188540 544882 188568 643175
rect 287704 643136 287756 643142
rect 287704 643078 287756 643084
rect 188618 642016 188674 642025
rect 188618 641951 188674 641960
rect 188528 544876 188580 544882
rect 188528 544818 188580 544824
rect 188632 544814 188660 641951
rect 286324 641776 286376 641782
rect 286324 641718 286376 641724
rect 188710 640384 188766 640393
rect 188710 640319 188766 640328
rect 284944 640348 284996 640354
rect 188620 544808 188672 544814
rect 188620 544750 188672 544756
rect 188724 544678 188752 640319
rect 284944 640290 284996 640296
rect 188802 639296 188858 639305
rect 188802 639231 188858 639240
rect 188712 544672 188764 544678
rect 188712 544614 188764 544620
rect 188816 544542 188844 639231
rect 188894 637664 188950 637673
rect 188894 637599 188950 637608
rect 188804 544536 188856 544542
rect 188804 544478 188856 544484
rect 188908 544474 188936 637599
rect 269118 589384 269174 589393
rect 269118 589319 269174 589328
rect 269132 587217 269160 589319
rect 269118 587208 269174 587217
rect 269118 587143 269174 587152
rect 270406 580408 270462 580417
rect 270406 580343 270462 580352
rect 270420 580310 270448 580343
rect 270408 580304 270460 580310
rect 270408 580246 270460 580252
rect 279148 580304 279200 580310
rect 279148 580246 279200 580252
rect 188986 579728 189042 579737
rect 188986 579663 189042 579672
rect 188896 544468 188948 544474
rect 188896 544410 188948 544416
rect 179236 543254 179288 543260
rect 188342 543280 188398 543289
rect 177212 542700 177264 542706
rect 177212 542642 177264 542648
rect 177224 539988 177252 542642
rect 179248 539988 179276 543254
rect 188342 543215 188398 543224
rect 183376 543176 183428 543182
rect 183376 543118 183428 543124
rect 181352 542632 181404 542638
rect 181352 542574 181404 542580
rect 181364 539988 181392 542574
rect 183388 539988 183416 543118
rect 187516 543108 187568 543114
rect 187516 543050 187568 543056
rect 185492 542768 185544 542774
rect 185492 542710 185544 542716
rect 185504 539988 185532 542710
rect 187528 539988 187556 543050
rect 189000 543017 189028 579663
rect 210974 560008 211030 560017
rect 210974 559943 211030 559952
rect 195978 558920 196034 558929
rect 194416 558884 194468 558890
rect 195978 558855 196034 558864
rect 200210 558920 200266 558929
rect 200210 558855 200266 558864
rect 202786 558920 202842 558929
rect 202786 558855 202842 558864
rect 203798 558920 203854 558929
rect 203798 558855 203854 558864
rect 204166 558920 204222 558929
rect 204166 558855 204222 558864
rect 205546 558920 205602 558929
rect 205546 558855 205602 558864
rect 206926 558920 206982 558929
rect 206926 558855 206982 558864
rect 208490 558920 208546 558929
rect 208490 558855 208546 558864
rect 210606 558920 210662 558929
rect 210606 558855 210662 558864
rect 194416 558826 194468 558832
rect 194428 558793 194456 558826
rect 194414 558784 194470 558793
rect 194414 558719 194470 558728
rect 189632 545080 189684 545086
rect 189632 545022 189684 545028
rect 188986 543008 189042 543017
rect 188986 542943 189042 542952
rect 189644 539988 189672 545022
rect 195992 544406 196020 558855
rect 200224 558822 200252 558855
rect 200212 558816 200264 558822
rect 200212 558758 200264 558764
rect 202142 558648 202198 558657
rect 202142 558583 202198 558592
rect 201498 557696 201554 557705
rect 202156 557666 202184 558583
rect 201498 557631 201554 557640
rect 202144 557660 202196 557666
rect 201512 557598 201540 557631
rect 202144 557602 202196 557608
rect 201500 557592 201552 557598
rect 201500 557534 201552 557540
rect 197912 544944 197964 544950
rect 197912 544886 197964 544892
rect 195980 544400 196032 544406
rect 195980 544342 196032 544348
rect 193772 543040 193824 543046
rect 193772 542982 193824 542988
rect 191748 542836 191800 542842
rect 191748 542778 191800 542784
rect 191760 539988 191788 542778
rect 193784 539988 193812 542982
rect 195888 542904 195940 542910
rect 195888 542846 195940 542852
rect 195900 539988 195928 542846
rect 197924 539988 197952 544886
rect 200026 543688 200082 543697
rect 200026 543623 200082 543632
rect 200040 539988 200068 543623
rect 202156 543250 202184 557602
rect 202144 543244 202196 543250
rect 202144 543186 202196 543192
rect 202050 543144 202106 543153
rect 202050 543079 202106 543088
rect 202064 539988 202092 543079
rect 202800 543046 202828 558855
rect 203812 558210 203840 558855
rect 203800 558204 203852 558210
rect 203800 558146 203852 558152
rect 203812 557734 203840 558146
rect 203800 557728 203852 557734
rect 203800 557670 203852 557676
rect 204180 543182 204208 558855
rect 204902 558648 204958 558657
rect 204902 558583 204958 558592
rect 204916 557734 204944 558583
rect 204904 557728 204956 557734
rect 204904 557670 204956 557676
rect 204916 543386 204944 557670
rect 205560 543726 205588 558855
rect 206940 558278 206968 558855
rect 208504 558550 208532 558855
rect 209042 558648 209098 558657
rect 209042 558583 209098 558592
rect 208492 558544 208544 558550
rect 208492 558486 208544 558492
rect 206928 558272 206980 558278
rect 206928 558214 206980 558220
rect 206940 557802 206968 558214
rect 208504 557870 208532 558486
rect 208492 557864 208544 557870
rect 208492 557806 208544 557812
rect 209056 557802 209084 558583
rect 210620 558414 210648 558855
rect 210608 558408 210660 558414
rect 210608 558350 210660 558356
rect 206928 557796 206980 557802
rect 206928 557738 206980 557744
rect 209044 557796 209096 557802
rect 209044 557738 209096 557744
rect 207662 557696 207718 557705
rect 207662 557631 207718 557640
rect 207676 557598 207704 557631
rect 207664 557592 207716 557598
rect 206926 557560 206982 557569
rect 207664 557534 207716 557540
rect 208306 557560 208362 557569
rect 206926 557495 206982 557504
rect 206192 544740 206244 544746
rect 206192 544682 206244 544688
rect 205548 543720 205600 543726
rect 205548 543662 205600 543668
rect 204904 543380 204956 543386
rect 204904 543322 204956 543328
rect 204168 543176 204220 543182
rect 204168 543118 204220 543124
rect 202788 543040 202840 543046
rect 202788 542982 202840 542988
rect 204168 542972 204220 542978
rect 204168 542914 204220 542920
rect 204180 539988 204208 542914
rect 206204 539988 206232 544682
rect 206940 543658 206968 557495
rect 206928 543652 206980 543658
rect 206928 543594 206980 543600
rect 207676 543454 207704 557534
rect 208306 557495 208362 557504
rect 208320 543590 208348 557495
rect 208308 543584 208360 543590
rect 208308 543526 208360 543532
rect 209056 543522 209084 557738
rect 209686 557560 209742 557569
rect 209686 557495 209742 557504
rect 209700 543522 209728 557495
rect 210422 543552 210478 543561
rect 209044 543516 209096 543522
rect 209044 543458 209096 543464
rect 209688 543516 209740 543522
rect 210422 543487 210478 543496
rect 209688 543458 209740 543464
rect 207664 543448 207716 543454
rect 207664 543390 207716 543396
rect 208306 543416 208362 543425
rect 208306 543351 208362 543360
rect 208320 539988 208348 543351
rect 210436 539988 210464 543487
rect 210988 542978 211016 559943
rect 211802 558920 211858 558929
rect 211802 558855 211858 558864
rect 213182 558920 213238 558929
rect 213182 558855 213238 558864
rect 214010 558920 214066 558929
rect 214010 558855 214066 558864
rect 215298 558920 215354 558929
rect 215298 558855 215354 558864
rect 217506 558920 217562 558929
rect 217506 558855 217562 558864
rect 218794 558920 218850 558929
rect 218794 558855 218850 558864
rect 220082 558920 220138 558929
rect 220082 558855 220138 558864
rect 221094 558920 221150 558929
rect 221094 558855 221150 558864
rect 222198 558920 222254 558929
rect 222198 558855 222254 558864
rect 224498 558920 224554 558929
rect 224498 558855 224554 558864
rect 225878 558920 225934 558929
rect 225878 558855 225934 558864
rect 226154 558920 226210 558929
rect 226154 558855 226210 558864
rect 227166 558920 227222 558929
rect 227166 558855 227222 558864
rect 227626 558920 227682 558929
rect 227626 558855 227682 558864
rect 227994 558920 228050 558929
rect 227994 558855 228050 558864
rect 229006 558920 229062 558929
rect 229006 558855 229062 558864
rect 229466 558920 229522 558929
rect 229466 558855 229522 558864
rect 230386 558920 230442 558929
rect 230386 558855 230442 558864
rect 231766 558920 231822 558929
rect 231766 558855 231822 558864
rect 233054 558920 233110 558929
rect 233054 558855 233110 558864
rect 233238 558920 233294 558929
rect 233238 558855 233294 558864
rect 234526 558920 234582 558929
rect 234526 558855 234582 558864
rect 235906 558920 235962 558929
rect 235906 558855 235962 558864
rect 237286 558920 237342 558929
rect 237286 558855 237342 558864
rect 240046 558920 240102 558929
rect 240046 558855 240102 558864
rect 211816 558346 211844 558855
rect 213196 558482 213224 558855
rect 213184 558476 213236 558482
rect 213184 558418 213236 558424
rect 211160 558340 211212 558346
rect 211160 558282 211212 558288
rect 211804 558340 211856 558346
rect 211804 558282 211856 558288
rect 211066 557696 211122 557705
rect 211172 557666 211200 558282
rect 213196 558210 213224 558418
rect 213184 558204 213236 558210
rect 213184 558146 213236 558152
rect 214024 557734 214052 558855
rect 215312 558822 215340 558855
rect 215300 558816 215352 558822
rect 215300 558758 215352 558764
rect 215312 558278 215340 558758
rect 217520 558618 217548 558855
rect 217598 558784 217654 558793
rect 218808 558754 218836 558855
rect 217598 558719 217654 558728
rect 218796 558748 218848 558754
rect 217508 558612 217560 558618
rect 217508 558554 217560 558560
rect 215300 558272 215352 558278
rect 215300 558214 215352 558220
rect 215208 558136 215260 558142
rect 215208 558078 215260 558084
rect 215220 557734 215248 558078
rect 214012 557728 214064 557734
rect 214012 557670 214064 557676
rect 215208 557728 215260 557734
rect 215208 557670 215260 557676
rect 211066 557631 211122 557640
rect 211160 557660 211212 557666
rect 211080 543454 211108 557631
rect 211160 557602 211212 557608
rect 217520 557598 217548 558554
rect 217612 558550 217640 558719
rect 218796 558690 218848 558696
rect 217600 558544 217652 558550
rect 217600 558486 217652 558492
rect 218808 557802 218836 558690
rect 220096 558414 220124 558855
rect 220084 558408 220136 558414
rect 220084 558350 220136 558356
rect 221108 558346 221136 558855
rect 222212 558686 222240 558855
rect 224512 558822 224540 558855
rect 224500 558816 224552 558822
rect 223578 558784 223634 558793
rect 224500 558758 224552 558764
rect 223578 558719 223634 558728
rect 222200 558680 222252 558686
rect 222200 558622 222252 558628
rect 222212 558482 222240 558622
rect 222200 558476 222252 558482
rect 222200 558418 222252 558424
rect 221096 558340 221148 558346
rect 221096 558282 221148 558288
rect 223592 557938 223620 558719
rect 224512 558278 224540 558758
rect 225892 558618 225920 558855
rect 225880 558612 225932 558618
rect 225880 558554 225932 558560
rect 224500 558272 224552 558278
rect 224500 558214 224552 558220
rect 223580 557932 223632 557938
rect 223580 557874 223632 557880
rect 218796 557796 218848 557802
rect 218796 557738 218848 557744
rect 217966 557696 218022 557705
rect 217966 557631 218022 557640
rect 217508 557592 217560 557598
rect 212446 557560 212502 557569
rect 212446 557495 212502 557504
rect 213826 557560 213882 557569
rect 213826 557495 213882 557504
rect 215206 557560 215262 557569
rect 215206 557495 215262 557504
rect 216586 557560 216642 557569
rect 217508 557534 217560 557540
rect 217874 557560 217930 557569
rect 216586 557495 216642 557504
rect 217874 557495 217930 557504
rect 212460 545578 212488 557495
rect 212368 545550 212488 545578
rect 211068 543448 211120 543454
rect 211068 543390 211120 543396
rect 212368 543386 212396 545550
rect 212448 544604 212500 544610
rect 212448 544546 212500 544552
rect 212356 543380 212408 543386
rect 212356 543322 212408 543328
rect 210976 542972 211028 542978
rect 210976 542914 211028 542920
rect 212460 539988 212488 544546
rect 213840 543114 213868 557495
rect 215220 543318 215248 557495
rect 216600 545578 216628 557495
rect 216508 545550 216628 545578
rect 215208 543312 215260 543318
rect 215208 543254 215260 543260
rect 216508 543250 216536 545550
rect 216496 543244 216548 543250
rect 216496 543186 216548 543192
rect 216588 543176 216640 543182
rect 216588 543118 216640 543124
rect 213828 543108 213880 543114
rect 213828 543050 213880 543056
rect 214564 543040 214616 543046
rect 214564 542982 214616 542988
rect 214576 539988 214604 542982
rect 216600 539988 216628 543118
rect 217888 542570 217916 557495
rect 217980 543046 218008 557631
rect 219346 557560 219402 557569
rect 219346 557495 219402 557504
rect 220726 557560 220782 557569
rect 220726 557495 220782 557504
rect 222106 557560 222162 557569
rect 222106 557495 222162 557504
rect 223486 557560 223542 557569
rect 223486 557495 223542 557504
rect 224866 557560 224922 557569
rect 224866 557495 224922 557504
rect 218704 543720 218756 543726
rect 218704 543662 218756 543668
rect 217968 543040 218020 543046
rect 217968 542982 218020 542988
rect 217876 542564 217928 542570
rect 217876 542506 217928 542512
rect 218716 539988 218744 543662
rect 219360 542502 219388 557495
rect 220740 543794 220768 557495
rect 220728 543788 220780 543794
rect 220728 543730 220780 543736
rect 220544 543720 220596 543726
rect 220544 543662 220596 543668
rect 220556 542706 220584 543662
rect 220728 543652 220780 543658
rect 220728 543594 220780 543600
rect 220544 542700 220596 542706
rect 220544 542642 220596 542648
rect 219348 542496 219400 542502
rect 219348 542438 219400 542444
rect 220740 539988 220768 543594
rect 222120 542638 222148 557495
rect 222844 543584 222896 543590
rect 222844 543526 222896 543532
rect 222108 542632 222160 542638
rect 222108 542574 222160 542580
rect 222856 539988 222884 543526
rect 223500 542842 223528 557495
rect 224880 545306 224908 557495
rect 224696 545278 224908 545306
rect 223488 542836 223540 542842
rect 223488 542778 223540 542784
rect 224696 542774 224724 545278
rect 224868 543516 224920 543522
rect 224868 543458 224920 543464
rect 224684 542768 224736 542774
rect 224684 542710 224736 542716
rect 224880 539988 224908 543458
rect 226168 542978 226196 558855
rect 226246 558784 226302 558793
rect 226246 558719 226302 558728
rect 226156 542972 226208 542978
rect 226156 542914 226208 542920
rect 226260 542910 226288 558719
rect 227180 558550 227208 558855
rect 227168 558544 227220 558550
rect 227168 558486 227220 558492
rect 227640 543658 227668 558855
rect 228008 558754 228036 558855
rect 227996 558748 228048 558754
rect 227996 558690 228048 558696
rect 229020 543726 229048 558855
rect 229480 558414 229508 558855
rect 229468 558408 229520 558414
rect 229468 558350 229520 558356
rect 229008 543720 229060 543726
rect 229008 543662 229060 543668
rect 227628 543652 227680 543658
rect 227628 543594 227680 543600
rect 230400 543590 230428 558855
rect 230478 558376 230534 558385
rect 230478 558311 230480 558320
rect 230532 558311 230534 558320
rect 230480 558282 230532 558288
rect 230388 543584 230440 543590
rect 230388 543526 230440 543532
rect 231780 543522 231808 558855
rect 231858 558784 231914 558793
rect 231858 558719 231914 558728
rect 231872 558686 231900 558719
rect 231860 558680 231912 558686
rect 231860 558622 231912 558628
rect 231858 558512 231914 558521
rect 231858 558447 231914 558456
rect 231872 558074 231900 558447
rect 231860 558068 231912 558074
rect 231860 558010 231912 558016
rect 231768 543516 231820 543522
rect 231768 543458 231820 543464
rect 226984 543448 227036 543454
rect 226984 543390 227036 543396
rect 226248 542904 226300 542910
rect 226248 542846 226300 542852
rect 226996 539988 227024 543390
rect 233068 543386 233096 558855
rect 233146 558784 233202 558793
rect 233146 558719 233202 558728
rect 233160 543454 233188 558719
rect 233252 558278 233280 558855
rect 233240 558272 233292 558278
rect 233240 558214 233292 558220
rect 233148 543448 233200 543454
rect 233148 543390 233200 543396
rect 231124 543380 231176 543386
rect 231124 543322 231176 543328
rect 233056 543380 233108 543386
rect 233056 543322 233108 543328
rect 229100 543244 229152 543250
rect 229100 543186 229152 543192
rect 229112 539988 229140 543186
rect 231136 539988 231164 543322
rect 234540 543250 234568 558855
rect 234618 558784 234674 558793
rect 234618 558719 234674 558728
rect 234632 558618 234660 558719
rect 234620 558612 234672 558618
rect 234620 558554 234672 558560
rect 235920 543318 235948 558855
rect 235998 558784 236054 558793
rect 235998 558719 236054 558728
rect 236012 558550 236040 558719
rect 236000 558544 236052 558550
rect 236000 558486 236052 558492
rect 235264 543312 235316 543318
rect 235264 543254 235316 543260
rect 235908 543312 235960 543318
rect 235908 543254 235960 543260
rect 234528 543244 234580 543250
rect 234528 543186 234580 543192
rect 233240 543108 233292 543114
rect 233240 543050 233292 543056
rect 233252 539988 233280 543050
rect 235276 539988 235304 543254
rect 237300 543114 237328 558855
rect 237378 558784 237434 558793
rect 237378 558719 237380 558728
rect 237432 558719 237434 558728
rect 237380 558690 237432 558696
rect 238758 558376 238814 558385
rect 238758 558311 238814 558320
rect 238772 558278 238800 558311
rect 238760 558272 238812 558278
rect 238760 558214 238812 558220
rect 238666 558104 238722 558113
rect 238666 558039 238722 558048
rect 238680 543182 238708 558039
rect 237380 543176 237432 543182
rect 237380 543118 237432 543124
rect 238668 543176 238720 543182
rect 238668 543118 238720 543124
rect 237288 543108 237340 543114
rect 237288 543050 237340 543056
rect 237392 539988 237420 543118
rect 240060 543046 240088 558855
rect 260196 543720 260248 543726
rect 260196 543662 260248 543668
rect 258080 543652 258132 543658
rect 258080 543594 258132 543600
rect 239404 543040 239456 543046
rect 239404 542982 239456 542988
rect 240048 543040 240100 543046
rect 240048 542982 240100 542988
rect 239416 539988 239444 542982
rect 256056 542972 256108 542978
rect 256056 542914 256108 542920
rect 253940 542904 253992 542910
rect 253940 542846 253992 542852
rect 249800 542836 249852 542842
rect 249800 542778 249852 542784
rect 245660 542700 245712 542706
rect 245660 542642 245712 542648
rect 241520 542564 241572 542570
rect 241520 542506 241572 542512
rect 241532 539988 241560 542506
rect 243544 542496 243596 542502
rect 243544 542438 243596 542444
rect 243556 539988 243584 542438
rect 245672 539988 245700 542642
rect 247776 542632 247828 542638
rect 247776 542574 247828 542580
rect 247788 539988 247816 542574
rect 249812 539988 249840 542778
rect 251916 542768 251968 542774
rect 251916 542710 251968 542716
rect 251928 539988 251956 542710
rect 253952 539988 253980 542846
rect 256068 539988 256096 542914
rect 258092 539988 258120 543594
rect 260208 539988 260236 543662
rect 262220 543584 262272 543590
rect 262220 543526 262272 543532
rect 262232 539988 262260 543526
rect 264336 543516 264388 543522
rect 264336 543458 264388 543464
rect 264348 539988 264376 543458
rect 266452 543448 266504 543454
rect 266452 543390 266504 543396
rect 266464 539988 266492 543390
rect 268476 543380 268528 543386
rect 268476 543322 268528 543328
rect 268488 539988 268516 543322
rect 272616 543312 272668 543318
rect 272616 543254 272668 543260
rect 270592 543244 270644 543250
rect 270592 543186 270644 543192
rect 270604 539988 270632 543186
rect 272628 539988 272656 543254
rect 276756 543176 276808 543182
rect 276756 543118 276808 543124
rect 274732 543108 274784 543114
rect 274732 543050 274784 543056
rect 274744 539988 274772 543050
rect 276768 539988 276796 543118
rect 278872 543040 278924 543046
rect 278872 542982 278924 542988
rect 278884 539988 278912 542982
rect 279160 320906 279188 580246
rect 281538 579048 281594 579057
rect 281538 578983 281594 578992
rect 281446 441008 281502 441017
rect 281446 440943 281502 440952
rect 281460 440298 281488 440943
rect 281448 440292 281500 440298
rect 281448 440234 281500 440240
rect 281446 429992 281502 430001
rect 281446 429927 281502 429936
rect 281460 429214 281488 429927
rect 281448 429208 281500 429214
rect 281448 429150 281500 429156
rect 281552 329882 281580 578983
rect 282274 539472 282330 539481
rect 282274 539407 282330 539416
rect 282288 538354 282316 539407
rect 282826 538520 282882 538529
rect 282826 538455 282882 538464
rect 282276 538348 282328 538354
rect 282276 538290 282328 538296
rect 282840 538286 282868 538455
rect 282828 538280 282880 538286
rect 282828 538222 282880 538228
rect 282826 537432 282882 537441
rect 282826 537367 282882 537376
rect 282840 536858 282868 537367
rect 282828 536852 282880 536858
rect 282828 536794 282880 536800
rect 282826 536480 282882 536489
rect 282826 536415 282882 536424
rect 282840 535498 282868 536415
rect 282828 535492 282880 535498
rect 282828 535434 282880 535440
rect 281722 535392 281778 535401
rect 281722 535327 281778 535336
rect 281736 534206 281764 535327
rect 282090 534440 282146 534449
rect 282090 534375 282146 534384
rect 281724 534200 281776 534206
rect 281724 534142 281776 534148
rect 282104 534138 282132 534375
rect 282092 534132 282144 534138
rect 282092 534074 282144 534080
rect 282090 533488 282146 533497
rect 282090 533423 282146 533432
rect 282104 532778 282132 533423
rect 282092 532772 282144 532778
rect 282092 532714 282144 532720
rect 282274 532400 282330 532409
rect 282274 532335 282330 532344
rect 282288 531418 282316 532335
rect 282826 531448 282882 531457
rect 282276 531412 282328 531418
rect 282826 531383 282882 531392
rect 282276 531354 282328 531360
rect 282840 531350 282868 531383
rect 282828 531344 282880 531350
rect 282828 531286 282880 531292
rect 282826 530360 282882 530369
rect 282826 530295 282882 530304
rect 282840 529990 282868 530295
rect 282828 529984 282880 529990
rect 282828 529926 282880 529932
rect 282826 529408 282882 529417
rect 282826 529343 282882 529352
rect 282840 528630 282868 529343
rect 282828 528624 282880 528630
rect 282828 528566 282880 528572
rect 282274 528320 282330 528329
rect 282274 528255 282330 528264
rect 282288 527202 282316 528255
rect 282826 527368 282882 527377
rect 282826 527303 282882 527312
rect 282840 527270 282868 527303
rect 282828 527264 282880 527270
rect 282828 527206 282880 527212
rect 282276 527196 282328 527202
rect 282276 527138 282328 527144
rect 281906 526416 281962 526425
rect 281906 526351 281962 526360
rect 281920 525842 281948 526351
rect 281908 525836 281960 525842
rect 281908 525778 281960 525784
rect 282826 525328 282882 525337
rect 282826 525263 282882 525272
rect 282840 524482 282868 525263
rect 282828 524476 282880 524482
rect 282828 524418 282880 524424
rect 282366 524376 282422 524385
rect 282366 524311 282422 524320
rect 282380 523054 282408 524311
rect 282826 523288 282882 523297
rect 282826 523223 282882 523232
rect 282840 523122 282868 523223
rect 282828 523116 282880 523122
rect 282828 523058 282880 523064
rect 282368 523048 282420 523054
rect 282368 522990 282420 522996
rect 282826 522336 282882 522345
rect 282826 522271 282882 522280
rect 282840 521694 282868 522271
rect 282828 521688 282880 521694
rect 282828 521630 282880 521636
rect 283562 521248 283618 521257
rect 283562 521183 283618 521192
rect 282828 520328 282880 520334
rect 282826 520296 282828 520305
rect 282880 520296 282882 520305
rect 282826 520231 282882 520240
rect 281722 519344 281778 519353
rect 281722 519279 281778 519288
rect 281736 519110 281764 519279
rect 281724 519104 281776 519110
rect 281724 519046 281776 519052
rect 282090 518256 282146 518265
rect 282090 518191 282146 518200
rect 282104 517546 282132 518191
rect 282092 517540 282144 517546
rect 282092 517482 282144 517488
rect 282274 517304 282330 517313
rect 282274 517239 282330 517248
rect 282288 516254 282316 517239
rect 282276 516248 282328 516254
rect 282276 516190 282328 516196
rect 282826 516216 282882 516225
rect 282826 516151 282828 516160
rect 282880 516151 282882 516160
rect 282828 516122 282880 516128
rect 282826 515264 282882 515273
rect 282826 515199 282882 515208
rect 282840 514826 282868 515199
rect 282828 514820 282880 514826
rect 282828 514762 282880 514768
rect 282274 514312 282330 514321
rect 282274 514247 282330 514256
rect 282288 513398 282316 514247
rect 282276 513392 282328 513398
rect 282276 513334 282328 513340
rect 282734 513224 282790 513233
rect 282734 513159 282790 513168
rect 282748 512106 282776 513159
rect 282826 512272 282882 512281
rect 282826 512207 282882 512216
rect 282736 512100 282788 512106
rect 282736 512042 282788 512048
rect 282840 512038 282868 512207
rect 282828 512032 282880 512038
rect 282828 511974 282880 511980
rect 281722 511184 281778 511193
rect 281722 511119 281778 511128
rect 281736 510678 281764 511119
rect 281724 510672 281776 510678
rect 281724 510614 281776 510620
rect 282274 510232 282330 510241
rect 282274 510167 282330 510176
rect 282288 509318 282316 510167
rect 282276 509312 282328 509318
rect 282276 509254 282328 509260
rect 282550 509144 282606 509153
rect 282550 509079 282606 509088
rect 282564 507958 282592 509079
rect 282826 508192 282882 508201
rect 282826 508127 282882 508136
rect 282552 507952 282604 507958
rect 282552 507894 282604 507900
rect 282840 507890 282868 508127
rect 282828 507884 282880 507890
rect 282828 507826 282880 507832
rect 282090 507240 282146 507249
rect 282090 507175 282146 507184
rect 282104 506530 282132 507175
rect 282092 506524 282144 506530
rect 282092 506466 282144 506472
rect 282734 506152 282790 506161
rect 282734 506087 282790 506096
rect 282748 505170 282776 506087
rect 282828 505232 282880 505238
rect 282826 505200 282828 505209
rect 282880 505200 282882 505209
rect 282736 505164 282788 505170
rect 282826 505135 282882 505144
rect 282736 505106 282788 505112
rect 282826 504112 282882 504121
rect 282826 504047 282882 504056
rect 282840 503742 282868 504047
rect 282828 503736 282880 503742
rect 282828 503678 282880 503684
rect 282826 503160 282882 503169
rect 282826 503095 282882 503104
rect 282840 502382 282868 503095
rect 282828 502376 282880 502382
rect 282828 502318 282880 502324
rect 282274 502072 282330 502081
rect 282274 502007 282330 502016
rect 282288 501022 282316 502007
rect 282826 501120 282882 501129
rect 282826 501055 282828 501064
rect 282880 501055 282882 501064
rect 282828 501026 282880 501032
rect 282276 501016 282328 501022
rect 282276 500958 282328 500964
rect 282826 499080 282882 499089
rect 282826 499015 282882 499024
rect 282840 498234 282868 499015
rect 282828 498228 282880 498234
rect 282828 498170 282880 498176
rect 282826 497040 282882 497049
rect 282826 496975 282882 496984
rect 282840 496874 282868 496975
rect 282828 496868 282880 496874
rect 282828 496810 282880 496816
rect 281906 496088 281962 496097
rect 281906 496023 281962 496032
rect 281920 495514 281948 496023
rect 281908 495508 281960 495514
rect 281908 495450 281960 495456
rect 282826 495136 282882 495145
rect 282826 495071 282882 495080
rect 282840 494086 282868 495071
rect 282828 494080 282880 494086
rect 282366 494048 282422 494057
rect 282828 494022 282880 494028
rect 282366 493983 282422 493992
rect 282380 492726 282408 493983
rect 282826 493096 282882 493105
rect 282826 493031 282882 493040
rect 282840 492794 282868 493031
rect 282828 492788 282880 492794
rect 282828 492730 282880 492736
rect 282368 492720 282420 492726
rect 282368 492662 282420 492668
rect 282826 492008 282882 492017
rect 282826 491943 282882 491952
rect 282840 491366 282868 491943
rect 282828 491360 282880 491366
rect 282828 491302 282880 491308
rect 282274 491056 282330 491065
rect 282274 490991 282330 491000
rect 282288 489938 282316 490991
rect 282828 490000 282880 490006
rect 282826 489968 282828 489977
rect 282880 489968 282882 489977
rect 282276 489932 282328 489938
rect 282826 489903 282882 489912
rect 282276 489874 282328 489880
rect 282274 489016 282330 489025
rect 282274 488951 282330 488960
rect 282288 488578 282316 488951
rect 282276 488572 282328 488578
rect 282276 488514 282328 488520
rect 282826 488064 282882 488073
rect 282826 487999 282882 488008
rect 282840 487218 282868 487999
rect 282828 487212 282880 487218
rect 282828 487154 282880 487160
rect 282274 486976 282330 486985
rect 282274 486911 282330 486920
rect 282288 485858 282316 486911
rect 282826 486024 282882 486033
rect 282826 485959 282882 485968
rect 282840 485926 282868 485959
rect 282828 485920 282880 485926
rect 282828 485862 282880 485868
rect 282276 485852 282328 485858
rect 282276 485794 282328 485800
rect 281722 484936 281778 484945
rect 281722 484871 281778 484880
rect 281736 484430 281764 484871
rect 281724 484424 281776 484430
rect 281724 484366 281776 484372
rect 282274 483984 282330 483993
rect 282274 483919 282330 483928
rect 282288 483070 282316 483919
rect 282276 483064 282328 483070
rect 282276 483006 282328 483012
rect 282550 482896 282606 482905
rect 282550 482831 282606 482840
rect 282564 481710 282592 482831
rect 282826 481944 282882 481953
rect 282826 481879 282882 481888
rect 282840 481778 282868 481879
rect 282828 481772 282880 481778
rect 282828 481714 282880 481720
rect 282552 481704 282604 481710
rect 282552 481646 282604 481652
rect 282090 480992 282146 481001
rect 282090 480927 282146 480936
rect 282104 480282 282132 480927
rect 282092 480276 282144 480282
rect 282092 480218 282144 480224
rect 282734 479904 282790 479913
rect 282734 479839 282790 479848
rect 282748 478922 282776 479839
rect 282828 478984 282880 478990
rect 282826 478952 282828 478961
rect 282880 478952 282882 478961
rect 282736 478916 282788 478922
rect 282826 478887 282882 478896
rect 282736 478858 282788 478864
rect 282826 477864 282882 477873
rect 282826 477799 282882 477808
rect 282840 477562 282868 477799
rect 282828 477556 282880 477562
rect 282828 477498 282880 477504
rect 282090 476912 282146 476921
rect 282090 476847 282146 476856
rect 282104 476134 282132 476847
rect 282092 476128 282144 476134
rect 282092 476070 282144 476076
rect 282274 475824 282330 475833
rect 282274 475759 282330 475768
rect 282288 474774 282316 475759
rect 282826 474872 282882 474881
rect 282826 474807 282828 474816
rect 282880 474807 282882 474816
rect 282828 474778 282880 474784
rect 282276 474768 282328 474774
rect 282276 474710 282328 474716
rect 281722 473920 281778 473929
rect 281722 473855 281778 473864
rect 281736 473414 281764 473855
rect 281724 473408 281776 473414
rect 281724 473350 281776 473356
rect 282090 472832 282146 472841
rect 282090 472767 282146 472776
rect 282104 472054 282132 472767
rect 282092 472048 282144 472054
rect 282092 471990 282144 471996
rect 282734 471880 282790 471889
rect 282734 471815 282790 471824
rect 282748 470626 282776 471815
rect 282826 470792 282882 470801
rect 282826 470727 282882 470736
rect 282840 470694 282868 470727
rect 282828 470688 282880 470694
rect 282828 470630 282880 470636
rect 282736 470620 282788 470626
rect 282736 470562 282788 470568
rect 281906 469840 281962 469849
rect 281906 469775 281962 469784
rect 281920 469266 281948 469775
rect 281908 469260 281960 469266
rect 281908 469202 281960 469208
rect 282826 468888 282882 468897
rect 282826 468823 282882 468832
rect 282840 467906 282868 468823
rect 282828 467900 282880 467906
rect 282828 467842 282880 467848
rect 282734 467800 282790 467809
rect 282734 467735 282790 467744
rect 282748 466546 282776 467735
rect 282826 466848 282882 466857
rect 282826 466783 282882 466792
rect 282736 466540 282788 466546
rect 282736 466482 282788 466488
rect 282840 466478 282868 466783
rect 282828 466472 282880 466478
rect 282828 466414 282880 466420
rect 282826 465760 282882 465769
rect 282826 465695 282882 465704
rect 282840 465118 282868 465695
rect 282828 465112 282880 465118
rect 282828 465054 282880 465060
rect 282734 464808 282790 464817
rect 282734 464743 282790 464752
rect 282748 463826 282776 464743
rect 282736 463820 282788 463826
rect 282736 463762 282788 463768
rect 282828 463752 282880 463758
rect 282826 463720 282828 463729
rect 282880 463720 282882 463729
rect 282826 463655 282882 463664
rect 282826 462768 282882 462777
rect 282826 462703 282882 462712
rect 282840 462398 282868 462703
rect 282828 462392 282880 462398
rect 282828 462334 282880 462340
rect 282826 461816 282882 461825
rect 282826 461751 282882 461760
rect 282840 460970 282868 461751
rect 282828 460964 282880 460970
rect 282828 460906 282880 460912
rect 282826 460728 282882 460737
rect 282826 460663 282882 460672
rect 282734 459776 282790 459785
rect 282734 459711 282790 459720
rect 282748 459678 282776 459711
rect 282736 459672 282788 459678
rect 282736 459614 282788 459620
rect 282840 459610 282868 460663
rect 282828 459604 282880 459610
rect 282828 459546 282880 459552
rect 281722 458688 281778 458697
rect 281722 458623 281778 458632
rect 281736 458250 281764 458623
rect 281724 458244 281776 458250
rect 281724 458186 281776 458192
rect 282090 457736 282146 457745
rect 282090 457671 282146 457680
rect 282104 456822 282132 457671
rect 282092 456816 282144 456822
rect 282092 456758 282144 456764
rect 281630 456648 281686 456657
rect 281630 456583 281686 456592
rect 281644 455530 281672 456583
rect 282826 455696 282882 455705
rect 282826 455631 282882 455640
rect 281632 455524 281684 455530
rect 281632 455466 281684 455472
rect 282840 455462 282868 455631
rect 282828 455456 282880 455462
rect 282828 455398 282880 455404
rect 281630 454744 281686 454753
rect 281630 454679 281686 454688
rect 281644 421394 281672 454679
rect 282458 453656 282514 453665
rect 282458 453591 282514 453600
rect 282274 452704 282330 452713
rect 282274 452639 282330 452648
rect 282090 446584 282146 446593
rect 282090 446519 282146 446528
rect 281814 445632 281870 445641
rect 281814 445567 281870 445576
rect 281722 442640 281778 442649
rect 281722 442575 281778 442584
rect 281632 421388 281684 421394
rect 281632 421330 281684 421336
rect 281632 421252 281684 421258
rect 281632 421194 281684 421200
rect 281644 413098 281672 421194
rect 281736 413846 281764 442575
rect 281724 413840 281776 413846
rect 281724 413782 281776 413788
rect 281828 413642 281856 445567
rect 281998 444544 282054 444553
rect 281998 444479 282054 444488
rect 281906 443592 281962 443601
rect 281906 443527 281962 443536
rect 281920 413778 281948 443527
rect 281908 413772 281960 413778
rect 281908 413714 281960 413720
rect 282012 413710 282040 444479
rect 282000 413704 282052 413710
rect 282000 413646 282052 413652
rect 281816 413636 281868 413642
rect 281816 413578 281868 413584
rect 282104 413574 282132 446519
rect 282182 440600 282238 440609
rect 282182 440535 282238 440544
rect 282196 440434 282224 440535
rect 282184 440428 282236 440434
rect 282184 440370 282236 440376
rect 282182 439512 282238 439521
rect 282182 439447 282238 439456
rect 282196 438938 282224 439447
rect 282184 438932 282236 438938
rect 282184 438874 282236 438880
rect 282182 437472 282238 437481
rect 282182 437407 282238 437416
rect 282196 436626 282224 437407
rect 282184 436620 282236 436626
rect 282184 436562 282236 436568
rect 282182 436520 282238 436529
rect 282182 436455 282238 436464
rect 282196 436218 282224 436455
rect 282184 436212 282236 436218
rect 282184 436154 282236 436160
rect 282182 435568 282238 435577
rect 282182 435503 282238 435512
rect 282196 434790 282224 435503
rect 282184 434784 282236 434790
rect 282184 434726 282236 434732
rect 282182 434480 282238 434489
rect 282182 434415 282238 434424
rect 282196 433362 282224 434415
rect 282184 433356 282236 433362
rect 282184 433298 282236 433304
rect 282182 432440 282238 432449
rect 282182 432375 282238 432384
rect 282196 413982 282224 432375
rect 282288 431594 282316 452639
rect 282366 451616 282422 451625
rect 282366 451551 282422 451560
rect 282276 431588 282328 431594
rect 282276 431530 282328 431536
rect 282274 431488 282330 431497
rect 282274 431423 282330 431432
rect 282288 430710 282316 431423
rect 282276 430704 282328 430710
rect 282276 430646 282328 430652
rect 282276 430568 282328 430574
rect 282276 430510 282328 430516
rect 282288 429457 282316 430510
rect 282274 429448 282330 429457
rect 282274 429383 282330 429392
rect 282276 429140 282328 429146
rect 282276 429082 282328 429088
rect 282288 428505 282316 429082
rect 282274 428496 282330 428505
rect 282274 428431 282330 428440
rect 282276 427780 282328 427786
rect 282276 427722 282328 427728
rect 282288 427417 282316 427722
rect 282274 427408 282330 427417
rect 282274 427343 282330 427352
rect 282276 427236 282328 427242
rect 282276 427178 282328 427184
rect 282288 427009 282316 427178
rect 282274 427000 282330 427009
rect 282274 426935 282330 426944
rect 282276 426420 282328 426426
rect 282276 426362 282328 426368
rect 282288 425377 282316 426362
rect 282274 425368 282330 425377
rect 282274 425303 282330 425312
rect 282276 425060 282328 425066
rect 282276 425002 282328 425008
rect 282288 424425 282316 425002
rect 282274 424416 282330 424425
rect 282274 424351 282330 424360
rect 282276 423632 282328 423638
rect 282276 423574 282328 423580
rect 282288 423473 282316 423574
rect 282274 423464 282330 423473
rect 282274 423399 282330 423408
rect 282276 423292 282328 423298
rect 282276 423234 282328 423240
rect 282288 422385 282316 423234
rect 282274 422376 282330 422385
rect 282274 422311 282330 422320
rect 282276 422272 282328 422278
rect 282276 422214 282328 422220
rect 282288 421433 282316 422214
rect 282274 421424 282330 421433
rect 282274 421359 282330 421368
rect 282380 421274 282408 451551
rect 282288 421246 282408 421274
rect 282472 421258 282500 453591
rect 282550 450664 282606 450673
rect 282550 450599 282606 450608
rect 282460 421252 282512 421258
rect 282288 417790 282316 421246
rect 282460 421194 282512 421200
rect 282564 421138 282592 450599
rect 282826 449712 282882 449721
rect 282826 449647 282882 449656
rect 282642 448624 282698 448633
rect 282642 448559 282698 448568
rect 282380 421110 282592 421138
rect 282276 417784 282328 417790
rect 282276 417726 282328 417732
rect 282276 417648 282328 417654
rect 282276 417590 282328 417596
rect 282288 415478 282316 417590
rect 282276 415472 282328 415478
rect 282276 415414 282328 415420
rect 282276 415336 282328 415342
rect 282276 415278 282328 415284
rect 282288 414361 282316 415278
rect 282274 414352 282330 414361
rect 282274 414287 282330 414296
rect 282184 413976 282236 413982
rect 282184 413918 282236 413924
rect 282276 413908 282328 413914
rect 282276 413850 282328 413856
rect 282092 413568 282144 413574
rect 282092 413510 282144 413516
rect 281632 413092 281684 413098
rect 281632 413034 281684 413040
rect 282288 413030 282316 413850
rect 282380 413370 282408 421110
rect 282460 421048 282512 421054
rect 282460 420990 282512 420996
rect 282368 413364 282420 413370
rect 282368 413306 282420 413312
rect 282472 413302 282500 420990
rect 282552 419484 282604 419490
rect 282552 419426 282604 419432
rect 282564 418305 282592 419426
rect 282550 418296 282606 418305
rect 282550 418231 282606 418240
rect 282552 417784 282604 417790
rect 282552 417726 282604 417732
rect 282460 413296 282512 413302
rect 282460 413238 282512 413244
rect 282564 413234 282592 417726
rect 282656 413438 282684 448559
rect 282734 447672 282790 447681
rect 282734 447607 282790 447616
rect 282748 413506 282776 447607
rect 282840 421054 282868 449647
rect 283470 438560 283526 438569
rect 283470 438495 283526 438504
rect 283378 433528 283434 433537
rect 283378 433463 283434 433472
rect 282828 421048 282880 421054
rect 282828 420990 282880 420996
rect 282828 420912 282880 420918
rect 282828 420854 282880 420860
rect 282840 420345 282868 420854
rect 282826 420336 282882 420345
rect 282826 420271 282882 420280
rect 282828 419416 282880 419422
rect 282826 419384 282828 419393
rect 282880 419384 282882 419393
rect 282826 419319 282882 419328
rect 282828 418124 282880 418130
rect 282828 418066 282880 418072
rect 282840 417353 282868 418066
rect 282826 417344 282882 417353
rect 282826 417279 282882 417288
rect 282828 416764 282880 416770
rect 282828 416706 282880 416712
rect 282840 416401 282868 416706
rect 282826 416392 282882 416401
rect 282826 416327 282882 416336
rect 283288 416220 283340 416226
rect 283288 416162 283340 416168
rect 283196 416152 283248 416158
rect 283196 416094 283248 416100
rect 283104 416084 283156 416090
rect 283104 416026 283156 416032
rect 282920 415472 282972 415478
rect 282920 415414 282972 415420
rect 282828 415404 282880 415410
rect 282828 415346 282880 415352
rect 282840 415313 282868 415346
rect 282826 415304 282882 415313
rect 282826 415239 282882 415248
rect 282932 415154 282960 415414
rect 282840 415126 282960 415154
rect 282736 413500 282788 413506
rect 282736 413442 282788 413448
rect 282644 413432 282696 413438
rect 282840 413386 282868 415126
rect 283012 414792 283064 414798
rect 283012 414734 283064 414740
rect 282920 414724 282972 414730
rect 282920 414666 282972 414672
rect 282644 413374 282696 413380
rect 282748 413358 282868 413386
rect 282552 413228 282604 413234
rect 282552 413170 282604 413176
rect 282748 413166 282776 413358
rect 282826 413264 282882 413273
rect 282932 413250 282960 414666
rect 282882 413222 282960 413250
rect 282826 413199 282882 413208
rect 282736 413160 282788 413166
rect 282736 413102 282788 413108
rect 282276 413024 282328 413030
rect 282276 412966 282328 412972
rect 282826 412312 282882 412321
rect 282826 412247 282882 412256
rect 282840 412162 282868 412247
rect 283024 412162 283052 414734
rect 282840 412134 283052 412162
rect 282736 411256 282788 411262
rect 282736 411198 282788 411204
rect 282826 411224 282882 411233
rect 281632 411120 281684 411126
rect 281632 411062 281684 411068
rect 281644 406994 281672 411062
rect 282000 411052 282052 411058
rect 282000 410994 282052 411000
rect 281724 409828 281776 409834
rect 281724 409770 281776 409776
rect 281736 409329 281764 409770
rect 281722 409320 281778 409329
rect 281722 409255 281778 409264
rect 281724 408468 281776 408474
rect 281724 408410 281776 408416
rect 281736 408241 281764 408410
rect 281722 408232 281778 408241
rect 281722 408167 281778 408176
rect 281644 406966 281764 406994
rect 281632 404048 281684 404054
rect 281632 403990 281684 403996
rect 281644 403209 281672 403990
rect 281630 403200 281686 403209
rect 281630 403135 281686 403144
rect 281632 398200 281684 398206
rect 281630 398168 281632 398177
rect 281684 398168 281686 398177
rect 281630 398103 281686 398112
rect 281632 397248 281684 397254
rect 281630 397216 281632 397225
rect 281684 397216 281686 397225
rect 281630 397151 281686 397160
rect 281632 396500 281684 396506
rect 281632 396442 281684 396448
rect 281644 396137 281672 396442
rect 281630 396128 281686 396137
rect 281630 396063 281686 396072
rect 281632 395820 281684 395826
rect 281632 395762 281684 395768
rect 281644 395185 281672 395762
rect 281630 395176 281686 395185
rect 281630 395111 281686 395120
rect 281632 394392 281684 394398
rect 281632 394334 281684 394340
rect 281644 394097 281672 394334
rect 281630 394088 281686 394097
rect 281630 394023 281686 394032
rect 281632 393236 281684 393242
rect 281632 393178 281684 393184
rect 281644 393145 281672 393178
rect 281630 393136 281686 393145
rect 281630 393071 281686 393080
rect 281632 392080 281684 392086
rect 281630 392048 281632 392057
rect 281684 392048 281686 392057
rect 281630 391983 281686 391992
rect 281632 391672 281684 391678
rect 281632 391614 281684 391620
rect 281644 391105 281672 391614
rect 281630 391096 281686 391105
rect 281630 391031 281686 391040
rect 281632 390176 281684 390182
rect 281630 390144 281632 390153
rect 281684 390144 281686 390153
rect 281630 390079 281686 390088
rect 281632 389088 281684 389094
rect 281630 389056 281632 389065
rect 281684 389056 281686 389065
rect 281630 388991 281686 389000
rect 281632 388340 281684 388346
rect 281632 388282 281684 388288
rect 281644 388113 281672 388282
rect 281630 388104 281686 388113
rect 281630 388039 281686 388048
rect 281632 387116 281684 387122
rect 281632 387058 281684 387064
rect 281644 387025 281672 387058
rect 281630 387016 281686 387025
rect 281630 386951 281686 386960
rect 281632 386096 281684 386102
rect 281630 386064 281632 386073
rect 281684 386064 281686 386073
rect 281630 385999 281686 386008
rect 281632 385280 281684 385286
rect 281632 385222 281684 385228
rect 281644 385121 281672 385222
rect 281630 385112 281686 385121
rect 281630 385047 281686 385056
rect 281632 384056 281684 384062
rect 281630 384024 281632 384033
rect 281684 384024 281686 384033
rect 281630 383959 281686 383968
rect 281632 383308 281684 383314
rect 281632 383250 281684 383256
rect 281644 383081 281672 383250
rect 281630 383072 281686 383081
rect 281630 383007 281686 383016
rect 281632 382152 281684 382158
rect 281632 382094 281684 382100
rect 281644 381993 281672 382094
rect 281630 381984 281686 381993
rect 281630 381919 281686 381928
rect 281632 380860 281684 380866
rect 281632 380802 281684 380808
rect 281644 379953 281672 380802
rect 281630 379944 281686 379953
rect 281630 379879 281686 379888
rect 281632 379500 281684 379506
rect 281632 379442 281684 379448
rect 281644 379001 281672 379442
rect 281630 378992 281686 379001
rect 281630 378927 281686 378936
rect 281632 378140 281684 378146
rect 281632 378082 281684 378088
rect 281644 378049 281672 378082
rect 281630 378040 281686 378049
rect 281630 377975 281686 377984
rect 281632 376712 281684 376718
rect 281632 376654 281684 376660
rect 281644 376009 281672 376654
rect 281630 376000 281686 376009
rect 281630 375935 281686 375944
rect 281632 375352 281684 375358
rect 281632 375294 281684 375300
rect 281644 374921 281672 375294
rect 281630 374912 281686 374921
rect 281630 374847 281686 374856
rect 281630 373960 281686 373969
rect 281630 373895 281686 373904
rect 281644 373182 281672 373895
rect 281632 373176 281684 373182
rect 281632 373118 281684 373124
rect 281632 371952 281684 371958
rect 281630 371920 281632 371929
rect 281684 371920 281686 371929
rect 281630 371855 281686 371864
rect 281632 371000 281684 371006
rect 281630 370968 281632 370977
rect 281684 370968 281686 370977
rect 281630 370903 281686 370912
rect 281632 369844 281684 369850
rect 281632 369786 281684 369792
rect 281644 368937 281672 369786
rect 281630 368928 281686 368937
rect 281630 368863 281686 368872
rect 281632 368484 281684 368490
rect 281632 368426 281684 368432
rect 281644 367849 281672 368426
rect 281630 367840 281686 367849
rect 281630 367775 281686 367784
rect 281632 365696 281684 365702
rect 281632 365638 281684 365644
rect 281644 364857 281672 365638
rect 281630 364848 281686 364857
rect 281630 364783 281686 364792
rect 281632 364336 281684 364342
rect 281632 364278 281684 364284
rect 281644 363905 281672 364278
rect 281630 363896 281686 363905
rect 281630 363831 281686 363840
rect 281632 362908 281684 362914
rect 281632 362850 281684 362856
rect 281644 362817 281672 362850
rect 281630 362808 281686 362817
rect 281630 362743 281686 362752
rect 281632 361548 281684 361554
rect 281632 361490 281684 361496
rect 281644 360777 281672 361490
rect 281630 360768 281686 360777
rect 281630 360703 281686 360712
rect 281632 360188 281684 360194
rect 281632 360130 281684 360136
rect 281644 359825 281672 360130
rect 281630 359816 281686 359825
rect 281630 359751 281686 359760
rect 281632 358760 281684 358766
rect 281632 358702 281684 358708
rect 281644 357785 281672 358702
rect 281630 357776 281686 357785
rect 281630 357711 281686 357720
rect 281632 351824 281684 351830
rect 281630 351792 281632 351801
rect 281684 351792 281686 351801
rect 281630 351727 281686 351736
rect 281632 350940 281684 350946
rect 281632 350882 281684 350888
rect 281644 350713 281672 350882
rect 281630 350704 281686 350713
rect 281630 350639 281686 350648
rect 281632 350328 281684 350334
rect 281632 350270 281684 350276
rect 281644 349761 281672 350270
rect 281630 349752 281686 349761
rect 281630 349687 281686 349696
rect 281632 349104 281684 349110
rect 281632 349046 281684 349052
rect 281644 348673 281672 349046
rect 281630 348664 281686 348673
rect 281630 348599 281686 348608
rect 281632 347744 281684 347750
rect 281630 347712 281632 347721
rect 281684 347712 281686 347721
rect 281630 347647 281686 347656
rect 281632 346792 281684 346798
rect 281632 346734 281684 346740
rect 281644 346633 281672 346734
rect 281630 346624 281686 346633
rect 281630 346559 281686 346568
rect 281632 345704 281684 345710
rect 281630 345672 281632 345681
rect 281684 345672 281686 345681
rect 281630 345607 281686 345616
rect 281632 344888 281684 344894
rect 281632 344830 281684 344836
rect 281644 344729 281672 344830
rect 281630 344720 281686 344729
rect 281630 344655 281686 344664
rect 281630 343632 281686 343641
rect 281630 343567 281632 343576
rect 281684 343567 281686 343576
rect 281632 343538 281684 343544
rect 281632 342236 281684 342242
rect 281632 342178 281684 342184
rect 281644 341601 281672 342178
rect 281630 341592 281686 341601
rect 281630 341527 281686 341536
rect 281632 340808 281684 340814
rect 281632 340750 281684 340756
rect 281736 340762 281764 406966
rect 282012 405770 282040 410994
rect 282184 410984 282236 410990
rect 282184 410926 282236 410932
rect 282196 405906 282224 410926
rect 282276 410916 282328 410922
rect 282276 410858 282328 410864
rect 282288 406042 282316 410858
rect 282644 410848 282696 410854
rect 282644 410790 282696 410796
rect 282552 410780 282604 410786
rect 282552 410722 282604 410728
rect 282460 410712 282512 410718
rect 282460 410654 282512 410660
rect 282368 410644 282420 410650
rect 282368 410586 282420 410592
rect 282380 406201 282408 410586
rect 282472 406586 282500 410654
rect 282564 406722 282592 410722
rect 282656 406858 282684 410790
rect 282748 410281 282776 411198
rect 282826 411159 282828 411168
rect 282880 411159 282882 411168
rect 282828 411130 282880 411136
rect 282828 410576 282880 410582
rect 282828 410518 282880 410524
rect 282734 410272 282790 410281
rect 282734 410207 282790 410216
rect 282840 407289 282868 410518
rect 282826 407280 282882 407289
rect 282826 407215 282882 407224
rect 282656 406830 282776 406858
rect 282564 406694 282684 406722
rect 282472 406558 282592 406586
rect 282366 406192 282422 406201
rect 282366 406127 282422 406136
rect 282288 406014 282500 406042
rect 282196 405878 282408 405906
rect 282012 405742 282224 405770
rect 282196 396030 282224 405742
rect 282276 400104 282328 400110
rect 282276 400046 282328 400052
rect 282288 399129 282316 400046
rect 282274 399120 282330 399129
rect 282274 399055 282330 399064
rect 282184 396024 282236 396030
rect 282184 395966 282236 395972
rect 282276 386436 282328 386442
rect 282276 386378 282328 386384
rect 281816 382220 281868 382226
rect 281816 382162 281868 382168
rect 281828 381041 281856 382162
rect 281814 381032 281870 381041
rect 281814 380967 281870 380976
rect 281816 378072 281868 378078
rect 281816 378014 281868 378020
rect 281828 376961 281856 378014
rect 281814 376952 281870 376961
rect 281814 376887 281870 376896
rect 281816 373992 281868 373998
rect 281816 373934 281868 373940
rect 281828 372881 281856 373934
rect 281814 372872 281870 372881
rect 281814 372807 281870 372816
rect 281816 371204 281868 371210
rect 281816 371146 281868 371152
rect 281828 369889 281856 371146
rect 282288 369918 282316 386378
rect 282276 369912 282328 369918
rect 281814 369880 281870 369889
rect 282276 369854 282328 369860
rect 281814 369815 281870 369824
rect 282184 367192 282236 367198
rect 282104 367140 282184 367146
rect 282104 367134 282236 367140
rect 282104 367118 282224 367134
rect 282104 367062 282132 367118
rect 282092 367056 282144 367062
rect 282092 366998 282144 367004
rect 282276 365016 282328 365022
rect 282276 364958 282328 364964
rect 281816 362840 281868 362846
rect 281816 362782 281868 362788
rect 281828 361865 281856 362782
rect 281814 361856 281870 361865
rect 281814 361791 281870 361800
rect 281816 360120 281868 360126
rect 281816 360062 281868 360068
rect 281828 358873 281856 360062
rect 281814 358864 281870 358873
rect 281814 358799 281870 358808
rect 282184 357468 282236 357474
rect 282184 357410 282236 357416
rect 282196 352594 282224 357410
rect 282288 354793 282316 364958
rect 282274 354784 282330 354793
rect 282274 354719 282330 354728
rect 282380 352753 282408 405878
rect 282472 353705 282500 406014
rect 282564 355745 282592 406558
rect 282656 356833 282684 406694
rect 282748 365022 282776 406830
rect 282826 405240 282882 405249
rect 283116 405226 283144 416026
rect 282882 405198 283144 405226
rect 282826 405175 282882 405184
rect 283208 404410 283236 416094
rect 282932 404382 283236 404410
rect 282826 404288 282882 404297
rect 282932 404274 282960 404382
rect 282882 404246 282960 404274
rect 282826 404223 282882 404232
rect 283300 404054 283328 416162
rect 283392 413409 283420 433463
rect 283484 413914 283512 438495
rect 283472 413908 283524 413914
rect 283472 413850 283524 413856
rect 283576 413681 283604 521183
rect 283748 519104 283800 519110
rect 283748 519046 283800 519052
rect 283656 462392 283708 462398
rect 283656 462334 283708 462340
rect 283562 413672 283618 413681
rect 283562 413607 283618 413616
rect 283378 413400 283434 413409
rect 283378 413335 283434 413344
rect 283668 412690 283696 462334
rect 283760 413545 283788 519046
rect 283932 498228 283984 498234
rect 283932 498170 283984 498176
rect 283840 459672 283892 459678
rect 283840 459614 283892 459620
rect 283746 413536 283802 413545
rect 283746 413471 283802 413480
rect 283852 412758 283880 459614
rect 283944 413273 283972 498170
rect 284024 458244 284076 458250
rect 284024 458186 284076 458192
rect 283930 413264 283986 413273
rect 283930 413199 283986 413208
rect 284036 412826 284064 458186
rect 284116 456816 284168 456822
rect 284116 456758 284168 456764
rect 284128 412962 284156 456758
rect 284208 455524 284260 455530
rect 284208 455466 284260 455472
rect 284116 412956 284168 412962
rect 284116 412898 284168 412904
rect 284220 412894 284248 455466
rect 284576 416424 284628 416430
rect 284576 416366 284628 416372
rect 284392 414452 284444 414458
rect 284392 414394 284444 414400
rect 284208 412888 284260 412894
rect 284208 412830 284260 412836
rect 284024 412820 284076 412826
rect 284024 412762 284076 412768
rect 283840 412752 283892 412758
rect 283840 412694 283892 412700
rect 283656 412684 283708 412690
rect 283656 412626 283708 412632
rect 283932 412616 283984 412622
rect 283932 412558 283984 412564
rect 283748 412548 283800 412554
rect 283748 412490 283800 412496
rect 283472 412276 283524 412282
rect 283472 412218 283524 412224
rect 283380 412004 283432 412010
rect 283380 411946 283432 411952
rect 283288 404048 283340 404054
rect 283288 403990 283340 403996
rect 282828 402280 282880 402286
rect 282826 402248 282828 402257
rect 282880 402248 282882 402257
rect 282826 402183 282882 402192
rect 282828 401192 282880 401198
rect 282826 401160 282828 401169
rect 282880 401160 282882 401169
rect 282826 401095 282882 401104
rect 282826 400208 282882 400217
rect 282826 400143 282828 400152
rect 282880 400143 282882 400152
rect 282828 400114 282880 400120
rect 283392 398206 283420 411946
rect 283380 398200 283432 398206
rect 283380 398142 283432 398148
rect 283484 396506 283512 412218
rect 283656 411868 283708 411874
rect 283656 411810 283708 411816
rect 283564 411800 283616 411806
rect 283564 411742 283616 411748
rect 283472 396500 283524 396506
rect 283472 396442 283524 396448
rect 283576 389094 283604 411742
rect 283668 390182 283696 411810
rect 283760 391678 283788 412490
rect 283840 412480 283892 412486
rect 283840 412422 283892 412428
rect 283852 393242 283880 412422
rect 283840 393236 283892 393242
rect 283840 393178 283892 393184
rect 283944 392086 283972 412558
rect 284024 412412 284076 412418
rect 284024 412354 284076 412360
rect 284036 394398 284064 412354
rect 284116 412344 284168 412350
rect 284116 412286 284168 412292
rect 284128 395826 284156 412286
rect 284208 412208 284260 412214
rect 284208 412150 284260 412156
rect 284220 397254 284248 412150
rect 284300 410508 284352 410514
rect 284300 410450 284352 410456
rect 284208 397248 284260 397254
rect 284208 397190 284260 397196
rect 284116 395820 284168 395826
rect 284116 395762 284168 395768
rect 284024 394392 284076 394398
rect 284024 394334 284076 394340
rect 283932 392080 283984 392086
rect 283932 392022 283984 392028
rect 283748 391672 283800 391678
rect 283748 391614 283800 391620
rect 283656 390176 283708 390182
rect 283656 390118 283708 390124
rect 283564 389088 283616 389094
rect 283564 389030 283616 389036
rect 284312 382158 284340 410450
rect 284404 384062 284432 414394
rect 284484 414384 284536 414390
rect 284484 414326 284536 414332
rect 284392 384056 284444 384062
rect 284392 383998 284444 384004
rect 284496 383314 284524 414326
rect 284484 383308 284536 383314
rect 284484 383250 284536 383256
rect 284300 382152 284352 382158
rect 284300 382094 284352 382100
rect 284484 367056 284536 367062
rect 284484 366998 284536 367004
rect 284496 366897 284524 366998
rect 284482 366888 284538 366897
rect 284482 366823 284538 366832
rect 282736 365016 282788 365022
rect 282736 364958 282788 364964
rect 282642 356824 282698 356833
rect 282642 356759 282698 356768
rect 282550 355736 282606 355745
rect 282550 355671 282606 355680
rect 282458 353696 282514 353705
rect 282458 353631 282514 353640
rect 282366 352744 282422 352753
rect 282366 352679 282422 352688
rect 282196 352566 282316 352594
rect 281816 343528 281868 343534
rect 281816 343470 281868 343476
rect 281828 342689 281856 343470
rect 281814 342680 281870 342689
rect 281814 342615 281870 342624
rect 282288 340882 282316 352566
rect 284588 350334 284616 416366
rect 284760 415132 284812 415138
rect 284760 415074 284812 415080
rect 284668 414996 284720 415002
rect 284668 414938 284720 414944
rect 284576 350328 284628 350334
rect 284576 350270 284628 350276
rect 282276 340876 282328 340882
rect 282276 340818 282328 340824
rect 282460 340876 282512 340882
rect 282460 340818 282512 340824
rect 281644 340649 281672 340750
rect 281736 340734 281948 340762
rect 281724 340672 281776 340678
rect 281630 340640 281686 340649
rect 281724 340614 281776 340620
rect 281630 340575 281686 340584
rect 281736 339697 281764 340614
rect 281722 339688 281778 339697
rect 281722 339623 281778 339632
rect 281632 338836 281684 338842
rect 281632 338778 281684 338784
rect 281644 338609 281672 338778
rect 281630 338600 281686 338609
rect 281630 338535 281686 338544
rect 281632 337952 281684 337958
rect 281632 337894 281684 337900
rect 281644 337657 281672 337894
rect 281630 337648 281686 337657
rect 281630 337583 281686 337592
rect 281724 336728 281776 336734
rect 281724 336670 281776 336676
rect 281632 336592 281684 336598
rect 281630 336560 281632 336569
rect 281684 336560 281686 336569
rect 281630 336495 281686 336504
rect 281736 335617 281764 336670
rect 281722 335608 281778 335617
rect 281722 335543 281778 335552
rect 281632 334620 281684 334626
rect 281632 334562 281684 334568
rect 281644 334529 281672 334562
rect 281630 334520 281686 334529
rect 281630 334455 281686 334464
rect 281724 333940 281776 333946
rect 281724 333882 281776 333888
rect 281632 333668 281684 333674
rect 281632 333610 281684 333616
rect 281644 333577 281672 333610
rect 281630 333568 281686 333577
rect 281630 333503 281686 333512
rect 281736 332625 281764 333882
rect 281722 332616 281778 332625
rect 281722 332551 281778 332560
rect 281920 331537 281948 340734
rect 282472 338094 282500 340818
rect 284680 340678 284708 414938
rect 284772 340814 284800 415074
rect 284852 415064 284904 415070
rect 284852 415006 284904 415012
rect 284760 340808 284812 340814
rect 284760 340750 284812 340756
rect 284668 340672 284720 340678
rect 284668 340614 284720 340620
rect 284864 338842 284892 415006
rect 284956 344894 284984 640290
rect 285128 558136 285180 558142
rect 285128 558078 285180 558084
rect 285036 557728 285088 557734
rect 285036 557670 285088 557676
rect 284944 344888 284996 344894
rect 284944 344830 284996 344836
rect 284852 338836 284904 338842
rect 284852 338778 284904 338784
rect 282460 338088 282512 338094
rect 282460 338030 282512 338036
rect 281906 331528 281962 331537
rect 281906 331463 281962 331472
rect 281632 331220 281684 331226
rect 281632 331162 281684 331168
rect 281644 330585 281672 331162
rect 281630 330576 281686 330585
rect 281630 330511 281686 330520
rect 281552 329854 281764 329882
rect 281540 329792 281592 329798
rect 281540 329734 281592 329740
rect 281552 329497 281580 329734
rect 281632 329724 281684 329730
rect 281632 329666 281684 329672
rect 281538 329488 281594 329497
rect 281538 329423 281594 329432
rect 281644 328545 281672 329666
rect 281630 328536 281686 328545
rect 281630 328471 281686 328480
rect 281540 328432 281592 328438
rect 281540 328374 281592 328380
rect 281552 327457 281580 328374
rect 281538 327448 281594 327457
rect 281538 327383 281594 327392
rect 281540 325576 281592 325582
rect 281538 325544 281540 325553
rect 281592 325544 281594 325553
rect 281538 325479 281594 325488
rect 281736 322425 281764 329854
rect 282368 328500 282420 328506
rect 282368 328442 282420 328448
rect 282380 326505 282408 328442
rect 282366 326496 282422 326505
rect 282366 326431 282422 326440
rect 285048 325582 285076 557670
rect 285140 371006 285168 558078
rect 286232 416356 286284 416362
rect 286232 416298 286284 416304
rect 286140 416288 286192 416294
rect 286140 416230 286192 416236
rect 285404 415268 285456 415274
rect 285404 415210 285456 415216
rect 285312 415200 285364 415206
rect 285312 415142 285364 415148
rect 285220 414928 285272 414934
rect 285220 414870 285272 414876
rect 285128 371000 285180 371006
rect 285128 370942 285180 370948
rect 285128 366988 285180 366994
rect 285128 366930 285180 366936
rect 285140 365809 285168 366930
rect 285126 365800 285182 365809
rect 285126 365735 285182 365744
rect 285232 333674 285260 414870
rect 285324 334626 285352 415142
rect 285416 336734 285444 415210
rect 285496 414656 285548 414662
rect 285496 414598 285548 414604
rect 285404 336728 285456 336734
rect 285404 336670 285456 336676
rect 285508 336598 285536 414598
rect 285588 414588 285640 414594
rect 285588 414530 285640 414536
rect 285600 337958 285628 414530
rect 286152 402286 286180 416230
rect 286140 402280 286192 402286
rect 286140 402222 286192 402228
rect 286244 401198 286272 416298
rect 286232 401192 286284 401198
rect 286232 401134 286284 401140
rect 286336 345710 286364 641718
rect 286416 558816 286468 558822
rect 286416 558758 286468 558764
rect 286428 350946 286456 558758
rect 286508 558748 286560 558754
rect 286508 558690 286560 558696
rect 286520 351830 286548 558690
rect 286600 557932 286652 557938
rect 286600 557874 286652 557880
rect 286612 371958 286640 557874
rect 287058 413400 287114 413409
rect 287058 413335 287114 413344
rect 287072 413137 287100 413335
rect 287150 413264 287206 413273
rect 287150 413199 287206 413208
rect 287058 413128 287114 413137
rect 287058 413063 287114 413072
rect 287060 413024 287112 413030
rect 287058 412992 287060 413001
rect 287112 412992 287114 413001
rect 287058 412927 287114 412936
rect 287164 412865 287192 413199
rect 287150 412856 287206 412865
rect 287150 412791 287206 412800
rect 286968 411732 287020 411738
rect 286968 411674 287020 411680
rect 286876 411664 286928 411670
rect 286876 411606 286928 411612
rect 286692 411596 286744 411602
rect 286692 411538 286744 411544
rect 286704 386102 286732 411538
rect 286784 411528 286836 411534
rect 286784 411470 286836 411476
rect 286692 386096 286744 386102
rect 286692 386038 286744 386044
rect 286796 385286 286824 411470
rect 286888 387122 286916 411606
rect 286980 388346 287008 411674
rect 286968 388340 287020 388346
rect 286968 388282 287020 388288
rect 286876 387116 286928 387122
rect 286876 387058 286928 387064
rect 286784 385280 286836 385286
rect 286784 385222 286836 385228
rect 286600 371952 286652 371958
rect 286600 371894 286652 371900
rect 286508 351824 286560 351830
rect 286508 351766 286560 351772
rect 286416 350940 286468 350946
rect 286416 350882 286468 350888
rect 287716 346798 287744 643078
rect 287796 557796 287848 557802
rect 287796 557738 287848 557744
rect 287808 373182 287836 557738
rect 287796 373176 287848 373182
rect 287796 373118 287848 373124
rect 290476 347750 290504 644438
rect 291856 349110 291884 645866
rect 307114 645008 307170 645017
rect 307114 644943 307170 644952
rect 307128 644502 307156 644943
rect 307116 644496 307168 644502
rect 307116 644438 307168 644444
rect 307114 643512 307170 643521
rect 307114 643447 307170 643456
rect 307128 643142 307156 643447
rect 307116 643136 307168 643142
rect 307116 643078 307168 643084
rect 307666 642152 307722 642161
rect 307666 642087 307722 642096
rect 307680 641782 307708 642087
rect 307668 641776 307720 641782
rect 307668 641718 307720 641724
rect 307666 640520 307722 640529
rect 307666 640455 307722 640464
rect 307680 640354 307708 640455
rect 307668 640348 307720 640354
rect 307668 640290 307720 640296
rect 307022 639296 307078 639305
rect 307022 639231 307078 639240
rect 306838 637936 306894 637945
rect 306838 637871 306894 637880
rect 306852 637634 306880 637871
rect 291936 637628 291988 637634
rect 291936 637570 291988 637576
rect 306840 637628 306892 637634
rect 306840 637570 306892 637576
rect 291844 349104 291896 349110
rect 291844 349046 291896 349052
rect 290464 347744 290516 347750
rect 290464 347686 290516 347692
rect 287704 346792 287756 346798
rect 287704 346734 287756 346740
rect 286324 345704 286376 345710
rect 286324 345646 286376 345652
rect 291948 343534 291976 637570
rect 302884 579692 302936 579698
rect 302884 579634 302936 579640
rect 292028 414860 292080 414866
rect 292028 414802 292080 414808
rect 292040 400110 292068 414802
rect 296626 413400 296682 413409
rect 296626 413335 296682 413344
rect 296534 413264 296590 413273
rect 296534 413199 296590 413208
rect 296548 412865 296576 413199
rect 296640 413137 296668 413335
rect 296626 413128 296682 413137
rect 296626 413063 296682 413072
rect 296628 413024 296680 413030
rect 296626 412992 296628 413001
rect 296680 412992 296682 413001
rect 296626 412927 296682 412936
rect 296534 412856 296590 412865
rect 296534 412791 296590 412800
rect 292580 411936 292632 411942
rect 292580 411878 292632 411884
rect 292592 409834 292620 411878
rect 292580 409828 292632 409834
rect 292580 409770 292632 409776
rect 292028 400104 292080 400110
rect 292028 400046 292080 400052
rect 291936 343528 291988 343534
rect 291936 343470 291988 343476
rect 285588 337952 285640 337958
rect 285588 337894 285640 337900
rect 285496 336592 285548 336598
rect 285496 336534 285548 336540
rect 285312 334620 285364 334626
rect 285312 334562 285364 334568
rect 302896 333946 302924 579634
rect 306378 413400 306434 413409
rect 306378 413335 306434 413344
rect 306392 413137 306420 413335
rect 306470 413264 306526 413273
rect 306470 413199 306526 413208
rect 306378 413128 306434 413137
rect 306378 413063 306434 413072
rect 306380 413024 306432 413030
rect 306378 412992 306380 413001
rect 306432 412992 306434 413001
rect 306378 412927 306434 412936
rect 306484 412865 306512 413199
rect 306470 412856 306526 412865
rect 306470 412791 306526 412800
rect 307036 343602 307064 639231
rect 307666 579864 307722 579873
rect 307666 579799 307722 579808
rect 307680 579698 307708 579799
rect 307668 579692 307720 579698
rect 307668 579634 307720 579640
rect 348422 559328 348478 559337
rect 348422 559263 348478 559272
rect 358174 559328 358230 559337
rect 358174 559263 358230 559272
rect 313832 558952 313884 558958
rect 313830 558920 313832 558929
rect 313884 558920 313886 558929
rect 313830 558855 313886 558864
rect 317418 558920 317474 558929
rect 317418 558855 317474 558864
rect 318798 558920 318854 558929
rect 318798 558855 318854 558864
rect 320178 558920 320234 558929
rect 320178 558855 320234 558864
rect 325698 558920 325754 558929
rect 325698 558855 325754 558864
rect 327078 558920 327134 558929
rect 327078 558855 327134 558864
rect 329286 558920 329342 558929
rect 329286 558855 329342 558864
rect 329930 558920 329986 558929
rect 329930 558855 329986 558864
rect 331770 558920 331826 558929
rect 331770 558855 331826 558864
rect 332598 558920 332654 558929
rect 332598 558855 332654 558864
rect 333978 558920 334034 558929
rect 333978 558855 334034 558864
rect 335358 558920 335414 558929
rect 335358 558855 335414 558864
rect 336738 558920 336794 558929
rect 336738 558855 336794 558864
rect 337566 558920 337622 558929
rect 337566 558855 337622 558864
rect 338118 558920 338174 558929
rect 338118 558855 338174 558864
rect 339498 558920 339554 558929
rect 339498 558855 339554 558864
rect 340878 558920 340934 558929
rect 340878 558855 340934 558864
rect 342258 558920 342314 558929
rect 342258 558855 342314 558864
rect 343730 558920 343786 558929
rect 343730 558855 343786 558864
rect 344282 558920 344338 558929
rect 344282 558855 344338 558864
rect 345018 558920 345074 558929
rect 345018 558855 345074 558864
rect 346398 558920 346454 558929
rect 347778 558920 347834 558929
rect 346398 558855 346454 558864
rect 347688 558884 347740 558890
rect 312544 558068 312596 558074
rect 312544 558010 312596 558016
rect 309784 558000 309836 558006
rect 309784 557942 309836 557948
rect 308404 557592 308456 557598
rect 308404 557534 308456 557540
rect 307024 343596 307076 343602
rect 307024 343538 307076 343544
rect 308416 342242 308444 557534
rect 309796 366994 309824 557942
rect 312556 367062 312584 558010
rect 316314 557832 316370 557841
rect 316314 557767 316370 557776
rect 315304 557660 315356 557666
rect 315304 557602 315356 557608
rect 315316 368490 315344 557602
rect 316328 557598 316356 557767
rect 316316 557592 316368 557598
rect 316316 557534 316368 557540
rect 315946 413400 316002 413409
rect 315946 413335 316002 413344
rect 315854 413264 315910 413273
rect 315854 413199 315910 413208
rect 315868 412865 315896 413199
rect 315960 413137 315988 413335
rect 315946 413128 316002 413137
rect 315946 413063 316002 413072
rect 315948 413024 316000 413030
rect 315946 412992 315948 413001
rect 316000 412992 316002 413001
rect 315946 412927 316002 412936
rect 315854 412856 315910 412865
rect 315854 412791 315910 412800
rect 315304 368484 315356 368490
rect 315304 368426 315356 368432
rect 312544 367056 312596 367062
rect 312544 366998 312596 367004
rect 309784 366988 309836 366994
rect 309784 366930 309836 366936
rect 308404 342236 308456 342242
rect 308404 342178 308456 342184
rect 302884 333940 302936 333946
rect 302884 333882 302936 333888
rect 285220 333668 285272 333674
rect 285220 333610 285272 333616
rect 317432 328438 317460 558855
rect 318812 329730 318840 558855
rect 320192 329798 320220 558855
rect 320270 558784 320326 558793
rect 320270 558719 320326 558728
rect 322202 558784 322258 558793
rect 322202 558719 322258 558728
rect 320284 331226 320312 558719
rect 321558 558104 321614 558113
rect 321558 558039 321614 558048
rect 321572 558006 321600 558039
rect 322216 558006 322244 558719
rect 323582 558648 323638 558657
rect 323582 558583 323638 558592
rect 324962 558648 325018 558657
rect 324962 558583 325018 558592
rect 322938 558104 322994 558113
rect 323596 558074 323624 558583
rect 322938 558039 322940 558048
rect 322992 558039 322994 558048
rect 323584 558068 323636 558074
rect 322940 558010 322992 558016
rect 323584 558010 323636 558016
rect 321560 558000 321612 558006
rect 321560 557942 321612 557948
rect 322204 558000 322256 558006
rect 322204 557942 322256 557948
rect 322216 358766 322244 557942
rect 323596 360126 323624 558010
rect 324976 557870 325004 558583
rect 324964 557864 325016 557870
rect 324964 557806 325016 557812
rect 324318 557696 324374 557705
rect 324318 557631 324320 557640
rect 324372 557631 324374 557640
rect 324320 557602 324372 557608
rect 324976 360194 325004 557806
rect 325712 369850 325740 558855
rect 326342 558784 326398 558793
rect 326342 558719 326398 558728
rect 326356 558686 326384 558719
rect 326344 558680 326396 558686
rect 326344 558622 326396 558628
rect 325700 369844 325752 369850
rect 325700 369786 325752 369792
rect 326356 361554 326384 558622
rect 327092 371210 327120 558855
rect 328458 558784 328514 558793
rect 328458 558719 328514 558728
rect 327722 558648 327778 558657
rect 327722 558583 327778 558592
rect 327736 557666 327764 558583
rect 328472 558142 328500 558719
rect 329102 558648 329158 558657
rect 329102 558583 329158 558592
rect 328460 558136 328512 558142
rect 328460 558078 328512 558084
rect 327724 557660 327776 557666
rect 327724 557602 327776 557608
rect 327080 371204 327132 371210
rect 327080 371146 327132 371152
rect 327736 362846 327764 557602
rect 329116 557598 329144 558583
rect 329300 558482 329328 558855
rect 329288 558476 329340 558482
rect 329288 558418 329340 558424
rect 329104 557592 329156 557598
rect 329104 557534 329156 557540
rect 329116 362914 329144 557534
rect 329300 364342 329328 558418
rect 329838 557968 329894 557977
rect 329838 557903 329840 557912
rect 329892 557903 329894 557912
rect 329840 557874 329892 557880
rect 329944 373998 329972 558855
rect 330482 558784 330538 558793
rect 330482 558719 330538 558728
rect 330496 558550 330524 558719
rect 330484 558544 330536 558550
rect 330484 558486 330536 558492
rect 329932 373992 329984 373998
rect 329932 373934 329984 373940
rect 330496 365702 330524 558486
rect 331784 558278 331812 558855
rect 331772 558272 331824 558278
rect 331772 558214 331824 558220
rect 331218 557832 331274 557841
rect 331218 557767 331220 557776
rect 331272 557767 331274 557776
rect 331220 557738 331272 557744
rect 331128 413024 331180 413030
rect 331126 412992 331128 413001
rect 331180 412992 331182 413001
rect 331126 412927 331182 412936
rect 332612 375358 332640 558855
rect 333150 558784 333206 558793
rect 333150 558719 333206 558728
rect 333164 558346 333192 558719
rect 333152 558340 333204 558346
rect 333152 558282 333204 558288
rect 333992 376718 334020 558855
rect 334070 558784 334126 558793
rect 334070 558719 334126 558728
rect 334084 558414 334112 558719
rect 334072 558408 334124 558414
rect 334072 558350 334124 558356
rect 335268 558408 335320 558414
rect 335268 558350 335320 558356
rect 335280 558210 335308 558350
rect 335268 558204 335320 558210
rect 335268 558146 335320 558152
rect 335266 413400 335322 413409
rect 335266 413335 335322 413344
rect 335174 413264 335230 413273
rect 335174 413199 335230 413208
rect 335188 412865 335216 413199
rect 335280 413137 335308 413335
rect 335266 413128 335322 413137
rect 335266 413063 335322 413072
rect 335268 413024 335320 413030
rect 335266 412992 335268 413001
rect 335320 412992 335322 413001
rect 335266 412927 335322 412936
rect 335174 412856 335230 412865
rect 335174 412791 335230 412800
rect 335372 378078 335400 558855
rect 335450 558784 335506 558793
rect 335450 558719 335506 558728
rect 336646 558784 336702 558793
rect 336646 558719 336702 558728
rect 335464 558686 335492 558719
rect 335452 558680 335504 558686
rect 335452 558622 335504 558628
rect 336660 558618 336688 558719
rect 336096 558612 336148 558618
rect 336096 558554 336148 558560
rect 336648 558612 336700 558618
rect 336648 558554 336700 558560
rect 336108 557666 336136 558554
rect 336096 557660 336148 557666
rect 336096 557602 336148 557608
rect 336752 378146 336780 558855
rect 336830 558784 336886 558793
rect 336830 558719 336886 558728
rect 336844 379506 336872 558719
rect 337580 558414 337608 558855
rect 337568 558408 337620 558414
rect 337568 558350 337620 558356
rect 337580 557598 337608 558350
rect 337568 557592 337620 557598
rect 337568 557534 337620 557540
rect 337384 414520 337436 414526
rect 337384 414462 337436 414468
rect 337396 400178 337424 414462
rect 338028 412072 338080 412078
rect 338028 412014 338080 412020
rect 338040 408474 338068 412014
rect 338028 408468 338080 408474
rect 338028 408410 338080 408416
rect 337384 400172 337436 400178
rect 337384 400114 337436 400120
rect 338132 380866 338160 558855
rect 339038 558784 339094 558793
rect 339038 558719 339094 558728
rect 339052 558482 339080 558719
rect 339040 558476 339092 558482
rect 339040 558418 339092 558424
rect 338764 411324 338816 411330
rect 338764 411266 338816 411272
rect 338120 380860 338172 380866
rect 338120 380802 338172 380808
rect 336832 379500 336884 379506
rect 336832 379442 336884 379448
rect 336740 378140 336792 378146
rect 336740 378082 336792 378088
rect 335360 378072 335412 378078
rect 335360 378014 335412 378020
rect 333980 376712 334032 376718
rect 333980 376654 334032 376660
rect 332600 375352 332652 375358
rect 332600 375294 332652 375300
rect 330484 365696 330536 365702
rect 330484 365638 330536 365644
rect 329288 364336 329340 364342
rect 329288 364278 329340 364284
rect 329104 362908 329156 362914
rect 329104 362850 329156 362856
rect 327724 362840 327776 362846
rect 327724 362782 327776 362788
rect 326344 361548 326396 361554
rect 326344 361490 326396 361496
rect 324964 360188 325016 360194
rect 324964 360130 325016 360136
rect 323584 360120 323636 360126
rect 323584 360062 323636 360068
rect 322204 358760 322256 358766
rect 322204 358702 322256 358708
rect 320272 331220 320324 331226
rect 320272 331162 320324 331168
rect 320180 329792 320232 329798
rect 320180 329734 320232 329740
rect 318800 329724 318852 329730
rect 318800 329666 318852 329672
rect 317420 328432 317472 328438
rect 317420 328374 317472 328380
rect 285036 325576 285088 325582
rect 285036 325518 285088 325524
rect 281722 322416 281778 322425
rect 281722 322351 281778 322360
rect 338776 321570 338804 411266
rect 339512 382226 339540 558855
rect 339866 558784 339922 558793
rect 339866 558719 339922 558728
rect 339880 558550 339908 558719
rect 339868 558544 339920 558550
rect 339868 558486 339920 558492
rect 340892 410514 340920 558855
rect 341246 558784 341302 558793
rect 341246 558719 341302 558728
rect 341260 558278 341288 558719
rect 341248 558272 341300 558278
rect 341248 558214 341300 558220
rect 342272 414390 342300 558855
rect 342534 558784 342590 558793
rect 342534 558719 342590 558728
rect 343638 558784 343694 558793
rect 343638 558719 343694 558728
rect 342548 558346 342576 558719
rect 342536 558340 342588 558346
rect 342536 558282 342588 558288
rect 343652 558210 343680 558719
rect 343640 558204 343692 558210
rect 343640 558146 343692 558152
rect 343638 557696 343694 557705
rect 343638 557631 343694 557640
rect 342260 414384 342312 414390
rect 342260 414326 342312 414332
rect 343088 412140 343140 412146
rect 343088 412082 343140 412088
rect 343100 411194 343128 412082
rect 343652 411534 343680 557631
rect 343744 414458 343772 558855
rect 344296 558686 344324 558855
rect 344284 558680 344336 558686
rect 344284 558622 344336 558628
rect 343732 414452 343784 414458
rect 343732 414394 343784 414400
rect 345032 411602 345060 558855
rect 346030 558784 346086 558793
rect 346030 558719 346086 558728
rect 346044 558618 346072 558719
rect 346032 558612 346084 558618
rect 346032 558554 346084 558560
rect 346412 411670 346440 558855
rect 347778 558855 347834 558864
rect 347688 558826 347740 558832
rect 347700 558793 347728 558826
rect 347686 558784 347742 558793
rect 347686 558719 347742 558728
rect 347700 558414 347728 558719
rect 347688 558408 347740 558414
rect 347688 558350 347740 558356
rect 347792 411738 347820 558855
rect 348238 558784 348294 558793
rect 348238 558719 348294 558728
rect 348252 558482 348280 558719
rect 348240 558476 348292 558482
rect 348240 558418 348292 558424
rect 348436 558346 348464 559263
rect 349158 558920 349214 558929
rect 349158 558855 349214 558864
rect 352010 558920 352066 558929
rect 352010 558855 352066 558864
rect 356058 558920 356114 558929
rect 356058 558855 356060 558864
rect 348424 558340 348476 558346
rect 348424 558282 348476 558288
rect 349172 411806 349200 558855
rect 349710 558784 349766 558793
rect 349710 558719 349766 558728
rect 349724 558550 349752 558719
rect 349712 558544 349764 558550
rect 349712 558486 349764 558492
rect 350538 558512 350594 558521
rect 350538 558447 350594 558456
rect 350552 558278 350580 558447
rect 350540 558272 350592 558278
rect 350540 558214 350592 558220
rect 352024 558210 352052 558855
rect 356112 558855 356114 558864
rect 356060 558826 356112 558832
rect 353298 558784 353354 558793
rect 353298 558719 353354 558728
rect 354678 558784 354734 558793
rect 354678 558719 354734 558728
rect 353312 558686 353340 558719
rect 353300 558680 353352 558686
rect 353300 558622 353352 558628
rect 354692 558618 354720 558719
rect 354680 558612 354732 558618
rect 354680 558554 354732 558560
rect 358188 558550 358216 559263
rect 358176 558544 358228 558550
rect 357438 558512 357494 558521
rect 358176 558486 358228 558492
rect 357438 558447 357440 558456
rect 357492 558447 357494 558456
rect 357440 558418 357492 558424
rect 352564 558408 352616 558414
rect 352564 558350 352616 558356
rect 352012 558204 352064 558210
rect 352012 558146 352064 558152
rect 352102 557696 352158 557705
rect 352102 557631 352158 557640
rect 350630 557560 350686 557569
rect 350630 557495 350686 557504
rect 350448 413024 350500 413030
rect 350446 412992 350448 413001
rect 350500 412992 350502 413001
rect 350446 412927 350502 412936
rect 350644 411874 350672 557495
rect 352010 555520 352066 555529
rect 352010 555455 352066 555464
rect 352024 412554 352052 555455
rect 352116 412622 352144 557631
rect 352576 419422 352604 558350
rect 352656 558340 352708 558346
rect 352656 558282 352708 558288
rect 352668 420918 352696 558282
rect 353944 558272 353996 558278
rect 353944 558214 353996 558220
rect 353298 557560 353354 557569
rect 353298 557495 353354 557504
rect 352656 420912 352708 420918
rect 352656 420854 352708 420860
rect 352564 419416 352616 419422
rect 352564 419358 352616 419364
rect 352104 412616 352156 412622
rect 352104 412558 352156 412564
rect 352012 412548 352064 412554
rect 352012 412490 352064 412496
rect 353312 412486 353340 557495
rect 353956 422278 353984 558214
rect 354036 558204 354088 558210
rect 354036 558146 354088 558152
rect 354048 423570 354076 558146
rect 356704 558136 356756 558142
rect 356704 558078 356756 558084
rect 355324 558068 355376 558074
rect 355324 558010 355376 558016
rect 354678 557560 354734 557569
rect 354678 557495 354734 557504
rect 354128 523116 354180 523122
rect 354128 523058 354180 523064
rect 354036 423564 354088 423570
rect 354036 423506 354088 423512
rect 353944 422272 353996 422278
rect 353944 422214 353996 422220
rect 354140 413817 354168 523058
rect 354126 413808 354182 413817
rect 354126 413743 354182 413752
rect 354586 413400 354642 413409
rect 354586 413335 354642 413344
rect 354494 413264 354550 413273
rect 354494 413199 354550 413208
rect 354508 412865 354536 413199
rect 354600 413137 354628 413335
rect 354586 413128 354642 413137
rect 354586 413063 354642 413072
rect 354588 413024 354640 413030
rect 354586 412992 354588 413001
rect 354640 412992 354642 413001
rect 354586 412927 354642 412936
rect 354494 412856 354550 412865
rect 354494 412791 354550 412800
rect 353300 412480 353352 412486
rect 353300 412422 353352 412428
rect 354692 412418 354720 557495
rect 355336 423638 355364 558010
rect 355416 557932 355468 557938
rect 355416 557874 355468 557880
rect 355428 425066 355456 557874
rect 356150 557560 356206 557569
rect 356150 557495 356206 557504
rect 355416 425060 355468 425066
rect 355416 425002 355468 425008
rect 355324 423632 355376 423638
rect 355324 423574 355376 423580
rect 354680 412412 354732 412418
rect 354680 412354 354732 412360
rect 356164 412350 356192 557495
rect 356716 426426 356744 558078
rect 356796 558000 356848 558006
rect 356796 557942 356848 557948
rect 356808 427718 356836 557942
rect 358084 557864 358136 557870
rect 358084 557806 358136 557812
rect 357530 557560 357586 557569
rect 357530 557495 357586 557504
rect 356796 427712 356848 427718
rect 356796 427654 356848 427660
rect 356704 426420 356756 426426
rect 356704 426362 356756 426368
rect 356152 412344 356204 412350
rect 356152 412286 356204 412292
rect 357544 412282 357572 557495
rect 358096 427786 358124 557806
rect 358176 557796 358228 557802
rect 358176 557738 358228 557744
rect 358188 429146 358216 557738
rect 358910 555520 358966 555529
rect 358910 555455 358966 555464
rect 358176 429140 358228 429146
rect 358176 429082 358228 429088
rect 358084 427780 358136 427786
rect 358084 427722 358136 427728
rect 357532 412276 357584 412282
rect 357532 412218 357584 412224
rect 358924 412214 358952 555455
rect 367100 538348 367152 538354
rect 367100 538290 367152 538296
rect 367112 413953 367140 538290
rect 368480 538280 368532 538286
rect 368480 538222 368532 538228
rect 367744 523048 367796 523054
rect 367744 522990 367796 522996
rect 367098 413944 367154 413953
rect 367098 413879 367154 413888
rect 364338 413400 364394 413409
rect 364338 413335 364394 413344
rect 364352 413137 364380 413335
rect 364338 413128 364394 413137
rect 364338 413063 364394 413072
rect 364340 413024 364392 413030
rect 364340 412966 364392 412972
rect 364352 412865 364380 412966
rect 364338 412856 364394 412865
rect 364338 412791 364394 412800
rect 367098 412720 367154 412729
rect 367756 412690 367784 522990
rect 368492 413137 368520 538222
rect 369860 536852 369912 536858
rect 369860 536794 369912 536800
rect 368572 460964 368624 460970
rect 368572 460906 368624 460912
rect 368584 413953 368612 460906
rect 368570 413944 368626 413953
rect 368570 413879 368626 413888
rect 369872 413137 369900 536794
rect 371240 535492 371292 535498
rect 371240 535434 371292 535440
rect 369952 459604 370004 459610
rect 369952 459546 370004 459552
rect 369964 413953 369992 459546
rect 371252 413953 371280 535434
rect 372620 534200 372672 534206
rect 372620 534142 372672 534148
rect 371884 524476 371936 524482
rect 371884 524418 371936 524424
rect 371896 414089 371924 524418
rect 371882 414080 371938 414089
rect 371882 414015 371938 414024
rect 372632 413953 372660 534142
rect 374000 534132 374052 534138
rect 374000 534074 374052 534080
rect 373264 433356 373316 433362
rect 373264 433298 373316 433304
rect 369950 413944 370006 413953
rect 369950 413879 370006 413888
rect 371238 413944 371294 413953
rect 371238 413879 371294 413888
rect 372618 413944 372674 413953
rect 372618 413879 372674 413888
rect 368294 413128 368350 413137
rect 368294 413063 368350 413072
rect 368478 413128 368534 413137
rect 368478 413063 368534 413072
rect 369858 413128 369914 413137
rect 369858 413063 369914 413072
rect 370962 413128 371018 413137
rect 370962 413063 371018 413072
rect 368308 412729 368336 413063
rect 370976 412729 371004 413063
rect 371330 412856 371386 412865
rect 373276 412826 373304 433298
rect 373906 413400 373962 413409
rect 373906 413335 373962 413344
rect 373920 413001 373948 413335
rect 374012 413273 374040 534074
rect 375380 532772 375432 532778
rect 375380 532714 375432 532720
rect 374644 525836 374696 525842
rect 374644 525778 374696 525784
rect 373998 413264 374054 413273
rect 373998 413199 374054 413208
rect 373906 412992 373962 413001
rect 373906 412927 373962 412936
rect 374000 412956 374052 412962
rect 374000 412898 374052 412904
rect 374012 412865 374040 412898
rect 374656 412894 374684 525778
rect 374736 434784 374788 434790
rect 374736 434726 374788 434732
rect 374184 412888 374236 412894
rect 373998 412856 374054 412865
rect 371330 412791 371386 412800
rect 372620 412820 372672 412826
rect 371344 412758 371372 412791
rect 372620 412762 372672 412768
rect 373264 412820 373316 412826
rect 374184 412830 374236 412836
rect 374644 412888 374696 412894
rect 374644 412830 374696 412836
rect 373998 412791 374054 412800
rect 373264 412762 373316 412768
rect 371240 412752 371292 412758
rect 368294 412720 368350 412729
rect 367098 412655 367100 412664
rect 367152 412655 367154 412664
rect 367744 412684 367796 412690
rect 367100 412626 367152 412632
rect 368294 412655 368350 412664
rect 370962 412720 371018 412729
rect 370962 412655 371018 412664
rect 371238 412720 371240 412729
rect 371332 412752 371384 412758
rect 371292 412720 371294 412729
rect 372632 412729 372660 412762
rect 374196 412729 374224 412830
rect 374748 412758 374776 434726
rect 375392 413273 375420 532714
rect 375472 531412 375524 531418
rect 375472 531354 375524 531360
rect 375378 413264 375434 413273
rect 375378 413199 375434 413208
rect 375484 413137 375512 531354
rect 376760 531344 376812 531350
rect 376760 531286 376812 531292
rect 376024 527264 376076 527270
rect 376024 527206 376076 527212
rect 375564 455456 375616 455462
rect 375564 455398 375616 455404
rect 375576 413273 375604 455398
rect 376036 413506 376064 527206
rect 376024 413500 376076 413506
rect 376024 413442 376076 413448
rect 376772 413273 376800 531286
rect 378232 529984 378284 529990
rect 378232 529926 378284 529932
rect 377404 436212 377456 436218
rect 377404 436154 377456 436160
rect 375562 413264 375618 413273
rect 375562 413199 375618 413208
rect 376758 413264 376814 413273
rect 376758 413199 376814 413208
rect 375470 413128 375526 413137
rect 375470 413063 375526 413072
rect 376760 413024 376812 413030
rect 376760 412966 376812 412972
rect 376772 412865 376800 412966
rect 376758 412856 376814 412865
rect 376758 412791 376814 412800
rect 377416 412758 377444 436154
rect 378244 413273 378272 529926
rect 379612 528624 379664 528630
rect 379612 528566 379664 528572
rect 378784 501084 378836 501090
rect 378784 501026 378836 501032
rect 378230 413264 378286 413273
rect 378796 413234 378824 501026
rect 379624 413953 379652 528566
rect 380992 527196 381044 527202
rect 380992 527138 381044 527144
rect 380164 436144 380216 436150
rect 380164 436086 380216 436092
rect 379610 413944 379666 413953
rect 379610 413879 379666 413888
rect 379794 413400 379850 413409
rect 379794 413335 379850 413344
rect 378230 413199 378286 413208
rect 378784 413228 378836 413234
rect 378784 413170 378836 413176
rect 378140 413092 378192 413098
rect 378140 413034 378192 413040
rect 379612 413092 379664 413098
rect 379612 413034 379664 413040
rect 378152 412865 378180 413034
rect 379624 412865 379652 413034
rect 379808 412865 379836 413335
rect 380176 413098 380204 436086
rect 380622 413808 380678 413817
rect 380622 413743 380678 413752
rect 380636 413273 380664 413743
rect 381004 413409 381032 527138
rect 387892 521688 387944 521694
rect 387892 521630 387944 521636
rect 387064 516248 387116 516254
rect 387064 516190 387116 516196
rect 385684 514820 385736 514826
rect 385684 514762 385736 514768
rect 384304 510672 384356 510678
rect 384304 510614 384356 510620
rect 382924 507952 382976 507958
rect 382924 507894 382976 507900
rect 381544 438932 381596 438938
rect 381544 438874 381596 438880
rect 381556 413574 381584 438874
rect 381544 413568 381596 413574
rect 381544 413510 381596 413516
rect 382280 413500 382332 413506
rect 382280 413442 382332 413448
rect 382292 413409 382320 413442
rect 380990 413400 381046 413409
rect 382278 413400 382334 413409
rect 380990 413335 381046 413344
rect 382188 413364 382240 413370
rect 382278 413335 382334 413344
rect 382188 413306 382240 413312
rect 380622 413264 380678 413273
rect 380622 413199 380678 413208
rect 382200 413137 382228 413306
rect 382372 413296 382424 413302
rect 382372 413238 382424 413244
rect 382384 413137 382412 413238
rect 382186 413128 382242 413137
rect 380164 413092 380216 413098
rect 382186 413063 382242 413072
rect 382370 413128 382426 413137
rect 382370 413063 382426 413072
rect 380164 413034 380216 413040
rect 380900 413024 380952 413030
rect 380900 412966 380952 412972
rect 378138 412856 378194 412865
rect 378138 412791 378194 412800
rect 379610 412856 379666 412865
rect 379610 412791 379666 412800
rect 379794 412856 379850 412865
rect 379794 412791 379850 412800
rect 374736 412752 374788 412758
rect 371332 412694 371384 412700
rect 372618 412720 372674 412729
rect 371238 412655 371294 412664
rect 372618 412655 372674 412664
rect 374182 412720 374238 412729
rect 374736 412694 374788 412700
rect 377404 412752 377456 412758
rect 380912 412729 380940 412966
rect 382936 412962 382964 507894
rect 383016 506524 383068 506530
rect 383016 506466 383068 506472
rect 383028 413302 383056 506466
rect 383108 505232 383160 505238
rect 383108 505174 383160 505180
rect 383120 414050 383148 505174
rect 383200 502376 383252 502382
rect 383200 502318 383252 502324
rect 383108 414044 383160 414050
rect 383108 413986 383160 413992
rect 383212 413506 383240 502318
rect 384316 413817 384344 510614
rect 384396 440428 384448 440434
rect 384396 440370 384448 440376
rect 384302 413808 384358 413817
rect 384302 413743 384358 413752
rect 383200 413500 383252 413506
rect 383200 413442 383252 413448
rect 383016 413296 383068 413302
rect 383016 413238 383068 413244
rect 384408 413234 384436 440370
rect 385314 413536 385370 413545
rect 385314 413471 385370 413480
rect 384304 413228 384356 413234
rect 384304 413170 384356 413176
rect 384396 413228 384448 413234
rect 384396 413170 384448 413176
rect 383660 413160 383712 413166
rect 383660 413102 383712 413108
rect 382924 412956 382976 412962
rect 382924 412898 382976 412904
rect 382280 412888 382332 412894
rect 382280 412830 382332 412836
rect 382292 412729 382320 412830
rect 383672 412729 383700 413102
rect 384316 412962 384344 413170
rect 385328 413137 385356 413471
rect 385038 413128 385094 413137
rect 385038 413063 385094 413072
rect 385314 413128 385370 413137
rect 385314 413063 385370 413072
rect 384304 412956 384356 412962
rect 384304 412898 384356 412904
rect 385052 412894 385080 413063
rect 385696 412894 385724 514762
rect 385776 512100 385828 512106
rect 385776 512042 385828 512048
rect 385788 413098 385816 512042
rect 386420 413636 386472 413642
rect 386420 413578 386472 413584
rect 386432 413545 386460 413578
rect 386418 413536 386474 413545
rect 386418 413471 386474 413480
rect 385776 413092 385828 413098
rect 385776 413034 385828 413040
rect 385040 412888 385092 412894
rect 385040 412830 385092 412836
rect 385684 412888 385736 412894
rect 385684 412830 385736 412836
rect 387076 412729 387104 516190
rect 387156 440292 387208 440298
rect 387156 440234 387208 440240
rect 387168 413846 387196 440234
rect 387904 413953 387932 521630
rect 390652 520328 390704 520334
rect 390652 520270 390704 520276
rect 388444 430704 388496 430710
rect 388444 430646 388496 430652
rect 388456 419370 388484 430646
rect 388456 419342 388576 419370
rect 387890 413944 387946 413953
rect 387890 413879 387946 413888
rect 387156 413840 387208 413846
rect 387156 413782 387208 413788
rect 388548 413642 388576 419342
rect 390664 413953 390692 520270
rect 392032 517540 392084 517546
rect 392032 517482 392084 517488
rect 392044 413953 392072 517482
rect 406384 466540 406436 466546
rect 406384 466482 406436 466488
rect 402980 413976 403032 413982
rect 390650 413944 390706 413953
rect 390650 413879 390706 413888
rect 392030 413944 392086 413953
rect 402978 413944 402980 413953
rect 403032 413944 403034 413953
rect 392030 413879 392086 413888
rect 396080 413908 396132 413914
rect 402978 413879 403034 413888
rect 396080 413850 396132 413856
rect 391940 413840 391992 413846
rect 391938 413808 391940 413817
rect 396092 413817 396120 413850
rect 391992 413808 391994 413817
rect 389272 413772 389324 413778
rect 391938 413743 391994 413752
rect 396078 413808 396134 413817
rect 406396 413778 406424 466482
rect 407776 413953 407804 650490
rect 516416 650480 516468 650486
rect 516416 650422 516468 650428
rect 516428 649913 516456 650422
rect 516414 649904 516470 649913
rect 516414 649839 516470 649848
rect 438122 646096 438178 646105
rect 438122 646031 438178 646040
rect 413928 558952 413980 558958
rect 413928 558894 413980 558900
rect 413940 558482 413968 558894
rect 413928 558476 413980 558482
rect 413928 558418 413980 558424
rect 410524 501016 410576 501022
rect 410524 500958 410576 500964
rect 409144 470688 409196 470694
rect 409144 470630 409196 470636
rect 407762 413944 407818 413953
rect 409156 413914 409184 470630
rect 410536 413953 410564 500958
rect 411904 470620 411956 470626
rect 411904 470562 411956 470568
rect 410522 413944 410578 413953
rect 407762 413879 407818 413888
rect 409144 413908 409196 413914
rect 410522 413879 410578 413888
rect 409144 413850 409196 413856
rect 396078 413743 396134 413752
rect 406384 413772 406436 413778
rect 389272 413714 389324 413720
rect 406384 413714 406436 413720
rect 389180 413704 389232 413710
rect 389180 413646 389232 413652
rect 388536 413636 388588 413642
rect 388536 413578 388588 413584
rect 389192 413545 389220 413646
rect 389178 413536 389234 413545
rect 389178 413471 389234 413480
rect 387800 413024 387852 413030
rect 389284 413001 389312 413714
rect 404360 413636 404412 413642
rect 404360 413578 404412 413584
rect 394700 413568 394752 413574
rect 389362 413536 389418 413545
rect 389362 413471 389418 413480
rect 394698 413536 394700 413545
rect 404372 413545 404400 413578
rect 394752 413536 394754 413545
rect 404358 413536 404414 413545
rect 394698 413471 394754 413480
rect 401600 413500 401652 413506
rect 387800 412966 387852 412972
rect 389086 412992 389142 413001
rect 387812 412729 387840 412966
rect 389086 412927 389142 412936
rect 389270 412992 389326 413001
rect 389270 412927 389326 412936
rect 389100 412842 389128 412927
rect 389376 412842 389404 413471
rect 404358 413471 404414 413480
rect 401600 413442 401652 413448
rect 397460 413432 397512 413438
rect 393226 413400 393282 413409
rect 393226 413335 393282 413344
rect 397458 413400 397460 413409
rect 401612 413409 401640 413442
rect 397512 413400 397514 413409
rect 401598 413400 401654 413409
rect 397458 413335 397514 413344
rect 397552 413364 397604 413370
rect 390560 413160 390612 413166
rect 390560 413102 390612 413108
rect 390572 413001 390600 413102
rect 390558 412992 390614 413001
rect 390558 412927 390614 412936
rect 393240 412865 393268 413335
rect 401598 413335 401654 413344
rect 397552 413306 397604 413312
rect 393320 413228 393372 413234
rect 393320 413170 393372 413176
rect 393332 413001 393360 413170
rect 397564 413137 397592 413306
rect 398840 413296 398892 413302
rect 398840 413238 398892 413244
rect 398852 413137 398880 413238
rect 397550 413128 397606 413137
rect 396080 413092 396132 413098
rect 397550 413063 397606 413072
rect 398838 413128 398894 413137
rect 398838 413063 398894 413072
rect 396080 413034 396132 413040
rect 396092 413001 396120 413034
rect 397460 413024 397512 413030
rect 393318 412992 393374 413001
rect 393318 412927 393374 412936
rect 396078 412992 396134 413001
rect 396078 412927 396134 412936
rect 397458 412992 397460 413001
rect 397512 412992 397514 413001
rect 397458 412927 397514 412936
rect 403164 412956 403216 412962
rect 403164 412898 403216 412904
rect 394700 412888 394752 412894
rect 389100 412814 389404 412842
rect 393226 412856 393282 412865
rect 393226 412791 393282 412800
rect 394698 412856 394700 412865
rect 403176 412865 403204 412898
rect 394752 412856 394754 412865
rect 394698 412791 394754 412800
rect 400218 412856 400274 412865
rect 400218 412791 400220 412800
rect 400272 412791 400274 412800
rect 403162 412856 403218 412865
rect 410536 412826 410564 413879
rect 411916 413846 411944 470562
rect 413940 413953 413968 558418
rect 419540 516180 419592 516186
rect 419540 516122 419592 516128
rect 416320 496868 416372 496874
rect 416320 496810 416372 496816
rect 416044 473408 416096 473414
rect 416044 473350 416096 473356
rect 413926 413944 413982 413953
rect 413926 413879 413982 413888
rect 411904 413840 411956 413846
rect 411904 413782 411956 413788
rect 413940 413642 413968 413879
rect 416056 413710 416084 473350
rect 416044 413704 416096 413710
rect 416044 413646 416096 413652
rect 413928 413636 413980 413642
rect 413928 413578 413980 413584
rect 403162 412791 403218 412800
rect 410524 412820 410576 412826
rect 400220 412762 400272 412768
rect 410524 412762 410576 412768
rect 398840 412752 398892 412758
rect 377404 412694 377456 412700
rect 380898 412720 380954 412729
rect 374182 412655 374238 412664
rect 380898 412655 380954 412664
rect 382278 412720 382334 412729
rect 382278 412655 382334 412664
rect 383658 412720 383714 412729
rect 383658 412655 383714 412664
rect 385038 412720 385094 412729
rect 385038 412655 385040 412664
rect 367744 412626 367796 412632
rect 385092 412655 385094 412664
rect 387062 412720 387118 412729
rect 387062 412655 387118 412664
rect 387798 412720 387854 412729
rect 387798 412655 387854 412664
rect 398838 412720 398840 412729
rect 398892 412720 398894 412729
rect 398838 412655 398894 412664
rect 400218 412720 400274 412729
rect 400218 412655 400220 412664
rect 385040 412626 385092 412632
rect 400272 412655 400274 412664
rect 400220 412626 400272 412632
rect 358912 412208 358964 412214
rect 358912 412150 358964 412156
rect 350632 411868 350684 411874
rect 350632 411810 350684 411816
rect 349160 411800 349212 411806
rect 349160 411742 349212 411748
rect 347780 411732 347832 411738
rect 347780 411674 347832 411680
rect 346400 411664 346452 411670
rect 346400 411606 346452 411612
rect 345020 411596 345072 411602
rect 345020 411538 345072 411544
rect 343640 411528 343692 411534
rect 343640 411470 343692 411476
rect 405738 411496 405794 411505
rect 405738 411431 405794 411440
rect 405752 411330 405780 411431
rect 405740 411324 405792 411330
rect 405740 411266 405792 411272
rect 343088 411188 343140 411194
rect 343088 411130 343140 411136
rect 340880 410508 340932 410514
rect 340880 410450 340932 410456
rect 416332 391354 416360 496810
rect 417424 463820 417476 463826
rect 417424 463762 417476 463768
rect 416780 429208 416832 429214
rect 416780 429150 416832 429156
rect 416792 393009 416820 429150
rect 417436 413166 417464 463762
rect 417424 413160 417476 413166
rect 417424 413102 417476 413108
rect 416778 393000 416834 393009
rect 416778 392935 416834 392944
rect 416410 391368 416466 391377
rect 416332 391326 416410 391354
rect 416410 391303 416466 391312
rect 339500 382220 339552 382226
rect 339500 382162 339552 382168
rect 419552 341057 419580 516122
rect 419632 513392 419684 513398
rect 419632 513334 419684 513340
rect 419644 341737 419672 513334
rect 419724 512032 419776 512038
rect 419724 511974 419776 511980
rect 419736 343777 419764 511974
rect 419816 509312 419868 509318
rect 419816 509254 419868 509260
rect 419828 344457 419856 509254
rect 419908 507884 419960 507890
rect 419908 507826 419960 507832
rect 419920 346633 419948 507826
rect 420000 505164 420052 505170
rect 420000 505106 420052 505112
rect 419906 346624 419962 346633
rect 419906 346559 419962 346568
rect 419814 344448 419870 344457
rect 419814 344383 419870 344392
rect 419722 343768 419778 343777
rect 419722 343703 419778 343712
rect 419630 341728 419686 341737
rect 419630 341663 419686 341672
rect 419538 341048 419594 341057
rect 419538 340983 419594 340992
rect 419552 325145 419580 340983
rect 419644 325825 419672 341663
rect 419736 328137 419764 343703
rect 419828 329225 419856 344383
rect 419920 330993 419948 346559
rect 420012 346497 420040 505106
rect 420092 503736 420144 503742
rect 420092 503678 420144 503684
rect 420104 349217 420132 503678
rect 435364 480276 435416 480282
rect 435364 480218 435416 480224
rect 431224 478984 431276 478990
rect 431224 478926 431276 478932
rect 429844 477556 429896 477562
rect 429844 477498 429896 477504
rect 428464 476128 428516 476134
rect 428464 476070 428516 476076
rect 424324 474836 424376 474842
rect 424324 474778 424376 474784
rect 424336 413642 424364 474778
rect 427084 474768 427136 474774
rect 427084 474710 427136 474716
rect 420184 413636 420236 413642
rect 420184 413578 420236 413584
rect 424324 413636 424376 413642
rect 424324 413578 424376 413584
rect 420196 412865 420224 413578
rect 427096 413438 427124 474710
rect 428476 413506 428504 476070
rect 428464 413500 428516 413506
rect 428464 413442 428516 413448
rect 427084 413432 427136 413438
rect 427084 413374 427136 413380
rect 429856 413370 429884 477498
rect 431236 413574 431264 478926
rect 433984 478916 434036 478922
rect 433984 478858 434036 478864
rect 431224 413568 431276 413574
rect 431224 413510 431276 413516
rect 429844 413364 429896 413370
rect 429844 413306 429896 413312
rect 433996 413234 434024 478858
rect 435376 413302 435404 480218
rect 438136 415138 438164 646031
rect 438214 645008 438270 645017
rect 438214 644943 438270 644952
rect 438124 415132 438176 415138
rect 438124 415074 438176 415080
rect 438228 415002 438256 644943
rect 438306 643240 438362 643249
rect 438306 643175 438362 643184
rect 438320 415070 438348 643175
rect 438398 642016 438454 642025
rect 438398 641951 438454 641960
rect 438308 415064 438360 415070
rect 438308 415006 438360 415012
rect 438216 414996 438268 415002
rect 438216 414938 438268 414944
rect 438412 414594 438440 641951
rect 438490 640384 438546 640393
rect 438490 640319 438546 640328
rect 438504 414662 438532 640319
rect 438582 639296 438638 639305
rect 438582 639231 438638 639240
rect 438596 415274 438624 639231
rect 438674 637664 438730 637673
rect 438674 637599 438730 637608
rect 438584 415268 438636 415274
rect 438584 415210 438636 415216
rect 438688 415206 438716 637599
rect 518912 589393 518940 652734
rect 518898 589384 518954 589393
rect 518898 589319 518954 589328
rect 518912 587761 518940 589319
rect 518898 587752 518954 587761
rect 518898 587687 518954 587696
rect 438766 579728 438822 579737
rect 438766 579663 438822 579672
rect 438676 415200 438728 415206
rect 438676 415142 438728 415148
rect 438492 414656 438544 414662
rect 438492 414598 438544 414604
rect 438400 414588 438452 414594
rect 438400 414530 438452 414536
rect 435364 413296 435416 413302
rect 435364 413238 435416 413244
rect 433984 413228 434036 413234
rect 433984 413170 434036 413176
rect 420182 412856 420238 412865
rect 420182 412791 420238 412800
rect 420090 349208 420146 349217
rect 420090 349143 420146 349152
rect 419998 346488 420054 346497
rect 419998 346423 420054 346432
rect 420012 332081 420040 346423
rect 420104 333713 420132 349143
rect 420090 333704 420146 333713
rect 420090 333639 420146 333648
rect 419998 332072 420054 332081
rect 419998 332007 420054 332016
rect 419906 330984 419962 330993
rect 419906 330919 419962 330928
rect 419814 329216 419870 329225
rect 419814 329151 419870 329160
rect 419722 328128 419778 328137
rect 419722 328063 419778 328072
rect 419630 325816 419686 325825
rect 419630 325751 419686 325760
rect 419538 325136 419594 325145
rect 419538 325071 419594 325080
rect 282828 321564 282880 321570
rect 282828 321506 282880 321512
rect 338764 321564 338816 321570
rect 338764 321506 338816 321512
rect 282840 321473 282868 321506
rect 282826 321464 282882 321473
rect 282826 321399 282882 321408
rect 279330 320920 279386 320929
rect 279160 320878 279330 320906
rect 279330 320855 279386 320864
rect 60950 320062 61424 320090
rect 44088 318776 44140 318782
rect 44088 318718 44140 318724
rect 20628 318708 20680 318714
rect 20628 318650 20680 318656
rect 16488 318028 16540 318034
rect 16488 317970 16540 317976
rect 12348 317960 12400 317966
rect 12348 317902 12400 317908
rect 5448 317892 5500 317898
rect 5448 317834 5500 317840
rect 1676 3188 1728 3194
rect 1676 3130 1728 3136
rect 572 2984 624 2990
rect 572 2926 624 2932
rect 584 480 612 2926
rect 1688 480 1716 3130
rect 4068 3052 4120 3058
rect 4068 2994 4120 3000
rect 2872 2848 2924 2854
rect 2872 2790 2924 2796
rect 2884 480 2912 2790
rect 4080 480 4108 2994
rect 5460 610 5488 317834
rect 12360 3534 12388 317902
rect 14832 4072 14884 4078
rect 14832 4014 14884 4020
rect 13636 4004 13688 4010
rect 13636 3946 13688 3952
rect 11244 3528 11296 3534
rect 11244 3470 11296 3476
rect 12348 3528 12400 3534
rect 12348 3470 12400 3476
rect 10048 3324 10100 3330
rect 10048 3266 10100 3272
rect 8852 3256 8904 3262
rect 8852 3198 8904 3204
rect 7656 3188 7708 3194
rect 7656 3130 7708 3136
rect 6460 3120 6512 3126
rect 6460 3062 6512 3068
rect 5264 604 5316 610
rect 5264 546 5316 552
rect 5448 604 5500 610
rect 5448 546 5500 552
rect 5276 480 5304 546
rect 6472 480 6500 3062
rect 7668 480 7696 3130
rect 8864 480 8892 3198
rect 10060 480 10088 3266
rect 11256 480 11284 3470
rect 12440 3392 12492 3398
rect 12440 3334 12492 3340
rect 12452 480 12480 3334
rect 13648 480 13676 3946
rect 14844 480 14872 4014
rect 16500 3534 16528 317970
rect 17224 4004 17276 4010
rect 17224 3946 17276 3952
rect 16028 3528 16080 3534
rect 16028 3470 16080 3476
rect 16488 3528 16540 3534
rect 16488 3470 16540 3476
rect 16040 480 16068 3470
rect 17236 480 17264 3946
rect 18328 3936 18380 3942
rect 18328 3878 18380 3884
rect 18340 480 18368 3878
rect 20640 3874 20668 318650
rect 22008 318640 22060 318646
rect 22008 318582 22060 318588
rect 22020 3874 22048 318582
rect 23388 318572 23440 318578
rect 23388 318514 23440 318520
rect 23400 4842 23428 318514
rect 30288 318504 30340 318510
rect 30288 318446 30340 318452
rect 28908 318436 28960 318442
rect 28908 318378 28960 318384
rect 23124 4814 23428 4842
rect 19524 3868 19576 3874
rect 19524 3810 19576 3816
rect 20628 3868 20680 3874
rect 20628 3810 20680 3816
rect 20720 3868 20772 3874
rect 20720 3810 20772 3816
rect 22008 3868 22060 3874
rect 22008 3810 22060 3816
rect 19536 480 19564 3810
rect 20732 480 20760 3810
rect 21916 3800 21968 3806
rect 21916 3742 21968 3748
rect 21928 480 21956 3742
rect 23124 480 23152 4814
rect 25504 3800 25556 3806
rect 25504 3742 25556 3748
rect 24308 3732 24360 3738
rect 24308 3674 24360 3680
rect 24320 480 24348 3674
rect 25516 480 25544 3742
rect 26700 3664 26752 3670
rect 26700 3606 26752 3612
rect 26712 480 26740 3606
rect 28920 3534 28948 318378
rect 30300 3534 30328 318446
rect 31668 318368 31720 318374
rect 31668 318310 31720 318316
rect 27896 3528 27948 3534
rect 27896 3470 27948 3476
rect 28908 3528 28960 3534
rect 28908 3470 28960 3476
rect 29092 3528 29144 3534
rect 29092 3470 29144 3476
rect 30288 3528 30340 3534
rect 31680 3482 31708 318310
rect 42708 318300 42760 318306
rect 42708 318242 42760 318248
rect 35808 318232 35860 318238
rect 35808 318174 35860 318180
rect 33048 317484 33100 317490
rect 33048 317426 33100 317432
rect 33060 3482 33088 317426
rect 35820 3602 35848 318174
rect 39948 318164 40000 318170
rect 39948 318106 40000 318112
rect 38476 317552 38528 317558
rect 38476 317494 38528 317500
rect 38488 4842 38516 317494
rect 39960 4842 39988 318106
rect 42720 4842 42748 318242
rect 44100 4842 44128 318718
rect 61396 318102 61424 320062
rect 62224 320062 62882 320090
rect 63696 320062 64814 320090
rect 66364 320062 66746 320090
rect 61384 318096 61436 318102
rect 61384 318038 61436 318044
rect 57888 317824 57940 317830
rect 57888 317766 57940 317772
rect 53748 317756 53800 317762
rect 53748 317698 53800 317704
rect 50988 317688 51040 317694
rect 50988 317630 51040 317636
rect 48136 317620 48188 317626
rect 48136 317562 48188 317568
rect 37372 4820 37424 4826
rect 38488 4814 38608 4842
rect 37372 4762 37424 4768
rect 34980 3596 35032 3602
rect 34980 3538 35032 3544
rect 35808 3596 35860 3602
rect 35808 3538 35860 3544
rect 30288 3470 30340 3476
rect 27908 480 27936 3470
rect 29104 480 29132 3470
rect 30196 3460 30248 3466
rect 30196 3402 30248 3408
rect 31496 3454 31708 3482
rect 32692 3454 33088 3482
rect 33876 3528 33928 3534
rect 33876 3470 33928 3476
rect 30208 1714 30236 3402
rect 30208 1686 30328 1714
rect 30300 480 30328 1686
rect 31496 480 31524 3454
rect 32692 480 32720 3454
rect 33888 480 33916 3470
rect 34992 480 35020 3538
rect 36176 3460 36228 3466
rect 36176 3402 36228 3408
rect 36188 480 36216 3402
rect 37384 480 37412 4762
rect 38580 480 38608 4814
rect 39776 4814 39988 4842
rect 42168 4814 42748 4842
rect 43364 4814 44128 4842
rect 39776 480 39804 4814
rect 40958 3904 41014 3913
rect 40958 3839 41014 3848
rect 40972 480 41000 3839
rect 42168 480 42196 4814
rect 43364 480 43392 4814
rect 48148 4214 48176 317562
rect 49332 6180 49384 6186
rect 49332 6122 49384 6128
rect 46940 4208 46992 4214
rect 46940 4150 46992 4156
rect 48136 4208 48188 4214
rect 48136 4150 48188 4156
rect 48228 4208 48280 4214
rect 48228 4150 48280 4156
rect 44546 4040 44602 4049
rect 44546 3975 44602 3984
rect 44560 480 44588 3975
rect 45742 3768 45798 3777
rect 45742 3703 45798 3712
rect 45756 480 45784 3703
rect 46952 480 46980 4150
rect 48240 2122 48268 4150
rect 48148 2094 48268 2122
rect 48148 480 48176 2094
rect 49344 480 49372 6122
rect 51000 3482 51028 317630
rect 51632 4276 51684 4282
rect 51632 4218 51684 4224
rect 50540 3454 51028 3482
rect 50540 480 50568 3454
rect 51644 480 51672 4218
rect 53760 3482 53788 317698
rect 55220 4344 55272 4350
rect 55220 4286 55272 4292
rect 54022 3632 54078 3641
rect 54022 3567 54078 3576
rect 52840 3454 53788 3482
rect 52840 480 52868 3454
rect 54036 480 54064 3567
rect 55232 480 55260 4286
rect 55310 4176 55366 4185
rect 55310 4111 55366 4120
rect 55324 4078 55352 4111
rect 55312 4072 55364 4078
rect 55312 4014 55364 4020
rect 56414 3496 56470 3505
rect 56414 3431 56470 3440
rect 56428 480 56456 3431
rect 57900 626 57928 317766
rect 60004 4888 60056 4894
rect 60004 4830 60056 4836
rect 58808 4412 58860 4418
rect 58808 4354 58860 4360
rect 57624 598 57928 626
rect 57624 480 57652 598
rect 58820 480 58848 4354
rect 60016 480 60044 4830
rect 61396 2990 61424 318038
rect 61384 2984 61436 2990
rect 61384 2926 61436 2932
rect 61200 2916 61252 2922
rect 61200 2858 61252 2864
rect 61212 480 61240 2858
rect 62224 2854 62252 320062
rect 62396 4480 62448 4486
rect 62396 4422 62448 4428
rect 62212 2848 62264 2854
rect 62212 2790 62264 2796
rect 62408 480 62436 4422
rect 63696 3398 63724 320062
rect 64786 318608 64842 318617
rect 64786 318543 64842 318552
rect 64694 4176 64750 4185
rect 64694 4111 64750 4120
rect 64708 4078 64736 4111
rect 64696 4072 64748 4078
rect 64696 4014 64748 4020
rect 63684 3392 63736 3398
rect 63684 3334 63736 3340
rect 63592 2848 63644 2854
rect 63592 2790 63644 2796
rect 63604 480 63632 2790
rect 64800 480 64828 318543
rect 65984 4548 66036 4554
rect 65984 4490 66036 4496
rect 65996 480 66024 4490
rect 66364 3058 66392 320062
rect 68664 317898 68692 320076
rect 70412 320062 70610 320090
rect 71976 320062 72542 320090
rect 68652 317892 68704 317898
rect 68652 317834 68704 317840
rect 67180 4956 67232 4962
rect 67180 4898 67232 4904
rect 66352 3052 66404 3058
rect 66352 2994 66404 3000
rect 67192 480 67220 4898
rect 69480 4616 69532 4622
rect 69480 4558 69532 4564
rect 68284 2984 68336 2990
rect 68284 2926 68336 2932
rect 68296 480 68324 2926
rect 69492 480 69520 4558
rect 70412 3126 70440 320062
rect 71872 3324 71924 3330
rect 71872 3266 71924 3272
rect 70400 3120 70452 3126
rect 70400 3062 70452 3068
rect 70676 3052 70728 3058
rect 70676 2994 70728 3000
rect 70688 480 70716 2994
rect 71884 480 71912 3266
rect 71976 3126 72004 320062
rect 74446 318472 74502 318481
rect 74446 318407 74502 318416
rect 72976 317892 73028 317898
rect 72976 317834 73028 317840
rect 72988 3330 73016 317834
rect 73068 4684 73120 4690
rect 73068 4626 73120 4632
rect 72976 3324 73028 3330
rect 72976 3266 73028 3272
rect 71964 3120 72016 3126
rect 71964 3062 72016 3068
rect 73080 480 73108 4626
rect 74460 610 74488 318407
rect 74552 3330 74580 320076
rect 76024 320062 76498 320090
rect 74540 3324 74592 3330
rect 74540 3266 74592 3272
rect 76024 3194 76052 320062
rect 78416 317966 78444 320076
rect 80164 320062 80362 320090
rect 81452 320062 82294 320090
rect 78404 317960 78456 317966
rect 78404 317902 78456 317908
rect 79968 317960 80020 317966
rect 79968 317902 80020 317908
rect 76656 4752 76708 4758
rect 76656 4694 76708 4700
rect 76012 3188 76064 3194
rect 76012 3130 76064 3136
rect 75460 3120 75512 3126
rect 75460 3062 75512 3068
rect 74264 604 74316 610
rect 74264 546 74316 552
rect 74448 604 74500 610
rect 74448 546 74500 552
rect 74276 480 74304 546
rect 75472 480 75500 3062
rect 76668 480 76696 4694
rect 79980 3398 80008 317902
rect 79048 3392 79100 3398
rect 79048 3334 79100 3340
rect 79968 3392 80020 3398
rect 79968 3334 80020 3340
rect 77852 3188 77904 3194
rect 77852 3130 77904 3136
rect 77864 480 77892 3130
rect 79060 480 79088 3334
rect 80164 3330 80192 320062
rect 80244 5500 80296 5506
rect 80244 5442 80296 5448
rect 80152 3324 80204 3330
rect 80152 3266 80204 3272
rect 80256 480 80284 5442
rect 81452 4162 81480 320062
rect 82634 318336 82690 318345
rect 82634 318271 82690 318280
rect 81360 4146 81480 4162
rect 81348 4140 81480 4146
rect 81400 4134 81480 4140
rect 81348 4082 81400 4088
rect 82648 4078 82676 318271
rect 82726 318200 82782 318209
rect 82726 318135 82782 318144
rect 81440 4072 81492 4078
rect 81440 4014 81492 4020
rect 82636 4072 82688 4078
rect 82636 4014 82688 4020
rect 81452 480 81480 4014
rect 82740 3482 82768 318135
rect 83832 5432 83884 5438
rect 83832 5374 83884 5380
rect 82648 3454 82768 3482
rect 82648 480 82676 3454
rect 83844 480 83872 5374
rect 84212 3398 84240 320076
rect 86236 318034 86264 320076
rect 86972 320062 88182 320090
rect 89732 320062 90114 320090
rect 86224 318028 86276 318034
rect 86224 317970 86276 317976
rect 86972 4010 87000 320062
rect 87328 5364 87380 5370
rect 87328 5306 87380 5312
rect 86960 4004 87012 4010
rect 86960 3946 87012 3952
rect 84936 3936 84988 3942
rect 84936 3878 84988 3884
rect 84200 3392 84252 3398
rect 84200 3334 84252 3340
rect 84948 480 84976 3878
rect 86132 3256 86184 3262
rect 86132 3198 86184 3204
rect 86144 480 86172 3198
rect 87340 480 87368 5306
rect 89732 4146 89760 320062
rect 92032 318714 92060 320076
rect 92020 318708 92072 318714
rect 92020 318650 92072 318656
rect 92388 318708 92440 318714
rect 92388 318650 92440 318656
rect 90916 318028 90968 318034
rect 90916 317970 90968 317976
rect 89720 4140 89772 4146
rect 89720 4082 89772 4088
rect 90928 3398 90956 317970
rect 91008 5296 91060 5302
rect 91008 5238 91060 5244
rect 89720 3392 89772 3398
rect 89720 3334 89772 3340
rect 90916 3392 90968 3398
rect 90916 3334 90968 3340
rect 88524 3324 88576 3330
rect 88524 3266 88576 3272
rect 88536 480 88564 3266
rect 89732 480 89760 3334
rect 91020 2666 91048 5238
rect 92400 3346 92428 318650
rect 93964 318646 93992 320076
rect 95252 320062 95910 320090
rect 93952 318640 94004 318646
rect 93952 318582 94004 318588
rect 94504 5228 94556 5234
rect 94504 5170 94556 5176
rect 93308 4140 93360 4146
rect 93308 4082 93360 4088
rect 90928 2638 91048 2666
rect 92124 3318 92428 3346
rect 90928 480 90956 2638
rect 92124 480 92152 3318
rect 93320 480 93348 4082
rect 94516 480 94544 5170
rect 95252 3874 95280 320062
rect 96528 318640 96580 318646
rect 96528 318582 96580 318588
rect 95240 3868 95292 3874
rect 95240 3810 95292 3816
rect 96540 3738 96568 318582
rect 97920 318578 97948 320076
rect 99392 320062 99866 320090
rect 100772 320062 101798 320090
rect 103532 320062 103730 320090
rect 97908 318572 97960 318578
rect 97908 318514 97960 318520
rect 98000 318572 98052 318578
rect 98000 318514 98052 318520
rect 98012 318458 98040 318514
rect 97920 318430 98040 318458
rect 97920 3738 97948 318430
rect 98092 5160 98144 5166
rect 98092 5102 98144 5108
rect 95700 3732 95752 3738
rect 95700 3674 95752 3680
rect 96528 3732 96580 3738
rect 96528 3674 96580 3680
rect 96896 3732 96948 3738
rect 96896 3674 96948 3680
rect 97908 3732 97960 3738
rect 97908 3674 97960 3680
rect 95712 480 95740 3674
rect 96908 480 96936 3674
rect 98104 480 98132 5102
rect 99288 4004 99340 4010
rect 99288 3946 99340 3952
rect 99300 480 99328 3946
rect 99392 3874 99420 320062
rect 99380 3868 99432 3874
rect 99380 3810 99432 3816
rect 100484 3868 100536 3874
rect 100484 3810 100536 3816
rect 100496 480 100524 3810
rect 100772 3806 100800 320062
rect 101588 5092 101640 5098
rect 101588 5034 101640 5040
rect 100760 3800 100812 3806
rect 100760 3742 100812 3748
rect 101600 480 101628 5034
rect 102784 3936 102836 3942
rect 102784 3878 102836 3884
rect 102796 480 102824 3878
rect 103532 3670 103560 320062
rect 105648 318442 105676 320076
rect 107580 318510 107608 320076
rect 109052 320062 109526 320090
rect 107568 318504 107620 318510
rect 107568 318446 107620 318452
rect 107660 318504 107712 318510
rect 107660 318446 107712 318452
rect 105636 318436 105688 318442
rect 105636 318378 105688 318384
rect 107672 318322 107700 318446
rect 107580 318294 107700 318322
rect 104806 318064 104862 318073
rect 104806 317999 104862 318008
rect 103520 3664 103572 3670
rect 103520 3606 103572 3612
rect 104820 3602 104848 317999
rect 105176 5024 105228 5030
rect 105176 4966 105228 4972
rect 103980 3596 104032 3602
rect 103980 3538 104032 3544
rect 104808 3596 104860 3602
rect 104808 3538 104860 3544
rect 103992 480 104020 3538
rect 105188 480 105216 4966
rect 107476 3800 107528 3806
rect 107476 3742 107528 3748
rect 106372 3596 106424 3602
rect 106372 3538 106424 3544
rect 106384 480 106412 3538
rect 107488 1986 107516 3742
rect 107580 3602 107608 318294
rect 108762 5536 108818 5545
rect 108762 5471 108818 5480
rect 107568 3596 107620 3602
rect 107568 3538 107620 3544
rect 107488 1958 107608 1986
rect 107580 480 107608 1958
rect 108776 480 108804 5471
rect 109052 3670 109080 320062
rect 110328 318436 110380 318442
rect 110328 318378 110380 318384
rect 109040 3664 109092 3670
rect 109040 3606 109092 3612
rect 110340 3346 110368 318378
rect 111536 318374 111564 320076
rect 111524 318368 111576 318374
rect 111524 318310 111576 318316
rect 111708 318368 111760 318374
rect 111708 318310 111760 318316
rect 111720 3602 111748 318310
rect 113468 317490 113496 320076
rect 114572 320062 115414 320090
rect 113456 317484 113508 317490
rect 113456 317426 113508 317432
rect 112350 5400 112406 5409
rect 112350 5335 112406 5344
rect 111156 3596 111208 3602
rect 111156 3538 111208 3544
rect 111708 3596 111760 3602
rect 111708 3538 111760 3544
rect 109972 3318 110368 3346
rect 109972 480 110000 3318
rect 111168 480 111196 3538
rect 112364 480 112392 5335
rect 113548 3732 113600 3738
rect 113548 3674 113600 3680
rect 113560 480 113588 3674
rect 114572 3534 114600 320062
rect 117332 318238 117360 320076
rect 118712 320062 119278 320090
rect 120092 320062 121210 320090
rect 117320 318232 117372 318238
rect 117320 318174 117372 318180
rect 118608 318232 118660 318238
rect 118608 318174 118660 318180
rect 115938 4856 115994 4865
rect 115938 4791 115994 4800
rect 114744 3800 114796 3806
rect 114744 3742 114796 3748
rect 114560 3528 114612 3534
rect 114560 3470 114612 3476
rect 114756 480 114784 3742
rect 115952 480 115980 4791
rect 117136 3664 117188 3670
rect 117136 3606 117188 3612
rect 117148 480 117176 3606
rect 118620 3346 118648 318174
rect 118712 3466 118740 320062
rect 120092 4826 120120 320062
rect 123220 317558 123248 320076
rect 125152 318170 125180 320076
rect 126992 320062 127098 320090
rect 125140 318164 125192 318170
rect 125140 318106 125192 318112
rect 125508 318164 125560 318170
rect 125508 318106 125560 318112
rect 123208 317552 123260 317558
rect 123208 317494 123260 317500
rect 123484 317552 123536 317558
rect 123484 317494 123536 317500
rect 120080 4820 120132 4826
rect 120080 4762 120132 4768
rect 123024 4820 123076 4826
rect 123024 4762 123076 4768
rect 119436 3596 119488 3602
rect 119436 3538 119488 3544
rect 118700 3460 118752 3466
rect 118700 3402 118752 3408
rect 118252 3318 118648 3346
rect 118252 480 118280 3318
rect 119448 480 119476 3538
rect 120632 3528 120684 3534
rect 120632 3470 120684 3476
rect 120644 480 120672 3470
rect 121826 3360 121882 3369
rect 121826 3295 121882 3304
rect 121840 480 121868 3295
rect 123036 480 123064 4762
rect 123496 4049 123524 317494
rect 124864 317484 124916 317490
rect 124864 317426 124916 317432
rect 124876 4894 124904 317426
rect 124864 4888 124916 4894
rect 124864 4830 124916 4836
rect 123482 4040 123538 4049
rect 123482 3975 123538 3984
rect 125520 3482 125548 318106
rect 126612 4888 126664 4894
rect 126612 4830 126664 4836
rect 124220 3460 124272 3466
rect 124220 3402 124272 3408
rect 125428 3454 125548 3482
rect 124232 480 124260 3402
rect 125428 480 125456 3454
rect 126624 480 126652 4830
rect 126992 3913 127020 320062
rect 129016 318306 129044 320076
rect 130948 318782 130976 320076
rect 132880 318782 132908 320076
rect 133892 320062 134918 320090
rect 130936 318776 130988 318782
rect 130936 318718 130988 318724
rect 132868 318776 132920 318782
rect 132868 318718 132920 318724
rect 133144 318776 133196 318782
rect 133144 318718 133196 318724
rect 129004 318300 129056 318306
rect 129004 318242 129056 318248
rect 130384 318300 130436 318306
rect 130384 318242 130436 318248
rect 129002 5264 129058 5273
rect 129002 5199 129058 5208
rect 127806 5128 127862 5137
rect 127806 5063 127862 5072
rect 126978 3904 127034 3913
rect 126978 3839 127034 3848
rect 127820 480 127848 5063
rect 129016 480 129044 5199
rect 130200 4888 130252 4894
rect 130200 4830 130252 4836
rect 130212 480 130240 4830
rect 130396 4826 130424 318242
rect 131764 317552 131816 317558
rect 131764 317494 131816 317500
rect 131776 4962 131804 317494
rect 132590 4992 132646 5001
rect 131764 4956 131816 4962
rect 132590 4927 132646 4936
rect 131764 4898 131816 4904
rect 130384 4820 130436 4826
rect 130384 4762 130436 4768
rect 131396 4820 131448 4826
rect 131396 4762 131448 4768
rect 131408 480 131436 4762
rect 132604 480 132632 4927
rect 133156 4865 133184 318718
rect 133142 4856 133198 4865
rect 133142 4791 133198 4800
rect 133892 3777 133920 320062
rect 136836 317626 136864 320076
rect 138032 320062 138782 320090
rect 139412 320062 140714 320090
rect 136824 317620 136876 317626
rect 136824 317562 136876 317568
rect 134890 4856 134946 4865
rect 134890 4791 134946 4800
rect 133878 3768 133934 3777
rect 133878 3703 133934 3712
rect 134904 480 134932 4791
rect 138032 4214 138060 320062
rect 139412 6186 139440 320062
rect 142632 317694 142660 320076
rect 143552 320062 144578 320090
rect 142620 317688 142672 317694
rect 142620 317630 142672 317636
rect 139400 6180 139452 6186
rect 139400 6122 139452 6128
rect 143552 4282 143580 320062
rect 146588 317762 146616 320076
rect 147692 320062 148534 320090
rect 146576 317756 146628 317762
rect 146576 317698 146628 317704
rect 143540 4276 143592 4282
rect 143540 4218 143592 4224
rect 138020 4208 138072 4214
rect 138020 4150 138072 4156
rect 147692 3641 147720 320062
rect 150452 4350 150480 320076
rect 151832 320062 152398 320090
rect 150440 4344 150492 4350
rect 150440 4286 150492 4292
rect 147678 3632 147734 3641
rect 147678 3567 147734 3576
rect 151832 3505 151860 320062
rect 154316 317830 154344 320076
rect 155972 320062 156262 320090
rect 154304 317824 154356 317830
rect 154304 317766 154356 317772
rect 155972 4418 156000 320062
rect 158180 317490 158208 320076
rect 160112 320062 160218 320090
rect 161492 320062 162150 320090
rect 162872 320062 164082 320090
rect 158168 317484 158220 317490
rect 158168 317426 158220 317432
rect 155960 4412 156012 4418
rect 155960 4354 156012 4360
rect 151818 3496 151874 3505
rect 151818 3431 151874 3440
rect 160112 2922 160140 320062
rect 161492 4486 161520 320062
rect 161480 4480 161532 4486
rect 161480 4422 161532 4428
rect 160100 2916 160152 2922
rect 160100 2858 160152 2864
rect 162872 2854 162900 320062
rect 166000 318617 166028 320076
rect 167012 320062 167946 320090
rect 165986 318608 166042 318617
rect 165986 318543 166042 318552
rect 167012 4554 167040 320062
rect 169864 317558 169892 320076
rect 171152 320062 171902 320090
rect 172532 320062 173834 320090
rect 175292 320062 175766 320090
rect 169852 317552 169904 317558
rect 169852 317494 169904 317500
rect 167000 4548 167052 4554
rect 167000 4490 167052 4496
rect 171152 2990 171180 320062
rect 172532 4622 172560 320062
rect 172520 4616 172572 4622
rect 172520 4558 172572 4564
rect 175292 3058 175320 320062
rect 177684 317898 177712 320076
rect 179432 320062 179630 320090
rect 177672 317892 177724 317898
rect 177672 317834 177724 317840
rect 179432 4690 179460 320062
rect 181548 318481 181576 320076
rect 181534 318472 181590 318481
rect 181534 318407 181590 318416
rect 179420 4684 179472 4690
rect 179420 4626 179472 4632
rect 183572 3126 183600 320076
rect 184952 320062 185518 320090
rect 186332 320062 187450 320090
rect 184952 4758 184980 320062
rect 184940 4752 184992 4758
rect 184940 4694 184992 4700
rect 186332 3194 186360 320062
rect 189368 317966 189396 320076
rect 190472 320062 191314 320090
rect 189356 317960 189408 317966
rect 189356 317902 189408 317908
rect 190472 5506 190500 320062
rect 193232 318345 193260 320076
rect 193218 318336 193274 318345
rect 193218 318271 193274 318280
rect 195164 318209 195192 320076
rect 195992 320062 197202 320090
rect 198752 320062 199134 320090
rect 200132 320062 201066 320090
rect 202892 320062 202998 320090
rect 204272 320062 204930 320090
rect 195150 318200 195206 318209
rect 195150 318135 195206 318144
rect 190460 5500 190512 5506
rect 190460 5442 190512 5448
rect 195992 5438 196020 320062
rect 195980 5432 196032 5438
rect 195980 5374 196032 5380
rect 198752 3262 198780 320062
rect 200132 3330 200160 320062
rect 202892 5370 202920 320062
rect 202880 5364 202932 5370
rect 202880 5306 202932 5312
rect 204272 3398 204300 320062
rect 206848 318034 206876 320076
rect 208412 320062 208886 320090
rect 206836 318028 206888 318034
rect 206836 317970 206888 317976
rect 208412 5302 208440 320062
rect 210804 318714 210832 320076
rect 212552 320062 212750 320090
rect 213932 320062 214682 320090
rect 210792 318708 210844 318714
rect 210792 318650 210844 318656
rect 208400 5296 208452 5302
rect 208400 5238 208452 5244
rect 212552 4146 212580 320062
rect 213932 5234 213960 320062
rect 216600 318646 216628 320076
rect 216588 318640 216640 318646
rect 216588 318582 216640 318588
rect 218532 318578 218560 320076
rect 219452 320062 220570 320090
rect 222212 320062 222502 320090
rect 223592 320062 224434 320090
rect 218520 318572 218572 318578
rect 218520 318514 218572 318520
rect 213920 5228 213972 5234
rect 213920 5170 213972 5176
rect 219452 5166 219480 320062
rect 219440 5160 219492 5166
rect 219440 5102 219492 5108
rect 212540 4140 212592 4146
rect 212540 4082 212592 4088
rect 222212 4010 222240 320062
rect 223592 4078 223620 320062
rect 226352 5098 226380 320076
rect 227732 320062 228298 320090
rect 226340 5092 226392 5098
rect 226340 5034 226392 5040
rect 223580 4072 223632 4078
rect 223580 4014 223632 4020
rect 222200 4004 222252 4010
rect 222200 3946 222252 3952
rect 227732 3942 227760 320062
rect 230216 318073 230244 320076
rect 231872 320062 232254 320090
rect 230202 318064 230258 318073
rect 230202 317999 230258 318008
rect 231872 5030 231900 320062
rect 234172 318510 234200 320076
rect 236012 320062 236118 320090
rect 237392 320062 238050 320090
rect 234160 318504 234212 318510
rect 234160 318446 234212 318452
rect 231860 5024 231912 5030
rect 231860 4966 231912 4972
rect 227720 3936 227772 3942
rect 227720 3878 227772 3884
rect 236012 3874 236040 320062
rect 237392 5545 237420 320062
rect 239968 318442 239996 320076
rect 239956 318436 240008 318442
rect 239956 318378 240008 318384
rect 241900 318374 241928 320076
rect 242912 320062 243846 320090
rect 245672 320062 245870 320090
rect 247052 320062 247802 320090
rect 241888 318368 241940 318374
rect 241888 318310 241940 318316
rect 237378 5536 237434 5545
rect 237378 5471 237434 5480
rect 242912 5409 242940 320062
rect 242898 5400 242954 5409
rect 242898 5335 242954 5344
rect 236000 3868 236052 3874
rect 236000 3810 236052 3816
rect 245672 3738 245700 320062
rect 247052 3806 247080 320062
rect 249720 318782 249748 320076
rect 251192 320062 251666 320090
rect 249708 318776 249760 318782
rect 249708 318718 249760 318724
rect 247040 3800 247092 3806
rect 247040 3742 247092 3748
rect 245660 3732 245712 3738
rect 245660 3674 245712 3680
rect 251192 3670 251220 320062
rect 253584 318238 253612 320076
rect 255332 320062 255530 320090
rect 256712 320062 257554 320090
rect 253572 318232 253624 318238
rect 253572 318174 253624 318180
rect 251180 3664 251232 3670
rect 251180 3606 251232 3612
rect 255332 3602 255360 320062
rect 255320 3596 255372 3602
rect 255320 3538 255372 3544
rect 256712 3534 256740 320062
rect 256700 3528 256752 3534
rect 256700 3470 256752 3476
rect 204260 3392 204312 3398
rect 259472 3369 259500 320076
rect 261404 318306 261432 320076
rect 262232 320062 263350 320090
rect 261392 318300 261444 318306
rect 261392 318242 261444 318248
rect 262232 3466 262260 320062
rect 265268 318170 265296 320076
rect 266372 320062 267214 320090
rect 269132 320062 269238 320090
rect 270512 320062 271170 320090
rect 271892 320062 273102 320090
rect 274652 320062 275034 320090
rect 276032 320062 276966 320090
rect 278792 320062 278898 320090
rect 265256 318164 265308 318170
rect 265256 318106 265308 318112
rect 266372 4962 266400 320062
rect 269132 5137 269160 320062
rect 270512 5273 270540 320062
rect 270498 5264 270554 5273
rect 270498 5199 270554 5208
rect 269118 5128 269174 5137
rect 269118 5063 269174 5072
rect 266360 4956 266412 4962
rect 266360 4898 266412 4904
rect 271892 4894 271920 320062
rect 271880 4888 271932 4894
rect 271880 4830 271932 4836
rect 274652 4826 274680 320062
rect 276032 5001 276060 320062
rect 276018 4992 276074 5001
rect 276018 4927 276074 4936
rect 278792 4865 278820 320062
rect 420196 318782 420224 412791
rect 438780 411126 438808 579663
rect 443090 558920 443146 558929
rect 443090 558855 443146 558864
rect 445758 558920 445814 558929
rect 445758 558855 445814 558864
rect 451278 558920 451334 558929
rect 451278 558855 451334 558864
rect 452658 558920 452714 558929
rect 452658 558855 452714 558864
rect 453670 558920 453726 558929
rect 453670 558855 453726 558864
rect 454038 558920 454094 558929
rect 454038 558855 454094 558864
rect 455418 558920 455474 558929
rect 455418 558855 455474 558864
rect 456798 558920 456854 558929
rect 456798 558855 456854 558864
rect 458178 558920 458234 558929
rect 458178 558855 458234 558864
rect 459558 558920 459614 558929
rect 459558 558855 459614 558864
rect 461030 558920 461086 558929
rect 461030 558855 461086 558864
rect 461674 558920 461730 558929
rect 461674 558855 461730 558864
rect 462318 558920 462374 558929
rect 462318 558855 462374 558864
rect 463698 558920 463754 558929
rect 463698 558855 463754 558864
rect 465078 558920 465134 558929
rect 465078 558855 465134 558864
rect 466458 558920 466514 558929
rect 466458 558855 466514 558864
rect 467838 558920 467894 558929
rect 468758 558920 468814 558929
rect 467838 558855 467894 558864
rect 468024 558884 468076 558890
rect 443104 558482 443132 558855
rect 443092 558476 443144 558482
rect 443092 558418 443144 558424
rect 442264 481772 442316 481778
rect 442264 481714 442316 481720
rect 442276 413098 442304 481714
rect 445024 481704 445076 481710
rect 445024 481646 445076 481652
rect 442264 413092 442316 413098
rect 442264 413034 442316 413040
rect 445036 413030 445064 481646
rect 445772 414934 445800 558855
rect 449898 557832 449954 557841
rect 449898 557767 449954 557776
rect 449912 557734 449940 557767
rect 449900 557728 449952 557734
rect 449900 557670 449952 557676
rect 449164 484424 449216 484430
rect 449164 484366 449216 484372
rect 446404 483064 446456 483070
rect 446404 483006 446456 483012
rect 445760 414928 445812 414934
rect 445760 414870 445812 414876
rect 445024 413024 445076 413030
rect 445024 412966 445076 412972
rect 446416 412962 446444 483006
rect 447784 465112 447836 465118
rect 447784 465054 447836 465060
rect 447796 413982 447824 465054
rect 447784 413976 447836 413982
rect 447784 413918 447836 413924
rect 446404 412956 446456 412962
rect 446404 412898 446456 412904
rect 449176 412894 449204 484366
rect 449164 412888 449216 412894
rect 449164 412830 449216 412836
rect 438768 411120 438820 411126
rect 438768 411062 438820 411068
rect 451292 411058 451320 558855
rect 452672 412010 452700 558855
rect 453684 558822 453712 558855
rect 453672 558816 453724 558822
rect 452750 558784 452806 558793
rect 453672 558758 453724 558764
rect 452750 558719 452806 558728
rect 452764 414866 452792 558719
rect 453302 558648 453358 558657
rect 453302 558583 453358 558592
rect 453316 558550 453344 558583
rect 453304 558544 453356 558550
rect 453304 558486 453356 558492
rect 453316 416430 453344 558486
rect 453304 416424 453356 416430
rect 453304 416366 453356 416372
rect 452752 414860 452804 414866
rect 452752 414802 452804 414808
rect 454052 414526 454080 558855
rect 454774 558784 454830 558793
rect 454774 558719 454776 558728
rect 454828 558719 454830 558728
rect 454776 558690 454828 558696
rect 454788 558482 454816 558690
rect 454776 558476 454828 558482
rect 454776 558418 454828 558424
rect 455432 416362 455460 558855
rect 456062 558784 456118 558793
rect 456062 558719 456118 558728
rect 456076 558686 456104 558719
rect 456064 558680 456116 558686
rect 456064 558622 456116 558628
rect 455420 416356 455472 416362
rect 455420 416298 455472 416304
rect 454040 414520 454092 414526
rect 454040 414462 454092 414468
rect 452660 412004 452712 412010
rect 452660 411946 452712 411952
rect 451280 411052 451332 411058
rect 451280 410994 451332 411000
rect 456076 410990 456104 558622
rect 456812 416294 456840 558855
rect 457456 558822 457484 558853
rect 457444 558816 457496 558822
rect 457442 558784 457444 558793
rect 457496 558784 457498 558793
rect 457442 558719 457498 558728
rect 456800 416288 456852 416294
rect 456800 416230 456852 416236
rect 456064 410984 456116 410990
rect 456064 410926 456116 410932
rect 457456 410922 457484 558719
rect 458192 416226 458220 558855
rect 458822 558784 458878 558793
rect 458822 558719 458824 558728
rect 458876 558719 458878 558728
rect 458824 558690 458876 558696
rect 458180 416220 458232 416226
rect 458180 416162 458232 416168
rect 457444 410916 457496 410922
rect 457444 410858 457496 410864
rect 458836 410854 458864 558690
rect 459572 416158 459600 558855
rect 460938 558784 460994 558793
rect 460938 558719 460994 558728
rect 460386 558648 460442 558657
rect 460386 558583 460442 558592
rect 460400 557734 460428 558583
rect 460388 557728 460440 557734
rect 460388 557670 460440 557676
rect 460846 557696 460902 557705
rect 460204 557660 460256 557666
rect 460204 557602 460256 557608
rect 459560 416152 459612 416158
rect 459560 416094 459612 416100
rect 458824 410848 458876 410854
rect 458824 410790 458876 410796
rect 460216 410786 460244 557602
rect 460204 410780 460256 410786
rect 460204 410722 460256 410728
rect 460400 410718 460428 557670
rect 460846 557631 460848 557640
rect 460900 557631 460902 557640
rect 460848 557602 460900 557608
rect 460388 410712 460440 410718
rect 460388 410654 460440 410660
rect 460952 410650 460980 558719
rect 461044 416090 461072 558855
rect 461688 558550 461716 558855
rect 461676 558544 461728 558550
rect 461676 558486 461728 558492
rect 461032 416084 461084 416090
rect 461032 416026 461084 416032
rect 460940 410644 460992 410650
rect 460940 410586 460992 410592
rect 462332 410582 462360 558855
rect 463054 558784 463110 558793
rect 463054 558719 463110 558728
rect 463068 558618 463096 558719
rect 463056 558612 463108 558618
rect 463056 558554 463108 558560
rect 463712 412078 463740 558855
rect 464250 558784 464306 558793
rect 464250 558719 464306 558728
rect 464264 558482 464292 558719
rect 464252 558476 464304 558482
rect 464252 558418 464304 558424
rect 464344 557592 464396 557598
rect 464344 557534 464396 557540
rect 464356 430574 464384 557534
rect 464344 430568 464396 430574
rect 464344 430510 464396 430516
rect 463700 412072 463752 412078
rect 463700 412014 463752 412020
rect 465092 411942 465120 558855
rect 465262 558784 465318 558793
rect 465262 558719 465318 558728
rect 465276 558686 465304 558719
rect 465264 558680 465316 558686
rect 465264 558622 465316 558628
rect 465724 485920 465776 485926
rect 465724 485862 465776 485868
rect 465736 412690 465764 485862
rect 465724 412684 465776 412690
rect 465724 412626 465776 412632
rect 465080 411936 465132 411942
rect 465080 411878 465132 411884
rect 466472 411262 466500 558855
rect 466552 558816 466604 558822
rect 466550 558784 466552 558793
rect 466604 558784 466606 558793
rect 466550 558719 466606 558728
rect 467104 485852 467156 485858
rect 467104 485794 467156 485800
rect 467116 412758 467144 485794
rect 467104 412752 467156 412758
rect 467104 412694 467156 412700
rect 467852 412146 467880 558855
rect 468758 558855 468814 558864
rect 469218 558920 469274 558929
rect 469218 558855 469274 558864
rect 470598 558920 470654 558929
rect 470598 558855 470654 558864
rect 471978 558920 472034 558929
rect 471978 558855 472034 558864
rect 473358 558920 473414 558929
rect 473358 558855 473414 558864
rect 474738 558920 474794 558929
rect 474738 558855 474794 558864
rect 475474 558920 475530 558929
rect 475474 558855 475530 558864
rect 476118 558920 476174 558929
rect 476118 558855 476174 558864
rect 476578 558920 476634 558929
rect 476578 558855 476580 558864
rect 468024 558826 468076 558832
rect 467930 558784 467986 558793
rect 468036 558754 468064 558826
rect 468772 558754 468800 558855
rect 467930 558719 467986 558728
rect 468024 558748 468076 558754
rect 467944 414798 467972 558719
rect 468024 558690 468076 558696
rect 468116 558748 468168 558754
rect 468116 558690 468168 558696
rect 468760 558748 468812 558754
rect 468760 558690 468812 558696
rect 468036 558657 468064 558690
rect 468022 558648 468078 558657
rect 468022 558583 468078 558592
rect 468128 557734 468156 558690
rect 468116 557728 468168 557734
rect 468116 557670 468168 557676
rect 467932 414792 467984 414798
rect 467932 414734 467984 414740
rect 469232 414730 469260 558855
rect 470046 558648 470102 558657
rect 470046 558583 470102 558592
rect 470060 557666 470088 558583
rect 470048 557660 470100 557666
rect 470048 557602 470100 557608
rect 470612 415342 470640 558855
rect 471334 558784 471390 558793
rect 471334 558719 471390 558728
rect 471348 558550 471376 558719
rect 471336 558544 471388 558550
rect 471336 558486 471388 558492
rect 470692 466472 470744 466478
rect 470692 466414 470744 466420
rect 470600 415336 470652 415342
rect 470600 415278 470652 415284
rect 469220 414724 469272 414730
rect 469220 414666 469272 414672
rect 469404 413976 469456 413982
rect 470704 413953 470732 466414
rect 471992 415410 472020 558855
rect 472162 558784 472218 558793
rect 472162 558719 472218 558728
rect 472176 558618 472204 558719
rect 472164 558612 472216 558618
rect 472164 558554 472216 558560
rect 473372 416770 473400 558855
rect 473450 558784 473506 558793
rect 473450 558719 473506 558728
rect 473464 558482 473492 558719
rect 473452 558476 473504 558482
rect 473452 558418 473504 558424
rect 473452 467900 473504 467906
rect 473452 467842 473504 467848
rect 473360 416764 473412 416770
rect 473360 416706 473412 416712
rect 471980 415404 472032 415410
rect 471980 415346 472032 415352
rect 469404 413918 469456 413924
rect 470690 413944 470746 413953
rect 468116 413160 468168 413166
rect 468116 413102 468168 413108
rect 468128 412729 468156 413102
rect 469416 412729 469444 413918
rect 470690 413879 470746 413888
rect 471980 413772 472032 413778
rect 471980 413714 472032 413720
rect 471992 412729 472020 413714
rect 468114 412720 468170 412729
rect 468114 412655 468170 412664
rect 469402 412720 469458 412729
rect 469402 412655 469458 412664
rect 471978 412720 472034 412729
rect 471978 412655 472034 412664
rect 467840 412140 467892 412146
rect 467840 412082 467892 412088
rect 466460 411256 466512 411262
rect 466460 411198 466512 411204
rect 462320 410576 462372 410582
rect 462320 410518 462372 410524
rect 473464 410417 473492 467842
rect 474752 418130 474780 558855
rect 475488 558822 475516 558855
rect 475476 558816 475528 558822
rect 474830 558784 474886 558793
rect 475476 558758 475528 558764
rect 474830 558719 474886 558728
rect 474844 558686 474872 558719
rect 474832 558680 474884 558686
rect 474832 558622 474884 558628
rect 474844 557734 474872 558622
rect 474832 557728 474884 557734
rect 474832 557670 474884 557676
rect 474832 469260 474884 469266
rect 474832 469202 474884 469208
rect 474740 418124 474792 418130
rect 474740 418066 474792 418072
rect 474844 413953 474872 469202
rect 476132 419490 476160 558855
rect 476632 558855 476634 558864
rect 477590 558920 477646 558929
rect 477590 558855 477646 558864
rect 478970 558920 479026 558929
rect 478970 558855 479026 558864
rect 480350 558920 480406 558929
rect 480350 558855 480406 558864
rect 476580 558826 476632 558832
rect 476210 558648 476266 558657
rect 476210 558583 476266 558592
rect 476224 558414 476252 558583
rect 476592 558414 476620 558826
rect 477604 558754 477632 558855
rect 477592 558748 477644 558754
rect 477592 558690 477644 558696
rect 476212 558408 476264 558414
rect 476212 558350 476264 558356
rect 476580 558408 476632 558414
rect 476580 558350 476632 558356
rect 477498 558376 477554 558385
rect 477604 558346 477632 558690
rect 478878 558512 478934 558521
rect 478878 558447 478934 558456
rect 477498 558311 477500 558320
rect 477552 558311 477554 558320
rect 477592 558340 477644 558346
rect 477500 558282 477552 558288
rect 477592 558282 477644 558288
rect 478892 558278 478920 558447
rect 478984 558278 479012 558855
rect 480364 558550 480392 558855
rect 484398 558784 484454 558793
rect 484398 558719 484454 558728
rect 484412 558686 484440 558719
rect 484400 558680 484452 558686
rect 481638 558648 481694 558657
rect 484400 558622 484452 558628
rect 481638 558583 481640 558592
rect 481692 558583 481694 558592
rect 481640 558554 481692 558560
rect 480352 558544 480404 558550
rect 480352 558486 480404 558492
rect 481638 558512 481694 558521
rect 481638 558447 481694 558456
rect 483018 558512 483074 558521
rect 483018 558447 483020 558456
rect 480350 558376 480406 558385
rect 480350 558311 480406 558320
rect 478880 558272 478932 558278
rect 478880 558214 478932 558220
rect 478972 558272 479024 558278
rect 478972 558214 479024 558220
rect 478984 557666 479012 558214
rect 480364 558210 480392 558311
rect 480352 558204 480404 558210
rect 480352 558146 480404 558152
rect 481652 558074 481680 558447
rect 483072 558447 483074 558456
rect 485778 558512 485834 558521
rect 485778 558447 485834 558456
rect 487158 558512 487214 558521
rect 487158 558447 487214 558456
rect 483020 558418 483072 558424
rect 485792 558414 485820 558447
rect 485780 558408 485832 558414
rect 485780 558350 485832 558356
rect 487172 558346 487200 558447
rect 488538 558376 488594 558385
rect 487160 558340 487212 558346
rect 488538 558311 488594 558320
rect 487160 558282 487212 558288
rect 488552 558278 488580 558311
rect 488540 558272 488592 558278
rect 483018 558240 483074 558249
rect 488540 558214 488592 558220
rect 483018 558175 483074 558184
rect 483032 558142 483060 558175
rect 483020 558136 483072 558142
rect 483020 558078 483072 558084
rect 484398 558104 484454 558113
rect 481640 558068 481692 558074
rect 484398 558039 484454 558048
rect 481640 558010 481692 558016
rect 484412 558006 484440 558039
rect 484400 558000 484452 558006
rect 483018 557968 483074 557977
rect 484400 557942 484452 557948
rect 485778 557968 485834 557977
rect 483018 557903 483020 557912
rect 483072 557903 483074 557912
rect 485778 557903 485834 557912
rect 483020 557874 483072 557880
rect 485792 557870 485820 557903
rect 485780 557864 485832 557870
rect 483018 557832 483074 557841
rect 485780 557806 485832 557812
rect 487158 557832 487214 557841
rect 483018 557767 483074 557776
rect 487158 557767 487160 557776
rect 483032 557734 483060 557767
rect 487212 557767 487214 557776
rect 487160 557738 487212 557744
rect 483020 557728 483072 557734
rect 483020 557670 483072 557676
rect 488538 557696 488594 557705
rect 478972 557660 479024 557666
rect 488538 557631 488594 557640
rect 478972 557602 479024 557608
rect 488552 557598 488580 557631
rect 488540 557592 488592 557598
rect 488540 557534 488592 557540
rect 498844 495508 498896 495514
rect 498844 495450 498896 495456
rect 496084 494080 496136 494086
rect 496084 494022 496136 494028
rect 491944 492788 491996 492794
rect 491944 492730 491996 492736
rect 489184 491360 489236 491366
rect 489184 491302 489236 491308
rect 483664 490000 483716 490006
rect 483664 489942 483716 489948
rect 482284 488572 482336 488578
rect 482284 488514 482336 488520
rect 480904 487212 480956 487218
rect 480904 487154 480956 487160
rect 477592 472048 477644 472054
rect 477592 471990 477644 471996
rect 476120 419484 476172 419490
rect 476120 419426 476172 419432
rect 477604 413953 477632 471990
rect 474830 413944 474886 413953
rect 477590 413944 477646 413953
rect 474830 413879 474886 413888
rect 476120 413908 476172 413914
rect 477590 413879 477646 413888
rect 476120 413850 476172 413856
rect 476132 413817 476160 413850
rect 477500 413840 477552 413846
rect 476118 413808 476174 413817
rect 476118 413743 476174 413752
rect 477498 413808 477500 413817
rect 477552 413808 477554 413817
rect 477498 413743 477554 413752
rect 478880 413704 478932 413710
rect 478878 413672 478880 413681
rect 478932 413672 478934 413681
rect 480916 413642 480944 487154
rect 482296 413710 482324 488514
rect 483676 413846 483704 489942
rect 485044 489932 485096 489938
rect 485044 489874 485096 489880
rect 483664 413840 483716 413846
rect 483664 413782 483716 413788
rect 482284 413704 482336 413710
rect 482284 413646 482336 413652
rect 478878 413607 478934 413616
rect 480444 413636 480496 413642
rect 480444 413578 480496 413584
rect 480904 413636 480956 413642
rect 480904 413578 480956 413584
rect 480456 413545 480484 413578
rect 480442 413536 480498 413545
rect 480442 413471 480498 413480
rect 483020 413500 483072 413506
rect 483020 413442 483072 413448
rect 481640 413432 481692 413438
rect 481638 413400 481640 413409
rect 483032 413409 483060 413442
rect 485056 413438 485084 489874
rect 489196 413914 489224 491302
rect 489184 413908 489236 413914
rect 489184 413850 489236 413856
rect 491956 413778 491984 492730
rect 493324 492720 493376 492726
rect 493324 492662 493376 492668
rect 491944 413772 491996 413778
rect 491944 413714 491996 413720
rect 485780 413568 485832 413574
rect 485778 413536 485780 413545
rect 485832 413536 485834 413545
rect 493336 413506 493364 492662
rect 496096 413982 496124 494022
rect 496084 413976 496136 413982
rect 496084 413918 496136 413924
rect 498856 413710 498884 495450
rect 526352 463752 526404 463758
rect 526352 463694 526404 463700
rect 505100 413976 505152 413982
rect 505100 413918 505152 413924
rect 502524 413908 502576 413914
rect 502524 413850 502576 413856
rect 499580 413840 499632 413846
rect 499580 413782 499632 413788
rect 498292 413704 498344 413710
rect 498292 413646 498344 413652
rect 498844 413704 498896 413710
rect 498844 413646 498896 413652
rect 496820 413636 496872 413642
rect 496820 413578 496872 413584
rect 485778 413471 485834 413480
rect 493324 413500 493376 413506
rect 493324 413442 493376 413448
rect 485044 413432 485096 413438
rect 481692 413400 481694 413409
rect 481638 413335 481694 413344
rect 483018 413400 483074 413409
rect 485044 413374 485096 413380
rect 483018 413335 483074 413344
rect 484400 413364 484452 413370
rect 484400 413306 484452 413312
rect 484412 413273 484440 413306
rect 488540 413296 488592 413302
rect 484398 413264 484454 413273
rect 488538 413264 488540 413273
rect 488592 413264 488594 413273
rect 484398 413199 484454 413208
rect 487160 413228 487212 413234
rect 488538 413199 488594 413208
rect 487160 413170 487212 413176
rect 487172 413137 487200 413170
rect 487158 413128 487214 413137
rect 487158 413063 487214 413072
rect 489920 413092 489972 413098
rect 489920 413034 489972 413040
rect 489932 413001 489960 413034
rect 491300 413024 491352 413030
rect 489918 412992 489974 413001
rect 489918 412927 489974 412936
rect 491298 412992 491300 413001
rect 491352 412992 491354 413001
rect 491298 412927 491354 412936
rect 491392 412956 491444 412962
rect 491392 412898 491444 412904
rect 491404 412729 491432 412898
rect 492680 412888 492732 412894
rect 492680 412830 492732 412836
rect 492692 412729 492720 412830
rect 495716 412752 495768 412758
rect 491390 412720 491446 412729
rect 491390 412655 491446 412664
rect 492678 412720 492734 412729
rect 492678 412655 492734 412664
rect 494058 412720 494114 412729
rect 494058 412655 494060 412664
rect 494112 412655 494114 412664
rect 495714 412720 495716 412729
rect 496832 412729 496860 413578
rect 498304 412729 498332 413646
rect 499592 412729 499620 413782
rect 501052 413432 501104 413438
rect 501052 413374 501104 413380
rect 501064 412729 501092 413374
rect 502536 412729 502564 413850
rect 505112 413817 505140 413918
rect 505098 413808 505154 413817
rect 503720 413772 503772 413778
rect 505098 413743 505154 413752
rect 503720 413714 503772 413720
rect 503732 412729 503760 413714
rect 506480 413704 506532 413710
rect 506478 413672 506480 413681
rect 506532 413672 506534 413681
rect 506478 413607 506534 413616
rect 503996 413500 504048 413506
rect 503996 413442 504048 413448
rect 504008 412729 504036 413442
rect 517520 412820 517572 412826
rect 517520 412762 517572 412768
rect 517532 412729 517560 412762
rect 495768 412720 495770 412729
rect 495714 412655 495770 412664
rect 496818 412720 496874 412729
rect 496818 412655 496874 412664
rect 498290 412720 498346 412729
rect 498290 412655 498346 412664
rect 499578 412720 499634 412729
rect 499578 412655 499634 412664
rect 501050 412720 501106 412729
rect 501050 412655 501106 412664
rect 502522 412720 502578 412729
rect 502522 412655 502578 412664
rect 503718 412720 503774 412729
rect 503718 412655 503774 412664
rect 503994 412720 504050 412729
rect 503994 412655 504050 412664
rect 517518 412720 517574 412729
rect 517518 412655 517574 412664
rect 494060 412626 494112 412632
rect 473450 410408 473506 410417
rect 473450 410343 473506 410352
rect 526364 409986 526392 463694
rect 526442 410000 526498 410009
rect 526364 409958 526442 409986
rect 526442 409935 526498 409944
rect 343640 318776 343692 318782
rect 343638 318744 343640 318753
rect 420184 318776 420236 318782
rect 343692 318744 343694 318753
rect 453120 318776 453172 318782
rect 420184 318718 420236 318724
rect 453118 318744 453120 318753
rect 453172 318744 453174 318753
rect 343638 318679 343694 318688
rect 453118 318679 453174 318688
rect 343652 318102 343680 318679
rect 343640 318096 343692 318102
rect 343640 318038 343692 318044
rect 278778 4856 278834 4865
rect 274640 4820 274692 4826
rect 278778 4791 278834 4800
rect 274640 4762 274692 4768
rect 262220 3460 262272 3466
rect 262220 3402 262272 3408
rect 204260 3334 204312 3340
rect 259458 3360 259514 3369
rect 200120 3324 200172 3330
rect 259458 3295 259514 3304
rect 200120 3266 200172 3272
rect 198740 3256 198792 3262
rect 198740 3198 198792 3204
rect 186320 3188 186372 3194
rect 186320 3130 186372 3136
rect 183560 3120 183612 3126
rect 183560 3062 183612 3068
rect 175280 3052 175332 3058
rect 175280 2994 175332 3000
rect 171140 2984 171192 2990
rect 171140 2926 171192 2932
rect 162860 2848 162912 2854
rect 162860 2790 162912 2796
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 13606 -960 13718 480
rect 14802 -960 14914 480
rect 15998 -960 16110 480
rect 17194 -960 17306 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 27866 -960 27978 480
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44518 -960 44630 480
rect 45714 -960 45826 480
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49302 -960 49414 480
rect 50498 -960 50610 480
rect 51602 -960 51714 480
rect 52798 -960 52910 480
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 56386 -960 56498 480
rect 57582 -960 57694 480
rect 58778 -960 58890 480
rect 59974 -960 60086 480
rect 61170 -960 61282 480
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64758 -960 64870 480
rect 65954 -960 66066 480
rect 67150 -960 67262 480
rect 68254 -960 68366 480
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 73038 -960 73150 480
rect 74234 -960 74346 480
rect 75430 -960 75542 480
rect 76626 -960 76738 480
rect 77822 -960 77934 480
rect 79018 -960 79130 480
rect 80214 -960 80326 480
rect 81410 -960 81522 480
rect 82606 -960 82718 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 88494 -960 88606 480
rect 89690 -960 89802 480
rect 90886 -960 90998 480
rect 92082 -960 92194 480
rect 93278 -960 93390 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 107538 -960 107650 480
rect 108734 -960 108846 480
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 151514 -960 151626 480
rect 152710 -960 152822 480
rect 153906 -960 154018 480
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157494 -960 157606 480
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 162278 -960 162390 480
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 189602 -960 189714 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197974 -960 198086 480
rect 199170 -960 199282 480
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246734 -960 246846 480
rect 247930 -960 248042 480
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 252622 -960 252734 480
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259798 -960 259910 480
rect 260994 -960 261106 480
rect 262190 -960 262302 480
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 268078 -960 268190 480
rect 269274 -960 269386 480
rect 270470 -960 270582 480
rect 271666 -960 271778 480
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 280038 -960 280150 480
rect 281234 -960 281346 480
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 289514 -960 289626 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436990 -960 437102 480
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441774 -960 441886 480
rect 442970 -960 443082 480
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 459622 -960 459734 480
rect 460818 -960 460930 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509578 -960 509690 480
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528622 -960 528734 480
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 569010 -960 569122 480
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 135074 651072 135130 651128
rect 137650 649655 137706 649711
rect 57886 646040 57942 646096
rect 57794 644952 57850 645008
rect 57702 643184 57758 643240
rect 57610 641960 57666 642016
rect 57518 640328 57574 640384
rect 57426 639240 57482 639296
rect 57334 637608 57390 637664
rect 57242 579672 57298 579728
rect 378138 652876 378140 652896
rect 378140 652876 378192 652896
rect 378192 652876 378194 652896
rect 378138 652840 378194 652876
rect 383566 652876 383568 652896
rect 383568 652876 383620 652896
rect 383620 652876 383622 652896
rect 383566 652840 383622 652876
rect 508410 652860 508466 652896
rect 508410 652840 508412 652860
rect 508412 652840 508464 652860
rect 508464 652840 508466 652860
rect 513378 652860 513434 652896
rect 513378 652840 513380 652860
rect 513380 652840 513432 652860
rect 513432 652840 513434 652860
rect 258538 651616 258594 651672
rect 263598 651616 263654 651672
rect 266634 649848 266690 649904
rect 387154 649848 387210 649904
rect 389178 649848 389234 649904
rect 188342 646040 188398 646096
rect 307390 646040 307446 646096
rect 139398 589600 139454 589656
rect 67546 558864 67602 558920
rect 68926 558864 68982 558920
rect 70306 558864 70362 558920
rect 71686 558864 71742 558920
rect 72514 558864 72570 558920
rect 73066 558864 73122 558920
rect 73710 558864 73766 558920
rect 74262 558864 74318 558920
rect 74998 558864 75054 558920
rect 75826 558864 75882 558920
rect 76838 558864 76894 558920
rect 77390 558884 77446 558920
rect 77390 558864 77392 558884
rect 77392 558864 77444 558884
rect 77444 558864 77446 558884
rect 62026 558320 62082 558376
rect 63406 558184 63462 558240
rect 70214 558592 70270 558648
rect 75918 558612 75974 558648
rect 75918 558592 75920 558612
rect 75920 558592 75972 558612
rect 75972 558592 75974 558612
rect 78586 558864 78642 558920
rect 79322 558864 79378 558920
rect 79874 558864 79930 558920
rect 80794 558864 80850 558920
rect 81254 558864 81310 558920
rect 81990 558864 82046 558920
rect 82910 558864 82966 558920
rect 83830 558864 83886 558920
rect 84198 558864 84254 558920
rect 85486 558864 85542 558920
rect 86314 558884 86370 558920
rect 86314 558864 86316 558884
rect 86316 558864 86368 558884
rect 86368 558864 86370 558884
rect 78494 558628 78496 558648
rect 78496 558628 78548 558648
rect 78548 558628 78550 558648
rect 78494 558592 78550 558628
rect 79414 558592 79470 558648
rect 85394 558612 85450 558648
rect 85394 558592 85396 558612
rect 85396 558592 85448 558612
rect 85448 558592 85450 558612
rect 82726 557912 82782 557968
rect 77574 542952 77630 543008
rect 86774 558864 86830 558920
rect 87878 558864 87934 558920
rect 88246 558864 88302 558920
rect 88890 558864 88946 558920
rect 89166 558864 89222 558920
rect 89810 558864 89866 558920
rect 91006 558864 91062 558920
rect 92202 558864 92258 558920
rect 92478 558864 92534 558920
rect 93306 558864 93362 558920
rect 93766 558884 93822 558920
rect 93766 558864 93768 558884
rect 93768 558864 93820 558884
rect 93820 558864 93822 558884
rect 86866 558592 86922 558648
rect 91098 558592 91154 558648
rect 95054 558864 95110 558920
rect 95698 558864 95754 558920
rect 96526 558864 96582 558920
rect 97170 558864 97226 558920
rect 97814 558864 97870 558920
rect 98366 558864 98422 558920
rect 99286 558864 99342 558920
rect 100022 558864 100078 558920
rect 102046 558864 102102 558920
rect 104806 558864 104862 558920
rect 107290 558864 107346 558920
rect 108486 558864 108542 558920
rect 93674 558592 93730 558648
rect 94778 558592 94834 558648
rect 96250 543224 96306 543280
rect 99470 558456 99526 558512
rect 100390 558456 100446 558512
rect 100022 557660 100078 557696
rect 100850 557796 100906 557832
rect 100850 557776 100852 557796
rect 100852 557776 100904 557796
rect 100904 557776 100906 557796
rect 101402 557776 101458 557832
rect 100022 557640 100024 557660
rect 100024 557640 100076 557660
rect 100076 557640 100078 557660
rect 106278 558592 106334 558648
rect 108486 558456 108542 558512
rect 110326 558456 110382 558512
rect 108302 557912 108358 557968
rect 106922 557640 106978 557696
rect 102046 557504 102102 557560
rect 102782 557504 102838 557560
rect 103426 557504 103482 557560
rect 104162 557504 104218 557560
rect 105542 557504 105598 557560
rect 106186 557504 106242 557560
rect 103426 543088 103482 543144
rect 140042 543632 140098 543688
rect 141422 543360 141478 543416
rect 148322 543496 148378 543552
rect 188434 644952 188490 645008
rect 188526 643184 188582 643240
rect 188618 641960 188674 642016
rect 188710 640328 188766 640384
rect 188802 639240 188858 639296
rect 188894 637608 188950 637664
rect 269118 589328 269174 589384
rect 269118 587152 269174 587208
rect 270406 580352 270462 580408
rect 188986 579672 189042 579728
rect 188342 543224 188398 543280
rect 210974 559952 211030 560008
rect 195978 558864 196034 558920
rect 200210 558864 200266 558920
rect 202786 558864 202842 558920
rect 203798 558864 203854 558920
rect 204166 558864 204222 558920
rect 205546 558864 205602 558920
rect 206926 558864 206982 558920
rect 208490 558864 208546 558920
rect 210606 558864 210662 558920
rect 194414 558728 194470 558784
rect 188986 542952 189042 543008
rect 202142 558592 202198 558648
rect 201498 557640 201554 557696
rect 200026 543632 200082 543688
rect 202050 543088 202106 543144
rect 204902 558592 204958 558648
rect 209042 558592 209098 558648
rect 207662 557640 207718 557696
rect 206926 557504 206982 557560
rect 208306 557504 208362 557560
rect 209686 557504 209742 557560
rect 210422 543496 210478 543552
rect 208306 543360 208362 543416
rect 211802 558864 211858 558920
rect 213182 558864 213238 558920
rect 214010 558864 214066 558920
rect 215298 558864 215354 558920
rect 217506 558864 217562 558920
rect 218794 558864 218850 558920
rect 220082 558864 220138 558920
rect 221094 558864 221150 558920
rect 222198 558864 222254 558920
rect 224498 558864 224554 558920
rect 225878 558864 225934 558920
rect 226154 558864 226210 558920
rect 227166 558864 227222 558920
rect 227626 558864 227682 558920
rect 227994 558864 228050 558920
rect 229006 558864 229062 558920
rect 229466 558864 229522 558920
rect 230386 558864 230442 558920
rect 231766 558864 231822 558920
rect 233054 558864 233110 558920
rect 233238 558864 233294 558920
rect 234526 558864 234582 558920
rect 235906 558864 235962 558920
rect 237286 558864 237342 558920
rect 240046 558864 240102 558920
rect 211066 557640 211122 557696
rect 217598 558728 217654 558784
rect 223578 558728 223634 558784
rect 217966 557640 218022 557696
rect 212446 557504 212502 557560
rect 213826 557504 213882 557560
rect 215206 557504 215262 557560
rect 216586 557504 216642 557560
rect 217874 557504 217930 557560
rect 219346 557504 219402 557560
rect 220726 557504 220782 557560
rect 222106 557504 222162 557560
rect 223486 557504 223542 557560
rect 224866 557504 224922 557560
rect 226246 558728 226302 558784
rect 230478 558340 230534 558376
rect 230478 558320 230480 558340
rect 230480 558320 230532 558340
rect 230532 558320 230534 558340
rect 231858 558728 231914 558784
rect 231858 558456 231914 558512
rect 233146 558728 233202 558784
rect 234618 558728 234674 558784
rect 235998 558728 236054 558784
rect 237378 558748 237434 558784
rect 237378 558728 237380 558748
rect 237380 558728 237432 558748
rect 237432 558728 237434 558748
rect 238758 558320 238814 558376
rect 238666 558048 238722 558104
rect 281538 578992 281594 579048
rect 281446 440952 281502 441008
rect 281446 429936 281502 429992
rect 282274 539416 282330 539472
rect 282826 538464 282882 538520
rect 282826 537376 282882 537432
rect 282826 536424 282882 536480
rect 281722 535336 281778 535392
rect 282090 534384 282146 534440
rect 282090 533432 282146 533488
rect 282274 532344 282330 532400
rect 282826 531392 282882 531448
rect 282826 530304 282882 530360
rect 282826 529352 282882 529408
rect 282274 528264 282330 528320
rect 282826 527312 282882 527368
rect 281906 526360 281962 526416
rect 282826 525272 282882 525328
rect 282366 524320 282422 524376
rect 282826 523232 282882 523288
rect 282826 522280 282882 522336
rect 283562 521192 283618 521248
rect 282826 520276 282828 520296
rect 282828 520276 282880 520296
rect 282880 520276 282882 520296
rect 282826 520240 282882 520276
rect 281722 519288 281778 519344
rect 282090 518200 282146 518256
rect 282274 517248 282330 517304
rect 282826 516180 282882 516216
rect 282826 516160 282828 516180
rect 282828 516160 282880 516180
rect 282880 516160 282882 516180
rect 282826 515208 282882 515264
rect 282274 514256 282330 514312
rect 282734 513168 282790 513224
rect 282826 512216 282882 512272
rect 281722 511128 281778 511184
rect 282274 510176 282330 510232
rect 282550 509088 282606 509144
rect 282826 508136 282882 508192
rect 282090 507184 282146 507240
rect 282734 506096 282790 506152
rect 282826 505180 282828 505200
rect 282828 505180 282880 505200
rect 282880 505180 282882 505200
rect 282826 505144 282882 505180
rect 282826 504056 282882 504112
rect 282826 503104 282882 503160
rect 282274 502016 282330 502072
rect 282826 501084 282882 501120
rect 282826 501064 282828 501084
rect 282828 501064 282880 501084
rect 282880 501064 282882 501084
rect 282826 499024 282882 499080
rect 282826 496984 282882 497040
rect 281906 496032 281962 496088
rect 282826 495080 282882 495136
rect 282366 493992 282422 494048
rect 282826 493040 282882 493096
rect 282826 491952 282882 492008
rect 282274 491000 282330 491056
rect 282826 489948 282828 489968
rect 282828 489948 282880 489968
rect 282880 489948 282882 489968
rect 282826 489912 282882 489948
rect 282274 488960 282330 489016
rect 282826 488008 282882 488064
rect 282274 486920 282330 486976
rect 282826 485968 282882 486024
rect 281722 484880 281778 484936
rect 282274 483928 282330 483984
rect 282550 482840 282606 482896
rect 282826 481888 282882 481944
rect 282090 480936 282146 480992
rect 282734 479848 282790 479904
rect 282826 478932 282828 478952
rect 282828 478932 282880 478952
rect 282880 478932 282882 478952
rect 282826 478896 282882 478932
rect 282826 477808 282882 477864
rect 282090 476856 282146 476912
rect 282274 475768 282330 475824
rect 282826 474836 282882 474872
rect 282826 474816 282828 474836
rect 282828 474816 282880 474836
rect 282880 474816 282882 474836
rect 281722 473864 281778 473920
rect 282090 472776 282146 472832
rect 282734 471824 282790 471880
rect 282826 470736 282882 470792
rect 281906 469784 281962 469840
rect 282826 468832 282882 468888
rect 282734 467744 282790 467800
rect 282826 466792 282882 466848
rect 282826 465704 282882 465760
rect 282734 464752 282790 464808
rect 282826 463700 282828 463720
rect 282828 463700 282880 463720
rect 282880 463700 282882 463720
rect 282826 463664 282882 463700
rect 282826 462712 282882 462768
rect 282826 461760 282882 461816
rect 282826 460672 282882 460728
rect 282734 459720 282790 459776
rect 281722 458632 281778 458688
rect 282090 457680 282146 457736
rect 281630 456592 281686 456648
rect 282826 455640 282882 455696
rect 281630 454688 281686 454744
rect 282458 453600 282514 453656
rect 282274 452648 282330 452704
rect 282090 446528 282146 446584
rect 281814 445576 281870 445632
rect 281722 442584 281778 442640
rect 281998 444488 282054 444544
rect 281906 443536 281962 443592
rect 282182 440544 282238 440600
rect 282182 439456 282238 439512
rect 282182 437416 282238 437472
rect 282182 436464 282238 436520
rect 282182 435512 282238 435568
rect 282182 434424 282238 434480
rect 282182 432384 282238 432440
rect 282366 451560 282422 451616
rect 282274 431432 282330 431488
rect 282274 429392 282330 429448
rect 282274 428440 282330 428496
rect 282274 427352 282330 427408
rect 282274 426944 282330 427000
rect 282274 425312 282330 425368
rect 282274 424360 282330 424416
rect 282274 423408 282330 423464
rect 282274 422320 282330 422376
rect 282274 421368 282330 421424
rect 282550 450608 282606 450664
rect 282826 449656 282882 449712
rect 282642 448568 282698 448624
rect 282274 414296 282330 414352
rect 282550 418240 282606 418296
rect 282734 447616 282790 447672
rect 283470 438504 283526 438560
rect 283378 433472 283434 433528
rect 282826 420280 282882 420336
rect 282826 419364 282828 419384
rect 282828 419364 282880 419384
rect 282880 419364 282882 419384
rect 282826 419328 282882 419364
rect 282826 417288 282882 417344
rect 282826 416336 282882 416392
rect 282826 415248 282882 415304
rect 282826 413208 282882 413264
rect 282826 412256 282882 412312
rect 281722 409264 281778 409320
rect 281722 408176 281778 408232
rect 281630 403144 281686 403200
rect 281630 398148 281632 398168
rect 281632 398148 281684 398168
rect 281684 398148 281686 398168
rect 281630 398112 281686 398148
rect 281630 397196 281632 397216
rect 281632 397196 281684 397216
rect 281684 397196 281686 397216
rect 281630 397160 281686 397196
rect 281630 396072 281686 396128
rect 281630 395120 281686 395176
rect 281630 394032 281686 394088
rect 281630 393080 281686 393136
rect 281630 392028 281632 392048
rect 281632 392028 281684 392048
rect 281684 392028 281686 392048
rect 281630 391992 281686 392028
rect 281630 391040 281686 391096
rect 281630 390124 281632 390144
rect 281632 390124 281684 390144
rect 281684 390124 281686 390144
rect 281630 390088 281686 390124
rect 281630 389036 281632 389056
rect 281632 389036 281684 389056
rect 281684 389036 281686 389056
rect 281630 389000 281686 389036
rect 281630 388048 281686 388104
rect 281630 386960 281686 387016
rect 281630 386044 281632 386064
rect 281632 386044 281684 386064
rect 281684 386044 281686 386064
rect 281630 386008 281686 386044
rect 281630 385056 281686 385112
rect 281630 384004 281632 384024
rect 281632 384004 281684 384024
rect 281684 384004 281686 384024
rect 281630 383968 281686 384004
rect 281630 383016 281686 383072
rect 281630 381928 281686 381984
rect 281630 379888 281686 379944
rect 281630 378936 281686 378992
rect 281630 377984 281686 378040
rect 281630 375944 281686 376000
rect 281630 374856 281686 374912
rect 281630 373904 281686 373960
rect 281630 371900 281632 371920
rect 281632 371900 281684 371920
rect 281684 371900 281686 371920
rect 281630 371864 281686 371900
rect 281630 370948 281632 370968
rect 281632 370948 281684 370968
rect 281684 370948 281686 370968
rect 281630 370912 281686 370948
rect 281630 368872 281686 368928
rect 281630 367784 281686 367840
rect 281630 364792 281686 364848
rect 281630 363840 281686 363896
rect 281630 362752 281686 362808
rect 281630 360712 281686 360768
rect 281630 359760 281686 359816
rect 281630 357720 281686 357776
rect 281630 351772 281632 351792
rect 281632 351772 281684 351792
rect 281684 351772 281686 351792
rect 281630 351736 281686 351772
rect 281630 350648 281686 350704
rect 281630 349696 281686 349752
rect 281630 348608 281686 348664
rect 281630 347692 281632 347712
rect 281632 347692 281684 347712
rect 281684 347692 281686 347712
rect 281630 347656 281686 347692
rect 281630 346568 281686 346624
rect 281630 345652 281632 345672
rect 281632 345652 281684 345672
rect 281684 345652 281686 345672
rect 281630 345616 281686 345652
rect 281630 344664 281686 344720
rect 281630 343596 281686 343632
rect 281630 343576 281632 343596
rect 281632 343576 281684 343596
rect 281684 343576 281686 343596
rect 281630 341536 281686 341592
rect 282826 411188 282882 411224
rect 282826 411168 282828 411188
rect 282828 411168 282880 411188
rect 282880 411168 282882 411188
rect 282734 410216 282790 410272
rect 282826 407224 282882 407280
rect 282366 406136 282422 406192
rect 282274 399064 282330 399120
rect 281814 380976 281870 381032
rect 281814 376896 281870 376952
rect 281814 372816 281870 372872
rect 281814 369824 281870 369880
rect 281814 361800 281870 361856
rect 281814 358808 281870 358864
rect 282274 354728 282330 354784
rect 282826 405184 282882 405240
rect 282826 404232 282882 404288
rect 283562 413616 283618 413672
rect 283378 413344 283434 413400
rect 283746 413480 283802 413536
rect 283930 413208 283986 413264
rect 282826 402228 282828 402248
rect 282828 402228 282880 402248
rect 282880 402228 282882 402248
rect 282826 402192 282882 402228
rect 282826 401140 282828 401160
rect 282828 401140 282880 401160
rect 282880 401140 282882 401160
rect 282826 401104 282882 401140
rect 282826 400172 282882 400208
rect 282826 400152 282828 400172
rect 282828 400152 282880 400172
rect 282880 400152 282882 400172
rect 284482 366832 284538 366888
rect 282642 356768 282698 356824
rect 282550 355680 282606 355736
rect 282458 353640 282514 353696
rect 282366 352688 282422 352744
rect 281814 342624 281870 342680
rect 281630 340584 281686 340640
rect 281722 339632 281778 339688
rect 281630 338544 281686 338600
rect 281630 337592 281686 337648
rect 281630 336540 281632 336560
rect 281632 336540 281684 336560
rect 281684 336540 281686 336560
rect 281630 336504 281686 336540
rect 281722 335552 281778 335608
rect 281630 334464 281686 334520
rect 281630 333512 281686 333568
rect 281722 332560 281778 332616
rect 281906 331472 281962 331528
rect 281630 330520 281686 330576
rect 281538 329432 281594 329488
rect 281630 328480 281686 328536
rect 281538 327392 281594 327448
rect 281538 325524 281540 325544
rect 281540 325524 281592 325544
rect 281592 325524 281594 325544
rect 281538 325488 281594 325524
rect 282366 326440 282422 326496
rect 285126 365744 285182 365800
rect 287058 413344 287114 413400
rect 287150 413208 287206 413264
rect 287058 413072 287114 413128
rect 287058 412972 287060 412992
rect 287060 412972 287112 412992
rect 287112 412972 287114 412992
rect 287058 412936 287114 412972
rect 287150 412800 287206 412856
rect 307114 644952 307170 645008
rect 307114 643456 307170 643512
rect 307666 642096 307722 642152
rect 307666 640464 307722 640520
rect 307022 639240 307078 639296
rect 306838 637880 306894 637936
rect 296626 413344 296682 413400
rect 296534 413208 296590 413264
rect 296626 413072 296682 413128
rect 296626 412972 296628 412992
rect 296628 412972 296680 412992
rect 296680 412972 296682 412992
rect 296626 412936 296682 412972
rect 296534 412800 296590 412856
rect 306378 413344 306434 413400
rect 306470 413208 306526 413264
rect 306378 413072 306434 413128
rect 306378 412972 306380 412992
rect 306380 412972 306432 412992
rect 306432 412972 306434 412992
rect 306378 412936 306434 412972
rect 306470 412800 306526 412856
rect 307666 579808 307722 579864
rect 348422 559272 348478 559328
rect 358174 559272 358230 559328
rect 313830 558900 313832 558920
rect 313832 558900 313884 558920
rect 313884 558900 313886 558920
rect 313830 558864 313886 558900
rect 317418 558864 317474 558920
rect 318798 558864 318854 558920
rect 320178 558864 320234 558920
rect 325698 558864 325754 558920
rect 327078 558864 327134 558920
rect 329286 558864 329342 558920
rect 329930 558864 329986 558920
rect 331770 558864 331826 558920
rect 332598 558864 332654 558920
rect 333978 558864 334034 558920
rect 335358 558864 335414 558920
rect 336738 558864 336794 558920
rect 337566 558864 337622 558920
rect 338118 558864 338174 558920
rect 339498 558864 339554 558920
rect 340878 558864 340934 558920
rect 342258 558864 342314 558920
rect 343730 558864 343786 558920
rect 344282 558864 344338 558920
rect 345018 558864 345074 558920
rect 346398 558864 346454 558920
rect 316314 557776 316370 557832
rect 315946 413344 316002 413400
rect 315854 413208 315910 413264
rect 315946 413072 316002 413128
rect 315946 412972 315948 412992
rect 315948 412972 316000 412992
rect 316000 412972 316002 412992
rect 315946 412936 316002 412972
rect 315854 412800 315910 412856
rect 320270 558728 320326 558784
rect 322202 558728 322258 558784
rect 321558 558048 321614 558104
rect 323582 558592 323638 558648
rect 324962 558592 325018 558648
rect 322938 558068 322994 558104
rect 322938 558048 322940 558068
rect 322940 558048 322992 558068
rect 322992 558048 322994 558068
rect 324318 557660 324374 557696
rect 324318 557640 324320 557660
rect 324320 557640 324372 557660
rect 324372 557640 324374 557660
rect 326342 558728 326398 558784
rect 328458 558728 328514 558784
rect 327722 558592 327778 558648
rect 329102 558592 329158 558648
rect 329838 557932 329894 557968
rect 329838 557912 329840 557932
rect 329840 557912 329892 557932
rect 329892 557912 329894 557932
rect 330482 558728 330538 558784
rect 331218 557796 331274 557832
rect 331218 557776 331220 557796
rect 331220 557776 331272 557796
rect 331272 557776 331274 557796
rect 331126 412972 331128 412992
rect 331128 412972 331180 412992
rect 331180 412972 331182 412992
rect 331126 412936 331182 412972
rect 333150 558728 333206 558784
rect 334070 558728 334126 558784
rect 335266 413344 335322 413400
rect 335174 413208 335230 413264
rect 335266 413072 335322 413128
rect 335266 412972 335268 412992
rect 335268 412972 335320 412992
rect 335320 412972 335322 412992
rect 335266 412936 335322 412972
rect 335174 412800 335230 412856
rect 335450 558728 335506 558784
rect 336646 558728 336702 558784
rect 336830 558728 336886 558784
rect 339038 558728 339094 558784
rect 281722 322360 281778 322416
rect 339866 558728 339922 558784
rect 341246 558728 341302 558784
rect 342534 558728 342590 558784
rect 343638 558728 343694 558784
rect 343638 557640 343694 557696
rect 346030 558728 346086 558784
rect 347778 558864 347834 558920
rect 347686 558728 347742 558784
rect 348238 558728 348294 558784
rect 349158 558864 349214 558920
rect 352010 558864 352066 558920
rect 356058 558884 356114 558920
rect 356058 558864 356060 558884
rect 356060 558864 356112 558884
rect 356112 558864 356114 558884
rect 349710 558728 349766 558784
rect 350538 558456 350594 558512
rect 353298 558728 353354 558784
rect 354678 558728 354734 558784
rect 357438 558476 357494 558512
rect 357438 558456 357440 558476
rect 357440 558456 357492 558476
rect 357492 558456 357494 558476
rect 352102 557640 352158 557696
rect 350630 557504 350686 557560
rect 350446 412972 350448 412992
rect 350448 412972 350500 412992
rect 350500 412972 350502 412992
rect 350446 412936 350502 412972
rect 352010 555464 352066 555520
rect 353298 557504 353354 557560
rect 354678 557504 354734 557560
rect 354126 413752 354182 413808
rect 354586 413344 354642 413400
rect 354494 413208 354550 413264
rect 354586 413072 354642 413128
rect 354586 412972 354588 412992
rect 354588 412972 354640 412992
rect 354640 412972 354642 412992
rect 354586 412936 354642 412972
rect 354494 412800 354550 412856
rect 356150 557504 356206 557560
rect 357530 557504 357586 557560
rect 358910 555464 358966 555520
rect 367098 413888 367154 413944
rect 364338 413344 364394 413400
rect 364338 413072 364394 413128
rect 364338 412800 364394 412856
rect 367098 412684 367154 412720
rect 368570 413888 368626 413944
rect 371882 414024 371938 414080
rect 369950 413888 370006 413944
rect 371238 413888 371294 413944
rect 372618 413888 372674 413944
rect 368294 413072 368350 413128
rect 368478 413072 368534 413128
rect 369858 413072 369914 413128
rect 370962 413072 371018 413128
rect 371330 412800 371386 412856
rect 373906 413344 373962 413400
rect 373998 413208 374054 413264
rect 373906 412936 373962 412992
rect 373998 412800 374054 412856
rect 367098 412664 367100 412684
rect 367100 412664 367152 412684
rect 367152 412664 367154 412684
rect 368294 412664 368350 412720
rect 370962 412664 371018 412720
rect 371238 412700 371240 412720
rect 371240 412700 371292 412720
rect 371292 412700 371294 412720
rect 371238 412664 371294 412700
rect 375378 413208 375434 413264
rect 375562 413208 375618 413264
rect 376758 413208 376814 413264
rect 375470 413072 375526 413128
rect 376758 412800 376814 412856
rect 378230 413208 378286 413264
rect 379610 413888 379666 413944
rect 379794 413344 379850 413400
rect 380622 413752 380678 413808
rect 380990 413344 381046 413400
rect 382278 413344 382334 413400
rect 380622 413208 380678 413264
rect 382186 413072 382242 413128
rect 382370 413072 382426 413128
rect 378138 412800 378194 412856
rect 379610 412800 379666 412856
rect 379794 412800 379850 412856
rect 372618 412664 372674 412720
rect 374182 412664 374238 412720
rect 384302 413752 384358 413808
rect 385314 413480 385370 413536
rect 385038 413072 385094 413128
rect 385314 413072 385370 413128
rect 386418 413480 386474 413536
rect 387890 413888 387946 413944
rect 390650 413888 390706 413944
rect 392030 413888 392086 413944
rect 402978 413924 402980 413944
rect 402980 413924 403032 413944
rect 403032 413924 403034 413944
rect 402978 413888 403034 413924
rect 391938 413788 391940 413808
rect 391940 413788 391992 413808
rect 391992 413788 391994 413808
rect 391938 413752 391994 413788
rect 396078 413752 396134 413808
rect 516414 649848 516470 649904
rect 438122 646040 438178 646096
rect 407762 413888 407818 413944
rect 410522 413888 410578 413944
rect 389178 413480 389234 413536
rect 389362 413480 389418 413536
rect 394698 413516 394700 413536
rect 394700 413516 394752 413536
rect 394752 413516 394754 413536
rect 394698 413480 394754 413516
rect 389086 412936 389142 412992
rect 389270 412936 389326 412992
rect 404358 413480 404414 413536
rect 393226 413344 393282 413400
rect 397458 413380 397460 413400
rect 397460 413380 397512 413400
rect 397512 413380 397514 413400
rect 397458 413344 397514 413380
rect 390558 412936 390614 412992
rect 401598 413344 401654 413400
rect 397550 413072 397606 413128
rect 398838 413072 398894 413128
rect 393318 412936 393374 412992
rect 396078 412936 396134 412992
rect 397458 412972 397460 412992
rect 397460 412972 397512 412992
rect 397512 412972 397514 412992
rect 397458 412936 397514 412972
rect 393226 412800 393282 412856
rect 394698 412836 394700 412856
rect 394700 412836 394752 412856
rect 394752 412836 394754 412856
rect 394698 412800 394754 412836
rect 400218 412820 400274 412856
rect 400218 412800 400220 412820
rect 400220 412800 400272 412820
rect 400272 412800 400274 412820
rect 403162 412800 403218 412856
rect 413926 413888 413982 413944
rect 380898 412664 380954 412720
rect 382278 412664 382334 412720
rect 383658 412664 383714 412720
rect 385038 412684 385094 412720
rect 385038 412664 385040 412684
rect 385040 412664 385092 412684
rect 385092 412664 385094 412684
rect 387062 412664 387118 412720
rect 387798 412664 387854 412720
rect 398838 412700 398840 412720
rect 398840 412700 398892 412720
rect 398892 412700 398894 412720
rect 398838 412664 398894 412700
rect 400218 412684 400274 412720
rect 400218 412664 400220 412684
rect 400220 412664 400272 412684
rect 400272 412664 400274 412684
rect 405738 411440 405794 411496
rect 416778 392944 416834 393000
rect 416410 391312 416466 391368
rect 419906 346568 419962 346624
rect 419814 344392 419870 344448
rect 419722 343712 419778 343768
rect 419630 341672 419686 341728
rect 419538 340992 419594 341048
rect 438214 644952 438270 645008
rect 438306 643184 438362 643240
rect 438398 641960 438454 642016
rect 438490 640328 438546 640384
rect 438582 639240 438638 639296
rect 438674 637608 438730 637664
rect 518898 589328 518954 589384
rect 518898 587696 518954 587752
rect 438766 579672 438822 579728
rect 420182 412800 420238 412856
rect 420090 349152 420146 349208
rect 419998 346432 420054 346488
rect 420090 333648 420146 333704
rect 419998 332016 420054 332072
rect 419906 330928 419962 330984
rect 419814 329160 419870 329216
rect 419722 328072 419778 328128
rect 419630 325760 419686 325816
rect 419538 325080 419594 325136
rect 282826 321408 282882 321464
rect 279330 320864 279386 320920
rect 40958 3848 41014 3904
rect 44546 3984 44602 4040
rect 45742 3712 45798 3768
rect 54022 3576 54078 3632
rect 55310 4120 55366 4176
rect 56414 3440 56470 3496
rect 64786 318552 64842 318608
rect 64694 4120 64750 4176
rect 74446 318416 74502 318472
rect 82634 318280 82690 318336
rect 82726 318144 82782 318200
rect 104806 318008 104862 318064
rect 108762 5480 108818 5536
rect 112350 5344 112406 5400
rect 115938 4800 115994 4856
rect 121826 3304 121882 3360
rect 123482 3984 123538 4040
rect 129002 5208 129058 5264
rect 127806 5072 127862 5128
rect 126978 3848 127034 3904
rect 132590 4936 132646 4992
rect 133142 4800 133198 4856
rect 134890 4800 134946 4856
rect 133878 3712 133934 3768
rect 147678 3576 147734 3632
rect 151818 3440 151874 3496
rect 165986 318552 166042 318608
rect 181534 318416 181590 318472
rect 193218 318280 193274 318336
rect 195150 318144 195206 318200
rect 230202 318008 230258 318064
rect 237378 5480 237434 5536
rect 242898 5344 242954 5400
rect 270498 5208 270554 5264
rect 269118 5072 269174 5128
rect 276018 4936 276074 4992
rect 443090 558864 443146 558920
rect 445758 558864 445814 558920
rect 451278 558864 451334 558920
rect 452658 558864 452714 558920
rect 453670 558864 453726 558920
rect 454038 558864 454094 558920
rect 455418 558864 455474 558920
rect 456798 558864 456854 558920
rect 458178 558864 458234 558920
rect 459558 558864 459614 558920
rect 461030 558864 461086 558920
rect 461674 558864 461730 558920
rect 462318 558864 462374 558920
rect 463698 558864 463754 558920
rect 465078 558864 465134 558920
rect 466458 558864 466514 558920
rect 467838 558864 467894 558920
rect 449898 557776 449954 557832
rect 452750 558728 452806 558784
rect 453302 558592 453358 558648
rect 454774 558748 454830 558784
rect 454774 558728 454776 558748
rect 454776 558728 454828 558748
rect 454828 558728 454830 558748
rect 456062 558728 456118 558784
rect 457442 558764 457444 558784
rect 457444 558764 457496 558784
rect 457496 558764 457498 558784
rect 457442 558728 457498 558764
rect 458822 558748 458878 558784
rect 458822 558728 458824 558748
rect 458824 558728 458876 558748
rect 458876 558728 458878 558748
rect 460938 558728 460994 558784
rect 460386 558592 460442 558648
rect 460846 557660 460902 557696
rect 460846 557640 460848 557660
rect 460848 557640 460900 557660
rect 460900 557640 460902 557660
rect 463054 558728 463110 558784
rect 464250 558728 464306 558784
rect 465262 558728 465318 558784
rect 466550 558764 466552 558784
rect 466552 558764 466604 558784
rect 466604 558764 466606 558784
rect 466550 558728 466606 558764
rect 468758 558864 468814 558920
rect 469218 558864 469274 558920
rect 470598 558864 470654 558920
rect 471978 558864 472034 558920
rect 473358 558864 473414 558920
rect 474738 558864 474794 558920
rect 475474 558864 475530 558920
rect 476118 558864 476174 558920
rect 476578 558884 476634 558920
rect 476578 558864 476580 558884
rect 476580 558864 476632 558884
rect 476632 558864 476634 558884
rect 467930 558728 467986 558784
rect 468022 558592 468078 558648
rect 470046 558592 470102 558648
rect 471334 558728 471390 558784
rect 472162 558728 472218 558784
rect 473450 558728 473506 558784
rect 470690 413888 470746 413944
rect 468114 412664 468170 412720
rect 469402 412664 469458 412720
rect 471978 412664 472034 412720
rect 474830 558728 474886 558784
rect 477590 558864 477646 558920
rect 478970 558864 479026 558920
rect 480350 558864 480406 558920
rect 476210 558592 476266 558648
rect 477498 558340 477554 558376
rect 478878 558456 478934 558512
rect 477498 558320 477500 558340
rect 477500 558320 477552 558340
rect 477552 558320 477554 558340
rect 484398 558728 484454 558784
rect 481638 558612 481694 558648
rect 481638 558592 481640 558612
rect 481640 558592 481692 558612
rect 481692 558592 481694 558612
rect 481638 558456 481694 558512
rect 483018 558476 483074 558512
rect 483018 558456 483020 558476
rect 483020 558456 483072 558476
rect 483072 558456 483074 558476
rect 480350 558320 480406 558376
rect 485778 558456 485834 558512
rect 487158 558456 487214 558512
rect 488538 558320 488594 558376
rect 483018 558184 483074 558240
rect 484398 558048 484454 558104
rect 483018 557932 483074 557968
rect 483018 557912 483020 557932
rect 483020 557912 483072 557932
rect 483072 557912 483074 557932
rect 485778 557912 485834 557968
rect 483018 557776 483074 557832
rect 487158 557796 487214 557832
rect 487158 557776 487160 557796
rect 487160 557776 487212 557796
rect 487212 557776 487214 557796
rect 488538 557640 488594 557696
rect 474830 413888 474886 413944
rect 477590 413888 477646 413944
rect 476118 413752 476174 413808
rect 477498 413788 477500 413808
rect 477500 413788 477552 413808
rect 477552 413788 477554 413808
rect 477498 413752 477554 413788
rect 478878 413652 478880 413672
rect 478880 413652 478932 413672
rect 478932 413652 478934 413672
rect 478878 413616 478934 413652
rect 480442 413480 480498 413536
rect 485778 413516 485780 413536
rect 485780 413516 485832 413536
rect 485832 413516 485834 413536
rect 485778 413480 485834 413516
rect 481638 413380 481640 413400
rect 481640 413380 481692 413400
rect 481692 413380 481694 413400
rect 481638 413344 481694 413380
rect 483018 413344 483074 413400
rect 484398 413208 484454 413264
rect 488538 413244 488540 413264
rect 488540 413244 488592 413264
rect 488592 413244 488594 413264
rect 488538 413208 488594 413244
rect 487158 413072 487214 413128
rect 489918 412936 489974 412992
rect 491298 412972 491300 412992
rect 491300 412972 491352 412992
rect 491352 412972 491354 412992
rect 491298 412936 491354 412972
rect 491390 412664 491446 412720
rect 492678 412664 492734 412720
rect 494058 412684 494114 412720
rect 494058 412664 494060 412684
rect 494060 412664 494112 412684
rect 494112 412664 494114 412684
rect 505098 413752 505154 413808
rect 506478 413652 506480 413672
rect 506480 413652 506532 413672
rect 506532 413652 506534 413672
rect 506478 413616 506534 413652
rect 495714 412700 495716 412720
rect 495716 412700 495768 412720
rect 495768 412700 495770 412720
rect 495714 412664 495770 412700
rect 496818 412664 496874 412720
rect 498290 412664 498346 412720
rect 499578 412664 499634 412720
rect 501050 412664 501106 412720
rect 502522 412664 502578 412720
rect 503718 412664 503774 412720
rect 503994 412664 504050 412720
rect 517518 412664 517574 412720
rect 473450 410352 473506 410408
rect 526442 409944 526498 410000
rect 343638 318724 343640 318744
rect 343640 318724 343692 318744
rect 343692 318724 343694 318744
rect 343638 318688 343694 318724
rect 453118 318724 453120 318744
rect 453120 318724 453172 318744
rect 453172 318724 453174 318744
rect 453118 318688 453174 318724
rect 278778 4800 278834 4856
rect 259458 3304 259514 3360
<< metal3 >>
rect 583520 697900 584960 698140
rect -960 696540 480 696780
rect 583520 686204 584960 686444
rect -960 682124 480 682364
rect 583520 674508 584960 674748
rect -960 667844 480 668084
rect 583520 662676 584960 662916
rect -960 653428 480 653668
rect 378133 652900 378199 652901
rect 383561 652900 383627 652901
rect 378133 652896 378180 652900
rect 378244 652898 378250 652900
rect 383510 652898 383516 652900
rect 378133 652840 378138 652896
rect 378133 652836 378180 652840
rect 378244 652838 378290 652898
rect 383470 652838 383516 652898
rect 383580 652896 383627 652900
rect 383622 652840 383627 652896
rect 378244 652836 378250 652838
rect 383510 652836 383516 652838
rect 383580 652836 383627 652840
rect 378133 652835 378199 652836
rect 383561 652835 383627 652836
rect 508405 652900 508471 652901
rect 513373 652900 513439 652901
rect 508405 652896 508452 652900
rect 508516 652898 508522 652900
rect 508405 652840 508410 652896
rect 508405 652836 508452 652840
rect 508516 652838 508562 652898
rect 513373 652896 513420 652900
rect 513484 652898 513490 652900
rect 513373 652840 513378 652896
rect 508516 652836 508522 652838
rect 513373 652836 513420 652840
rect 513484 652838 513530 652898
rect 513484 652836 513490 652838
rect 508405 652835 508471 652836
rect 513373 652835 513439 652836
rect 258533 651676 258599 651677
rect 263593 651676 263659 651677
rect 258533 651672 258576 651676
rect 258640 651674 258646 651676
rect 263565 651674 263571 651676
rect 258533 651616 258538 651672
rect 258533 651612 258576 651616
rect 258640 651614 258690 651674
rect 263502 651614 263571 651674
rect 263635 651672 263659 651676
rect 263654 651616 263659 651672
rect 258640 651612 258646 651614
rect 263565 651612 263571 651614
rect 263635 651612 263659 651616
rect 258533 651611 258599 651612
rect 263593 651611 263659 651612
rect 129222 651068 129228 651132
rect 129292 651130 129298 651132
rect 133822 651130 133828 651132
rect 129292 651070 133828 651130
rect 129292 651068 129298 651070
rect 133822 651068 133828 651070
rect 133892 651130 133898 651132
rect 135069 651130 135135 651133
rect 133892 651128 135135 651130
rect 133892 651072 135074 651128
rect 135130 651072 135135 651128
rect 133892 651070 135135 651072
rect 133892 651068 133898 651070
rect 135069 651067 135135 651070
rect 583520 650980 584960 651220
rect 266629 649906 266695 649909
rect 387149 649906 387215 649909
rect 389173 649906 389239 649909
rect 266629 649904 266738 649906
rect 266629 649848 266634 649904
rect 266690 649848 266738 649904
rect 266629 649843 266738 649848
rect 387068 649904 389239 649906
rect 387068 649848 387154 649904
rect 387210 649848 389178 649904
rect 389234 649848 389239 649904
rect 387068 649846 389239 649848
rect 387149 649843 387258 649846
rect 389173 649843 389239 649846
rect 516409 649906 516475 649909
rect 516409 649904 516610 649906
rect 516409 649848 516414 649904
rect 516470 649848 516610 649904
rect 516409 649846 516610 649848
rect 516409 649843 516475 649846
rect 137645 649713 137711 649716
rect 137172 649711 137711 649713
rect 137172 649655 137650 649711
rect 137706 649655 137711 649711
rect 266678 649683 266738 649843
rect 387198 649683 387258 649843
rect 516550 649683 516610 649846
rect 137172 649653 137711 649655
rect 137645 649650 137711 649653
rect 57881 646098 57947 646101
rect 60046 646098 60106 646587
rect 57881 646096 60106 646098
rect 57881 646040 57886 646096
rect 57942 646040 60106 646096
rect 57881 646038 60106 646040
rect 188337 646098 188403 646101
rect 190134 646098 190194 646587
rect 188337 646096 190194 646098
rect 188337 646040 188342 646096
rect 188398 646040 190194 646096
rect 188337 646038 190194 646040
rect 307385 646098 307451 646101
rect 310102 646098 310162 646587
rect 307385 646096 310162 646098
rect 307385 646040 307390 646096
rect 307446 646040 310162 646096
rect 307385 646038 310162 646040
rect 438117 646098 438183 646101
rect 440006 646098 440066 646587
rect 438117 646096 440066 646098
rect 438117 646040 438122 646096
rect 438178 646040 440066 646096
rect 438117 646038 440066 646040
rect 57881 646035 57947 646038
rect 188337 646035 188403 646038
rect 307385 646035 307451 646038
rect 438117 646035 438183 646038
rect 57789 645010 57855 645013
rect 60046 645010 60106 645459
rect 57789 645008 60106 645010
rect 57789 644952 57794 645008
rect 57850 644952 60106 645008
rect 57789 644950 60106 644952
rect 188429 645010 188495 645013
rect 190134 645010 190194 645459
rect 188429 645008 190194 645010
rect 188429 644952 188434 645008
rect 188490 644952 190194 645008
rect 188429 644950 190194 644952
rect 307109 645010 307175 645013
rect 310102 645010 310162 645459
rect 307109 645008 310162 645010
rect 307109 644952 307114 645008
rect 307170 644952 310162 645008
rect 307109 644950 310162 644952
rect 438209 645010 438275 645013
rect 440006 645010 440066 645459
rect 438209 645008 440066 645010
rect 438209 644952 438214 645008
rect 438270 644952 440066 645008
rect 438209 644950 440066 644952
rect 57789 644947 57855 644950
rect 188429 644947 188495 644950
rect 307109 644947 307175 644950
rect 438209 644947 438275 644950
rect 57697 643242 57763 643245
rect 60046 643242 60106 643759
rect 57697 643240 60106 643242
rect 57697 643184 57702 643240
rect 57758 643184 60106 643240
rect 57697 643182 60106 643184
rect 188521 643242 188587 643245
rect 190134 643242 190194 643759
rect 307109 643514 307175 643517
rect 310102 643514 310162 643759
rect 307109 643512 310162 643514
rect 307109 643456 307114 643512
rect 307170 643456 310162 643512
rect 307109 643454 310162 643456
rect 307109 643451 307175 643454
rect 188521 643240 190194 643242
rect 188521 643184 188526 643240
rect 188582 643184 190194 643240
rect 188521 643182 190194 643184
rect 438301 643242 438367 643245
rect 440006 643242 440066 643759
rect 438301 643240 440066 643242
rect 438301 643184 438306 643240
rect 438362 643184 440066 643240
rect 438301 643182 440066 643184
rect 57697 643179 57763 643182
rect 188521 643179 188587 643182
rect 438301 643179 438367 643182
rect 57605 642018 57671 642021
rect 60046 642018 60106 642631
rect 57605 642016 60106 642018
rect 57605 641960 57610 642016
rect 57666 641960 60106 642016
rect 57605 641958 60106 641960
rect 188613 642018 188679 642021
rect 190134 642018 190194 642631
rect 307661 642154 307727 642157
rect 310102 642154 310162 642631
rect 307661 642152 310162 642154
rect 307661 642096 307666 642152
rect 307722 642096 310162 642152
rect 307661 642094 310162 642096
rect 307661 642091 307727 642094
rect 188613 642016 190194 642018
rect 188613 641960 188618 642016
rect 188674 641960 190194 642016
rect 188613 641958 190194 641960
rect 438393 642018 438459 642021
rect 440006 642018 440066 642631
rect 438393 642016 440066 642018
rect 438393 641960 438398 642016
rect 438454 641960 440066 642016
rect 438393 641958 440066 641960
rect 57605 641955 57671 641958
rect 188613 641955 188679 641958
rect 438393 641955 438459 641958
rect 57513 640386 57579 640389
rect 60046 640386 60106 640931
rect 57513 640384 60106 640386
rect 57513 640328 57518 640384
rect 57574 640328 60106 640384
rect 57513 640326 60106 640328
rect 188705 640386 188771 640389
rect 190134 640386 190194 640931
rect 307661 640522 307727 640525
rect 310102 640522 310162 640931
rect 307661 640520 310162 640522
rect 307661 640464 307666 640520
rect 307722 640464 310162 640520
rect 307661 640462 310162 640464
rect 307661 640459 307727 640462
rect 188705 640384 190194 640386
rect 188705 640328 188710 640384
rect 188766 640328 190194 640384
rect 188705 640326 190194 640328
rect 438485 640386 438551 640389
rect 440006 640386 440066 640931
rect 438485 640384 440066 640386
rect 438485 640328 438490 640384
rect 438546 640328 440066 640384
rect 438485 640326 440066 640328
rect 57513 640323 57579 640326
rect 188705 640323 188771 640326
rect 438485 640323 438551 640326
rect 57421 639298 57487 639301
rect 60046 639298 60106 639803
rect 57421 639296 60106 639298
rect -960 639012 480 639252
rect 57421 639240 57426 639296
rect 57482 639240 60106 639296
rect 57421 639238 60106 639240
rect 188797 639298 188863 639301
rect 190134 639298 190194 639803
rect 188797 639296 190194 639298
rect 188797 639240 188802 639296
rect 188858 639240 190194 639296
rect 188797 639238 190194 639240
rect 307017 639298 307083 639301
rect 310102 639298 310162 639803
rect 307017 639296 310162 639298
rect 307017 639240 307022 639296
rect 307078 639240 310162 639296
rect 307017 639238 310162 639240
rect 438577 639298 438643 639301
rect 440006 639298 440066 639803
rect 438577 639296 440066 639298
rect 438577 639240 438582 639296
rect 438638 639240 440066 639296
rect 583520 639284 584960 639524
rect 438577 639238 440066 639240
rect 57421 639235 57487 639238
rect 188797 639235 188863 639238
rect 307017 639235 307083 639238
rect 438577 639235 438643 639238
rect 57329 637666 57395 637669
rect 60046 637666 60106 638103
rect 57329 637664 60106 637666
rect 57329 637608 57334 637664
rect 57390 637608 60106 637664
rect 57329 637606 60106 637608
rect 188889 637666 188955 637669
rect 190134 637666 190194 638103
rect 306833 637938 306899 637941
rect 310102 637938 310162 638103
rect 306833 637936 310162 637938
rect 306833 637880 306838 637936
rect 306894 637880 310162 637936
rect 306833 637878 310162 637880
rect 306833 637875 306899 637878
rect 188889 637664 190194 637666
rect 188889 637608 188894 637664
rect 188950 637608 190194 637664
rect 188889 637606 190194 637608
rect 438669 637666 438735 637669
rect 440006 637666 440066 638103
rect 438669 637664 440066 637666
rect 438669 637608 438674 637664
rect 438730 637608 440066 637664
rect 438669 637606 440066 637608
rect 57329 637603 57395 637606
rect 188889 637603 188955 637606
rect 438669 637603 438735 637606
rect 583520 627588 584960 627828
rect -960 624732 480 624972
rect 583520 615756 584960 615996
rect -960 610316 480 610556
rect 583520 604060 584960 604300
rect -960 595900 480 596140
rect 583520 592364 584960 592604
rect 139393 589658 139459 589661
rect 136958 589656 139459 589658
rect 136958 589600 139398 589656
rect 139454 589600 139459 589656
rect 136958 589598 139459 589600
rect 136958 586614 137018 589598
rect 139393 589595 139459 589598
rect 267230 589386 267290 589412
rect 269113 589386 269179 589389
rect 267230 589384 269179 589386
rect 267230 589328 269118 589384
rect 269174 589328 269179 589384
rect 267230 589326 269179 589328
rect 269113 589323 269179 589326
rect 267230 587210 267290 587712
rect 269113 587210 269179 587213
rect 270350 587210 270356 587212
rect 267230 587208 270356 587210
rect 267230 587152 269118 587208
rect 269174 587152 270356 587208
rect 267230 587150 270356 587152
rect 136958 586584 137172 586614
rect 136988 586554 137202 586584
rect -960 581620 480 581860
rect 137142 580928 137202 586554
rect 267230 580410 267290 587150
rect 269113 587147 269179 587150
rect 270350 587148 270356 587150
rect 270420 587148 270426 587212
rect 387198 587210 387258 589412
rect 517102 589386 517162 589412
rect 518893 589386 518959 589389
rect 517102 589384 518959 589386
rect 517102 589328 518898 589384
rect 518954 589328 518959 589384
rect 517102 589326 518959 589328
rect 518893 589323 518959 589326
rect 518893 587754 518959 587757
rect 517102 587752 518959 587754
rect 517102 587696 518898 587752
rect 518954 587696 518959 587752
rect 517102 587694 518959 587696
rect 387558 587210 387564 587212
rect 387198 587150 387564 587210
rect 387198 580954 387258 587150
rect 387558 587148 387564 587150
rect 387628 587148 387634 587212
rect 389214 580954 389220 580956
rect 387198 580894 389220 580954
rect 389214 580892 389220 580894
rect 389284 580892 389290 580956
rect 517102 580954 517162 587694
rect 518893 587691 518959 587694
rect 518934 580954 518940 580956
rect 517102 580894 518940 580954
rect 518934 580892 518940 580894
rect 519004 580892 519010 580956
rect 583520 580668 584960 580908
rect 270401 580410 270467 580413
rect 267230 580408 270467 580410
rect 267230 580352 270406 580408
rect 270462 580352 270467 580408
rect 267230 580350 270467 580352
rect 270401 580347 270467 580350
rect 57237 579730 57303 579733
rect 60046 579730 60106 580255
rect 57237 579728 60106 579730
rect 57237 579672 57242 579728
rect 57298 579672 60106 579728
rect 57237 579670 60106 579672
rect 188981 579730 189047 579733
rect 190134 579730 190194 580255
rect 307661 579866 307727 579869
rect 310102 579866 310162 580255
rect 307661 579864 310162 579866
rect 307661 579808 307666 579864
rect 307722 579808 310162 579864
rect 307661 579806 310162 579808
rect 307661 579803 307727 579806
rect 188981 579728 190194 579730
rect 188981 579672 188986 579728
rect 189042 579672 190194 579728
rect 188981 579670 190194 579672
rect 438761 579730 438827 579733
rect 440006 579730 440066 580255
rect 438761 579728 440066 579730
rect 438761 579672 438766 579728
rect 438822 579672 440066 579728
rect 438761 579670 440066 579672
rect 57237 579667 57303 579670
rect 188981 579667 189047 579670
rect 438761 579667 438827 579670
rect 60590 578988 60596 579052
rect 60660 578988 60666 579052
rect 188838 578988 188844 579052
rect 188908 579050 188914 579052
rect 281533 579050 281599 579053
rect 282494 579050 282500 579052
rect 188908 578990 190194 579050
rect 188908 578988 188914 578990
rect 60598 578555 60658 578988
rect 190134 578555 190194 578990
rect 281533 579048 282500 579050
rect 281533 578992 281538 579048
rect 281594 578992 282500 579048
rect 281533 578990 282500 578992
rect 281533 578987 281599 578990
rect 282494 578988 282500 578990
rect 282564 578988 282570 579052
rect 310278 578988 310284 579052
rect 310348 578988 310354 579052
rect 437422 578988 437428 579052
rect 437492 579050 437498 579052
rect 437492 578990 440066 579050
rect 437492 578988 437498 578990
rect 310286 578555 310346 578988
rect 440006 578555 440066 578990
rect 583520 568836 584960 569076
rect -960 567204 480 567444
rect 210969 560010 211035 560013
rect 211102 560010 211108 560012
rect 210969 560008 211108 560010
rect 210969 559952 210974 560008
rect 211030 559952 211108 560008
rect 210969 559950 211108 559952
rect 210969 559947 211035 559950
rect 211102 559948 211108 559950
rect 211172 559948 211178 560012
rect 348417 559330 348483 559333
rect 351862 559330 351868 559332
rect 348417 559328 351868 559330
rect 348417 559272 348422 559328
rect 348478 559272 351868 559328
rect 348417 559270 351868 559272
rect 348417 559267 348483 559270
rect 351862 559268 351868 559270
rect 351932 559268 351938 559332
rect 358169 559330 358235 559333
rect 358854 559330 358860 559332
rect 358169 559328 358860 559330
rect 358169 559272 358174 559328
rect 358230 559272 358860 559328
rect 358169 559270 358860 559272
rect 358169 559267 358235 559270
rect 358854 559268 358860 559270
rect 358924 559268 358930 559332
rect 67398 558860 67404 558924
rect 67468 558922 67474 558924
rect 67541 558922 67607 558925
rect 67468 558920 67607 558922
rect 67468 558864 67546 558920
rect 67602 558864 67607 558920
rect 67468 558862 67607 558864
rect 67468 558860 67474 558862
rect 67541 558859 67607 558862
rect 68502 558860 68508 558924
rect 68572 558922 68578 558924
rect 68921 558922 68987 558925
rect 68572 558920 68987 558922
rect 68572 558864 68926 558920
rect 68982 558864 68987 558920
rect 68572 558862 68987 558864
rect 68572 558860 68578 558862
rect 68921 558859 68987 558862
rect 70158 558860 70164 558924
rect 70228 558922 70234 558924
rect 70301 558922 70367 558925
rect 71681 558924 71747 558925
rect 70228 558920 70367 558922
rect 70228 558864 70306 558920
rect 70362 558864 70367 558920
rect 70228 558862 70367 558864
rect 70228 558860 70234 558862
rect 70301 558859 70367 558862
rect 71630 558860 71636 558924
rect 71700 558922 71747 558924
rect 71700 558920 71792 558922
rect 71742 558864 71792 558920
rect 71700 558862 71792 558864
rect 71700 558860 71747 558862
rect 72366 558860 72372 558924
rect 72436 558922 72442 558924
rect 72509 558922 72575 558925
rect 72436 558920 72575 558922
rect 72436 558864 72514 558920
rect 72570 558864 72575 558920
rect 72436 558862 72575 558864
rect 72436 558860 72442 558862
rect 71681 558859 71747 558860
rect 72509 558859 72575 558862
rect 72918 558860 72924 558924
rect 72988 558922 72994 558924
rect 73061 558922 73127 558925
rect 73705 558924 73771 558925
rect 74257 558924 74323 558925
rect 74993 558924 75059 558925
rect 73654 558922 73660 558924
rect 72988 558920 73127 558922
rect 72988 558864 73066 558920
rect 73122 558864 73127 558920
rect 72988 558862 73127 558864
rect 73614 558862 73660 558922
rect 73724 558920 73771 558924
rect 74206 558922 74212 558924
rect 73766 558864 73771 558920
rect 72988 558860 72994 558862
rect 73061 558859 73127 558862
rect 73654 558860 73660 558862
rect 73724 558860 73771 558864
rect 74166 558862 74212 558922
rect 74276 558920 74323 558924
rect 74942 558922 74948 558924
rect 74318 558864 74323 558920
rect 74206 558860 74212 558862
rect 74276 558860 74323 558864
rect 74902 558862 74948 558922
rect 75012 558920 75059 558924
rect 75054 558864 75059 558920
rect 74942 558860 74948 558862
rect 75012 558860 75059 558864
rect 75678 558860 75684 558924
rect 75748 558922 75754 558924
rect 75821 558922 75887 558925
rect 76833 558924 76899 558925
rect 77385 558924 77451 558925
rect 76782 558922 76788 558924
rect 75748 558920 75887 558922
rect 75748 558864 75826 558920
rect 75882 558864 75887 558920
rect 75748 558862 75887 558864
rect 76742 558862 76788 558922
rect 76852 558920 76899 558924
rect 77334 558922 77340 558924
rect 76894 558864 76899 558920
rect 75748 558860 75754 558862
rect 73705 558859 73771 558860
rect 74257 558859 74323 558860
rect 74993 558859 75059 558860
rect 75821 558859 75887 558862
rect 76782 558860 76788 558862
rect 76852 558860 76899 558864
rect 77294 558862 77340 558922
rect 77404 558920 77451 558924
rect 77446 558864 77451 558920
rect 77334 558860 77340 558862
rect 77404 558860 77451 558864
rect 78070 558860 78076 558924
rect 78140 558922 78146 558924
rect 78581 558922 78647 558925
rect 78140 558920 78647 558922
rect 78140 558864 78586 558920
rect 78642 558864 78647 558920
rect 78140 558862 78647 558864
rect 78140 558860 78146 558862
rect 76833 558859 76899 558860
rect 77385 558859 77451 558860
rect 78581 558859 78647 558862
rect 79174 558860 79180 558924
rect 79244 558922 79250 558924
rect 79317 558922 79383 558925
rect 79869 558924 79935 558925
rect 79869 558922 79916 558924
rect 79244 558920 79383 558922
rect 79244 558864 79322 558920
rect 79378 558864 79383 558920
rect 79244 558862 79383 558864
rect 79824 558920 79916 558922
rect 79824 558864 79874 558920
rect 79824 558862 79916 558864
rect 79244 558860 79250 558862
rect 79317 558859 79383 558862
rect 79869 558860 79916 558862
rect 79980 558860 79986 558924
rect 80646 558860 80652 558924
rect 80716 558922 80722 558924
rect 80789 558922 80855 558925
rect 81249 558924 81315 558925
rect 81985 558924 82051 558925
rect 82905 558924 82971 558925
rect 83825 558924 83891 558925
rect 84193 558924 84259 558925
rect 81198 558922 81204 558924
rect 80716 558920 80855 558922
rect 80716 558864 80794 558920
rect 80850 558864 80855 558920
rect 80716 558862 80855 558864
rect 81158 558862 81204 558922
rect 81268 558920 81315 558924
rect 81934 558922 81940 558924
rect 81310 558864 81315 558920
rect 80716 558860 80722 558862
rect 79869 558859 79935 558860
rect 80789 558859 80855 558862
rect 81198 558860 81204 558862
rect 81268 558860 81315 558864
rect 81894 558862 81940 558922
rect 82004 558920 82051 558924
rect 82854 558922 82860 558924
rect 82046 558864 82051 558920
rect 81934 558860 81940 558862
rect 82004 558860 82051 558864
rect 82814 558862 82860 558922
rect 82924 558920 82971 558924
rect 83774 558922 83780 558924
rect 82966 558864 82971 558920
rect 82854 558860 82860 558862
rect 82924 558860 82971 558864
rect 83734 558862 83780 558922
rect 83844 558920 83891 558924
rect 83886 558864 83891 558920
rect 83774 558860 83780 558862
rect 83844 558860 83891 558864
rect 84142 558860 84148 558924
rect 84212 558922 84259 558924
rect 84212 558920 84304 558922
rect 84254 558864 84304 558920
rect 84212 558862 84304 558864
rect 84212 558860 84259 558862
rect 85062 558860 85068 558924
rect 85132 558922 85138 558924
rect 85481 558922 85547 558925
rect 85132 558920 85547 558922
rect 85132 558864 85486 558920
rect 85542 558864 85547 558920
rect 85132 558862 85547 558864
rect 85132 558860 85138 558862
rect 81249 558859 81315 558860
rect 81985 558859 82051 558860
rect 82905 558859 82971 558860
rect 83825 558859 83891 558860
rect 84193 558859 84259 558860
rect 85481 558859 85547 558862
rect 86309 558924 86375 558925
rect 86769 558924 86835 558925
rect 87873 558924 87939 558925
rect 88241 558924 88307 558925
rect 86309 558920 86356 558924
rect 86420 558922 86426 558924
rect 86309 558864 86314 558920
rect 86309 558860 86356 558864
rect 86420 558862 86466 558922
rect 86420 558860 86426 558862
rect 86718 558860 86724 558924
rect 86788 558922 86835 558924
rect 87822 558922 87828 558924
rect 86788 558920 86880 558922
rect 86830 558864 86880 558920
rect 86788 558862 86880 558864
rect 87782 558862 87828 558922
rect 87892 558920 87939 558924
rect 87934 558864 87939 558920
rect 86788 558860 86835 558862
rect 87822 558860 87828 558862
rect 87892 558860 87939 558864
rect 88190 558860 88196 558924
rect 88260 558922 88307 558924
rect 88885 558924 88951 558925
rect 89161 558924 89227 558925
rect 88885 558922 88932 558924
rect 88260 558920 88352 558922
rect 88302 558864 88352 558920
rect 88260 558862 88352 558864
rect 88840 558920 88932 558922
rect 88840 558864 88890 558920
rect 88840 558862 88932 558864
rect 88260 558860 88307 558862
rect 86309 558859 86375 558860
rect 86769 558859 86835 558860
rect 87873 558859 87939 558860
rect 88241 558859 88307 558860
rect 88885 558860 88932 558862
rect 88996 558860 89002 558924
rect 89110 558922 89116 558924
rect 89070 558862 89116 558922
rect 89180 558920 89227 558924
rect 89222 558864 89227 558920
rect 89110 558860 89116 558862
rect 89180 558860 89227 558864
rect 88885 558859 88951 558860
rect 89161 558859 89227 558860
rect 89805 558924 89871 558925
rect 91001 558924 91067 558925
rect 89805 558920 89852 558924
rect 89916 558922 89922 558924
rect 89805 558864 89810 558920
rect 89805 558860 89852 558864
rect 89916 558862 89962 558922
rect 89916 558860 89922 558862
rect 90950 558860 90956 558924
rect 91020 558922 91067 558924
rect 91020 558920 91112 558922
rect 91062 558864 91112 558920
rect 91020 558862 91112 558864
rect 91020 558860 91067 558862
rect 91870 558860 91876 558924
rect 91940 558922 91946 558924
rect 92197 558922 92263 558925
rect 92473 558924 92539 558925
rect 92422 558922 92428 558924
rect 91940 558920 92263 558922
rect 91940 558864 92202 558920
rect 92258 558864 92263 558920
rect 91940 558862 92263 558864
rect 92382 558862 92428 558922
rect 92492 558920 92539 558924
rect 92534 558864 92539 558920
rect 91940 558860 91946 558862
rect 89805 558859 89871 558860
rect 91001 558859 91067 558860
rect 92197 558859 92263 558862
rect 92422 558860 92428 558862
rect 92492 558860 92539 558864
rect 92473 558859 92539 558860
rect 93301 558924 93367 558925
rect 93761 558924 93827 558925
rect 95049 558924 95115 558925
rect 93301 558920 93348 558924
rect 93412 558922 93418 558924
rect 93710 558922 93716 558924
rect 93301 558864 93306 558920
rect 93301 558860 93348 558864
rect 93412 558862 93458 558922
rect 93670 558862 93716 558922
rect 93780 558920 93827 558924
rect 93822 558864 93827 558920
rect 93412 558860 93418 558862
rect 93710 558860 93716 558862
rect 93780 558860 93827 558864
rect 94998 558860 95004 558924
rect 95068 558922 95115 558924
rect 95693 558924 95759 558925
rect 96521 558924 96587 558925
rect 95068 558920 95160 558922
rect 95110 558864 95160 558920
rect 95068 558862 95160 558864
rect 95693 558920 95740 558924
rect 95804 558922 95810 558924
rect 95693 558864 95698 558920
rect 95068 558860 95115 558862
rect 93301 558859 93367 558860
rect 93761 558859 93827 558860
rect 95049 558859 95115 558860
rect 95693 558860 95740 558864
rect 95804 558862 95850 558922
rect 95804 558860 95810 558862
rect 96470 558860 96476 558924
rect 96540 558922 96587 558924
rect 96540 558920 96632 558922
rect 96582 558864 96632 558920
rect 96540 558862 96632 558864
rect 96540 558860 96587 558862
rect 97022 558860 97028 558924
rect 97092 558922 97098 558924
rect 97165 558922 97231 558925
rect 97809 558924 97875 558925
rect 98361 558924 98427 558925
rect 97758 558922 97764 558924
rect 97092 558920 97231 558922
rect 97092 558864 97170 558920
rect 97226 558864 97231 558920
rect 97092 558862 97231 558864
rect 97718 558862 97764 558922
rect 97828 558920 97875 558924
rect 98310 558922 98316 558924
rect 97870 558864 97875 558920
rect 97092 558860 97098 558862
rect 95693 558859 95759 558860
rect 96521 558859 96587 558860
rect 97165 558859 97231 558862
rect 97758 558860 97764 558862
rect 97828 558860 97875 558864
rect 98270 558862 98316 558922
rect 98380 558920 98427 558924
rect 98422 558864 98427 558920
rect 98310 558860 98316 558862
rect 98380 558860 98427 558864
rect 99046 558860 99052 558924
rect 99116 558922 99122 558924
rect 99281 558922 99347 558925
rect 100017 558924 100083 558925
rect 102041 558924 102107 558925
rect 104801 558924 104867 558925
rect 99966 558922 99972 558924
rect 99116 558920 99347 558922
rect 99116 558864 99286 558920
rect 99342 558864 99347 558920
rect 99116 558862 99347 558864
rect 99926 558862 99972 558922
rect 100036 558920 100083 558924
rect 101990 558922 101996 558924
rect 100078 558864 100083 558920
rect 99116 558860 99122 558862
rect 97809 558859 97875 558860
rect 98361 558859 98427 558860
rect 99281 558859 99347 558862
rect 99966 558860 99972 558862
rect 100036 558860 100083 558864
rect 101950 558862 101996 558922
rect 102060 558920 102107 558924
rect 104750 558922 104756 558924
rect 102102 558864 102107 558920
rect 101990 558860 101996 558862
rect 102060 558860 102107 558864
rect 104710 558862 104756 558922
rect 104820 558920 104867 558924
rect 104862 558864 104867 558920
rect 104750 558860 104756 558862
rect 104820 558860 104867 558864
rect 107142 558860 107148 558924
rect 107212 558922 107218 558924
rect 107285 558922 107351 558925
rect 108481 558924 108547 558925
rect 108430 558922 108436 558924
rect 107212 558920 107351 558922
rect 107212 558864 107290 558920
rect 107346 558864 107351 558920
rect 107212 558862 107351 558864
rect 108390 558862 108436 558922
rect 108500 558920 108547 558924
rect 108542 558864 108547 558920
rect 107212 558860 107218 558862
rect 100017 558859 100083 558860
rect 102041 558859 102107 558860
rect 104801 558859 104867 558860
rect 107285 558859 107351 558862
rect 108430 558860 108436 558862
rect 108500 558860 108547 558864
rect 108481 558859 108547 558860
rect 195973 558922 196039 558925
rect 200205 558924 200271 558925
rect 196198 558922 196204 558924
rect 195973 558920 196204 558922
rect 195973 558864 195978 558920
rect 196034 558864 196204 558920
rect 195973 558862 196204 558864
rect 195973 558859 196039 558862
rect 196198 558860 196204 558862
rect 196268 558860 196274 558924
rect 200205 558922 200252 558924
rect 200160 558920 200252 558922
rect 200160 558864 200210 558920
rect 200160 558862 200252 558864
rect 200205 558860 200252 558862
rect 200316 558860 200322 558924
rect 202638 558860 202644 558924
rect 202708 558922 202714 558924
rect 202781 558922 202847 558925
rect 203793 558924 203859 558925
rect 203742 558922 203748 558924
rect 202708 558920 202847 558922
rect 202708 558864 202786 558920
rect 202842 558864 202847 558920
rect 202708 558862 202847 558864
rect 203702 558862 203748 558922
rect 203812 558920 203859 558924
rect 203854 558864 203859 558920
rect 202708 558860 202714 558862
rect 200205 558859 200271 558860
rect 202781 558859 202847 558862
rect 203742 558860 203748 558862
rect 203812 558860 203859 558864
rect 203926 558860 203932 558924
rect 203996 558922 204002 558924
rect 204161 558922 204227 558925
rect 203996 558920 204227 558922
rect 203996 558864 204166 558920
rect 204222 558864 204227 558920
rect 203996 558862 204227 558864
rect 203996 558860 204002 558862
rect 203793 558859 203859 558860
rect 204161 558859 204227 558862
rect 205398 558860 205404 558924
rect 205468 558922 205474 558924
rect 205541 558922 205607 558925
rect 205468 558920 205607 558922
rect 205468 558864 205546 558920
rect 205602 558864 205607 558920
rect 205468 558862 205607 558864
rect 205468 558860 205474 558862
rect 205541 558859 205607 558862
rect 206134 558860 206140 558924
rect 206204 558922 206210 558924
rect 206921 558922 206987 558925
rect 206204 558920 206987 558922
rect 206204 558864 206926 558920
rect 206982 558864 206987 558920
rect 206204 558862 206987 558864
rect 206204 558860 206210 558862
rect 206921 558859 206987 558862
rect 208342 558860 208348 558924
rect 208412 558922 208418 558924
rect 208485 558922 208551 558925
rect 210601 558924 210667 558925
rect 210550 558922 210556 558924
rect 208412 558920 208551 558922
rect 208412 558864 208490 558920
rect 208546 558864 208551 558920
rect 208412 558862 208551 558864
rect 210510 558862 210556 558922
rect 210620 558920 210667 558924
rect 210662 558864 210667 558920
rect 208412 558860 208418 558862
rect 208485 558859 208551 558862
rect 210550 558860 210556 558862
rect 210620 558860 210667 558864
rect 210601 558859 210667 558860
rect 211797 558924 211863 558925
rect 213177 558924 213243 558925
rect 211797 558920 211844 558924
rect 211908 558922 211914 558924
rect 213126 558922 213132 558924
rect 211797 558864 211802 558920
rect 211797 558860 211844 558864
rect 211908 558862 211954 558922
rect 213086 558862 213132 558922
rect 213196 558920 213243 558924
rect 213238 558864 213243 558920
rect 211908 558860 211914 558862
rect 213126 558860 213132 558862
rect 213196 558860 213243 558864
rect 211797 558859 211863 558860
rect 213177 558859 213243 558860
rect 214005 558924 214071 558925
rect 215293 558924 215359 558925
rect 214005 558920 214052 558924
rect 214116 558922 214122 558924
rect 214005 558864 214010 558920
rect 214005 558860 214052 558864
rect 214116 558862 214162 558922
rect 215293 558920 215340 558924
rect 215404 558922 215410 558924
rect 215293 558864 215298 558920
rect 214116 558860 214122 558862
rect 215293 558860 215340 558864
rect 215404 558862 215450 558922
rect 215404 558860 215410 558862
rect 216622 558860 216628 558924
rect 216692 558922 216698 558924
rect 217501 558922 217567 558925
rect 216692 558920 217567 558922
rect 216692 558864 217506 558920
rect 217562 558864 217567 558920
rect 216692 558862 217567 558864
rect 216692 558860 216698 558862
rect 214005 558859 214071 558860
rect 215293 558859 215359 558860
rect 217501 558859 217567 558862
rect 218789 558924 218855 558925
rect 220077 558924 220143 558925
rect 221089 558924 221155 558925
rect 218789 558920 218836 558924
rect 218900 558922 218906 558924
rect 218789 558864 218794 558920
rect 218789 558860 218836 558864
rect 218900 558862 218946 558922
rect 220077 558920 220124 558924
rect 220188 558922 220194 558924
rect 221038 558922 221044 558924
rect 220077 558864 220082 558920
rect 218900 558860 218906 558862
rect 220077 558860 220124 558864
rect 220188 558862 220234 558922
rect 220998 558862 221044 558922
rect 221108 558920 221155 558924
rect 221150 558864 221155 558920
rect 220188 558860 220194 558862
rect 221038 558860 221044 558862
rect 221108 558860 221155 558864
rect 218789 558859 218855 558860
rect 220077 558859 220143 558860
rect 221089 558859 221155 558860
rect 222193 558922 222259 558925
rect 224493 558924 224559 558925
rect 225873 558924 225939 558925
rect 222326 558922 222332 558924
rect 222193 558920 222332 558922
rect 222193 558864 222198 558920
rect 222254 558864 222332 558920
rect 222193 558862 222332 558864
rect 222193 558859 222259 558862
rect 222326 558860 222332 558862
rect 222396 558860 222402 558924
rect 224493 558920 224540 558924
rect 224604 558922 224610 558924
rect 225822 558922 225828 558924
rect 224493 558864 224498 558920
rect 224493 558860 224540 558864
rect 224604 558862 224650 558922
rect 225782 558862 225828 558922
rect 225892 558920 225939 558924
rect 226149 558924 226215 558925
rect 227161 558924 227227 558925
rect 226149 558922 226196 558924
rect 225934 558864 225939 558920
rect 224604 558860 224610 558862
rect 225822 558860 225828 558862
rect 225892 558860 225939 558864
rect 226104 558920 226196 558922
rect 226104 558864 226154 558920
rect 226104 558862 226196 558864
rect 224493 558859 224559 558860
rect 225873 558859 225939 558860
rect 226149 558860 226196 558862
rect 226260 558860 226266 558924
rect 227110 558922 227116 558924
rect 227070 558862 227116 558922
rect 227180 558920 227227 558924
rect 227222 558864 227227 558920
rect 227110 558860 227116 558862
rect 227180 558860 227227 558864
rect 227478 558860 227484 558924
rect 227548 558922 227554 558924
rect 227621 558922 227687 558925
rect 227548 558920 227687 558922
rect 227548 558864 227626 558920
rect 227682 558864 227687 558920
rect 227548 558862 227687 558864
rect 227548 558860 227554 558862
rect 226149 558859 226215 558860
rect 227161 558859 227227 558860
rect 227621 558859 227687 558862
rect 227989 558924 228055 558925
rect 227989 558920 228036 558924
rect 228100 558922 228106 558924
rect 227989 558864 227994 558920
rect 227989 558860 228036 558864
rect 228100 558862 228146 558922
rect 228100 558860 228106 558862
rect 228766 558860 228772 558924
rect 228836 558922 228842 558924
rect 229001 558922 229067 558925
rect 228836 558920 229067 558922
rect 228836 558864 229006 558920
rect 229062 558864 229067 558920
rect 228836 558862 229067 558864
rect 228836 558860 228842 558862
rect 227989 558859 228055 558860
rect 229001 558859 229067 558862
rect 229461 558924 229527 558925
rect 229461 558920 229508 558924
rect 229572 558922 229578 558924
rect 229461 558864 229466 558920
rect 229461 558860 229508 558864
rect 229572 558862 229618 558922
rect 229572 558860 229578 558862
rect 230238 558860 230244 558924
rect 230308 558922 230314 558924
rect 230381 558922 230447 558925
rect 230308 558920 230447 558922
rect 230308 558864 230386 558920
rect 230442 558864 230447 558920
rect 230308 558862 230447 558864
rect 230308 558860 230314 558862
rect 229461 558859 229527 558860
rect 230381 558859 230447 558862
rect 230790 558860 230796 558924
rect 230860 558922 230866 558924
rect 231761 558922 231827 558925
rect 233049 558924 233115 558925
rect 230860 558920 231827 558922
rect 230860 558864 231766 558920
rect 231822 558864 231827 558920
rect 230860 558862 231827 558864
rect 230860 558860 230866 558862
rect 231761 558859 231827 558862
rect 232998 558860 233004 558924
rect 233068 558922 233115 558924
rect 233233 558922 233299 558925
rect 234521 558924 234587 558925
rect 233550 558922 233556 558924
rect 233068 558920 233160 558922
rect 233110 558864 233160 558920
rect 233068 558862 233160 558864
rect 233233 558920 233556 558922
rect 233233 558864 233238 558920
rect 233294 558864 233556 558920
rect 233233 558862 233556 558864
rect 233068 558860 233115 558862
rect 233049 558859 233115 558860
rect 233233 558859 233299 558862
rect 233550 558860 233556 558862
rect 233620 558860 233626 558924
rect 234470 558860 234476 558924
rect 234540 558922 234587 558924
rect 234540 558920 234632 558922
rect 234582 558864 234632 558920
rect 234540 558862 234632 558864
rect 234540 558860 234587 558862
rect 235758 558860 235764 558924
rect 235828 558922 235834 558924
rect 235901 558922 235967 558925
rect 237281 558924 237347 558925
rect 235828 558920 235967 558922
rect 235828 558864 235906 558920
rect 235962 558864 235967 558920
rect 235828 558862 235967 558864
rect 235828 558860 235834 558862
rect 234521 558859 234587 558860
rect 235901 558859 235967 558862
rect 237230 558860 237236 558924
rect 237300 558922 237347 558924
rect 237300 558920 237392 558922
rect 237342 558864 237392 558920
rect 237300 558862 237392 558864
rect 237300 558860 237347 558862
rect 239622 558860 239628 558924
rect 239692 558922 239698 558924
rect 240041 558922 240107 558925
rect 313825 558924 313891 558925
rect 313774 558922 313780 558924
rect 239692 558920 240107 558922
rect 239692 558864 240046 558920
rect 240102 558864 240107 558920
rect 239692 558862 240107 558864
rect 313734 558862 313780 558922
rect 313844 558920 313891 558924
rect 317413 558924 317479 558925
rect 317413 558922 317460 558924
rect 313886 558864 313891 558920
rect 239692 558860 239698 558862
rect 237281 558859 237347 558860
rect 240041 558859 240107 558862
rect 313774 558860 313780 558862
rect 313844 558860 313891 558864
rect 317368 558920 317460 558922
rect 317368 558864 317418 558920
rect 317368 558862 317460 558864
rect 313825 558859 313891 558860
rect 317413 558860 317460 558862
rect 317524 558860 317530 558924
rect 318793 558922 318859 558925
rect 320173 558924 320239 558925
rect 318926 558922 318932 558924
rect 318793 558920 318932 558922
rect 318793 558864 318798 558920
rect 318854 558864 318932 558920
rect 318793 558862 318932 558864
rect 317413 558859 317479 558860
rect 318793 558859 318859 558862
rect 318926 558860 318932 558862
rect 318996 558860 319002 558924
rect 320173 558922 320220 558924
rect 320128 558920 320220 558922
rect 320128 558864 320178 558920
rect 320128 558862 320220 558864
rect 320173 558860 320220 558862
rect 320284 558860 320290 558924
rect 325693 558922 325759 558925
rect 326286 558922 326292 558924
rect 325693 558920 326292 558922
rect 325693 558864 325698 558920
rect 325754 558864 326292 558920
rect 325693 558862 326292 558864
rect 320173 558859 320239 558860
rect 325693 558859 325759 558862
rect 326286 558860 326292 558862
rect 326356 558860 326362 558924
rect 327073 558922 327139 558925
rect 327574 558922 327580 558924
rect 327073 558920 327580 558922
rect 327073 558864 327078 558920
rect 327134 558864 327580 558920
rect 327073 558862 327580 558864
rect 327073 558859 327139 558862
rect 327574 558860 327580 558862
rect 327644 558860 327650 558924
rect 329281 558922 329347 558925
rect 329598 558922 329604 558924
rect 329281 558920 329604 558922
rect 329281 558864 329286 558920
rect 329342 558864 329604 558920
rect 329281 558862 329604 558864
rect 329281 558859 329347 558862
rect 329598 558860 329604 558862
rect 329668 558860 329674 558924
rect 329925 558922 329991 558925
rect 331765 558924 331831 558925
rect 331070 558922 331076 558924
rect 329925 558920 331076 558922
rect 329925 558864 329930 558920
rect 329986 558864 331076 558920
rect 329925 558862 331076 558864
rect 329925 558859 329991 558862
rect 331070 558860 331076 558862
rect 331140 558860 331146 558924
rect 331765 558920 331812 558924
rect 331876 558922 331882 558924
rect 332593 558922 332659 558925
rect 333278 558922 333284 558924
rect 331765 558864 331770 558920
rect 331765 558860 331812 558864
rect 331876 558862 331922 558922
rect 332593 558920 333284 558922
rect 332593 558864 332598 558920
rect 332654 558864 333284 558920
rect 332593 558862 333284 558864
rect 331876 558860 331882 558862
rect 331765 558859 331831 558860
rect 332593 558859 332659 558862
rect 333278 558860 333284 558862
rect 333348 558860 333354 558924
rect 333973 558922 334039 558925
rect 334566 558922 334572 558924
rect 333973 558920 334572 558922
rect 333973 558864 333978 558920
rect 334034 558864 334572 558920
rect 333973 558862 334572 558864
rect 333973 558859 334039 558862
rect 334566 558860 334572 558862
rect 334636 558860 334642 558924
rect 335353 558922 335419 558925
rect 336733 558924 336799 558925
rect 335854 558922 335860 558924
rect 335353 558920 335860 558922
rect 335353 558864 335358 558920
rect 335414 558864 335860 558920
rect 335353 558862 335860 558864
rect 335353 558859 335419 558862
rect 335854 558860 335860 558862
rect 335924 558860 335930 558924
rect 336733 558922 336780 558924
rect 336688 558920 336780 558922
rect 336688 558864 336738 558920
rect 336688 558862 336780 558864
rect 336733 558860 336780 558862
rect 336844 558860 336850 558924
rect 337561 558922 337627 558925
rect 337694 558922 337700 558924
rect 337561 558920 337700 558922
rect 337561 558864 337566 558920
rect 337622 558864 337700 558920
rect 337561 558862 337700 558864
rect 336733 558859 336799 558860
rect 337561 558859 337627 558862
rect 337694 558860 337700 558862
rect 337764 558860 337770 558924
rect 338113 558922 338179 558925
rect 339166 558922 339172 558924
rect 338113 558920 339172 558922
rect 338113 558864 338118 558920
rect 338174 558864 339172 558920
rect 338113 558862 339172 558864
rect 338113 558859 338179 558862
rect 339166 558860 339172 558862
rect 339236 558860 339242 558924
rect 339493 558922 339559 558925
rect 340454 558922 340460 558924
rect 339493 558920 340460 558922
rect 339493 558864 339498 558920
rect 339554 558864 340460 558920
rect 339493 558862 340460 558864
rect 339493 558859 339559 558862
rect 340454 558860 340460 558862
rect 340524 558860 340530 558924
rect 340873 558922 340939 558925
rect 341742 558922 341748 558924
rect 340873 558920 341748 558922
rect 340873 558864 340878 558920
rect 340934 558864 341748 558920
rect 340873 558862 341748 558864
rect 340873 558859 340939 558862
rect 341742 558860 341748 558862
rect 341812 558860 341818 558924
rect 342253 558922 342319 558925
rect 342662 558922 342668 558924
rect 342253 558920 342668 558922
rect 342253 558864 342258 558920
rect 342314 558864 342668 558920
rect 342253 558862 342668 558864
rect 342253 558859 342319 558862
rect 342662 558860 342668 558862
rect 342732 558860 342738 558924
rect 343725 558922 343791 558925
rect 344277 558924 344343 558925
rect 343950 558922 343956 558924
rect 343725 558920 343956 558922
rect 343725 558864 343730 558920
rect 343786 558864 343956 558920
rect 343725 558862 343956 558864
rect 343725 558859 343791 558862
rect 343950 558860 343956 558862
rect 344020 558860 344026 558924
rect 344277 558920 344324 558924
rect 344388 558922 344394 558924
rect 345013 558922 345079 558925
rect 346158 558922 346164 558924
rect 344277 558864 344282 558920
rect 344277 558860 344324 558864
rect 344388 558862 344434 558922
rect 345013 558920 346164 558922
rect 345013 558864 345018 558920
rect 345074 558864 346164 558920
rect 345013 558862 346164 558864
rect 344388 558860 344394 558862
rect 344277 558859 344343 558860
rect 345013 558859 345079 558862
rect 346158 558860 346164 558862
rect 346228 558860 346234 558924
rect 346393 558922 346459 558925
rect 347446 558922 347452 558924
rect 346393 558920 347452 558922
rect 346393 558864 346398 558920
rect 346454 558864 347452 558920
rect 346393 558862 347452 558864
rect 346393 558859 346459 558862
rect 347446 558860 347452 558862
rect 347516 558860 347522 558924
rect 347773 558922 347839 558925
rect 348734 558922 348740 558924
rect 347773 558920 348740 558922
rect 347773 558864 347778 558920
rect 347834 558864 348740 558920
rect 347773 558862 348740 558864
rect 347773 558859 347839 558862
rect 348734 558860 348740 558862
rect 348804 558860 348810 558924
rect 349153 558922 349219 558925
rect 349654 558922 349660 558924
rect 349153 558920 349660 558922
rect 349153 558864 349158 558920
rect 349214 558864 349660 558920
rect 349153 558862 349660 558864
rect 349153 558859 349219 558862
rect 349654 558860 349660 558862
rect 349724 558860 349730 558924
rect 352005 558922 352071 558925
rect 356053 558924 356119 558925
rect 443085 558924 443151 558925
rect 352414 558922 352420 558924
rect 352005 558920 352420 558922
rect 352005 558864 352010 558920
rect 352066 558864 352420 558920
rect 352005 558862 352420 558864
rect 352005 558859 352071 558862
rect 352414 558860 352420 558862
rect 352484 558860 352490 558924
rect 356053 558922 356100 558924
rect 356008 558920 356100 558922
rect 356008 558864 356058 558920
rect 356008 558862 356100 558864
rect 356053 558860 356100 558862
rect 356164 558860 356170 558924
rect 443085 558920 443132 558924
rect 443196 558922 443202 558924
rect 445753 558922 445819 558925
rect 446254 558922 446260 558924
rect 443085 558864 443090 558920
rect 443085 558860 443132 558864
rect 443196 558862 443242 558922
rect 445753 558920 446260 558922
rect 445753 558864 445758 558920
rect 445814 558864 446260 558920
rect 445753 558862 446260 558864
rect 443196 558860 443202 558862
rect 356053 558859 356119 558860
rect 443085 558859 443151 558860
rect 445753 558859 445819 558862
rect 446254 558860 446260 558862
rect 446324 558860 446330 558924
rect 451273 558922 451339 558925
rect 451406 558922 451412 558924
rect 451273 558920 451412 558922
rect 451273 558864 451278 558920
rect 451334 558864 451412 558920
rect 451273 558862 451412 558864
rect 451273 558859 451339 558862
rect 451406 558860 451412 558862
rect 451476 558860 451482 558924
rect 452653 558922 452719 558925
rect 453665 558924 453731 558925
rect 452878 558922 452884 558924
rect 452653 558920 452884 558922
rect 452653 558864 452658 558920
rect 452714 558864 452884 558920
rect 452653 558862 452884 558864
rect 452653 558859 452719 558862
rect 452878 558860 452884 558862
rect 452948 558860 452954 558924
rect 453614 558922 453620 558924
rect 453574 558862 453620 558922
rect 453684 558920 453731 558924
rect 453726 558864 453731 558920
rect 453614 558860 453620 558862
rect 453684 558860 453731 558864
rect 453665 558859 453731 558860
rect 454033 558922 454099 558925
rect 455270 558922 455276 558924
rect 454033 558920 455276 558922
rect 454033 558864 454038 558920
rect 454094 558864 455276 558920
rect 454033 558862 455276 558864
rect 454033 558859 454099 558862
rect 455270 558860 455276 558862
rect 455340 558860 455346 558924
rect 455413 558922 455479 558925
rect 456558 558922 456564 558924
rect 455413 558920 456564 558922
rect 455413 558864 455418 558920
rect 455474 558864 456564 558920
rect 455413 558862 456564 558864
rect 455413 558859 455479 558862
rect 456558 558860 456564 558862
rect 456628 558860 456634 558924
rect 456793 558922 456859 558925
rect 457478 558922 457484 558924
rect 456793 558920 457484 558922
rect 456793 558864 456798 558920
rect 456854 558864 457484 558920
rect 456793 558862 457484 558864
rect 456793 558859 456859 558862
rect 457478 558860 457484 558862
rect 457548 558860 457554 558924
rect 458173 558922 458239 558925
rect 458766 558922 458772 558924
rect 458173 558920 458772 558922
rect 458173 558864 458178 558920
rect 458234 558864 458772 558920
rect 458173 558862 458772 558864
rect 458173 558859 458239 558862
rect 458766 558860 458772 558862
rect 458836 558860 458842 558924
rect 459553 558922 459619 558925
rect 461025 558924 461091 558925
rect 460054 558922 460060 558924
rect 459553 558920 460060 558922
rect 459553 558864 459558 558920
rect 459614 558864 460060 558920
rect 459553 558862 460060 558864
rect 459553 558859 459619 558862
rect 460054 558860 460060 558862
rect 460124 558860 460130 558924
rect 460974 558860 460980 558924
rect 461044 558922 461091 558924
rect 461669 558924 461735 558925
rect 461044 558920 461136 558922
rect 461086 558864 461136 558920
rect 461044 558862 461136 558864
rect 461669 558920 461716 558924
rect 461780 558922 461786 558924
rect 462313 558922 462379 558925
rect 463366 558922 463372 558924
rect 461669 558864 461674 558920
rect 461044 558860 461091 558862
rect 461025 558859 461091 558860
rect 461669 558860 461716 558864
rect 461780 558862 461826 558922
rect 462313 558920 463372 558922
rect 462313 558864 462318 558920
rect 462374 558864 463372 558920
rect 462313 558862 463372 558864
rect 461780 558860 461786 558862
rect 461669 558859 461735 558860
rect 462313 558859 462379 558862
rect 463366 558860 463372 558862
rect 463436 558860 463442 558924
rect 463693 558922 463759 558925
rect 464470 558922 464476 558924
rect 463693 558920 464476 558922
rect 463693 558864 463698 558920
rect 463754 558864 464476 558920
rect 463693 558862 464476 558864
rect 463693 558859 463759 558862
rect 464470 558860 464476 558862
rect 464540 558860 464546 558924
rect 465073 558922 465139 558925
rect 465758 558922 465764 558924
rect 465073 558920 465764 558922
rect 465073 558864 465078 558920
rect 465134 558864 465764 558920
rect 465073 558862 465764 558864
rect 465073 558859 465139 558862
rect 465758 558860 465764 558862
rect 465828 558860 465834 558924
rect 466453 558922 466519 558925
rect 466862 558922 466868 558924
rect 466453 558920 466868 558922
rect 466453 558864 466458 558920
rect 466514 558864 466868 558920
rect 466453 558862 466868 558864
rect 466453 558859 466519 558862
rect 466862 558860 466868 558862
rect 466932 558860 466938 558924
rect 467833 558922 467899 558925
rect 468753 558924 468819 558925
rect 467966 558922 467972 558924
rect 467833 558920 467972 558922
rect 467833 558864 467838 558920
rect 467894 558864 467972 558920
rect 467833 558862 467972 558864
rect 467833 558859 467899 558862
rect 467966 558860 467972 558862
rect 468036 558860 468042 558924
rect 468702 558922 468708 558924
rect 468662 558862 468708 558922
rect 468772 558920 468819 558924
rect 468814 558864 468819 558920
rect 468702 558860 468708 558862
rect 468772 558860 468819 558864
rect 468753 558859 468819 558860
rect 469213 558922 469279 558925
rect 470358 558922 470364 558924
rect 469213 558920 470364 558922
rect 469213 558864 469218 558920
rect 469274 558864 470364 558920
rect 469213 558862 470364 558864
rect 469213 558859 469279 558862
rect 470358 558860 470364 558862
rect 470428 558860 470434 558924
rect 470593 558922 470659 558925
rect 471462 558922 471468 558924
rect 470593 558920 471468 558922
rect 470593 558864 470598 558920
rect 470654 558864 471468 558920
rect 470593 558862 471468 558864
rect 470593 558859 470659 558862
rect 471462 558860 471468 558862
rect 471532 558860 471538 558924
rect 471973 558922 472039 558925
rect 472750 558922 472756 558924
rect 471973 558920 472756 558922
rect 471973 558864 471978 558920
rect 472034 558864 472756 558920
rect 471973 558862 472756 558864
rect 471973 558859 472039 558862
rect 472750 558860 472756 558862
rect 472820 558860 472826 558924
rect 473353 558922 473419 558925
rect 474038 558922 474044 558924
rect 473353 558920 474044 558922
rect 473353 558864 473358 558920
rect 473414 558864 474044 558920
rect 473353 558862 474044 558864
rect 473353 558859 473419 558862
rect 474038 558860 474044 558862
rect 474108 558860 474114 558924
rect 474733 558922 474799 558925
rect 475469 558924 475535 558925
rect 474958 558922 474964 558924
rect 474733 558920 474964 558922
rect 474733 558864 474738 558920
rect 474794 558864 474964 558920
rect 474733 558862 474964 558864
rect 474733 558859 474799 558862
rect 474958 558860 474964 558862
rect 475028 558860 475034 558924
rect 475469 558920 475516 558924
rect 475580 558922 475586 558924
rect 476113 558922 476179 558925
rect 476573 558924 476639 558925
rect 476246 558922 476252 558924
rect 475469 558864 475474 558920
rect 475469 558860 475516 558864
rect 475580 558862 475626 558922
rect 476113 558920 476252 558922
rect 476113 558864 476118 558920
rect 476174 558864 476252 558920
rect 476113 558862 476252 558864
rect 475580 558860 475586 558862
rect 475469 558859 475535 558860
rect 476113 558859 476179 558862
rect 476246 558860 476252 558862
rect 476316 558860 476322 558924
rect 476573 558920 476620 558924
rect 476684 558922 476690 558924
rect 477585 558922 477651 558925
rect 478965 558924 479031 558925
rect 477902 558922 477908 558924
rect 476573 558864 476578 558920
rect 476573 558860 476620 558864
rect 476684 558862 476730 558922
rect 477585 558920 477908 558922
rect 477585 558864 477590 558920
rect 477646 558864 477908 558920
rect 477585 558862 477908 558864
rect 476684 558860 476690 558862
rect 476573 558859 476639 558860
rect 477585 558859 477651 558862
rect 477902 558860 477908 558862
rect 477972 558860 477978 558924
rect 478965 558920 479012 558924
rect 479076 558922 479082 558924
rect 480345 558922 480411 558925
rect 480478 558922 480484 558924
rect 478965 558864 478970 558920
rect 478965 558860 479012 558864
rect 479076 558862 479122 558922
rect 480345 558920 480484 558922
rect 480345 558864 480350 558920
rect 480406 558864 480484 558920
rect 480345 558862 480484 558864
rect 479076 558860 479082 558862
rect 478965 558859 479031 558860
rect 480345 558859 480411 558862
rect 480478 558860 480484 558862
rect 480548 558860 480554 558924
rect 194409 558788 194475 558789
rect 217593 558788 217659 558789
rect 64270 558724 64276 558788
rect 64340 558786 64346 558788
rect 194358 558786 194364 558788
rect 64340 558726 194364 558786
rect 194428 558784 194475 558788
rect 217542 558786 217548 558788
rect 194470 558728 194475 558784
rect 64340 558724 64346 558726
rect 194358 558724 194364 558726
rect 194428 558724 194475 558728
rect 217502 558726 217548 558786
rect 217612 558784 217659 558788
rect 217654 558728 217659 558784
rect 217542 558724 217548 558726
rect 217612 558724 217659 558728
rect 194409 558723 194475 558724
rect 217593 558723 217659 558724
rect 223573 558788 223639 558789
rect 223573 558784 223620 558788
rect 223684 558786 223690 558788
rect 223573 558728 223578 558784
rect 223573 558724 223620 558728
rect 223684 558726 223730 558786
rect 223684 558724 223690 558726
rect 225638 558724 225644 558788
rect 225708 558786 225714 558788
rect 226241 558786 226307 558789
rect 231853 558788 231919 558789
rect 231853 558786 231900 558788
rect 225708 558784 226307 558786
rect 225708 558728 226246 558784
rect 226302 558728 226307 558784
rect 225708 558726 226307 558728
rect 231808 558784 231900 558786
rect 231808 558728 231858 558784
rect 231808 558726 231900 558728
rect 225708 558724 225714 558726
rect 223573 558723 223639 558724
rect 226241 558723 226307 558726
rect 231853 558724 231900 558726
rect 231964 558724 231970 558788
rect 232630 558724 232636 558788
rect 232700 558786 232706 558788
rect 233141 558786 233207 558789
rect 234613 558788 234679 558789
rect 234613 558786 234660 558788
rect 232700 558784 233207 558786
rect 232700 558728 233146 558784
rect 233202 558728 233207 558784
rect 232700 558726 233207 558728
rect 234568 558784 234660 558786
rect 234568 558728 234618 558784
rect 234568 558726 234660 558728
rect 232700 558724 232706 558726
rect 231853 558723 231919 558724
rect 233141 558723 233207 558726
rect 234613 558724 234660 558726
rect 234724 558724 234730 558788
rect 235993 558786 236059 558789
rect 237373 558788 237439 558789
rect 236126 558786 236132 558788
rect 235993 558784 236132 558786
rect 235993 558728 235998 558784
rect 236054 558728 236132 558784
rect 235993 558726 236132 558728
rect 234613 558723 234679 558724
rect 235993 558723 236059 558726
rect 236126 558724 236132 558726
rect 236196 558724 236202 558788
rect 237373 558786 237420 558788
rect 237328 558784 237420 558786
rect 237328 558728 237378 558784
rect 237328 558726 237420 558728
rect 237373 558724 237420 558726
rect 237484 558724 237490 558788
rect 320265 558786 320331 558789
rect 320950 558786 320956 558788
rect 320265 558784 320956 558786
rect 320265 558728 320270 558784
rect 320326 558728 320956 558784
rect 320265 558726 320956 558728
rect 237373 558723 237439 558724
rect 320265 558723 320331 558726
rect 320950 558724 320956 558726
rect 321020 558724 321026 558788
rect 322197 558786 322263 558789
rect 322606 558786 322612 558788
rect 322197 558784 322612 558786
rect 322197 558728 322202 558784
rect 322258 558728 322612 558784
rect 322197 558726 322612 558728
rect 322197 558723 322263 558726
rect 322606 558724 322612 558726
rect 322676 558724 322682 558788
rect 326102 558724 326108 558788
rect 326172 558786 326178 558788
rect 326337 558786 326403 558789
rect 326172 558784 326403 558786
rect 326172 558728 326342 558784
rect 326398 558728 326403 558784
rect 326172 558726 326403 558728
rect 326172 558724 326178 558726
rect 326337 558723 326403 558726
rect 328453 558786 328519 558789
rect 330477 558788 330543 558789
rect 333145 558788 333211 558789
rect 334065 558788 334131 558789
rect 328862 558786 328868 558788
rect 328453 558784 328868 558786
rect 328453 558728 328458 558784
rect 328514 558728 328868 558784
rect 328453 558726 328868 558728
rect 328453 558723 328519 558726
rect 328862 558724 328868 558726
rect 328932 558724 328938 558788
rect 330477 558784 330524 558788
rect 330588 558786 330594 558788
rect 333094 558786 333100 558788
rect 330477 558728 330482 558784
rect 330477 558724 330524 558728
rect 330588 558726 330634 558786
rect 333054 558726 333100 558786
rect 333164 558784 333211 558788
rect 334014 558786 334020 558788
rect 333206 558728 333211 558784
rect 330588 558724 330594 558726
rect 333094 558724 333100 558726
rect 333164 558724 333211 558728
rect 333974 558726 334020 558786
rect 334084 558784 334131 558788
rect 334126 558728 334131 558784
rect 334014 558724 334020 558726
rect 334084 558724 334131 558728
rect 330477 558723 330543 558724
rect 333145 558723 333211 558724
rect 334065 558723 334131 558724
rect 335445 558788 335511 558789
rect 336641 558788 336707 558789
rect 335445 558784 335492 558788
rect 335556 558786 335562 558788
rect 336590 558786 336596 558788
rect 335445 558728 335450 558784
rect 335445 558724 335492 558728
rect 335556 558726 335602 558786
rect 336550 558726 336596 558786
rect 336660 558784 336707 558788
rect 336702 558728 336707 558784
rect 335556 558724 335562 558726
rect 336590 558724 336596 558726
rect 336660 558724 336707 558728
rect 335445 558723 335511 558724
rect 336641 558723 336707 558724
rect 336825 558786 336891 558789
rect 339033 558788 339099 558789
rect 337878 558786 337884 558788
rect 336825 558784 337884 558786
rect 336825 558728 336830 558784
rect 336886 558728 337884 558784
rect 336825 558726 337884 558728
rect 336825 558723 336891 558726
rect 337878 558724 337884 558726
rect 337948 558724 337954 558788
rect 338982 558786 338988 558788
rect 338942 558726 338988 558786
rect 339052 558784 339099 558788
rect 339094 558728 339099 558784
rect 338982 558724 338988 558726
rect 339052 558724 339099 558728
rect 339033 558723 339099 558724
rect 339861 558788 339927 558789
rect 341241 558788 341307 558789
rect 342529 558788 342595 558789
rect 343633 558788 343699 558789
rect 346025 558788 346091 558789
rect 339861 558784 339908 558788
rect 339972 558786 339978 558788
rect 341190 558786 341196 558788
rect 339861 558728 339866 558784
rect 339861 558724 339908 558728
rect 339972 558726 340018 558786
rect 341150 558726 341196 558786
rect 341260 558784 341307 558788
rect 342478 558786 342484 558788
rect 341302 558728 341307 558784
rect 339972 558724 339978 558726
rect 341190 558724 341196 558726
rect 341260 558724 341307 558728
rect 342438 558726 342484 558786
rect 342548 558784 342595 558788
rect 343582 558786 343588 558788
rect 342590 558728 342595 558784
rect 342478 558724 342484 558726
rect 342548 558724 342595 558728
rect 343542 558726 343588 558786
rect 343652 558784 343699 558788
rect 345974 558786 345980 558788
rect 343694 558728 343699 558784
rect 343582 558724 343588 558726
rect 343652 558724 343699 558728
rect 345934 558726 345980 558786
rect 346044 558784 346091 558788
rect 346086 558728 346091 558784
rect 345974 558724 345980 558726
rect 346044 558724 346091 558728
rect 346894 558724 346900 558788
rect 346964 558786 346970 558788
rect 347681 558786 347747 558789
rect 348233 558788 348299 558789
rect 348182 558786 348188 558788
rect 346964 558784 347747 558786
rect 346964 558728 347686 558784
rect 347742 558728 347747 558784
rect 346964 558726 347747 558728
rect 348142 558726 348188 558786
rect 348252 558784 348299 558788
rect 348294 558728 348299 558784
rect 346964 558724 346970 558726
rect 339861 558723 339927 558724
rect 341241 558723 341307 558724
rect 342529 558723 342595 558724
rect 343633 558723 343699 558724
rect 346025 558723 346091 558724
rect 347681 558723 347747 558726
rect 348182 558724 348188 558726
rect 348252 558724 348299 558728
rect 349470 558724 349476 558788
rect 349540 558786 349546 558788
rect 349705 558786 349771 558789
rect 349540 558784 349771 558786
rect 349540 558728 349710 558784
rect 349766 558728 349771 558784
rect 349540 558726 349771 558728
rect 349540 558724 349546 558726
rect 348233 558723 348299 558724
rect 349705 558723 349771 558726
rect 353293 558786 353359 558789
rect 353518 558786 353524 558788
rect 353293 558784 353524 558786
rect 353293 558728 353298 558784
rect 353354 558728 353524 558784
rect 353293 558726 353524 558728
rect 353293 558723 353359 558726
rect 353518 558724 353524 558726
rect 353588 558724 353594 558788
rect 354673 558786 354739 558789
rect 354806 558786 354812 558788
rect 354673 558784 354812 558786
rect 354673 558728 354678 558784
rect 354734 558728 354812 558784
rect 354673 558726 354812 558728
rect 354673 558723 354739 558726
rect 354806 558724 354812 558726
rect 354876 558724 354882 558788
rect 452745 558786 452811 558789
rect 454769 558788 454835 558789
rect 456057 558788 456123 558789
rect 453798 558786 453804 558788
rect 452745 558784 453804 558786
rect 452745 558728 452750 558784
rect 452806 558728 453804 558784
rect 452745 558726 453804 558728
rect 452745 558723 452811 558726
rect 453798 558724 453804 558726
rect 453868 558724 453874 558788
rect 454718 558786 454724 558788
rect 454678 558726 454724 558786
rect 454788 558784 454835 558788
rect 454830 558728 454835 558784
rect 454718 558724 454724 558726
rect 454788 558724 454835 558728
rect 456006 558724 456012 558788
rect 456076 558786 456123 558788
rect 456076 558784 456168 558786
rect 456118 558728 456168 558784
rect 456076 558726 456168 558728
rect 456076 558724 456123 558726
rect 457294 558724 457300 558788
rect 457364 558786 457370 558788
rect 457437 558786 457503 558789
rect 457364 558784 457503 558786
rect 457364 558728 457442 558784
rect 457498 558728 457503 558784
rect 457364 558726 457503 558728
rect 457364 558724 457370 558726
rect 454769 558723 454835 558724
rect 456057 558723 456123 558724
rect 457437 558723 457503 558726
rect 458398 558724 458404 558788
rect 458468 558786 458474 558788
rect 458817 558786 458883 558789
rect 458468 558784 458883 558786
rect 458468 558728 458822 558784
rect 458878 558728 458883 558784
rect 458468 558726 458883 558728
rect 458468 558724 458474 558726
rect 458817 558723 458883 558726
rect 460933 558786 460999 558789
rect 463049 558788 463115 558789
rect 462078 558786 462084 558788
rect 460933 558784 462084 558786
rect 460933 558728 460938 558784
rect 460994 558728 462084 558784
rect 460933 558726 462084 558728
rect 460933 558723 460999 558726
rect 462078 558724 462084 558726
rect 462148 558724 462154 558788
rect 462998 558786 463004 558788
rect 462958 558726 463004 558786
rect 463068 558784 463115 558788
rect 463110 558728 463115 558784
rect 462998 558724 463004 558726
rect 463068 558724 463115 558728
rect 463049 558723 463115 558724
rect 464245 558788 464311 558789
rect 465257 558788 465323 558789
rect 466545 558788 466611 558789
rect 464245 558784 464292 558788
rect 464356 558786 464362 558788
rect 465206 558786 465212 558788
rect 464245 558728 464250 558784
rect 464245 558724 464292 558728
rect 464356 558726 464402 558786
rect 465166 558726 465212 558786
rect 465276 558784 465323 558788
rect 466494 558786 466500 558788
rect 465318 558728 465323 558784
rect 464356 558724 464362 558726
rect 465206 558724 465212 558726
rect 465276 558724 465323 558728
rect 466454 558726 466500 558786
rect 466564 558784 466611 558788
rect 466606 558728 466611 558784
rect 466494 558724 466500 558726
rect 466564 558724 466611 558728
rect 464245 558723 464311 558724
rect 465257 558723 465323 558724
rect 466545 558723 466611 558724
rect 467925 558786 467991 558789
rect 471329 558788 471395 558789
rect 469070 558786 469076 558788
rect 467925 558784 469076 558786
rect 467925 558728 467930 558784
rect 467986 558728 469076 558784
rect 467925 558726 469076 558728
rect 467925 558723 467991 558726
rect 469070 558724 469076 558726
rect 469140 558724 469146 558788
rect 471278 558786 471284 558788
rect 471238 558726 471284 558786
rect 471348 558784 471395 558788
rect 471390 558728 471395 558784
rect 471278 558724 471284 558726
rect 471348 558724 471395 558728
rect 471329 558723 471395 558724
rect 472157 558788 472223 558789
rect 473445 558788 473511 558789
rect 474825 558788 474891 558789
rect 472157 558784 472204 558788
rect 472268 558786 472274 558788
rect 472157 558728 472162 558784
rect 472157 558724 472204 558728
rect 472268 558726 472314 558786
rect 473445 558784 473492 558788
rect 473556 558786 473562 558788
rect 474774 558786 474780 558788
rect 473445 558728 473450 558784
rect 472268 558724 472274 558726
rect 473445 558724 473492 558728
rect 473556 558726 473602 558786
rect 474734 558726 474780 558786
rect 474844 558784 474891 558788
rect 474886 558728 474891 558784
rect 473556 558724 473562 558726
rect 474774 558724 474780 558726
rect 474844 558724 474891 558728
rect 472157 558723 472223 558724
rect 473445 558723 473511 558724
rect 474825 558723 474891 558724
rect 484393 558786 484459 558789
rect 484710 558786 484716 558788
rect 484393 558784 484716 558786
rect 484393 558728 484398 558784
rect 484454 558728 484716 558784
rect 484393 558726 484716 558728
rect 484393 558723 484459 558726
rect 484710 558724 484716 558726
rect 484780 558724 484786 558788
rect 69790 558588 69796 558652
rect 69860 558650 69866 558652
rect 70209 558650 70275 558653
rect 75913 558652 75979 558653
rect 78489 558652 78555 558653
rect 79409 558652 79475 558653
rect 75862 558650 75868 558652
rect 69860 558648 70275 558650
rect 69860 558592 70214 558648
rect 70270 558592 70275 558648
rect 69860 558590 70275 558592
rect 75822 558590 75868 558650
rect 75932 558648 75979 558652
rect 78438 558650 78444 558652
rect 75974 558592 75979 558648
rect 69860 558588 69866 558590
rect 70209 558587 70275 558590
rect 75862 558588 75868 558590
rect 75932 558588 75979 558592
rect 78398 558590 78444 558650
rect 78508 558648 78555 558652
rect 79358 558650 79364 558652
rect 78550 558592 78555 558648
rect 78438 558588 78444 558590
rect 78508 558588 78555 558592
rect 79318 558590 79364 558650
rect 79428 558648 79475 558652
rect 79470 558592 79475 558648
rect 79358 558588 79364 558590
rect 79428 558588 79475 558592
rect 75913 558587 75979 558588
rect 78489 558587 78555 558588
rect 79409 558587 79475 558588
rect 85389 558652 85455 558653
rect 85389 558648 85436 558652
rect 85500 558650 85506 558652
rect 85389 558592 85394 558648
rect 85389 558588 85436 558592
rect 85500 558590 85546 558650
rect 85500 558588 85506 558590
rect 86166 558588 86172 558652
rect 86236 558650 86242 558652
rect 86861 558650 86927 558653
rect 86236 558648 86927 558650
rect 86236 558592 86866 558648
rect 86922 558592 86927 558648
rect 86236 558590 86927 558592
rect 86236 558588 86242 558590
rect 85389 558587 85455 558588
rect 86861 558587 86927 558590
rect 91093 558652 91159 558653
rect 91093 558648 91140 558652
rect 91204 558650 91210 558652
rect 91093 558592 91098 558648
rect 91093 558588 91140 558592
rect 91204 558590 91250 558650
rect 91204 558588 91210 558590
rect 93158 558588 93164 558652
rect 93228 558650 93234 558652
rect 93669 558650 93735 558653
rect 93228 558648 93735 558650
rect 93228 558592 93674 558648
rect 93730 558592 93735 558648
rect 93228 558590 93735 558592
rect 93228 558588 93234 558590
rect 91093 558587 91159 558588
rect 93669 558587 93735 558590
rect 94773 558652 94839 558653
rect 106273 558652 106339 558653
rect 94773 558648 94820 558652
rect 94884 558650 94890 558652
rect 94773 558592 94778 558648
rect 94773 558588 94820 558592
rect 94884 558590 94930 558650
rect 94884 558588 94890 558590
rect 106222 558588 106228 558652
rect 106292 558650 106339 558652
rect 202137 558650 202203 558653
rect 204897 558652 204963 558653
rect 202454 558650 202460 558652
rect 106292 558648 106384 558650
rect 106334 558592 106384 558648
rect 106292 558590 106384 558592
rect 202137 558648 202460 558650
rect 202137 558592 202142 558648
rect 202198 558592 202460 558648
rect 202137 558590 202460 558592
rect 106292 558588 106339 558590
rect 94773 558587 94839 558588
rect 106273 558587 106339 558588
rect 202137 558587 202203 558590
rect 202454 558588 202460 558590
rect 202524 558588 202530 558652
rect 204846 558650 204852 558652
rect 204806 558590 204852 558650
rect 204916 558648 204963 558652
rect 204958 558592 204963 558648
rect 204846 558588 204852 558590
rect 204916 558588 204963 558592
rect 204897 558587 204963 558588
rect 209037 558650 209103 558653
rect 323577 558652 323643 558653
rect 209630 558650 209636 558652
rect 209037 558648 209636 558650
rect 209037 558592 209042 558648
rect 209098 558592 209636 558648
rect 209037 558590 209636 558592
rect 209037 558587 209103 558590
rect 209630 558588 209636 558590
rect 209700 558588 209706 558652
rect 323526 558588 323532 558652
rect 323596 558650 323643 558652
rect 323596 558648 323688 558650
rect 323638 558592 323688 558648
rect 323596 558590 323688 558592
rect 323596 558588 323643 558590
rect 324814 558588 324820 558652
rect 324884 558650 324890 558652
rect 324957 558650 325023 558653
rect 324884 558648 325023 558650
rect 324884 558592 324962 558648
rect 325018 558592 325023 558648
rect 324884 558590 325023 558592
rect 324884 558588 324890 558590
rect 323577 558587 323643 558588
rect 324957 558587 325023 558590
rect 327022 558588 327028 558652
rect 327092 558650 327098 558652
rect 327717 558650 327783 558653
rect 327092 558648 327783 558650
rect 327092 558592 327722 558648
rect 327778 558592 327783 558648
rect 327092 558590 327783 558592
rect 327092 558588 327098 558590
rect 327717 558587 327783 558590
rect 328494 558588 328500 558652
rect 328564 558650 328570 558652
rect 329097 558650 329163 558653
rect 328564 558648 329163 558650
rect 328564 558592 329102 558648
rect 329158 558592 329163 558648
rect 328564 558590 329163 558592
rect 328564 558588 328570 558590
rect 329097 558587 329163 558590
rect 452694 558588 452700 558652
rect 452764 558650 452770 558652
rect 453297 558650 453363 558653
rect 452764 558648 453363 558650
rect 452764 558592 453302 558648
rect 453358 558592 453363 558648
rect 452764 558590 453363 558592
rect 452764 558588 452770 558590
rect 453297 558587 453363 558590
rect 459502 558588 459508 558652
rect 459572 558650 459578 558652
rect 460381 558650 460447 558653
rect 459572 558648 460447 558650
rect 459572 558592 460386 558648
rect 460442 558592 460447 558648
rect 459572 558590 460447 558592
rect 459572 558588 459578 558590
rect 460381 558587 460447 558590
rect 467782 558588 467788 558652
rect 467852 558650 467858 558652
rect 468017 558650 468083 558653
rect 470041 558652 470107 558653
rect 469990 558650 469996 558652
rect 467852 558648 468083 558650
rect 467852 558592 468022 558648
rect 468078 558592 468083 558648
rect 467852 558590 468083 558592
rect 469950 558590 469996 558650
rect 470060 558648 470107 558652
rect 470102 558592 470107 558648
rect 467852 558588 467858 558590
rect 468017 558587 468083 558590
rect 469990 558588 469996 558590
rect 470060 558588 470107 558592
rect 470041 558587 470107 558588
rect 476205 558650 476271 558653
rect 481633 558652 481699 558653
rect 477350 558650 477356 558652
rect 476205 558648 477356 558650
rect 476205 558592 476210 558648
rect 476266 558592 477356 558648
rect 476205 558590 477356 558592
rect 476205 558587 476271 558590
rect 477350 558588 477356 558590
rect 477420 558588 477426 558652
rect 481582 558588 481588 558652
rect 481652 558650 481699 558652
rect 481652 558648 481744 558650
rect 481694 558592 481744 558648
rect 481652 558590 481744 558592
rect 481652 558588 481699 558590
rect 481633 558587 481699 558588
rect 99465 558514 99531 558517
rect 99598 558514 99604 558516
rect 99465 558512 99604 558514
rect 99465 558456 99470 558512
rect 99526 558456 99604 558512
rect 99465 558454 99604 558456
rect 99465 558451 99531 558454
rect 99598 558452 99604 558454
rect 99668 558514 99674 558516
rect 100385 558514 100451 558517
rect 99668 558512 100451 558514
rect 99668 558456 100390 558512
rect 100446 558456 100451 558512
rect 99668 558454 100451 558456
rect 99668 558452 99674 558454
rect 100385 558451 100451 558454
rect 108481 558514 108547 558517
rect 108614 558514 108620 558516
rect 108481 558512 108620 558514
rect 108481 558456 108486 558512
rect 108542 558456 108620 558512
rect 108481 558454 108620 558456
rect 108481 558451 108547 558454
rect 108614 558452 108620 558454
rect 108684 558452 108690 558516
rect 108982 558452 108988 558516
rect 109052 558514 109058 558516
rect 110321 558514 110387 558517
rect 109052 558512 110387 558514
rect 109052 558456 110326 558512
rect 110382 558456 110387 558512
rect 109052 558454 110387 558456
rect 109052 558452 109058 558454
rect 110321 558451 110387 558454
rect 231853 558514 231919 558517
rect 350533 558516 350599 558517
rect 232814 558514 232820 558516
rect 231853 558512 232820 558514
rect 231853 558456 231858 558512
rect 231914 558456 232820 558512
rect 231853 558454 232820 558456
rect 231853 558451 231919 558454
rect 232814 558452 232820 558454
rect 232884 558452 232890 558516
rect 350533 558512 350580 558516
rect 350644 558514 350650 558516
rect 357433 558514 357499 558517
rect 357566 558514 357572 558516
rect 350533 558456 350538 558512
rect 350533 558452 350580 558456
rect 350644 558454 350690 558514
rect 357433 558512 357572 558514
rect 357433 558456 357438 558512
rect 357494 558456 357572 558512
rect 357433 558454 357572 558456
rect 350644 558452 350650 558454
rect 350533 558451 350599 558452
rect 357433 558451 357499 558454
rect 357566 558452 357572 558454
rect 357636 558452 357642 558516
rect 478873 558514 478939 558517
rect 479742 558514 479748 558516
rect 478873 558512 479748 558514
rect 478873 558456 478878 558512
rect 478934 558456 479748 558512
rect 478873 558454 479748 558456
rect 478873 558451 478939 558454
rect 479742 558452 479748 558454
rect 479812 558452 479818 558516
rect 481633 558514 481699 558517
rect 483013 558516 483079 558517
rect 482134 558514 482140 558516
rect 481633 558512 482140 558514
rect 481633 558456 481638 558512
rect 481694 558456 482140 558512
rect 481633 558454 482140 558456
rect 481633 558451 481699 558454
rect 482134 558452 482140 558454
rect 482204 558452 482210 558516
rect 483013 558514 483060 558516
rect 482968 558512 483060 558514
rect 482968 558456 483018 558512
rect 482968 558454 483060 558456
rect 483013 558452 483060 558454
rect 483124 558452 483130 558516
rect 485773 558514 485839 558517
rect 485998 558514 486004 558516
rect 485773 558512 486004 558514
rect 485773 558456 485778 558512
rect 485834 558456 486004 558512
rect 485773 558454 486004 558456
rect 483013 558451 483079 558452
rect 485773 558451 485839 558454
rect 485998 558452 486004 558454
rect 486068 558452 486074 558516
rect 487153 558514 487219 558517
rect 487286 558514 487292 558516
rect 487153 558512 487292 558514
rect 487153 558456 487158 558512
rect 487214 558456 487292 558512
rect 487153 558454 487292 558456
rect 487153 558451 487219 558454
rect 487286 558452 487292 558454
rect 487356 558452 487362 558516
rect 62021 558378 62087 558381
rect 197302 558378 197308 558380
rect 62021 558376 197308 558378
rect 62021 558320 62026 558376
rect 62082 558320 197308 558376
rect 62021 558318 197308 558320
rect 62021 558315 62087 558318
rect 197302 558316 197308 558318
rect 197372 558316 197378 558380
rect 230473 558378 230539 558381
rect 238753 558380 238819 558381
rect 230606 558378 230612 558380
rect 230473 558376 230612 558378
rect 230473 558320 230478 558376
rect 230534 558320 230612 558376
rect 230473 558318 230612 558320
rect 230473 558315 230539 558318
rect 230606 558316 230612 558318
rect 230676 558316 230682 558380
rect 238702 558316 238708 558380
rect 238772 558378 238819 558380
rect 238772 558376 238864 558378
rect 238814 558320 238864 558376
rect 238772 558318 238864 558320
rect 238772 558316 238819 558318
rect 282310 558316 282316 558380
rect 282380 558378 282386 558380
rect 447358 558378 447364 558380
rect 282380 558318 447364 558378
rect 282380 558316 282386 558318
rect 447358 558316 447364 558318
rect 447428 558316 447434 558380
rect 477493 558378 477559 558381
rect 478454 558378 478460 558380
rect 477493 558376 478460 558378
rect 477493 558320 477498 558376
rect 477554 558320 478460 558376
rect 477493 558318 478460 558320
rect 238753 558315 238819 558316
rect 477493 558315 477559 558318
rect 478454 558316 478460 558318
rect 478524 558316 478530 558380
rect 480345 558378 480411 558381
rect 488533 558380 488599 558381
rect 480846 558378 480852 558380
rect 480345 558376 480852 558378
rect 480345 558320 480350 558376
rect 480406 558320 480852 558376
rect 480345 558318 480852 558320
rect 480345 558315 480411 558318
rect 480846 558316 480852 558318
rect 480916 558316 480922 558380
rect 488533 558378 488580 558380
rect 488488 558376 488580 558378
rect 488488 558320 488538 558376
rect 488488 558318 488580 558320
rect 488533 558316 488580 558318
rect 488644 558316 488650 558380
rect 488533 558315 488599 558316
rect 63401 558242 63467 558245
rect 198774 558242 198780 558244
rect 63401 558240 198780 558242
rect 63401 558184 63406 558240
rect 63462 558184 198780 558240
rect 63401 558182 198780 558184
rect 63401 558179 63467 558182
rect 198774 558180 198780 558182
rect 198844 558180 198850 558244
rect 283414 558180 283420 558244
rect 283484 558242 283490 558244
rect 448462 558242 448468 558244
rect 283484 558182 448468 558242
rect 283484 558180 283490 558182
rect 448462 558180 448468 558182
rect 448532 558180 448538 558244
rect 483013 558242 483079 558245
rect 484158 558242 484164 558244
rect 483013 558240 484164 558242
rect 483013 558184 483018 558240
rect 483074 558184 484164 558240
rect 483013 558182 484164 558184
rect 483013 558179 483079 558182
rect 484158 558180 484164 558182
rect 484228 558180 484234 558244
rect 238334 558044 238340 558108
rect 238404 558106 238410 558108
rect 238661 558106 238727 558109
rect 238404 558104 238727 558106
rect 238404 558048 238666 558104
rect 238722 558048 238727 558104
rect 238404 558046 238727 558048
rect 238404 558044 238410 558046
rect 238661 558043 238727 558046
rect 321553 558106 321619 558109
rect 322790 558106 322796 558108
rect 321553 558104 322796 558106
rect 321553 558048 321558 558104
rect 321614 558048 322796 558104
rect 321553 558046 322796 558048
rect 321553 558043 321619 558046
rect 322790 558044 322796 558046
rect 322860 558044 322866 558108
rect 322933 558106 322999 558109
rect 324078 558106 324084 558108
rect 322933 558104 324084 558106
rect 322933 558048 322938 558104
rect 322994 558048 324084 558104
rect 322933 558046 324084 558048
rect 322933 558043 322999 558046
rect 324078 558044 324084 558046
rect 324148 558044 324154 558108
rect 484393 558106 484459 558109
rect 485630 558106 485636 558108
rect 484393 558104 485636 558106
rect 484393 558048 484398 558104
rect 484454 558048 485636 558104
rect 484393 558046 485636 558048
rect 484393 558043 484459 558046
rect 485630 558044 485636 558046
rect 485700 558044 485706 558108
rect 82721 557972 82787 557973
rect 82670 557908 82676 557972
rect 82740 557970 82787 557972
rect 82740 557968 82832 557970
rect 82782 557912 82832 557968
rect 82740 557910 82832 557912
rect 82740 557908 82787 557910
rect 107694 557908 107700 557972
rect 107764 557970 107770 557972
rect 108297 557970 108363 557973
rect 329833 557972 329899 557973
rect 107764 557968 108363 557970
rect 107764 557912 108302 557968
rect 108358 557912 108363 557968
rect 107764 557910 108363 557912
rect 107764 557908 107770 557910
rect 82721 557907 82787 557908
rect 108297 557907 108363 557910
rect 329782 557908 329788 557972
rect 329852 557970 329899 557972
rect 483013 557970 483079 557973
rect 483422 557970 483428 557972
rect 329852 557968 329944 557970
rect 329894 557912 329944 557968
rect 329852 557910 329944 557912
rect 483013 557968 483428 557970
rect 483013 557912 483018 557968
rect 483074 557912 483428 557968
rect 483013 557910 483428 557912
rect 329852 557908 329899 557910
rect 329833 557907 329899 557908
rect 483013 557907 483079 557910
rect 483422 557908 483428 557910
rect 483492 557908 483498 557972
rect 485773 557970 485839 557973
rect 486918 557970 486924 557972
rect 485773 557968 486924 557970
rect 485773 557912 485778 557968
rect 485834 557912 486924 557968
rect 485773 557910 486924 557912
rect 485773 557907 485839 557910
rect 486918 557908 486924 557910
rect 486988 557908 486994 557972
rect 100845 557834 100911 557837
rect 101397 557834 101463 557837
rect 316309 557836 316375 557837
rect 101622 557834 101628 557836
rect 100845 557832 101628 557834
rect 100845 557776 100850 557832
rect 100906 557776 101402 557832
rect 101458 557776 101628 557832
rect 100845 557774 101628 557776
rect 100845 557771 100911 557774
rect 101397 557771 101463 557774
rect 101622 557772 101628 557774
rect 101692 557772 101698 557836
rect 316309 557834 316356 557836
rect 316264 557832 316356 557834
rect 316264 557776 316314 557832
rect 316264 557774 316356 557776
rect 316309 557772 316356 557774
rect 316420 557772 316426 557836
rect 331213 557834 331279 557837
rect 449893 557836 449959 557837
rect 332358 557834 332364 557836
rect 331213 557832 332364 557834
rect 331213 557776 331218 557832
rect 331274 557776 332364 557832
rect 331213 557774 332364 557776
rect 316309 557771 316375 557772
rect 331213 557771 331279 557774
rect 332358 557772 332364 557774
rect 332428 557772 332434 557836
rect 449893 557834 449940 557836
rect 449848 557832 449940 557834
rect 449848 557776 449898 557832
rect 449848 557774 449940 557776
rect 449893 557772 449940 557774
rect 450004 557772 450010 557836
rect 483013 557834 483079 557837
rect 483606 557834 483612 557836
rect 483013 557832 483612 557834
rect 483013 557776 483018 557832
rect 483074 557776 483612 557832
rect 483013 557774 483612 557776
rect 449893 557771 449959 557772
rect 483013 557771 483079 557774
rect 483606 557772 483612 557774
rect 483676 557772 483682 557836
rect 487153 557834 487219 557837
rect 487838 557834 487844 557836
rect 487153 557832 487844 557834
rect 487153 557776 487158 557832
rect 487214 557776 487844 557832
rect 487153 557774 487844 557776
rect 487153 557771 487219 557774
rect 487838 557772 487844 557774
rect 487908 557772 487914 557836
rect 100017 557698 100083 557701
rect 100150 557698 100156 557700
rect 100017 557696 100156 557698
rect 100017 557640 100022 557696
rect 100078 557640 100156 557696
rect 100017 557638 100156 557640
rect 100017 557635 100083 557638
rect 100150 557636 100156 557638
rect 100220 557636 100226 557700
rect 106222 557636 106228 557700
rect 106292 557698 106298 557700
rect 106917 557698 106983 557701
rect 201493 557700 201559 557701
rect 201493 557698 201540 557700
rect 106292 557696 106983 557698
rect 106292 557640 106922 557696
rect 106978 557640 106983 557696
rect 106292 557638 106983 557640
rect 201448 557696 201540 557698
rect 201448 557640 201498 557696
rect 201448 557638 201540 557640
rect 106292 557636 106298 557638
rect 106917 557635 106983 557638
rect 201493 557636 201540 557638
rect 201604 557636 201610 557700
rect 207054 557636 207060 557700
rect 207124 557698 207130 557700
rect 207657 557698 207723 557701
rect 207124 557696 207723 557698
rect 207124 557640 207662 557696
rect 207718 557640 207723 557696
rect 207124 557638 207723 557640
rect 207124 557636 207130 557638
rect 201493 557635 201559 557636
rect 207657 557635 207723 557638
rect 210366 557636 210372 557700
rect 210436 557698 210442 557700
rect 211061 557698 211127 557701
rect 210436 557696 211127 557698
rect 210436 557640 211066 557696
rect 211122 557640 211127 557696
rect 210436 557638 211127 557640
rect 210436 557636 210442 557638
rect 211061 557635 211127 557638
rect 217358 557636 217364 557700
rect 217428 557698 217434 557700
rect 217961 557698 218027 557701
rect 217428 557696 218027 557698
rect 217428 557640 217966 557696
rect 218022 557640 218027 557696
rect 217428 557638 218027 557640
rect 217428 557636 217434 557638
rect 217961 557635 218027 557638
rect 324313 557698 324379 557701
rect 325366 557698 325372 557700
rect 324313 557696 325372 557698
rect 324313 557640 324318 557696
rect 324374 557640 325372 557696
rect 324313 557638 325372 557640
rect 324313 557635 324379 557638
rect 325366 557636 325372 557638
rect 325436 557636 325442 557700
rect 343633 557698 343699 557701
rect 344870 557698 344876 557700
rect 343633 557696 344876 557698
rect 343633 557640 343638 557696
rect 343694 557640 344876 557696
rect 343633 557638 344876 557640
rect 343633 557635 343699 557638
rect 344870 557636 344876 557638
rect 344940 557636 344946 557700
rect 352097 557698 352163 557701
rect 460841 557700 460907 557701
rect 353150 557698 353156 557700
rect 352097 557696 353156 557698
rect 352097 557640 352102 557696
rect 352158 557640 353156 557696
rect 352097 557638 353156 557640
rect 352097 557635 352163 557638
rect 353150 557636 353156 557638
rect 353220 557636 353226 557700
rect 460790 557698 460796 557700
rect 460750 557638 460796 557698
rect 460860 557696 460907 557700
rect 460902 557640 460907 557696
rect 460790 557636 460796 557638
rect 460860 557636 460907 557640
rect 460841 557635 460907 557636
rect 488533 557698 488599 557701
rect 489126 557698 489132 557700
rect 488533 557696 489132 557698
rect 488533 557640 488538 557696
rect 488594 557640 489132 557696
rect 488533 557638 489132 557640
rect 488533 557635 488599 557638
rect 489126 557636 489132 557638
rect 489196 557636 489202 557700
rect 101438 557500 101444 557564
rect 101508 557562 101514 557564
rect 102041 557562 102107 557565
rect 102777 557564 102843 557565
rect 102726 557562 102732 557564
rect 101508 557560 102107 557562
rect 101508 557504 102046 557560
rect 102102 557504 102107 557560
rect 101508 557502 102107 557504
rect 102686 557502 102732 557562
rect 102796 557560 102843 557564
rect 102838 557504 102843 557560
rect 101508 557500 101514 557502
rect 102041 557499 102107 557502
rect 102726 557500 102732 557502
rect 102796 557500 102843 557504
rect 103278 557500 103284 557564
rect 103348 557562 103354 557564
rect 103421 557562 103487 557565
rect 103348 557560 103487 557562
rect 103348 557504 103426 557560
rect 103482 557504 103487 557560
rect 103348 557502 103487 557504
rect 103348 557500 103354 557502
rect 102777 557499 102843 557500
rect 103421 557499 103487 557502
rect 104014 557500 104020 557564
rect 104084 557562 104090 557564
rect 104157 557562 104223 557565
rect 104084 557560 104223 557562
rect 104084 557504 104162 557560
rect 104218 557504 104223 557560
rect 104084 557502 104223 557504
rect 104084 557500 104090 557502
rect 104157 557499 104223 557502
rect 105302 557500 105308 557564
rect 105372 557562 105378 557564
rect 105537 557562 105603 557565
rect 105372 557560 105603 557562
rect 105372 557504 105542 557560
rect 105598 557504 105603 557560
rect 105372 557502 105603 557504
rect 105372 557500 105378 557502
rect 105537 557499 105603 557502
rect 106038 557500 106044 557564
rect 106108 557562 106114 557564
rect 106181 557562 106247 557565
rect 206921 557564 206987 557565
rect 106108 557560 106247 557562
rect 106108 557504 106186 557560
rect 106242 557504 106247 557560
rect 106108 557502 106247 557504
rect 106108 557500 106114 557502
rect 106181 557499 106247 557502
rect 206870 557500 206876 557564
rect 206940 557562 206987 557564
rect 206940 557560 207032 557562
rect 206982 557504 207032 557560
rect 206940 557502 207032 557504
rect 206940 557500 206987 557502
rect 207974 557500 207980 557564
rect 208044 557562 208050 557564
rect 208301 557562 208367 557565
rect 208044 557560 208367 557562
rect 208044 557504 208306 557560
rect 208362 557504 208367 557560
rect 208044 557502 208367 557504
rect 208044 557500 208050 557502
rect 206921 557499 206987 557500
rect 208301 557499 208367 557502
rect 209262 557500 209268 557564
rect 209332 557562 209338 557564
rect 209681 557562 209747 557565
rect 212441 557564 212507 557565
rect 209332 557560 209747 557562
rect 209332 557504 209686 557560
rect 209742 557504 209747 557560
rect 209332 557502 209747 557504
rect 209332 557500 209338 557502
rect 209681 557499 209747 557502
rect 212390 557500 212396 557564
rect 212460 557562 212507 557564
rect 212460 557560 212552 557562
rect 212502 557504 212552 557560
rect 212460 557502 212552 557504
rect 212460 557500 212507 557502
rect 213494 557500 213500 557564
rect 213564 557562 213570 557564
rect 213821 557562 213887 557565
rect 213564 557560 213887 557562
rect 213564 557504 213826 557560
rect 213882 557504 213887 557560
rect 213564 557502 213887 557504
rect 213564 557500 213570 557502
rect 212441 557499 212507 557500
rect 213821 557499 213887 557502
rect 214782 557500 214788 557564
rect 214852 557562 214858 557564
rect 215201 557562 215267 557565
rect 214852 557560 215267 557562
rect 214852 557504 215206 557560
rect 215262 557504 215267 557560
rect 214852 557502 215267 557504
rect 214852 557500 214858 557502
rect 215201 557499 215267 557502
rect 216254 557500 216260 557564
rect 216324 557562 216330 557564
rect 216581 557562 216647 557565
rect 217869 557564 217935 557565
rect 217869 557562 217916 557564
rect 216324 557560 216647 557562
rect 216324 557504 216586 557560
rect 216642 557504 216647 557560
rect 216324 557502 216647 557504
rect 217824 557560 217916 557562
rect 217824 557504 217874 557560
rect 217824 557502 217916 557504
rect 216324 557500 216330 557502
rect 216581 557499 216647 557502
rect 217869 557500 217916 557502
rect 217980 557500 217986 557564
rect 219198 557500 219204 557564
rect 219268 557562 219274 557564
rect 219341 557562 219407 557565
rect 220721 557564 220787 557565
rect 219268 557560 219407 557562
rect 219268 557504 219346 557560
rect 219402 557504 219407 557560
rect 219268 557502 219407 557504
rect 219268 557500 219274 557502
rect 217869 557499 217935 557500
rect 219341 557499 219407 557502
rect 220670 557500 220676 557564
rect 220740 557562 220787 557564
rect 220740 557560 220832 557562
rect 220782 557504 220832 557560
rect 220740 557502 220832 557504
rect 220740 557500 220787 557502
rect 221958 557500 221964 557564
rect 222028 557562 222034 557564
rect 222101 557562 222167 557565
rect 222028 557560 222167 557562
rect 222028 557504 222106 557560
rect 222162 557504 222167 557560
rect 222028 557502 222167 557504
rect 222028 557500 222034 557502
rect 220721 557499 220787 557500
rect 222101 557499 222167 557502
rect 223246 557500 223252 557564
rect 223316 557562 223322 557564
rect 223481 557562 223547 557565
rect 223316 557560 223547 557562
rect 223316 557504 223486 557560
rect 223542 557504 223547 557560
rect 223316 557502 223547 557504
rect 223316 557500 223322 557502
rect 223481 557499 223547 557502
rect 224350 557500 224356 557564
rect 224420 557562 224426 557564
rect 224861 557562 224927 557565
rect 224420 557560 224927 557562
rect 224420 557504 224866 557560
rect 224922 557504 224927 557560
rect 224420 557502 224927 557504
rect 224420 557500 224426 557502
rect 224861 557499 224927 557502
rect 350625 557562 350691 557565
rect 350942 557562 350948 557564
rect 350625 557560 350948 557562
rect 350625 557504 350630 557560
rect 350686 557504 350948 557560
rect 350625 557502 350948 557504
rect 350625 557499 350691 557502
rect 350942 557500 350948 557502
rect 351012 557500 351018 557564
rect 353293 557562 353359 557565
rect 354438 557562 354444 557564
rect 353293 557560 354444 557562
rect 353293 557504 353298 557560
rect 353354 557504 354444 557560
rect 353293 557502 354444 557504
rect 353293 557499 353359 557502
rect 354438 557500 354444 557502
rect 354508 557500 354514 557564
rect 354673 557562 354739 557565
rect 355726 557562 355732 557564
rect 354673 557560 355732 557562
rect 354673 557504 354678 557560
rect 354734 557504 355732 557560
rect 354673 557502 355732 557504
rect 354673 557499 354739 557502
rect 355726 557500 355732 557502
rect 355796 557500 355802 557564
rect 356145 557562 356211 557565
rect 356646 557562 356652 557564
rect 356145 557560 356652 557562
rect 356145 557504 356150 557560
rect 356206 557504 356652 557560
rect 356145 557502 356652 557504
rect 356145 557499 356211 557502
rect 356646 557500 356652 557502
rect 356716 557500 356722 557564
rect 357525 557562 357591 557565
rect 357934 557562 357940 557564
rect 357525 557560 357940 557562
rect 357525 557504 357530 557560
rect 357586 557504 357940 557560
rect 357525 557502 357940 557504
rect 357525 557499 357591 557502
rect 357934 557500 357940 557502
rect 358004 557500 358010 557564
rect 583520 557140 584960 557380
rect 352005 555522 352071 555525
rect 352230 555522 352236 555524
rect 352005 555520 352236 555522
rect 352005 555464 352010 555520
rect 352066 555464 352236 555520
rect 352005 555462 352236 555464
rect 352005 555459 352071 555462
rect 352230 555460 352236 555462
rect 352300 555460 352306 555524
rect 358905 555522 358971 555525
rect 359222 555522 359228 555524
rect 358905 555520 359228 555522
rect 358905 555464 358910 555520
rect 358966 555464 359228 555520
rect 358905 555462 359228 555464
rect 358905 555459 358971 555462
rect 359222 555460 359228 555462
rect 359292 555460 359298 555524
rect -960 552924 480 553164
rect 583520 545444 584960 545684
rect 140037 543690 140103 543693
rect 200021 543690 200087 543693
rect 140037 543688 200087 543690
rect 140037 543632 140042 543688
rect 140098 543632 200026 543688
rect 200082 543632 200087 543688
rect 140037 543630 200087 543632
rect 140037 543627 140103 543630
rect 200021 543627 200087 543630
rect 148317 543554 148383 543557
rect 210417 543554 210483 543557
rect 148317 543552 210483 543554
rect 148317 543496 148322 543552
rect 148378 543496 210422 543552
rect 210478 543496 210483 543552
rect 148317 543494 210483 543496
rect 148317 543491 148383 543494
rect 210417 543491 210483 543494
rect 141417 543418 141483 543421
rect 208301 543418 208367 543421
rect 141417 543416 208367 543418
rect 141417 543360 141422 543416
rect 141478 543360 208306 543416
rect 208362 543360 208367 543416
rect 141417 543358 208367 543360
rect 141417 543355 141483 543358
rect 208301 543355 208367 543358
rect 96245 543282 96311 543285
rect 188337 543282 188403 543285
rect 96245 543280 188403 543282
rect 96245 543224 96250 543280
rect 96306 543224 188342 543280
rect 188398 543224 188403 543280
rect 96245 543222 188403 543224
rect 96245 543219 96311 543222
rect 188337 543219 188403 543222
rect 103421 543146 103487 543149
rect 202045 543146 202111 543149
rect 103421 543144 202111 543146
rect 103421 543088 103426 543144
rect 103482 543088 202050 543144
rect 202106 543088 202111 543144
rect 103421 543086 202111 543088
rect 103421 543083 103487 543086
rect 202045 543083 202111 543086
rect 77569 543010 77635 543013
rect 188981 543010 189047 543013
rect 77569 543008 189047 543010
rect 77569 542952 77574 543008
rect 77630 542952 188986 543008
rect 189042 542952 189047 543008
rect 77569 542950 189047 542952
rect 77569 542947 77635 542950
rect 188981 542947 189047 542950
rect 282269 539474 282335 539477
rect 279956 539472 282335 539474
rect 279956 539416 282274 539472
rect 282330 539416 282335 539472
rect 279956 539414 282335 539416
rect 282269 539411 282335 539414
rect -960 538508 480 538748
rect 282821 538522 282887 538525
rect 279956 538520 282887 538522
rect 279956 538464 282826 538520
rect 282882 538464 282887 538520
rect 279956 538462 282887 538464
rect 282821 538459 282887 538462
rect 282821 537434 282887 537437
rect 279956 537432 282887 537434
rect 279956 537376 282826 537432
rect 282882 537376 282887 537432
rect 279956 537374 282887 537376
rect 282821 537371 282887 537374
rect 282821 536482 282887 536485
rect 279956 536480 282887 536482
rect 279956 536424 282826 536480
rect 282882 536424 282887 536480
rect 279956 536422 282887 536424
rect 282821 536419 282887 536422
rect 281717 535394 281783 535397
rect 279956 535392 281783 535394
rect 279956 535336 281722 535392
rect 281778 535336 281783 535392
rect 279956 535334 281783 535336
rect 281717 535331 281783 535334
rect 282085 534442 282151 534445
rect 279956 534440 282151 534442
rect 279956 534384 282090 534440
rect 282146 534384 282151 534440
rect 279956 534382 282151 534384
rect 282085 534379 282151 534382
rect 583520 533748 584960 533988
rect 282085 533490 282151 533493
rect 279956 533488 282151 533490
rect 279956 533432 282090 533488
rect 282146 533432 282151 533488
rect 279956 533430 282151 533432
rect 282085 533427 282151 533430
rect 282269 532402 282335 532405
rect 279956 532400 282335 532402
rect 279956 532344 282274 532400
rect 282330 532344 282335 532400
rect 279956 532342 282335 532344
rect 282269 532339 282335 532342
rect 282821 531450 282887 531453
rect 279956 531448 282887 531450
rect 279956 531392 282826 531448
rect 282882 531392 282887 531448
rect 279956 531390 282887 531392
rect 282821 531387 282887 531390
rect 282821 530362 282887 530365
rect 279956 530360 282887 530362
rect 279956 530304 282826 530360
rect 282882 530304 282887 530360
rect 279956 530302 282887 530304
rect 282821 530299 282887 530302
rect 282821 529410 282887 529413
rect 279956 529408 282887 529410
rect 279956 529352 282826 529408
rect 282882 529352 282887 529408
rect 279956 529350 282887 529352
rect 282821 529347 282887 529350
rect 282269 528322 282335 528325
rect 279956 528320 282335 528322
rect 279956 528264 282274 528320
rect 282330 528264 282335 528320
rect 279956 528262 282335 528264
rect 282269 528259 282335 528262
rect 282821 527370 282887 527373
rect 279956 527368 282887 527370
rect 279956 527312 282826 527368
rect 282882 527312 282887 527368
rect 279956 527310 282887 527312
rect 282821 527307 282887 527310
rect 281901 526418 281967 526421
rect 279956 526416 281967 526418
rect 279956 526360 281906 526416
rect 281962 526360 281967 526416
rect 279956 526358 281967 526360
rect 281901 526355 281967 526358
rect 282821 525330 282887 525333
rect 279956 525328 282887 525330
rect 279956 525272 282826 525328
rect 282882 525272 282887 525328
rect 279956 525270 282887 525272
rect 282821 525267 282887 525270
rect 282361 524378 282427 524381
rect 279956 524376 282427 524378
rect -960 524092 480 524332
rect 279956 524320 282366 524376
rect 282422 524320 282427 524376
rect 279956 524318 282427 524320
rect 282361 524315 282427 524318
rect 282821 523290 282887 523293
rect 279956 523288 282887 523290
rect 279956 523232 282826 523288
rect 282882 523232 282887 523288
rect 279956 523230 282887 523232
rect 282821 523227 282887 523230
rect 282821 522338 282887 522341
rect 279956 522336 282887 522338
rect 279956 522280 282826 522336
rect 282882 522280 282887 522336
rect 279956 522278 282887 522280
rect 282821 522275 282887 522278
rect 583520 521916 584960 522156
rect 283557 521250 283623 521253
rect 279956 521248 283623 521250
rect 279956 521192 283562 521248
rect 283618 521192 283623 521248
rect 279956 521190 283623 521192
rect 283557 521187 283623 521190
rect 282821 520298 282887 520301
rect 279956 520296 282887 520298
rect 279956 520240 282826 520296
rect 282882 520240 282887 520296
rect 279956 520238 282887 520240
rect 282821 520235 282887 520238
rect 281717 519346 281783 519349
rect 279956 519344 281783 519346
rect 279956 519288 281722 519344
rect 281778 519288 281783 519344
rect 279956 519286 281783 519288
rect 281717 519283 281783 519286
rect 282085 518258 282151 518261
rect 279956 518256 282151 518258
rect 279956 518200 282090 518256
rect 282146 518200 282151 518256
rect 279956 518198 282151 518200
rect 282085 518195 282151 518198
rect 282269 517306 282335 517309
rect 279956 517304 282335 517306
rect 279956 517248 282274 517304
rect 282330 517248 282335 517304
rect 279956 517246 282335 517248
rect 282269 517243 282335 517246
rect 282821 516218 282887 516221
rect 279956 516216 282887 516218
rect 279956 516160 282826 516216
rect 282882 516160 282887 516216
rect 279956 516158 282887 516160
rect 282821 516155 282887 516158
rect 282821 515266 282887 515269
rect 279956 515264 282887 515266
rect 279956 515208 282826 515264
rect 282882 515208 282887 515264
rect 279956 515206 282887 515208
rect 282821 515203 282887 515206
rect 282269 514314 282335 514317
rect 279956 514312 282335 514314
rect 279956 514256 282274 514312
rect 282330 514256 282335 514312
rect 279956 514254 282335 514256
rect 282269 514251 282335 514254
rect 282729 513226 282795 513229
rect 279956 513224 282795 513226
rect 279956 513168 282734 513224
rect 282790 513168 282795 513224
rect 279956 513166 282795 513168
rect 282729 513163 282795 513166
rect 282821 512274 282887 512277
rect 279956 512272 282887 512274
rect 279956 512216 282826 512272
rect 282882 512216 282887 512272
rect 279956 512214 282887 512216
rect 282821 512211 282887 512214
rect 281717 511186 281783 511189
rect 279956 511184 281783 511186
rect 279956 511128 281722 511184
rect 281778 511128 281783 511184
rect 279956 511126 281783 511128
rect 281717 511123 281783 511126
rect 282269 510234 282335 510237
rect 279956 510232 282335 510234
rect 279956 510176 282274 510232
rect 282330 510176 282335 510232
rect 583520 510220 584960 510460
rect 279956 510174 282335 510176
rect 282269 510171 282335 510174
rect -960 509812 480 510052
rect 282545 509146 282611 509149
rect 279956 509144 282611 509146
rect 279956 509088 282550 509144
rect 282606 509088 282611 509144
rect 279956 509086 282611 509088
rect 282545 509083 282611 509086
rect 282821 508194 282887 508197
rect 279956 508192 282887 508194
rect 279956 508136 282826 508192
rect 282882 508136 282887 508192
rect 279956 508134 282887 508136
rect 282821 508131 282887 508134
rect 282085 507242 282151 507245
rect 279956 507240 282151 507242
rect 279956 507184 282090 507240
rect 282146 507184 282151 507240
rect 279956 507182 282151 507184
rect 282085 507179 282151 507182
rect 282729 506154 282795 506157
rect 279956 506152 282795 506154
rect 279956 506096 282734 506152
rect 282790 506096 282795 506152
rect 279956 506094 282795 506096
rect 282729 506091 282795 506094
rect 282821 505202 282887 505205
rect 279956 505200 282887 505202
rect 279956 505144 282826 505200
rect 282882 505144 282887 505200
rect 279956 505142 282887 505144
rect 282821 505139 282887 505142
rect 282821 504114 282887 504117
rect 279956 504112 282887 504114
rect 279956 504056 282826 504112
rect 282882 504056 282887 504112
rect 279956 504054 282887 504056
rect 282821 504051 282887 504054
rect 282821 503162 282887 503165
rect 279956 503160 282887 503162
rect 279956 503104 282826 503160
rect 282882 503104 282887 503160
rect 279956 503102 282887 503104
rect 282821 503099 282887 503102
rect 282269 502074 282335 502077
rect 279956 502072 282335 502074
rect 279956 502016 282274 502072
rect 282330 502016 282335 502072
rect 279956 502014 282335 502016
rect 282269 502011 282335 502014
rect 282821 501122 282887 501125
rect 279956 501120 282887 501122
rect 279956 501064 282826 501120
rect 282882 501064 282887 501120
rect 279956 501062 282887 501064
rect 282821 501059 282887 501062
rect 282821 499082 282887 499085
rect 279956 499080 282887 499082
rect 279956 499024 282826 499080
rect 282882 499024 282887 499080
rect 279956 499022 282887 499024
rect 282821 499019 282887 499022
rect 583520 498524 584960 498764
rect 282821 497042 282887 497045
rect 279956 497040 282887 497042
rect 279956 496984 282826 497040
rect 282882 496984 282887 497040
rect 279956 496982 282887 496984
rect 282821 496979 282887 496982
rect 281901 496090 281967 496093
rect 279956 496088 281967 496090
rect 279956 496032 281906 496088
rect 281962 496032 281967 496088
rect 279956 496030 281967 496032
rect 281901 496027 281967 496030
rect -960 495396 480 495636
rect 282821 495138 282887 495141
rect 279956 495136 282887 495138
rect 279956 495080 282826 495136
rect 282882 495080 282887 495136
rect 279956 495078 282887 495080
rect 282821 495075 282887 495078
rect 282361 494050 282427 494053
rect 279956 494048 282427 494050
rect 279956 493992 282366 494048
rect 282422 493992 282427 494048
rect 279956 493990 282427 493992
rect 282361 493987 282427 493990
rect 282821 493098 282887 493101
rect 279956 493096 282887 493098
rect 279956 493040 282826 493096
rect 282882 493040 282887 493096
rect 279956 493038 282887 493040
rect 282821 493035 282887 493038
rect 282821 492010 282887 492013
rect 279956 492008 282887 492010
rect 279956 491952 282826 492008
rect 282882 491952 282887 492008
rect 279956 491950 282887 491952
rect 282821 491947 282887 491950
rect 282269 491058 282335 491061
rect 279956 491056 282335 491058
rect 279956 491000 282274 491056
rect 282330 491000 282335 491056
rect 279956 490998 282335 491000
rect 282269 490995 282335 490998
rect 282821 489970 282887 489973
rect 279956 489968 282887 489970
rect 279956 489912 282826 489968
rect 282882 489912 282887 489968
rect 279956 489910 282887 489912
rect 282821 489907 282887 489910
rect 282269 489018 282335 489021
rect 279956 489016 282335 489018
rect 279956 488960 282274 489016
rect 282330 488960 282335 489016
rect 279956 488958 282335 488960
rect 282269 488955 282335 488958
rect 282821 488066 282887 488069
rect 279956 488064 282887 488066
rect 279956 488008 282826 488064
rect 282882 488008 282887 488064
rect 279956 488006 282887 488008
rect 282821 488003 282887 488006
rect 282269 486978 282335 486981
rect 279956 486976 282335 486978
rect 279956 486920 282274 486976
rect 282330 486920 282335 486976
rect 279956 486918 282335 486920
rect 282269 486915 282335 486918
rect 583520 486692 584960 486932
rect 282821 486026 282887 486029
rect 279956 486024 282887 486026
rect 279956 485968 282826 486024
rect 282882 485968 282887 486024
rect 279956 485966 282887 485968
rect 282821 485963 282887 485966
rect 281717 484938 281783 484941
rect 279956 484936 281783 484938
rect 279956 484880 281722 484936
rect 281778 484880 281783 484936
rect 279956 484878 281783 484880
rect 281717 484875 281783 484878
rect 282269 483986 282335 483989
rect 279956 483984 282335 483986
rect 279956 483928 282274 483984
rect 282330 483928 282335 483984
rect 279956 483926 282335 483928
rect 282269 483923 282335 483926
rect 282545 482898 282611 482901
rect 279956 482896 282611 482898
rect 279956 482840 282550 482896
rect 282606 482840 282611 482896
rect 279956 482838 282611 482840
rect 282545 482835 282611 482838
rect 282821 481946 282887 481949
rect 279956 481944 282887 481946
rect 279956 481888 282826 481944
rect 282882 481888 282887 481944
rect 279956 481886 282887 481888
rect 282821 481883 282887 481886
rect -960 480980 480 481220
rect 282085 480994 282151 480997
rect 279956 480992 282151 480994
rect 279956 480936 282090 480992
rect 282146 480936 282151 480992
rect 279956 480934 282151 480936
rect 282085 480931 282151 480934
rect 282729 479906 282795 479909
rect 279956 479904 282795 479906
rect 279956 479848 282734 479904
rect 282790 479848 282795 479904
rect 279956 479846 282795 479848
rect 282729 479843 282795 479846
rect 282821 478954 282887 478957
rect 279956 478952 282887 478954
rect 279956 478896 282826 478952
rect 282882 478896 282887 478952
rect 279956 478894 282887 478896
rect 282821 478891 282887 478894
rect 282821 477866 282887 477869
rect 279956 477864 282887 477866
rect 279956 477808 282826 477864
rect 282882 477808 282887 477864
rect 279956 477806 282887 477808
rect 282821 477803 282887 477806
rect 282085 476914 282151 476917
rect 279956 476912 282151 476914
rect 279956 476856 282090 476912
rect 282146 476856 282151 476912
rect 279956 476854 282151 476856
rect 282085 476851 282151 476854
rect 282269 475826 282335 475829
rect 279956 475824 282335 475826
rect 279956 475768 282274 475824
rect 282330 475768 282335 475824
rect 279956 475766 282335 475768
rect 282269 475763 282335 475766
rect 583520 474996 584960 475236
rect 282821 474874 282887 474877
rect 279956 474872 282887 474874
rect 279956 474816 282826 474872
rect 282882 474816 282887 474872
rect 279956 474814 282887 474816
rect 282821 474811 282887 474814
rect 281717 473922 281783 473925
rect 279956 473920 281783 473922
rect 279956 473864 281722 473920
rect 281778 473864 281783 473920
rect 279956 473862 281783 473864
rect 281717 473859 281783 473862
rect 282085 472834 282151 472837
rect 279956 472832 282151 472834
rect 279956 472776 282090 472832
rect 282146 472776 282151 472832
rect 279956 472774 282151 472776
rect 282085 472771 282151 472774
rect 282729 471882 282795 471885
rect 279956 471880 282795 471882
rect 279956 471824 282734 471880
rect 282790 471824 282795 471880
rect 279956 471822 282795 471824
rect 282729 471819 282795 471822
rect 282821 470794 282887 470797
rect 279956 470792 282887 470794
rect 279956 470736 282826 470792
rect 282882 470736 282887 470792
rect 279956 470734 282887 470736
rect 282821 470731 282887 470734
rect 281901 469842 281967 469845
rect 279956 469840 281967 469842
rect 279956 469784 281906 469840
rect 281962 469784 281967 469840
rect 279956 469782 281967 469784
rect 281901 469779 281967 469782
rect 282821 468890 282887 468893
rect 279956 468888 282887 468890
rect 279956 468832 282826 468888
rect 282882 468832 282887 468888
rect 279956 468830 282887 468832
rect 282821 468827 282887 468830
rect 282729 467802 282795 467805
rect 279956 467800 282795 467802
rect 279956 467744 282734 467800
rect 282790 467744 282795 467800
rect 279956 467742 282795 467744
rect 282729 467739 282795 467742
rect -960 466700 480 466940
rect 282821 466850 282887 466853
rect 279956 466848 282887 466850
rect 279956 466792 282826 466848
rect 282882 466792 282887 466848
rect 279956 466790 282887 466792
rect 282821 466787 282887 466790
rect 282821 465762 282887 465765
rect 279956 465760 282887 465762
rect 279956 465704 282826 465760
rect 282882 465704 282887 465760
rect 279956 465702 282887 465704
rect 282821 465699 282887 465702
rect 282729 464810 282795 464813
rect 279956 464808 282795 464810
rect 279956 464752 282734 464808
rect 282790 464752 282795 464808
rect 279956 464750 282795 464752
rect 282729 464747 282795 464750
rect 282821 463722 282887 463725
rect 279956 463720 282887 463722
rect 279956 463664 282826 463720
rect 282882 463664 282887 463720
rect 279956 463662 282887 463664
rect 282821 463659 282887 463662
rect 583520 463300 584960 463540
rect 282821 462770 282887 462773
rect 279956 462768 282887 462770
rect 279956 462712 282826 462768
rect 282882 462712 282887 462768
rect 279956 462710 282887 462712
rect 282821 462707 282887 462710
rect 282821 461818 282887 461821
rect 279956 461816 282887 461818
rect 279956 461760 282826 461816
rect 282882 461760 282887 461816
rect 279956 461758 282887 461760
rect 282821 461755 282887 461758
rect 282821 460730 282887 460733
rect 279956 460728 282887 460730
rect 279956 460672 282826 460728
rect 282882 460672 282887 460728
rect 279956 460670 282887 460672
rect 282821 460667 282887 460670
rect 282729 459778 282795 459781
rect 279956 459776 282795 459778
rect 279956 459720 282734 459776
rect 282790 459720 282795 459776
rect 279956 459718 282795 459720
rect 282729 459715 282795 459718
rect 281717 458690 281783 458693
rect 279956 458688 281783 458690
rect 279956 458632 281722 458688
rect 281778 458632 281783 458688
rect 279956 458630 281783 458632
rect 281717 458627 281783 458630
rect 282085 457738 282151 457741
rect 279956 457736 282151 457738
rect 279956 457680 282090 457736
rect 282146 457680 282151 457736
rect 279956 457678 282151 457680
rect 282085 457675 282151 457678
rect 281625 456650 281691 456653
rect 279956 456648 281691 456650
rect 279956 456592 281630 456648
rect 281686 456592 281691 456648
rect 279956 456590 281691 456592
rect 281625 456587 281691 456590
rect 282821 455698 282887 455701
rect 279956 455696 282887 455698
rect 279956 455640 282826 455696
rect 282882 455640 282887 455696
rect 279956 455638 282887 455640
rect 282821 455635 282887 455638
rect 281625 454746 281691 454749
rect 279956 454744 281691 454746
rect 279956 454688 281630 454744
rect 281686 454688 281691 454744
rect 279956 454686 281691 454688
rect 281625 454683 281691 454686
rect 282453 453658 282519 453661
rect 279956 453656 282519 453658
rect 279956 453600 282458 453656
rect 282514 453600 282519 453656
rect 279956 453598 282519 453600
rect 282453 453595 282519 453598
rect 282269 452706 282335 452709
rect 279956 452704 282335 452706
rect 279956 452648 282274 452704
rect 282330 452648 282335 452704
rect 279956 452646 282335 452648
rect 282269 452643 282335 452646
rect -960 452284 480 452524
rect 282361 451618 282427 451621
rect 279956 451616 282427 451618
rect 279956 451560 282366 451616
rect 282422 451560 282427 451616
rect 583520 451604 584960 451844
rect 279956 451558 282427 451560
rect 282361 451555 282427 451558
rect 282545 450666 282611 450669
rect 279956 450664 282611 450666
rect 279956 450608 282550 450664
rect 282606 450608 282611 450664
rect 279956 450606 282611 450608
rect 282545 450603 282611 450606
rect 282821 449714 282887 449717
rect 279956 449712 282887 449714
rect 279956 449656 282826 449712
rect 282882 449656 282887 449712
rect 279956 449654 282887 449656
rect 282821 449651 282887 449654
rect 282637 448626 282703 448629
rect 279956 448624 282703 448626
rect 279956 448568 282642 448624
rect 282698 448568 282703 448624
rect 279956 448566 282703 448568
rect 282637 448563 282703 448566
rect 282729 447674 282795 447677
rect 279956 447672 282795 447674
rect 279956 447616 282734 447672
rect 282790 447616 282795 447672
rect 279956 447614 282795 447616
rect 282729 447611 282795 447614
rect 282085 446586 282151 446589
rect 279956 446584 282151 446586
rect 279956 446528 282090 446584
rect 282146 446528 282151 446584
rect 279956 446526 282151 446528
rect 282085 446523 282151 446526
rect 281809 445634 281875 445637
rect 279956 445632 281875 445634
rect 279956 445576 281814 445632
rect 281870 445576 281875 445632
rect 279956 445574 281875 445576
rect 281809 445571 281875 445574
rect 281993 444546 282059 444549
rect 279956 444544 282059 444546
rect 279956 444488 281998 444544
rect 282054 444488 282059 444544
rect 279956 444486 282059 444488
rect 281993 444483 282059 444486
rect 281901 443594 281967 443597
rect 279956 443592 281967 443594
rect 279956 443536 281906 443592
rect 281962 443536 281967 443592
rect 279956 443534 281967 443536
rect 281901 443531 281967 443534
rect 281717 442642 281783 442645
rect 279956 442640 281783 442642
rect 279956 442584 281722 442640
rect 281778 442584 281783 442640
rect 279956 442582 281783 442584
rect 281717 442579 281783 442582
rect 279926 441010 279986 441524
rect 281441 441010 281507 441013
rect 279926 441008 281507 441010
rect 279926 440952 281446 441008
rect 281502 440952 281507 441008
rect 279926 440950 281507 440952
rect 281441 440947 281507 440950
rect 282177 440602 282243 440605
rect 279956 440600 282243 440602
rect 279956 440544 282182 440600
rect 282238 440544 282243 440600
rect 279956 440542 282243 440544
rect 282177 440539 282243 440542
rect 583520 439772 584960 440012
rect 282177 439514 282243 439517
rect 279956 439512 282243 439514
rect 279956 439456 282182 439512
rect 282238 439456 282243 439512
rect 279956 439454 282243 439456
rect 282177 439451 282243 439454
rect 283465 438562 283531 438565
rect 279956 438560 283531 438562
rect 279956 438504 283470 438560
rect 283526 438504 283531 438560
rect 279956 438502 283531 438504
rect 283465 438499 283531 438502
rect -960 437868 480 438108
rect 282177 437474 282243 437477
rect 279956 437472 282243 437474
rect 279956 437416 282182 437472
rect 282238 437416 282243 437472
rect 279956 437414 282243 437416
rect 282177 437411 282243 437414
rect 282177 436522 282243 436525
rect 279956 436520 282243 436522
rect 279956 436464 282182 436520
rect 282238 436464 282243 436520
rect 279956 436462 282243 436464
rect 282177 436459 282243 436462
rect 282177 435570 282243 435573
rect 279956 435568 282243 435570
rect 279956 435512 282182 435568
rect 282238 435512 282243 435568
rect 279956 435510 282243 435512
rect 282177 435507 282243 435510
rect 282177 434482 282243 434485
rect 279956 434480 282243 434482
rect 279956 434424 282182 434480
rect 282238 434424 282243 434480
rect 279956 434422 282243 434424
rect 282177 434419 282243 434422
rect 283373 433530 283439 433533
rect 279956 433528 283439 433530
rect 279956 433472 283378 433528
rect 283434 433472 283439 433528
rect 279956 433470 283439 433472
rect 283373 433467 283439 433470
rect 282177 432442 282243 432445
rect 279956 432440 282243 432442
rect 279956 432384 282182 432440
rect 282238 432384 282243 432440
rect 279956 432382 282243 432384
rect 282177 432379 282243 432382
rect 282269 431490 282335 431493
rect 279956 431488 282335 431490
rect 279956 431432 282274 431488
rect 282330 431432 282335 431488
rect 279956 431430 282335 431432
rect 282269 431427 282335 431430
rect 279926 429994 279986 430508
rect 281441 429994 281507 429997
rect 279926 429992 281507 429994
rect 279926 429936 281446 429992
rect 281502 429936 281507 429992
rect 279926 429934 281507 429936
rect 281441 429931 281507 429934
rect 282269 429450 282335 429453
rect 279956 429448 282335 429450
rect 279956 429392 282274 429448
rect 282330 429392 282335 429448
rect 279956 429390 282335 429392
rect 282269 429387 282335 429390
rect 282269 428498 282335 428501
rect 279956 428496 282335 428498
rect 279956 428440 282274 428496
rect 282330 428440 282335 428496
rect 279956 428438 282335 428440
rect 282269 428435 282335 428438
rect 583520 428076 584960 428316
rect 282269 427410 282335 427413
rect 279956 427408 282335 427410
rect 279956 427352 282274 427408
rect 282330 427352 282335 427408
rect 279956 427350 282335 427352
rect 282269 427347 282335 427350
rect 282269 427002 282335 427005
rect 279926 427000 282335 427002
rect 279926 426944 282274 427000
rect 282330 426944 282335 427000
rect 279926 426942 282335 426944
rect 279926 426428 279986 426942
rect 282269 426939 282335 426942
rect 282269 425370 282335 425373
rect 279956 425368 282335 425370
rect 279956 425312 282274 425368
rect 282330 425312 282335 425368
rect 279956 425310 282335 425312
rect 282269 425307 282335 425310
rect 282269 424418 282335 424421
rect 279956 424416 282335 424418
rect 279956 424360 282274 424416
rect 282330 424360 282335 424416
rect 279956 424358 282335 424360
rect 282269 424355 282335 424358
rect -960 423588 480 423828
rect 282269 423466 282335 423469
rect 279956 423464 282335 423466
rect 279956 423408 282274 423464
rect 282330 423408 282335 423464
rect 279956 423406 282335 423408
rect 282269 423403 282335 423406
rect 282269 422378 282335 422381
rect 279956 422376 282335 422378
rect 279956 422320 282274 422376
rect 282330 422320 282335 422376
rect 279956 422318 282335 422320
rect 282269 422315 282335 422318
rect 282269 421426 282335 421429
rect 279956 421424 282335 421426
rect 279956 421368 282274 421424
rect 282330 421368 282335 421424
rect 279956 421366 282335 421368
rect 282269 421363 282335 421366
rect 282821 420338 282887 420341
rect 279956 420336 282887 420338
rect 279956 420280 282826 420336
rect 282882 420280 282887 420336
rect 279956 420278 282887 420280
rect 282821 420275 282887 420278
rect 282821 419386 282887 419389
rect 279956 419384 282887 419386
rect 279956 419328 282826 419384
rect 282882 419328 282887 419384
rect 279956 419326 282887 419328
rect 282821 419323 282887 419326
rect 282545 418298 282611 418301
rect 279956 418296 282611 418298
rect 279956 418240 282550 418296
rect 282606 418240 282611 418296
rect 279956 418238 282611 418240
rect 282545 418235 282611 418238
rect 282821 417346 282887 417349
rect 279956 417344 282887 417346
rect 279956 417288 282826 417344
rect 282882 417288 282887 417344
rect 279956 417286 282887 417288
rect 282821 417283 282887 417286
rect 282821 416394 282887 416397
rect 279956 416392 282887 416394
rect 279956 416336 282826 416392
rect 282882 416336 282887 416392
rect 583520 416380 584960 416620
rect 279956 416334 282887 416336
rect 282821 416331 282887 416334
rect 282821 415306 282887 415309
rect 279956 415304 282887 415306
rect 279956 415248 282826 415304
rect 282882 415248 282887 415304
rect 279956 415246 282887 415248
rect 282821 415243 282887 415246
rect 282269 414354 282335 414357
rect 279956 414352 282335 414354
rect 279956 414296 282274 414352
rect 282330 414296 282335 414352
rect 279956 414294 282335 414296
rect 282269 414291 282335 414294
rect 371877 414082 371943 414085
rect 371877 414080 373274 414082
rect 371877 414024 371882 414080
rect 371938 414024 373274 414080
rect 371877 414022 373274 414024
rect 371877 414019 371943 414022
rect 367093 413946 367159 413949
rect 368238 413946 368244 413948
rect 367093 413944 368244 413946
rect 367093 413888 367098 413944
rect 367154 413888 368244 413944
rect 367093 413886 368244 413888
rect 367093 413883 367159 413886
rect 368238 413884 368244 413886
rect 368308 413884 368314 413948
rect 368565 413946 368631 413949
rect 368974 413946 368980 413948
rect 368565 413944 368980 413946
rect 368565 413888 368570 413944
rect 368626 413888 368980 413944
rect 368565 413886 368980 413888
rect 368565 413883 368631 413886
rect 368974 413884 368980 413886
rect 369044 413884 369050 413948
rect 369945 413946 370011 413949
rect 370262 413946 370268 413948
rect 369945 413944 370268 413946
rect 369945 413888 369950 413944
rect 370006 413888 370268 413944
rect 369945 413886 370268 413888
rect 369945 413883 370011 413886
rect 370262 413884 370268 413886
rect 370332 413884 370338 413948
rect 371233 413946 371299 413949
rect 371918 413946 371924 413948
rect 371233 413944 371924 413946
rect 371233 413888 371238 413944
rect 371294 413888 371924 413944
rect 371233 413886 371924 413888
rect 371233 413883 371299 413886
rect 371918 413884 371924 413886
rect 371988 413884 371994 413948
rect 372613 413946 372679 413949
rect 373022 413946 373028 413948
rect 372613 413944 373028 413946
rect 372613 413888 372618 413944
rect 372674 413888 373028 413944
rect 372613 413886 373028 413888
rect 372613 413883 372679 413886
rect 373022 413884 373028 413886
rect 373092 413884 373098 413948
rect 373214 413946 373274 414022
rect 379470 414022 380450 414082
rect 379470 413946 379530 414022
rect 373214 413886 379530 413946
rect 379605 413946 379671 413949
rect 380198 413946 380204 413948
rect 379605 413944 380204 413946
rect 379605 413888 379610 413944
rect 379666 413888 380204 413944
rect 379605 413886 380204 413888
rect 379605 413883 379671 413886
rect 380198 413884 380204 413886
rect 380268 413884 380274 413948
rect 380390 413946 380450 414022
rect 384614 413946 384620 413948
rect 380390 413886 380818 413946
rect 354121 413810 354187 413813
rect 380617 413810 380683 413813
rect 354121 413808 380683 413810
rect 354121 413752 354126 413808
rect 354182 413752 380622 413808
rect 380678 413752 380683 413808
rect 354121 413750 380683 413752
rect 380758 413810 380818 413886
rect 381494 413886 384620 413946
rect 381494 413810 381554 413886
rect 384614 413884 384620 413886
rect 384684 413884 384690 413948
rect 387885 413946 387951 413949
rect 390645 413948 390711 413949
rect 388294 413946 388300 413948
rect 387885 413944 388300 413946
rect 387885 413888 387890 413944
rect 387946 413888 388300 413944
rect 387885 413886 388300 413888
rect 387885 413883 387951 413886
rect 388294 413884 388300 413886
rect 388364 413884 388370 413948
rect 390645 413946 390692 413948
rect 390600 413944 390692 413946
rect 390600 413888 390650 413944
rect 390600 413886 390692 413888
rect 390645 413884 390692 413886
rect 390756 413884 390762 413948
rect 392025 413946 392091 413949
rect 402973 413948 403039 413949
rect 407757 413948 407823 413949
rect 410517 413948 410583 413949
rect 413921 413948 413987 413949
rect 392894 413946 392900 413948
rect 392025 413944 392900 413946
rect 392025 413888 392030 413944
rect 392086 413888 392900 413944
rect 392025 413886 392900 413888
rect 390645 413883 390711 413884
rect 392025 413883 392091 413886
rect 392894 413884 392900 413886
rect 392964 413884 392970 413948
rect 397862 413946 397868 413948
rect 393086 413886 397868 413946
rect 380758 413750 381554 413810
rect 384297 413810 384363 413813
rect 391933 413810 391999 413813
rect 392158 413810 392164 413812
rect 384297 413808 389650 413810
rect 384297 413752 384302 413808
rect 384358 413752 389650 413808
rect 384297 413750 389650 413752
rect 354121 413747 354187 413750
rect 380617 413747 380683 413750
rect 384297 413747 384363 413750
rect 283557 413674 283623 413677
rect 389398 413674 389404 413676
rect 283557 413672 389404 413674
rect 283557 413616 283562 413672
rect 283618 413616 389404 413672
rect 283557 413614 389404 413616
rect 283557 413611 283623 413614
rect 389398 413612 389404 413614
rect 389468 413612 389474 413676
rect 389590 413674 389650 413750
rect 391933 413808 392164 413810
rect 391933 413752 391938 413808
rect 391994 413752 392164 413808
rect 391933 413750 392164 413752
rect 391933 413747 391999 413750
rect 392158 413748 392164 413750
rect 392228 413748 392234 413812
rect 393086 413674 393146 413886
rect 397862 413884 397868 413886
rect 397932 413884 397938 413948
rect 402973 413944 403020 413948
rect 403084 413946 403090 413948
rect 407757 413946 407804 413948
rect 402973 413888 402978 413944
rect 402973 413884 403020 413888
rect 403084 413886 403130 413946
rect 407712 413944 407804 413946
rect 407712 413888 407762 413944
rect 407712 413886 407804 413888
rect 403084 413884 403090 413886
rect 407757 413884 407804 413886
rect 407868 413884 407874 413948
rect 410517 413944 410564 413948
rect 410628 413946 410634 413948
rect 413870 413946 413876 413948
rect 410517 413888 410522 413944
rect 410517 413884 410564 413888
rect 410628 413886 410674 413946
rect 413830 413886 413876 413946
rect 413940 413944 413987 413948
rect 413982 413888 413987 413944
rect 410628 413884 410634 413886
rect 413870 413884 413876 413886
rect 413940 413884 413987 413888
rect 402973 413883 403039 413884
rect 407757 413883 407823 413884
rect 410517 413883 410583 413884
rect 413921 413883 413987 413884
rect 470685 413946 470751 413949
rect 474825 413948 474891 413949
rect 470910 413946 470916 413948
rect 470685 413944 470916 413946
rect 470685 413888 470690 413944
rect 470746 413888 470916 413944
rect 470685 413886 470916 413888
rect 470685 413883 470751 413886
rect 470910 413884 470916 413886
rect 470980 413884 470986 413948
rect 474774 413946 474780 413948
rect 474734 413886 474780 413946
rect 474844 413944 474891 413948
rect 474886 413888 474891 413944
rect 474774 413884 474780 413886
rect 474844 413884 474891 413888
rect 474825 413883 474891 413884
rect 477585 413946 477651 413949
rect 478270 413946 478276 413948
rect 477585 413944 478276 413946
rect 477585 413888 477590 413944
rect 477646 413888 478276 413944
rect 477585 413886 478276 413888
rect 477585 413883 477651 413886
rect 478270 413884 478276 413886
rect 478340 413884 478346 413948
rect 396073 413812 396139 413813
rect 396022 413748 396028 413812
rect 396092 413810 396139 413812
rect 476113 413810 476179 413813
rect 477493 413812 477559 413813
rect 476246 413810 476252 413812
rect 396092 413808 396184 413810
rect 396134 413752 396184 413808
rect 396092 413750 396184 413752
rect 476113 413808 476252 413810
rect 476113 413752 476118 413808
rect 476174 413752 476252 413808
rect 476113 413750 476252 413752
rect 396092 413748 396139 413750
rect 396073 413747 396139 413748
rect 476113 413747 476179 413750
rect 476246 413748 476252 413750
rect 476316 413748 476322 413812
rect 477493 413810 477540 413812
rect 477448 413808 477540 413810
rect 477448 413752 477498 413808
rect 477448 413750 477540 413752
rect 477493 413748 477540 413750
rect 477604 413748 477610 413812
rect 505093 413810 505159 413813
rect 505686 413810 505692 413812
rect 505093 413808 505692 413810
rect 505093 413752 505098 413808
rect 505154 413752 505692 413808
rect 505093 413750 505692 413752
rect 477493 413747 477559 413748
rect 505093 413747 505159 413750
rect 505686 413748 505692 413750
rect 505756 413748 505762 413812
rect 389590 413614 393146 413674
rect 478873 413674 478939 413677
rect 479374 413674 479380 413676
rect 478873 413672 479380 413674
rect 478873 413616 478878 413672
rect 478934 413616 479380 413672
rect 478873 413614 479380 413616
rect 478873 413611 478939 413614
rect 479374 413612 479380 413614
rect 479444 413612 479450 413676
rect 506473 413674 506539 413677
rect 506974 413674 506980 413676
rect 506473 413672 506980 413674
rect 506473 413616 506478 413672
rect 506534 413616 506980 413672
rect 506473 413614 506980 413616
rect 506473 413611 506539 413614
rect 506974 413612 506980 413614
rect 507044 413612 507050 413676
rect 283741 413538 283807 413541
rect 385309 413538 385375 413541
rect 386413 413540 386479 413541
rect 389173 413540 389239 413541
rect 386413 413538 386460 413540
rect 283741 413536 385375 413538
rect 283741 413480 283746 413536
rect 283802 413480 385314 413536
rect 385370 413480 385375 413536
rect 283741 413478 385375 413480
rect 386368 413536 386460 413538
rect 386368 413480 386418 413536
rect 386368 413478 386460 413480
rect 283741 413475 283807 413478
rect 385309 413475 385375 413478
rect 386413 413476 386460 413478
rect 386524 413476 386530 413540
rect 389173 413538 389220 413540
rect 389128 413536 389220 413538
rect 389128 413480 389178 413536
rect 389128 413478 389220 413480
rect 389173 413476 389220 413478
rect 389284 413476 389290 413540
rect 389357 413538 389423 413541
rect 394693 413540 394759 413541
rect 404353 413540 404419 413541
rect 394693 413538 394740 413540
rect 389357 413536 393146 413538
rect 389357 413480 389362 413536
rect 389418 413480 393146 413536
rect 389357 413478 393146 413480
rect 394648 413536 394740 413538
rect 394648 413480 394698 413536
rect 394648 413478 394740 413480
rect 386413 413475 386479 413476
rect 389173 413475 389239 413476
rect 389357 413475 389423 413478
rect 283373 413402 283439 413405
rect 287053 413402 287119 413405
rect 283373 413400 287119 413402
rect 283373 413344 283378 413400
rect 283434 413344 287058 413400
rect 287114 413344 287119 413400
rect 283373 413342 287119 413344
rect 283373 413339 283439 413342
rect 287053 413339 287119 413342
rect 296621 413402 296687 413405
rect 306373 413402 306439 413405
rect 296621 413400 306439 413402
rect 296621 413344 296626 413400
rect 296682 413344 306378 413400
rect 306434 413344 306439 413400
rect 296621 413342 306439 413344
rect 296621 413339 296687 413342
rect 306373 413339 306439 413342
rect 315941 413402 316007 413405
rect 335261 413402 335327 413405
rect 354581 413402 354647 413405
rect 364333 413402 364399 413405
rect 315941 413400 321018 413402
rect 315941 413344 315946 413400
rect 316002 413344 321018 413400
rect 315941 413342 321018 413344
rect 315941 413339 316007 413342
rect 282821 413266 282887 413269
rect 279956 413264 282887 413266
rect 279956 413208 282826 413264
rect 282882 413208 282887 413264
rect 279956 413206 282887 413208
rect 282821 413203 282887 413206
rect 283925 413266 283991 413269
rect 287145 413266 287211 413269
rect 283925 413264 287211 413266
rect 283925 413208 283930 413264
rect 283986 413208 287150 413264
rect 287206 413208 287211 413264
rect 283925 413206 287211 413208
rect 283925 413203 283991 413206
rect 287145 413203 287211 413206
rect 296529 413266 296595 413269
rect 306465 413266 306531 413269
rect 296529 413264 306531 413266
rect 296529 413208 296534 413264
rect 296590 413208 306470 413264
rect 306526 413208 306531 413264
rect 296529 413206 306531 413208
rect 296529 413203 296595 413206
rect 306465 413203 306531 413206
rect 315849 413266 315915 413269
rect 315849 413264 320650 413266
rect 315849 413208 315854 413264
rect 315910 413208 320650 413264
rect 315849 413206 320650 413208
rect 315849 413203 315915 413206
rect 287053 413130 287119 413133
rect 296621 413130 296687 413133
rect 287053 413128 296687 413130
rect 287053 413072 287058 413128
rect 287114 413072 296626 413128
rect 296682 413072 296687 413128
rect 287053 413070 296687 413072
rect 287053 413067 287119 413070
rect 296621 413067 296687 413070
rect 306373 413130 306439 413133
rect 315941 413130 316007 413133
rect 306373 413128 316007 413130
rect 306373 413072 306378 413128
rect 306434 413072 315946 413128
rect 316002 413072 316007 413128
rect 306373 413070 316007 413072
rect 306373 413067 306439 413070
rect 315941 413067 316007 413070
rect 287053 412994 287119 412997
rect 296621 412994 296687 412997
rect 287053 412992 296687 412994
rect 287053 412936 287058 412992
rect 287114 412936 296626 412992
rect 296682 412936 296687 412992
rect 287053 412934 296687 412936
rect 287053 412931 287119 412934
rect 296621 412931 296687 412934
rect 306373 412994 306439 412997
rect 315941 412994 316007 412997
rect 306373 412992 316007 412994
rect 306373 412936 306378 412992
rect 306434 412936 315946 412992
rect 316002 412936 316007 412992
rect 306373 412934 316007 412936
rect 306373 412931 306439 412934
rect 315941 412931 316007 412934
rect 287145 412858 287211 412861
rect 296529 412858 296595 412861
rect 287145 412856 296595 412858
rect 287145 412800 287150 412856
rect 287206 412800 296534 412856
rect 296590 412800 296595 412856
rect 287145 412798 296595 412800
rect 287145 412795 287211 412798
rect 296529 412795 296595 412798
rect 306465 412858 306531 412861
rect 315849 412858 315915 412861
rect 306465 412856 315915 412858
rect 306465 412800 306470 412856
rect 306526 412800 315854 412856
rect 315910 412800 315915 412856
rect 306465 412798 315915 412800
rect 320590 412858 320650 413206
rect 320958 413130 321018 413342
rect 335261 413400 340522 413402
rect 335261 413344 335266 413400
rect 335322 413344 340522 413400
rect 335261 413342 340522 413344
rect 335261 413339 335327 413342
rect 335169 413266 335235 413269
rect 335169 413264 340154 413266
rect 335169 413208 335174 413264
rect 335230 413208 340154 413264
rect 335169 413206 340154 413208
rect 335169 413203 335235 413206
rect 335261 413130 335327 413133
rect 320958 413128 335327 413130
rect 320958 413072 335266 413128
rect 335322 413072 335327 413128
rect 320958 413070 335327 413072
rect 335261 413067 335327 413070
rect 331121 412994 331187 412997
rect 335261 412994 335327 412997
rect 331121 412992 335327 412994
rect 331121 412936 331126 412992
rect 331182 412936 335266 412992
rect 335322 412936 335327 412992
rect 331121 412934 335327 412936
rect 340094 412994 340154 413206
rect 340462 413130 340522 413342
rect 354581 413400 364399 413402
rect 354581 413344 354586 413400
rect 354642 413344 364338 413400
rect 364394 413344 364399 413400
rect 354581 413342 364399 413344
rect 354581 413339 354647 413342
rect 364333 413339 364399 413342
rect 373901 413402 373967 413405
rect 379789 413402 379855 413405
rect 373901 413400 379855 413402
rect 373901 413344 373906 413400
rect 373962 413344 379794 413400
rect 379850 413344 379855 413400
rect 373901 413342 379855 413344
rect 373901 413339 373967 413342
rect 379789 413339 379855 413342
rect 380985 413402 381051 413405
rect 381486 413402 381492 413404
rect 380985 413400 381492 413402
rect 380985 413344 380990 413400
rect 381046 413344 381492 413400
rect 380985 413342 381492 413344
rect 380985 413339 381051 413342
rect 381486 413340 381492 413342
rect 381556 413340 381562 413404
rect 382273 413402 382339 413405
rect 382406 413402 382412 413404
rect 382273 413400 382412 413402
rect 382273 413344 382278 413400
rect 382334 413344 382412 413400
rect 382273 413342 382412 413344
rect 382273 413339 382339 413342
rect 382406 413340 382412 413342
rect 382476 413340 382482 413404
rect 354489 413266 354555 413269
rect 373993 413266 374059 413269
rect 375373 413268 375439 413269
rect 374310 413266 374316 413268
rect 354489 413264 364626 413266
rect 354489 413208 354494 413264
rect 354550 413208 364626 413264
rect 354489 413206 364626 413208
rect 354489 413203 354555 413206
rect 354581 413130 354647 413133
rect 340462 413128 354647 413130
rect 340462 413072 354586 413128
rect 354642 413072 354647 413128
rect 340462 413070 354647 413072
rect 354581 413067 354647 413070
rect 364333 413130 364399 413133
rect 364566 413130 364626 413206
rect 373993 413264 374316 413266
rect 373993 413208 373998 413264
rect 374054 413208 374316 413264
rect 373993 413206 374316 413208
rect 373993 413203 374059 413206
rect 374310 413204 374316 413206
rect 374380 413204 374386 413268
rect 375373 413266 375420 413268
rect 375328 413264 375420 413266
rect 375328 413208 375378 413264
rect 375328 413206 375420 413208
rect 375373 413204 375420 413206
rect 375484 413204 375490 413268
rect 375557 413266 375623 413269
rect 375966 413266 375972 413268
rect 375557 413264 375972 413266
rect 375557 413208 375562 413264
rect 375618 413208 375972 413264
rect 375557 413206 375972 413208
rect 375373 413203 375439 413204
rect 375557 413203 375623 413206
rect 375966 413204 375972 413206
rect 376036 413204 376042 413268
rect 376753 413266 376819 413269
rect 377806 413266 377812 413268
rect 376753 413264 377812 413266
rect 376753 413208 376758 413264
rect 376814 413208 377812 413264
rect 376753 413206 377812 413208
rect 376753 413203 376819 413206
rect 377806 413204 377812 413206
rect 377876 413204 377882 413268
rect 378225 413266 378291 413269
rect 378910 413266 378916 413268
rect 378225 413264 378916 413266
rect 378225 413208 378230 413264
rect 378286 413208 378916 413264
rect 378225 413206 378916 413208
rect 378225 413203 378291 413206
rect 378910 413204 378916 413206
rect 378980 413204 378986 413268
rect 380617 413266 380683 413269
rect 387190 413266 387196 413268
rect 380617 413264 387196 413266
rect 380617 413208 380622 413264
rect 380678 413208 387196 413264
rect 380617 413206 387196 413208
rect 380617 413203 380683 413206
rect 387190 413204 387196 413206
rect 387260 413204 387266 413268
rect 393086 413266 393146 413478
rect 394693 413476 394740 413478
rect 394804 413476 394810 413540
rect 401542 413538 401548 413540
rect 397134 413478 401548 413538
rect 394693 413475 394759 413476
rect 393221 413402 393287 413405
rect 397134 413402 397194 413478
rect 401542 413476 401548 413478
rect 401612 413476 401618 413540
rect 404302 413476 404308 413540
rect 404372 413538 404419 413540
rect 480437 413538 480503 413541
rect 485773 413540 485839 413541
rect 480662 413538 480668 413540
rect 404372 413536 404464 413538
rect 404414 413480 404464 413536
rect 404372 413478 404464 413480
rect 480437 413536 480668 413538
rect 480437 413480 480442 413536
rect 480498 413480 480668 413536
rect 480437 413478 480668 413480
rect 404372 413476 404419 413478
rect 404353 413475 404419 413476
rect 480437 413475 480503 413478
rect 480662 413476 480668 413478
rect 480732 413476 480738 413540
rect 485773 413538 485820 413540
rect 485728 413536 485820 413538
rect 485728 413480 485778 413536
rect 485728 413478 485820 413480
rect 485773 413476 485820 413478
rect 485884 413476 485890 413540
rect 485773 413475 485839 413476
rect 397453 413404 397519 413405
rect 397453 413402 397500 413404
rect 393221 413400 397194 413402
rect 393221 413344 393226 413400
rect 393282 413344 397194 413400
rect 393221 413342 397194 413344
rect 397408 413400 397500 413402
rect 397408 413344 397458 413400
rect 397408 413342 397500 413344
rect 393221 413339 393287 413342
rect 397453 413340 397500 413342
rect 397564 413340 397570 413404
rect 401593 413402 401659 413405
rect 402278 413402 402284 413404
rect 401593 413400 402284 413402
rect 401593 413344 401598 413400
rect 401654 413344 402284 413400
rect 401593 413342 402284 413344
rect 397453 413339 397519 413340
rect 401593 413339 401659 413342
rect 402278 413340 402284 413342
rect 402348 413340 402354 413404
rect 481633 413402 481699 413405
rect 481950 413402 481956 413404
rect 481633 413400 481956 413402
rect 481633 413344 481638 413400
rect 481694 413344 481956 413400
rect 481633 413342 481956 413344
rect 481633 413339 481699 413342
rect 481950 413340 481956 413342
rect 482020 413340 482026 413404
rect 483013 413402 483079 413405
rect 483422 413402 483428 413404
rect 483013 413400 483428 413402
rect 483013 413344 483018 413400
rect 483074 413344 483428 413400
rect 483013 413342 483428 413344
rect 483013 413339 483079 413342
rect 483422 413340 483428 413342
rect 483492 413340 483498 413404
rect 404670 413266 404676 413268
rect 393086 413206 404676 413266
rect 404670 413204 404676 413206
rect 404740 413204 404746 413268
rect 484393 413266 484459 413269
rect 488533 413268 488599 413269
rect 484526 413266 484532 413268
rect 484393 413264 484532 413266
rect 484393 413208 484398 413264
rect 484454 413208 484532 413264
rect 484393 413206 484532 413208
rect 484393 413203 484459 413206
rect 484526 413204 484532 413206
rect 484596 413204 484602 413268
rect 488533 413266 488580 413268
rect 488488 413264 488580 413266
rect 488488 413208 488538 413264
rect 488488 413206 488580 413208
rect 488533 413204 488580 413206
rect 488644 413204 488650 413268
rect 488533 413203 488599 413204
rect 368289 413130 368355 413133
rect 364333 413128 364442 413130
rect 364333 413072 364338 413128
rect 364394 413072 364442 413128
rect 364333 413067 364442 413072
rect 364566 413128 368355 413130
rect 364566 413072 368294 413128
rect 368350 413072 368355 413128
rect 364566 413070 368355 413072
rect 368289 413067 368355 413070
rect 368473 413130 368539 413133
rect 369526 413130 369532 413132
rect 368473 413128 369532 413130
rect 368473 413072 368478 413128
rect 368534 413072 369532 413128
rect 368473 413070 369532 413072
rect 368473 413067 368539 413070
rect 369526 413068 369532 413070
rect 369596 413068 369602 413132
rect 369853 413130 369919 413133
rect 370814 413130 370820 413132
rect 369853 413128 370820 413130
rect 369853 413072 369858 413128
rect 369914 413072 370820 413128
rect 369853 413070 370820 413072
rect 369853 413067 369919 413070
rect 370814 413068 370820 413070
rect 370884 413068 370890 413132
rect 370957 413130 371023 413133
rect 375465 413130 375531 413133
rect 382181 413132 382247 413133
rect 376518 413130 376524 413132
rect 370957 413128 375298 413130
rect 370957 413072 370962 413128
rect 371018 413072 375298 413128
rect 370957 413070 375298 413072
rect 370957 413067 371023 413070
rect 350441 412994 350507 412997
rect 354581 412994 354647 412997
rect 340094 412934 345674 412994
rect 331121 412931 331187 412934
rect 335261 412931 335327 412934
rect 335169 412858 335235 412861
rect 320590 412856 335235 412858
rect 320590 412800 335174 412856
rect 335230 412800 335235 412856
rect 320590 412798 335235 412800
rect 345614 412858 345674 412934
rect 350441 412992 354647 412994
rect 350441 412936 350446 412992
rect 350502 412936 354586 412992
rect 354642 412936 354647 412992
rect 350441 412934 354647 412936
rect 364382 412994 364442 413067
rect 373901 412994 373967 412997
rect 364382 412992 373967 412994
rect 364382 412936 373906 412992
rect 373962 412936 373967 412992
rect 364382 412934 373967 412936
rect 375238 412994 375298 413070
rect 375465 413128 376524 413130
rect 375465 413072 375470 413128
rect 375526 413072 376524 413128
rect 375465 413070 376524 413072
rect 375465 413067 375531 413070
rect 376518 413068 376524 413070
rect 376588 413068 376594 413132
rect 382181 413130 382228 413132
rect 382136 413128 382228 413130
rect 382136 413072 382186 413128
rect 382136 413070 382228 413072
rect 382181 413068 382228 413070
rect 382292 413068 382298 413132
rect 382365 413130 382431 413133
rect 382774 413130 382780 413132
rect 382365 413128 382780 413130
rect 382365 413072 382370 413128
rect 382426 413072 382780 413128
rect 382365 413070 382780 413072
rect 382181 413067 382247 413068
rect 382365 413067 382431 413070
rect 382774 413068 382780 413070
rect 382844 413068 382850 413132
rect 385033 413130 385099 413133
rect 385166 413130 385172 413132
rect 385033 413128 385172 413130
rect 385033 413072 385038 413128
rect 385094 413072 385172 413128
rect 385033 413070 385172 413072
rect 385033 413067 385099 413070
rect 385166 413068 385172 413070
rect 385236 413068 385242 413132
rect 385309 413130 385375 413133
rect 391790 413130 391796 413132
rect 385309 413128 391796 413130
rect 385309 413072 385314 413128
rect 385370 413072 391796 413128
rect 385309 413070 391796 413072
rect 385309 413067 385375 413070
rect 391790 413068 391796 413070
rect 391860 413068 391866 413132
rect 397545 413130 397611 413133
rect 398046 413130 398052 413132
rect 397545 413128 398052 413130
rect 397545 413072 397550 413128
rect 397606 413072 398052 413128
rect 397545 413070 398052 413072
rect 397545 413067 397611 413070
rect 398046 413068 398052 413070
rect 398116 413068 398122 413132
rect 398833 413130 398899 413133
rect 399886 413130 399892 413132
rect 398833 413128 399892 413130
rect 398833 413072 398838 413128
rect 398894 413072 399892 413128
rect 398833 413070 399892 413072
rect 398833 413067 398899 413070
rect 399886 413068 399892 413070
rect 399956 413068 399962 413132
rect 487153 413130 487219 413133
rect 487286 413130 487292 413132
rect 487153 413128 487292 413130
rect 487153 413072 487158 413128
rect 487214 413072 487292 413128
rect 487153 413070 487292 413072
rect 487153 413067 487219 413070
rect 487286 413068 487292 413070
rect 487356 413068 487362 413132
rect 389081 412994 389147 412997
rect 375238 412992 389147 412994
rect 375238 412936 389086 412992
rect 389142 412936 389147 412992
rect 375238 412934 389147 412936
rect 350441 412931 350507 412934
rect 354581 412931 354647 412934
rect 373901 412931 373967 412934
rect 389081 412931 389147 412934
rect 389265 412994 389331 412997
rect 389766 412994 389772 412996
rect 389265 412992 389772 412994
rect 389265 412936 389270 412992
rect 389326 412936 389772 412992
rect 389265 412934 389772 412936
rect 389265 412931 389331 412934
rect 389766 412932 389772 412934
rect 389836 412932 389842 412996
rect 390553 412994 390619 412997
rect 391054 412994 391060 412996
rect 390553 412992 391060 412994
rect 390553 412936 390558 412992
rect 390614 412936 391060 412992
rect 390553 412934 391060 412936
rect 390553 412931 390619 412934
rect 391054 412932 391060 412934
rect 391124 412932 391130 412996
rect 393313 412994 393379 412997
rect 393446 412994 393452 412996
rect 393313 412992 393452 412994
rect 393313 412936 393318 412992
rect 393374 412936 393452 412992
rect 393313 412934 393452 412936
rect 393313 412931 393379 412934
rect 393446 412932 393452 412934
rect 393516 412932 393522 412996
rect 396073 412994 396139 412997
rect 396390 412994 396396 412996
rect 396073 412992 396396 412994
rect 396073 412936 396078 412992
rect 396134 412936 396396 412992
rect 396073 412934 396396 412936
rect 396073 412931 396139 412934
rect 396390 412932 396396 412934
rect 396460 412932 396466 412996
rect 397453 412994 397519 412997
rect 398598 412994 398604 412996
rect 397453 412992 398604 412994
rect 397453 412936 397458 412992
rect 397514 412936 398604 412992
rect 397453 412934 398604 412936
rect 397453 412931 397519 412934
rect 398598 412932 398604 412934
rect 398668 412932 398674 412996
rect 489913 412994 489979 412997
rect 491293 412996 491359 412997
rect 490046 412994 490052 412996
rect 489913 412992 490052 412994
rect 489913 412936 489918 412992
rect 489974 412936 490052 412992
rect 489913 412934 490052 412936
rect 489913 412931 489979 412934
rect 490046 412932 490052 412934
rect 490116 412932 490122 412996
rect 491293 412994 491340 412996
rect 491248 412992 491340 412994
rect 491248 412936 491298 412992
rect 491248 412934 491340 412936
rect 491293 412932 491340 412934
rect 491404 412932 491410 412996
rect 491293 412931 491359 412932
rect 354489 412858 354555 412861
rect 345614 412856 354555 412858
rect 345614 412800 354494 412856
rect 354550 412800 354555 412856
rect 345614 412798 354555 412800
rect 306465 412795 306531 412798
rect 315849 412795 315915 412798
rect 335169 412795 335235 412798
rect 354489 412795 354555 412798
rect 364333 412858 364399 412861
rect 371325 412858 371391 412861
rect 373993 412860 374059 412861
rect 364333 412856 371391 412858
rect 364333 412800 364338 412856
rect 364394 412800 371330 412856
rect 371386 412800 371391 412856
rect 364333 412798 371391 412800
rect 364333 412795 364399 412798
rect 371325 412795 371391 412798
rect 373942 412796 373948 412860
rect 374012 412858 374059 412860
rect 376753 412858 376819 412861
rect 378133 412860 378199 412861
rect 379605 412860 379671 412861
rect 377254 412858 377260 412860
rect 374012 412856 374104 412858
rect 374054 412800 374104 412856
rect 374012 412798 374104 412800
rect 376753 412856 377260 412858
rect 376753 412800 376758 412856
rect 376814 412800 377260 412856
rect 376753 412798 377260 412800
rect 374012 412796 374059 412798
rect 373993 412795 374059 412796
rect 376753 412795 376819 412798
rect 377254 412796 377260 412798
rect 377324 412796 377330 412860
rect 378133 412858 378180 412860
rect 378088 412856 378180 412858
rect 378088 412800 378138 412856
rect 378088 412798 378180 412800
rect 378133 412796 378180 412798
rect 378244 412796 378250 412860
rect 379605 412858 379652 412860
rect 379560 412856 379652 412858
rect 379560 412800 379610 412856
rect 379560 412798 379652 412800
rect 379605 412796 379652 412798
rect 379716 412796 379722 412860
rect 379789 412858 379855 412861
rect 393221 412858 393287 412861
rect 379789 412856 393287 412858
rect 379789 412800 379794 412856
rect 379850 412800 393226 412856
rect 393282 412800 393287 412856
rect 379789 412798 393287 412800
rect 378133 412795 378199 412796
rect 379605 412795 379671 412796
rect 379789 412795 379855 412798
rect 393221 412795 393287 412798
rect 394693 412858 394759 412861
rect 395286 412858 395292 412860
rect 394693 412856 395292 412858
rect 394693 412800 394698 412856
rect 394754 412800 395292 412856
rect 394693 412798 395292 412800
rect 394693 412795 394759 412798
rect 395286 412796 395292 412798
rect 395356 412796 395362 412860
rect 400213 412858 400279 412861
rect 400438 412858 400444 412860
rect 400213 412856 400444 412858
rect 400213 412800 400218 412856
rect 400274 412800 400444 412856
rect 400213 412798 400444 412800
rect 400213 412795 400279 412798
rect 400438 412796 400444 412798
rect 400508 412796 400514 412860
rect 403157 412858 403223 412861
rect 403382 412858 403388 412860
rect 403157 412856 403388 412858
rect 403157 412800 403162 412856
rect 403218 412800 403388 412856
rect 403157 412798 403388 412800
rect 403157 412795 403223 412798
rect 403382 412796 403388 412798
rect 403452 412796 403458 412860
rect 420177 412858 420243 412861
rect 522982 412858 522988 412860
rect 420177 412856 522988 412858
rect 420177 412800 420182 412856
rect 420238 412800 522988 412856
rect 420177 412798 522988 412800
rect 420177 412795 420243 412798
rect 522982 412796 522988 412798
rect 523052 412796 523058 412860
rect 367093 412722 367159 412725
rect 367686 412722 367692 412724
rect 367093 412720 367692 412722
rect 367093 412664 367098 412720
rect 367154 412664 367692 412720
rect 367093 412662 367692 412664
rect 367093 412659 367159 412662
rect 367686 412660 367692 412662
rect 367756 412660 367762 412724
rect 368289 412722 368355 412725
rect 370957 412722 371023 412725
rect 368289 412720 371023 412722
rect 368289 412664 368294 412720
rect 368350 412664 370962 412720
rect 371018 412664 371023 412720
rect 368289 412662 371023 412664
rect 368289 412659 368355 412662
rect 370957 412659 371023 412662
rect 371233 412722 371299 412725
rect 372613 412724 372679 412725
rect 371366 412722 371372 412724
rect 371233 412720 371372 412722
rect 371233 412664 371238 412720
rect 371294 412664 371372 412720
rect 371233 412662 371372 412664
rect 371233 412659 371299 412662
rect 371366 412660 371372 412662
rect 371436 412660 371442 412724
rect 372613 412722 372660 412724
rect 372568 412720 372660 412722
rect 372568 412664 372618 412720
rect 372568 412662 372660 412664
rect 372613 412660 372660 412662
rect 372724 412660 372730 412724
rect 374177 412722 374243 412725
rect 380893 412724 380959 412725
rect 374678 412722 374684 412724
rect 374177 412720 374684 412722
rect 374177 412664 374182 412720
rect 374238 412664 374684 412720
rect 374177 412662 374684 412664
rect 372613 412659 372679 412660
rect 374177 412659 374243 412662
rect 374678 412660 374684 412662
rect 374748 412660 374754 412724
rect 380893 412722 380940 412724
rect 380848 412720 380940 412722
rect 380848 412664 380898 412720
rect 380848 412662 380940 412664
rect 380893 412660 380940 412662
rect 381004 412660 381010 412724
rect 382273 412722 382339 412725
rect 383510 412722 383516 412724
rect 382273 412720 383516 412722
rect 382273 412664 382278 412720
rect 382334 412664 383516 412720
rect 382273 412662 383516 412664
rect 380893 412659 380959 412660
rect 382273 412659 382339 412662
rect 383510 412660 383516 412662
rect 383580 412660 383586 412724
rect 383653 412722 383719 412725
rect 384062 412722 384068 412724
rect 383653 412720 384068 412722
rect 383653 412664 383658 412720
rect 383714 412664 384068 412720
rect 383653 412662 384068 412664
rect 383653 412659 383719 412662
rect 384062 412660 384068 412662
rect 384132 412660 384138 412724
rect 385033 412722 385099 412725
rect 385902 412722 385908 412724
rect 385033 412720 385908 412722
rect 385033 412664 385038 412720
rect 385094 412664 385908 412720
rect 385033 412662 385908 412664
rect 385033 412659 385099 412662
rect 385902 412660 385908 412662
rect 385972 412660 385978 412724
rect 387057 412722 387123 412725
rect 387793 412722 387859 412725
rect 388110 412722 388116 412724
rect 387057 412720 387626 412722
rect 387057 412664 387062 412720
rect 387118 412664 387626 412720
rect 387057 412662 387626 412664
rect 387057 412659 387123 412662
rect 387566 412586 387626 412662
rect 387793 412720 388116 412722
rect 387793 412664 387798 412720
rect 387854 412664 388116 412720
rect 387793 412662 388116 412664
rect 387793 412659 387859 412662
rect 388110 412660 388116 412662
rect 388180 412660 388186 412724
rect 394182 412722 394188 412724
rect 388302 412662 394188 412722
rect 388302 412586 388362 412662
rect 394182 412660 394188 412662
rect 394252 412660 394258 412724
rect 398833 412722 398899 412725
rect 399150 412722 399156 412724
rect 398833 412720 399156 412722
rect 398833 412664 398838 412720
rect 398894 412664 399156 412720
rect 398833 412662 399156 412664
rect 398833 412659 398899 412662
rect 399150 412660 399156 412662
rect 399220 412660 399226 412724
rect 400213 412722 400279 412725
rect 468109 412724 468175 412725
rect 469397 412724 469463 412725
rect 471973 412724 472039 412725
rect 401174 412722 401180 412724
rect 400213 412720 401180 412722
rect 400213 412664 400218 412720
rect 400274 412664 401180 412720
rect 400213 412662 401180 412664
rect 400213 412659 400279 412662
rect 401174 412660 401180 412662
rect 401244 412660 401250 412724
rect 468109 412720 468156 412724
rect 468220 412722 468226 412724
rect 468109 412664 468114 412720
rect 468109 412660 468156 412664
rect 468220 412662 468266 412722
rect 469397 412720 469444 412724
rect 469508 412722 469514 412724
rect 469397 412664 469402 412720
rect 468220 412660 468226 412662
rect 469397 412660 469444 412664
rect 469508 412662 469554 412722
rect 471973 412720 472020 412724
rect 472084 412722 472090 412724
rect 491385 412722 491451 412725
rect 491886 412722 491892 412724
rect 471973 412664 471978 412720
rect 469508 412660 469514 412662
rect 471973 412660 472020 412664
rect 472084 412662 472130 412722
rect 491385 412720 491892 412722
rect 491385 412664 491390 412720
rect 491446 412664 491892 412720
rect 491385 412662 491892 412664
rect 472084 412660 472090 412662
rect 468109 412659 468175 412660
rect 469397 412659 469463 412660
rect 471973 412659 472039 412660
rect 491385 412659 491451 412662
rect 491886 412660 491892 412662
rect 491956 412660 491962 412724
rect 492673 412722 492739 412725
rect 493174 412722 493180 412724
rect 492673 412720 493180 412722
rect 492673 412664 492678 412720
rect 492734 412664 493180 412720
rect 492673 412662 493180 412664
rect 492673 412659 492739 412662
rect 493174 412660 493180 412662
rect 493244 412660 493250 412724
rect 494053 412722 494119 412725
rect 495709 412724 495775 412725
rect 496813 412724 496879 412725
rect 498285 412724 498351 412725
rect 499573 412724 499639 412725
rect 501045 412724 501111 412725
rect 494462 412722 494468 412724
rect 494053 412720 494468 412722
rect 494053 412664 494058 412720
rect 494114 412664 494468 412720
rect 494053 412662 494468 412664
rect 494053 412659 494119 412662
rect 494462 412660 494468 412662
rect 494532 412660 494538 412724
rect 495709 412720 495756 412724
rect 495820 412722 495826 412724
rect 495709 412664 495714 412720
rect 495709 412660 495756 412664
rect 495820 412662 495866 412722
rect 496813 412720 496860 412724
rect 496924 412722 496930 412724
rect 496813 412664 496818 412720
rect 495820 412660 495826 412662
rect 496813 412660 496860 412664
rect 496924 412662 496970 412722
rect 498285 412720 498332 412724
rect 498396 412722 498402 412724
rect 498285 412664 498290 412720
rect 496924 412660 496930 412662
rect 498285 412660 498332 412664
rect 498396 412662 498442 412722
rect 499573 412720 499620 412724
rect 499684 412722 499690 412724
rect 499573 412664 499578 412720
rect 498396 412660 498402 412662
rect 499573 412660 499620 412664
rect 499684 412662 499730 412722
rect 501045 412720 501092 412724
rect 501156 412722 501162 412724
rect 502517 412722 502583 412725
rect 503713 412724 503779 412725
rect 502742 412722 502748 412724
rect 501045 412664 501050 412720
rect 499684 412660 499690 412662
rect 501045 412660 501092 412664
rect 501156 412662 501202 412722
rect 502517 412720 502748 412722
rect 502517 412664 502522 412720
rect 502578 412664 502748 412720
rect 502517 412662 502748 412664
rect 501156 412660 501162 412662
rect 495709 412659 495775 412660
rect 496813 412659 496879 412660
rect 498285 412659 498351 412660
rect 499573 412659 499639 412660
rect 501045 412659 501111 412660
rect 502517 412659 502583 412662
rect 502742 412660 502748 412662
rect 502812 412660 502818 412724
rect 503662 412722 503668 412724
rect 503622 412662 503668 412722
rect 503732 412720 503779 412724
rect 503774 412664 503779 412720
rect 503662 412660 503668 412662
rect 503732 412660 503779 412664
rect 503713 412659 503779 412660
rect 503989 412722 504055 412725
rect 504398 412722 504404 412724
rect 503989 412720 504404 412722
rect 503989 412664 503994 412720
rect 504050 412664 504404 412720
rect 503989 412662 504404 412664
rect 503989 412659 504055 412662
rect 504398 412660 504404 412662
rect 504468 412660 504474 412724
rect 517513 412722 517579 412725
rect 518014 412722 518020 412724
rect 517513 412720 518020 412722
rect 517513 412664 517518 412720
rect 517574 412664 518020 412720
rect 517513 412662 518020 412664
rect 517513 412659 517579 412662
rect 518014 412660 518020 412662
rect 518084 412660 518090 412724
rect 387566 412526 388362 412586
rect 282821 412314 282887 412317
rect 279956 412312 282887 412314
rect 279956 412256 282826 412312
rect 282882 412256 282887 412312
rect 279956 412254 282887 412256
rect 282821 412251 282887 412254
rect 405733 411500 405799 411501
rect 405733 411496 405760 411500
rect 405824 411498 405830 411500
rect 405733 411440 405738 411496
rect 405733 411436 405760 411440
rect 405824 411438 405890 411498
rect 405824 411436 405830 411438
rect 405733 411435 405799 411436
rect 282821 411226 282887 411229
rect 279956 411224 282887 411226
rect 279956 411168 282826 411224
rect 282882 411168 282887 411224
rect 279956 411166 282887 411168
rect 282821 411163 282887 411166
rect 473445 410412 473511 410413
rect 473440 410410 473446 410412
rect 473354 410350 473446 410410
rect 473440 410348 473446 410350
rect 473510 410348 473516 410412
rect 473445 410347 473511 410348
rect 282729 410274 282795 410277
rect 279956 410272 282795 410274
rect 279956 410216 282734 410272
rect 282790 410216 282795 410272
rect 279956 410214 282795 410216
rect 282729 410211 282795 410214
rect 526437 410002 526503 410005
rect 526437 410000 526546 410002
rect 526437 409944 526442 410000
rect 526498 409944 526546 410000
rect 526437 409939 526546 409944
rect 526486 409683 526546 409939
rect -960 409172 480 409412
rect 281717 409322 281783 409325
rect 279956 409320 281783 409322
rect 279956 409264 281722 409320
rect 281778 409264 281783 409320
rect 279956 409262 281783 409264
rect 281717 409259 281783 409262
rect 281717 408234 281783 408237
rect 279956 408232 281783 408234
rect 279956 408176 281722 408232
rect 281778 408176 281783 408232
rect 279956 408174 281783 408176
rect 281717 408171 281783 408174
rect 282821 407282 282887 407285
rect 279956 407280 282887 407282
rect 279956 407224 282826 407280
rect 282882 407224 282887 407280
rect 279956 407222 282887 407224
rect 282821 407219 282887 407222
rect 282361 406194 282427 406197
rect 279956 406192 282427 406194
rect 279956 406136 282366 406192
rect 282422 406136 282427 406192
rect 279956 406134 282427 406136
rect 282361 406131 282427 406134
rect 282821 405242 282887 405245
rect 279956 405240 282887 405242
rect 279956 405184 282826 405240
rect 282882 405184 282887 405240
rect 279956 405182 282887 405184
rect 282821 405179 282887 405182
rect 583520 404684 584960 404924
rect 282821 404290 282887 404293
rect 279956 404288 282887 404290
rect 279956 404232 282826 404288
rect 282882 404232 282887 404288
rect 279956 404230 282887 404232
rect 282821 404227 282887 404230
rect 281625 403202 281691 403205
rect 279956 403200 281691 403202
rect 279956 403144 281630 403200
rect 281686 403144 281691 403200
rect 279956 403142 281691 403144
rect 281625 403139 281691 403142
rect 282821 402250 282887 402253
rect 279956 402248 282887 402250
rect 279956 402192 282826 402248
rect 282882 402192 282887 402248
rect 279956 402190 282887 402192
rect 282821 402187 282887 402190
rect 282821 401162 282887 401165
rect 279956 401160 282887 401162
rect 279956 401104 282826 401160
rect 282882 401104 282887 401160
rect 279956 401102 282887 401104
rect 282821 401099 282887 401102
rect 282821 400210 282887 400213
rect 279956 400208 282887 400210
rect 279956 400152 282826 400208
rect 282882 400152 282887 400208
rect 279956 400150 282887 400152
rect 282821 400147 282887 400150
rect 282269 399122 282335 399125
rect 279956 399120 282335 399122
rect 279956 399064 282274 399120
rect 282330 399064 282335 399120
rect 279956 399062 282335 399064
rect 282269 399059 282335 399062
rect 281625 398170 281691 398173
rect 279956 398168 281691 398170
rect 279956 398112 281630 398168
rect 281686 398112 281691 398168
rect 279956 398110 281691 398112
rect 281625 398107 281691 398110
rect 281625 397218 281691 397221
rect 279956 397216 281691 397218
rect 279956 397160 281630 397216
rect 281686 397160 281691 397216
rect 279956 397158 281691 397160
rect 281625 397155 281691 397158
rect 281625 396130 281691 396133
rect 279956 396128 281691 396130
rect 279956 396072 281630 396128
rect 281686 396072 281691 396128
rect 279956 396070 281691 396072
rect 281625 396067 281691 396070
rect 281625 395178 281691 395181
rect 279956 395176 281691 395178
rect -960 394892 480 395132
rect 279956 395120 281630 395176
rect 281686 395120 281691 395176
rect 279956 395118 281691 395120
rect 281625 395115 281691 395118
rect 281625 394090 281691 394093
rect 279956 394088 281691 394090
rect 279956 394032 281630 394088
rect 281686 394032 281691 394088
rect 279956 394030 281691 394032
rect 281625 394027 281691 394030
rect 281625 393138 281691 393141
rect 279956 393136 281691 393138
rect 279956 393080 281630 393136
rect 281686 393080 281691 393136
rect 279956 393078 281691 393080
rect 281625 393075 281691 393078
rect 416773 393002 416839 393005
rect 416773 393000 416882 393002
rect 416773 392944 416778 393000
rect 416834 392944 416882 393000
rect 416773 392939 416882 392944
rect 416822 392692 416882 392939
rect 583520 392852 584960 393092
rect 281625 392050 281691 392053
rect 279956 392048 281691 392050
rect 279956 391992 281630 392048
rect 281686 391992 281691 392048
rect 279956 391990 281691 391992
rect 281625 391987 281691 391990
rect 416405 391370 416471 391373
rect 416405 391368 416514 391370
rect 416405 391312 416410 391368
rect 416466 391312 416514 391368
rect 416405 391307 416514 391312
rect 281625 391098 281691 391101
rect 279956 391096 281691 391098
rect 279956 391040 281630 391096
rect 281686 391040 281691 391096
rect 279956 391038 281691 391040
rect 281625 391035 281691 391038
rect 416454 390992 416514 391307
rect 281625 390146 281691 390149
rect 279956 390144 281691 390146
rect 279956 390088 281630 390144
rect 281686 390088 281691 390144
rect 279956 390086 281691 390088
rect 281625 390083 281691 390086
rect 281625 389058 281691 389061
rect 279956 389056 281691 389058
rect 279956 389000 281630 389056
rect 281686 389000 281691 389056
rect 279956 388998 281691 389000
rect 281625 388995 281691 388998
rect 281625 388106 281691 388109
rect 279956 388104 281691 388106
rect 279956 388048 281630 388104
rect 281686 388048 281691 388104
rect 279956 388046 281691 388048
rect 281625 388043 281691 388046
rect 281625 387018 281691 387021
rect 279956 387016 281691 387018
rect 279956 386960 281630 387016
rect 281686 386960 281691 387016
rect 279956 386958 281691 386960
rect 281625 386955 281691 386958
rect 281625 386066 281691 386069
rect 279956 386064 281691 386066
rect 279956 386008 281630 386064
rect 281686 386008 281691 386064
rect 279956 386006 281691 386008
rect 281625 386003 281691 386006
rect 281625 385114 281691 385117
rect 279956 385112 281691 385114
rect 279956 385056 281630 385112
rect 281686 385056 281691 385112
rect 279956 385054 281691 385056
rect 281625 385051 281691 385054
rect 281625 384026 281691 384029
rect 279956 384024 281691 384026
rect 279956 383968 281630 384024
rect 281686 383968 281691 384024
rect 279956 383966 281691 383968
rect 281625 383963 281691 383966
rect 281625 383074 281691 383077
rect 279956 383072 281691 383074
rect 279956 383016 281630 383072
rect 281686 383016 281691 383072
rect 279956 383014 281691 383016
rect 281625 383011 281691 383014
rect 281625 381986 281691 381989
rect 279956 381984 281691 381986
rect 279956 381928 281630 381984
rect 281686 381928 281691 381984
rect 279956 381926 281691 381928
rect 281625 381923 281691 381926
rect 583520 381156 584960 381396
rect 281809 381034 281875 381037
rect 279956 381032 281875 381034
rect 279956 380976 281814 381032
rect 281870 380976 281875 381032
rect 279956 380974 281875 380976
rect 281809 380971 281875 380974
rect -960 380476 480 380716
rect 281625 379946 281691 379949
rect 279956 379944 281691 379946
rect 279956 379888 281630 379944
rect 281686 379888 281691 379944
rect 279956 379886 281691 379888
rect 281625 379883 281691 379886
rect 281625 378994 281691 378997
rect 279956 378992 281691 378994
rect 279956 378936 281630 378992
rect 281686 378936 281691 378992
rect 279956 378934 281691 378936
rect 281625 378931 281691 378934
rect 281625 378042 281691 378045
rect 279956 378040 281691 378042
rect 279956 377984 281630 378040
rect 281686 377984 281691 378040
rect 279956 377982 281691 377984
rect 281625 377979 281691 377982
rect 281809 376954 281875 376957
rect 279956 376952 281875 376954
rect 279956 376896 281814 376952
rect 281870 376896 281875 376952
rect 279956 376894 281875 376896
rect 281809 376891 281875 376894
rect 281625 376002 281691 376005
rect 279956 376000 281691 376002
rect 279956 375944 281630 376000
rect 281686 375944 281691 376000
rect 279956 375942 281691 375944
rect 281625 375939 281691 375942
rect 281625 374914 281691 374917
rect 279956 374912 281691 374914
rect 279956 374856 281630 374912
rect 281686 374856 281691 374912
rect 279956 374854 281691 374856
rect 281625 374851 281691 374854
rect 281625 373962 281691 373965
rect 279956 373960 281691 373962
rect 279956 373904 281630 373960
rect 281686 373904 281691 373960
rect 279956 373902 281691 373904
rect 281625 373899 281691 373902
rect 281809 372874 281875 372877
rect 279956 372872 281875 372874
rect 279956 372816 281814 372872
rect 281870 372816 281875 372872
rect 279956 372814 281875 372816
rect 281809 372811 281875 372814
rect 281625 371922 281691 371925
rect 279956 371920 281691 371922
rect 279956 371864 281630 371920
rect 281686 371864 281691 371920
rect 279956 371862 281691 371864
rect 281625 371859 281691 371862
rect 281625 370970 281691 370973
rect 279956 370968 281691 370970
rect 279956 370912 281630 370968
rect 281686 370912 281691 370968
rect 279956 370910 281691 370912
rect 281625 370907 281691 370910
rect 281809 369882 281875 369885
rect 279956 369880 281875 369882
rect 279956 369824 281814 369880
rect 281870 369824 281875 369880
rect 279956 369822 281875 369824
rect 281809 369819 281875 369822
rect 583520 369460 584960 369700
rect 281625 368930 281691 368933
rect 279956 368928 281691 368930
rect 279956 368872 281630 368928
rect 281686 368872 281691 368928
rect 279956 368870 281691 368872
rect 281625 368867 281691 368870
rect 281625 367842 281691 367845
rect 279956 367840 281691 367842
rect 279956 367784 281630 367840
rect 281686 367784 281691 367840
rect 279956 367782 281691 367784
rect 281625 367779 281691 367782
rect 284477 366890 284543 366893
rect 279956 366888 284543 366890
rect 279956 366832 284482 366888
rect 284538 366832 284543 366888
rect 279956 366830 284543 366832
rect 284477 366827 284543 366830
rect -960 366060 480 366300
rect 285121 365802 285187 365805
rect 279956 365800 285187 365802
rect 279956 365744 285126 365800
rect 285182 365744 285187 365800
rect 279956 365742 285187 365744
rect 285121 365739 285187 365742
rect 281625 364850 281691 364853
rect 279956 364848 281691 364850
rect 279956 364792 281630 364848
rect 281686 364792 281691 364848
rect 279956 364790 281691 364792
rect 281625 364787 281691 364790
rect 281625 363898 281691 363901
rect 279956 363896 281691 363898
rect 279956 363840 281630 363896
rect 281686 363840 281691 363896
rect 279956 363838 281691 363840
rect 281625 363835 281691 363838
rect 281625 362810 281691 362813
rect 279956 362808 281691 362810
rect 279956 362752 281630 362808
rect 281686 362752 281691 362808
rect 279956 362750 281691 362752
rect 281625 362747 281691 362750
rect 281809 361858 281875 361861
rect 279956 361856 281875 361858
rect 279956 361800 281814 361856
rect 281870 361800 281875 361856
rect 279956 361798 281875 361800
rect 281809 361795 281875 361798
rect 281625 360770 281691 360773
rect 279956 360768 281691 360770
rect 279956 360712 281630 360768
rect 281686 360712 281691 360768
rect 279956 360710 281691 360712
rect 281625 360707 281691 360710
rect 281625 359818 281691 359821
rect 279956 359816 281691 359818
rect 279956 359760 281630 359816
rect 281686 359760 281691 359816
rect 279956 359758 281691 359760
rect 281625 359755 281691 359758
rect 281809 358866 281875 358869
rect 279956 358864 281875 358866
rect 279956 358808 281814 358864
rect 281870 358808 281875 358864
rect 279956 358806 281875 358808
rect 281809 358803 281875 358806
rect 281625 357778 281691 357781
rect 279956 357776 281691 357778
rect 279956 357720 281630 357776
rect 281686 357720 281691 357776
rect 583520 357764 584960 358004
rect 279956 357718 281691 357720
rect 281625 357715 281691 357718
rect 282637 356826 282703 356829
rect 279956 356824 282703 356826
rect 279956 356768 282642 356824
rect 282698 356768 282703 356824
rect 279956 356766 282703 356768
rect 282637 356763 282703 356766
rect 282545 355738 282611 355741
rect 279956 355736 282611 355738
rect 279956 355680 282550 355736
rect 282606 355680 282611 355736
rect 279956 355678 282611 355680
rect 282545 355675 282611 355678
rect 282269 354786 282335 354789
rect 279956 354784 282335 354786
rect 279956 354728 282274 354784
rect 282330 354728 282335 354784
rect 279956 354726 282335 354728
rect 282269 354723 282335 354726
rect 282453 353698 282519 353701
rect 279956 353696 282519 353698
rect 279956 353640 282458 353696
rect 282514 353640 282519 353696
rect 279956 353638 282519 353640
rect 282453 353635 282519 353638
rect 282361 352746 282427 352749
rect 279956 352744 282427 352746
rect 279956 352688 282366 352744
rect 282422 352688 282427 352744
rect 279956 352686 282427 352688
rect 282361 352683 282427 352686
rect -960 351780 480 352020
rect 281625 351794 281691 351797
rect 279956 351792 281691 351794
rect 279956 351736 281630 351792
rect 281686 351736 281691 351792
rect 279956 351734 281691 351736
rect 281625 351731 281691 351734
rect 281625 350706 281691 350709
rect 279956 350704 281691 350706
rect 279956 350648 281630 350704
rect 281686 350648 281691 350704
rect 279956 350646 281691 350648
rect 281625 350643 281691 350646
rect 281625 349754 281691 349757
rect 279956 349752 281691 349754
rect 279956 349696 281630 349752
rect 281686 349696 281691 349752
rect 279956 349694 281691 349696
rect 281625 349691 281691 349694
rect 420085 349210 420151 349213
rect 420678 349210 420684 349212
rect 420085 349208 420684 349210
rect 420085 349152 420090 349208
rect 420146 349152 420684 349208
rect 420085 349150 420684 349152
rect 420085 349147 420151 349150
rect 420678 349148 420684 349150
rect 420748 349148 420754 349212
rect 527222 349210 527282 349412
rect 527582 349210 527588 349212
rect 527222 349150 527588 349210
rect 527582 349148 527588 349150
rect 527652 349148 527658 349212
rect 281625 348666 281691 348669
rect 279956 348664 281691 348666
rect 279956 348608 281630 348664
rect 281686 348608 281691 348664
rect 279956 348606 281691 348608
rect 281625 348603 281691 348606
rect 281625 347714 281691 347717
rect 279956 347712 281691 347714
rect 279956 347656 281630 347712
rect 281686 347656 281691 347712
rect 279956 347654 281691 347656
rect 281625 347651 281691 347654
rect 527222 347170 527282 347712
rect 527950 347170 527956 347172
rect 527222 347110 527956 347170
rect 527950 347108 527956 347110
rect 528020 347108 528026 347172
rect 281625 346626 281691 346629
rect 279956 346624 281691 346626
rect 279956 346568 281630 346624
rect 281686 346568 281691 346624
rect 279956 346566 281691 346568
rect 281625 346563 281691 346566
rect 419901 346628 419967 346629
rect 419901 346624 419948 346628
rect 420012 346626 420018 346628
rect 419901 346568 419906 346624
rect 419901 346564 419948 346568
rect 420012 346566 420058 346626
rect 420012 346564 420018 346566
rect 419901 346563 419967 346564
rect 419993 346490 420059 346493
rect 420678 346490 420684 346492
rect 419993 346488 420684 346490
rect 419993 346432 419998 346488
rect 420054 346432 420684 346488
rect 419993 346430 420684 346432
rect 419993 346427 420059 346430
rect 420678 346428 420684 346430
rect 420748 346428 420754 346492
rect 422886 346428 422892 346492
rect 422956 346490 422962 346492
rect 427854 346490 427860 346492
rect 422956 346430 427860 346490
rect 422956 346428 422962 346430
rect 427854 346428 427860 346430
rect 427924 346428 427930 346492
rect 446806 346428 446812 346492
rect 446876 346490 446882 346492
rect 447726 346490 447732 346492
rect 446876 346430 447732 346490
rect 446876 346428 446882 346430
rect 447726 346428 447732 346430
rect 447796 346428 447802 346492
rect 527222 346490 527282 346584
rect 527582 346490 527588 346492
rect 527222 346430 527588 346490
rect 527582 346428 527588 346430
rect 527652 346428 527658 346492
rect 583520 345932 584960 346172
rect 437974 345748 437980 345812
rect 438044 345810 438050 345812
rect 447174 345810 447180 345812
rect 438044 345750 447180 345810
rect 438044 345748 438050 345750
rect 447174 345748 447180 345750
rect 447244 345748 447250 345812
rect 281625 345674 281691 345677
rect 279956 345672 281691 345674
rect 279956 345616 281630 345672
rect 281686 345616 281691 345672
rect 279956 345614 281691 345616
rect 281625 345611 281691 345614
rect 527582 344914 527588 344916
rect 527252 344854 527588 344914
rect 527582 344852 527588 344854
rect 527652 344852 527658 344916
rect 281625 344722 281691 344725
rect 279956 344720 281691 344722
rect 279956 344664 281630 344720
rect 281686 344664 281691 344720
rect 279956 344662 281691 344664
rect 281625 344659 281691 344662
rect 419809 344450 419875 344453
rect 437790 344450 437796 344452
rect 419809 344448 437796 344450
rect 419809 344392 419814 344448
rect 419870 344392 437796 344448
rect 419809 344390 437796 344392
rect 419809 344387 419875 344390
rect 437790 344388 437796 344390
rect 437860 344388 437866 344452
rect 419717 343770 419783 343773
rect 420678 343770 420684 343772
rect 419717 343768 420684 343770
rect 419717 343712 419722 343768
rect 419778 343712 420684 343768
rect 419717 343710 420684 343712
rect 419717 343707 419783 343710
rect 420678 343708 420684 343710
rect 420748 343708 420754 343772
rect 281625 343634 281691 343637
rect 279956 343632 281691 343634
rect 279956 343576 281630 343632
rect 281686 343576 281691 343632
rect 279956 343574 281691 343576
rect 281625 343571 281691 343574
rect 527222 343226 527282 343756
rect 527950 343226 527956 343228
rect 527222 343166 527956 343226
rect 527950 343164 527956 343166
rect 528020 343164 528026 343228
rect 437606 343028 437612 343092
rect 437676 343090 437682 343092
rect 448094 343090 448100 343092
rect 437676 343030 448100 343090
rect 437676 343028 437682 343030
rect 448094 343028 448100 343030
rect 448164 343028 448170 343092
rect 449566 343028 449572 343092
rect 449636 343090 449642 343092
rect 450670 343090 450676 343092
rect 449636 343030 450676 343090
rect 449636 343028 449642 343030
rect 450670 343028 450676 343030
rect 450740 343028 450746 343092
rect 281809 342682 281875 342685
rect 279956 342680 281875 342682
rect 279956 342624 281814 342680
rect 281870 342624 281875 342680
rect 279956 342622 281875 342624
rect 281809 342619 281875 342622
rect 419625 341730 419691 341733
rect 420494 341730 420500 341732
rect 419625 341728 420500 341730
rect 419625 341672 419630 341728
rect 419686 341672 420500 341728
rect 419625 341670 420500 341672
rect 419625 341667 419691 341670
rect 420494 341668 420500 341670
rect 420564 341668 420570 341732
rect 527222 341730 527282 342056
rect 527582 341940 527588 342004
rect 527652 342002 527658 342004
rect 527652 341942 527834 342002
rect 527652 341940 527658 341942
rect 527582 341730 527588 341732
rect 527222 341670 527588 341730
rect 527582 341668 527588 341670
rect 527652 341668 527658 341732
rect 281625 341594 281691 341597
rect 527774 341594 527834 341942
rect 279956 341592 281691 341594
rect 279956 341536 281630 341592
rect 281686 341536 281691 341592
rect 279956 341534 281691 341536
rect 281625 341531 281691 341534
rect 527222 341534 527834 341594
rect 427854 341124 427860 341188
rect 427924 341186 427930 341188
rect 439446 341186 439452 341188
rect 427924 341126 439452 341186
rect 427924 341124 427930 341126
rect 439446 341124 439452 341126
rect 439516 341124 439522 341188
rect 419533 341050 419599 341053
rect 420494 341050 420500 341052
rect 419533 341048 420500 341050
rect 419533 340992 419538 341048
rect 419594 340992 420500 341048
rect 419533 340990 420500 340992
rect 419533 340987 419599 340990
rect 420494 340988 420500 340990
rect 420564 340988 420570 341052
rect 527222 340928 527282 341534
rect 281625 340642 281691 340645
rect 279956 340640 281691 340642
rect 279956 340584 281630 340640
rect 281686 340584 281691 340640
rect 279956 340582 281691 340584
rect 281625 340579 281691 340582
rect 444414 340308 444420 340372
rect 444484 340370 444490 340372
rect 445518 340370 445524 340372
rect 444484 340310 445524 340370
rect 444484 340308 444490 340310
rect 445518 340308 445524 340310
rect 445588 340308 445594 340372
rect 281717 339690 281783 339693
rect 279956 339688 281783 339690
rect 279956 339632 281722 339688
rect 281778 339632 281783 339688
rect 279956 339630 281783 339632
rect 281717 339627 281783 339630
rect 281625 338602 281691 338605
rect 279956 338600 281691 338602
rect 279956 338544 281630 338600
rect 281686 338544 281691 338600
rect 279956 338542 281691 338544
rect 281625 338539 281691 338542
rect 281625 337650 281691 337653
rect 279956 337648 281691 337650
rect -960 337364 480 337604
rect 279956 337592 281630 337648
rect 281686 337592 281691 337648
rect 279956 337590 281691 337592
rect 281625 337587 281691 337590
rect 281625 336562 281691 336565
rect 279956 336560 281691 336562
rect 279956 336504 281630 336560
rect 281686 336504 281691 336560
rect 279956 336502 281691 336504
rect 281625 336499 281691 336502
rect 281717 335610 281783 335613
rect 279956 335608 281783 335610
rect 279956 335552 281722 335608
rect 281778 335552 281783 335608
rect 279956 335550 281783 335552
rect 281717 335547 281783 335550
rect 281625 334522 281691 334525
rect 279956 334520 281691 334522
rect 279956 334464 281630 334520
rect 281686 334464 281691 334520
rect 279956 334462 281691 334464
rect 281625 334459 281691 334462
rect 583520 334236 584960 334476
rect 420085 333706 420151 333709
rect 417190 333704 420151 333706
rect 417190 333648 420090 333704
rect 420146 333648 420151 333704
rect 417190 333646 420151 333648
rect 281625 333570 281691 333573
rect 279956 333568 281691 333570
rect 279956 333512 281630 333568
rect 281686 333512 281691 333568
rect 279956 333510 281691 333512
rect 281625 333507 281691 333510
rect 417190 333144 417250 333646
rect 420085 333643 420151 333646
rect 281717 332618 281783 332621
rect 279956 332616 281783 332618
rect 279956 332560 281722 332616
rect 281778 332560 281783 332616
rect 279956 332558 281783 332560
rect 281717 332555 281783 332558
rect 419993 332074 420059 332077
rect 417190 332072 420059 332074
rect 417190 332016 419998 332072
rect 420054 332016 420059 332072
rect 417190 332014 420059 332016
rect 281901 331530 281967 331533
rect 279956 331528 281967 331530
rect 279956 331472 281906 331528
rect 281962 331472 281967 331528
rect 279956 331470 281967 331472
rect 281901 331467 281967 331470
rect 417190 331444 417250 332014
rect 419993 332011 420059 332014
rect 419901 330986 419967 330989
rect 417190 330984 419967 330986
rect 417190 330928 419906 330984
rect 419962 330928 419967 330984
rect 417190 330926 419967 330928
rect 281625 330578 281691 330581
rect 279956 330576 281691 330578
rect 279956 330520 281630 330576
rect 281686 330520 281691 330576
rect 279956 330518 281691 330520
rect 281625 330515 281691 330518
rect 417190 330316 417250 330926
rect 419901 330923 419967 330926
rect 281533 329490 281599 329493
rect 279956 329488 281599 329490
rect 279956 329432 281538 329488
rect 281594 329432 281599 329488
rect 279956 329430 281599 329432
rect 281533 329427 281599 329430
rect 419809 329218 419875 329221
rect 417190 329216 419875 329218
rect 417190 329160 419814 329216
rect 419870 329160 419875 329216
rect 417190 329158 419875 329160
rect 417190 328616 417250 329158
rect 419809 329155 419875 329158
rect 281625 328538 281691 328541
rect 279956 328536 281691 328538
rect 279956 328480 281630 328536
rect 281686 328480 281691 328536
rect 279956 328478 281691 328480
rect 281625 328475 281691 328478
rect 419717 328130 419783 328133
rect 417190 328128 419783 328130
rect 417190 328072 419722 328128
rect 419778 328072 419783 328128
rect 417190 328070 419783 328072
rect 417190 327488 417250 328070
rect 419717 328067 419783 328070
rect 281533 327450 281599 327453
rect 279956 327448 281599 327450
rect 279956 327392 281538 327448
rect 281594 327392 281599 327448
rect 279956 327390 281599 327392
rect 281533 327387 281599 327390
rect 282361 326498 282427 326501
rect 279956 326496 282427 326498
rect 279956 326440 282366 326496
rect 282422 326440 282427 326496
rect 279956 326438 282427 326440
rect 282361 326435 282427 326438
rect 419625 325818 419691 325821
rect 417220 325816 419691 325818
rect 417220 325760 419630 325816
rect 419686 325760 419691 325816
rect 417220 325758 419691 325760
rect 419625 325755 419691 325758
rect 281533 325546 281599 325549
rect 279956 325544 281599 325546
rect 279956 325488 281538 325544
rect 281594 325488 281599 325544
rect 279956 325486 281599 325488
rect 281533 325483 281599 325486
rect 419533 325138 419599 325141
rect 417190 325136 419599 325138
rect 417190 325080 419538 325136
rect 419594 325080 419599 325136
rect 417190 325078 419599 325080
rect 417190 324660 417250 325078
rect 419533 325075 419599 325078
rect 283414 324458 283420 324460
rect 279956 324398 283420 324458
rect 283414 324396 283420 324398
rect 283484 324396 283490 324460
rect 282310 323506 282316 323508
rect 279956 323446 282316 323506
rect 282310 323444 282316 323446
rect 282380 323444 282386 323508
rect -960 322948 480 323188
rect 583520 322540 584960 322780
rect 281717 322418 281783 322421
rect 279956 322416 281783 322418
rect 279956 322360 281722 322416
rect 281778 322360 281783 322416
rect 279956 322358 281783 322360
rect 281717 322355 281783 322358
rect 282821 321466 282887 321469
rect 279956 321464 282887 321466
rect 279956 321408 282826 321464
rect 282882 321408 282887 321464
rect 279956 321406 282887 321408
rect 282821 321403 282887 321406
rect 279325 320922 279391 320925
rect 279325 320920 279434 320922
rect 279325 320864 279330 320920
rect 279386 320864 279434 320920
rect 279325 320859 279434 320864
rect 279374 320484 279434 320859
rect 343633 318746 343699 318749
rect 343950 318746 343956 318748
rect 343633 318744 343956 318746
rect 343633 318688 343638 318744
rect 343694 318688 343956 318744
rect 343633 318686 343956 318688
rect 343633 318683 343699 318686
rect 343950 318684 343956 318686
rect 344020 318684 344026 318748
rect 453113 318746 453179 318749
rect 453246 318746 453252 318748
rect 453113 318744 453252 318746
rect 453113 318688 453118 318744
rect 453174 318688 453252 318744
rect 453113 318686 453252 318688
rect 453113 318683 453179 318686
rect 453246 318684 453252 318686
rect 453316 318684 453322 318748
rect 64781 318610 64847 318613
rect 165981 318610 166047 318613
rect 64781 318608 166047 318610
rect 64781 318552 64786 318608
rect 64842 318552 165986 318608
rect 166042 318552 166047 318608
rect 64781 318550 166047 318552
rect 64781 318547 64847 318550
rect 165981 318547 166047 318550
rect 74441 318474 74507 318477
rect 181529 318474 181595 318477
rect 74441 318472 181595 318474
rect 74441 318416 74446 318472
rect 74502 318416 181534 318472
rect 181590 318416 181595 318472
rect 74441 318414 181595 318416
rect 74441 318411 74507 318414
rect 181529 318411 181595 318414
rect 82629 318338 82695 318341
rect 193213 318338 193279 318341
rect 82629 318336 193279 318338
rect 82629 318280 82634 318336
rect 82690 318280 193218 318336
rect 193274 318280 193279 318336
rect 82629 318278 193279 318280
rect 82629 318275 82695 318278
rect 193213 318275 193279 318278
rect 82721 318202 82787 318205
rect 195145 318202 195211 318205
rect 82721 318200 195211 318202
rect 82721 318144 82726 318200
rect 82782 318144 195150 318200
rect 195206 318144 195211 318200
rect 82721 318142 195211 318144
rect 82721 318139 82787 318142
rect 195145 318139 195211 318142
rect 104801 318066 104867 318069
rect 230197 318066 230263 318069
rect 104801 318064 230263 318066
rect 104801 318008 104806 318064
rect 104862 318008 230202 318064
rect 230258 318008 230263 318064
rect 104801 318006 230263 318008
rect 104801 318003 104867 318006
rect 230197 318003 230263 318006
rect 583520 310708 584960 310948
rect -960 308668 480 308908
rect 583520 299012 584960 299252
rect -960 294252 480 294492
rect 583520 287316 584960 287556
rect -960 279972 480 280212
rect 583520 275620 584960 275860
rect -960 265556 480 265796
rect 583520 263788 584960 264028
rect 583520 252092 584960 252332
rect -960 251140 480 251380
rect 583520 240396 584960 240636
rect -960 236860 480 237100
rect 583520 228700 584960 228940
rect -960 222444 480 222684
rect 583520 216868 584960 217108
rect -960 208028 480 208268
rect 583520 205172 584960 205412
rect -960 193748 480 193988
rect 583520 193476 584960 193716
rect 583520 181780 584960 182020
rect -960 179332 480 179572
rect 583520 169948 584960 170188
rect -960 164916 480 165156
rect 583520 158252 584960 158492
rect -960 150636 480 150876
rect 583520 146556 584960 146796
rect -960 136220 480 136460
rect 583520 134724 584960 134964
rect 583520 123028 584960 123268
rect -960 121940 480 122180
rect 583520 111332 584960 111572
rect -960 107524 480 107764
rect 583520 99636 584960 99876
rect -960 93108 480 93348
rect 583520 87804 584960 88044
rect -960 78828 480 79068
rect 583520 76108 584960 76348
rect -960 64412 480 64652
rect 583520 64412 584960 64652
rect 583520 52716 584960 52956
rect -960 49996 480 50236
rect 583520 40884 584960 41124
rect -960 35716 480 35956
rect 583520 29188 584960 29428
rect -960 21300 480 21540
rect 583520 17492 584960 17732
rect -960 7020 480 7260
rect 583520 5796 584960 6036
rect 108757 5538 108823 5541
rect 237373 5538 237439 5541
rect 108757 5536 237439 5538
rect 108757 5480 108762 5536
rect 108818 5480 237378 5536
rect 237434 5480 237439 5536
rect 108757 5478 237439 5480
rect 108757 5475 108823 5478
rect 237373 5475 237439 5478
rect 112345 5402 112411 5405
rect 242893 5402 242959 5405
rect 112345 5400 242959 5402
rect 112345 5344 112350 5400
rect 112406 5344 242898 5400
rect 242954 5344 242959 5400
rect 112345 5342 242959 5344
rect 112345 5339 112411 5342
rect 242893 5339 242959 5342
rect 128997 5266 129063 5269
rect 270493 5266 270559 5269
rect 128997 5264 270559 5266
rect 128997 5208 129002 5264
rect 129058 5208 270498 5264
rect 270554 5208 270559 5264
rect 128997 5206 270559 5208
rect 128997 5203 129063 5206
rect 270493 5203 270559 5206
rect 127801 5130 127867 5133
rect 269113 5130 269179 5133
rect 127801 5128 269179 5130
rect 127801 5072 127806 5128
rect 127862 5072 269118 5128
rect 269174 5072 269179 5128
rect 127801 5070 269179 5072
rect 127801 5067 127867 5070
rect 269113 5067 269179 5070
rect 132585 4994 132651 4997
rect 276013 4994 276079 4997
rect 132585 4992 276079 4994
rect 132585 4936 132590 4992
rect 132646 4936 276018 4992
rect 276074 4936 276079 4992
rect 132585 4934 276079 4936
rect 132585 4931 132651 4934
rect 276013 4931 276079 4934
rect 115933 4858 115999 4861
rect 133137 4858 133203 4861
rect 115933 4856 133203 4858
rect 115933 4800 115938 4856
rect 115994 4800 133142 4856
rect 133198 4800 133203 4856
rect 115933 4798 133203 4800
rect 115933 4795 115999 4798
rect 133137 4795 133203 4798
rect 134885 4858 134951 4861
rect 278773 4858 278839 4861
rect 134885 4856 278839 4858
rect 134885 4800 134890 4856
rect 134946 4800 278778 4856
rect 278834 4800 278839 4856
rect 134885 4798 278839 4800
rect 134885 4795 134951 4798
rect 278773 4795 278839 4798
rect 55305 4178 55371 4181
rect 64689 4178 64755 4181
rect 55305 4176 64755 4178
rect 55305 4120 55310 4176
rect 55366 4120 64694 4176
rect 64750 4120 64755 4176
rect 55305 4118 64755 4120
rect 55305 4115 55371 4118
rect 64689 4115 64755 4118
rect 44541 4042 44607 4045
rect 123477 4042 123543 4045
rect 44541 4040 123543 4042
rect 44541 3984 44546 4040
rect 44602 3984 123482 4040
rect 123538 3984 123543 4040
rect 44541 3982 123543 3984
rect 44541 3979 44607 3982
rect 123477 3979 123543 3982
rect 40953 3906 41019 3909
rect 126973 3906 127039 3909
rect 40953 3904 127039 3906
rect 40953 3848 40958 3904
rect 41014 3848 126978 3904
rect 127034 3848 127039 3904
rect 40953 3846 127039 3848
rect 40953 3843 41019 3846
rect 126973 3843 127039 3846
rect 45737 3770 45803 3773
rect 133873 3770 133939 3773
rect 45737 3768 133939 3770
rect 45737 3712 45742 3768
rect 45798 3712 133878 3768
rect 133934 3712 133939 3768
rect 45737 3710 133939 3712
rect 45737 3707 45803 3710
rect 133873 3707 133939 3710
rect 54017 3634 54083 3637
rect 147673 3634 147739 3637
rect 54017 3632 147739 3634
rect 54017 3576 54022 3632
rect 54078 3576 147678 3632
rect 147734 3576 147739 3632
rect 54017 3574 147739 3576
rect 54017 3571 54083 3574
rect 147673 3571 147739 3574
rect 56409 3498 56475 3501
rect 151813 3498 151879 3501
rect 56409 3496 151879 3498
rect 56409 3440 56414 3496
rect 56470 3440 151818 3496
rect 151874 3440 151879 3496
rect 56409 3438 151879 3440
rect 56409 3435 56475 3438
rect 151813 3435 151879 3438
rect 121821 3362 121887 3365
rect 259453 3362 259519 3365
rect 121821 3360 259519 3362
rect 121821 3304 121826 3360
rect 121882 3304 259458 3360
rect 259514 3304 259519 3360
rect 121821 3302 259519 3304
rect 121821 3299 121887 3302
rect 259453 3299 259519 3302
<< via3 >>
rect 378180 652896 378244 652900
rect 378180 652840 378194 652896
rect 378194 652840 378244 652896
rect 378180 652836 378244 652840
rect 383516 652896 383580 652900
rect 383516 652840 383566 652896
rect 383566 652840 383580 652896
rect 383516 652836 383580 652840
rect 508452 652896 508516 652900
rect 508452 652840 508466 652896
rect 508466 652840 508516 652896
rect 508452 652836 508516 652840
rect 513420 652896 513484 652900
rect 513420 652840 513434 652896
rect 513434 652840 513484 652896
rect 513420 652836 513484 652840
rect 258576 651672 258640 651676
rect 258576 651616 258594 651672
rect 258594 651616 258640 651672
rect 258576 651612 258640 651616
rect 263571 651672 263635 651676
rect 263571 651616 263598 651672
rect 263598 651616 263635 651672
rect 263571 651612 263635 651616
rect 129228 651068 129292 651132
rect 133828 651068 133892 651132
rect 270356 587148 270420 587212
rect 387564 587148 387628 587212
rect 389220 580892 389284 580956
rect 518940 580892 519004 580956
rect 60596 578988 60660 579052
rect 188844 578988 188908 579052
rect 282500 578988 282564 579052
rect 310284 578988 310348 579052
rect 437428 578988 437492 579052
rect 211108 559948 211172 560012
rect 351868 559268 351932 559332
rect 358860 559268 358924 559332
rect 67404 558860 67468 558924
rect 68508 558860 68572 558924
rect 70164 558860 70228 558924
rect 71636 558920 71700 558924
rect 71636 558864 71686 558920
rect 71686 558864 71700 558920
rect 71636 558860 71700 558864
rect 72372 558860 72436 558924
rect 72924 558860 72988 558924
rect 73660 558920 73724 558924
rect 73660 558864 73710 558920
rect 73710 558864 73724 558920
rect 73660 558860 73724 558864
rect 74212 558920 74276 558924
rect 74212 558864 74262 558920
rect 74262 558864 74276 558920
rect 74212 558860 74276 558864
rect 74948 558920 75012 558924
rect 74948 558864 74998 558920
rect 74998 558864 75012 558920
rect 74948 558860 75012 558864
rect 75684 558860 75748 558924
rect 76788 558920 76852 558924
rect 76788 558864 76838 558920
rect 76838 558864 76852 558920
rect 76788 558860 76852 558864
rect 77340 558920 77404 558924
rect 77340 558864 77390 558920
rect 77390 558864 77404 558920
rect 77340 558860 77404 558864
rect 78076 558860 78140 558924
rect 79180 558860 79244 558924
rect 79916 558920 79980 558924
rect 79916 558864 79930 558920
rect 79930 558864 79980 558920
rect 79916 558860 79980 558864
rect 80652 558860 80716 558924
rect 81204 558920 81268 558924
rect 81204 558864 81254 558920
rect 81254 558864 81268 558920
rect 81204 558860 81268 558864
rect 81940 558920 82004 558924
rect 81940 558864 81990 558920
rect 81990 558864 82004 558920
rect 81940 558860 82004 558864
rect 82860 558920 82924 558924
rect 82860 558864 82910 558920
rect 82910 558864 82924 558920
rect 82860 558860 82924 558864
rect 83780 558920 83844 558924
rect 83780 558864 83830 558920
rect 83830 558864 83844 558920
rect 83780 558860 83844 558864
rect 84148 558920 84212 558924
rect 84148 558864 84198 558920
rect 84198 558864 84212 558920
rect 84148 558860 84212 558864
rect 85068 558860 85132 558924
rect 86356 558920 86420 558924
rect 86356 558864 86370 558920
rect 86370 558864 86420 558920
rect 86356 558860 86420 558864
rect 86724 558920 86788 558924
rect 86724 558864 86774 558920
rect 86774 558864 86788 558920
rect 86724 558860 86788 558864
rect 87828 558920 87892 558924
rect 87828 558864 87878 558920
rect 87878 558864 87892 558920
rect 87828 558860 87892 558864
rect 88196 558920 88260 558924
rect 88196 558864 88246 558920
rect 88246 558864 88260 558920
rect 88196 558860 88260 558864
rect 88932 558920 88996 558924
rect 88932 558864 88946 558920
rect 88946 558864 88996 558920
rect 88932 558860 88996 558864
rect 89116 558920 89180 558924
rect 89116 558864 89166 558920
rect 89166 558864 89180 558920
rect 89116 558860 89180 558864
rect 89852 558920 89916 558924
rect 89852 558864 89866 558920
rect 89866 558864 89916 558920
rect 89852 558860 89916 558864
rect 90956 558920 91020 558924
rect 90956 558864 91006 558920
rect 91006 558864 91020 558920
rect 90956 558860 91020 558864
rect 91876 558860 91940 558924
rect 92428 558920 92492 558924
rect 92428 558864 92478 558920
rect 92478 558864 92492 558920
rect 92428 558860 92492 558864
rect 93348 558920 93412 558924
rect 93348 558864 93362 558920
rect 93362 558864 93412 558920
rect 93348 558860 93412 558864
rect 93716 558920 93780 558924
rect 93716 558864 93766 558920
rect 93766 558864 93780 558920
rect 93716 558860 93780 558864
rect 95004 558920 95068 558924
rect 95004 558864 95054 558920
rect 95054 558864 95068 558920
rect 95004 558860 95068 558864
rect 95740 558920 95804 558924
rect 95740 558864 95754 558920
rect 95754 558864 95804 558920
rect 95740 558860 95804 558864
rect 96476 558920 96540 558924
rect 96476 558864 96526 558920
rect 96526 558864 96540 558920
rect 96476 558860 96540 558864
rect 97028 558860 97092 558924
rect 97764 558920 97828 558924
rect 97764 558864 97814 558920
rect 97814 558864 97828 558920
rect 97764 558860 97828 558864
rect 98316 558920 98380 558924
rect 98316 558864 98366 558920
rect 98366 558864 98380 558920
rect 98316 558860 98380 558864
rect 99052 558860 99116 558924
rect 99972 558920 100036 558924
rect 99972 558864 100022 558920
rect 100022 558864 100036 558920
rect 99972 558860 100036 558864
rect 101996 558920 102060 558924
rect 101996 558864 102046 558920
rect 102046 558864 102060 558920
rect 101996 558860 102060 558864
rect 104756 558920 104820 558924
rect 104756 558864 104806 558920
rect 104806 558864 104820 558920
rect 104756 558860 104820 558864
rect 107148 558860 107212 558924
rect 108436 558920 108500 558924
rect 108436 558864 108486 558920
rect 108486 558864 108500 558920
rect 108436 558860 108500 558864
rect 196204 558860 196268 558924
rect 200252 558920 200316 558924
rect 200252 558864 200266 558920
rect 200266 558864 200316 558920
rect 200252 558860 200316 558864
rect 202644 558860 202708 558924
rect 203748 558920 203812 558924
rect 203748 558864 203798 558920
rect 203798 558864 203812 558920
rect 203748 558860 203812 558864
rect 203932 558860 203996 558924
rect 205404 558860 205468 558924
rect 206140 558860 206204 558924
rect 208348 558860 208412 558924
rect 210556 558920 210620 558924
rect 210556 558864 210606 558920
rect 210606 558864 210620 558920
rect 210556 558860 210620 558864
rect 211844 558920 211908 558924
rect 211844 558864 211858 558920
rect 211858 558864 211908 558920
rect 211844 558860 211908 558864
rect 213132 558920 213196 558924
rect 213132 558864 213182 558920
rect 213182 558864 213196 558920
rect 213132 558860 213196 558864
rect 214052 558920 214116 558924
rect 214052 558864 214066 558920
rect 214066 558864 214116 558920
rect 214052 558860 214116 558864
rect 215340 558920 215404 558924
rect 215340 558864 215354 558920
rect 215354 558864 215404 558920
rect 215340 558860 215404 558864
rect 216628 558860 216692 558924
rect 218836 558920 218900 558924
rect 218836 558864 218850 558920
rect 218850 558864 218900 558920
rect 218836 558860 218900 558864
rect 220124 558920 220188 558924
rect 220124 558864 220138 558920
rect 220138 558864 220188 558920
rect 220124 558860 220188 558864
rect 221044 558920 221108 558924
rect 221044 558864 221094 558920
rect 221094 558864 221108 558920
rect 221044 558860 221108 558864
rect 222332 558860 222396 558924
rect 224540 558920 224604 558924
rect 224540 558864 224554 558920
rect 224554 558864 224604 558920
rect 224540 558860 224604 558864
rect 225828 558920 225892 558924
rect 225828 558864 225878 558920
rect 225878 558864 225892 558920
rect 225828 558860 225892 558864
rect 226196 558920 226260 558924
rect 226196 558864 226210 558920
rect 226210 558864 226260 558920
rect 226196 558860 226260 558864
rect 227116 558920 227180 558924
rect 227116 558864 227166 558920
rect 227166 558864 227180 558920
rect 227116 558860 227180 558864
rect 227484 558860 227548 558924
rect 228036 558920 228100 558924
rect 228036 558864 228050 558920
rect 228050 558864 228100 558920
rect 228036 558860 228100 558864
rect 228772 558860 228836 558924
rect 229508 558920 229572 558924
rect 229508 558864 229522 558920
rect 229522 558864 229572 558920
rect 229508 558860 229572 558864
rect 230244 558860 230308 558924
rect 230796 558860 230860 558924
rect 233004 558920 233068 558924
rect 233004 558864 233054 558920
rect 233054 558864 233068 558920
rect 233004 558860 233068 558864
rect 233556 558860 233620 558924
rect 234476 558920 234540 558924
rect 234476 558864 234526 558920
rect 234526 558864 234540 558920
rect 234476 558860 234540 558864
rect 235764 558860 235828 558924
rect 237236 558920 237300 558924
rect 237236 558864 237286 558920
rect 237286 558864 237300 558920
rect 237236 558860 237300 558864
rect 239628 558860 239692 558924
rect 313780 558920 313844 558924
rect 313780 558864 313830 558920
rect 313830 558864 313844 558920
rect 313780 558860 313844 558864
rect 317460 558920 317524 558924
rect 317460 558864 317474 558920
rect 317474 558864 317524 558920
rect 317460 558860 317524 558864
rect 318932 558860 318996 558924
rect 320220 558920 320284 558924
rect 320220 558864 320234 558920
rect 320234 558864 320284 558920
rect 320220 558860 320284 558864
rect 326292 558860 326356 558924
rect 327580 558860 327644 558924
rect 329604 558860 329668 558924
rect 331076 558860 331140 558924
rect 331812 558920 331876 558924
rect 331812 558864 331826 558920
rect 331826 558864 331876 558920
rect 331812 558860 331876 558864
rect 333284 558860 333348 558924
rect 334572 558860 334636 558924
rect 335860 558860 335924 558924
rect 336780 558920 336844 558924
rect 336780 558864 336794 558920
rect 336794 558864 336844 558920
rect 336780 558860 336844 558864
rect 337700 558860 337764 558924
rect 339172 558860 339236 558924
rect 340460 558860 340524 558924
rect 341748 558860 341812 558924
rect 342668 558860 342732 558924
rect 343956 558860 344020 558924
rect 344324 558920 344388 558924
rect 344324 558864 344338 558920
rect 344338 558864 344388 558920
rect 344324 558860 344388 558864
rect 346164 558860 346228 558924
rect 347452 558860 347516 558924
rect 348740 558860 348804 558924
rect 349660 558860 349724 558924
rect 352420 558860 352484 558924
rect 356100 558920 356164 558924
rect 356100 558864 356114 558920
rect 356114 558864 356164 558920
rect 356100 558860 356164 558864
rect 443132 558920 443196 558924
rect 443132 558864 443146 558920
rect 443146 558864 443196 558920
rect 443132 558860 443196 558864
rect 446260 558860 446324 558924
rect 451412 558860 451476 558924
rect 452884 558860 452948 558924
rect 453620 558920 453684 558924
rect 453620 558864 453670 558920
rect 453670 558864 453684 558920
rect 453620 558860 453684 558864
rect 455276 558860 455340 558924
rect 456564 558860 456628 558924
rect 457484 558860 457548 558924
rect 458772 558860 458836 558924
rect 460060 558860 460124 558924
rect 460980 558920 461044 558924
rect 460980 558864 461030 558920
rect 461030 558864 461044 558920
rect 460980 558860 461044 558864
rect 461716 558920 461780 558924
rect 461716 558864 461730 558920
rect 461730 558864 461780 558920
rect 461716 558860 461780 558864
rect 463372 558860 463436 558924
rect 464476 558860 464540 558924
rect 465764 558860 465828 558924
rect 466868 558860 466932 558924
rect 467972 558860 468036 558924
rect 468708 558920 468772 558924
rect 468708 558864 468758 558920
rect 468758 558864 468772 558920
rect 468708 558860 468772 558864
rect 470364 558860 470428 558924
rect 471468 558860 471532 558924
rect 472756 558860 472820 558924
rect 474044 558860 474108 558924
rect 474964 558860 475028 558924
rect 475516 558920 475580 558924
rect 475516 558864 475530 558920
rect 475530 558864 475580 558920
rect 475516 558860 475580 558864
rect 476252 558860 476316 558924
rect 476620 558920 476684 558924
rect 476620 558864 476634 558920
rect 476634 558864 476684 558920
rect 476620 558860 476684 558864
rect 477908 558860 477972 558924
rect 479012 558920 479076 558924
rect 479012 558864 479026 558920
rect 479026 558864 479076 558920
rect 479012 558860 479076 558864
rect 480484 558860 480548 558924
rect 64276 558724 64340 558788
rect 194364 558784 194428 558788
rect 194364 558728 194414 558784
rect 194414 558728 194428 558784
rect 194364 558724 194428 558728
rect 217548 558784 217612 558788
rect 217548 558728 217598 558784
rect 217598 558728 217612 558784
rect 217548 558724 217612 558728
rect 223620 558784 223684 558788
rect 223620 558728 223634 558784
rect 223634 558728 223684 558784
rect 223620 558724 223684 558728
rect 225644 558724 225708 558788
rect 231900 558784 231964 558788
rect 231900 558728 231914 558784
rect 231914 558728 231964 558784
rect 231900 558724 231964 558728
rect 232636 558724 232700 558788
rect 234660 558784 234724 558788
rect 234660 558728 234674 558784
rect 234674 558728 234724 558784
rect 234660 558724 234724 558728
rect 236132 558724 236196 558788
rect 237420 558784 237484 558788
rect 237420 558728 237434 558784
rect 237434 558728 237484 558784
rect 237420 558724 237484 558728
rect 320956 558724 321020 558788
rect 322612 558724 322676 558788
rect 326108 558724 326172 558788
rect 328868 558724 328932 558788
rect 330524 558784 330588 558788
rect 330524 558728 330538 558784
rect 330538 558728 330588 558784
rect 330524 558724 330588 558728
rect 333100 558784 333164 558788
rect 333100 558728 333150 558784
rect 333150 558728 333164 558784
rect 333100 558724 333164 558728
rect 334020 558784 334084 558788
rect 334020 558728 334070 558784
rect 334070 558728 334084 558784
rect 334020 558724 334084 558728
rect 335492 558784 335556 558788
rect 335492 558728 335506 558784
rect 335506 558728 335556 558784
rect 335492 558724 335556 558728
rect 336596 558784 336660 558788
rect 336596 558728 336646 558784
rect 336646 558728 336660 558784
rect 336596 558724 336660 558728
rect 337884 558724 337948 558788
rect 338988 558784 339052 558788
rect 338988 558728 339038 558784
rect 339038 558728 339052 558784
rect 338988 558724 339052 558728
rect 339908 558784 339972 558788
rect 339908 558728 339922 558784
rect 339922 558728 339972 558784
rect 339908 558724 339972 558728
rect 341196 558784 341260 558788
rect 341196 558728 341246 558784
rect 341246 558728 341260 558784
rect 341196 558724 341260 558728
rect 342484 558784 342548 558788
rect 342484 558728 342534 558784
rect 342534 558728 342548 558784
rect 342484 558724 342548 558728
rect 343588 558784 343652 558788
rect 343588 558728 343638 558784
rect 343638 558728 343652 558784
rect 343588 558724 343652 558728
rect 345980 558784 346044 558788
rect 345980 558728 346030 558784
rect 346030 558728 346044 558784
rect 345980 558724 346044 558728
rect 346900 558724 346964 558788
rect 348188 558784 348252 558788
rect 348188 558728 348238 558784
rect 348238 558728 348252 558784
rect 348188 558724 348252 558728
rect 349476 558724 349540 558788
rect 353524 558724 353588 558788
rect 354812 558724 354876 558788
rect 453804 558724 453868 558788
rect 454724 558784 454788 558788
rect 454724 558728 454774 558784
rect 454774 558728 454788 558784
rect 454724 558724 454788 558728
rect 456012 558784 456076 558788
rect 456012 558728 456062 558784
rect 456062 558728 456076 558784
rect 456012 558724 456076 558728
rect 457300 558724 457364 558788
rect 458404 558724 458468 558788
rect 462084 558724 462148 558788
rect 463004 558784 463068 558788
rect 463004 558728 463054 558784
rect 463054 558728 463068 558784
rect 463004 558724 463068 558728
rect 464292 558784 464356 558788
rect 464292 558728 464306 558784
rect 464306 558728 464356 558784
rect 464292 558724 464356 558728
rect 465212 558784 465276 558788
rect 465212 558728 465262 558784
rect 465262 558728 465276 558784
rect 465212 558724 465276 558728
rect 466500 558784 466564 558788
rect 466500 558728 466550 558784
rect 466550 558728 466564 558784
rect 466500 558724 466564 558728
rect 469076 558724 469140 558788
rect 471284 558784 471348 558788
rect 471284 558728 471334 558784
rect 471334 558728 471348 558784
rect 471284 558724 471348 558728
rect 472204 558784 472268 558788
rect 472204 558728 472218 558784
rect 472218 558728 472268 558784
rect 472204 558724 472268 558728
rect 473492 558784 473556 558788
rect 473492 558728 473506 558784
rect 473506 558728 473556 558784
rect 473492 558724 473556 558728
rect 474780 558784 474844 558788
rect 474780 558728 474830 558784
rect 474830 558728 474844 558784
rect 474780 558724 474844 558728
rect 484716 558724 484780 558788
rect 69796 558588 69860 558652
rect 75868 558648 75932 558652
rect 75868 558592 75918 558648
rect 75918 558592 75932 558648
rect 75868 558588 75932 558592
rect 78444 558648 78508 558652
rect 78444 558592 78494 558648
rect 78494 558592 78508 558648
rect 78444 558588 78508 558592
rect 79364 558648 79428 558652
rect 79364 558592 79414 558648
rect 79414 558592 79428 558648
rect 79364 558588 79428 558592
rect 85436 558648 85500 558652
rect 85436 558592 85450 558648
rect 85450 558592 85500 558648
rect 85436 558588 85500 558592
rect 86172 558588 86236 558652
rect 91140 558648 91204 558652
rect 91140 558592 91154 558648
rect 91154 558592 91204 558648
rect 91140 558588 91204 558592
rect 93164 558588 93228 558652
rect 94820 558648 94884 558652
rect 94820 558592 94834 558648
rect 94834 558592 94884 558648
rect 94820 558588 94884 558592
rect 106228 558648 106292 558652
rect 106228 558592 106278 558648
rect 106278 558592 106292 558648
rect 106228 558588 106292 558592
rect 202460 558588 202524 558652
rect 204852 558648 204916 558652
rect 204852 558592 204902 558648
rect 204902 558592 204916 558648
rect 204852 558588 204916 558592
rect 209636 558588 209700 558652
rect 323532 558648 323596 558652
rect 323532 558592 323582 558648
rect 323582 558592 323596 558648
rect 323532 558588 323596 558592
rect 324820 558588 324884 558652
rect 327028 558588 327092 558652
rect 328500 558588 328564 558652
rect 452700 558588 452764 558652
rect 459508 558588 459572 558652
rect 467788 558588 467852 558652
rect 469996 558648 470060 558652
rect 469996 558592 470046 558648
rect 470046 558592 470060 558648
rect 469996 558588 470060 558592
rect 477356 558588 477420 558652
rect 481588 558648 481652 558652
rect 481588 558592 481638 558648
rect 481638 558592 481652 558648
rect 481588 558588 481652 558592
rect 99604 558452 99668 558516
rect 108620 558452 108684 558516
rect 108988 558452 109052 558516
rect 232820 558452 232884 558516
rect 350580 558512 350644 558516
rect 350580 558456 350594 558512
rect 350594 558456 350644 558512
rect 350580 558452 350644 558456
rect 357572 558452 357636 558516
rect 479748 558452 479812 558516
rect 482140 558452 482204 558516
rect 483060 558512 483124 558516
rect 483060 558456 483074 558512
rect 483074 558456 483124 558512
rect 483060 558452 483124 558456
rect 486004 558452 486068 558516
rect 487292 558452 487356 558516
rect 197308 558316 197372 558380
rect 230612 558316 230676 558380
rect 238708 558376 238772 558380
rect 238708 558320 238758 558376
rect 238758 558320 238772 558376
rect 238708 558316 238772 558320
rect 282316 558316 282380 558380
rect 447364 558316 447428 558380
rect 478460 558316 478524 558380
rect 480852 558316 480916 558380
rect 488580 558376 488644 558380
rect 488580 558320 488594 558376
rect 488594 558320 488644 558376
rect 488580 558316 488644 558320
rect 198780 558180 198844 558244
rect 283420 558180 283484 558244
rect 448468 558180 448532 558244
rect 484164 558180 484228 558244
rect 238340 558044 238404 558108
rect 322796 558044 322860 558108
rect 324084 558044 324148 558108
rect 485636 558044 485700 558108
rect 82676 557968 82740 557972
rect 82676 557912 82726 557968
rect 82726 557912 82740 557968
rect 82676 557908 82740 557912
rect 107700 557908 107764 557972
rect 329788 557968 329852 557972
rect 329788 557912 329838 557968
rect 329838 557912 329852 557968
rect 329788 557908 329852 557912
rect 483428 557908 483492 557972
rect 486924 557908 486988 557972
rect 101628 557772 101692 557836
rect 316356 557832 316420 557836
rect 316356 557776 316370 557832
rect 316370 557776 316420 557832
rect 316356 557772 316420 557776
rect 332364 557772 332428 557836
rect 449940 557832 450004 557836
rect 449940 557776 449954 557832
rect 449954 557776 450004 557832
rect 449940 557772 450004 557776
rect 483612 557772 483676 557836
rect 487844 557772 487908 557836
rect 100156 557636 100220 557700
rect 106228 557636 106292 557700
rect 201540 557696 201604 557700
rect 201540 557640 201554 557696
rect 201554 557640 201604 557696
rect 201540 557636 201604 557640
rect 207060 557636 207124 557700
rect 210372 557636 210436 557700
rect 217364 557636 217428 557700
rect 325372 557636 325436 557700
rect 344876 557636 344940 557700
rect 353156 557636 353220 557700
rect 460796 557696 460860 557700
rect 460796 557640 460846 557696
rect 460846 557640 460860 557696
rect 460796 557636 460860 557640
rect 489132 557636 489196 557700
rect 101444 557500 101508 557564
rect 102732 557560 102796 557564
rect 102732 557504 102782 557560
rect 102782 557504 102796 557560
rect 102732 557500 102796 557504
rect 103284 557500 103348 557564
rect 104020 557500 104084 557564
rect 105308 557500 105372 557564
rect 106044 557500 106108 557564
rect 206876 557560 206940 557564
rect 206876 557504 206926 557560
rect 206926 557504 206940 557560
rect 206876 557500 206940 557504
rect 207980 557500 208044 557564
rect 209268 557500 209332 557564
rect 212396 557560 212460 557564
rect 212396 557504 212446 557560
rect 212446 557504 212460 557560
rect 212396 557500 212460 557504
rect 213500 557500 213564 557564
rect 214788 557500 214852 557564
rect 216260 557500 216324 557564
rect 217916 557560 217980 557564
rect 217916 557504 217930 557560
rect 217930 557504 217980 557560
rect 217916 557500 217980 557504
rect 219204 557500 219268 557564
rect 220676 557560 220740 557564
rect 220676 557504 220726 557560
rect 220726 557504 220740 557560
rect 220676 557500 220740 557504
rect 221964 557500 222028 557564
rect 223252 557500 223316 557564
rect 224356 557500 224420 557564
rect 350948 557500 351012 557564
rect 354444 557500 354508 557564
rect 355732 557500 355796 557564
rect 356652 557500 356716 557564
rect 357940 557500 358004 557564
rect 352236 555460 352300 555524
rect 359228 555460 359292 555524
rect 368244 413884 368308 413948
rect 368980 413884 369044 413948
rect 370268 413884 370332 413948
rect 371924 413884 371988 413948
rect 373028 413884 373092 413948
rect 380204 413884 380268 413948
rect 384620 413884 384684 413948
rect 388300 413884 388364 413948
rect 390692 413944 390756 413948
rect 390692 413888 390706 413944
rect 390706 413888 390756 413944
rect 390692 413884 390756 413888
rect 392900 413884 392964 413948
rect 389404 413612 389468 413676
rect 392164 413748 392228 413812
rect 397868 413884 397932 413948
rect 403020 413944 403084 413948
rect 403020 413888 403034 413944
rect 403034 413888 403084 413944
rect 403020 413884 403084 413888
rect 407804 413944 407868 413948
rect 407804 413888 407818 413944
rect 407818 413888 407868 413944
rect 407804 413884 407868 413888
rect 410564 413944 410628 413948
rect 410564 413888 410578 413944
rect 410578 413888 410628 413944
rect 410564 413884 410628 413888
rect 413876 413944 413940 413948
rect 413876 413888 413926 413944
rect 413926 413888 413940 413944
rect 413876 413884 413940 413888
rect 470916 413884 470980 413948
rect 474780 413944 474844 413948
rect 474780 413888 474830 413944
rect 474830 413888 474844 413944
rect 474780 413884 474844 413888
rect 478276 413884 478340 413948
rect 396028 413808 396092 413812
rect 396028 413752 396078 413808
rect 396078 413752 396092 413808
rect 396028 413748 396092 413752
rect 476252 413748 476316 413812
rect 477540 413808 477604 413812
rect 477540 413752 477554 413808
rect 477554 413752 477604 413808
rect 477540 413748 477604 413752
rect 505692 413748 505756 413812
rect 479380 413612 479444 413676
rect 506980 413612 507044 413676
rect 386460 413536 386524 413540
rect 386460 413480 386474 413536
rect 386474 413480 386524 413536
rect 386460 413476 386524 413480
rect 389220 413536 389284 413540
rect 389220 413480 389234 413536
rect 389234 413480 389284 413536
rect 389220 413476 389284 413480
rect 394740 413536 394804 413540
rect 394740 413480 394754 413536
rect 394754 413480 394804 413536
rect 381492 413340 381556 413404
rect 382412 413340 382476 413404
rect 374316 413204 374380 413268
rect 375420 413264 375484 413268
rect 375420 413208 375434 413264
rect 375434 413208 375484 413264
rect 375420 413204 375484 413208
rect 375972 413204 376036 413268
rect 377812 413204 377876 413268
rect 378916 413204 378980 413268
rect 387196 413204 387260 413268
rect 394740 413476 394804 413480
rect 401548 413476 401612 413540
rect 404308 413536 404372 413540
rect 404308 413480 404358 413536
rect 404358 413480 404372 413536
rect 404308 413476 404372 413480
rect 480668 413476 480732 413540
rect 485820 413536 485884 413540
rect 485820 413480 485834 413536
rect 485834 413480 485884 413536
rect 485820 413476 485884 413480
rect 397500 413400 397564 413404
rect 397500 413344 397514 413400
rect 397514 413344 397564 413400
rect 397500 413340 397564 413344
rect 402284 413340 402348 413404
rect 481956 413340 482020 413404
rect 483428 413340 483492 413404
rect 404676 413204 404740 413268
rect 484532 413204 484596 413268
rect 488580 413264 488644 413268
rect 488580 413208 488594 413264
rect 488594 413208 488644 413264
rect 488580 413204 488644 413208
rect 369532 413068 369596 413132
rect 370820 413068 370884 413132
rect 376524 413068 376588 413132
rect 382228 413128 382292 413132
rect 382228 413072 382242 413128
rect 382242 413072 382292 413128
rect 382228 413068 382292 413072
rect 382780 413068 382844 413132
rect 385172 413068 385236 413132
rect 391796 413068 391860 413132
rect 398052 413068 398116 413132
rect 399892 413068 399956 413132
rect 487292 413068 487356 413132
rect 389772 412932 389836 412996
rect 391060 412932 391124 412996
rect 393452 412932 393516 412996
rect 396396 412932 396460 412996
rect 398604 412932 398668 412996
rect 490052 412932 490116 412996
rect 491340 412992 491404 412996
rect 491340 412936 491354 412992
rect 491354 412936 491404 412992
rect 491340 412932 491404 412936
rect 373948 412856 374012 412860
rect 373948 412800 373998 412856
rect 373998 412800 374012 412856
rect 373948 412796 374012 412800
rect 377260 412796 377324 412860
rect 378180 412856 378244 412860
rect 378180 412800 378194 412856
rect 378194 412800 378244 412856
rect 378180 412796 378244 412800
rect 379652 412856 379716 412860
rect 379652 412800 379666 412856
rect 379666 412800 379716 412856
rect 379652 412796 379716 412800
rect 395292 412796 395356 412860
rect 400444 412796 400508 412860
rect 403388 412796 403452 412860
rect 522988 412796 523052 412860
rect 367692 412660 367756 412724
rect 371372 412660 371436 412724
rect 372660 412720 372724 412724
rect 372660 412664 372674 412720
rect 372674 412664 372724 412720
rect 372660 412660 372724 412664
rect 374684 412660 374748 412724
rect 380940 412720 381004 412724
rect 380940 412664 380954 412720
rect 380954 412664 381004 412720
rect 380940 412660 381004 412664
rect 383516 412660 383580 412724
rect 384068 412660 384132 412724
rect 385908 412660 385972 412724
rect 388116 412660 388180 412724
rect 394188 412660 394252 412724
rect 399156 412660 399220 412724
rect 401180 412660 401244 412724
rect 468156 412720 468220 412724
rect 468156 412664 468170 412720
rect 468170 412664 468220 412720
rect 468156 412660 468220 412664
rect 469444 412720 469508 412724
rect 469444 412664 469458 412720
rect 469458 412664 469508 412720
rect 469444 412660 469508 412664
rect 472020 412720 472084 412724
rect 472020 412664 472034 412720
rect 472034 412664 472084 412720
rect 472020 412660 472084 412664
rect 491892 412660 491956 412724
rect 493180 412660 493244 412724
rect 494468 412660 494532 412724
rect 495756 412720 495820 412724
rect 495756 412664 495770 412720
rect 495770 412664 495820 412720
rect 495756 412660 495820 412664
rect 496860 412720 496924 412724
rect 496860 412664 496874 412720
rect 496874 412664 496924 412720
rect 496860 412660 496924 412664
rect 498332 412720 498396 412724
rect 498332 412664 498346 412720
rect 498346 412664 498396 412720
rect 498332 412660 498396 412664
rect 499620 412720 499684 412724
rect 499620 412664 499634 412720
rect 499634 412664 499684 412720
rect 499620 412660 499684 412664
rect 501092 412720 501156 412724
rect 501092 412664 501106 412720
rect 501106 412664 501156 412720
rect 501092 412660 501156 412664
rect 502748 412660 502812 412724
rect 503668 412720 503732 412724
rect 503668 412664 503718 412720
rect 503718 412664 503732 412720
rect 503668 412660 503732 412664
rect 504404 412660 504468 412724
rect 518020 412660 518084 412724
rect 405760 411496 405824 411500
rect 405760 411440 405794 411496
rect 405794 411440 405824 411496
rect 405760 411436 405824 411440
rect 473446 410408 473510 410412
rect 473446 410352 473450 410408
rect 473450 410352 473506 410408
rect 473506 410352 473510 410408
rect 473446 410348 473510 410352
rect 420684 349148 420748 349212
rect 527588 349148 527652 349212
rect 527956 347108 528020 347172
rect 419948 346624 420012 346628
rect 419948 346568 419962 346624
rect 419962 346568 420012 346624
rect 419948 346564 420012 346568
rect 420684 346428 420748 346492
rect 422892 346428 422956 346492
rect 427860 346428 427924 346492
rect 446812 346428 446876 346492
rect 447732 346428 447796 346492
rect 527588 346428 527652 346492
rect 437980 345748 438044 345812
rect 447180 345748 447244 345812
rect 527588 344852 527652 344916
rect 437796 344388 437860 344452
rect 420684 343708 420748 343772
rect 527956 343164 528020 343228
rect 437612 343028 437676 343092
rect 448100 343028 448164 343092
rect 449572 343028 449636 343092
rect 450676 343028 450740 343092
rect 420500 341668 420564 341732
rect 527588 341940 527652 342004
rect 527588 341668 527652 341732
rect 427860 341124 427924 341188
rect 439452 341124 439516 341188
rect 420500 340988 420564 341052
rect 444420 340308 444484 340372
rect 445524 340308 445588 340372
rect 283420 324396 283484 324460
rect 282316 323444 282380 323508
rect 343956 318684 344020 318748
rect 453252 318684 453316 318748
<< metal4 >>
rect -8576 711418 -7976 711440
rect -8576 711182 -8394 711418
rect -8158 711182 -7976 711418
rect -8576 711098 -7976 711182
rect -8576 710862 -8394 711098
rect -8158 710862 -7976 711098
rect -8576 679254 -7976 710862
rect -8576 679018 -8394 679254
rect -8158 679018 -7976 679254
rect -8576 678934 -7976 679018
rect -8576 678698 -8394 678934
rect -8158 678698 -7976 678934
rect -8576 643254 -7976 678698
rect -8576 643018 -8394 643254
rect -8158 643018 -7976 643254
rect -8576 642934 -7976 643018
rect -8576 642698 -8394 642934
rect -8158 642698 -7976 642934
rect -8576 607254 -7976 642698
rect -8576 607018 -8394 607254
rect -8158 607018 -7976 607254
rect -8576 606934 -7976 607018
rect -8576 606698 -8394 606934
rect -8158 606698 -7976 606934
rect -8576 571254 -7976 606698
rect -8576 571018 -8394 571254
rect -8158 571018 -7976 571254
rect -8576 570934 -7976 571018
rect -8576 570698 -8394 570934
rect -8158 570698 -7976 570934
rect -8576 535254 -7976 570698
rect -8576 535018 -8394 535254
rect -8158 535018 -7976 535254
rect -8576 534934 -7976 535018
rect -8576 534698 -8394 534934
rect -8158 534698 -7976 534934
rect -8576 499254 -7976 534698
rect -8576 499018 -8394 499254
rect -8158 499018 -7976 499254
rect -8576 498934 -7976 499018
rect -8576 498698 -8394 498934
rect -8158 498698 -7976 498934
rect -8576 463254 -7976 498698
rect -8576 463018 -8394 463254
rect -8158 463018 -7976 463254
rect -8576 462934 -7976 463018
rect -8576 462698 -8394 462934
rect -8158 462698 -7976 462934
rect -8576 427254 -7976 462698
rect -8576 427018 -8394 427254
rect -8158 427018 -7976 427254
rect -8576 426934 -7976 427018
rect -8576 426698 -8394 426934
rect -8158 426698 -7976 426934
rect -8576 391254 -7976 426698
rect -8576 391018 -8394 391254
rect -8158 391018 -7976 391254
rect -8576 390934 -7976 391018
rect -8576 390698 -8394 390934
rect -8158 390698 -7976 390934
rect -8576 355254 -7976 390698
rect -8576 355018 -8394 355254
rect -8158 355018 -7976 355254
rect -8576 354934 -7976 355018
rect -8576 354698 -8394 354934
rect -8158 354698 -7976 354934
rect -8576 319254 -7976 354698
rect -8576 319018 -8394 319254
rect -8158 319018 -7976 319254
rect -8576 318934 -7976 319018
rect -8576 318698 -8394 318934
rect -8158 318698 -7976 318934
rect -8576 283254 -7976 318698
rect -8576 283018 -8394 283254
rect -8158 283018 -7976 283254
rect -8576 282934 -7976 283018
rect -8576 282698 -8394 282934
rect -8158 282698 -7976 282934
rect -8576 247254 -7976 282698
rect -8576 247018 -8394 247254
rect -8158 247018 -7976 247254
rect -8576 246934 -7976 247018
rect -8576 246698 -8394 246934
rect -8158 246698 -7976 246934
rect -8576 211254 -7976 246698
rect -8576 211018 -8394 211254
rect -8158 211018 -7976 211254
rect -8576 210934 -7976 211018
rect -8576 210698 -8394 210934
rect -8158 210698 -7976 210934
rect -8576 175254 -7976 210698
rect -8576 175018 -8394 175254
rect -8158 175018 -7976 175254
rect -8576 174934 -7976 175018
rect -8576 174698 -8394 174934
rect -8158 174698 -7976 174934
rect -8576 139254 -7976 174698
rect -8576 139018 -8394 139254
rect -8158 139018 -7976 139254
rect -8576 138934 -7976 139018
rect -8576 138698 -8394 138934
rect -8158 138698 -7976 138934
rect -8576 103254 -7976 138698
rect -8576 103018 -8394 103254
rect -8158 103018 -7976 103254
rect -8576 102934 -7976 103018
rect -8576 102698 -8394 102934
rect -8158 102698 -7976 102934
rect -8576 67254 -7976 102698
rect -8576 67018 -8394 67254
rect -8158 67018 -7976 67254
rect -8576 66934 -7976 67018
rect -8576 66698 -8394 66934
rect -8158 66698 -7976 66934
rect -8576 31254 -7976 66698
rect -8576 31018 -8394 31254
rect -8158 31018 -7976 31254
rect -8576 30934 -7976 31018
rect -8576 30698 -8394 30934
rect -8158 30698 -7976 30934
rect -8576 -6926 -7976 30698
rect -7636 710478 -7036 710500
rect -7636 710242 -7454 710478
rect -7218 710242 -7036 710478
rect -7636 710158 -7036 710242
rect -7636 709922 -7454 710158
rect -7218 709922 -7036 710158
rect -7636 697254 -7036 709922
rect 11604 710478 12204 711440
rect 11604 710242 11786 710478
rect 12022 710242 12204 710478
rect 11604 710158 12204 710242
rect 11604 709922 11786 710158
rect 12022 709922 12204 710158
rect -7636 697018 -7454 697254
rect -7218 697018 -7036 697254
rect -7636 696934 -7036 697018
rect -7636 696698 -7454 696934
rect -7218 696698 -7036 696934
rect -7636 661254 -7036 696698
rect -7636 661018 -7454 661254
rect -7218 661018 -7036 661254
rect -7636 660934 -7036 661018
rect -7636 660698 -7454 660934
rect -7218 660698 -7036 660934
rect -7636 625254 -7036 660698
rect -7636 625018 -7454 625254
rect -7218 625018 -7036 625254
rect -7636 624934 -7036 625018
rect -7636 624698 -7454 624934
rect -7218 624698 -7036 624934
rect -7636 589254 -7036 624698
rect -7636 589018 -7454 589254
rect -7218 589018 -7036 589254
rect -7636 588934 -7036 589018
rect -7636 588698 -7454 588934
rect -7218 588698 -7036 588934
rect -7636 553254 -7036 588698
rect -7636 553018 -7454 553254
rect -7218 553018 -7036 553254
rect -7636 552934 -7036 553018
rect -7636 552698 -7454 552934
rect -7218 552698 -7036 552934
rect -7636 517254 -7036 552698
rect -7636 517018 -7454 517254
rect -7218 517018 -7036 517254
rect -7636 516934 -7036 517018
rect -7636 516698 -7454 516934
rect -7218 516698 -7036 516934
rect -7636 481254 -7036 516698
rect -7636 481018 -7454 481254
rect -7218 481018 -7036 481254
rect -7636 480934 -7036 481018
rect -7636 480698 -7454 480934
rect -7218 480698 -7036 480934
rect -7636 445254 -7036 480698
rect -7636 445018 -7454 445254
rect -7218 445018 -7036 445254
rect -7636 444934 -7036 445018
rect -7636 444698 -7454 444934
rect -7218 444698 -7036 444934
rect -7636 409254 -7036 444698
rect -7636 409018 -7454 409254
rect -7218 409018 -7036 409254
rect -7636 408934 -7036 409018
rect -7636 408698 -7454 408934
rect -7218 408698 -7036 408934
rect -7636 373254 -7036 408698
rect -7636 373018 -7454 373254
rect -7218 373018 -7036 373254
rect -7636 372934 -7036 373018
rect -7636 372698 -7454 372934
rect -7218 372698 -7036 372934
rect -7636 337254 -7036 372698
rect -7636 337018 -7454 337254
rect -7218 337018 -7036 337254
rect -7636 336934 -7036 337018
rect -7636 336698 -7454 336934
rect -7218 336698 -7036 336934
rect -7636 301254 -7036 336698
rect -7636 301018 -7454 301254
rect -7218 301018 -7036 301254
rect -7636 300934 -7036 301018
rect -7636 300698 -7454 300934
rect -7218 300698 -7036 300934
rect -7636 265254 -7036 300698
rect -7636 265018 -7454 265254
rect -7218 265018 -7036 265254
rect -7636 264934 -7036 265018
rect -7636 264698 -7454 264934
rect -7218 264698 -7036 264934
rect -7636 229254 -7036 264698
rect -7636 229018 -7454 229254
rect -7218 229018 -7036 229254
rect -7636 228934 -7036 229018
rect -7636 228698 -7454 228934
rect -7218 228698 -7036 228934
rect -7636 193254 -7036 228698
rect -7636 193018 -7454 193254
rect -7218 193018 -7036 193254
rect -7636 192934 -7036 193018
rect -7636 192698 -7454 192934
rect -7218 192698 -7036 192934
rect -7636 157254 -7036 192698
rect -7636 157018 -7454 157254
rect -7218 157018 -7036 157254
rect -7636 156934 -7036 157018
rect -7636 156698 -7454 156934
rect -7218 156698 -7036 156934
rect -7636 121254 -7036 156698
rect -7636 121018 -7454 121254
rect -7218 121018 -7036 121254
rect -7636 120934 -7036 121018
rect -7636 120698 -7454 120934
rect -7218 120698 -7036 120934
rect -7636 85254 -7036 120698
rect -7636 85018 -7454 85254
rect -7218 85018 -7036 85254
rect -7636 84934 -7036 85018
rect -7636 84698 -7454 84934
rect -7218 84698 -7036 84934
rect -7636 49254 -7036 84698
rect -7636 49018 -7454 49254
rect -7218 49018 -7036 49254
rect -7636 48934 -7036 49018
rect -7636 48698 -7454 48934
rect -7218 48698 -7036 48934
rect -7636 13254 -7036 48698
rect -7636 13018 -7454 13254
rect -7218 13018 -7036 13254
rect -7636 12934 -7036 13018
rect -7636 12698 -7454 12934
rect -7218 12698 -7036 12934
rect -7636 -5986 -7036 12698
rect -6696 709538 -6096 709560
rect -6696 709302 -6514 709538
rect -6278 709302 -6096 709538
rect -6696 709218 -6096 709302
rect -6696 708982 -6514 709218
rect -6278 708982 -6096 709218
rect -6696 675654 -6096 708982
rect -6696 675418 -6514 675654
rect -6278 675418 -6096 675654
rect -6696 675334 -6096 675418
rect -6696 675098 -6514 675334
rect -6278 675098 -6096 675334
rect -6696 639654 -6096 675098
rect -6696 639418 -6514 639654
rect -6278 639418 -6096 639654
rect -6696 639334 -6096 639418
rect -6696 639098 -6514 639334
rect -6278 639098 -6096 639334
rect -6696 603654 -6096 639098
rect -6696 603418 -6514 603654
rect -6278 603418 -6096 603654
rect -6696 603334 -6096 603418
rect -6696 603098 -6514 603334
rect -6278 603098 -6096 603334
rect -6696 567654 -6096 603098
rect -6696 567418 -6514 567654
rect -6278 567418 -6096 567654
rect -6696 567334 -6096 567418
rect -6696 567098 -6514 567334
rect -6278 567098 -6096 567334
rect -6696 531654 -6096 567098
rect -6696 531418 -6514 531654
rect -6278 531418 -6096 531654
rect -6696 531334 -6096 531418
rect -6696 531098 -6514 531334
rect -6278 531098 -6096 531334
rect -6696 495654 -6096 531098
rect -6696 495418 -6514 495654
rect -6278 495418 -6096 495654
rect -6696 495334 -6096 495418
rect -6696 495098 -6514 495334
rect -6278 495098 -6096 495334
rect -6696 459654 -6096 495098
rect -6696 459418 -6514 459654
rect -6278 459418 -6096 459654
rect -6696 459334 -6096 459418
rect -6696 459098 -6514 459334
rect -6278 459098 -6096 459334
rect -6696 423654 -6096 459098
rect -6696 423418 -6514 423654
rect -6278 423418 -6096 423654
rect -6696 423334 -6096 423418
rect -6696 423098 -6514 423334
rect -6278 423098 -6096 423334
rect -6696 387654 -6096 423098
rect -6696 387418 -6514 387654
rect -6278 387418 -6096 387654
rect -6696 387334 -6096 387418
rect -6696 387098 -6514 387334
rect -6278 387098 -6096 387334
rect -6696 351654 -6096 387098
rect -6696 351418 -6514 351654
rect -6278 351418 -6096 351654
rect -6696 351334 -6096 351418
rect -6696 351098 -6514 351334
rect -6278 351098 -6096 351334
rect -6696 315654 -6096 351098
rect -6696 315418 -6514 315654
rect -6278 315418 -6096 315654
rect -6696 315334 -6096 315418
rect -6696 315098 -6514 315334
rect -6278 315098 -6096 315334
rect -6696 279654 -6096 315098
rect -6696 279418 -6514 279654
rect -6278 279418 -6096 279654
rect -6696 279334 -6096 279418
rect -6696 279098 -6514 279334
rect -6278 279098 -6096 279334
rect -6696 243654 -6096 279098
rect -6696 243418 -6514 243654
rect -6278 243418 -6096 243654
rect -6696 243334 -6096 243418
rect -6696 243098 -6514 243334
rect -6278 243098 -6096 243334
rect -6696 207654 -6096 243098
rect -6696 207418 -6514 207654
rect -6278 207418 -6096 207654
rect -6696 207334 -6096 207418
rect -6696 207098 -6514 207334
rect -6278 207098 -6096 207334
rect -6696 171654 -6096 207098
rect -6696 171418 -6514 171654
rect -6278 171418 -6096 171654
rect -6696 171334 -6096 171418
rect -6696 171098 -6514 171334
rect -6278 171098 -6096 171334
rect -6696 135654 -6096 171098
rect -6696 135418 -6514 135654
rect -6278 135418 -6096 135654
rect -6696 135334 -6096 135418
rect -6696 135098 -6514 135334
rect -6278 135098 -6096 135334
rect -6696 99654 -6096 135098
rect -6696 99418 -6514 99654
rect -6278 99418 -6096 99654
rect -6696 99334 -6096 99418
rect -6696 99098 -6514 99334
rect -6278 99098 -6096 99334
rect -6696 63654 -6096 99098
rect -6696 63418 -6514 63654
rect -6278 63418 -6096 63654
rect -6696 63334 -6096 63418
rect -6696 63098 -6514 63334
rect -6278 63098 -6096 63334
rect -6696 27654 -6096 63098
rect -6696 27418 -6514 27654
rect -6278 27418 -6096 27654
rect -6696 27334 -6096 27418
rect -6696 27098 -6514 27334
rect -6278 27098 -6096 27334
rect -6696 -5046 -6096 27098
rect -5756 708598 -5156 708620
rect -5756 708362 -5574 708598
rect -5338 708362 -5156 708598
rect -5756 708278 -5156 708362
rect -5756 708042 -5574 708278
rect -5338 708042 -5156 708278
rect -5756 693654 -5156 708042
rect 8004 708598 8604 709560
rect 8004 708362 8186 708598
rect 8422 708362 8604 708598
rect 8004 708278 8604 708362
rect 8004 708042 8186 708278
rect 8422 708042 8604 708278
rect -5756 693418 -5574 693654
rect -5338 693418 -5156 693654
rect -5756 693334 -5156 693418
rect -5756 693098 -5574 693334
rect -5338 693098 -5156 693334
rect -5756 657654 -5156 693098
rect -5756 657418 -5574 657654
rect -5338 657418 -5156 657654
rect -5756 657334 -5156 657418
rect -5756 657098 -5574 657334
rect -5338 657098 -5156 657334
rect -5756 621654 -5156 657098
rect -5756 621418 -5574 621654
rect -5338 621418 -5156 621654
rect -5756 621334 -5156 621418
rect -5756 621098 -5574 621334
rect -5338 621098 -5156 621334
rect -5756 585654 -5156 621098
rect -5756 585418 -5574 585654
rect -5338 585418 -5156 585654
rect -5756 585334 -5156 585418
rect -5756 585098 -5574 585334
rect -5338 585098 -5156 585334
rect -5756 549654 -5156 585098
rect -5756 549418 -5574 549654
rect -5338 549418 -5156 549654
rect -5756 549334 -5156 549418
rect -5756 549098 -5574 549334
rect -5338 549098 -5156 549334
rect -5756 513654 -5156 549098
rect -5756 513418 -5574 513654
rect -5338 513418 -5156 513654
rect -5756 513334 -5156 513418
rect -5756 513098 -5574 513334
rect -5338 513098 -5156 513334
rect -5756 477654 -5156 513098
rect -5756 477418 -5574 477654
rect -5338 477418 -5156 477654
rect -5756 477334 -5156 477418
rect -5756 477098 -5574 477334
rect -5338 477098 -5156 477334
rect -5756 441654 -5156 477098
rect -5756 441418 -5574 441654
rect -5338 441418 -5156 441654
rect -5756 441334 -5156 441418
rect -5756 441098 -5574 441334
rect -5338 441098 -5156 441334
rect -5756 405654 -5156 441098
rect -5756 405418 -5574 405654
rect -5338 405418 -5156 405654
rect -5756 405334 -5156 405418
rect -5756 405098 -5574 405334
rect -5338 405098 -5156 405334
rect -5756 369654 -5156 405098
rect -5756 369418 -5574 369654
rect -5338 369418 -5156 369654
rect -5756 369334 -5156 369418
rect -5756 369098 -5574 369334
rect -5338 369098 -5156 369334
rect -5756 333654 -5156 369098
rect -5756 333418 -5574 333654
rect -5338 333418 -5156 333654
rect -5756 333334 -5156 333418
rect -5756 333098 -5574 333334
rect -5338 333098 -5156 333334
rect -5756 297654 -5156 333098
rect -5756 297418 -5574 297654
rect -5338 297418 -5156 297654
rect -5756 297334 -5156 297418
rect -5756 297098 -5574 297334
rect -5338 297098 -5156 297334
rect -5756 261654 -5156 297098
rect -5756 261418 -5574 261654
rect -5338 261418 -5156 261654
rect -5756 261334 -5156 261418
rect -5756 261098 -5574 261334
rect -5338 261098 -5156 261334
rect -5756 225654 -5156 261098
rect -5756 225418 -5574 225654
rect -5338 225418 -5156 225654
rect -5756 225334 -5156 225418
rect -5756 225098 -5574 225334
rect -5338 225098 -5156 225334
rect -5756 189654 -5156 225098
rect -5756 189418 -5574 189654
rect -5338 189418 -5156 189654
rect -5756 189334 -5156 189418
rect -5756 189098 -5574 189334
rect -5338 189098 -5156 189334
rect -5756 153654 -5156 189098
rect -5756 153418 -5574 153654
rect -5338 153418 -5156 153654
rect -5756 153334 -5156 153418
rect -5756 153098 -5574 153334
rect -5338 153098 -5156 153334
rect -5756 117654 -5156 153098
rect -5756 117418 -5574 117654
rect -5338 117418 -5156 117654
rect -5756 117334 -5156 117418
rect -5756 117098 -5574 117334
rect -5338 117098 -5156 117334
rect -5756 81654 -5156 117098
rect -5756 81418 -5574 81654
rect -5338 81418 -5156 81654
rect -5756 81334 -5156 81418
rect -5756 81098 -5574 81334
rect -5338 81098 -5156 81334
rect -5756 45654 -5156 81098
rect -5756 45418 -5574 45654
rect -5338 45418 -5156 45654
rect -5756 45334 -5156 45418
rect -5756 45098 -5574 45334
rect -5338 45098 -5156 45334
rect -5756 9654 -5156 45098
rect -5756 9418 -5574 9654
rect -5338 9418 -5156 9654
rect -5756 9334 -5156 9418
rect -5756 9098 -5574 9334
rect -5338 9098 -5156 9334
rect -5756 -4106 -5156 9098
rect -4816 707658 -4216 707680
rect -4816 707422 -4634 707658
rect -4398 707422 -4216 707658
rect -4816 707338 -4216 707422
rect -4816 707102 -4634 707338
rect -4398 707102 -4216 707338
rect -4816 672054 -4216 707102
rect -4816 671818 -4634 672054
rect -4398 671818 -4216 672054
rect -4816 671734 -4216 671818
rect -4816 671498 -4634 671734
rect -4398 671498 -4216 671734
rect -4816 636054 -4216 671498
rect -4816 635818 -4634 636054
rect -4398 635818 -4216 636054
rect -4816 635734 -4216 635818
rect -4816 635498 -4634 635734
rect -4398 635498 -4216 635734
rect -4816 600054 -4216 635498
rect -4816 599818 -4634 600054
rect -4398 599818 -4216 600054
rect -4816 599734 -4216 599818
rect -4816 599498 -4634 599734
rect -4398 599498 -4216 599734
rect -4816 564054 -4216 599498
rect -4816 563818 -4634 564054
rect -4398 563818 -4216 564054
rect -4816 563734 -4216 563818
rect -4816 563498 -4634 563734
rect -4398 563498 -4216 563734
rect -4816 528054 -4216 563498
rect -4816 527818 -4634 528054
rect -4398 527818 -4216 528054
rect -4816 527734 -4216 527818
rect -4816 527498 -4634 527734
rect -4398 527498 -4216 527734
rect -4816 492054 -4216 527498
rect -4816 491818 -4634 492054
rect -4398 491818 -4216 492054
rect -4816 491734 -4216 491818
rect -4816 491498 -4634 491734
rect -4398 491498 -4216 491734
rect -4816 456054 -4216 491498
rect -4816 455818 -4634 456054
rect -4398 455818 -4216 456054
rect -4816 455734 -4216 455818
rect -4816 455498 -4634 455734
rect -4398 455498 -4216 455734
rect -4816 420054 -4216 455498
rect -4816 419818 -4634 420054
rect -4398 419818 -4216 420054
rect -4816 419734 -4216 419818
rect -4816 419498 -4634 419734
rect -4398 419498 -4216 419734
rect -4816 384054 -4216 419498
rect -4816 383818 -4634 384054
rect -4398 383818 -4216 384054
rect -4816 383734 -4216 383818
rect -4816 383498 -4634 383734
rect -4398 383498 -4216 383734
rect -4816 348054 -4216 383498
rect -4816 347818 -4634 348054
rect -4398 347818 -4216 348054
rect -4816 347734 -4216 347818
rect -4816 347498 -4634 347734
rect -4398 347498 -4216 347734
rect -4816 312054 -4216 347498
rect -4816 311818 -4634 312054
rect -4398 311818 -4216 312054
rect -4816 311734 -4216 311818
rect -4816 311498 -4634 311734
rect -4398 311498 -4216 311734
rect -4816 276054 -4216 311498
rect -4816 275818 -4634 276054
rect -4398 275818 -4216 276054
rect -4816 275734 -4216 275818
rect -4816 275498 -4634 275734
rect -4398 275498 -4216 275734
rect -4816 240054 -4216 275498
rect -4816 239818 -4634 240054
rect -4398 239818 -4216 240054
rect -4816 239734 -4216 239818
rect -4816 239498 -4634 239734
rect -4398 239498 -4216 239734
rect -4816 204054 -4216 239498
rect -4816 203818 -4634 204054
rect -4398 203818 -4216 204054
rect -4816 203734 -4216 203818
rect -4816 203498 -4634 203734
rect -4398 203498 -4216 203734
rect -4816 168054 -4216 203498
rect -4816 167818 -4634 168054
rect -4398 167818 -4216 168054
rect -4816 167734 -4216 167818
rect -4816 167498 -4634 167734
rect -4398 167498 -4216 167734
rect -4816 132054 -4216 167498
rect -4816 131818 -4634 132054
rect -4398 131818 -4216 132054
rect -4816 131734 -4216 131818
rect -4816 131498 -4634 131734
rect -4398 131498 -4216 131734
rect -4816 96054 -4216 131498
rect -4816 95818 -4634 96054
rect -4398 95818 -4216 96054
rect -4816 95734 -4216 95818
rect -4816 95498 -4634 95734
rect -4398 95498 -4216 95734
rect -4816 60054 -4216 95498
rect -4816 59818 -4634 60054
rect -4398 59818 -4216 60054
rect -4816 59734 -4216 59818
rect -4816 59498 -4634 59734
rect -4398 59498 -4216 59734
rect -4816 24054 -4216 59498
rect -4816 23818 -4634 24054
rect -4398 23818 -4216 24054
rect -4816 23734 -4216 23818
rect -4816 23498 -4634 23734
rect -4398 23498 -4216 23734
rect -4816 -3166 -4216 23498
rect -3876 706718 -3276 706740
rect -3876 706482 -3694 706718
rect -3458 706482 -3276 706718
rect -3876 706398 -3276 706482
rect -3876 706162 -3694 706398
rect -3458 706162 -3276 706398
rect -3876 690054 -3276 706162
rect 4404 706718 5004 707680
rect 4404 706482 4586 706718
rect 4822 706482 5004 706718
rect 4404 706398 5004 706482
rect 4404 706162 4586 706398
rect 4822 706162 5004 706398
rect -3876 689818 -3694 690054
rect -3458 689818 -3276 690054
rect -3876 689734 -3276 689818
rect -3876 689498 -3694 689734
rect -3458 689498 -3276 689734
rect -3876 654054 -3276 689498
rect -3876 653818 -3694 654054
rect -3458 653818 -3276 654054
rect -3876 653734 -3276 653818
rect -3876 653498 -3694 653734
rect -3458 653498 -3276 653734
rect -3876 618054 -3276 653498
rect -3876 617818 -3694 618054
rect -3458 617818 -3276 618054
rect -3876 617734 -3276 617818
rect -3876 617498 -3694 617734
rect -3458 617498 -3276 617734
rect -3876 582054 -3276 617498
rect -3876 581818 -3694 582054
rect -3458 581818 -3276 582054
rect -3876 581734 -3276 581818
rect -3876 581498 -3694 581734
rect -3458 581498 -3276 581734
rect -3876 546054 -3276 581498
rect -3876 545818 -3694 546054
rect -3458 545818 -3276 546054
rect -3876 545734 -3276 545818
rect -3876 545498 -3694 545734
rect -3458 545498 -3276 545734
rect -3876 510054 -3276 545498
rect -3876 509818 -3694 510054
rect -3458 509818 -3276 510054
rect -3876 509734 -3276 509818
rect -3876 509498 -3694 509734
rect -3458 509498 -3276 509734
rect -3876 474054 -3276 509498
rect -3876 473818 -3694 474054
rect -3458 473818 -3276 474054
rect -3876 473734 -3276 473818
rect -3876 473498 -3694 473734
rect -3458 473498 -3276 473734
rect -3876 438054 -3276 473498
rect -3876 437818 -3694 438054
rect -3458 437818 -3276 438054
rect -3876 437734 -3276 437818
rect -3876 437498 -3694 437734
rect -3458 437498 -3276 437734
rect -3876 402054 -3276 437498
rect -3876 401818 -3694 402054
rect -3458 401818 -3276 402054
rect -3876 401734 -3276 401818
rect -3876 401498 -3694 401734
rect -3458 401498 -3276 401734
rect -3876 366054 -3276 401498
rect -3876 365818 -3694 366054
rect -3458 365818 -3276 366054
rect -3876 365734 -3276 365818
rect -3876 365498 -3694 365734
rect -3458 365498 -3276 365734
rect -3876 330054 -3276 365498
rect -3876 329818 -3694 330054
rect -3458 329818 -3276 330054
rect -3876 329734 -3276 329818
rect -3876 329498 -3694 329734
rect -3458 329498 -3276 329734
rect -3876 294054 -3276 329498
rect -3876 293818 -3694 294054
rect -3458 293818 -3276 294054
rect -3876 293734 -3276 293818
rect -3876 293498 -3694 293734
rect -3458 293498 -3276 293734
rect -3876 258054 -3276 293498
rect -3876 257818 -3694 258054
rect -3458 257818 -3276 258054
rect -3876 257734 -3276 257818
rect -3876 257498 -3694 257734
rect -3458 257498 -3276 257734
rect -3876 222054 -3276 257498
rect -3876 221818 -3694 222054
rect -3458 221818 -3276 222054
rect -3876 221734 -3276 221818
rect -3876 221498 -3694 221734
rect -3458 221498 -3276 221734
rect -3876 186054 -3276 221498
rect -3876 185818 -3694 186054
rect -3458 185818 -3276 186054
rect -3876 185734 -3276 185818
rect -3876 185498 -3694 185734
rect -3458 185498 -3276 185734
rect -3876 150054 -3276 185498
rect -3876 149818 -3694 150054
rect -3458 149818 -3276 150054
rect -3876 149734 -3276 149818
rect -3876 149498 -3694 149734
rect -3458 149498 -3276 149734
rect -3876 114054 -3276 149498
rect -3876 113818 -3694 114054
rect -3458 113818 -3276 114054
rect -3876 113734 -3276 113818
rect -3876 113498 -3694 113734
rect -3458 113498 -3276 113734
rect -3876 78054 -3276 113498
rect -3876 77818 -3694 78054
rect -3458 77818 -3276 78054
rect -3876 77734 -3276 77818
rect -3876 77498 -3694 77734
rect -3458 77498 -3276 77734
rect -3876 42054 -3276 77498
rect -3876 41818 -3694 42054
rect -3458 41818 -3276 42054
rect -3876 41734 -3276 41818
rect -3876 41498 -3694 41734
rect -3458 41498 -3276 41734
rect -3876 6054 -3276 41498
rect -3876 5818 -3694 6054
rect -3458 5818 -3276 6054
rect -3876 5734 -3276 5818
rect -3876 5498 -3694 5734
rect -3458 5498 -3276 5734
rect -3876 -2226 -3276 5498
rect -2936 705778 -2336 705800
rect -2936 705542 -2754 705778
rect -2518 705542 -2336 705778
rect -2936 705458 -2336 705542
rect -2936 705222 -2754 705458
rect -2518 705222 -2336 705458
rect -2936 668454 -2336 705222
rect -2936 668218 -2754 668454
rect -2518 668218 -2336 668454
rect -2936 668134 -2336 668218
rect -2936 667898 -2754 668134
rect -2518 667898 -2336 668134
rect -2936 632454 -2336 667898
rect -2936 632218 -2754 632454
rect -2518 632218 -2336 632454
rect -2936 632134 -2336 632218
rect -2936 631898 -2754 632134
rect -2518 631898 -2336 632134
rect -2936 596454 -2336 631898
rect -2936 596218 -2754 596454
rect -2518 596218 -2336 596454
rect -2936 596134 -2336 596218
rect -2936 595898 -2754 596134
rect -2518 595898 -2336 596134
rect -2936 560454 -2336 595898
rect -2936 560218 -2754 560454
rect -2518 560218 -2336 560454
rect -2936 560134 -2336 560218
rect -2936 559898 -2754 560134
rect -2518 559898 -2336 560134
rect -2936 524454 -2336 559898
rect -2936 524218 -2754 524454
rect -2518 524218 -2336 524454
rect -2936 524134 -2336 524218
rect -2936 523898 -2754 524134
rect -2518 523898 -2336 524134
rect -2936 488454 -2336 523898
rect -2936 488218 -2754 488454
rect -2518 488218 -2336 488454
rect -2936 488134 -2336 488218
rect -2936 487898 -2754 488134
rect -2518 487898 -2336 488134
rect -2936 452454 -2336 487898
rect -2936 452218 -2754 452454
rect -2518 452218 -2336 452454
rect -2936 452134 -2336 452218
rect -2936 451898 -2754 452134
rect -2518 451898 -2336 452134
rect -2936 416454 -2336 451898
rect -2936 416218 -2754 416454
rect -2518 416218 -2336 416454
rect -2936 416134 -2336 416218
rect -2936 415898 -2754 416134
rect -2518 415898 -2336 416134
rect -2936 380454 -2336 415898
rect -2936 380218 -2754 380454
rect -2518 380218 -2336 380454
rect -2936 380134 -2336 380218
rect -2936 379898 -2754 380134
rect -2518 379898 -2336 380134
rect -2936 344454 -2336 379898
rect -2936 344218 -2754 344454
rect -2518 344218 -2336 344454
rect -2936 344134 -2336 344218
rect -2936 343898 -2754 344134
rect -2518 343898 -2336 344134
rect -2936 308454 -2336 343898
rect -2936 308218 -2754 308454
rect -2518 308218 -2336 308454
rect -2936 308134 -2336 308218
rect -2936 307898 -2754 308134
rect -2518 307898 -2336 308134
rect -2936 272454 -2336 307898
rect -2936 272218 -2754 272454
rect -2518 272218 -2336 272454
rect -2936 272134 -2336 272218
rect -2936 271898 -2754 272134
rect -2518 271898 -2336 272134
rect -2936 236454 -2336 271898
rect -2936 236218 -2754 236454
rect -2518 236218 -2336 236454
rect -2936 236134 -2336 236218
rect -2936 235898 -2754 236134
rect -2518 235898 -2336 236134
rect -2936 200454 -2336 235898
rect -2936 200218 -2754 200454
rect -2518 200218 -2336 200454
rect -2936 200134 -2336 200218
rect -2936 199898 -2754 200134
rect -2518 199898 -2336 200134
rect -2936 164454 -2336 199898
rect -2936 164218 -2754 164454
rect -2518 164218 -2336 164454
rect -2936 164134 -2336 164218
rect -2936 163898 -2754 164134
rect -2518 163898 -2336 164134
rect -2936 128454 -2336 163898
rect -2936 128218 -2754 128454
rect -2518 128218 -2336 128454
rect -2936 128134 -2336 128218
rect -2936 127898 -2754 128134
rect -2518 127898 -2336 128134
rect -2936 92454 -2336 127898
rect -2936 92218 -2754 92454
rect -2518 92218 -2336 92454
rect -2936 92134 -2336 92218
rect -2936 91898 -2754 92134
rect -2518 91898 -2336 92134
rect -2936 56454 -2336 91898
rect -2936 56218 -2754 56454
rect -2518 56218 -2336 56454
rect -2936 56134 -2336 56218
rect -2936 55898 -2754 56134
rect -2518 55898 -2336 56134
rect -2936 20454 -2336 55898
rect -2936 20218 -2754 20454
rect -2518 20218 -2336 20454
rect -2936 20134 -2336 20218
rect -2936 19898 -2754 20134
rect -2518 19898 -2336 20134
rect -2936 -1286 -2336 19898
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 686454 -1396 704282
rect -1996 686218 -1814 686454
rect -1578 686218 -1396 686454
rect -1996 686134 -1396 686218
rect -1996 685898 -1814 686134
rect -1578 685898 -1396 686134
rect -1996 650454 -1396 685898
rect -1996 650218 -1814 650454
rect -1578 650218 -1396 650454
rect -1996 650134 -1396 650218
rect -1996 649898 -1814 650134
rect -1578 649898 -1396 650134
rect -1996 614454 -1396 649898
rect -1996 614218 -1814 614454
rect -1578 614218 -1396 614454
rect -1996 614134 -1396 614218
rect -1996 613898 -1814 614134
rect -1578 613898 -1396 614134
rect -1996 578454 -1396 613898
rect -1996 578218 -1814 578454
rect -1578 578218 -1396 578454
rect -1996 578134 -1396 578218
rect -1996 577898 -1814 578134
rect -1578 577898 -1396 578134
rect -1996 542454 -1396 577898
rect -1996 542218 -1814 542454
rect -1578 542218 -1396 542454
rect -1996 542134 -1396 542218
rect -1996 541898 -1814 542134
rect -1578 541898 -1396 542134
rect -1996 506454 -1396 541898
rect -1996 506218 -1814 506454
rect -1578 506218 -1396 506454
rect -1996 506134 -1396 506218
rect -1996 505898 -1814 506134
rect -1578 505898 -1396 506134
rect -1996 470454 -1396 505898
rect -1996 470218 -1814 470454
rect -1578 470218 -1396 470454
rect -1996 470134 -1396 470218
rect -1996 469898 -1814 470134
rect -1578 469898 -1396 470134
rect -1996 434454 -1396 469898
rect -1996 434218 -1814 434454
rect -1578 434218 -1396 434454
rect -1996 434134 -1396 434218
rect -1996 433898 -1814 434134
rect -1578 433898 -1396 434134
rect -1996 398454 -1396 433898
rect -1996 398218 -1814 398454
rect -1578 398218 -1396 398454
rect -1996 398134 -1396 398218
rect -1996 397898 -1814 398134
rect -1578 397898 -1396 398134
rect -1996 362454 -1396 397898
rect -1996 362218 -1814 362454
rect -1578 362218 -1396 362454
rect -1996 362134 -1396 362218
rect -1996 361898 -1814 362134
rect -1578 361898 -1396 362134
rect -1996 326454 -1396 361898
rect -1996 326218 -1814 326454
rect -1578 326218 -1396 326454
rect -1996 326134 -1396 326218
rect -1996 325898 -1814 326134
rect -1578 325898 -1396 326134
rect -1996 290454 -1396 325898
rect -1996 290218 -1814 290454
rect -1578 290218 -1396 290454
rect -1996 290134 -1396 290218
rect -1996 289898 -1814 290134
rect -1578 289898 -1396 290134
rect -1996 254454 -1396 289898
rect -1996 254218 -1814 254454
rect -1578 254218 -1396 254454
rect -1996 254134 -1396 254218
rect -1996 253898 -1814 254134
rect -1578 253898 -1396 254134
rect -1996 218454 -1396 253898
rect -1996 218218 -1814 218454
rect -1578 218218 -1396 218454
rect -1996 218134 -1396 218218
rect -1996 217898 -1814 218134
rect -1578 217898 -1396 218134
rect -1996 182454 -1396 217898
rect -1996 182218 -1814 182454
rect -1578 182218 -1396 182454
rect -1996 182134 -1396 182218
rect -1996 181898 -1814 182134
rect -1578 181898 -1396 182134
rect -1996 146454 -1396 181898
rect -1996 146218 -1814 146454
rect -1578 146218 -1396 146454
rect -1996 146134 -1396 146218
rect -1996 145898 -1814 146134
rect -1578 145898 -1396 146134
rect -1996 110454 -1396 145898
rect -1996 110218 -1814 110454
rect -1578 110218 -1396 110454
rect -1996 110134 -1396 110218
rect -1996 109898 -1814 110134
rect -1578 109898 -1396 110134
rect -1996 74454 -1396 109898
rect -1996 74218 -1814 74454
rect -1578 74218 -1396 74454
rect -1996 74134 -1396 74218
rect -1996 73898 -1814 74134
rect -1578 73898 -1396 74134
rect -1996 38454 -1396 73898
rect -1996 38218 -1814 38454
rect -1578 38218 -1396 38454
rect -1996 38134 -1396 38218
rect -1996 37898 -1814 38134
rect -1578 37898 -1396 38134
rect -1996 2454 -1396 37898
rect -1996 2218 -1814 2454
rect -1578 2218 -1396 2454
rect -1996 2134 -1396 2218
rect -1996 1898 -1814 2134
rect -1578 1898 -1396 2134
rect -1996 -346 -1396 1898
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 804 704838 1404 705800
rect 804 704602 986 704838
rect 1222 704602 1404 704838
rect 804 704518 1404 704602
rect 804 704282 986 704518
rect 1222 704282 1404 704518
rect 804 686454 1404 704282
rect 804 686218 986 686454
rect 1222 686218 1404 686454
rect 804 686134 1404 686218
rect 804 685898 986 686134
rect 1222 685898 1404 686134
rect 804 650454 1404 685898
rect 804 650218 986 650454
rect 1222 650218 1404 650454
rect 804 650134 1404 650218
rect 804 649898 986 650134
rect 1222 649898 1404 650134
rect 804 614454 1404 649898
rect 804 614218 986 614454
rect 1222 614218 1404 614454
rect 804 614134 1404 614218
rect 804 613898 986 614134
rect 1222 613898 1404 614134
rect 804 578454 1404 613898
rect 804 578218 986 578454
rect 1222 578218 1404 578454
rect 804 578134 1404 578218
rect 804 577898 986 578134
rect 1222 577898 1404 578134
rect 804 542454 1404 577898
rect 804 542218 986 542454
rect 1222 542218 1404 542454
rect 804 542134 1404 542218
rect 804 541898 986 542134
rect 1222 541898 1404 542134
rect 804 506454 1404 541898
rect 804 506218 986 506454
rect 1222 506218 1404 506454
rect 804 506134 1404 506218
rect 804 505898 986 506134
rect 1222 505898 1404 506134
rect 804 470454 1404 505898
rect 804 470218 986 470454
rect 1222 470218 1404 470454
rect 804 470134 1404 470218
rect 804 469898 986 470134
rect 1222 469898 1404 470134
rect 804 434454 1404 469898
rect 804 434218 986 434454
rect 1222 434218 1404 434454
rect 804 434134 1404 434218
rect 804 433898 986 434134
rect 1222 433898 1404 434134
rect 804 398454 1404 433898
rect 804 398218 986 398454
rect 1222 398218 1404 398454
rect 804 398134 1404 398218
rect 804 397898 986 398134
rect 1222 397898 1404 398134
rect 804 362454 1404 397898
rect 804 362218 986 362454
rect 1222 362218 1404 362454
rect 804 362134 1404 362218
rect 804 361898 986 362134
rect 1222 361898 1404 362134
rect 804 326454 1404 361898
rect 804 326218 986 326454
rect 1222 326218 1404 326454
rect 804 326134 1404 326218
rect 804 325898 986 326134
rect 1222 325898 1404 326134
rect 804 290454 1404 325898
rect 804 290218 986 290454
rect 1222 290218 1404 290454
rect 804 290134 1404 290218
rect 804 289898 986 290134
rect 1222 289898 1404 290134
rect 804 254454 1404 289898
rect 804 254218 986 254454
rect 1222 254218 1404 254454
rect 804 254134 1404 254218
rect 804 253898 986 254134
rect 1222 253898 1404 254134
rect 804 218454 1404 253898
rect 804 218218 986 218454
rect 1222 218218 1404 218454
rect 804 218134 1404 218218
rect 804 217898 986 218134
rect 1222 217898 1404 218134
rect 804 182454 1404 217898
rect 804 182218 986 182454
rect 1222 182218 1404 182454
rect 804 182134 1404 182218
rect 804 181898 986 182134
rect 1222 181898 1404 182134
rect 804 146454 1404 181898
rect 804 146218 986 146454
rect 1222 146218 1404 146454
rect 804 146134 1404 146218
rect 804 145898 986 146134
rect 1222 145898 1404 146134
rect 804 110454 1404 145898
rect 804 110218 986 110454
rect 1222 110218 1404 110454
rect 804 110134 1404 110218
rect 804 109898 986 110134
rect 1222 109898 1404 110134
rect 804 74454 1404 109898
rect 804 74218 986 74454
rect 1222 74218 1404 74454
rect 804 74134 1404 74218
rect 804 73898 986 74134
rect 1222 73898 1404 74134
rect 804 38454 1404 73898
rect 804 38218 986 38454
rect 1222 38218 1404 38454
rect 804 38134 1404 38218
rect 804 37898 986 38134
rect 1222 37898 1404 38134
rect 804 2454 1404 37898
rect 804 2218 986 2454
rect 1222 2218 1404 2454
rect 804 2134 1404 2218
rect 804 1898 986 2134
rect 1222 1898 1404 2134
rect 804 -346 1404 1898
rect 804 -582 986 -346
rect 1222 -582 1404 -346
rect 804 -666 1404 -582
rect 804 -902 986 -666
rect 1222 -902 1404 -666
rect -2936 -1522 -2754 -1286
rect -2518 -1522 -2336 -1286
rect -2936 -1606 -2336 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 -2336 -1606
rect -2936 -1864 -2336 -1842
rect 804 -1864 1404 -902
rect 4404 690054 5004 706162
rect 4404 689818 4586 690054
rect 4822 689818 5004 690054
rect 4404 689734 5004 689818
rect 4404 689498 4586 689734
rect 4822 689498 5004 689734
rect 4404 654054 5004 689498
rect 4404 653818 4586 654054
rect 4822 653818 5004 654054
rect 4404 653734 5004 653818
rect 4404 653498 4586 653734
rect 4822 653498 5004 653734
rect 4404 618054 5004 653498
rect 4404 617818 4586 618054
rect 4822 617818 5004 618054
rect 4404 617734 5004 617818
rect 4404 617498 4586 617734
rect 4822 617498 5004 617734
rect 4404 582054 5004 617498
rect 4404 581818 4586 582054
rect 4822 581818 5004 582054
rect 4404 581734 5004 581818
rect 4404 581498 4586 581734
rect 4822 581498 5004 581734
rect 4404 546054 5004 581498
rect 4404 545818 4586 546054
rect 4822 545818 5004 546054
rect 4404 545734 5004 545818
rect 4404 545498 4586 545734
rect 4822 545498 5004 545734
rect 4404 510054 5004 545498
rect 4404 509818 4586 510054
rect 4822 509818 5004 510054
rect 4404 509734 5004 509818
rect 4404 509498 4586 509734
rect 4822 509498 5004 509734
rect 4404 474054 5004 509498
rect 4404 473818 4586 474054
rect 4822 473818 5004 474054
rect 4404 473734 5004 473818
rect 4404 473498 4586 473734
rect 4822 473498 5004 473734
rect 4404 438054 5004 473498
rect 4404 437818 4586 438054
rect 4822 437818 5004 438054
rect 4404 437734 5004 437818
rect 4404 437498 4586 437734
rect 4822 437498 5004 437734
rect 4404 402054 5004 437498
rect 4404 401818 4586 402054
rect 4822 401818 5004 402054
rect 4404 401734 5004 401818
rect 4404 401498 4586 401734
rect 4822 401498 5004 401734
rect 4404 366054 5004 401498
rect 4404 365818 4586 366054
rect 4822 365818 5004 366054
rect 4404 365734 5004 365818
rect 4404 365498 4586 365734
rect 4822 365498 5004 365734
rect 4404 330054 5004 365498
rect 4404 329818 4586 330054
rect 4822 329818 5004 330054
rect 4404 329734 5004 329818
rect 4404 329498 4586 329734
rect 4822 329498 5004 329734
rect 4404 294054 5004 329498
rect 4404 293818 4586 294054
rect 4822 293818 5004 294054
rect 4404 293734 5004 293818
rect 4404 293498 4586 293734
rect 4822 293498 5004 293734
rect 4404 258054 5004 293498
rect 4404 257818 4586 258054
rect 4822 257818 5004 258054
rect 4404 257734 5004 257818
rect 4404 257498 4586 257734
rect 4822 257498 5004 257734
rect 4404 222054 5004 257498
rect 4404 221818 4586 222054
rect 4822 221818 5004 222054
rect 4404 221734 5004 221818
rect 4404 221498 4586 221734
rect 4822 221498 5004 221734
rect 4404 186054 5004 221498
rect 4404 185818 4586 186054
rect 4822 185818 5004 186054
rect 4404 185734 5004 185818
rect 4404 185498 4586 185734
rect 4822 185498 5004 185734
rect 4404 150054 5004 185498
rect 4404 149818 4586 150054
rect 4822 149818 5004 150054
rect 4404 149734 5004 149818
rect 4404 149498 4586 149734
rect 4822 149498 5004 149734
rect 4404 114054 5004 149498
rect 4404 113818 4586 114054
rect 4822 113818 5004 114054
rect 4404 113734 5004 113818
rect 4404 113498 4586 113734
rect 4822 113498 5004 113734
rect 4404 78054 5004 113498
rect 4404 77818 4586 78054
rect 4822 77818 5004 78054
rect 4404 77734 5004 77818
rect 4404 77498 4586 77734
rect 4822 77498 5004 77734
rect 4404 42054 5004 77498
rect 4404 41818 4586 42054
rect 4822 41818 5004 42054
rect 4404 41734 5004 41818
rect 4404 41498 4586 41734
rect 4822 41498 5004 41734
rect 4404 6054 5004 41498
rect 4404 5818 4586 6054
rect 4822 5818 5004 6054
rect 4404 5734 5004 5818
rect 4404 5498 4586 5734
rect 4822 5498 5004 5734
rect -3876 -2462 -3694 -2226
rect -3458 -2462 -3276 -2226
rect -3876 -2546 -3276 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 -3276 -2546
rect -3876 -2804 -3276 -2782
rect 4404 -2226 5004 5498
rect 4404 -2462 4586 -2226
rect 4822 -2462 5004 -2226
rect 4404 -2546 5004 -2462
rect 4404 -2782 4586 -2546
rect 4822 -2782 5004 -2546
rect -4816 -3402 -4634 -3166
rect -4398 -3402 -4216 -3166
rect -4816 -3486 -4216 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 -4216 -3486
rect -4816 -3744 -4216 -3722
rect 4404 -3744 5004 -2782
rect 8004 693654 8604 708042
rect 8004 693418 8186 693654
rect 8422 693418 8604 693654
rect 8004 693334 8604 693418
rect 8004 693098 8186 693334
rect 8422 693098 8604 693334
rect 8004 657654 8604 693098
rect 8004 657418 8186 657654
rect 8422 657418 8604 657654
rect 8004 657334 8604 657418
rect 8004 657098 8186 657334
rect 8422 657098 8604 657334
rect 8004 621654 8604 657098
rect 8004 621418 8186 621654
rect 8422 621418 8604 621654
rect 8004 621334 8604 621418
rect 8004 621098 8186 621334
rect 8422 621098 8604 621334
rect 8004 585654 8604 621098
rect 8004 585418 8186 585654
rect 8422 585418 8604 585654
rect 8004 585334 8604 585418
rect 8004 585098 8186 585334
rect 8422 585098 8604 585334
rect 8004 549654 8604 585098
rect 8004 549418 8186 549654
rect 8422 549418 8604 549654
rect 8004 549334 8604 549418
rect 8004 549098 8186 549334
rect 8422 549098 8604 549334
rect 8004 513654 8604 549098
rect 8004 513418 8186 513654
rect 8422 513418 8604 513654
rect 8004 513334 8604 513418
rect 8004 513098 8186 513334
rect 8422 513098 8604 513334
rect 8004 477654 8604 513098
rect 8004 477418 8186 477654
rect 8422 477418 8604 477654
rect 8004 477334 8604 477418
rect 8004 477098 8186 477334
rect 8422 477098 8604 477334
rect 8004 441654 8604 477098
rect 8004 441418 8186 441654
rect 8422 441418 8604 441654
rect 8004 441334 8604 441418
rect 8004 441098 8186 441334
rect 8422 441098 8604 441334
rect 8004 405654 8604 441098
rect 8004 405418 8186 405654
rect 8422 405418 8604 405654
rect 8004 405334 8604 405418
rect 8004 405098 8186 405334
rect 8422 405098 8604 405334
rect 8004 369654 8604 405098
rect 8004 369418 8186 369654
rect 8422 369418 8604 369654
rect 8004 369334 8604 369418
rect 8004 369098 8186 369334
rect 8422 369098 8604 369334
rect 8004 333654 8604 369098
rect 8004 333418 8186 333654
rect 8422 333418 8604 333654
rect 8004 333334 8604 333418
rect 8004 333098 8186 333334
rect 8422 333098 8604 333334
rect 8004 297654 8604 333098
rect 8004 297418 8186 297654
rect 8422 297418 8604 297654
rect 8004 297334 8604 297418
rect 8004 297098 8186 297334
rect 8422 297098 8604 297334
rect 8004 261654 8604 297098
rect 8004 261418 8186 261654
rect 8422 261418 8604 261654
rect 8004 261334 8604 261418
rect 8004 261098 8186 261334
rect 8422 261098 8604 261334
rect 8004 225654 8604 261098
rect 8004 225418 8186 225654
rect 8422 225418 8604 225654
rect 8004 225334 8604 225418
rect 8004 225098 8186 225334
rect 8422 225098 8604 225334
rect 8004 189654 8604 225098
rect 8004 189418 8186 189654
rect 8422 189418 8604 189654
rect 8004 189334 8604 189418
rect 8004 189098 8186 189334
rect 8422 189098 8604 189334
rect 8004 153654 8604 189098
rect 8004 153418 8186 153654
rect 8422 153418 8604 153654
rect 8004 153334 8604 153418
rect 8004 153098 8186 153334
rect 8422 153098 8604 153334
rect 8004 117654 8604 153098
rect 8004 117418 8186 117654
rect 8422 117418 8604 117654
rect 8004 117334 8604 117418
rect 8004 117098 8186 117334
rect 8422 117098 8604 117334
rect 8004 81654 8604 117098
rect 8004 81418 8186 81654
rect 8422 81418 8604 81654
rect 8004 81334 8604 81418
rect 8004 81098 8186 81334
rect 8422 81098 8604 81334
rect 8004 45654 8604 81098
rect 8004 45418 8186 45654
rect 8422 45418 8604 45654
rect 8004 45334 8604 45418
rect 8004 45098 8186 45334
rect 8422 45098 8604 45334
rect 8004 9654 8604 45098
rect 8004 9418 8186 9654
rect 8422 9418 8604 9654
rect 8004 9334 8604 9418
rect 8004 9098 8186 9334
rect 8422 9098 8604 9334
rect -5756 -4342 -5574 -4106
rect -5338 -4342 -5156 -4106
rect -5756 -4426 -5156 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 -5156 -4426
rect -5756 -4684 -5156 -4662
rect 8004 -4106 8604 9098
rect 8004 -4342 8186 -4106
rect 8422 -4342 8604 -4106
rect 8004 -4426 8604 -4342
rect 8004 -4662 8186 -4426
rect 8422 -4662 8604 -4426
rect -6696 -5282 -6514 -5046
rect -6278 -5282 -6096 -5046
rect -6696 -5366 -6096 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 -6096 -5366
rect -6696 -5624 -6096 -5602
rect 8004 -5624 8604 -4662
rect 11604 697254 12204 709922
rect 29604 711418 30204 711440
rect 29604 711182 29786 711418
rect 30022 711182 30204 711418
rect 29604 711098 30204 711182
rect 29604 710862 29786 711098
rect 30022 710862 30204 711098
rect 26004 709538 26604 709560
rect 26004 709302 26186 709538
rect 26422 709302 26604 709538
rect 26004 709218 26604 709302
rect 26004 708982 26186 709218
rect 26422 708982 26604 709218
rect 22404 707658 23004 707680
rect 22404 707422 22586 707658
rect 22822 707422 23004 707658
rect 22404 707338 23004 707422
rect 22404 707102 22586 707338
rect 22822 707102 23004 707338
rect 11604 697018 11786 697254
rect 12022 697018 12204 697254
rect 11604 696934 12204 697018
rect 11604 696698 11786 696934
rect 12022 696698 12204 696934
rect 11604 661254 12204 696698
rect 11604 661018 11786 661254
rect 12022 661018 12204 661254
rect 11604 660934 12204 661018
rect 11604 660698 11786 660934
rect 12022 660698 12204 660934
rect 11604 625254 12204 660698
rect 11604 625018 11786 625254
rect 12022 625018 12204 625254
rect 11604 624934 12204 625018
rect 11604 624698 11786 624934
rect 12022 624698 12204 624934
rect 11604 589254 12204 624698
rect 11604 589018 11786 589254
rect 12022 589018 12204 589254
rect 11604 588934 12204 589018
rect 11604 588698 11786 588934
rect 12022 588698 12204 588934
rect 11604 553254 12204 588698
rect 11604 553018 11786 553254
rect 12022 553018 12204 553254
rect 11604 552934 12204 553018
rect 11604 552698 11786 552934
rect 12022 552698 12204 552934
rect 11604 517254 12204 552698
rect 11604 517018 11786 517254
rect 12022 517018 12204 517254
rect 11604 516934 12204 517018
rect 11604 516698 11786 516934
rect 12022 516698 12204 516934
rect 11604 481254 12204 516698
rect 11604 481018 11786 481254
rect 12022 481018 12204 481254
rect 11604 480934 12204 481018
rect 11604 480698 11786 480934
rect 12022 480698 12204 480934
rect 11604 445254 12204 480698
rect 11604 445018 11786 445254
rect 12022 445018 12204 445254
rect 11604 444934 12204 445018
rect 11604 444698 11786 444934
rect 12022 444698 12204 444934
rect 11604 409254 12204 444698
rect 11604 409018 11786 409254
rect 12022 409018 12204 409254
rect 11604 408934 12204 409018
rect 11604 408698 11786 408934
rect 12022 408698 12204 408934
rect 11604 373254 12204 408698
rect 11604 373018 11786 373254
rect 12022 373018 12204 373254
rect 11604 372934 12204 373018
rect 11604 372698 11786 372934
rect 12022 372698 12204 372934
rect 11604 337254 12204 372698
rect 11604 337018 11786 337254
rect 12022 337018 12204 337254
rect 11604 336934 12204 337018
rect 11604 336698 11786 336934
rect 12022 336698 12204 336934
rect 11604 301254 12204 336698
rect 11604 301018 11786 301254
rect 12022 301018 12204 301254
rect 11604 300934 12204 301018
rect 11604 300698 11786 300934
rect 12022 300698 12204 300934
rect 11604 265254 12204 300698
rect 11604 265018 11786 265254
rect 12022 265018 12204 265254
rect 11604 264934 12204 265018
rect 11604 264698 11786 264934
rect 12022 264698 12204 264934
rect 11604 229254 12204 264698
rect 11604 229018 11786 229254
rect 12022 229018 12204 229254
rect 11604 228934 12204 229018
rect 11604 228698 11786 228934
rect 12022 228698 12204 228934
rect 11604 193254 12204 228698
rect 11604 193018 11786 193254
rect 12022 193018 12204 193254
rect 11604 192934 12204 193018
rect 11604 192698 11786 192934
rect 12022 192698 12204 192934
rect 11604 157254 12204 192698
rect 11604 157018 11786 157254
rect 12022 157018 12204 157254
rect 11604 156934 12204 157018
rect 11604 156698 11786 156934
rect 12022 156698 12204 156934
rect 11604 121254 12204 156698
rect 11604 121018 11786 121254
rect 12022 121018 12204 121254
rect 11604 120934 12204 121018
rect 11604 120698 11786 120934
rect 12022 120698 12204 120934
rect 11604 85254 12204 120698
rect 11604 85018 11786 85254
rect 12022 85018 12204 85254
rect 11604 84934 12204 85018
rect 11604 84698 11786 84934
rect 12022 84698 12204 84934
rect 11604 49254 12204 84698
rect 11604 49018 11786 49254
rect 12022 49018 12204 49254
rect 11604 48934 12204 49018
rect 11604 48698 11786 48934
rect 12022 48698 12204 48934
rect 11604 13254 12204 48698
rect 11604 13018 11786 13254
rect 12022 13018 12204 13254
rect 11604 12934 12204 13018
rect 11604 12698 11786 12934
rect 12022 12698 12204 12934
rect -7636 -6222 -7454 -5986
rect -7218 -6222 -7036 -5986
rect -7636 -6306 -7036 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 -7036 -6306
rect -7636 -6564 -7036 -6542
rect 11604 -5986 12204 12698
rect 18804 705778 19404 705800
rect 18804 705542 18986 705778
rect 19222 705542 19404 705778
rect 18804 705458 19404 705542
rect 18804 705222 18986 705458
rect 19222 705222 19404 705458
rect 18804 668454 19404 705222
rect 18804 668218 18986 668454
rect 19222 668218 19404 668454
rect 18804 668134 19404 668218
rect 18804 667898 18986 668134
rect 19222 667898 19404 668134
rect 18804 632454 19404 667898
rect 18804 632218 18986 632454
rect 19222 632218 19404 632454
rect 18804 632134 19404 632218
rect 18804 631898 18986 632134
rect 19222 631898 19404 632134
rect 18804 596454 19404 631898
rect 18804 596218 18986 596454
rect 19222 596218 19404 596454
rect 18804 596134 19404 596218
rect 18804 595898 18986 596134
rect 19222 595898 19404 596134
rect 18804 560454 19404 595898
rect 18804 560218 18986 560454
rect 19222 560218 19404 560454
rect 18804 560134 19404 560218
rect 18804 559898 18986 560134
rect 19222 559898 19404 560134
rect 18804 524454 19404 559898
rect 18804 524218 18986 524454
rect 19222 524218 19404 524454
rect 18804 524134 19404 524218
rect 18804 523898 18986 524134
rect 19222 523898 19404 524134
rect 18804 488454 19404 523898
rect 18804 488218 18986 488454
rect 19222 488218 19404 488454
rect 18804 488134 19404 488218
rect 18804 487898 18986 488134
rect 19222 487898 19404 488134
rect 18804 452454 19404 487898
rect 18804 452218 18986 452454
rect 19222 452218 19404 452454
rect 18804 452134 19404 452218
rect 18804 451898 18986 452134
rect 19222 451898 19404 452134
rect 18804 416454 19404 451898
rect 18804 416218 18986 416454
rect 19222 416218 19404 416454
rect 18804 416134 19404 416218
rect 18804 415898 18986 416134
rect 19222 415898 19404 416134
rect 18804 380454 19404 415898
rect 18804 380218 18986 380454
rect 19222 380218 19404 380454
rect 18804 380134 19404 380218
rect 18804 379898 18986 380134
rect 19222 379898 19404 380134
rect 18804 344454 19404 379898
rect 18804 344218 18986 344454
rect 19222 344218 19404 344454
rect 18804 344134 19404 344218
rect 18804 343898 18986 344134
rect 19222 343898 19404 344134
rect 18804 308454 19404 343898
rect 18804 308218 18986 308454
rect 19222 308218 19404 308454
rect 18804 308134 19404 308218
rect 18804 307898 18986 308134
rect 19222 307898 19404 308134
rect 18804 272454 19404 307898
rect 18804 272218 18986 272454
rect 19222 272218 19404 272454
rect 18804 272134 19404 272218
rect 18804 271898 18986 272134
rect 19222 271898 19404 272134
rect 18804 236454 19404 271898
rect 18804 236218 18986 236454
rect 19222 236218 19404 236454
rect 18804 236134 19404 236218
rect 18804 235898 18986 236134
rect 19222 235898 19404 236134
rect 18804 200454 19404 235898
rect 18804 200218 18986 200454
rect 19222 200218 19404 200454
rect 18804 200134 19404 200218
rect 18804 199898 18986 200134
rect 19222 199898 19404 200134
rect 18804 164454 19404 199898
rect 18804 164218 18986 164454
rect 19222 164218 19404 164454
rect 18804 164134 19404 164218
rect 18804 163898 18986 164134
rect 19222 163898 19404 164134
rect 18804 128454 19404 163898
rect 18804 128218 18986 128454
rect 19222 128218 19404 128454
rect 18804 128134 19404 128218
rect 18804 127898 18986 128134
rect 19222 127898 19404 128134
rect 18804 92454 19404 127898
rect 18804 92218 18986 92454
rect 19222 92218 19404 92454
rect 18804 92134 19404 92218
rect 18804 91898 18986 92134
rect 19222 91898 19404 92134
rect 18804 56454 19404 91898
rect 18804 56218 18986 56454
rect 19222 56218 19404 56454
rect 18804 56134 19404 56218
rect 18804 55898 18986 56134
rect 19222 55898 19404 56134
rect 18804 20454 19404 55898
rect 18804 20218 18986 20454
rect 19222 20218 19404 20454
rect 18804 20134 19404 20218
rect 18804 19898 18986 20134
rect 19222 19898 19404 20134
rect 18804 -1286 19404 19898
rect 18804 -1522 18986 -1286
rect 19222 -1522 19404 -1286
rect 18804 -1606 19404 -1522
rect 18804 -1842 18986 -1606
rect 19222 -1842 19404 -1606
rect 18804 -1864 19404 -1842
rect 22404 672054 23004 707102
rect 22404 671818 22586 672054
rect 22822 671818 23004 672054
rect 22404 671734 23004 671818
rect 22404 671498 22586 671734
rect 22822 671498 23004 671734
rect 22404 636054 23004 671498
rect 22404 635818 22586 636054
rect 22822 635818 23004 636054
rect 22404 635734 23004 635818
rect 22404 635498 22586 635734
rect 22822 635498 23004 635734
rect 22404 600054 23004 635498
rect 22404 599818 22586 600054
rect 22822 599818 23004 600054
rect 22404 599734 23004 599818
rect 22404 599498 22586 599734
rect 22822 599498 23004 599734
rect 22404 564054 23004 599498
rect 22404 563818 22586 564054
rect 22822 563818 23004 564054
rect 22404 563734 23004 563818
rect 22404 563498 22586 563734
rect 22822 563498 23004 563734
rect 22404 528054 23004 563498
rect 22404 527818 22586 528054
rect 22822 527818 23004 528054
rect 22404 527734 23004 527818
rect 22404 527498 22586 527734
rect 22822 527498 23004 527734
rect 22404 492054 23004 527498
rect 22404 491818 22586 492054
rect 22822 491818 23004 492054
rect 22404 491734 23004 491818
rect 22404 491498 22586 491734
rect 22822 491498 23004 491734
rect 22404 456054 23004 491498
rect 22404 455818 22586 456054
rect 22822 455818 23004 456054
rect 22404 455734 23004 455818
rect 22404 455498 22586 455734
rect 22822 455498 23004 455734
rect 22404 420054 23004 455498
rect 22404 419818 22586 420054
rect 22822 419818 23004 420054
rect 22404 419734 23004 419818
rect 22404 419498 22586 419734
rect 22822 419498 23004 419734
rect 22404 384054 23004 419498
rect 22404 383818 22586 384054
rect 22822 383818 23004 384054
rect 22404 383734 23004 383818
rect 22404 383498 22586 383734
rect 22822 383498 23004 383734
rect 22404 348054 23004 383498
rect 22404 347818 22586 348054
rect 22822 347818 23004 348054
rect 22404 347734 23004 347818
rect 22404 347498 22586 347734
rect 22822 347498 23004 347734
rect 22404 312054 23004 347498
rect 22404 311818 22586 312054
rect 22822 311818 23004 312054
rect 22404 311734 23004 311818
rect 22404 311498 22586 311734
rect 22822 311498 23004 311734
rect 22404 276054 23004 311498
rect 22404 275818 22586 276054
rect 22822 275818 23004 276054
rect 22404 275734 23004 275818
rect 22404 275498 22586 275734
rect 22822 275498 23004 275734
rect 22404 240054 23004 275498
rect 22404 239818 22586 240054
rect 22822 239818 23004 240054
rect 22404 239734 23004 239818
rect 22404 239498 22586 239734
rect 22822 239498 23004 239734
rect 22404 204054 23004 239498
rect 22404 203818 22586 204054
rect 22822 203818 23004 204054
rect 22404 203734 23004 203818
rect 22404 203498 22586 203734
rect 22822 203498 23004 203734
rect 22404 168054 23004 203498
rect 22404 167818 22586 168054
rect 22822 167818 23004 168054
rect 22404 167734 23004 167818
rect 22404 167498 22586 167734
rect 22822 167498 23004 167734
rect 22404 132054 23004 167498
rect 22404 131818 22586 132054
rect 22822 131818 23004 132054
rect 22404 131734 23004 131818
rect 22404 131498 22586 131734
rect 22822 131498 23004 131734
rect 22404 96054 23004 131498
rect 22404 95818 22586 96054
rect 22822 95818 23004 96054
rect 22404 95734 23004 95818
rect 22404 95498 22586 95734
rect 22822 95498 23004 95734
rect 22404 60054 23004 95498
rect 22404 59818 22586 60054
rect 22822 59818 23004 60054
rect 22404 59734 23004 59818
rect 22404 59498 22586 59734
rect 22822 59498 23004 59734
rect 22404 24054 23004 59498
rect 22404 23818 22586 24054
rect 22822 23818 23004 24054
rect 22404 23734 23004 23818
rect 22404 23498 22586 23734
rect 22822 23498 23004 23734
rect 22404 -3166 23004 23498
rect 22404 -3402 22586 -3166
rect 22822 -3402 23004 -3166
rect 22404 -3486 23004 -3402
rect 22404 -3722 22586 -3486
rect 22822 -3722 23004 -3486
rect 22404 -3744 23004 -3722
rect 26004 675654 26604 708982
rect 26004 675418 26186 675654
rect 26422 675418 26604 675654
rect 26004 675334 26604 675418
rect 26004 675098 26186 675334
rect 26422 675098 26604 675334
rect 26004 639654 26604 675098
rect 26004 639418 26186 639654
rect 26422 639418 26604 639654
rect 26004 639334 26604 639418
rect 26004 639098 26186 639334
rect 26422 639098 26604 639334
rect 26004 603654 26604 639098
rect 26004 603418 26186 603654
rect 26422 603418 26604 603654
rect 26004 603334 26604 603418
rect 26004 603098 26186 603334
rect 26422 603098 26604 603334
rect 26004 567654 26604 603098
rect 26004 567418 26186 567654
rect 26422 567418 26604 567654
rect 26004 567334 26604 567418
rect 26004 567098 26186 567334
rect 26422 567098 26604 567334
rect 26004 531654 26604 567098
rect 26004 531418 26186 531654
rect 26422 531418 26604 531654
rect 26004 531334 26604 531418
rect 26004 531098 26186 531334
rect 26422 531098 26604 531334
rect 26004 495654 26604 531098
rect 26004 495418 26186 495654
rect 26422 495418 26604 495654
rect 26004 495334 26604 495418
rect 26004 495098 26186 495334
rect 26422 495098 26604 495334
rect 26004 459654 26604 495098
rect 26004 459418 26186 459654
rect 26422 459418 26604 459654
rect 26004 459334 26604 459418
rect 26004 459098 26186 459334
rect 26422 459098 26604 459334
rect 26004 423654 26604 459098
rect 26004 423418 26186 423654
rect 26422 423418 26604 423654
rect 26004 423334 26604 423418
rect 26004 423098 26186 423334
rect 26422 423098 26604 423334
rect 26004 387654 26604 423098
rect 26004 387418 26186 387654
rect 26422 387418 26604 387654
rect 26004 387334 26604 387418
rect 26004 387098 26186 387334
rect 26422 387098 26604 387334
rect 26004 351654 26604 387098
rect 26004 351418 26186 351654
rect 26422 351418 26604 351654
rect 26004 351334 26604 351418
rect 26004 351098 26186 351334
rect 26422 351098 26604 351334
rect 26004 315654 26604 351098
rect 26004 315418 26186 315654
rect 26422 315418 26604 315654
rect 26004 315334 26604 315418
rect 26004 315098 26186 315334
rect 26422 315098 26604 315334
rect 26004 279654 26604 315098
rect 26004 279418 26186 279654
rect 26422 279418 26604 279654
rect 26004 279334 26604 279418
rect 26004 279098 26186 279334
rect 26422 279098 26604 279334
rect 26004 243654 26604 279098
rect 26004 243418 26186 243654
rect 26422 243418 26604 243654
rect 26004 243334 26604 243418
rect 26004 243098 26186 243334
rect 26422 243098 26604 243334
rect 26004 207654 26604 243098
rect 26004 207418 26186 207654
rect 26422 207418 26604 207654
rect 26004 207334 26604 207418
rect 26004 207098 26186 207334
rect 26422 207098 26604 207334
rect 26004 171654 26604 207098
rect 26004 171418 26186 171654
rect 26422 171418 26604 171654
rect 26004 171334 26604 171418
rect 26004 171098 26186 171334
rect 26422 171098 26604 171334
rect 26004 135654 26604 171098
rect 26004 135418 26186 135654
rect 26422 135418 26604 135654
rect 26004 135334 26604 135418
rect 26004 135098 26186 135334
rect 26422 135098 26604 135334
rect 26004 99654 26604 135098
rect 26004 99418 26186 99654
rect 26422 99418 26604 99654
rect 26004 99334 26604 99418
rect 26004 99098 26186 99334
rect 26422 99098 26604 99334
rect 26004 63654 26604 99098
rect 26004 63418 26186 63654
rect 26422 63418 26604 63654
rect 26004 63334 26604 63418
rect 26004 63098 26186 63334
rect 26422 63098 26604 63334
rect 26004 27654 26604 63098
rect 26004 27418 26186 27654
rect 26422 27418 26604 27654
rect 26004 27334 26604 27418
rect 26004 27098 26186 27334
rect 26422 27098 26604 27334
rect 26004 -5046 26604 27098
rect 26004 -5282 26186 -5046
rect 26422 -5282 26604 -5046
rect 26004 -5366 26604 -5282
rect 26004 -5602 26186 -5366
rect 26422 -5602 26604 -5366
rect 26004 -5624 26604 -5602
rect 29604 679254 30204 710862
rect 47604 710478 48204 711440
rect 47604 710242 47786 710478
rect 48022 710242 48204 710478
rect 47604 710158 48204 710242
rect 47604 709922 47786 710158
rect 48022 709922 48204 710158
rect 44004 708598 44604 709560
rect 44004 708362 44186 708598
rect 44422 708362 44604 708598
rect 44004 708278 44604 708362
rect 44004 708042 44186 708278
rect 44422 708042 44604 708278
rect 40404 706718 41004 707680
rect 40404 706482 40586 706718
rect 40822 706482 41004 706718
rect 40404 706398 41004 706482
rect 40404 706162 40586 706398
rect 40822 706162 41004 706398
rect 29604 679018 29786 679254
rect 30022 679018 30204 679254
rect 29604 678934 30204 679018
rect 29604 678698 29786 678934
rect 30022 678698 30204 678934
rect 29604 643254 30204 678698
rect 29604 643018 29786 643254
rect 30022 643018 30204 643254
rect 29604 642934 30204 643018
rect 29604 642698 29786 642934
rect 30022 642698 30204 642934
rect 29604 607254 30204 642698
rect 29604 607018 29786 607254
rect 30022 607018 30204 607254
rect 29604 606934 30204 607018
rect 29604 606698 29786 606934
rect 30022 606698 30204 606934
rect 29604 571254 30204 606698
rect 29604 571018 29786 571254
rect 30022 571018 30204 571254
rect 29604 570934 30204 571018
rect 29604 570698 29786 570934
rect 30022 570698 30204 570934
rect 29604 535254 30204 570698
rect 29604 535018 29786 535254
rect 30022 535018 30204 535254
rect 29604 534934 30204 535018
rect 29604 534698 29786 534934
rect 30022 534698 30204 534934
rect 29604 499254 30204 534698
rect 29604 499018 29786 499254
rect 30022 499018 30204 499254
rect 29604 498934 30204 499018
rect 29604 498698 29786 498934
rect 30022 498698 30204 498934
rect 29604 463254 30204 498698
rect 29604 463018 29786 463254
rect 30022 463018 30204 463254
rect 29604 462934 30204 463018
rect 29604 462698 29786 462934
rect 30022 462698 30204 462934
rect 29604 427254 30204 462698
rect 29604 427018 29786 427254
rect 30022 427018 30204 427254
rect 29604 426934 30204 427018
rect 29604 426698 29786 426934
rect 30022 426698 30204 426934
rect 29604 391254 30204 426698
rect 29604 391018 29786 391254
rect 30022 391018 30204 391254
rect 29604 390934 30204 391018
rect 29604 390698 29786 390934
rect 30022 390698 30204 390934
rect 29604 355254 30204 390698
rect 29604 355018 29786 355254
rect 30022 355018 30204 355254
rect 29604 354934 30204 355018
rect 29604 354698 29786 354934
rect 30022 354698 30204 354934
rect 29604 319254 30204 354698
rect 29604 319018 29786 319254
rect 30022 319018 30204 319254
rect 29604 318934 30204 319018
rect 29604 318698 29786 318934
rect 30022 318698 30204 318934
rect 29604 283254 30204 318698
rect 29604 283018 29786 283254
rect 30022 283018 30204 283254
rect 29604 282934 30204 283018
rect 29604 282698 29786 282934
rect 30022 282698 30204 282934
rect 29604 247254 30204 282698
rect 29604 247018 29786 247254
rect 30022 247018 30204 247254
rect 29604 246934 30204 247018
rect 29604 246698 29786 246934
rect 30022 246698 30204 246934
rect 29604 211254 30204 246698
rect 29604 211018 29786 211254
rect 30022 211018 30204 211254
rect 29604 210934 30204 211018
rect 29604 210698 29786 210934
rect 30022 210698 30204 210934
rect 29604 175254 30204 210698
rect 29604 175018 29786 175254
rect 30022 175018 30204 175254
rect 29604 174934 30204 175018
rect 29604 174698 29786 174934
rect 30022 174698 30204 174934
rect 29604 139254 30204 174698
rect 29604 139018 29786 139254
rect 30022 139018 30204 139254
rect 29604 138934 30204 139018
rect 29604 138698 29786 138934
rect 30022 138698 30204 138934
rect 29604 103254 30204 138698
rect 29604 103018 29786 103254
rect 30022 103018 30204 103254
rect 29604 102934 30204 103018
rect 29604 102698 29786 102934
rect 30022 102698 30204 102934
rect 29604 67254 30204 102698
rect 29604 67018 29786 67254
rect 30022 67018 30204 67254
rect 29604 66934 30204 67018
rect 29604 66698 29786 66934
rect 30022 66698 30204 66934
rect 29604 31254 30204 66698
rect 29604 31018 29786 31254
rect 30022 31018 30204 31254
rect 29604 30934 30204 31018
rect 29604 30698 29786 30934
rect 30022 30698 30204 30934
rect 11604 -6222 11786 -5986
rect 12022 -6222 12204 -5986
rect 11604 -6306 12204 -6222
rect 11604 -6542 11786 -6306
rect 12022 -6542 12204 -6306
rect -8576 -7162 -8394 -6926
rect -8158 -7162 -7976 -6926
rect -8576 -7246 -7976 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 -7976 -7246
rect -8576 -7504 -7976 -7482
rect 11604 -7504 12204 -6542
rect 29604 -6926 30204 30698
rect 36804 704838 37404 705800
rect 36804 704602 36986 704838
rect 37222 704602 37404 704838
rect 36804 704518 37404 704602
rect 36804 704282 36986 704518
rect 37222 704282 37404 704518
rect 36804 686454 37404 704282
rect 36804 686218 36986 686454
rect 37222 686218 37404 686454
rect 36804 686134 37404 686218
rect 36804 685898 36986 686134
rect 37222 685898 37404 686134
rect 36804 650454 37404 685898
rect 36804 650218 36986 650454
rect 37222 650218 37404 650454
rect 36804 650134 37404 650218
rect 36804 649898 36986 650134
rect 37222 649898 37404 650134
rect 36804 614454 37404 649898
rect 36804 614218 36986 614454
rect 37222 614218 37404 614454
rect 36804 614134 37404 614218
rect 36804 613898 36986 614134
rect 37222 613898 37404 614134
rect 36804 578454 37404 613898
rect 36804 578218 36986 578454
rect 37222 578218 37404 578454
rect 36804 578134 37404 578218
rect 36804 577898 36986 578134
rect 37222 577898 37404 578134
rect 36804 542454 37404 577898
rect 36804 542218 36986 542454
rect 37222 542218 37404 542454
rect 36804 542134 37404 542218
rect 36804 541898 36986 542134
rect 37222 541898 37404 542134
rect 36804 506454 37404 541898
rect 36804 506218 36986 506454
rect 37222 506218 37404 506454
rect 36804 506134 37404 506218
rect 36804 505898 36986 506134
rect 37222 505898 37404 506134
rect 36804 470454 37404 505898
rect 36804 470218 36986 470454
rect 37222 470218 37404 470454
rect 36804 470134 37404 470218
rect 36804 469898 36986 470134
rect 37222 469898 37404 470134
rect 36804 434454 37404 469898
rect 36804 434218 36986 434454
rect 37222 434218 37404 434454
rect 36804 434134 37404 434218
rect 36804 433898 36986 434134
rect 37222 433898 37404 434134
rect 36804 398454 37404 433898
rect 36804 398218 36986 398454
rect 37222 398218 37404 398454
rect 36804 398134 37404 398218
rect 36804 397898 36986 398134
rect 37222 397898 37404 398134
rect 36804 362454 37404 397898
rect 36804 362218 36986 362454
rect 37222 362218 37404 362454
rect 36804 362134 37404 362218
rect 36804 361898 36986 362134
rect 37222 361898 37404 362134
rect 36804 326454 37404 361898
rect 36804 326218 36986 326454
rect 37222 326218 37404 326454
rect 36804 326134 37404 326218
rect 36804 325898 36986 326134
rect 37222 325898 37404 326134
rect 36804 290454 37404 325898
rect 36804 290218 36986 290454
rect 37222 290218 37404 290454
rect 36804 290134 37404 290218
rect 36804 289898 36986 290134
rect 37222 289898 37404 290134
rect 36804 254454 37404 289898
rect 36804 254218 36986 254454
rect 37222 254218 37404 254454
rect 36804 254134 37404 254218
rect 36804 253898 36986 254134
rect 37222 253898 37404 254134
rect 36804 218454 37404 253898
rect 36804 218218 36986 218454
rect 37222 218218 37404 218454
rect 36804 218134 37404 218218
rect 36804 217898 36986 218134
rect 37222 217898 37404 218134
rect 36804 182454 37404 217898
rect 36804 182218 36986 182454
rect 37222 182218 37404 182454
rect 36804 182134 37404 182218
rect 36804 181898 36986 182134
rect 37222 181898 37404 182134
rect 36804 146454 37404 181898
rect 36804 146218 36986 146454
rect 37222 146218 37404 146454
rect 36804 146134 37404 146218
rect 36804 145898 36986 146134
rect 37222 145898 37404 146134
rect 36804 110454 37404 145898
rect 36804 110218 36986 110454
rect 37222 110218 37404 110454
rect 36804 110134 37404 110218
rect 36804 109898 36986 110134
rect 37222 109898 37404 110134
rect 36804 74454 37404 109898
rect 36804 74218 36986 74454
rect 37222 74218 37404 74454
rect 36804 74134 37404 74218
rect 36804 73898 36986 74134
rect 37222 73898 37404 74134
rect 36804 38454 37404 73898
rect 36804 38218 36986 38454
rect 37222 38218 37404 38454
rect 36804 38134 37404 38218
rect 36804 37898 36986 38134
rect 37222 37898 37404 38134
rect 36804 2454 37404 37898
rect 36804 2218 36986 2454
rect 37222 2218 37404 2454
rect 36804 2134 37404 2218
rect 36804 1898 36986 2134
rect 37222 1898 37404 2134
rect 36804 -346 37404 1898
rect 36804 -582 36986 -346
rect 37222 -582 37404 -346
rect 36804 -666 37404 -582
rect 36804 -902 36986 -666
rect 37222 -902 37404 -666
rect 36804 -1864 37404 -902
rect 40404 690054 41004 706162
rect 40404 689818 40586 690054
rect 40822 689818 41004 690054
rect 40404 689734 41004 689818
rect 40404 689498 40586 689734
rect 40822 689498 41004 689734
rect 40404 654054 41004 689498
rect 40404 653818 40586 654054
rect 40822 653818 41004 654054
rect 40404 653734 41004 653818
rect 40404 653498 40586 653734
rect 40822 653498 41004 653734
rect 40404 618054 41004 653498
rect 40404 617818 40586 618054
rect 40822 617818 41004 618054
rect 40404 617734 41004 617818
rect 40404 617498 40586 617734
rect 40822 617498 41004 617734
rect 40404 582054 41004 617498
rect 40404 581818 40586 582054
rect 40822 581818 41004 582054
rect 40404 581734 41004 581818
rect 40404 581498 40586 581734
rect 40822 581498 41004 581734
rect 40404 546054 41004 581498
rect 40404 545818 40586 546054
rect 40822 545818 41004 546054
rect 40404 545734 41004 545818
rect 40404 545498 40586 545734
rect 40822 545498 41004 545734
rect 40404 510054 41004 545498
rect 40404 509818 40586 510054
rect 40822 509818 41004 510054
rect 40404 509734 41004 509818
rect 40404 509498 40586 509734
rect 40822 509498 41004 509734
rect 40404 474054 41004 509498
rect 40404 473818 40586 474054
rect 40822 473818 41004 474054
rect 40404 473734 41004 473818
rect 40404 473498 40586 473734
rect 40822 473498 41004 473734
rect 40404 438054 41004 473498
rect 40404 437818 40586 438054
rect 40822 437818 41004 438054
rect 40404 437734 41004 437818
rect 40404 437498 40586 437734
rect 40822 437498 41004 437734
rect 40404 402054 41004 437498
rect 40404 401818 40586 402054
rect 40822 401818 41004 402054
rect 40404 401734 41004 401818
rect 40404 401498 40586 401734
rect 40822 401498 41004 401734
rect 40404 366054 41004 401498
rect 40404 365818 40586 366054
rect 40822 365818 41004 366054
rect 40404 365734 41004 365818
rect 40404 365498 40586 365734
rect 40822 365498 41004 365734
rect 40404 330054 41004 365498
rect 40404 329818 40586 330054
rect 40822 329818 41004 330054
rect 40404 329734 41004 329818
rect 40404 329498 40586 329734
rect 40822 329498 41004 329734
rect 40404 294054 41004 329498
rect 40404 293818 40586 294054
rect 40822 293818 41004 294054
rect 40404 293734 41004 293818
rect 40404 293498 40586 293734
rect 40822 293498 41004 293734
rect 40404 258054 41004 293498
rect 40404 257818 40586 258054
rect 40822 257818 41004 258054
rect 40404 257734 41004 257818
rect 40404 257498 40586 257734
rect 40822 257498 41004 257734
rect 40404 222054 41004 257498
rect 40404 221818 40586 222054
rect 40822 221818 41004 222054
rect 40404 221734 41004 221818
rect 40404 221498 40586 221734
rect 40822 221498 41004 221734
rect 40404 186054 41004 221498
rect 40404 185818 40586 186054
rect 40822 185818 41004 186054
rect 40404 185734 41004 185818
rect 40404 185498 40586 185734
rect 40822 185498 41004 185734
rect 40404 150054 41004 185498
rect 40404 149818 40586 150054
rect 40822 149818 41004 150054
rect 40404 149734 41004 149818
rect 40404 149498 40586 149734
rect 40822 149498 41004 149734
rect 40404 114054 41004 149498
rect 40404 113818 40586 114054
rect 40822 113818 41004 114054
rect 40404 113734 41004 113818
rect 40404 113498 40586 113734
rect 40822 113498 41004 113734
rect 40404 78054 41004 113498
rect 40404 77818 40586 78054
rect 40822 77818 41004 78054
rect 40404 77734 41004 77818
rect 40404 77498 40586 77734
rect 40822 77498 41004 77734
rect 40404 42054 41004 77498
rect 40404 41818 40586 42054
rect 40822 41818 41004 42054
rect 40404 41734 41004 41818
rect 40404 41498 40586 41734
rect 40822 41498 41004 41734
rect 40404 6054 41004 41498
rect 40404 5818 40586 6054
rect 40822 5818 41004 6054
rect 40404 5734 41004 5818
rect 40404 5498 40586 5734
rect 40822 5498 41004 5734
rect 40404 -2226 41004 5498
rect 40404 -2462 40586 -2226
rect 40822 -2462 41004 -2226
rect 40404 -2546 41004 -2462
rect 40404 -2782 40586 -2546
rect 40822 -2782 41004 -2546
rect 40404 -3744 41004 -2782
rect 44004 693654 44604 708042
rect 44004 693418 44186 693654
rect 44422 693418 44604 693654
rect 44004 693334 44604 693418
rect 44004 693098 44186 693334
rect 44422 693098 44604 693334
rect 44004 657654 44604 693098
rect 44004 657418 44186 657654
rect 44422 657418 44604 657654
rect 44004 657334 44604 657418
rect 44004 657098 44186 657334
rect 44422 657098 44604 657334
rect 44004 621654 44604 657098
rect 44004 621418 44186 621654
rect 44422 621418 44604 621654
rect 44004 621334 44604 621418
rect 44004 621098 44186 621334
rect 44422 621098 44604 621334
rect 44004 585654 44604 621098
rect 44004 585418 44186 585654
rect 44422 585418 44604 585654
rect 44004 585334 44604 585418
rect 44004 585098 44186 585334
rect 44422 585098 44604 585334
rect 44004 549654 44604 585098
rect 44004 549418 44186 549654
rect 44422 549418 44604 549654
rect 44004 549334 44604 549418
rect 44004 549098 44186 549334
rect 44422 549098 44604 549334
rect 44004 513654 44604 549098
rect 44004 513418 44186 513654
rect 44422 513418 44604 513654
rect 44004 513334 44604 513418
rect 44004 513098 44186 513334
rect 44422 513098 44604 513334
rect 44004 477654 44604 513098
rect 44004 477418 44186 477654
rect 44422 477418 44604 477654
rect 44004 477334 44604 477418
rect 44004 477098 44186 477334
rect 44422 477098 44604 477334
rect 44004 441654 44604 477098
rect 44004 441418 44186 441654
rect 44422 441418 44604 441654
rect 44004 441334 44604 441418
rect 44004 441098 44186 441334
rect 44422 441098 44604 441334
rect 44004 405654 44604 441098
rect 44004 405418 44186 405654
rect 44422 405418 44604 405654
rect 44004 405334 44604 405418
rect 44004 405098 44186 405334
rect 44422 405098 44604 405334
rect 44004 369654 44604 405098
rect 44004 369418 44186 369654
rect 44422 369418 44604 369654
rect 44004 369334 44604 369418
rect 44004 369098 44186 369334
rect 44422 369098 44604 369334
rect 44004 333654 44604 369098
rect 44004 333418 44186 333654
rect 44422 333418 44604 333654
rect 44004 333334 44604 333418
rect 44004 333098 44186 333334
rect 44422 333098 44604 333334
rect 44004 297654 44604 333098
rect 44004 297418 44186 297654
rect 44422 297418 44604 297654
rect 44004 297334 44604 297418
rect 44004 297098 44186 297334
rect 44422 297098 44604 297334
rect 44004 261654 44604 297098
rect 44004 261418 44186 261654
rect 44422 261418 44604 261654
rect 44004 261334 44604 261418
rect 44004 261098 44186 261334
rect 44422 261098 44604 261334
rect 44004 225654 44604 261098
rect 44004 225418 44186 225654
rect 44422 225418 44604 225654
rect 44004 225334 44604 225418
rect 44004 225098 44186 225334
rect 44422 225098 44604 225334
rect 44004 189654 44604 225098
rect 44004 189418 44186 189654
rect 44422 189418 44604 189654
rect 44004 189334 44604 189418
rect 44004 189098 44186 189334
rect 44422 189098 44604 189334
rect 44004 153654 44604 189098
rect 44004 153418 44186 153654
rect 44422 153418 44604 153654
rect 44004 153334 44604 153418
rect 44004 153098 44186 153334
rect 44422 153098 44604 153334
rect 44004 117654 44604 153098
rect 44004 117418 44186 117654
rect 44422 117418 44604 117654
rect 44004 117334 44604 117418
rect 44004 117098 44186 117334
rect 44422 117098 44604 117334
rect 44004 81654 44604 117098
rect 44004 81418 44186 81654
rect 44422 81418 44604 81654
rect 44004 81334 44604 81418
rect 44004 81098 44186 81334
rect 44422 81098 44604 81334
rect 44004 45654 44604 81098
rect 44004 45418 44186 45654
rect 44422 45418 44604 45654
rect 44004 45334 44604 45418
rect 44004 45098 44186 45334
rect 44422 45098 44604 45334
rect 44004 9654 44604 45098
rect 44004 9418 44186 9654
rect 44422 9418 44604 9654
rect 44004 9334 44604 9418
rect 44004 9098 44186 9334
rect 44422 9098 44604 9334
rect 44004 -4106 44604 9098
rect 44004 -4342 44186 -4106
rect 44422 -4342 44604 -4106
rect 44004 -4426 44604 -4342
rect 44004 -4662 44186 -4426
rect 44422 -4662 44604 -4426
rect 44004 -5624 44604 -4662
rect 47604 697254 48204 709922
rect 65604 711418 66204 711440
rect 65604 711182 65786 711418
rect 66022 711182 66204 711418
rect 65604 711098 66204 711182
rect 65604 710862 65786 711098
rect 66022 710862 66204 711098
rect 62004 709538 62604 709560
rect 62004 709302 62186 709538
rect 62422 709302 62604 709538
rect 62004 709218 62604 709302
rect 62004 708982 62186 709218
rect 62422 708982 62604 709218
rect 58404 707658 59004 707680
rect 58404 707422 58586 707658
rect 58822 707422 59004 707658
rect 58404 707338 59004 707422
rect 58404 707102 58586 707338
rect 58822 707102 59004 707338
rect 47604 697018 47786 697254
rect 48022 697018 48204 697254
rect 47604 696934 48204 697018
rect 47604 696698 47786 696934
rect 48022 696698 48204 696934
rect 47604 661254 48204 696698
rect 47604 661018 47786 661254
rect 48022 661018 48204 661254
rect 47604 660934 48204 661018
rect 47604 660698 47786 660934
rect 48022 660698 48204 660934
rect 47604 625254 48204 660698
rect 47604 625018 47786 625254
rect 48022 625018 48204 625254
rect 47604 624934 48204 625018
rect 47604 624698 47786 624934
rect 48022 624698 48204 624934
rect 47604 589254 48204 624698
rect 47604 589018 47786 589254
rect 48022 589018 48204 589254
rect 47604 588934 48204 589018
rect 47604 588698 47786 588934
rect 48022 588698 48204 588934
rect 47604 553254 48204 588698
rect 47604 553018 47786 553254
rect 48022 553018 48204 553254
rect 47604 552934 48204 553018
rect 47604 552698 47786 552934
rect 48022 552698 48204 552934
rect 47604 517254 48204 552698
rect 47604 517018 47786 517254
rect 48022 517018 48204 517254
rect 47604 516934 48204 517018
rect 47604 516698 47786 516934
rect 48022 516698 48204 516934
rect 47604 481254 48204 516698
rect 47604 481018 47786 481254
rect 48022 481018 48204 481254
rect 47604 480934 48204 481018
rect 47604 480698 47786 480934
rect 48022 480698 48204 480934
rect 47604 445254 48204 480698
rect 47604 445018 47786 445254
rect 48022 445018 48204 445254
rect 47604 444934 48204 445018
rect 47604 444698 47786 444934
rect 48022 444698 48204 444934
rect 47604 409254 48204 444698
rect 47604 409018 47786 409254
rect 48022 409018 48204 409254
rect 47604 408934 48204 409018
rect 47604 408698 47786 408934
rect 48022 408698 48204 408934
rect 47604 373254 48204 408698
rect 47604 373018 47786 373254
rect 48022 373018 48204 373254
rect 47604 372934 48204 373018
rect 47604 372698 47786 372934
rect 48022 372698 48204 372934
rect 47604 337254 48204 372698
rect 47604 337018 47786 337254
rect 48022 337018 48204 337254
rect 47604 336934 48204 337018
rect 47604 336698 47786 336934
rect 48022 336698 48204 336934
rect 47604 301254 48204 336698
rect 47604 301018 47786 301254
rect 48022 301018 48204 301254
rect 47604 300934 48204 301018
rect 47604 300698 47786 300934
rect 48022 300698 48204 300934
rect 47604 265254 48204 300698
rect 47604 265018 47786 265254
rect 48022 265018 48204 265254
rect 47604 264934 48204 265018
rect 47604 264698 47786 264934
rect 48022 264698 48204 264934
rect 47604 229254 48204 264698
rect 47604 229018 47786 229254
rect 48022 229018 48204 229254
rect 47604 228934 48204 229018
rect 47604 228698 47786 228934
rect 48022 228698 48204 228934
rect 47604 193254 48204 228698
rect 47604 193018 47786 193254
rect 48022 193018 48204 193254
rect 47604 192934 48204 193018
rect 47604 192698 47786 192934
rect 48022 192698 48204 192934
rect 47604 157254 48204 192698
rect 47604 157018 47786 157254
rect 48022 157018 48204 157254
rect 47604 156934 48204 157018
rect 47604 156698 47786 156934
rect 48022 156698 48204 156934
rect 47604 121254 48204 156698
rect 47604 121018 47786 121254
rect 48022 121018 48204 121254
rect 47604 120934 48204 121018
rect 47604 120698 47786 120934
rect 48022 120698 48204 120934
rect 47604 85254 48204 120698
rect 47604 85018 47786 85254
rect 48022 85018 48204 85254
rect 47604 84934 48204 85018
rect 47604 84698 47786 84934
rect 48022 84698 48204 84934
rect 47604 49254 48204 84698
rect 47604 49018 47786 49254
rect 48022 49018 48204 49254
rect 47604 48934 48204 49018
rect 47604 48698 47786 48934
rect 48022 48698 48204 48934
rect 47604 13254 48204 48698
rect 47604 13018 47786 13254
rect 48022 13018 48204 13254
rect 47604 12934 48204 13018
rect 47604 12698 47786 12934
rect 48022 12698 48204 12934
rect 29604 -7162 29786 -6926
rect 30022 -7162 30204 -6926
rect 29604 -7246 30204 -7162
rect 29604 -7482 29786 -7246
rect 30022 -7482 30204 -7246
rect 29604 -7504 30204 -7482
rect 47604 -5986 48204 12698
rect 54804 705778 55404 705800
rect 54804 705542 54986 705778
rect 55222 705542 55404 705778
rect 54804 705458 55404 705542
rect 54804 705222 54986 705458
rect 55222 705222 55404 705458
rect 54804 668454 55404 705222
rect 54804 668218 54986 668454
rect 55222 668218 55404 668454
rect 54804 668134 55404 668218
rect 54804 667898 54986 668134
rect 55222 667898 55404 668134
rect 54804 632454 55404 667898
rect 58404 672054 59004 707102
rect 58404 671818 58586 672054
rect 58822 671818 59004 672054
rect 58404 671734 59004 671818
rect 58404 671498 58586 671734
rect 58822 671498 59004 671734
rect 58404 654247 59004 671498
rect 62004 675654 62604 708982
rect 62004 675418 62186 675654
rect 62422 675418 62604 675654
rect 62004 675334 62604 675418
rect 62004 675098 62186 675334
rect 62422 675098 62604 675334
rect 62004 654247 62604 675098
rect 65604 679254 66204 710862
rect 83604 710478 84204 711440
rect 83604 710242 83786 710478
rect 84022 710242 84204 710478
rect 83604 710158 84204 710242
rect 83604 709922 83786 710158
rect 84022 709922 84204 710158
rect 80004 708598 80604 709560
rect 80004 708362 80186 708598
rect 80422 708362 80604 708598
rect 80004 708278 80604 708362
rect 80004 708042 80186 708278
rect 80422 708042 80604 708278
rect 76404 706718 77004 707680
rect 76404 706482 76586 706718
rect 76822 706482 77004 706718
rect 76404 706398 77004 706482
rect 76404 706162 76586 706398
rect 76822 706162 77004 706398
rect 65604 679018 65786 679254
rect 66022 679018 66204 679254
rect 65604 678934 66204 679018
rect 65604 678698 65786 678934
rect 66022 678698 66204 678934
rect 65604 654247 66204 678698
rect 72804 704838 73404 705800
rect 72804 704602 72986 704838
rect 73222 704602 73404 704838
rect 72804 704518 73404 704602
rect 72804 704282 72986 704518
rect 73222 704282 73404 704518
rect 72804 686454 73404 704282
rect 72804 686218 72986 686454
rect 73222 686218 73404 686454
rect 72804 686134 73404 686218
rect 72804 685898 72986 686134
rect 73222 685898 73404 686134
rect 72804 654247 73404 685898
rect 76404 690054 77004 706162
rect 76404 689818 76586 690054
rect 76822 689818 77004 690054
rect 76404 689734 77004 689818
rect 76404 689498 76586 689734
rect 76822 689498 77004 689734
rect 76404 654247 77004 689498
rect 80004 693654 80604 708042
rect 80004 693418 80186 693654
rect 80422 693418 80604 693654
rect 80004 693334 80604 693418
rect 80004 693098 80186 693334
rect 80422 693098 80604 693334
rect 80004 657654 80604 693098
rect 80004 657418 80186 657654
rect 80422 657418 80604 657654
rect 80004 657334 80604 657418
rect 80004 657098 80186 657334
rect 80422 657098 80604 657334
rect 80004 654247 80604 657098
rect 83604 697254 84204 709922
rect 101604 711418 102204 711440
rect 101604 711182 101786 711418
rect 102022 711182 102204 711418
rect 101604 711098 102204 711182
rect 101604 710862 101786 711098
rect 102022 710862 102204 711098
rect 98004 709538 98604 709560
rect 98004 709302 98186 709538
rect 98422 709302 98604 709538
rect 98004 709218 98604 709302
rect 98004 708982 98186 709218
rect 98422 708982 98604 709218
rect 94404 707658 95004 707680
rect 94404 707422 94586 707658
rect 94822 707422 95004 707658
rect 94404 707338 95004 707422
rect 94404 707102 94586 707338
rect 94822 707102 95004 707338
rect 83604 697018 83786 697254
rect 84022 697018 84204 697254
rect 83604 696934 84204 697018
rect 83604 696698 83786 696934
rect 84022 696698 84204 696934
rect 83604 661254 84204 696698
rect 83604 661018 83786 661254
rect 84022 661018 84204 661254
rect 83604 660934 84204 661018
rect 83604 660698 83786 660934
rect 84022 660698 84204 660934
rect 83604 654247 84204 660698
rect 90804 705778 91404 705800
rect 90804 705542 90986 705778
rect 91222 705542 91404 705778
rect 90804 705458 91404 705542
rect 90804 705222 90986 705458
rect 91222 705222 91404 705458
rect 90804 668454 91404 705222
rect 90804 668218 90986 668454
rect 91222 668218 91404 668454
rect 90804 668134 91404 668218
rect 90804 667898 90986 668134
rect 91222 667898 91404 668134
rect 90804 654247 91404 667898
rect 94404 672054 95004 707102
rect 94404 671818 94586 672054
rect 94822 671818 95004 672054
rect 94404 671734 95004 671818
rect 94404 671498 94586 671734
rect 94822 671498 95004 671734
rect 94404 654247 95004 671498
rect 98004 675654 98604 708982
rect 98004 675418 98186 675654
rect 98422 675418 98604 675654
rect 98004 675334 98604 675418
rect 98004 675098 98186 675334
rect 98422 675098 98604 675334
rect 98004 654247 98604 675098
rect 101604 679254 102204 710862
rect 119604 710478 120204 711440
rect 119604 710242 119786 710478
rect 120022 710242 120204 710478
rect 119604 710158 120204 710242
rect 119604 709922 119786 710158
rect 120022 709922 120204 710158
rect 116004 708598 116604 709560
rect 116004 708362 116186 708598
rect 116422 708362 116604 708598
rect 116004 708278 116604 708362
rect 116004 708042 116186 708278
rect 116422 708042 116604 708278
rect 112404 706718 113004 707680
rect 112404 706482 112586 706718
rect 112822 706482 113004 706718
rect 112404 706398 113004 706482
rect 112404 706162 112586 706398
rect 112822 706162 113004 706398
rect 101604 679018 101786 679254
rect 102022 679018 102204 679254
rect 101604 678934 102204 679018
rect 101604 678698 101786 678934
rect 102022 678698 102204 678934
rect 101604 654247 102204 678698
rect 108804 704838 109404 705800
rect 108804 704602 108986 704838
rect 109222 704602 109404 704838
rect 108804 704518 109404 704602
rect 108804 704282 108986 704518
rect 109222 704282 109404 704518
rect 108804 686454 109404 704282
rect 108804 686218 108986 686454
rect 109222 686218 109404 686454
rect 108804 686134 109404 686218
rect 108804 685898 108986 686134
rect 109222 685898 109404 686134
rect 108804 654247 109404 685898
rect 112404 690054 113004 706162
rect 112404 689818 112586 690054
rect 112822 689818 113004 690054
rect 112404 689734 113004 689818
rect 112404 689498 112586 689734
rect 112822 689498 113004 689734
rect 112404 654247 113004 689498
rect 116004 693654 116604 708042
rect 116004 693418 116186 693654
rect 116422 693418 116604 693654
rect 116004 693334 116604 693418
rect 116004 693098 116186 693334
rect 116422 693098 116604 693334
rect 116004 657654 116604 693098
rect 116004 657418 116186 657654
rect 116422 657418 116604 657654
rect 116004 657334 116604 657418
rect 116004 657098 116186 657334
rect 116422 657098 116604 657334
rect 116004 654247 116604 657098
rect 119604 697254 120204 709922
rect 137604 711418 138204 711440
rect 137604 711182 137786 711418
rect 138022 711182 138204 711418
rect 137604 711098 138204 711182
rect 137604 710862 137786 711098
rect 138022 710862 138204 711098
rect 134004 709538 134604 709560
rect 134004 709302 134186 709538
rect 134422 709302 134604 709538
rect 134004 709218 134604 709302
rect 134004 708982 134186 709218
rect 134422 708982 134604 709218
rect 130404 707658 131004 707680
rect 130404 707422 130586 707658
rect 130822 707422 131004 707658
rect 130404 707338 131004 707422
rect 130404 707102 130586 707338
rect 130822 707102 131004 707338
rect 119604 697018 119786 697254
rect 120022 697018 120204 697254
rect 119604 696934 120204 697018
rect 119604 696698 119786 696934
rect 120022 696698 120204 696934
rect 119604 661254 120204 696698
rect 119604 661018 119786 661254
rect 120022 661018 120204 661254
rect 119604 660934 120204 661018
rect 119604 660698 119786 660934
rect 120022 660698 120204 660934
rect 119604 654247 120204 660698
rect 126804 705778 127404 705800
rect 126804 705542 126986 705778
rect 127222 705542 127404 705778
rect 126804 705458 127404 705542
rect 126804 705222 126986 705458
rect 127222 705222 127404 705458
rect 126804 668454 127404 705222
rect 126804 668218 126986 668454
rect 127222 668218 127404 668454
rect 126804 668134 127404 668218
rect 126804 667898 126986 668134
rect 127222 667898 127404 668134
rect 126804 654247 127404 667898
rect 130404 672054 131004 707102
rect 130404 671818 130586 672054
rect 130822 671818 131004 672054
rect 130404 671734 131004 671818
rect 130404 671498 130586 671734
rect 130822 671498 131004 671734
rect 130404 654247 131004 671498
rect 134004 675654 134604 708982
rect 134004 675418 134186 675654
rect 134422 675418 134604 675654
rect 134004 675334 134604 675418
rect 134004 675098 134186 675334
rect 134422 675098 134604 675334
rect 134004 654247 134604 675098
rect 137604 679254 138204 710862
rect 155604 710478 156204 711440
rect 155604 710242 155786 710478
rect 156022 710242 156204 710478
rect 155604 710158 156204 710242
rect 155604 709922 155786 710158
rect 156022 709922 156204 710158
rect 152004 708598 152604 709560
rect 152004 708362 152186 708598
rect 152422 708362 152604 708598
rect 152004 708278 152604 708362
rect 152004 708042 152186 708278
rect 152422 708042 152604 708278
rect 148404 706718 149004 707680
rect 148404 706482 148586 706718
rect 148822 706482 149004 706718
rect 148404 706398 149004 706482
rect 148404 706162 148586 706398
rect 148822 706162 149004 706398
rect 137604 679018 137786 679254
rect 138022 679018 138204 679254
rect 137604 678934 138204 679018
rect 137604 678698 137786 678934
rect 138022 678698 138204 678934
rect 137604 654247 138204 678698
rect 144804 704838 145404 705800
rect 144804 704602 144986 704838
rect 145222 704602 145404 704838
rect 144804 704518 145404 704602
rect 144804 704282 144986 704518
rect 145222 704282 145404 704518
rect 144804 686454 145404 704282
rect 144804 686218 144986 686454
rect 145222 686218 145404 686454
rect 144804 686134 145404 686218
rect 144804 685898 144986 686134
rect 145222 685898 145404 686134
rect 129227 651132 129293 651133
rect 129227 651130 129228 651132
rect 128608 651070 129228 651130
rect 129227 651068 129228 651070
rect 129292 651068 129293 651132
rect 129227 651067 129293 651068
rect 133827 651132 133893 651133
rect 133827 651068 133828 651132
rect 133892 651068 133893 651132
rect 133827 651067 133893 651068
rect 133830 650790 133890 651067
rect 133603 650730 133890 650790
rect 144804 650454 145404 685898
rect 144804 650218 144986 650454
rect 145222 650218 145404 650454
rect 144804 650134 145404 650218
rect 144804 649898 144986 650134
rect 145222 649898 145404 650134
rect 136938 643254 137262 643276
rect 136938 643018 136982 643254
rect 137218 643018 137262 643254
rect 136938 642934 137262 643018
rect 136938 642698 136982 642934
rect 137218 642698 137262 642934
rect 136938 642676 137262 642698
rect 136938 639654 137262 639676
rect 136938 639418 136982 639654
rect 137218 639418 137262 639654
rect 136938 639334 137262 639418
rect 136938 639098 136982 639334
rect 137218 639098 137262 639334
rect 136938 639076 137262 639098
rect 136938 636054 137262 636076
rect 136938 635818 136982 636054
rect 137218 635818 137262 636054
rect 136938 635734 137262 635818
rect 136938 635498 136982 635734
rect 137218 635498 137262 635734
rect 136938 635476 137262 635498
rect 54804 632218 54986 632454
rect 55222 632218 55404 632454
rect 54804 632134 55404 632218
rect 54804 631898 54986 632134
rect 55222 631898 55404 632134
rect 54804 596454 55404 631898
rect 136938 632454 137262 632476
rect 136938 632218 136982 632454
rect 137218 632218 137262 632454
rect 136938 632134 137262 632218
rect 136938 631898 136982 632134
rect 137218 631898 137262 632134
rect 136938 631876 137262 631898
rect 136494 625254 136814 625276
rect 136494 625018 136536 625254
rect 136772 625018 136814 625254
rect 136494 624934 136814 625018
rect 136494 624698 136536 624934
rect 136772 624698 136814 624934
rect 136494 624676 136814 624698
rect 136494 621654 136814 621676
rect 136494 621418 136536 621654
rect 136772 621418 136814 621654
rect 136494 621334 136814 621418
rect 136494 621098 136536 621334
rect 136772 621098 136814 621334
rect 136494 621076 136814 621098
rect 136494 618054 136814 618076
rect 136494 617818 136536 618054
rect 136772 617818 136814 618054
rect 136494 617734 136814 617818
rect 136494 617498 136536 617734
rect 136772 617498 136814 617734
rect 136494 617476 136814 617498
rect 136494 614454 136814 614476
rect 136494 614218 136536 614454
rect 136772 614218 136814 614454
rect 136494 614134 136814 614218
rect 136494 613898 136536 614134
rect 136772 613898 136814 614134
rect 136494 613876 136814 613898
rect 144804 614454 145404 649898
rect 144804 614218 144986 614454
rect 145222 614218 145404 614454
rect 144804 614134 145404 614218
rect 144804 613898 144986 614134
rect 145222 613898 145404 614134
rect 136938 607254 137262 607276
rect 136938 607018 136982 607254
rect 137218 607018 137262 607254
rect 136938 606934 137262 607018
rect 136938 606698 136982 606934
rect 137218 606698 137262 606934
rect 136938 606676 137262 606698
rect 136938 603654 137262 603676
rect 136938 603418 136982 603654
rect 137218 603418 137262 603654
rect 136938 603334 137262 603418
rect 136938 603098 136982 603334
rect 137218 603098 137262 603334
rect 136938 603076 137262 603098
rect 136938 600054 137262 600076
rect 136938 599818 136982 600054
rect 137218 599818 137262 600054
rect 136938 599734 137262 599818
rect 136938 599498 136982 599734
rect 137218 599498 137262 599734
rect 136938 599476 137262 599498
rect 54804 596218 54986 596454
rect 55222 596218 55404 596454
rect 54804 596134 55404 596218
rect 54804 595898 54986 596134
rect 55222 595898 55404 596134
rect 54804 560454 55404 595898
rect 136938 596454 137262 596476
rect 136938 596218 136982 596454
rect 137218 596218 137262 596454
rect 136938 596134 137262 596218
rect 136938 595898 136982 596134
rect 137218 595898 137262 596134
rect 136938 595876 137262 595898
rect 136494 589254 136814 589276
rect 136494 589018 136536 589254
rect 136772 589018 136814 589254
rect 136494 588934 136814 589018
rect 136494 588698 136536 588934
rect 136772 588698 136814 588934
rect 136494 588676 136814 588698
rect 136494 585654 136814 585676
rect 136494 585418 136536 585654
rect 136772 585418 136814 585654
rect 136494 585334 136814 585418
rect 136494 585098 136536 585334
rect 136772 585098 136814 585334
rect 136494 585076 136814 585098
rect 136494 582054 136814 582076
rect 136494 581818 136536 582054
rect 136772 581818 136814 582054
rect 136494 581734 136814 581818
rect 136494 581498 136536 581734
rect 136772 581498 136814 581734
rect 136494 581476 136814 581498
rect 136494 578454 136814 578476
rect 136494 578218 136536 578454
rect 136772 578218 136814 578454
rect 136494 578134 136814 578218
rect 136494 577898 136536 578134
rect 136772 577898 136814 578134
rect 136494 577876 136814 577898
rect 144804 578454 145404 613898
rect 144804 578218 144986 578454
rect 145222 578218 145404 578454
rect 144804 578134 145404 578218
rect 144804 577898 144986 578134
rect 145222 577898 145404 578134
rect 136938 571254 137262 571276
rect 136938 571018 136982 571254
rect 137218 571018 137262 571254
rect 136938 570934 137262 571018
rect 136938 570698 136982 570934
rect 137218 570698 137262 570934
rect 136938 570676 137262 570698
rect 136938 567654 137262 567676
rect 136938 567418 136982 567654
rect 137218 567418 137262 567654
rect 136938 567334 137262 567418
rect 136938 567098 136982 567334
rect 137218 567098 137262 567334
rect 136938 567076 137262 567098
rect 136938 564054 137262 564076
rect 136938 563818 136982 564054
rect 137218 563818 137262 564054
rect 136938 563734 137262 563818
rect 136938 563498 136982 563734
rect 137218 563498 137262 563734
rect 136938 563476 137262 563498
rect 54804 560218 54986 560454
rect 55222 560218 55404 560454
rect 72374 560430 72672 560490
rect 79366 560430 79680 560490
rect 82862 560430 83184 560490
rect 86358 560430 86688 560490
rect 102734 560430 103040 560490
rect 106230 560430 106544 560490
rect 63833 560290 64338 560350
rect 66832 560290 67466 560350
rect 68000 560290 68570 560350
rect 69168 560290 69858 560350
rect 54804 560134 55404 560218
rect 54804 559898 54986 560134
rect 55222 559898 55404 560134
rect 54804 524454 55404 559898
rect 64278 558789 64338 560290
rect 67406 558925 67466 560290
rect 68510 558925 68570 560290
rect 67403 558924 67469 558925
rect 67403 558860 67404 558924
rect 67468 558860 67469 558924
rect 67403 558859 67469 558860
rect 68507 558924 68573 558925
rect 68507 558860 68508 558924
rect 68572 558860 68573 558924
rect 68507 558859 68573 558860
rect 64275 558788 64341 558789
rect 64275 558724 64276 558788
rect 64340 558724 64341 558788
rect 64275 558723 64341 558724
rect 69798 558653 69858 560290
rect 70166 560290 70336 560350
rect 71504 560290 71698 560350
rect 70166 558925 70226 560290
rect 71638 558925 71698 560290
rect 72374 558925 72434 560430
rect 72796 560290 72986 560350
rect 72926 558925 72986 560290
rect 73662 560290 73840 560350
rect 73964 560290 74274 560350
rect 73662 558925 73722 560290
rect 74214 558925 74274 560290
rect 74950 558925 75010 560350
rect 75132 560290 75746 560350
rect 75686 558925 75746 560290
rect 75870 560290 76176 560350
rect 76300 560290 76850 560350
rect 70163 558924 70229 558925
rect 70163 558860 70164 558924
rect 70228 558860 70229 558924
rect 70163 558859 70229 558860
rect 71635 558924 71701 558925
rect 71635 558860 71636 558924
rect 71700 558860 71701 558924
rect 71635 558859 71701 558860
rect 72371 558924 72437 558925
rect 72371 558860 72372 558924
rect 72436 558860 72437 558924
rect 72371 558859 72437 558860
rect 72923 558924 72989 558925
rect 72923 558860 72924 558924
rect 72988 558860 72989 558924
rect 72923 558859 72989 558860
rect 73659 558924 73725 558925
rect 73659 558860 73660 558924
rect 73724 558860 73725 558924
rect 73659 558859 73725 558860
rect 74211 558924 74277 558925
rect 74211 558860 74212 558924
rect 74276 558860 74277 558924
rect 74211 558859 74277 558860
rect 74947 558924 75013 558925
rect 74947 558860 74948 558924
rect 75012 558860 75013 558924
rect 74947 558859 75013 558860
rect 75683 558924 75749 558925
rect 75683 558860 75684 558924
rect 75748 558860 75749 558924
rect 75683 558859 75749 558860
rect 75870 558653 75930 560290
rect 76790 558925 76850 560290
rect 77314 559330 77374 560320
rect 77468 560290 78138 560350
rect 77314 559270 77402 559330
rect 77342 558925 77402 559270
rect 78078 558925 78138 560290
rect 78446 560290 78512 560350
rect 78636 560290 79242 560350
rect 76787 558924 76853 558925
rect 76787 558860 76788 558924
rect 76852 558860 76853 558924
rect 76787 558859 76853 558860
rect 77339 558924 77405 558925
rect 77339 558860 77340 558924
rect 77404 558860 77405 558924
rect 77339 558859 77405 558860
rect 78075 558924 78141 558925
rect 78075 558860 78076 558924
rect 78140 558860 78141 558924
rect 78075 558859 78141 558860
rect 78446 558653 78506 560290
rect 79182 558925 79242 560290
rect 79179 558924 79245 558925
rect 79179 558860 79180 558924
rect 79244 558860 79245 558924
rect 79179 558859 79245 558860
rect 79366 558653 79426 560430
rect 79804 560290 79978 560350
rect 79918 558925 79978 560290
rect 80654 560290 80848 560350
rect 80972 560290 81266 560350
rect 80654 558925 80714 560290
rect 81206 558925 81266 560290
rect 81942 560290 82016 560350
rect 82140 560290 82738 560350
rect 81942 558925 82002 560290
rect 79915 558924 79981 558925
rect 79915 558860 79916 558924
rect 79980 558860 79981 558924
rect 79915 558859 79981 558860
rect 80651 558924 80717 558925
rect 80651 558860 80652 558924
rect 80716 558860 80717 558924
rect 80651 558859 80717 558860
rect 81203 558924 81269 558925
rect 81203 558860 81204 558924
rect 81268 558860 81269 558924
rect 81203 558859 81269 558860
rect 81939 558924 82005 558925
rect 81939 558860 81940 558924
rect 82004 558860 82005 558924
rect 81939 558859 82005 558860
rect 69795 558652 69861 558653
rect 69795 558588 69796 558652
rect 69860 558588 69861 558652
rect 69795 558587 69861 558588
rect 75867 558652 75933 558653
rect 75867 558588 75868 558652
rect 75932 558588 75933 558652
rect 75867 558587 75933 558588
rect 78443 558652 78509 558653
rect 78443 558588 78444 558652
rect 78508 558588 78509 558652
rect 78443 558587 78509 558588
rect 79363 558652 79429 558653
rect 79363 558588 79364 558652
rect 79428 558588 79429 558652
rect 79363 558587 79429 558588
rect 82678 557973 82738 560290
rect 82862 558925 82922 560430
rect 83308 560290 83842 560350
rect 83782 558925 83842 560290
rect 84150 560290 84352 560350
rect 84476 560290 85130 560350
rect 84150 558925 84210 560290
rect 85070 558925 85130 560290
rect 85438 560290 85520 560350
rect 85644 560290 86234 560350
rect 82859 558924 82925 558925
rect 82859 558860 82860 558924
rect 82924 558860 82925 558924
rect 82859 558859 82925 558860
rect 83779 558924 83845 558925
rect 83779 558860 83780 558924
rect 83844 558860 83845 558924
rect 83779 558859 83845 558860
rect 84147 558924 84213 558925
rect 84147 558860 84148 558924
rect 84212 558860 84213 558924
rect 84147 558859 84213 558860
rect 85067 558924 85133 558925
rect 85067 558860 85068 558924
rect 85132 558860 85133 558924
rect 85067 558859 85133 558860
rect 85438 558653 85498 560290
rect 86174 558653 86234 560290
rect 86358 558925 86418 560430
rect 86782 559330 86842 560320
rect 87826 560010 87886 560320
rect 87980 560290 88258 560350
rect 87826 559950 87890 560010
rect 86726 559270 86842 559330
rect 86726 558925 86786 559270
rect 87830 558925 87890 559950
rect 88198 558925 88258 560290
rect 88934 560290 89024 560350
rect 88934 558925 88994 560290
rect 89118 558925 89178 560320
rect 89854 560290 90192 560350
rect 90316 560290 91018 560350
rect 89854 558925 89914 560290
rect 90958 558925 91018 560290
rect 91142 560290 91360 560350
rect 91484 560290 91938 560350
rect 86355 558924 86421 558925
rect 86355 558860 86356 558924
rect 86420 558860 86421 558924
rect 86355 558859 86421 558860
rect 86723 558924 86789 558925
rect 86723 558860 86724 558924
rect 86788 558860 86789 558924
rect 86723 558859 86789 558860
rect 87827 558924 87893 558925
rect 87827 558860 87828 558924
rect 87892 558860 87893 558924
rect 87827 558859 87893 558860
rect 88195 558924 88261 558925
rect 88195 558860 88196 558924
rect 88260 558860 88261 558924
rect 88195 558859 88261 558860
rect 88931 558924 88997 558925
rect 88931 558860 88932 558924
rect 88996 558860 88997 558924
rect 88931 558859 88997 558860
rect 89115 558924 89181 558925
rect 89115 558860 89116 558924
rect 89180 558860 89181 558924
rect 89115 558859 89181 558860
rect 89851 558924 89917 558925
rect 89851 558860 89852 558924
rect 89916 558860 89917 558924
rect 89851 558859 89917 558860
rect 90955 558924 91021 558925
rect 90955 558860 90956 558924
rect 91020 558860 91021 558924
rect 90955 558859 91021 558860
rect 91142 558653 91202 560290
rect 91878 558925 91938 560290
rect 92498 560010 92558 560320
rect 92652 560290 93226 560350
rect 92430 559950 92558 560010
rect 92430 558925 92490 559950
rect 91875 558924 91941 558925
rect 91875 558860 91876 558924
rect 91940 558860 91941 558924
rect 91875 558859 91941 558860
rect 92427 558924 92493 558925
rect 92427 558860 92428 558924
rect 92492 558860 92493 558924
rect 92427 558859 92493 558860
rect 93166 558653 93226 560290
rect 93350 560290 93696 560350
rect 93350 558925 93410 560290
rect 93790 559330 93850 560320
rect 93718 559270 93850 559330
rect 93718 558925 93778 559270
rect 93347 558924 93413 558925
rect 93347 558860 93348 558924
rect 93412 558860 93413 558924
rect 93347 558859 93413 558860
rect 93715 558924 93781 558925
rect 93715 558860 93716 558924
rect 93780 558860 93781 558924
rect 93715 558859 93781 558860
rect 94822 558653 94882 560350
rect 94988 560290 95066 560350
rect 95006 558925 95066 560290
rect 95742 560290 96032 560350
rect 96156 560290 96538 560350
rect 95742 558925 95802 560290
rect 96478 558925 96538 560290
rect 97030 560290 97200 560350
rect 97324 560290 97826 560350
rect 97030 558925 97090 560290
rect 97766 558925 97826 560290
rect 98318 558925 98378 560350
rect 98492 560290 99114 560350
rect 99054 558925 99114 560290
rect 99506 559330 99566 560320
rect 99660 560290 100034 560350
rect 99506 559270 99666 559330
rect 95003 558924 95069 558925
rect 95003 558860 95004 558924
rect 95068 558860 95069 558924
rect 95003 558859 95069 558860
rect 95739 558924 95805 558925
rect 95739 558860 95740 558924
rect 95804 558860 95805 558924
rect 95739 558859 95805 558860
rect 96475 558924 96541 558925
rect 96475 558860 96476 558924
rect 96540 558860 96541 558924
rect 96475 558859 96541 558860
rect 97027 558924 97093 558925
rect 97027 558860 97028 558924
rect 97092 558860 97093 558924
rect 97027 558859 97093 558860
rect 97763 558924 97829 558925
rect 97763 558860 97764 558924
rect 97828 558860 97829 558924
rect 97763 558859 97829 558860
rect 98315 558924 98381 558925
rect 98315 558860 98316 558924
rect 98380 558860 98381 558924
rect 98315 558859 98381 558860
rect 99051 558924 99117 558925
rect 99051 558860 99052 558924
rect 99116 558860 99117 558924
rect 99051 558859 99117 558860
rect 85435 558652 85501 558653
rect 85435 558588 85436 558652
rect 85500 558588 85501 558652
rect 85435 558587 85501 558588
rect 86171 558652 86237 558653
rect 86171 558588 86172 558652
rect 86236 558588 86237 558652
rect 86171 558587 86237 558588
rect 91139 558652 91205 558653
rect 91139 558588 91140 558652
rect 91204 558588 91205 558652
rect 91139 558587 91205 558588
rect 93163 558652 93229 558653
rect 93163 558588 93164 558652
rect 93228 558588 93229 558652
rect 93163 558587 93229 558588
rect 94819 558652 94885 558653
rect 94819 558588 94820 558652
rect 94884 558588 94885 558652
rect 94819 558587 94885 558588
rect 99606 558517 99666 559270
rect 99974 558925 100034 560290
rect 100158 560290 100704 560350
rect 100828 560290 101506 560350
rect 99971 558924 100037 558925
rect 99971 558860 99972 558924
rect 100036 558860 100037 558924
rect 99971 558859 100037 558860
rect 99603 558516 99669 558517
rect 99603 558452 99604 558516
rect 99668 558452 99669 558516
rect 99603 558451 99669 558452
rect 82675 557972 82741 557973
rect 82675 557908 82676 557972
rect 82740 557908 82741 557972
rect 82675 557907 82741 557908
rect 100158 557701 100218 560290
rect 100155 557700 100221 557701
rect 100155 557636 100156 557700
rect 100220 557636 100221 557700
rect 100155 557635 100221 557636
rect 101446 557565 101506 560290
rect 101630 560290 101872 560350
rect 101996 560290 102058 560350
rect 101630 557837 101690 560290
rect 101998 558925 102058 560290
rect 101995 558924 102061 558925
rect 101995 558860 101996 558924
rect 102060 558860 102061 558924
rect 101995 558859 102061 558860
rect 101627 557836 101693 557837
rect 101627 557772 101628 557836
rect 101692 557772 101693 557836
rect 101627 557771 101693 557772
rect 102734 557565 102794 560430
rect 103164 560290 103346 560350
rect 103286 557565 103346 560290
rect 104022 560290 104208 560350
rect 104332 560290 104818 560350
rect 104022 557565 104082 560290
rect 104758 558925 104818 560290
rect 105310 560290 105376 560350
rect 105500 560290 106106 560350
rect 104755 558924 104821 558925
rect 104755 558860 104756 558924
rect 104820 558860 104821 558924
rect 104755 558859 104821 558860
rect 105310 557565 105370 560290
rect 106046 557565 106106 560290
rect 106230 558653 106290 560430
rect 106668 560290 107210 560350
rect 107150 558925 107210 560290
rect 107682 559330 107742 560320
rect 107836 560290 108498 560350
rect 107682 559270 107762 559330
rect 107147 558924 107213 558925
rect 107147 558860 107148 558924
rect 107212 558860 107213 558924
rect 107147 558859 107213 558860
rect 106227 558652 106293 558653
rect 106227 558588 106228 558652
rect 106292 558588 106293 558652
rect 106227 558587 106293 558588
rect 106230 557701 106290 558587
rect 107702 557973 107762 559270
rect 108438 558925 108498 560290
rect 108622 560290 108880 560350
rect 108435 558924 108501 558925
rect 108435 558860 108436 558924
rect 108500 558860 108501 558924
rect 108435 558859 108501 558860
rect 108622 558517 108682 560290
rect 108990 558517 109050 560350
rect 108619 558516 108685 558517
rect 108619 558452 108620 558516
rect 108684 558452 108685 558516
rect 108619 558451 108685 558452
rect 108987 558516 109053 558517
rect 108987 558452 108988 558516
rect 109052 558452 109053 558516
rect 108987 558451 109053 558452
rect 107699 557972 107765 557973
rect 107699 557908 107700 557972
rect 107764 557908 107765 557972
rect 107699 557907 107765 557908
rect 106227 557700 106293 557701
rect 106227 557636 106228 557700
rect 106292 557636 106293 557700
rect 106227 557635 106293 557636
rect 101443 557564 101509 557565
rect 101443 557500 101444 557564
rect 101508 557500 101509 557564
rect 101443 557499 101509 557500
rect 102731 557564 102797 557565
rect 102731 557500 102732 557564
rect 102796 557500 102797 557564
rect 102731 557499 102797 557500
rect 103283 557564 103349 557565
rect 103283 557500 103284 557564
rect 103348 557500 103349 557564
rect 103283 557499 103349 557500
rect 104019 557564 104085 557565
rect 104019 557500 104020 557564
rect 104084 557500 104085 557564
rect 104019 557499 104085 557500
rect 105307 557564 105373 557565
rect 105307 557500 105308 557564
rect 105372 557500 105373 557564
rect 105307 557499 105373 557500
rect 106043 557564 106109 557565
rect 106043 557500 106044 557564
rect 106108 557500 106109 557564
rect 106043 557499 106109 557500
rect 58404 543000 59004 557000
rect 62004 543000 62604 557000
rect 65604 543000 66204 557000
rect 72804 543000 73404 557000
rect 76404 546054 77004 557000
rect 76404 545818 76586 546054
rect 76822 545818 77004 546054
rect 76404 545734 77004 545818
rect 76404 545498 76586 545734
rect 76822 545498 77004 545734
rect 76404 543000 77004 545498
rect 80004 549654 80604 557000
rect 80004 549418 80186 549654
rect 80422 549418 80604 549654
rect 80004 549334 80604 549418
rect 80004 549098 80186 549334
rect 80422 549098 80604 549334
rect 80004 543000 80604 549098
rect 83604 553254 84204 557000
rect 83604 553018 83786 553254
rect 84022 553018 84204 553254
rect 83604 552934 84204 553018
rect 83604 552698 83786 552934
rect 84022 552698 84204 552934
rect 83604 543000 84204 552698
rect 90804 543000 91404 557000
rect 94404 543000 95004 557000
rect 98004 543000 98604 557000
rect 101604 543000 102204 557000
rect 108804 543000 109404 557000
rect 112404 546054 113004 557000
rect 112404 545818 112586 546054
rect 112822 545818 113004 546054
rect 112404 545734 113004 545818
rect 112404 545498 112586 545734
rect 112822 545498 113004 545734
rect 112404 543000 113004 545498
rect 116004 549654 116604 557000
rect 116004 549418 116186 549654
rect 116422 549418 116604 549654
rect 116004 549334 116604 549418
rect 116004 549098 116186 549334
rect 116422 549098 116604 549334
rect 116004 543000 116604 549098
rect 119604 553254 120204 557000
rect 119604 553018 119786 553254
rect 120022 553018 120204 553254
rect 119604 552934 120204 553018
rect 119604 552698 119786 552934
rect 120022 552698 120204 552934
rect 119604 543000 120204 552698
rect 126804 543000 127404 557000
rect 130404 543000 131004 557000
rect 134004 543000 134604 557000
rect 137604 543000 138204 557000
rect 144804 543000 145404 577898
rect 148404 690054 149004 706162
rect 148404 689818 148586 690054
rect 148822 689818 149004 690054
rect 148404 689734 149004 689818
rect 148404 689498 148586 689734
rect 148822 689498 149004 689734
rect 148404 654054 149004 689498
rect 148404 653818 148586 654054
rect 148822 653818 149004 654054
rect 148404 653734 149004 653818
rect 148404 653498 148586 653734
rect 148822 653498 149004 653734
rect 148404 618054 149004 653498
rect 148404 617818 148586 618054
rect 148822 617818 149004 618054
rect 148404 617734 149004 617818
rect 148404 617498 148586 617734
rect 148822 617498 149004 617734
rect 148404 582054 149004 617498
rect 148404 581818 148586 582054
rect 148822 581818 149004 582054
rect 148404 581734 149004 581818
rect 148404 581498 148586 581734
rect 148822 581498 149004 581734
rect 148404 546054 149004 581498
rect 148404 545818 148586 546054
rect 148822 545818 149004 546054
rect 148404 545734 149004 545818
rect 148404 545498 148586 545734
rect 148822 545498 149004 545734
rect 148404 543000 149004 545498
rect 152004 693654 152604 708042
rect 152004 693418 152186 693654
rect 152422 693418 152604 693654
rect 152004 693334 152604 693418
rect 152004 693098 152186 693334
rect 152422 693098 152604 693334
rect 152004 657654 152604 693098
rect 152004 657418 152186 657654
rect 152422 657418 152604 657654
rect 152004 657334 152604 657418
rect 152004 657098 152186 657334
rect 152422 657098 152604 657334
rect 152004 621654 152604 657098
rect 152004 621418 152186 621654
rect 152422 621418 152604 621654
rect 152004 621334 152604 621418
rect 152004 621098 152186 621334
rect 152422 621098 152604 621334
rect 152004 585654 152604 621098
rect 152004 585418 152186 585654
rect 152422 585418 152604 585654
rect 152004 585334 152604 585418
rect 152004 585098 152186 585334
rect 152422 585098 152604 585334
rect 152004 549654 152604 585098
rect 152004 549418 152186 549654
rect 152422 549418 152604 549654
rect 152004 549334 152604 549418
rect 152004 549098 152186 549334
rect 152422 549098 152604 549334
rect 152004 543000 152604 549098
rect 155604 697254 156204 709922
rect 173604 711418 174204 711440
rect 173604 711182 173786 711418
rect 174022 711182 174204 711418
rect 173604 711098 174204 711182
rect 173604 710862 173786 711098
rect 174022 710862 174204 711098
rect 170004 709538 170604 709560
rect 170004 709302 170186 709538
rect 170422 709302 170604 709538
rect 170004 709218 170604 709302
rect 170004 708982 170186 709218
rect 170422 708982 170604 709218
rect 166404 707658 167004 707680
rect 166404 707422 166586 707658
rect 166822 707422 167004 707658
rect 166404 707338 167004 707422
rect 166404 707102 166586 707338
rect 166822 707102 167004 707338
rect 155604 697018 155786 697254
rect 156022 697018 156204 697254
rect 155604 696934 156204 697018
rect 155604 696698 155786 696934
rect 156022 696698 156204 696934
rect 155604 661254 156204 696698
rect 155604 661018 155786 661254
rect 156022 661018 156204 661254
rect 155604 660934 156204 661018
rect 155604 660698 155786 660934
rect 156022 660698 156204 660934
rect 155604 625254 156204 660698
rect 155604 625018 155786 625254
rect 156022 625018 156204 625254
rect 155604 624934 156204 625018
rect 155604 624698 155786 624934
rect 156022 624698 156204 624934
rect 155604 589254 156204 624698
rect 155604 589018 155786 589254
rect 156022 589018 156204 589254
rect 155604 588934 156204 589018
rect 155604 588698 155786 588934
rect 156022 588698 156204 588934
rect 155604 553254 156204 588698
rect 155604 553018 155786 553254
rect 156022 553018 156204 553254
rect 155604 552934 156204 553018
rect 155604 552698 155786 552934
rect 156022 552698 156204 552934
rect 155604 543000 156204 552698
rect 162804 705778 163404 705800
rect 162804 705542 162986 705778
rect 163222 705542 163404 705778
rect 162804 705458 163404 705542
rect 162804 705222 162986 705458
rect 163222 705222 163404 705458
rect 162804 668454 163404 705222
rect 162804 668218 162986 668454
rect 163222 668218 163404 668454
rect 162804 668134 163404 668218
rect 162804 667898 162986 668134
rect 163222 667898 163404 668134
rect 162804 632454 163404 667898
rect 162804 632218 162986 632454
rect 163222 632218 163404 632454
rect 162804 632134 163404 632218
rect 162804 631898 162986 632134
rect 163222 631898 163404 632134
rect 162804 596454 163404 631898
rect 162804 596218 162986 596454
rect 163222 596218 163404 596454
rect 162804 596134 163404 596218
rect 162804 595898 162986 596134
rect 163222 595898 163404 596134
rect 162804 560454 163404 595898
rect 162804 560218 162986 560454
rect 163222 560218 163404 560454
rect 162804 560134 163404 560218
rect 162804 559898 162986 560134
rect 163222 559898 163404 560134
rect 162804 543000 163404 559898
rect 166404 672054 167004 707102
rect 166404 671818 166586 672054
rect 166822 671818 167004 672054
rect 166404 671734 167004 671818
rect 166404 671498 166586 671734
rect 166822 671498 167004 671734
rect 166404 636054 167004 671498
rect 166404 635818 166586 636054
rect 166822 635818 167004 636054
rect 166404 635734 167004 635818
rect 166404 635498 166586 635734
rect 166822 635498 167004 635734
rect 166404 600054 167004 635498
rect 166404 599818 166586 600054
rect 166822 599818 167004 600054
rect 166404 599734 167004 599818
rect 166404 599498 166586 599734
rect 166822 599498 167004 599734
rect 166404 564054 167004 599498
rect 166404 563818 166586 564054
rect 166822 563818 167004 564054
rect 166404 563734 167004 563818
rect 166404 563498 166586 563734
rect 166822 563498 167004 563734
rect 166404 543000 167004 563498
rect 170004 675654 170604 708982
rect 170004 675418 170186 675654
rect 170422 675418 170604 675654
rect 170004 675334 170604 675418
rect 170004 675098 170186 675334
rect 170422 675098 170604 675334
rect 170004 639654 170604 675098
rect 170004 639418 170186 639654
rect 170422 639418 170604 639654
rect 170004 639334 170604 639418
rect 170004 639098 170186 639334
rect 170422 639098 170604 639334
rect 170004 603654 170604 639098
rect 170004 603418 170186 603654
rect 170422 603418 170604 603654
rect 170004 603334 170604 603418
rect 170004 603098 170186 603334
rect 170422 603098 170604 603334
rect 170004 567654 170604 603098
rect 170004 567418 170186 567654
rect 170422 567418 170604 567654
rect 170004 567334 170604 567418
rect 170004 567098 170186 567334
rect 170422 567098 170604 567334
rect 170004 543000 170604 567098
rect 173604 679254 174204 710862
rect 191604 710478 192204 711440
rect 191604 710242 191786 710478
rect 192022 710242 192204 710478
rect 191604 710158 192204 710242
rect 191604 709922 191786 710158
rect 192022 709922 192204 710158
rect 188004 708598 188604 709560
rect 188004 708362 188186 708598
rect 188422 708362 188604 708598
rect 188004 708278 188604 708362
rect 188004 708042 188186 708278
rect 188422 708042 188604 708278
rect 184404 706718 185004 707680
rect 184404 706482 184586 706718
rect 184822 706482 185004 706718
rect 184404 706398 185004 706482
rect 184404 706162 184586 706398
rect 184822 706162 185004 706398
rect 173604 679018 173786 679254
rect 174022 679018 174204 679254
rect 173604 678934 174204 679018
rect 173604 678698 173786 678934
rect 174022 678698 174204 678934
rect 173604 643254 174204 678698
rect 173604 643018 173786 643254
rect 174022 643018 174204 643254
rect 173604 642934 174204 643018
rect 173604 642698 173786 642934
rect 174022 642698 174204 642934
rect 173604 607254 174204 642698
rect 173604 607018 173786 607254
rect 174022 607018 174204 607254
rect 173604 606934 174204 607018
rect 173604 606698 173786 606934
rect 174022 606698 174204 606934
rect 173604 571254 174204 606698
rect 173604 571018 173786 571254
rect 174022 571018 174204 571254
rect 173604 570934 174204 571018
rect 173604 570698 173786 570934
rect 174022 570698 174204 570934
rect 173604 543000 174204 570698
rect 180804 704838 181404 705800
rect 180804 704602 180986 704838
rect 181222 704602 181404 704838
rect 180804 704518 181404 704602
rect 180804 704282 180986 704518
rect 181222 704282 181404 704518
rect 180804 686454 181404 704282
rect 180804 686218 180986 686454
rect 181222 686218 181404 686454
rect 180804 686134 181404 686218
rect 180804 685898 180986 686134
rect 181222 685898 181404 686134
rect 180804 650454 181404 685898
rect 180804 650218 180986 650454
rect 181222 650218 181404 650454
rect 180804 650134 181404 650218
rect 180804 649898 180986 650134
rect 181222 649898 181404 650134
rect 180804 614454 181404 649898
rect 180804 614218 180986 614454
rect 181222 614218 181404 614454
rect 180804 614134 181404 614218
rect 180804 613898 180986 614134
rect 181222 613898 181404 614134
rect 180804 578454 181404 613898
rect 180804 578218 180986 578454
rect 181222 578218 181404 578454
rect 180804 578134 181404 578218
rect 180804 577898 180986 578134
rect 181222 577898 181404 578134
rect 180804 543000 181404 577898
rect 184404 690054 185004 706162
rect 184404 689818 184586 690054
rect 184822 689818 185004 690054
rect 184404 689734 185004 689818
rect 184404 689498 184586 689734
rect 184822 689498 185004 689734
rect 184404 654054 185004 689498
rect 188004 693654 188604 708042
rect 188004 693418 188186 693654
rect 188422 693418 188604 693654
rect 188004 693334 188604 693418
rect 188004 693098 188186 693334
rect 188422 693098 188604 693334
rect 188004 657654 188604 693098
rect 188004 657418 188186 657654
rect 188422 657418 188604 657654
rect 188004 657334 188604 657418
rect 188004 657098 188186 657334
rect 188422 657098 188604 657334
rect 188004 654247 188604 657098
rect 191604 697254 192204 709922
rect 209604 711418 210204 711440
rect 209604 711182 209786 711418
rect 210022 711182 210204 711418
rect 209604 711098 210204 711182
rect 209604 710862 209786 711098
rect 210022 710862 210204 711098
rect 206004 709538 206604 709560
rect 206004 709302 206186 709538
rect 206422 709302 206604 709538
rect 206004 709218 206604 709302
rect 206004 708982 206186 709218
rect 206422 708982 206604 709218
rect 202404 707658 203004 707680
rect 202404 707422 202586 707658
rect 202822 707422 203004 707658
rect 202404 707338 203004 707422
rect 202404 707102 202586 707338
rect 202822 707102 203004 707338
rect 191604 697018 191786 697254
rect 192022 697018 192204 697254
rect 191604 696934 192204 697018
rect 191604 696698 191786 696934
rect 192022 696698 192204 696934
rect 191604 661254 192204 696698
rect 191604 661018 191786 661254
rect 192022 661018 192204 661254
rect 191604 660934 192204 661018
rect 191604 660698 191786 660934
rect 192022 660698 192204 660934
rect 191604 654247 192204 660698
rect 198804 705778 199404 705800
rect 198804 705542 198986 705778
rect 199222 705542 199404 705778
rect 198804 705458 199404 705542
rect 198804 705222 198986 705458
rect 199222 705222 199404 705458
rect 198804 668454 199404 705222
rect 198804 668218 198986 668454
rect 199222 668218 199404 668454
rect 198804 668134 199404 668218
rect 198804 667898 198986 668134
rect 199222 667898 199404 668134
rect 198804 654247 199404 667898
rect 202404 672054 203004 707102
rect 202404 671818 202586 672054
rect 202822 671818 203004 672054
rect 202404 671734 203004 671818
rect 202404 671498 202586 671734
rect 202822 671498 203004 671734
rect 202404 654247 203004 671498
rect 206004 675654 206604 708982
rect 206004 675418 206186 675654
rect 206422 675418 206604 675654
rect 206004 675334 206604 675418
rect 206004 675098 206186 675334
rect 206422 675098 206604 675334
rect 206004 654247 206604 675098
rect 209604 679254 210204 710862
rect 227604 710478 228204 711440
rect 227604 710242 227786 710478
rect 228022 710242 228204 710478
rect 227604 710158 228204 710242
rect 227604 709922 227786 710158
rect 228022 709922 228204 710158
rect 224004 708598 224604 709560
rect 224004 708362 224186 708598
rect 224422 708362 224604 708598
rect 224004 708278 224604 708362
rect 224004 708042 224186 708278
rect 224422 708042 224604 708278
rect 220404 706718 221004 707680
rect 220404 706482 220586 706718
rect 220822 706482 221004 706718
rect 220404 706398 221004 706482
rect 220404 706162 220586 706398
rect 220822 706162 221004 706398
rect 209604 679018 209786 679254
rect 210022 679018 210204 679254
rect 209604 678934 210204 679018
rect 209604 678698 209786 678934
rect 210022 678698 210204 678934
rect 209604 654247 210204 678698
rect 216804 704838 217404 705800
rect 216804 704602 216986 704838
rect 217222 704602 217404 704838
rect 216804 704518 217404 704602
rect 216804 704282 216986 704518
rect 217222 704282 217404 704518
rect 216804 686454 217404 704282
rect 216804 686218 216986 686454
rect 217222 686218 217404 686454
rect 216804 686134 217404 686218
rect 216804 685898 216986 686134
rect 217222 685898 217404 686134
rect 216804 654247 217404 685898
rect 220404 690054 221004 706162
rect 220404 689818 220586 690054
rect 220822 689818 221004 690054
rect 220404 689734 221004 689818
rect 220404 689498 220586 689734
rect 220822 689498 221004 689734
rect 220404 654247 221004 689498
rect 224004 693654 224604 708042
rect 224004 693418 224186 693654
rect 224422 693418 224604 693654
rect 224004 693334 224604 693418
rect 224004 693098 224186 693334
rect 224422 693098 224604 693334
rect 224004 657654 224604 693098
rect 224004 657418 224186 657654
rect 224422 657418 224604 657654
rect 224004 657334 224604 657418
rect 224004 657098 224186 657334
rect 224422 657098 224604 657334
rect 224004 654247 224604 657098
rect 227604 697254 228204 709922
rect 245604 711418 246204 711440
rect 245604 711182 245786 711418
rect 246022 711182 246204 711418
rect 245604 711098 246204 711182
rect 245604 710862 245786 711098
rect 246022 710862 246204 711098
rect 242004 709538 242604 709560
rect 242004 709302 242186 709538
rect 242422 709302 242604 709538
rect 242004 709218 242604 709302
rect 242004 708982 242186 709218
rect 242422 708982 242604 709218
rect 238404 707658 239004 707680
rect 238404 707422 238586 707658
rect 238822 707422 239004 707658
rect 238404 707338 239004 707422
rect 238404 707102 238586 707338
rect 238822 707102 239004 707338
rect 227604 697018 227786 697254
rect 228022 697018 228204 697254
rect 227604 696934 228204 697018
rect 227604 696698 227786 696934
rect 228022 696698 228204 696934
rect 227604 661254 228204 696698
rect 227604 661018 227786 661254
rect 228022 661018 228204 661254
rect 227604 660934 228204 661018
rect 227604 660698 227786 660934
rect 228022 660698 228204 660934
rect 227604 654247 228204 660698
rect 234804 705778 235404 705800
rect 234804 705542 234986 705778
rect 235222 705542 235404 705778
rect 234804 705458 235404 705542
rect 234804 705222 234986 705458
rect 235222 705222 235404 705458
rect 234804 668454 235404 705222
rect 234804 668218 234986 668454
rect 235222 668218 235404 668454
rect 234804 668134 235404 668218
rect 234804 667898 234986 668134
rect 235222 667898 235404 668134
rect 234804 654247 235404 667898
rect 238404 672054 239004 707102
rect 238404 671818 238586 672054
rect 238822 671818 239004 672054
rect 238404 671734 239004 671818
rect 238404 671498 238586 671734
rect 238822 671498 239004 671734
rect 238404 654247 239004 671498
rect 242004 675654 242604 708982
rect 242004 675418 242186 675654
rect 242422 675418 242604 675654
rect 242004 675334 242604 675418
rect 242004 675098 242186 675334
rect 242422 675098 242604 675334
rect 242004 654247 242604 675098
rect 245604 679254 246204 710862
rect 263604 710478 264204 711440
rect 263604 710242 263786 710478
rect 264022 710242 264204 710478
rect 263604 710158 264204 710242
rect 263604 709922 263786 710158
rect 264022 709922 264204 710158
rect 260004 708598 260604 709560
rect 260004 708362 260186 708598
rect 260422 708362 260604 708598
rect 260004 708278 260604 708362
rect 260004 708042 260186 708278
rect 260422 708042 260604 708278
rect 256404 706718 257004 707680
rect 256404 706482 256586 706718
rect 256822 706482 257004 706718
rect 256404 706398 257004 706482
rect 256404 706162 256586 706398
rect 256822 706162 257004 706398
rect 245604 679018 245786 679254
rect 246022 679018 246204 679254
rect 245604 678934 246204 679018
rect 245604 678698 245786 678934
rect 246022 678698 246204 678934
rect 245604 654247 246204 678698
rect 252804 704838 253404 705800
rect 252804 704602 252986 704838
rect 253222 704602 253404 704838
rect 252804 704518 253404 704602
rect 252804 704282 252986 704518
rect 253222 704282 253404 704518
rect 252804 686454 253404 704282
rect 252804 686218 252986 686454
rect 253222 686218 253404 686454
rect 252804 686134 253404 686218
rect 252804 685898 252986 686134
rect 253222 685898 253404 686134
rect 252804 654247 253404 685898
rect 256404 690054 257004 706162
rect 256404 689818 256586 690054
rect 256822 689818 257004 690054
rect 256404 689734 257004 689818
rect 256404 689498 256586 689734
rect 256822 689498 257004 689734
rect 256404 654247 257004 689498
rect 260004 693654 260604 708042
rect 260004 693418 260186 693654
rect 260422 693418 260604 693654
rect 260004 693334 260604 693418
rect 260004 693098 260186 693334
rect 260422 693098 260604 693334
rect 260004 657654 260604 693098
rect 260004 657418 260186 657654
rect 260422 657418 260604 657654
rect 260004 657334 260604 657418
rect 260004 657098 260186 657334
rect 260422 657098 260604 657334
rect 260004 654247 260604 657098
rect 263604 697254 264204 709922
rect 281604 711418 282204 711440
rect 281604 711182 281786 711418
rect 282022 711182 282204 711418
rect 281604 711098 282204 711182
rect 281604 710862 281786 711098
rect 282022 710862 282204 711098
rect 278004 709538 278604 709560
rect 278004 709302 278186 709538
rect 278422 709302 278604 709538
rect 278004 709218 278604 709302
rect 278004 708982 278186 709218
rect 278422 708982 278604 709218
rect 274404 707658 275004 707680
rect 274404 707422 274586 707658
rect 274822 707422 275004 707658
rect 274404 707338 275004 707422
rect 274404 707102 274586 707338
rect 274822 707102 275004 707338
rect 263604 697018 263786 697254
rect 264022 697018 264204 697254
rect 263604 696934 264204 697018
rect 263604 696698 263786 696934
rect 264022 696698 264204 696934
rect 263604 661254 264204 696698
rect 263604 661018 263786 661254
rect 264022 661018 264204 661254
rect 263604 660934 264204 661018
rect 263604 660698 263786 660934
rect 264022 660698 264204 660934
rect 263604 654247 264204 660698
rect 270804 705778 271404 705800
rect 270804 705542 270986 705778
rect 271222 705542 271404 705778
rect 270804 705458 271404 705542
rect 270804 705222 270986 705458
rect 271222 705222 271404 705458
rect 270804 668454 271404 705222
rect 270804 668218 270986 668454
rect 271222 668218 271404 668454
rect 270804 668134 271404 668218
rect 270804 667898 270986 668134
rect 271222 667898 271404 668134
rect 184404 653818 184586 654054
rect 184822 653818 185004 654054
rect 184404 653734 185004 653818
rect 184404 653498 184586 653734
rect 184822 653498 185004 653734
rect 184404 618054 185004 653498
rect 258575 651676 258641 651677
rect 258575 651612 258576 651676
rect 258640 651612 258641 651676
rect 258575 651611 258641 651612
rect 263570 651676 263636 651677
rect 263570 651612 263571 651676
rect 263635 651612 263636 651676
rect 263570 651611 263636 651612
rect 258578 651100 258638 651611
rect 263573 651100 263633 651611
rect 266938 643254 267262 643276
rect 266938 643018 266982 643254
rect 267218 643018 267262 643254
rect 266938 642934 267262 643018
rect 266938 642698 266982 642934
rect 267218 642698 267262 642934
rect 266938 642676 267262 642698
rect 266938 639654 267262 639676
rect 266938 639418 266982 639654
rect 267218 639418 267262 639654
rect 266938 639334 267262 639418
rect 266938 639098 266982 639334
rect 267218 639098 267262 639334
rect 266938 639076 267262 639098
rect 266938 636054 267262 636076
rect 266938 635818 266982 636054
rect 267218 635818 267262 636054
rect 266938 635734 267262 635818
rect 266938 635498 266982 635734
rect 267218 635498 267262 635734
rect 266938 635476 267262 635498
rect 266938 632454 267262 632476
rect 266938 632218 266982 632454
rect 267218 632218 267262 632454
rect 266938 632134 267262 632218
rect 266938 631898 266982 632134
rect 267218 631898 267262 632134
rect 266938 631876 267262 631898
rect 270804 632454 271404 667898
rect 270804 632218 270986 632454
rect 271222 632218 271404 632454
rect 270804 632134 271404 632218
rect 270804 631898 270986 632134
rect 271222 631898 271404 632134
rect 266494 625254 266814 625276
rect 266494 625018 266536 625254
rect 266772 625018 266814 625254
rect 266494 624934 266814 625018
rect 266494 624698 266536 624934
rect 266772 624698 266814 624934
rect 266494 624676 266814 624698
rect 266494 621654 266814 621676
rect 266494 621418 266536 621654
rect 266772 621418 266814 621654
rect 266494 621334 266814 621418
rect 266494 621098 266536 621334
rect 266772 621098 266814 621334
rect 266494 621076 266814 621098
rect 184404 617818 184586 618054
rect 184822 617818 185004 618054
rect 184404 617734 185004 617818
rect 184404 617498 184586 617734
rect 184822 617498 185004 617734
rect 184404 582054 185004 617498
rect 266494 618054 266814 618076
rect 266494 617818 266536 618054
rect 266772 617818 266814 618054
rect 266494 617734 266814 617818
rect 266494 617498 266536 617734
rect 266772 617498 266814 617734
rect 266494 617476 266814 617498
rect 266494 614454 266814 614476
rect 266494 614218 266536 614454
rect 266772 614218 266814 614454
rect 266494 614134 266814 614218
rect 266494 613898 266536 614134
rect 266772 613898 266814 614134
rect 266494 613876 266814 613898
rect 266938 607254 267262 607276
rect 266938 607018 266982 607254
rect 267218 607018 267262 607254
rect 266938 606934 267262 607018
rect 266938 606698 266982 606934
rect 267218 606698 267262 606934
rect 266938 606676 267262 606698
rect 266938 603654 267262 603676
rect 266938 603418 266982 603654
rect 267218 603418 267262 603654
rect 266938 603334 267262 603418
rect 266938 603098 266982 603334
rect 267218 603098 267262 603334
rect 266938 603076 267262 603098
rect 266938 600054 267262 600076
rect 266938 599818 266982 600054
rect 267218 599818 267262 600054
rect 266938 599734 267262 599818
rect 266938 599498 266982 599734
rect 267218 599498 267262 599734
rect 266938 599476 267262 599498
rect 266938 596454 267262 596476
rect 266938 596218 266982 596454
rect 267218 596218 267262 596454
rect 266938 596134 267262 596218
rect 266938 595898 266982 596134
rect 267218 595898 267262 596134
rect 266938 595876 267262 595898
rect 270804 596454 271404 631898
rect 270804 596218 270986 596454
rect 271222 596218 271404 596454
rect 270804 596134 271404 596218
rect 270804 595898 270986 596134
rect 271222 595898 271404 596134
rect 266494 589254 266814 589276
rect 266494 589018 266536 589254
rect 266772 589018 266814 589254
rect 266494 588934 266814 589018
rect 266494 588698 266536 588934
rect 266772 588698 266814 588934
rect 266494 588676 266814 588698
rect 266494 585654 266814 585676
rect 266494 585418 266536 585654
rect 266772 585418 266814 585654
rect 266494 585334 266814 585418
rect 266494 585098 266536 585334
rect 266772 585098 266814 585334
rect 266494 585076 266814 585098
rect 184404 581818 184586 582054
rect 184822 581818 185004 582054
rect 184404 581734 185004 581818
rect 184404 581498 184586 581734
rect 184822 581498 185004 581734
rect 184404 546054 185004 581498
rect 266494 582054 266814 582076
rect 266494 581818 266536 582054
rect 266772 581818 266814 582054
rect 266494 581734 266814 581818
rect 266494 581498 266536 581734
rect 266772 581498 266814 581734
rect 266494 581476 266814 581498
rect 266494 578454 266814 578476
rect 266494 578218 266536 578454
rect 266772 578218 266814 578454
rect 266494 578134 266814 578218
rect 266494 577898 266536 578134
rect 266772 577898 266814 578134
rect 266494 577876 266814 577898
rect 266938 571254 267262 571276
rect 266938 571018 266982 571254
rect 267218 571018 267262 571254
rect 266938 570934 267262 571018
rect 266938 570698 266982 570934
rect 267218 570698 267262 570934
rect 266938 570676 267262 570698
rect 266938 567654 267262 567676
rect 266938 567418 266982 567654
rect 267218 567418 267262 567654
rect 266938 567334 267262 567418
rect 266938 567098 266982 567334
rect 267218 567098 267262 567334
rect 266938 567076 267262 567098
rect 266938 564054 267262 564076
rect 266938 563818 266982 564054
rect 267218 563818 267262 564054
rect 266938 563734 267262 563818
rect 266938 563498 266982 563734
rect 267218 563498 267262 563734
rect 266938 563476 267262 563498
rect 207062 560430 207344 560490
rect 214054 560430 214352 560490
rect 217550 560430 217856 560490
rect 221046 560430 221360 560490
rect 228038 560430 228368 560490
rect 270804 560454 271404 595898
rect 193833 560290 194426 560350
rect 194366 558789 194426 560290
rect 196206 560290 196832 560350
rect 197310 560290 198000 560350
rect 198782 560290 199168 560350
rect 200254 560290 200336 560350
rect 196206 558925 196266 560290
rect 196203 558924 196269 558925
rect 196203 558860 196204 558924
rect 196268 558860 196269 558924
rect 196203 558859 196269 558860
rect 194363 558788 194429 558789
rect 194363 558724 194364 558788
rect 194428 558724 194429 558788
rect 194363 558723 194429 558724
rect 197310 558381 197370 560290
rect 197307 558380 197373 558381
rect 197307 558316 197308 558380
rect 197372 558316 197373 558380
rect 197307 558315 197373 558316
rect 198782 558245 198842 560290
rect 200254 558925 200314 560290
rect 201474 560010 201534 560320
rect 202462 560290 202672 560350
rect 201474 559950 201602 560010
rect 200251 558924 200317 558925
rect 200251 558860 200252 558924
rect 200316 558860 200317 558924
rect 200251 558859 200317 558860
rect 198779 558244 198845 558245
rect 198779 558180 198780 558244
rect 198844 558180 198845 558244
rect 198779 558179 198845 558180
rect 201542 557701 201602 559950
rect 202462 558653 202522 560290
rect 202766 559330 202826 560320
rect 202646 559270 202826 559330
rect 203750 560290 203840 560350
rect 202646 558925 202706 559270
rect 203750 558925 203810 560290
rect 203934 558925 203994 560320
rect 204854 560290 205008 560350
rect 205132 560290 205466 560350
rect 202643 558924 202709 558925
rect 202643 558860 202644 558924
rect 202708 558860 202709 558924
rect 202643 558859 202709 558860
rect 203747 558924 203813 558925
rect 203747 558860 203748 558924
rect 203812 558860 203813 558924
rect 203747 558859 203813 558860
rect 203931 558924 203997 558925
rect 203931 558860 203932 558924
rect 203996 558860 203997 558924
rect 203931 558859 203997 558860
rect 204854 558653 204914 560290
rect 205406 558925 205466 560290
rect 206142 558925 206202 560350
rect 206300 560290 206938 560350
rect 205403 558924 205469 558925
rect 205403 558860 205404 558924
rect 205468 558860 205469 558924
rect 205403 558859 205469 558860
rect 206139 558924 206205 558925
rect 206139 558860 206140 558924
rect 206204 558860 206205 558924
rect 206139 558859 206205 558860
rect 202459 558652 202525 558653
rect 202459 558588 202460 558652
rect 202524 558588 202525 558652
rect 202459 558587 202525 558588
rect 204851 558652 204917 558653
rect 204851 558588 204852 558652
rect 204916 558588 204917 558652
rect 204851 558587 204917 558588
rect 201539 557700 201605 557701
rect 201539 557636 201540 557700
rect 201604 557636 201605 557700
rect 201539 557635 201605 557636
rect 206878 557565 206938 560290
rect 207062 557701 207122 560430
rect 207468 560290 208042 560350
rect 207059 557700 207125 557701
rect 207059 557636 207060 557700
rect 207124 557636 207125 557700
rect 207059 557635 207125 557636
rect 207982 557565 208042 560290
rect 208350 560290 208512 560350
rect 208636 560290 209330 560350
rect 208350 558925 208410 560290
rect 208347 558924 208413 558925
rect 208347 558860 208348 558924
rect 208412 558860 208413 558924
rect 208347 558859 208413 558860
rect 209270 557565 209330 560290
rect 209638 558653 209698 560350
rect 209804 560290 210434 560350
rect 209635 558652 209701 558653
rect 209635 558588 209636 558652
rect 209700 558588 209701 558652
rect 209635 558587 209701 558588
rect 210374 557701 210434 560290
rect 210558 560290 210848 560350
rect 210558 558925 210618 560290
rect 210942 560010 211002 560320
rect 211846 560290 212016 560350
rect 212140 560290 212458 560350
rect 211107 560012 211173 560013
rect 211107 560010 211108 560012
rect 210942 559950 211108 560010
rect 211107 559948 211108 559950
rect 211172 559948 211173 560012
rect 211107 559947 211173 559948
rect 211846 558925 211906 560290
rect 210555 558924 210621 558925
rect 210555 558860 210556 558924
rect 210620 558860 210621 558924
rect 210555 558859 210621 558860
rect 211843 558924 211909 558925
rect 211843 558860 211844 558924
rect 211908 558860 211909 558924
rect 211843 558859 211909 558860
rect 210371 557700 210437 557701
rect 210371 557636 210372 557700
rect 210436 557636 210437 557700
rect 210371 557635 210437 557636
rect 212398 557565 212458 560290
rect 213134 558925 213194 560350
rect 213308 560290 213562 560350
rect 213131 558924 213197 558925
rect 213131 558860 213132 558924
rect 213196 558860 213197 558924
rect 213131 558859 213197 558860
rect 213502 557565 213562 560290
rect 214054 558925 214114 560430
rect 214476 560290 214850 560350
rect 214051 558924 214117 558925
rect 214051 558860 214052 558924
rect 214116 558860 214117 558924
rect 214051 558859 214117 558860
rect 214790 557565 214850 560290
rect 215342 560290 215520 560350
rect 215644 560290 216322 560350
rect 215342 558925 215402 560290
rect 215339 558924 215405 558925
rect 215339 558860 215340 558924
rect 215404 558860 215405 558924
rect 215339 558859 215405 558860
rect 216262 557565 216322 560290
rect 216630 558925 216690 560350
rect 216812 560290 217426 560350
rect 216627 558924 216693 558925
rect 216627 558860 216628 558924
rect 216692 558860 216693 558924
rect 216627 558859 216693 558860
rect 217366 557701 217426 560290
rect 217550 558789 217610 560430
rect 217950 559330 218010 560320
rect 217918 559270 218010 559330
rect 218838 560290 219024 560350
rect 217547 558788 217613 558789
rect 217547 558724 217548 558788
rect 217612 558724 217613 558788
rect 217547 558723 217613 558724
rect 217363 557700 217429 557701
rect 217363 557636 217364 557700
rect 217428 557636 217429 557700
rect 217363 557635 217429 557636
rect 217918 557565 217978 559270
rect 218838 558925 218898 560290
rect 219118 560010 219178 560320
rect 220126 560290 220192 560350
rect 220316 560290 220738 560350
rect 219118 559950 219266 560010
rect 218835 558924 218901 558925
rect 218835 558860 218836 558924
rect 218900 558860 218901 558924
rect 218835 558859 218901 558860
rect 219206 557565 219266 559950
rect 220126 558925 220186 560290
rect 220123 558924 220189 558925
rect 220123 558860 220124 558924
rect 220188 558860 220189 558924
rect 220123 558859 220189 558860
rect 220678 557565 220738 560290
rect 221046 558925 221106 560430
rect 221484 560290 222026 560350
rect 221043 558924 221109 558925
rect 221043 558860 221044 558924
rect 221108 558860 221109 558924
rect 221043 558859 221109 558860
rect 221966 557565 222026 560290
rect 222334 560290 222528 560350
rect 222652 560290 223314 560350
rect 222334 558925 222394 560290
rect 222331 558924 222397 558925
rect 222331 558860 222332 558924
rect 222396 558860 222397 558924
rect 222331 558859 222397 558860
rect 223254 557565 223314 560290
rect 223622 560290 223696 560350
rect 223820 560290 224418 560350
rect 223622 558789 223682 560290
rect 223619 558788 223685 558789
rect 223619 558724 223620 558788
rect 223684 558724 223685 558788
rect 223619 558723 223685 558724
rect 224358 557565 224418 560290
rect 224542 560290 224864 560350
rect 224988 560290 225706 560350
rect 224542 558925 224602 560290
rect 224539 558924 224605 558925
rect 224539 558860 224540 558924
rect 224604 558860 224605 558924
rect 224539 558859 224605 558860
rect 225646 558789 225706 560290
rect 225830 560290 226032 560350
rect 225830 558925 225890 560290
rect 226126 560010 226186 560320
rect 227118 560290 227200 560350
rect 227324 560290 227546 560350
rect 226126 559950 226258 560010
rect 226198 558925 226258 559950
rect 227118 558925 227178 560290
rect 227486 558925 227546 560290
rect 228038 558925 228098 560430
rect 228492 560290 228834 560350
rect 228774 558925 228834 560290
rect 229506 560010 229566 560320
rect 229660 560290 230306 560350
rect 229506 559950 229570 560010
rect 229510 558925 229570 559950
rect 230246 558925 230306 560290
rect 230614 560290 230704 560350
rect 225827 558924 225893 558925
rect 225827 558860 225828 558924
rect 225892 558860 225893 558924
rect 225827 558859 225893 558860
rect 226195 558924 226261 558925
rect 226195 558860 226196 558924
rect 226260 558860 226261 558924
rect 226195 558859 226261 558860
rect 227115 558924 227181 558925
rect 227115 558860 227116 558924
rect 227180 558860 227181 558924
rect 227115 558859 227181 558860
rect 227483 558924 227549 558925
rect 227483 558860 227484 558924
rect 227548 558860 227549 558924
rect 227483 558859 227549 558860
rect 228035 558924 228101 558925
rect 228035 558860 228036 558924
rect 228100 558860 228101 558924
rect 228035 558859 228101 558860
rect 228771 558924 228837 558925
rect 228771 558860 228772 558924
rect 228836 558860 228837 558924
rect 228771 558859 228837 558860
rect 229507 558924 229573 558925
rect 229507 558860 229508 558924
rect 229572 558860 229573 558924
rect 229507 558859 229573 558860
rect 230243 558924 230309 558925
rect 230243 558860 230244 558924
rect 230308 558860 230309 558924
rect 230243 558859 230309 558860
rect 225643 558788 225709 558789
rect 225643 558724 225644 558788
rect 225708 558724 225709 558788
rect 225643 558723 225709 558724
rect 230614 558381 230674 560290
rect 230798 558925 230858 560320
rect 231842 559330 231902 560320
rect 231996 560290 232698 560350
rect 231842 559270 231962 559330
rect 230795 558924 230861 558925
rect 230795 558860 230796 558924
rect 230860 558860 230861 558924
rect 230795 558859 230861 558860
rect 231902 558789 231962 559270
rect 232638 558789 232698 560290
rect 232822 560290 233040 560350
rect 231899 558788 231965 558789
rect 231899 558724 231900 558788
rect 231964 558724 231965 558788
rect 231899 558723 231965 558724
rect 232635 558788 232701 558789
rect 232635 558724 232636 558788
rect 232700 558724 232701 558788
rect 232635 558723 232701 558724
rect 232822 558517 232882 560290
rect 233134 559330 233194 560320
rect 233006 559270 233194 559330
rect 233558 560290 234208 560350
rect 234332 560290 234538 560350
rect 233006 558925 233066 559270
rect 233558 558925 233618 560290
rect 234478 558925 234538 560290
rect 234662 560290 235376 560350
rect 235500 560290 235826 560350
rect 233003 558924 233069 558925
rect 233003 558860 233004 558924
rect 233068 558860 233069 558924
rect 233003 558859 233069 558860
rect 233555 558924 233621 558925
rect 233555 558860 233556 558924
rect 233620 558860 233621 558924
rect 233555 558859 233621 558860
rect 234475 558924 234541 558925
rect 234475 558860 234476 558924
rect 234540 558860 234541 558924
rect 234475 558859 234541 558860
rect 234662 558789 234722 560290
rect 235766 558925 235826 560290
rect 236134 560290 236544 560350
rect 236668 560290 237298 560350
rect 235763 558924 235829 558925
rect 235763 558860 235764 558924
rect 235828 558860 235829 558924
rect 235763 558859 235829 558860
rect 236134 558789 236194 560290
rect 237238 558925 237298 560290
rect 237422 560290 237712 560350
rect 237836 560290 238402 560350
rect 237235 558924 237301 558925
rect 237235 558860 237236 558924
rect 237300 558860 237301 558924
rect 237235 558859 237301 558860
rect 237422 558789 237482 560290
rect 234659 558788 234725 558789
rect 234659 558724 234660 558788
rect 234724 558724 234725 558788
rect 234659 558723 234725 558724
rect 236131 558788 236197 558789
rect 236131 558724 236132 558788
rect 236196 558724 236197 558788
rect 236131 558723 236197 558724
rect 237419 558788 237485 558789
rect 237419 558724 237420 558788
rect 237484 558724 237485 558788
rect 237419 558723 237485 558724
rect 232819 558516 232885 558517
rect 232819 558452 232820 558516
rect 232884 558452 232885 558516
rect 232819 558451 232885 558452
rect 230611 558380 230677 558381
rect 230611 558316 230612 558380
rect 230676 558316 230677 558380
rect 230611 558315 230677 558316
rect 238342 558109 238402 560290
rect 238710 560290 238880 560350
rect 239004 560290 239690 560350
rect 238710 558381 238770 560290
rect 239630 558925 239690 560290
rect 270804 560218 270986 560454
rect 271222 560218 271404 560454
rect 270804 560134 271404 560218
rect 270804 559898 270986 560134
rect 271222 559898 271404 560134
rect 239627 558924 239693 558925
rect 239627 558860 239628 558924
rect 239692 558860 239693 558924
rect 239627 558859 239693 558860
rect 238707 558380 238773 558381
rect 238707 558316 238708 558380
rect 238772 558316 238773 558380
rect 238707 558315 238773 558316
rect 238339 558108 238405 558109
rect 238339 558044 238340 558108
rect 238404 558044 238405 558108
rect 238339 558043 238405 558044
rect 206875 557564 206941 557565
rect 206875 557500 206876 557564
rect 206940 557500 206941 557564
rect 206875 557499 206941 557500
rect 207979 557564 208045 557565
rect 207979 557500 207980 557564
rect 208044 557500 208045 557564
rect 207979 557499 208045 557500
rect 209267 557564 209333 557565
rect 209267 557500 209268 557564
rect 209332 557500 209333 557564
rect 209267 557499 209333 557500
rect 212395 557564 212461 557565
rect 212395 557500 212396 557564
rect 212460 557500 212461 557564
rect 212395 557499 212461 557500
rect 213499 557564 213565 557565
rect 213499 557500 213500 557564
rect 213564 557500 213565 557564
rect 213499 557499 213565 557500
rect 214787 557564 214853 557565
rect 214787 557500 214788 557564
rect 214852 557500 214853 557564
rect 214787 557499 214853 557500
rect 216259 557564 216325 557565
rect 216259 557500 216260 557564
rect 216324 557500 216325 557564
rect 216259 557499 216325 557500
rect 217915 557564 217981 557565
rect 217915 557500 217916 557564
rect 217980 557500 217981 557564
rect 217915 557499 217981 557500
rect 219203 557564 219269 557565
rect 219203 557500 219204 557564
rect 219268 557500 219269 557564
rect 219203 557499 219269 557500
rect 220675 557564 220741 557565
rect 220675 557500 220676 557564
rect 220740 557500 220741 557564
rect 220675 557499 220741 557500
rect 221963 557564 222029 557565
rect 221963 557500 221964 557564
rect 222028 557500 222029 557564
rect 221963 557499 222029 557500
rect 223251 557564 223317 557565
rect 223251 557500 223252 557564
rect 223316 557500 223317 557564
rect 223251 557499 223317 557500
rect 224355 557564 224421 557565
rect 224355 557500 224356 557564
rect 224420 557500 224421 557564
rect 224355 557499 224421 557500
rect 184404 545818 184586 546054
rect 184822 545818 185004 546054
rect 184404 545734 185004 545818
rect 184404 545498 184586 545734
rect 184822 545498 185004 545734
rect 184404 543000 185004 545498
rect 188004 549654 188604 557000
rect 188004 549418 188186 549654
rect 188422 549418 188604 549654
rect 188004 549334 188604 549418
rect 188004 549098 188186 549334
rect 188422 549098 188604 549334
rect 188004 543000 188604 549098
rect 191604 553254 192204 557000
rect 191604 553018 191786 553254
rect 192022 553018 192204 553254
rect 191604 552934 192204 553018
rect 191604 552698 191786 552934
rect 192022 552698 192204 552934
rect 191604 543000 192204 552698
rect 198804 543000 199404 557000
rect 202404 543000 203004 557000
rect 206004 543000 206604 557000
rect 209604 543000 210204 557000
rect 216804 543000 217404 557000
rect 220404 546054 221004 557000
rect 220404 545818 220586 546054
rect 220822 545818 221004 546054
rect 220404 545734 221004 545818
rect 220404 545498 220586 545734
rect 220822 545498 221004 545734
rect 220404 543000 221004 545498
rect 224004 549654 224604 557000
rect 224004 549418 224186 549654
rect 224422 549418 224604 549654
rect 224004 549334 224604 549418
rect 224004 549098 224186 549334
rect 224422 549098 224604 549334
rect 224004 543000 224604 549098
rect 227604 553254 228204 557000
rect 227604 553018 227786 553254
rect 228022 553018 228204 553254
rect 227604 552934 228204 553018
rect 227604 552698 227786 552934
rect 228022 552698 228204 552934
rect 227604 543000 228204 552698
rect 234804 543000 235404 557000
rect 238404 543000 239004 557000
rect 242004 543000 242604 557000
rect 245604 543000 246204 557000
rect 252804 543000 253404 557000
rect 256404 546054 257004 557000
rect 256404 545818 256586 546054
rect 256822 545818 257004 546054
rect 256404 545734 257004 545818
rect 256404 545498 256586 545734
rect 256822 545498 257004 545734
rect 256404 543000 257004 545498
rect 260004 549654 260604 557000
rect 260004 549418 260186 549654
rect 260422 549418 260604 549654
rect 260004 549334 260604 549418
rect 260004 549098 260186 549334
rect 260422 549098 260604 549334
rect 260004 543000 260604 549098
rect 263604 553254 264204 557000
rect 263604 553018 263786 553254
rect 264022 553018 264204 553254
rect 263604 552934 264204 553018
rect 263604 552698 263786 552934
rect 264022 552698 264204 552934
rect 263604 543000 264204 552698
rect 270804 543000 271404 559898
rect 274404 672054 275004 707102
rect 274404 671818 274586 672054
rect 274822 671818 275004 672054
rect 274404 671734 275004 671818
rect 274404 671498 274586 671734
rect 274822 671498 275004 671734
rect 274404 636054 275004 671498
rect 274404 635818 274586 636054
rect 274822 635818 275004 636054
rect 274404 635734 275004 635818
rect 274404 635498 274586 635734
rect 274822 635498 275004 635734
rect 274404 600054 275004 635498
rect 274404 599818 274586 600054
rect 274822 599818 275004 600054
rect 274404 599734 275004 599818
rect 274404 599498 274586 599734
rect 274822 599498 275004 599734
rect 274404 564054 275004 599498
rect 274404 563818 274586 564054
rect 274822 563818 275004 564054
rect 274404 563734 275004 563818
rect 274404 563498 274586 563734
rect 274822 563498 275004 563734
rect 274404 543000 275004 563498
rect 278004 675654 278604 708982
rect 278004 675418 278186 675654
rect 278422 675418 278604 675654
rect 278004 675334 278604 675418
rect 278004 675098 278186 675334
rect 278422 675098 278604 675334
rect 278004 639654 278604 675098
rect 278004 639418 278186 639654
rect 278422 639418 278604 639654
rect 278004 639334 278604 639418
rect 278004 639098 278186 639334
rect 278422 639098 278604 639334
rect 278004 603654 278604 639098
rect 278004 603418 278186 603654
rect 278422 603418 278604 603654
rect 278004 603334 278604 603418
rect 278004 603098 278186 603334
rect 278422 603098 278604 603334
rect 278004 567654 278604 603098
rect 278004 567418 278186 567654
rect 278422 567418 278604 567654
rect 278004 567334 278604 567418
rect 278004 567098 278186 567334
rect 278422 567098 278604 567334
rect 278004 543000 278604 567098
rect 281604 679254 282204 710862
rect 299604 710478 300204 711440
rect 299604 710242 299786 710478
rect 300022 710242 300204 710478
rect 299604 710158 300204 710242
rect 299604 709922 299786 710158
rect 300022 709922 300204 710158
rect 296004 708598 296604 709560
rect 296004 708362 296186 708598
rect 296422 708362 296604 708598
rect 296004 708278 296604 708362
rect 296004 708042 296186 708278
rect 296422 708042 296604 708278
rect 292404 706718 293004 707680
rect 292404 706482 292586 706718
rect 292822 706482 293004 706718
rect 292404 706398 293004 706482
rect 292404 706162 292586 706398
rect 292822 706162 293004 706398
rect 281604 679018 281786 679254
rect 282022 679018 282204 679254
rect 281604 678934 282204 679018
rect 281604 678698 281786 678934
rect 282022 678698 282204 678934
rect 281604 643254 282204 678698
rect 281604 643018 281786 643254
rect 282022 643018 282204 643254
rect 281604 642934 282204 643018
rect 281604 642698 281786 642934
rect 282022 642698 282204 642934
rect 281604 607254 282204 642698
rect 281604 607018 281786 607254
rect 282022 607018 282204 607254
rect 281604 606934 282204 607018
rect 281604 606698 281786 606934
rect 282022 606698 282204 606934
rect 281604 571254 282204 606698
rect 288804 704838 289404 705800
rect 288804 704602 288986 704838
rect 289222 704602 289404 704838
rect 288804 704518 289404 704602
rect 288804 704282 288986 704518
rect 289222 704282 289404 704518
rect 288804 686454 289404 704282
rect 288804 686218 288986 686454
rect 289222 686218 289404 686454
rect 288804 686134 289404 686218
rect 288804 685898 288986 686134
rect 289222 685898 289404 686134
rect 288804 650454 289404 685898
rect 288804 650218 288986 650454
rect 289222 650218 289404 650454
rect 288804 650134 289404 650218
rect 288804 649898 288986 650134
rect 289222 649898 289404 650134
rect 288804 614454 289404 649898
rect 288804 614218 288986 614454
rect 289222 614218 289404 614454
rect 288804 614134 289404 614218
rect 288804 613898 288986 614134
rect 289222 613898 289404 614134
rect 281604 571018 281786 571254
rect 282022 571018 282204 571254
rect 281604 570934 282204 571018
rect 281604 570698 281786 570934
rect 282022 570698 282204 570934
rect 281604 543000 282204 570698
rect 288804 578454 289404 613898
rect 288804 578218 288986 578454
rect 289222 578218 289404 578454
rect 288804 578134 289404 578218
rect 288804 577898 288986 578134
rect 289222 577898 289404 578134
rect 282315 558380 282381 558381
rect 282315 558316 282316 558380
rect 282380 558316 282381 558380
rect 282315 558315 282381 558316
rect 79568 535254 79888 535276
rect 79568 535018 79610 535254
rect 79846 535018 79888 535254
rect 79568 534934 79888 535018
rect 79568 534698 79610 534934
rect 79846 534698 79888 534934
rect 79568 534676 79888 534698
rect 79568 531654 79888 531676
rect 79568 531418 79610 531654
rect 79846 531418 79888 531654
rect 79568 531334 79888 531418
rect 79568 531098 79610 531334
rect 79846 531098 79888 531334
rect 79568 531076 79888 531098
rect 79568 528054 79888 528076
rect 79568 527818 79610 528054
rect 79846 527818 79888 528054
rect 79568 527734 79888 527818
rect 79568 527498 79610 527734
rect 79846 527498 79888 527734
rect 79568 527476 79888 527498
rect 54804 524218 54986 524454
rect 55222 524218 55404 524454
rect 54804 524134 55404 524218
rect 54804 523898 54986 524134
rect 55222 523898 55404 524134
rect 54804 488454 55404 523898
rect 79568 524454 79888 524476
rect 79568 524218 79610 524454
rect 79846 524218 79888 524454
rect 79568 524134 79888 524218
rect 79568 523898 79610 524134
rect 79846 523898 79888 524134
rect 79568 523876 79888 523898
rect 64208 517254 64528 517276
rect 64208 517018 64250 517254
rect 64486 517018 64528 517254
rect 64208 516934 64528 517018
rect 64208 516698 64250 516934
rect 64486 516698 64528 516934
rect 64208 516676 64528 516698
rect 64208 513654 64528 513676
rect 64208 513418 64250 513654
rect 64486 513418 64528 513654
rect 64208 513334 64528 513418
rect 64208 513098 64250 513334
rect 64486 513098 64528 513334
rect 64208 513076 64528 513098
rect 64208 510054 64528 510076
rect 64208 509818 64250 510054
rect 64486 509818 64528 510054
rect 64208 509734 64528 509818
rect 64208 509498 64250 509734
rect 64486 509498 64528 509734
rect 64208 509476 64528 509498
rect 64208 506454 64528 506476
rect 64208 506218 64250 506454
rect 64486 506218 64528 506454
rect 64208 506134 64528 506218
rect 64208 505898 64250 506134
rect 64486 505898 64528 506134
rect 64208 505876 64528 505898
rect 79568 499254 79888 499276
rect 79568 499018 79610 499254
rect 79846 499018 79888 499254
rect 79568 498934 79888 499018
rect 79568 498698 79610 498934
rect 79846 498698 79888 498934
rect 79568 498676 79888 498698
rect 79568 495654 79888 495676
rect 79568 495418 79610 495654
rect 79846 495418 79888 495654
rect 79568 495334 79888 495418
rect 79568 495098 79610 495334
rect 79846 495098 79888 495334
rect 79568 495076 79888 495098
rect 79568 492054 79888 492076
rect 79568 491818 79610 492054
rect 79846 491818 79888 492054
rect 79568 491734 79888 491818
rect 79568 491498 79610 491734
rect 79846 491498 79888 491734
rect 79568 491476 79888 491498
rect 54804 488218 54986 488454
rect 55222 488218 55404 488454
rect 54804 488134 55404 488218
rect 54804 487898 54986 488134
rect 55222 487898 55404 488134
rect 54804 452454 55404 487898
rect 79568 488454 79888 488476
rect 79568 488218 79610 488454
rect 79846 488218 79888 488454
rect 79568 488134 79888 488218
rect 79568 487898 79610 488134
rect 79846 487898 79888 488134
rect 79568 487876 79888 487898
rect 64208 481254 64528 481276
rect 64208 481018 64250 481254
rect 64486 481018 64528 481254
rect 64208 480934 64528 481018
rect 64208 480698 64250 480934
rect 64486 480698 64528 480934
rect 64208 480676 64528 480698
rect 64208 477654 64528 477676
rect 64208 477418 64250 477654
rect 64486 477418 64528 477654
rect 64208 477334 64528 477418
rect 64208 477098 64250 477334
rect 64486 477098 64528 477334
rect 64208 477076 64528 477098
rect 64208 474054 64528 474076
rect 64208 473818 64250 474054
rect 64486 473818 64528 474054
rect 64208 473734 64528 473818
rect 64208 473498 64250 473734
rect 64486 473498 64528 473734
rect 64208 473476 64528 473498
rect 64208 470454 64528 470476
rect 64208 470218 64250 470454
rect 64486 470218 64528 470454
rect 64208 470134 64528 470218
rect 64208 469898 64250 470134
rect 64486 469898 64528 470134
rect 64208 469876 64528 469898
rect 79568 463254 79888 463276
rect 79568 463018 79610 463254
rect 79846 463018 79888 463254
rect 79568 462934 79888 463018
rect 79568 462698 79610 462934
rect 79846 462698 79888 462934
rect 79568 462676 79888 462698
rect 79568 459654 79888 459676
rect 79568 459418 79610 459654
rect 79846 459418 79888 459654
rect 79568 459334 79888 459418
rect 79568 459098 79610 459334
rect 79846 459098 79888 459334
rect 79568 459076 79888 459098
rect 79568 456054 79888 456076
rect 79568 455818 79610 456054
rect 79846 455818 79888 456054
rect 79568 455734 79888 455818
rect 79568 455498 79610 455734
rect 79846 455498 79888 455734
rect 79568 455476 79888 455498
rect 54804 452218 54986 452454
rect 55222 452218 55404 452454
rect 54804 452134 55404 452218
rect 54804 451898 54986 452134
rect 55222 451898 55404 452134
rect 54804 416454 55404 451898
rect 79568 452454 79888 452476
rect 79568 452218 79610 452454
rect 79846 452218 79888 452454
rect 79568 452134 79888 452218
rect 79568 451898 79610 452134
rect 79846 451898 79888 452134
rect 79568 451876 79888 451898
rect 64208 445254 64528 445276
rect 64208 445018 64250 445254
rect 64486 445018 64528 445254
rect 64208 444934 64528 445018
rect 64208 444698 64250 444934
rect 64486 444698 64528 444934
rect 64208 444676 64528 444698
rect 64208 441654 64528 441676
rect 64208 441418 64250 441654
rect 64486 441418 64528 441654
rect 64208 441334 64528 441418
rect 64208 441098 64250 441334
rect 64486 441098 64528 441334
rect 64208 441076 64528 441098
rect 64208 438054 64528 438076
rect 64208 437818 64250 438054
rect 64486 437818 64528 438054
rect 64208 437734 64528 437818
rect 64208 437498 64250 437734
rect 64486 437498 64528 437734
rect 64208 437476 64528 437498
rect 64208 434454 64528 434476
rect 64208 434218 64250 434454
rect 64486 434218 64528 434454
rect 64208 434134 64528 434218
rect 64208 433898 64250 434134
rect 64486 433898 64528 434134
rect 64208 433876 64528 433898
rect 79568 427254 79888 427276
rect 79568 427018 79610 427254
rect 79846 427018 79888 427254
rect 79568 426934 79888 427018
rect 79568 426698 79610 426934
rect 79846 426698 79888 426934
rect 79568 426676 79888 426698
rect 79568 423654 79888 423676
rect 79568 423418 79610 423654
rect 79846 423418 79888 423654
rect 79568 423334 79888 423418
rect 79568 423098 79610 423334
rect 79846 423098 79888 423334
rect 79568 423076 79888 423098
rect 79568 420054 79888 420076
rect 79568 419818 79610 420054
rect 79846 419818 79888 420054
rect 79568 419734 79888 419818
rect 79568 419498 79610 419734
rect 79846 419498 79888 419734
rect 79568 419476 79888 419498
rect 54804 416218 54986 416454
rect 55222 416218 55404 416454
rect 54804 416134 55404 416218
rect 54804 415898 54986 416134
rect 55222 415898 55404 416134
rect 54804 380454 55404 415898
rect 79568 416454 79888 416476
rect 79568 416218 79610 416454
rect 79846 416218 79888 416454
rect 79568 416134 79888 416218
rect 79568 415898 79610 416134
rect 79846 415898 79888 416134
rect 79568 415876 79888 415898
rect 64208 409254 64528 409276
rect 64208 409018 64250 409254
rect 64486 409018 64528 409254
rect 64208 408934 64528 409018
rect 64208 408698 64250 408934
rect 64486 408698 64528 408934
rect 64208 408676 64528 408698
rect 64208 405654 64528 405676
rect 64208 405418 64250 405654
rect 64486 405418 64528 405654
rect 64208 405334 64528 405418
rect 64208 405098 64250 405334
rect 64486 405098 64528 405334
rect 64208 405076 64528 405098
rect 64208 402054 64528 402076
rect 64208 401818 64250 402054
rect 64486 401818 64528 402054
rect 64208 401734 64528 401818
rect 64208 401498 64250 401734
rect 64486 401498 64528 401734
rect 64208 401476 64528 401498
rect 64208 398454 64528 398476
rect 64208 398218 64250 398454
rect 64486 398218 64528 398454
rect 64208 398134 64528 398218
rect 64208 397898 64250 398134
rect 64486 397898 64528 398134
rect 64208 397876 64528 397898
rect 79568 391254 79888 391276
rect 79568 391018 79610 391254
rect 79846 391018 79888 391254
rect 79568 390934 79888 391018
rect 79568 390698 79610 390934
rect 79846 390698 79888 390934
rect 79568 390676 79888 390698
rect 79568 387654 79888 387676
rect 79568 387418 79610 387654
rect 79846 387418 79888 387654
rect 79568 387334 79888 387418
rect 79568 387098 79610 387334
rect 79846 387098 79888 387334
rect 79568 387076 79888 387098
rect 79568 384054 79888 384076
rect 79568 383818 79610 384054
rect 79846 383818 79888 384054
rect 79568 383734 79888 383818
rect 79568 383498 79610 383734
rect 79846 383498 79888 383734
rect 79568 383476 79888 383498
rect 54804 380218 54986 380454
rect 55222 380218 55404 380454
rect 54804 380134 55404 380218
rect 54804 379898 54986 380134
rect 55222 379898 55404 380134
rect 54804 344454 55404 379898
rect 79568 380454 79888 380476
rect 79568 380218 79610 380454
rect 79846 380218 79888 380454
rect 79568 380134 79888 380218
rect 79568 379898 79610 380134
rect 79846 379898 79888 380134
rect 79568 379876 79888 379898
rect 64208 373254 64528 373276
rect 64208 373018 64250 373254
rect 64486 373018 64528 373254
rect 64208 372934 64528 373018
rect 64208 372698 64250 372934
rect 64486 372698 64528 372934
rect 64208 372676 64528 372698
rect 64208 369654 64528 369676
rect 64208 369418 64250 369654
rect 64486 369418 64528 369654
rect 64208 369334 64528 369418
rect 64208 369098 64250 369334
rect 64486 369098 64528 369334
rect 64208 369076 64528 369098
rect 64208 366054 64528 366076
rect 64208 365818 64250 366054
rect 64486 365818 64528 366054
rect 64208 365734 64528 365818
rect 64208 365498 64250 365734
rect 64486 365498 64528 365734
rect 64208 365476 64528 365498
rect 64208 362454 64528 362476
rect 64208 362218 64250 362454
rect 64486 362218 64528 362454
rect 64208 362134 64528 362218
rect 64208 361898 64250 362134
rect 64486 361898 64528 362134
rect 64208 361876 64528 361898
rect 79568 355254 79888 355276
rect 79568 355018 79610 355254
rect 79846 355018 79888 355254
rect 79568 354934 79888 355018
rect 79568 354698 79610 354934
rect 79846 354698 79888 354934
rect 79568 354676 79888 354698
rect 79568 351654 79888 351676
rect 79568 351418 79610 351654
rect 79846 351418 79888 351654
rect 79568 351334 79888 351418
rect 79568 351098 79610 351334
rect 79846 351098 79888 351334
rect 79568 351076 79888 351098
rect 79568 348054 79888 348076
rect 79568 347818 79610 348054
rect 79846 347818 79888 348054
rect 79568 347734 79888 347818
rect 79568 347498 79610 347734
rect 79846 347498 79888 347734
rect 79568 347476 79888 347498
rect 54804 344218 54986 344454
rect 55222 344218 55404 344454
rect 54804 344134 55404 344218
rect 54804 343898 54986 344134
rect 55222 343898 55404 344134
rect 54804 308454 55404 343898
rect 79568 344454 79888 344476
rect 79568 344218 79610 344454
rect 79846 344218 79888 344454
rect 79568 344134 79888 344218
rect 79568 343898 79610 344134
rect 79846 343898 79888 344134
rect 79568 343876 79888 343898
rect 64208 337254 64528 337276
rect 64208 337018 64250 337254
rect 64486 337018 64528 337254
rect 64208 336934 64528 337018
rect 64208 336698 64250 336934
rect 64486 336698 64528 336934
rect 64208 336676 64528 336698
rect 64208 333654 64528 333676
rect 64208 333418 64250 333654
rect 64486 333418 64528 333654
rect 64208 333334 64528 333418
rect 64208 333098 64250 333334
rect 64486 333098 64528 333334
rect 64208 333076 64528 333098
rect 64208 330054 64528 330076
rect 64208 329818 64250 330054
rect 64486 329818 64528 330054
rect 64208 329734 64528 329818
rect 64208 329498 64250 329734
rect 64486 329498 64528 329734
rect 64208 329476 64528 329498
rect 64208 326454 64528 326476
rect 64208 326218 64250 326454
rect 64486 326218 64528 326454
rect 64208 326134 64528 326218
rect 64208 325898 64250 326134
rect 64486 325898 64528 326134
rect 64208 325876 64528 325898
rect 282318 323509 282378 558315
rect 283419 558244 283485 558245
rect 283419 558180 283420 558244
rect 283484 558180 283485 558244
rect 283419 558179 283485 558180
rect 283422 324461 283482 558179
rect 288804 542454 289404 577898
rect 288804 542218 288986 542454
rect 289222 542218 289404 542454
rect 288804 542134 289404 542218
rect 288804 541898 288986 542134
rect 289222 541898 289404 542134
rect 288804 506454 289404 541898
rect 288804 506218 288986 506454
rect 289222 506218 289404 506454
rect 288804 506134 289404 506218
rect 288804 505898 288986 506134
rect 289222 505898 289404 506134
rect 288804 470454 289404 505898
rect 288804 470218 288986 470454
rect 289222 470218 289404 470454
rect 288804 470134 289404 470218
rect 288804 469898 288986 470134
rect 289222 469898 289404 470134
rect 288804 434454 289404 469898
rect 288804 434218 288986 434454
rect 289222 434218 289404 434454
rect 288804 434134 289404 434218
rect 288804 433898 288986 434134
rect 289222 433898 289404 434134
rect 288804 398454 289404 433898
rect 288804 398218 288986 398454
rect 289222 398218 289404 398454
rect 288804 398134 289404 398218
rect 288804 397898 288986 398134
rect 289222 397898 289404 398134
rect 288804 362454 289404 397898
rect 288804 362218 288986 362454
rect 289222 362218 289404 362454
rect 288804 362134 289404 362218
rect 288804 361898 288986 362134
rect 289222 361898 289404 362134
rect 288804 326454 289404 361898
rect 288804 326218 288986 326454
rect 289222 326218 289404 326454
rect 288804 326134 289404 326218
rect 288804 325898 288986 326134
rect 289222 325898 289404 326134
rect 283419 324460 283485 324461
rect 283419 324396 283420 324460
rect 283484 324396 283485 324460
rect 283419 324395 283485 324396
rect 282315 323508 282381 323509
rect 282315 323444 282316 323508
rect 282380 323444 282381 323508
rect 282315 323443 282381 323444
rect 54804 308218 54986 308454
rect 55222 308218 55404 308454
rect 54804 308134 55404 308218
rect 54804 307898 54986 308134
rect 55222 307898 55404 308134
rect 54804 272454 55404 307898
rect 54804 272218 54986 272454
rect 55222 272218 55404 272454
rect 54804 272134 55404 272218
rect 54804 271898 54986 272134
rect 55222 271898 55404 272134
rect 54804 236454 55404 271898
rect 54804 236218 54986 236454
rect 55222 236218 55404 236454
rect 54804 236134 55404 236218
rect 54804 235898 54986 236134
rect 55222 235898 55404 236134
rect 54804 200454 55404 235898
rect 54804 200218 54986 200454
rect 55222 200218 55404 200454
rect 54804 200134 55404 200218
rect 54804 199898 54986 200134
rect 55222 199898 55404 200134
rect 54804 164454 55404 199898
rect 54804 164218 54986 164454
rect 55222 164218 55404 164454
rect 54804 164134 55404 164218
rect 54804 163898 54986 164134
rect 55222 163898 55404 164134
rect 54804 128454 55404 163898
rect 54804 128218 54986 128454
rect 55222 128218 55404 128454
rect 54804 128134 55404 128218
rect 54804 127898 54986 128134
rect 55222 127898 55404 128134
rect 54804 92454 55404 127898
rect 54804 92218 54986 92454
rect 55222 92218 55404 92454
rect 54804 92134 55404 92218
rect 54804 91898 54986 92134
rect 55222 91898 55404 92134
rect 54804 56454 55404 91898
rect 54804 56218 54986 56454
rect 55222 56218 55404 56454
rect 54804 56134 55404 56218
rect 54804 55898 54986 56134
rect 55222 55898 55404 56134
rect 54804 20454 55404 55898
rect 54804 20218 54986 20454
rect 55222 20218 55404 20454
rect 54804 20134 55404 20218
rect 54804 19898 54986 20134
rect 55222 19898 55404 20134
rect 54804 -1286 55404 19898
rect 54804 -1522 54986 -1286
rect 55222 -1522 55404 -1286
rect 54804 -1606 55404 -1522
rect 54804 -1842 54986 -1606
rect 55222 -1842 55404 -1606
rect 54804 -1864 55404 -1842
rect 58404 312054 59004 317000
rect 58404 311818 58586 312054
rect 58822 311818 59004 312054
rect 58404 311734 59004 311818
rect 58404 311498 58586 311734
rect 58822 311498 59004 311734
rect 58404 276054 59004 311498
rect 58404 275818 58586 276054
rect 58822 275818 59004 276054
rect 58404 275734 59004 275818
rect 58404 275498 58586 275734
rect 58822 275498 59004 275734
rect 58404 240054 59004 275498
rect 58404 239818 58586 240054
rect 58822 239818 59004 240054
rect 58404 239734 59004 239818
rect 58404 239498 58586 239734
rect 58822 239498 59004 239734
rect 58404 204054 59004 239498
rect 58404 203818 58586 204054
rect 58822 203818 59004 204054
rect 58404 203734 59004 203818
rect 58404 203498 58586 203734
rect 58822 203498 59004 203734
rect 58404 168054 59004 203498
rect 58404 167818 58586 168054
rect 58822 167818 59004 168054
rect 58404 167734 59004 167818
rect 58404 167498 58586 167734
rect 58822 167498 59004 167734
rect 58404 132054 59004 167498
rect 58404 131818 58586 132054
rect 58822 131818 59004 132054
rect 58404 131734 59004 131818
rect 58404 131498 58586 131734
rect 58822 131498 59004 131734
rect 58404 96054 59004 131498
rect 58404 95818 58586 96054
rect 58822 95818 59004 96054
rect 58404 95734 59004 95818
rect 58404 95498 58586 95734
rect 58822 95498 59004 95734
rect 58404 60054 59004 95498
rect 58404 59818 58586 60054
rect 58822 59818 59004 60054
rect 58404 59734 59004 59818
rect 58404 59498 58586 59734
rect 58822 59498 59004 59734
rect 58404 24054 59004 59498
rect 58404 23818 58586 24054
rect 58822 23818 59004 24054
rect 58404 23734 59004 23818
rect 58404 23498 58586 23734
rect 58822 23498 59004 23734
rect 58404 -3166 59004 23498
rect 58404 -3402 58586 -3166
rect 58822 -3402 59004 -3166
rect 58404 -3486 59004 -3402
rect 58404 -3722 58586 -3486
rect 58822 -3722 59004 -3486
rect 58404 -3744 59004 -3722
rect 62004 315654 62604 317000
rect 62004 315418 62186 315654
rect 62422 315418 62604 315654
rect 62004 315334 62604 315418
rect 62004 315098 62186 315334
rect 62422 315098 62604 315334
rect 62004 279654 62604 315098
rect 62004 279418 62186 279654
rect 62422 279418 62604 279654
rect 62004 279334 62604 279418
rect 62004 279098 62186 279334
rect 62422 279098 62604 279334
rect 62004 243654 62604 279098
rect 62004 243418 62186 243654
rect 62422 243418 62604 243654
rect 62004 243334 62604 243418
rect 62004 243098 62186 243334
rect 62422 243098 62604 243334
rect 62004 207654 62604 243098
rect 62004 207418 62186 207654
rect 62422 207418 62604 207654
rect 62004 207334 62604 207418
rect 62004 207098 62186 207334
rect 62422 207098 62604 207334
rect 62004 171654 62604 207098
rect 62004 171418 62186 171654
rect 62422 171418 62604 171654
rect 62004 171334 62604 171418
rect 62004 171098 62186 171334
rect 62422 171098 62604 171334
rect 62004 135654 62604 171098
rect 62004 135418 62186 135654
rect 62422 135418 62604 135654
rect 62004 135334 62604 135418
rect 62004 135098 62186 135334
rect 62422 135098 62604 135334
rect 62004 99654 62604 135098
rect 62004 99418 62186 99654
rect 62422 99418 62604 99654
rect 62004 99334 62604 99418
rect 62004 99098 62186 99334
rect 62422 99098 62604 99334
rect 62004 63654 62604 99098
rect 62004 63418 62186 63654
rect 62422 63418 62604 63654
rect 62004 63334 62604 63418
rect 62004 63098 62186 63334
rect 62422 63098 62604 63334
rect 62004 27654 62604 63098
rect 62004 27418 62186 27654
rect 62422 27418 62604 27654
rect 62004 27334 62604 27418
rect 62004 27098 62186 27334
rect 62422 27098 62604 27334
rect 62004 -5046 62604 27098
rect 62004 -5282 62186 -5046
rect 62422 -5282 62604 -5046
rect 62004 -5366 62604 -5282
rect 62004 -5602 62186 -5366
rect 62422 -5602 62604 -5366
rect 62004 -5624 62604 -5602
rect 65604 283254 66204 317000
rect 65604 283018 65786 283254
rect 66022 283018 66204 283254
rect 65604 282934 66204 283018
rect 65604 282698 65786 282934
rect 66022 282698 66204 282934
rect 65604 247254 66204 282698
rect 65604 247018 65786 247254
rect 66022 247018 66204 247254
rect 65604 246934 66204 247018
rect 65604 246698 65786 246934
rect 66022 246698 66204 246934
rect 65604 211254 66204 246698
rect 65604 211018 65786 211254
rect 66022 211018 66204 211254
rect 65604 210934 66204 211018
rect 65604 210698 65786 210934
rect 66022 210698 66204 210934
rect 65604 175254 66204 210698
rect 65604 175018 65786 175254
rect 66022 175018 66204 175254
rect 65604 174934 66204 175018
rect 65604 174698 65786 174934
rect 66022 174698 66204 174934
rect 65604 139254 66204 174698
rect 65604 139018 65786 139254
rect 66022 139018 66204 139254
rect 65604 138934 66204 139018
rect 65604 138698 65786 138934
rect 66022 138698 66204 138934
rect 65604 103254 66204 138698
rect 65604 103018 65786 103254
rect 66022 103018 66204 103254
rect 65604 102934 66204 103018
rect 65604 102698 65786 102934
rect 66022 102698 66204 102934
rect 65604 67254 66204 102698
rect 65604 67018 65786 67254
rect 66022 67018 66204 67254
rect 65604 66934 66204 67018
rect 65604 66698 65786 66934
rect 66022 66698 66204 66934
rect 65604 31254 66204 66698
rect 65604 31018 65786 31254
rect 66022 31018 66204 31254
rect 65604 30934 66204 31018
rect 65604 30698 65786 30934
rect 66022 30698 66204 30934
rect 47604 -6222 47786 -5986
rect 48022 -6222 48204 -5986
rect 47604 -6306 48204 -6222
rect 47604 -6542 47786 -6306
rect 48022 -6542 48204 -6306
rect 47604 -7504 48204 -6542
rect 65604 -6926 66204 30698
rect 72804 290454 73404 317000
rect 72804 290218 72986 290454
rect 73222 290218 73404 290454
rect 72804 290134 73404 290218
rect 72804 289898 72986 290134
rect 73222 289898 73404 290134
rect 72804 254454 73404 289898
rect 72804 254218 72986 254454
rect 73222 254218 73404 254454
rect 72804 254134 73404 254218
rect 72804 253898 72986 254134
rect 73222 253898 73404 254134
rect 72804 218454 73404 253898
rect 72804 218218 72986 218454
rect 73222 218218 73404 218454
rect 72804 218134 73404 218218
rect 72804 217898 72986 218134
rect 73222 217898 73404 218134
rect 72804 182454 73404 217898
rect 72804 182218 72986 182454
rect 73222 182218 73404 182454
rect 72804 182134 73404 182218
rect 72804 181898 72986 182134
rect 73222 181898 73404 182134
rect 72804 146454 73404 181898
rect 72804 146218 72986 146454
rect 73222 146218 73404 146454
rect 72804 146134 73404 146218
rect 72804 145898 72986 146134
rect 73222 145898 73404 146134
rect 72804 110454 73404 145898
rect 72804 110218 72986 110454
rect 73222 110218 73404 110454
rect 72804 110134 73404 110218
rect 72804 109898 72986 110134
rect 73222 109898 73404 110134
rect 72804 74454 73404 109898
rect 72804 74218 72986 74454
rect 73222 74218 73404 74454
rect 72804 74134 73404 74218
rect 72804 73898 72986 74134
rect 73222 73898 73404 74134
rect 72804 38454 73404 73898
rect 72804 38218 72986 38454
rect 73222 38218 73404 38454
rect 72804 38134 73404 38218
rect 72804 37898 72986 38134
rect 73222 37898 73404 38134
rect 72804 2454 73404 37898
rect 72804 2218 72986 2454
rect 73222 2218 73404 2454
rect 72804 2134 73404 2218
rect 72804 1898 72986 2134
rect 73222 1898 73404 2134
rect 72804 -346 73404 1898
rect 72804 -582 72986 -346
rect 73222 -582 73404 -346
rect 72804 -666 73404 -582
rect 72804 -902 72986 -666
rect 73222 -902 73404 -666
rect 72804 -1864 73404 -902
rect 76404 294054 77004 317000
rect 76404 293818 76586 294054
rect 76822 293818 77004 294054
rect 76404 293734 77004 293818
rect 76404 293498 76586 293734
rect 76822 293498 77004 293734
rect 76404 258054 77004 293498
rect 76404 257818 76586 258054
rect 76822 257818 77004 258054
rect 76404 257734 77004 257818
rect 76404 257498 76586 257734
rect 76822 257498 77004 257734
rect 76404 222054 77004 257498
rect 76404 221818 76586 222054
rect 76822 221818 77004 222054
rect 76404 221734 77004 221818
rect 76404 221498 76586 221734
rect 76822 221498 77004 221734
rect 76404 186054 77004 221498
rect 76404 185818 76586 186054
rect 76822 185818 77004 186054
rect 76404 185734 77004 185818
rect 76404 185498 76586 185734
rect 76822 185498 77004 185734
rect 76404 150054 77004 185498
rect 76404 149818 76586 150054
rect 76822 149818 77004 150054
rect 76404 149734 77004 149818
rect 76404 149498 76586 149734
rect 76822 149498 77004 149734
rect 76404 114054 77004 149498
rect 76404 113818 76586 114054
rect 76822 113818 77004 114054
rect 76404 113734 77004 113818
rect 76404 113498 76586 113734
rect 76822 113498 77004 113734
rect 76404 78054 77004 113498
rect 76404 77818 76586 78054
rect 76822 77818 77004 78054
rect 76404 77734 77004 77818
rect 76404 77498 76586 77734
rect 76822 77498 77004 77734
rect 76404 42054 77004 77498
rect 76404 41818 76586 42054
rect 76822 41818 77004 42054
rect 76404 41734 77004 41818
rect 76404 41498 76586 41734
rect 76822 41498 77004 41734
rect 76404 6054 77004 41498
rect 76404 5818 76586 6054
rect 76822 5818 77004 6054
rect 76404 5734 77004 5818
rect 76404 5498 76586 5734
rect 76822 5498 77004 5734
rect 76404 -2226 77004 5498
rect 76404 -2462 76586 -2226
rect 76822 -2462 77004 -2226
rect 76404 -2546 77004 -2462
rect 76404 -2782 76586 -2546
rect 76822 -2782 77004 -2546
rect 76404 -3744 77004 -2782
rect 80004 297654 80604 317000
rect 80004 297418 80186 297654
rect 80422 297418 80604 297654
rect 80004 297334 80604 297418
rect 80004 297098 80186 297334
rect 80422 297098 80604 297334
rect 80004 261654 80604 297098
rect 80004 261418 80186 261654
rect 80422 261418 80604 261654
rect 80004 261334 80604 261418
rect 80004 261098 80186 261334
rect 80422 261098 80604 261334
rect 80004 225654 80604 261098
rect 80004 225418 80186 225654
rect 80422 225418 80604 225654
rect 80004 225334 80604 225418
rect 80004 225098 80186 225334
rect 80422 225098 80604 225334
rect 80004 189654 80604 225098
rect 80004 189418 80186 189654
rect 80422 189418 80604 189654
rect 80004 189334 80604 189418
rect 80004 189098 80186 189334
rect 80422 189098 80604 189334
rect 80004 153654 80604 189098
rect 80004 153418 80186 153654
rect 80422 153418 80604 153654
rect 80004 153334 80604 153418
rect 80004 153098 80186 153334
rect 80422 153098 80604 153334
rect 80004 117654 80604 153098
rect 80004 117418 80186 117654
rect 80422 117418 80604 117654
rect 80004 117334 80604 117418
rect 80004 117098 80186 117334
rect 80422 117098 80604 117334
rect 80004 81654 80604 117098
rect 80004 81418 80186 81654
rect 80422 81418 80604 81654
rect 80004 81334 80604 81418
rect 80004 81098 80186 81334
rect 80422 81098 80604 81334
rect 80004 45654 80604 81098
rect 80004 45418 80186 45654
rect 80422 45418 80604 45654
rect 80004 45334 80604 45418
rect 80004 45098 80186 45334
rect 80422 45098 80604 45334
rect 80004 9654 80604 45098
rect 80004 9418 80186 9654
rect 80422 9418 80604 9654
rect 80004 9334 80604 9418
rect 80004 9098 80186 9334
rect 80422 9098 80604 9334
rect 80004 -4106 80604 9098
rect 80004 -4342 80186 -4106
rect 80422 -4342 80604 -4106
rect 80004 -4426 80604 -4342
rect 80004 -4662 80186 -4426
rect 80422 -4662 80604 -4426
rect 80004 -5624 80604 -4662
rect 83604 301254 84204 317000
rect 83604 301018 83786 301254
rect 84022 301018 84204 301254
rect 83604 300934 84204 301018
rect 83604 300698 83786 300934
rect 84022 300698 84204 300934
rect 83604 265254 84204 300698
rect 83604 265018 83786 265254
rect 84022 265018 84204 265254
rect 83604 264934 84204 265018
rect 83604 264698 83786 264934
rect 84022 264698 84204 264934
rect 83604 229254 84204 264698
rect 83604 229018 83786 229254
rect 84022 229018 84204 229254
rect 83604 228934 84204 229018
rect 83604 228698 83786 228934
rect 84022 228698 84204 228934
rect 83604 193254 84204 228698
rect 83604 193018 83786 193254
rect 84022 193018 84204 193254
rect 83604 192934 84204 193018
rect 83604 192698 83786 192934
rect 84022 192698 84204 192934
rect 83604 157254 84204 192698
rect 83604 157018 83786 157254
rect 84022 157018 84204 157254
rect 83604 156934 84204 157018
rect 83604 156698 83786 156934
rect 84022 156698 84204 156934
rect 83604 121254 84204 156698
rect 83604 121018 83786 121254
rect 84022 121018 84204 121254
rect 83604 120934 84204 121018
rect 83604 120698 83786 120934
rect 84022 120698 84204 120934
rect 83604 85254 84204 120698
rect 83604 85018 83786 85254
rect 84022 85018 84204 85254
rect 83604 84934 84204 85018
rect 83604 84698 83786 84934
rect 84022 84698 84204 84934
rect 83604 49254 84204 84698
rect 83604 49018 83786 49254
rect 84022 49018 84204 49254
rect 83604 48934 84204 49018
rect 83604 48698 83786 48934
rect 84022 48698 84204 48934
rect 83604 13254 84204 48698
rect 83604 13018 83786 13254
rect 84022 13018 84204 13254
rect 83604 12934 84204 13018
rect 83604 12698 83786 12934
rect 84022 12698 84204 12934
rect 65604 -7162 65786 -6926
rect 66022 -7162 66204 -6926
rect 65604 -7246 66204 -7162
rect 65604 -7482 65786 -7246
rect 66022 -7482 66204 -7246
rect 65604 -7504 66204 -7482
rect 83604 -5986 84204 12698
rect 90804 308454 91404 317000
rect 90804 308218 90986 308454
rect 91222 308218 91404 308454
rect 90804 308134 91404 308218
rect 90804 307898 90986 308134
rect 91222 307898 91404 308134
rect 90804 272454 91404 307898
rect 90804 272218 90986 272454
rect 91222 272218 91404 272454
rect 90804 272134 91404 272218
rect 90804 271898 90986 272134
rect 91222 271898 91404 272134
rect 90804 236454 91404 271898
rect 90804 236218 90986 236454
rect 91222 236218 91404 236454
rect 90804 236134 91404 236218
rect 90804 235898 90986 236134
rect 91222 235898 91404 236134
rect 90804 200454 91404 235898
rect 90804 200218 90986 200454
rect 91222 200218 91404 200454
rect 90804 200134 91404 200218
rect 90804 199898 90986 200134
rect 91222 199898 91404 200134
rect 90804 164454 91404 199898
rect 90804 164218 90986 164454
rect 91222 164218 91404 164454
rect 90804 164134 91404 164218
rect 90804 163898 90986 164134
rect 91222 163898 91404 164134
rect 90804 128454 91404 163898
rect 90804 128218 90986 128454
rect 91222 128218 91404 128454
rect 90804 128134 91404 128218
rect 90804 127898 90986 128134
rect 91222 127898 91404 128134
rect 90804 92454 91404 127898
rect 90804 92218 90986 92454
rect 91222 92218 91404 92454
rect 90804 92134 91404 92218
rect 90804 91898 90986 92134
rect 91222 91898 91404 92134
rect 90804 56454 91404 91898
rect 90804 56218 90986 56454
rect 91222 56218 91404 56454
rect 90804 56134 91404 56218
rect 90804 55898 90986 56134
rect 91222 55898 91404 56134
rect 90804 20454 91404 55898
rect 90804 20218 90986 20454
rect 91222 20218 91404 20454
rect 90804 20134 91404 20218
rect 90804 19898 90986 20134
rect 91222 19898 91404 20134
rect 90804 -1286 91404 19898
rect 90804 -1522 90986 -1286
rect 91222 -1522 91404 -1286
rect 90804 -1606 91404 -1522
rect 90804 -1842 90986 -1606
rect 91222 -1842 91404 -1606
rect 90804 -1864 91404 -1842
rect 94404 312054 95004 317000
rect 94404 311818 94586 312054
rect 94822 311818 95004 312054
rect 94404 311734 95004 311818
rect 94404 311498 94586 311734
rect 94822 311498 95004 311734
rect 94404 276054 95004 311498
rect 94404 275818 94586 276054
rect 94822 275818 95004 276054
rect 94404 275734 95004 275818
rect 94404 275498 94586 275734
rect 94822 275498 95004 275734
rect 94404 240054 95004 275498
rect 94404 239818 94586 240054
rect 94822 239818 95004 240054
rect 94404 239734 95004 239818
rect 94404 239498 94586 239734
rect 94822 239498 95004 239734
rect 94404 204054 95004 239498
rect 94404 203818 94586 204054
rect 94822 203818 95004 204054
rect 94404 203734 95004 203818
rect 94404 203498 94586 203734
rect 94822 203498 95004 203734
rect 94404 168054 95004 203498
rect 94404 167818 94586 168054
rect 94822 167818 95004 168054
rect 94404 167734 95004 167818
rect 94404 167498 94586 167734
rect 94822 167498 95004 167734
rect 94404 132054 95004 167498
rect 94404 131818 94586 132054
rect 94822 131818 95004 132054
rect 94404 131734 95004 131818
rect 94404 131498 94586 131734
rect 94822 131498 95004 131734
rect 94404 96054 95004 131498
rect 94404 95818 94586 96054
rect 94822 95818 95004 96054
rect 94404 95734 95004 95818
rect 94404 95498 94586 95734
rect 94822 95498 95004 95734
rect 94404 60054 95004 95498
rect 94404 59818 94586 60054
rect 94822 59818 95004 60054
rect 94404 59734 95004 59818
rect 94404 59498 94586 59734
rect 94822 59498 95004 59734
rect 94404 24054 95004 59498
rect 94404 23818 94586 24054
rect 94822 23818 95004 24054
rect 94404 23734 95004 23818
rect 94404 23498 94586 23734
rect 94822 23498 95004 23734
rect 94404 -3166 95004 23498
rect 94404 -3402 94586 -3166
rect 94822 -3402 95004 -3166
rect 94404 -3486 95004 -3402
rect 94404 -3722 94586 -3486
rect 94822 -3722 95004 -3486
rect 94404 -3744 95004 -3722
rect 98004 315654 98604 317000
rect 98004 315418 98186 315654
rect 98422 315418 98604 315654
rect 98004 315334 98604 315418
rect 98004 315098 98186 315334
rect 98422 315098 98604 315334
rect 98004 279654 98604 315098
rect 98004 279418 98186 279654
rect 98422 279418 98604 279654
rect 98004 279334 98604 279418
rect 98004 279098 98186 279334
rect 98422 279098 98604 279334
rect 98004 243654 98604 279098
rect 98004 243418 98186 243654
rect 98422 243418 98604 243654
rect 98004 243334 98604 243418
rect 98004 243098 98186 243334
rect 98422 243098 98604 243334
rect 98004 207654 98604 243098
rect 98004 207418 98186 207654
rect 98422 207418 98604 207654
rect 98004 207334 98604 207418
rect 98004 207098 98186 207334
rect 98422 207098 98604 207334
rect 98004 171654 98604 207098
rect 98004 171418 98186 171654
rect 98422 171418 98604 171654
rect 98004 171334 98604 171418
rect 98004 171098 98186 171334
rect 98422 171098 98604 171334
rect 98004 135654 98604 171098
rect 98004 135418 98186 135654
rect 98422 135418 98604 135654
rect 98004 135334 98604 135418
rect 98004 135098 98186 135334
rect 98422 135098 98604 135334
rect 98004 99654 98604 135098
rect 98004 99418 98186 99654
rect 98422 99418 98604 99654
rect 98004 99334 98604 99418
rect 98004 99098 98186 99334
rect 98422 99098 98604 99334
rect 98004 63654 98604 99098
rect 98004 63418 98186 63654
rect 98422 63418 98604 63654
rect 98004 63334 98604 63418
rect 98004 63098 98186 63334
rect 98422 63098 98604 63334
rect 98004 27654 98604 63098
rect 98004 27418 98186 27654
rect 98422 27418 98604 27654
rect 98004 27334 98604 27418
rect 98004 27098 98186 27334
rect 98422 27098 98604 27334
rect 98004 -5046 98604 27098
rect 98004 -5282 98186 -5046
rect 98422 -5282 98604 -5046
rect 98004 -5366 98604 -5282
rect 98004 -5602 98186 -5366
rect 98422 -5602 98604 -5366
rect 98004 -5624 98604 -5602
rect 101604 283254 102204 317000
rect 101604 283018 101786 283254
rect 102022 283018 102204 283254
rect 101604 282934 102204 283018
rect 101604 282698 101786 282934
rect 102022 282698 102204 282934
rect 101604 247254 102204 282698
rect 101604 247018 101786 247254
rect 102022 247018 102204 247254
rect 101604 246934 102204 247018
rect 101604 246698 101786 246934
rect 102022 246698 102204 246934
rect 101604 211254 102204 246698
rect 101604 211018 101786 211254
rect 102022 211018 102204 211254
rect 101604 210934 102204 211018
rect 101604 210698 101786 210934
rect 102022 210698 102204 210934
rect 101604 175254 102204 210698
rect 101604 175018 101786 175254
rect 102022 175018 102204 175254
rect 101604 174934 102204 175018
rect 101604 174698 101786 174934
rect 102022 174698 102204 174934
rect 101604 139254 102204 174698
rect 101604 139018 101786 139254
rect 102022 139018 102204 139254
rect 101604 138934 102204 139018
rect 101604 138698 101786 138934
rect 102022 138698 102204 138934
rect 101604 103254 102204 138698
rect 101604 103018 101786 103254
rect 102022 103018 102204 103254
rect 101604 102934 102204 103018
rect 101604 102698 101786 102934
rect 102022 102698 102204 102934
rect 101604 67254 102204 102698
rect 101604 67018 101786 67254
rect 102022 67018 102204 67254
rect 101604 66934 102204 67018
rect 101604 66698 101786 66934
rect 102022 66698 102204 66934
rect 101604 31254 102204 66698
rect 101604 31018 101786 31254
rect 102022 31018 102204 31254
rect 101604 30934 102204 31018
rect 101604 30698 101786 30934
rect 102022 30698 102204 30934
rect 83604 -6222 83786 -5986
rect 84022 -6222 84204 -5986
rect 83604 -6306 84204 -6222
rect 83604 -6542 83786 -6306
rect 84022 -6542 84204 -6306
rect 83604 -7504 84204 -6542
rect 101604 -6926 102204 30698
rect 108804 290454 109404 317000
rect 108804 290218 108986 290454
rect 109222 290218 109404 290454
rect 108804 290134 109404 290218
rect 108804 289898 108986 290134
rect 109222 289898 109404 290134
rect 108804 254454 109404 289898
rect 108804 254218 108986 254454
rect 109222 254218 109404 254454
rect 108804 254134 109404 254218
rect 108804 253898 108986 254134
rect 109222 253898 109404 254134
rect 108804 218454 109404 253898
rect 108804 218218 108986 218454
rect 109222 218218 109404 218454
rect 108804 218134 109404 218218
rect 108804 217898 108986 218134
rect 109222 217898 109404 218134
rect 108804 182454 109404 217898
rect 108804 182218 108986 182454
rect 109222 182218 109404 182454
rect 108804 182134 109404 182218
rect 108804 181898 108986 182134
rect 109222 181898 109404 182134
rect 108804 146454 109404 181898
rect 108804 146218 108986 146454
rect 109222 146218 109404 146454
rect 108804 146134 109404 146218
rect 108804 145898 108986 146134
rect 109222 145898 109404 146134
rect 108804 110454 109404 145898
rect 108804 110218 108986 110454
rect 109222 110218 109404 110454
rect 108804 110134 109404 110218
rect 108804 109898 108986 110134
rect 109222 109898 109404 110134
rect 108804 74454 109404 109898
rect 108804 74218 108986 74454
rect 109222 74218 109404 74454
rect 108804 74134 109404 74218
rect 108804 73898 108986 74134
rect 109222 73898 109404 74134
rect 108804 38454 109404 73898
rect 108804 38218 108986 38454
rect 109222 38218 109404 38454
rect 108804 38134 109404 38218
rect 108804 37898 108986 38134
rect 109222 37898 109404 38134
rect 108804 2454 109404 37898
rect 108804 2218 108986 2454
rect 109222 2218 109404 2454
rect 108804 2134 109404 2218
rect 108804 1898 108986 2134
rect 109222 1898 109404 2134
rect 108804 -346 109404 1898
rect 108804 -582 108986 -346
rect 109222 -582 109404 -346
rect 108804 -666 109404 -582
rect 108804 -902 108986 -666
rect 109222 -902 109404 -666
rect 108804 -1864 109404 -902
rect 112404 294054 113004 317000
rect 112404 293818 112586 294054
rect 112822 293818 113004 294054
rect 112404 293734 113004 293818
rect 112404 293498 112586 293734
rect 112822 293498 113004 293734
rect 112404 258054 113004 293498
rect 112404 257818 112586 258054
rect 112822 257818 113004 258054
rect 112404 257734 113004 257818
rect 112404 257498 112586 257734
rect 112822 257498 113004 257734
rect 112404 222054 113004 257498
rect 112404 221818 112586 222054
rect 112822 221818 113004 222054
rect 112404 221734 113004 221818
rect 112404 221498 112586 221734
rect 112822 221498 113004 221734
rect 112404 186054 113004 221498
rect 112404 185818 112586 186054
rect 112822 185818 113004 186054
rect 112404 185734 113004 185818
rect 112404 185498 112586 185734
rect 112822 185498 113004 185734
rect 112404 150054 113004 185498
rect 112404 149818 112586 150054
rect 112822 149818 113004 150054
rect 112404 149734 113004 149818
rect 112404 149498 112586 149734
rect 112822 149498 113004 149734
rect 112404 114054 113004 149498
rect 112404 113818 112586 114054
rect 112822 113818 113004 114054
rect 112404 113734 113004 113818
rect 112404 113498 112586 113734
rect 112822 113498 113004 113734
rect 112404 78054 113004 113498
rect 112404 77818 112586 78054
rect 112822 77818 113004 78054
rect 112404 77734 113004 77818
rect 112404 77498 112586 77734
rect 112822 77498 113004 77734
rect 112404 42054 113004 77498
rect 112404 41818 112586 42054
rect 112822 41818 113004 42054
rect 112404 41734 113004 41818
rect 112404 41498 112586 41734
rect 112822 41498 113004 41734
rect 112404 6054 113004 41498
rect 112404 5818 112586 6054
rect 112822 5818 113004 6054
rect 112404 5734 113004 5818
rect 112404 5498 112586 5734
rect 112822 5498 113004 5734
rect 112404 -2226 113004 5498
rect 112404 -2462 112586 -2226
rect 112822 -2462 113004 -2226
rect 112404 -2546 113004 -2462
rect 112404 -2782 112586 -2546
rect 112822 -2782 113004 -2546
rect 112404 -3744 113004 -2782
rect 116004 297654 116604 317000
rect 116004 297418 116186 297654
rect 116422 297418 116604 297654
rect 116004 297334 116604 297418
rect 116004 297098 116186 297334
rect 116422 297098 116604 297334
rect 116004 261654 116604 297098
rect 116004 261418 116186 261654
rect 116422 261418 116604 261654
rect 116004 261334 116604 261418
rect 116004 261098 116186 261334
rect 116422 261098 116604 261334
rect 116004 225654 116604 261098
rect 116004 225418 116186 225654
rect 116422 225418 116604 225654
rect 116004 225334 116604 225418
rect 116004 225098 116186 225334
rect 116422 225098 116604 225334
rect 116004 189654 116604 225098
rect 116004 189418 116186 189654
rect 116422 189418 116604 189654
rect 116004 189334 116604 189418
rect 116004 189098 116186 189334
rect 116422 189098 116604 189334
rect 116004 153654 116604 189098
rect 116004 153418 116186 153654
rect 116422 153418 116604 153654
rect 116004 153334 116604 153418
rect 116004 153098 116186 153334
rect 116422 153098 116604 153334
rect 116004 117654 116604 153098
rect 116004 117418 116186 117654
rect 116422 117418 116604 117654
rect 116004 117334 116604 117418
rect 116004 117098 116186 117334
rect 116422 117098 116604 117334
rect 116004 81654 116604 117098
rect 116004 81418 116186 81654
rect 116422 81418 116604 81654
rect 116004 81334 116604 81418
rect 116004 81098 116186 81334
rect 116422 81098 116604 81334
rect 116004 45654 116604 81098
rect 116004 45418 116186 45654
rect 116422 45418 116604 45654
rect 116004 45334 116604 45418
rect 116004 45098 116186 45334
rect 116422 45098 116604 45334
rect 116004 9654 116604 45098
rect 116004 9418 116186 9654
rect 116422 9418 116604 9654
rect 116004 9334 116604 9418
rect 116004 9098 116186 9334
rect 116422 9098 116604 9334
rect 116004 -4106 116604 9098
rect 116004 -4342 116186 -4106
rect 116422 -4342 116604 -4106
rect 116004 -4426 116604 -4342
rect 116004 -4662 116186 -4426
rect 116422 -4662 116604 -4426
rect 116004 -5624 116604 -4662
rect 119604 301254 120204 317000
rect 119604 301018 119786 301254
rect 120022 301018 120204 301254
rect 119604 300934 120204 301018
rect 119604 300698 119786 300934
rect 120022 300698 120204 300934
rect 119604 265254 120204 300698
rect 119604 265018 119786 265254
rect 120022 265018 120204 265254
rect 119604 264934 120204 265018
rect 119604 264698 119786 264934
rect 120022 264698 120204 264934
rect 119604 229254 120204 264698
rect 119604 229018 119786 229254
rect 120022 229018 120204 229254
rect 119604 228934 120204 229018
rect 119604 228698 119786 228934
rect 120022 228698 120204 228934
rect 119604 193254 120204 228698
rect 119604 193018 119786 193254
rect 120022 193018 120204 193254
rect 119604 192934 120204 193018
rect 119604 192698 119786 192934
rect 120022 192698 120204 192934
rect 119604 157254 120204 192698
rect 119604 157018 119786 157254
rect 120022 157018 120204 157254
rect 119604 156934 120204 157018
rect 119604 156698 119786 156934
rect 120022 156698 120204 156934
rect 119604 121254 120204 156698
rect 119604 121018 119786 121254
rect 120022 121018 120204 121254
rect 119604 120934 120204 121018
rect 119604 120698 119786 120934
rect 120022 120698 120204 120934
rect 119604 85254 120204 120698
rect 119604 85018 119786 85254
rect 120022 85018 120204 85254
rect 119604 84934 120204 85018
rect 119604 84698 119786 84934
rect 120022 84698 120204 84934
rect 119604 49254 120204 84698
rect 119604 49018 119786 49254
rect 120022 49018 120204 49254
rect 119604 48934 120204 49018
rect 119604 48698 119786 48934
rect 120022 48698 120204 48934
rect 119604 13254 120204 48698
rect 119604 13018 119786 13254
rect 120022 13018 120204 13254
rect 119604 12934 120204 13018
rect 119604 12698 119786 12934
rect 120022 12698 120204 12934
rect 101604 -7162 101786 -6926
rect 102022 -7162 102204 -6926
rect 101604 -7246 102204 -7162
rect 101604 -7482 101786 -7246
rect 102022 -7482 102204 -7246
rect 101604 -7504 102204 -7482
rect 119604 -5986 120204 12698
rect 126804 308454 127404 317000
rect 126804 308218 126986 308454
rect 127222 308218 127404 308454
rect 126804 308134 127404 308218
rect 126804 307898 126986 308134
rect 127222 307898 127404 308134
rect 126804 272454 127404 307898
rect 126804 272218 126986 272454
rect 127222 272218 127404 272454
rect 126804 272134 127404 272218
rect 126804 271898 126986 272134
rect 127222 271898 127404 272134
rect 126804 236454 127404 271898
rect 126804 236218 126986 236454
rect 127222 236218 127404 236454
rect 126804 236134 127404 236218
rect 126804 235898 126986 236134
rect 127222 235898 127404 236134
rect 126804 200454 127404 235898
rect 126804 200218 126986 200454
rect 127222 200218 127404 200454
rect 126804 200134 127404 200218
rect 126804 199898 126986 200134
rect 127222 199898 127404 200134
rect 126804 164454 127404 199898
rect 126804 164218 126986 164454
rect 127222 164218 127404 164454
rect 126804 164134 127404 164218
rect 126804 163898 126986 164134
rect 127222 163898 127404 164134
rect 126804 128454 127404 163898
rect 126804 128218 126986 128454
rect 127222 128218 127404 128454
rect 126804 128134 127404 128218
rect 126804 127898 126986 128134
rect 127222 127898 127404 128134
rect 126804 92454 127404 127898
rect 126804 92218 126986 92454
rect 127222 92218 127404 92454
rect 126804 92134 127404 92218
rect 126804 91898 126986 92134
rect 127222 91898 127404 92134
rect 126804 56454 127404 91898
rect 126804 56218 126986 56454
rect 127222 56218 127404 56454
rect 126804 56134 127404 56218
rect 126804 55898 126986 56134
rect 127222 55898 127404 56134
rect 126804 20454 127404 55898
rect 126804 20218 126986 20454
rect 127222 20218 127404 20454
rect 126804 20134 127404 20218
rect 126804 19898 126986 20134
rect 127222 19898 127404 20134
rect 126804 -1286 127404 19898
rect 126804 -1522 126986 -1286
rect 127222 -1522 127404 -1286
rect 126804 -1606 127404 -1522
rect 126804 -1842 126986 -1606
rect 127222 -1842 127404 -1606
rect 126804 -1864 127404 -1842
rect 130404 312054 131004 317000
rect 130404 311818 130586 312054
rect 130822 311818 131004 312054
rect 130404 311734 131004 311818
rect 130404 311498 130586 311734
rect 130822 311498 131004 311734
rect 130404 276054 131004 311498
rect 130404 275818 130586 276054
rect 130822 275818 131004 276054
rect 130404 275734 131004 275818
rect 130404 275498 130586 275734
rect 130822 275498 131004 275734
rect 130404 240054 131004 275498
rect 130404 239818 130586 240054
rect 130822 239818 131004 240054
rect 130404 239734 131004 239818
rect 130404 239498 130586 239734
rect 130822 239498 131004 239734
rect 130404 204054 131004 239498
rect 130404 203818 130586 204054
rect 130822 203818 131004 204054
rect 130404 203734 131004 203818
rect 130404 203498 130586 203734
rect 130822 203498 131004 203734
rect 130404 168054 131004 203498
rect 130404 167818 130586 168054
rect 130822 167818 131004 168054
rect 130404 167734 131004 167818
rect 130404 167498 130586 167734
rect 130822 167498 131004 167734
rect 130404 132054 131004 167498
rect 130404 131818 130586 132054
rect 130822 131818 131004 132054
rect 130404 131734 131004 131818
rect 130404 131498 130586 131734
rect 130822 131498 131004 131734
rect 130404 96054 131004 131498
rect 130404 95818 130586 96054
rect 130822 95818 131004 96054
rect 130404 95734 131004 95818
rect 130404 95498 130586 95734
rect 130822 95498 131004 95734
rect 130404 60054 131004 95498
rect 130404 59818 130586 60054
rect 130822 59818 131004 60054
rect 130404 59734 131004 59818
rect 130404 59498 130586 59734
rect 130822 59498 131004 59734
rect 130404 24054 131004 59498
rect 130404 23818 130586 24054
rect 130822 23818 131004 24054
rect 130404 23734 131004 23818
rect 130404 23498 130586 23734
rect 130822 23498 131004 23734
rect 130404 -3166 131004 23498
rect 130404 -3402 130586 -3166
rect 130822 -3402 131004 -3166
rect 130404 -3486 131004 -3402
rect 130404 -3722 130586 -3486
rect 130822 -3722 131004 -3486
rect 130404 -3744 131004 -3722
rect 134004 315654 134604 317000
rect 134004 315418 134186 315654
rect 134422 315418 134604 315654
rect 134004 315334 134604 315418
rect 134004 315098 134186 315334
rect 134422 315098 134604 315334
rect 134004 279654 134604 315098
rect 134004 279418 134186 279654
rect 134422 279418 134604 279654
rect 134004 279334 134604 279418
rect 134004 279098 134186 279334
rect 134422 279098 134604 279334
rect 134004 243654 134604 279098
rect 134004 243418 134186 243654
rect 134422 243418 134604 243654
rect 134004 243334 134604 243418
rect 134004 243098 134186 243334
rect 134422 243098 134604 243334
rect 134004 207654 134604 243098
rect 134004 207418 134186 207654
rect 134422 207418 134604 207654
rect 134004 207334 134604 207418
rect 134004 207098 134186 207334
rect 134422 207098 134604 207334
rect 134004 171654 134604 207098
rect 134004 171418 134186 171654
rect 134422 171418 134604 171654
rect 134004 171334 134604 171418
rect 134004 171098 134186 171334
rect 134422 171098 134604 171334
rect 134004 135654 134604 171098
rect 134004 135418 134186 135654
rect 134422 135418 134604 135654
rect 134004 135334 134604 135418
rect 134004 135098 134186 135334
rect 134422 135098 134604 135334
rect 134004 99654 134604 135098
rect 134004 99418 134186 99654
rect 134422 99418 134604 99654
rect 134004 99334 134604 99418
rect 134004 99098 134186 99334
rect 134422 99098 134604 99334
rect 134004 63654 134604 99098
rect 134004 63418 134186 63654
rect 134422 63418 134604 63654
rect 134004 63334 134604 63418
rect 134004 63098 134186 63334
rect 134422 63098 134604 63334
rect 134004 27654 134604 63098
rect 134004 27418 134186 27654
rect 134422 27418 134604 27654
rect 134004 27334 134604 27418
rect 134004 27098 134186 27334
rect 134422 27098 134604 27334
rect 134004 -5046 134604 27098
rect 134004 -5282 134186 -5046
rect 134422 -5282 134604 -5046
rect 134004 -5366 134604 -5282
rect 134004 -5602 134186 -5366
rect 134422 -5602 134604 -5366
rect 134004 -5624 134604 -5602
rect 137604 283254 138204 317000
rect 137604 283018 137786 283254
rect 138022 283018 138204 283254
rect 137604 282934 138204 283018
rect 137604 282698 137786 282934
rect 138022 282698 138204 282934
rect 137604 247254 138204 282698
rect 137604 247018 137786 247254
rect 138022 247018 138204 247254
rect 137604 246934 138204 247018
rect 137604 246698 137786 246934
rect 138022 246698 138204 246934
rect 137604 211254 138204 246698
rect 137604 211018 137786 211254
rect 138022 211018 138204 211254
rect 137604 210934 138204 211018
rect 137604 210698 137786 210934
rect 138022 210698 138204 210934
rect 137604 175254 138204 210698
rect 137604 175018 137786 175254
rect 138022 175018 138204 175254
rect 137604 174934 138204 175018
rect 137604 174698 137786 174934
rect 138022 174698 138204 174934
rect 137604 139254 138204 174698
rect 137604 139018 137786 139254
rect 138022 139018 138204 139254
rect 137604 138934 138204 139018
rect 137604 138698 137786 138934
rect 138022 138698 138204 138934
rect 137604 103254 138204 138698
rect 137604 103018 137786 103254
rect 138022 103018 138204 103254
rect 137604 102934 138204 103018
rect 137604 102698 137786 102934
rect 138022 102698 138204 102934
rect 137604 67254 138204 102698
rect 137604 67018 137786 67254
rect 138022 67018 138204 67254
rect 137604 66934 138204 67018
rect 137604 66698 137786 66934
rect 138022 66698 138204 66934
rect 137604 31254 138204 66698
rect 137604 31018 137786 31254
rect 138022 31018 138204 31254
rect 137604 30934 138204 31018
rect 137604 30698 137786 30934
rect 138022 30698 138204 30934
rect 119604 -6222 119786 -5986
rect 120022 -6222 120204 -5986
rect 119604 -6306 120204 -6222
rect 119604 -6542 119786 -6306
rect 120022 -6542 120204 -6306
rect 119604 -7504 120204 -6542
rect 137604 -6926 138204 30698
rect 144804 290454 145404 317000
rect 144804 290218 144986 290454
rect 145222 290218 145404 290454
rect 144804 290134 145404 290218
rect 144804 289898 144986 290134
rect 145222 289898 145404 290134
rect 144804 254454 145404 289898
rect 144804 254218 144986 254454
rect 145222 254218 145404 254454
rect 144804 254134 145404 254218
rect 144804 253898 144986 254134
rect 145222 253898 145404 254134
rect 144804 218454 145404 253898
rect 144804 218218 144986 218454
rect 145222 218218 145404 218454
rect 144804 218134 145404 218218
rect 144804 217898 144986 218134
rect 145222 217898 145404 218134
rect 144804 182454 145404 217898
rect 144804 182218 144986 182454
rect 145222 182218 145404 182454
rect 144804 182134 145404 182218
rect 144804 181898 144986 182134
rect 145222 181898 145404 182134
rect 144804 146454 145404 181898
rect 144804 146218 144986 146454
rect 145222 146218 145404 146454
rect 144804 146134 145404 146218
rect 144804 145898 144986 146134
rect 145222 145898 145404 146134
rect 144804 110454 145404 145898
rect 144804 110218 144986 110454
rect 145222 110218 145404 110454
rect 144804 110134 145404 110218
rect 144804 109898 144986 110134
rect 145222 109898 145404 110134
rect 144804 74454 145404 109898
rect 144804 74218 144986 74454
rect 145222 74218 145404 74454
rect 144804 74134 145404 74218
rect 144804 73898 144986 74134
rect 145222 73898 145404 74134
rect 144804 38454 145404 73898
rect 144804 38218 144986 38454
rect 145222 38218 145404 38454
rect 144804 38134 145404 38218
rect 144804 37898 144986 38134
rect 145222 37898 145404 38134
rect 144804 2454 145404 37898
rect 144804 2218 144986 2454
rect 145222 2218 145404 2454
rect 144804 2134 145404 2218
rect 144804 1898 144986 2134
rect 145222 1898 145404 2134
rect 144804 -346 145404 1898
rect 144804 -582 144986 -346
rect 145222 -582 145404 -346
rect 144804 -666 145404 -582
rect 144804 -902 144986 -666
rect 145222 -902 145404 -666
rect 144804 -1864 145404 -902
rect 148404 294054 149004 317000
rect 148404 293818 148586 294054
rect 148822 293818 149004 294054
rect 148404 293734 149004 293818
rect 148404 293498 148586 293734
rect 148822 293498 149004 293734
rect 148404 258054 149004 293498
rect 148404 257818 148586 258054
rect 148822 257818 149004 258054
rect 148404 257734 149004 257818
rect 148404 257498 148586 257734
rect 148822 257498 149004 257734
rect 148404 222054 149004 257498
rect 148404 221818 148586 222054
rect 148822 221818 149004 222054
rect 148404 221734 149004 221818
rect 148404 221498 148586 221734
rect 148822 221498 149004 221734
rect 148404 186054 149004 221498
rect 148404 185818 148586 186054
rect 148822 185818 149004 186054
rect 148404 185734 149004 185818
rect 148404 185498 148586 185734
rect 148822 185498 149004 185734
rect 148404 150054 149004 185498
rect 148404 149818 148586 150054
rect 148822 149818 149004 150054
rect 148404 149734 149004 149818
rect 148404 149498 148586 149734
rect 148822 149498 149004 149734
rect 148404 114054 149004 149498
rect 148404 113818 148586 114054
rect 148822 113818 149004 114054
rect 148404 113734 149004 113818
rect 148404 113498 148586 113734
rect 148822 113498 149004 113734
rect 148404 78054 149004 113498
rect 148404 77818 148586 78054
rect 148822 77818 149004 78054
rect 148404 77734 149004 77818
rect 148404 77498 148586 77734
rect 148822 77498 149004 77734
rect 148404 42054 149004 77498
rect 148404 41818 148586 42054
rect 148822 41818 149004 42054
rect 148404 41734 149004 41818
rect 148404 41498 148586 41734
rect 148822 41498 149004 41734
rect 148404 6054 149004 41498
rect 148404 5818 148586 6054
rect 148822 5818 149004 6054
rect 148404 5734 149004 5818
rect 148404 5498 148586 5734
rect 148822 5498 149004 5734
rect 148404 -2226 149004 5498
rect 148404 -2462 148586 -2226
rect 148822 -2462 149004 -2226
rect 148404 -2546 149004 -2462
rect 148404 -2782 148586 -2546
rect 148822 -2782 149004 -2546
rect 148404 -3744 149004 -2782
rect 152004 297654 152604 317000
rect 152004 297418 152186 297654
rect 152422 297418 152604 297654
rect 152004 297334 152604 297418
rect 152004 297098 152186 297334
rect 152422 297098 152604 297334
rect 152004 261654 152604 297098
rect 152004 261418 152186 261654
rect 152422 261418 152604 261654
rect 152004 261334 152604 261418
rect 152004 261098 152186 261334
rect 152422 261098 152604 261334
rect 152004 225654 152604 261098
rect 152004 225418 152186 225654
rect 152422 225418 152604 225654
rect 152004 225334 152604 225418
rect 152004 225098 152186 225334
rect 152422 225098 152604 225334
rect 152004 189654 152604 225098
rect 152004 189418 152186 189654
rect 152422 189418 152604 189654
rect 152004 189334 152604 189418
rect 152004 189098 152186 189334
rect 152422 189098 152604 189334
rect 152004 153654 152604 189098
rect 152004 153418 152186 153654
rect 152422 153418 152604 153654
rect 152004 153334 152604 153418
rect 152004 153098 152186 153334
rect 152422 153098 152604 153334
rect 152004 117654 152604 153098
rect 152004 117418 152186 117654
rect 152422 117418 152604 117654
rect 152004 117334 152604 117418
rect 152004 117098 152186 117334
rect 152422 117098 152604 117334
rect 152004 81654 152604 117098
rect 152004 81418 152186 81654
rect 152422 81418 152604 81654
rect 152004 81334 152604 81418
rect 152004 81098 152186 81334
rect 152422 81098 152604 81334
rect 152004 45654 152604 81098
rect 152004 45418 152186 45654
rect 152422 45418 152604 45654
rect 152004 45334 152604 45418
rect 152004 45098 152186 45334
rect 152422 45098 152604 45334
rect 152004 9654 152604 45098
rect 152004 9418 152186 9654
rect 152422 9418 152604 9654
rect 152004 9334 152604 9418
rect 152004 9098 152186 9334
rect 152422 9098 152604 9334
rect 152004 -4106 152604 9098
rect 152004 -4342 152186 -4106
rect 152422 -4342 152604 -4106
rect 152004 -4426 152604 -4342
rect 152004 -4662 152186 -4426
rect 152422 -4662 152604 -4426
rect 152004 -5624 152604 -4662
rect 155604 301254 156204 317000
rect 155604 301018 155786 301254
rect 156022 301018 156204 301254
rect 155604 300934 156204 301018
rect 155604 300698 155786 300934
rect 156022 300698 156204 300934
rect 155604 265254 156204 300698
rect 155604 265018 155786 265254
rect 156022 265018 156204 265254
rect 155604 264934 156204 265018
rect 155604 264698 155786 264934
rect 156022 264698 156204 264934
rect 155604 229254 156204 264698
rect 155604 229018 155786 229254
rect 156022 229018 156204 229254
rect 155604 228934 156204 229018
rect 155604 228698 155786 228934
rect 156022 228698 156204 228934
rect 155604 193254 156204 228698
rect 155604 193018 155786 193254
rect 156022 193018 156204 193254
rect 155604 192934 156204 193018
rect 155604 192698 155786 192934
rect 156022 192698 156204 192934
rect 155604 157254 156204 192698
rect 155604 157018 155786 157254
rect 156022 157018 156204 157254
rect 155604 156934 156204 157018
rect 155604 156698 155786 156934
rect 156022 156698 156204 156934
rect 155604 121254 156204 156698
rect 155604 121018 155786 121254
rect 156022 121018 156204 121254
rect 155604 120934 156204 121018
rect 155604 120698 155786 120934
rect 156022 120698 156204 120934
rect 155604 85254 156204 120698
rect 155604 85018 155786 85254
rect 156022 85018 156204 85254
rect 155604 84934 156204 85018
rect 155604 84698 155786 84934
rect 156022 84698 156204 84934
rect 155604 49254 156204 84698
rect 155604 49018 155786 49254
rect 156022 49018 156204 49254
rect 155604 48934 156204 49018
rect 155604 48698 155786 48934
rect 156022 48698 156204 48934
rect 155604 13254 156204 48698
rect 155604 13018 155786 13254
rect 156022 13018 156204 13254
rect 155604 12934 156204 13018
rect 155604 12698 155786 12934
rect 156022 12698 156204 12934
rect 137604 -7162 137786 -6926
rect 138022 -7162 138204 -6926
rect 137604 -7246 138204 -7162
rect 137604 -7482 137786 -7246
rect 138022 -7482 138204 -7246
rect 137604 -7504 138204 -7482
rect 155604 -5986 156204 12698
rect 162804 308454 163404 317000
rect 162804 308218 162986 308454
rect 163222 308218 163404 308454
rect 162804 308134 163404 308218
rect 162804 307898 162986 308134
rect 163222 307898 163404 308134
rect 162804 272454 163404 307898
rect 162804 272218 162986 272454
rect 163222 272218 163404 272454
rect 162804 272134 163404 272218
rect 162804 271898 162986 272134
rect 163222 271898 163404 272134
rect 162804 236454 163404 271898
rect 162804 236218 162986 236454
rect 163222 236218 163404 236454
rect 162804 236134 163404 236218
rect 162804 235898 162986 236134
rect 163222 235898 163404 236134
rect 162804 200454 163404 235898
rect 162804 200218 162986 200454
rect 163222 200218 163404 200454
rect 162804 200134 163404 200218
rect 162804 199898 162986 200134
rect 163222 199898 163404 200134
rect 162804 164454 163404 199898
rect 162804 164218 162986 164454
rect 163222 164218 163404 164454
rect 162804 164134 163404 164218
rect 162804 163898 162986 164134
rect 163222 163898 163404 164134
rect 162804 128454 163404 163898
rect 162804 128218 162986 128454
rect 163222 128218 163404 128454
rect 162804 128134 163404 128218
rect 162804 127898 162986 128134
rect 163222 127898 163404 128134
rect 162804 92454 163404 127898
rect 162804 92218 162986 92454
rect 163222 92218 163404 92454
rect 162804 92134 163404 92218
rect 162804 91898 162986 92134
rect 163222 91898 163404 92134
rect 162804 56454 163404 91898
rect 162804 56218 162986 56454
rect 163222 56218 163404 56454
rect 162804 56134 163404 56218
rect 162804 55898 162986 56134
rect 163222 55898 163404 56134
rect 162804 20454 163404 55898
rect 162804 20218 162986 20454
rect 163222 20218 163404 20454
rect 162804 20134 163404 20218
rect 162804 19898 162986 20134
rect 163222 19898 163404 20134
rect 162804 -1286 163404 19898
rect 162804 -1522 162986 -1286
rect 163222 -1522 163404 -1286
rect 162804 -1606 163404 -1522
rect 162804 -1842 162986 -1606
rect 163222 -1842 163404 -1606
rect 162804 -1864 163404 -1842
rect 166404 312054 167004 317000
rect 166404 311818 166586 312054
rect 166822 311818 167004 312054
rect 166404 311734 167004 311818
rect 166404 311498 166586 311734
rect 166822 311498 167004 311734
rect 166404 276054 167004 311498
rect 166404 275818 166586 276054
rect 166822 275818 167004 276054
rect 166404 275734 167004 275818
rect 166404 275498 166586 275734
rect 166822 275498 167004 275734
rect 166404 240054 167004 275498
rect 166404 239818 166586 240054
rect 166822 239818 167004 240054
rect 166404 239734 167004 239818
rect 166404 239498 166586 239734
rect 166822 239498 167004 239734
rect 166404 204054 167004 239498
rect 166404 203818 166586 204054
rect 166822 203818 167004 204054
rect 166404 203734 167004 203818
rect 166404 203498 166586 203734
rect 166822 203498 167004 203734
rect 166404 168054 167004 203498
rect 166404 167818 166586 168054
rect 166822 167818 167004 168054
rect 166404 167734 167004 167818
rect 166404 167498 166586 167734
rect 166822 167498 167004 167734
rect 166404 132054 167004 167498
rect 166404 131818 166586 132054
rect 166822 131818 167004 132054
rect 166404 131734 167004 131818
rect 166404 131498 166586 131734
rect 166822 131498 167004 131734
rect 166404 96054 167004 131498
rect 166404 95818 166586 96054
rect 166822 95818 167004 96054
rect 166404 95734 167004 95818
rect 166404 95498 166586 95734
rect 166822 95498 167004 95734
rect 166404 60054 167004 95498
rect 166404 59818 166586 60054
rect 166822 59818 167004 60054
rect 166404 59734 167004 59818
rect 166404 59498 166586 59734
rect 166822 59498 167004 59734
rect 166404 24054 167004 59498
rect 166404 23818 166586 24054
rect 166822 23818 167004 24054
rect 166404 23734 167004 23818
rect 166404 23498 166586 23734
rect 166822 23498 167004 23734
rect 166404 -3166 167004 23498
rect 166404 -3402 166586 -3166
rect 166822 -3402 167004 -3166
rect 166404 -3486 167004 -3402
rect 166404 -3722 166586 -3486
rect 166822 -3722 167004 -3486
rect 166404 -3744 167004 -3722
rect 170004 315654 170604 317000
rect 170004 315418 170186 315654
rect 170422 315418 170604 315654
rect 170004 315334 170604 315418
rect 170004 315098 170186 315334
rect 170422 315098 170604 315334
rect 170004 279654 170604 315098
rect 170004 279418 170186 279654
rect 170422 279418 170604 279654
rect 170004 279334 170604 279418
rect 170004 279098 170186 279334
rect 170422 279098 170604 279334
rect 170004 243654 170604 279098
rect 170004 243418 170186 243654
rect 170422 243418 170604 243654
rect 170004 243334 170604 243418
rect 170004 243098 170186 243334
rect 170422 243098 170604 243334
rect 170004 207654 170604 243098
rect 170004 207418 170186 207654
rect 170422 207418 170604 207654
rect 170004 207334 170604 207418
rect 170004 207098 170186 207334
rect 170422 207098 170604 207334
rect 170004 171654 170604 207098
rect 170004 171418 170186 171654
rect 170422 171418 170604 171654
rect 170004 171334 170604 171418
rect 170004 171098 170186 171334
rect 170422 171098 170604 171334
rect 170004 135654 170604 171098
rect 170004 135418 170186 135654
rect 170422 135418 170604 135654
rect 170004 135334 170604 135418
rect 170004 135098 170186 135334
rect 170422 135098 170604 135334
rect 170004 99654 170604 135098
rect 170004 99418 170186 99654
rect 170422 99418 170604 99654
rect 170004 99334 170604 99418
rect 170004 99098 170186 99334
rect 170422 99098 170604 99334
rect 170004 63654 170604 99098
rect 170004 63418 170186 63654
rect 170422 63418 170604 63654
rect 170004 63334 170604 63418
rect 170004 63098 170186 63334
rect 170422 63098 170604 63334
rect 170004 27654 170604 63098
rect 170004 27418 170186 27654
rect 170422 27418 170604 27654
rect 170004 27334 170604 27418
rect 170004 27098 170186 27334
rect 170422 27098 170604 27334
rect 170004 -5046 170604 27098
rect 170004 -5282 170186 -5046
rect 170422 -5282 170604 -5046
rect 170004 -5366 170604 -5282
rect 170004 -5602 170186 -5366
rect 170422 -5602 170604 -5366
rect 170004 -5624 170604 -5602
rect 173604 283254 174204 317000
rect 173604 283018 173786 283254
rect 174022 283018 174204 283254
rect 173604 282934 174204 283018
rect 173604 282698 173786 282934
rect 174022 282698 174204 282934
rect 173604 247254 174204 282698
rect 173604 247018 173786 247254
rect 174022 247018 174204 247254
rect 173604 246934 174204 247018
rect 173604 246698 173786 246934
rect 174022 246698 174204 246934
rect 173604 211254 174204 246698
rect 173604 211018 173786 211254
rect 174022 211018 174204 211254
rect 173604 210934 174204 211018
rect 173604 210698 173786 210934
rect 174022 210698 174204 210934
rect 173604 175254 174204 210698
rect 173604 175018 173786 175254
rect 174022 175018 174204 175254
rect 173604 174934 174204 175018
rect 173604 174698 173786 174934
rect 174022 174698 174204 174934
rect 173604 139254 174204 174698
rect 173604 139018 173786 139254
rect 174022 139018 174204 139254
rect 173604 138934 174204 139018
rect 173604 138698 173786 138934
rect 174022 138698 174204 138934
rect 173604 103254 174204 138698
rect 173604 103018 173786 103254
rect 174022 103018 174204 103254
rect 173604 102934 174204 103018
rect 173604 102698 173786 102934
rect 174022 102698 174204 102934
rect 173604 67254 174204 102698
rect 173604 67018 173786 67254
rect 174022 67018 174204 67254
rect 173604 66934 174204 67018
rect 173604 66698 173786 66934
rect 174022 66698 174204 66934
rect 173604 31254 174204 66698
rect 173604 31018 173786 31254
rect 174022 31018 174204 31254
rect 173604 30934 174204 31018
rect 173604 30698 173786 30934
rect 174022 30698 174204 30934
rect 155604 -6222 155786 -5986
rect 156022 -6222 156204 -5986
rect 155604 -6306 156204 -6222
rect 155604 -6542 155786 -6306
rect 156022 -6542 156204 -6306
rect 155604 -7504 156204 -6542
rect 173604 -6926 174204 30698
rect 180804 290454 181404 317000
rect 180804 290218 180986 290454
rect 181222 290218 181404 290454
rect 180804 290134 181404 290218
rect 180804 289898 180986 290134
rect 181222 289898 181404 290134
rect 180804 254454 181404 289898
rect 180804 254218 180986 254454
rect 181222 254218 181404 254454
rect 180804 254134 181404 254218
rect 180804 253898 180986 254134
rect 181222 253898 181404 254134
rect 180804 218454 181404 253898
rect 180804 218218 180986 218454
rect 181222 218218 181404 218454
rect 180804 218134 181404 218218
rect 180804 217898 180986 218134
rect 181222 217898 181404 218134
rect 180804 182454 181404 217898
rect 180804 182218 180986 182454
rect 181222 182218 181404 182454
rect 180804 182134 181404 182218
rect 180804 181898 180986 182134
rect 181222 181898 181404 182134
rect 180804 146454 181404 181898
rect 180804 146218 180986 146454
rect 181222 146218 181404 146454
rect 180804 146134 181404 146218
rect 180804 145898 180986 146134
rect 181222 145898 181404 146134
rect 180804 110454 181404 145898
rect 180804 110218 180986 110454
rect 181222 110218 181404 110454
rect 180804 110134 181404 110218
rect 180804 109898 180986 110134
rect 181222 109898 181404 110134
rect 180804 74454 181404 109898
rect 180804 74218 180986 74454
rect 181222 74218 181404 74454
rect 180804 74134 181404 74218
rect 180804 73898 180986 74134
rect 181222 73898 181404 74134
rect 180804 38454 181404 73898
rect 180804 38218 180986 38454
rect 181222 38218 181404 38454
rect 180804 38134 181404 38218
rect 180804 37898 180986 38134
rect 181222 37898 181404 38134
rect 180804 2454 181404 37898
rect 180804 2218 180986 2454
rect 181222 2218 181404 2454
rect 180804 2134 181404 2218
rect 180804 1898 180986 2134
rect 181222 1898 181404 2134
rect 180804 -346 181404 1898
rect 180804 -582 180986 -346
rect 181222 -582 181404 -346
rect 180804 -666 181404 -582
rect 180804 -902 180986 -666
rect 181222 -902 181404 -666
rect 180804 -1864 181404 -902
rect 184404 294054 185004 317000
rect 184404 293818 184586 294054
rect 184822 293818 185004 294054
rect 184404 293734 185004 293818
rect 184404 293498 184586 293734
rect 184822 293498 185004 293734
rect 184404 258054 185004 293498
rect 184404 257818 184586 258054
rect 184822 257818 185004 258054
rect 184404 257734 185004 257818
rect 184404 257498 184586 257734
rect 184822 257498 185004 257734
rect 184404 222054 185004 257498
rect 184404 221818 184586 222054
rect 184822 221818 185004 222054
rect 184404 221734 185004 221818
rect 184404 221498 184586 221734
rect 184822 221498 185004 221734
rect 184404 186054 185004 221498
rect 184404 185818 184586 186054
rect 184822 185818 185004 186054
rect 184404 185734 185004 185818
rect 184404 185498 184586 185734
rect 184822 185498 185004 185734
rect 184404 150054 185004 185498
rect 184404 149818 184586 150054
rect 184822 149818 185004 150054
rect 184404 149734 185004 149818
rect 184404 149498 184586 149734
rect 184822 149498 185004 149734
rect 184404 114054 185004 149498
rect 184404 113818 184586 114054
rect 184822 113818 185004 114054
rect 184404 113734 185004 113818
rect 184404 113498 184586 113734
rect 184822 113498 185004 113734
rect 184404 78054 185004 113498
rect 184404 77818 184586 78054
rect 184822 77818 185004 78054
rect 184404 77734 185004 77818
rect 184404 77498 184586 77734
rect 184822 77498 185004 77734
rect 184404 42054 185004 77498
rect 184404 41818 184586 42054
rect 184822 41818 185004 42054
rect 184404 41734 185004 41818
rect 184404 41498 184586 41734
rect 184822 41498 185004 41734
rect 184404 6054 185004 41498
rect 184404 5818 184586 6054
rect 184822 5818 185004 6054
rect 184404 5734 185004 5818
rect 184404 5498 184586 5734
rect 184822 5498 185004 5734
rect 184404 -2226 185004 5498
rect 184404 -2462 184586 -2226
rect 184822 -2462 185004 -2226
rect 184404 -2546 185004 -2462
rect 184404 -2782 184586 -2546
rect 184822 -2782 185004 -2546
rect 184404 -3744 185004 -2782
rect 188004 297654 188604 317000
rect 188004 297418 188186 297654
rect 188422 297418 188604 297654
rect 188004 297334 188604 297418
rect 188004 297098 188186 297334
rect 188422 297098 188604 297334
rect 188004 261654 188604 297098
rect 188004 261418 188186 261654
rect 188422 261418 188604 261654
rect 188004 261334 188604 261418
rect 188004 261098 188186 261334
rect 188422 261098 188604 261334
rect 188004 225654 188604 261098
rect 188004 225418 188186 225654
rect 188422 225418 188604 225654
rect 188004 225334 188604 225418
rect 188004 225098 188186 225334
rect 188422 225098 188604 225334
rect 188004 189654 188604 225098
rect 188004 189418 188186 189654
rect 188422 189418 188604 189654
rect 188004 189334 188604 189418
rect 188004 189098 188186 189334
rect 188422 189098 188604 189334
rect 188004 153654 188604 189098
rect 188004 153418 188186 153654
rect 188422 153418 188604 153654
rect 188004 153334 188604 153418
rect 188004 153098 188186 153334
rect 188422 153098 188604 153334
rect 188004 117654 188604 153098
rect 188004 117418 188186 117654
rect 188422 117418 188604 117654
rect 188004 117334 188604 117418
rect 188004 117098 188186 117334
rect 188422 117098 188604 117334
rect 188004 81654 188604 117098
rect 188004 81418 188186 81654
rect 188422 81418 188604 81654
rect 188004 81334 188604 81418
rect 188004 81098 188186 81334
rect 188422 81098 188604 81334
rect 188004 45654 188604 81098
rect 188004 45418 188186 45654
rect 188422 45418 188604 45654
rect 188004 45334 188604 45418
rect 188004 45098 188186 45334
rect 188422 45098 188604 45334
rect 188004 9654 188604 45098
rect 188004 9418 188186 9654
rect 188422 9418 188604 9654
rect 188004 9334 188604 9418
rect 188004 9098 188186 9334
rect 188422 9098 188604 9334
rect 188004 -4106 188604 9098
rect 188004 -4342 188186 -4106
rect 188422 -4342 188604 -4106
rect 188004 -4426 188604 -4342
rect 188004 -4662 188186 -4426
rect 188422 -4662 188604 -4426
rect 188004 -5624 188604 -4662
rect 191604 301254 192204 317000
rect 191604 301018 191786 301254
rect 192022 301018 192204 301254
rect 191604 300934 192204 301018
rect 191604 300698 191786 300934
rect 192022 300698 192204 300934
rect 191604 265254 192204 300698
rect 191604 265018 191786 265254
rect 192022 265018 192204 265254
rect 191604 264934 192204 265018
rect 191604 264698 191786 264934
rect 192022 264698 192204 264934
rect 191604 229254 192204 264698
rect 191604 229018 191786 229254
rect 192022 229018 192204 229254
rect 191604 228934 192204 229018
rect 191604 228698 191786 228934
rect 192022 228698 192204 228934
rect 191604 193254 192204 228698
rect 191604 193018 191786 193254
rect 192022 193018 192204 193254
rect 191604 192934 192204 193018
rect 191604 192698 191786 192934
rect 192022 192698 192204 192934
rect 191604 157254 192204 192698
rect 191604 157018 191786 157254
rect 192022 157018 192204 157254
rect 191604 156934 192204 157018
rect 191604 156698 191786 156934
rect 192022 156698 192204 156934
rect 191604 121254 192204 156698
rect 191604 121018 191786 121254
rect 192022 121018 192204 121254
rect 191604 120934 192204 121018
rect 191604 120698 191786 120934
rect 192022 120698 192204 120934
rect 191604 85254 192204 120698
rect 191604 85018 191786 85254
rect 192022 85018 192204 85254
rect 191604 84934 192204 85018
rect 191604 84698 191786 84934
rect 192022 84698 192204 84934
rect 191604 49254 192204 84698
rect 191604 49018 191786 49254
rect 192022 49018 192204 49254
rect 191604 48934 192204 49018
rect 191604 48698 191786 48934
rect 192022 48698 192204 48934
rect 191604 13254 192204 48698
rect 191604 13018 191786 13254
rect 192022 13018 192204 13254
rect 191604 12934 192204 13018
rect 191604 12698 191786 12934
rect 192022 12698 192204 12934
rect 173604 -7162 173786 -6926
rect 174022 -7162 174204 -6926
rect 173604 -7246 174204 -7162
rect 173604 -7482 173786 -7246
rect 174022 -7482 174204 -7246
rect 173604 -7504 174204 -7482
rect 191604 -5986 192204 12698
rect 198804 308454 199404 317000
rect 198804 308218 198986 308454
rect 199222 308218 199404 308454
rect 198804 308134 199404 308218
rect 198804 307898 198986 308134
rect 199222 307898 199404 308134
rect 198804 272454 199404 307898
rect 198804 272218 198986 272454
rect 199222 272218 199404 272454
rect 198804 272134 199404 272218
rect 198804 271898 198986 272134
rect 199222 271898 199404 272134
rect 198804 236454 199404 271898
rect 198804 236218 198986 236454
rect 199222 236218 199404 236454
rect 198804 236134 199404 236218
rect 198804 235898 198986 236134
rect 199222 235898 199404 236134
rect 198804 200454 199404 235898
rect 198804 200218 198986 200454
rect 199222 200218 199404 200454
rect 198804 200134 199404 200218
rect 198804 199898 198986 200134
rect 199222 199898 199404 200134
rect 198804 164454 199404 199898
rect 198804 164218 198986 164454
rect 199222 164218 199404 164454
rect 198804 164134 199404 164218
rect 198804 163898 198986 164134
rect 199222 163898 199404 164134
rect 198804 128454 199404 163898
rect 198804 128218 198986 128454
rect 199222 128218 199404 128454
rect 198804 128134 199404 128218
rect 198804 127898 198986 128134
rect 199222 127898 199404 128134
rect 198804 92454 199404 127898
rect 198804 92218 198986 92454
rect 199222 92218 199404 92454
rect 198804 92134 199404 92218
rect 198804 91898 198986 92134
rect 199222 91898 199404 92134
rect 198804 56454 199404 91898
rect 198804 56218 198986 56454
rect 199222 56218 199404 56454
rect 198804 56134 199404 56218
rect 198804 55898 198986 56134
rect 199222 55898 199404 56134
rect 198804 20454 199404 55898
rect 198804 20218 198986 20454
rect 199222 20218 199404 20454
rect 198804 20134 199404 20218
rect 198804 19898 198986 20134
rect 199222 19898 199404 20134
rect 198804 -1286 199404 19898
rect 198804 -1522 198986 -1286
rect 199222 -1522 199404 -1286
rect 198804 -1606 199404 -1522
rect 198804 -1842 198986 -1606
rect 199222 -1842 199404 -1606
rect 198804 -1864 199404 -1842
rect 202404 312054 203004 317000
rect 202404 311818 202586 312054
rect 202822 311818 203004 312054
rect 202404 311734 203004 311818
rect 202404 311498 202586 311734
rect 202822 311498 203004 311734
rect 202404 276054 203004 311498
rect 202404 275818 202586 276054
rect 202822 275818 203004 276054
rect 202404 275734 203004 275818
rect 202404 275498 202586 275734
rect 202822 275498 203004 275734
rect 202404 240054 203004 275498
rect 202404 239818 202586 240054
rect 202822 239818 203004 240054
rect 202404 239734 203004 239818
rect 202404 239498 202586 239734
rect 202822 239498 203004 239734
rect 202404 204054 203004 239498
rect 202404 203818 202586 204054
rect 202822 203818 203004 204054
rect 202404 203734 203004 203818
rect 202404 203498 202586 203734
rect 202822 203498 203004 203734
rect 202404 168054 203004 203498
rect 202404 167818 202586 168054
rect 202822 167818 203004 168054
rect 202404 167734 203004 167818
rect 202404 167498 202586 167734
rect 202822 167498 203004 167734
rect 202404 132054 203004 167498
rect 202404 131818 202586 132054
rect 202822 131818 203004 132054
rect 202404 131734 203004 131818
rect 202404 131498 202586 131734
rect 202822 131498 203004 131734
rect 202404 96054 203004 131498
rect 202404 95818 202586 96054
rect 202822 95818 203004 96054
rect 202404 95734 203004 95818
rect 202404 95498 202586 95734
rect 202822 95498 203004 95734
rect 202404 60054 203004 95498
rect 202404 59818 202586 60054
rect 202822 59818 203004 60054
rect 202404 59734 203004 59818
rect 202404 59498 202586 59734
rect 202822 59498 203004 59734
rect 202404 24054 203004 59498
rect 202404 23818 202586 24054
rect 202822 23818 203004 24054
rect 202404 23734 203004 23818
rect 202404 23498 202586 23734
rect 202822 23498 203004 23734
rect 202404 -3166 203004 23498
rect 202404 -3402 202586 -3166
rect 202822 -3402 203004 -3166
rect 202404 -3486 203004 -3402
rect 202404 -3722 202586 -3486
rect 202822 -3722 203004 -3486
rect 202404 -3744 203004 -3722
rect 206004 315654 206604 317000
rect 206004 315418 206186 315654
rect 206422 315418 206604 315654
rect 206004 315334 206604 315418
rect 206004 315098 206186 315334
rect 206422 315098 206604 315334
rect 206004 279654 206604 315098
rect 206004 279418 206186 279654
rect 206422 279418 206604 279654
rect 206004 279334 206604 279418
rect 206004 279098 206186 279334
rect 206422 279098 206604 279334
rect 206004 243654 206604 279098
rect 206004 243418 206186 243654
rect 206422 243418 206604 243654
rect 206004 243334 206604 243418
rect 206004 243098 206186 243334
rect 206422 243098 206604 243334
rect 206004 207654 206604 243098
rect 206004 207418 206186 207654
rect 206422 207418 206604 207654
rect 206004 207334 206604 207418
rect 206004 207098 206186 207334
rect 206422 207098 206604 207334
rect 206004 171654 206604 207098
rect 206004 171418 206186 171654
rect 206422 171418 206604 171654
rect 206004 171334 206604 171418
rect 206004 171098 206186 171334
rect 206422 171098 206604 171334
rect 206004 135654 206604 171098
rect 206004 135418 206186 135654
rect 206422 135418 206604 135654
rect 206004 135334 206604 135418
rect 206004 135098 206186 135334
rect 206422 135098 206604 135334
rect 206004 99654 206604 135098
rect 206004 99418 206186 99654
rect 206422 99418 206604 99654
rect 206004 99334 206604 99418
rect 206004 99098 206186 99334
rect 206422 99098 206604 99334
rect 206004 63654 206604 99098
rect 206004 63418 206186 63654
rect 206422 63418 206604 63654
rect 206004 63334 206604 63418
rect 206004 63098 206186 63334
rect 206422 63098 206604 63334
rect 206004 27654 206604 63098
rect 206004 27418 206186 27654
rect 206422 27418 206604 27654
rect 206004 27334 206604 27418
rect 206004 27098 206186 27334
rect 206422 27098 206604 27334
rect 206004 -5046 206604 27098
rect 206004 -5282 206186 -5046
rect 206422 -5282 206604 -5046
rect 206004 -5366 206604 -5282
rect 206004 -5602 206186 -5366
rect 206422 -5602 206604 -5366
rect 206004 -5624 206604 -5602
rect 209604 283254 210204 317000
rect 209604 283018 209786 283254
rect 210022 283018 210204 283254
rect 209604 282934 210204 283018
rect 209604 282698 209786 282934
rect 210022 282698 210204 282934
rect 209604 247254 210204 282698
rect 209604 247018 209786 247254
rect 210022 247018 210204 247254
rect 209604 246934 210204 247018
rect 209604 246698 209786 246934
rect 210022 246698 210204 246934
rect 209604 211254 210204 246698
rect 209604 211018 209786 211254
rect 210022 211018 210204 211254
rect 209604 210934 210204 211018
rect 209604 210698 209786 210934
rect 210022 210698 210204 210934
rect 209604 175254 210204 210698
rect 209604 175018 209786 175254
rect 210022 175018 210204 175254
rect 209604 174934 210204 175018
rect 209604 174698 209786 174934
rect 210022 174698 210204 174934
rect 209604 139254 210204 174698
rect 209604 139018 209786 139254
rect 210022 139018 210204 139254
rect 209604 138934 210204 139018
rect 209604 138698 209786 138934
rect 210022 138698 210204 138934
rect 209604 103254 210204 138698
rect 209604 103018 209786 103254
rect 210022 103018 210204 103254
rect 209604 102934 210204 103018
rect 209604 102698 209786 102934
rect 210022 102698 210204 102934
rect 209604 67254 210204 102698
rect 209604 67018 209786 67254
rect 210022 67018 210204 67254
rect 209604 66934 210204 67018
rect 209604 66698 209786 66934
rect 210022 66698 210204 66934
rect 209604 31254 210204 66698
rect 209604 31018 209786 31254
rect 210022 31018 210204 31254
rect 209604 30934 210204 31018
rect 209604 30698 209786 30934
rect 210022 30698 210204 30934
rect 191604 -6222 191786 -5986
rect 192022 -6222 192204 -5986
rect 191604 -6306 192204 -6222
rect 191604 -6542 191786 -6306
rect 192022 -6542 192204 -6306
rect 191604 -7504 192204 -6542
rect 209604 -6926 210204 30698
rect 216804 290454 217404 317000
rect 216804 290218 216986 290454
rect 217222 290218 217404 290454
rect 216804 290134 217404 290218
rect 216804 289898 216986 290134
rect 217222 289898 217404 290134
rect 216804 254454 217404 289898
rect 216804 254218 216986 254454
rect 217222 254218 217404 254454
rect 216804 254134 217404 254218
rect 216804 253898 216986 254134
rect 217222 253898 217404 254134
rect 216804 218454 217404 253898
rect 216804 218218 216986 218454
rect 217222 218218 217404 218454
rect 216804 218134 217404 218218
rect 216804 217898 216986 218134
rect 217222 217898 217404 218134
rect 216804 182454 217404 217898
rect 216804 182218 216986 182454
rect 217222 182218 217404 182454
rect 216804 182134 217404 182218
rect 216804 181898 216986 182134
rect 217222 181898 217404 182134
rect 216804 146454 217404 181898
rect 216804 146218 216986 146454
rect 217222 146218 217404 146454
rect 216804 146134 217404 146218
rect 216804 145898 216986 146134
rect 217222 145898 217404 146134
rect 216804 110454 217404 145898
rect 216804 110218 216986 110454
rect 217222 110218 217404 110454
rect 216804 110134 217404 110218
rect 216804 109898 216986 110134
rect 217222 109898 217404 110134
rect 216804 74454 217404 109898
rect 216804 74218 216986 74454
rect 217222 74218 217404 74454
rect 216804 74134 217404 74218
rect 216804 73898 216986 74134
rect 217222 73898 217404 74134
rect 216804 38454 217404 73898
rect 216804 38218 216986 38454
rect 217222 38218 217404 38454
rect 216804 38134 217404 38218
rect 216804 37898 216986 38134
rect 217222 37898 217404 38134
rect 216804 2454 217404 37898
rect 216804 2218 216986 2454
rect 217222 2218 217404 2454
rect 216804 2134 217404 2218
rect 216804 1898 216986 2134
rect 217222 1898 217404 2134
rect 216804 -346 217404 1898
rect 216804 -582 216986 -346
rect 217222 -582 217404 -346
rect 216804 -666 217404 -582
rect 216804 -902 216986 -666
rect 217222 -902 217404 -666
rect 216804 -1864 217404 -902
rect 220404 294054 221004 317000
rect 220404 293818 220586 294054
rect 220822 293818 221004 294054
rect 220404 293734 221004 293818
rect 220404 293498 220586 293734
rect 220822 293498 221004 293734
rect 220404 258054 221004 293498
rect 220404 257818 220586 258054
rect 220822 257818 221004 258054
rect 220404 257734 221004 257818
rect 220404 257498 220586 257734
rect 220822 257498 221004 257734
rect 220404 222054 221004 257498
rect 220404 221818 220586 222054
rect 220822 221818 221004 222054
rect 220404 221734 221004 221818
rect 220404 221498 220586 221734
rect 220822 221498 221004 221734
rect 220404 186054 221004 221498
rect 220404 185818 220586 186054
rect 220822 185818 221004 186054
rect 220404 185734 221004 185818
rect 220404 185498 220586 185734
rect 220822 185498 221004 185734
rect 220404 150054 221004 185498
rect 220404 149818 220586 150054
rect 220822 149818 221004 150054
rect 220404 149734 221004 149818
rect 220404 149498 220586 149734
rect 220822 149498 221004 149734
rect 220404 114054 221004 149498
rect 220404 113818 220586 114054
rect 220822 113818 221004 114054
rect 220404 113734 221004 113818
rect 220404 113498 220586 113734
rect 220822 113498 221004 113734
rect 220404 78054 221004 113498
rect 220404 77818 220586 78054
rect 220822 77818 221004 78054
rect 220404 77734 221004 77818
rect 220404 77498 220586 77734
rect 220822 77498 221004 77734
rect 220404 42054 221004 77498
rect 220404 41818 220586 42054
rect 220822 41818 221004 42054
rect 220404 41734 221004 41818
rect 220404 41498 220586 41734
rect 220822 41498 221004 41734
rect 220404 6054 221004 41498
rect 220404 5818 220586 6054
rect 220822 5818 221004 6054
rect 220404 5734 221004 5818
rect 220404 5498 220586 5734
rect 220822 5498 221004 5734
rect 220404 -2226 221004 5498
rect 220404 -2462 220586 -2226
rect 220822 -2462 221004 -2226
rect 220404 -2546 221004 -2462
rect 220404 -2782 220586 -2546
rect 220822 -2782 221004 -2546
rect 220404 -3744 221004 -2782
rect 224004 297654 224604 317000
rect 224004 297418 224186 297654
rect 224422 297418 224604 297654
rect 224004 297334 224604 297418
rect 224004 297098 224186 297334
rect 224422 297098 224604 297334
rect 224004 261654 224604 297098
rect 224004 261418 224186 261654
rect 224422 261418 224604 261654
rect 224004 261334 224604 261418
rect 224004 261098 224186 261334
rect 224422 261098 224604 261334
rect 224004 225654 224604 261098
rect 224004 225418 224186 225654
rect 224422 225418 224604 225654
rect 224004 225334 224604 225418
rect 224004 225098 224186 225334
rect 224422 225098 224604 225334
rect 224004 189654 224604 225098
rect 224004 189418 224186 189654
rect 224422 189418 224604 189654
rect 224004 189334 224604 189418
rect 224004 189098 224186 189334
rect 224422 189098 224604 189334
rect 224004 153654 224604 189098
rect 224004 153418 224186 153654
rect 224422 153418 224604 153654
rect 224004 153334 224604 153418
rect 224004 153098 224186 153334
rect 224422 153098 224604 153334
rect 224004 117654 224604 153098
rect 224004 117418 224186 117654
rect 224422 117418 224604 117654
rect 224004 117334 224604 117418
rect 224004 117098 224186 117334
rect 224422 117098 224604 117334
rect 224004 81654 224604 117098
rect 224004 81418 224186 81654
rect 224422 81418 224604 81654
rect 224004 81334 224604 81418
rect 224004 81098 224186 81334
rect 224422 81098 224604 81334
rect 224004 45654 224604 81098
rect 224004 45418 224186 45654
rect 224422 45418 224604 45654
rect 224004 45334 224604 45418
rect 224004 45098 224186 45334
rect 224422 45098 224604 45334
rect 224004 9654 224604 45098
rect 224004 9418 224186 9654
rect 224422 9418 224604 9654
rect 224004 9334 224604 9418
rect 224004 9098 224186 9334
rect 224422 9098 224604 9334
rect 224004 -4106 224604 9098
rect 224004 -4342 224186 -4106
rect 224422 -4342 224604 -4106
rect 224004 -4426 224604 -4342
rect 224004 -4662 224186 -4426
rect 224422 -4662 224604 -4426
rect 224004 -5624 224604 -4662
rect 227604 301254 228204 317000
rect 227604 301018 227786 301254
rect 228022 301018 228204 301254
rect 227604 300934 228204 301018
rect 227604 300698 227786 300934
rect 228022 300698 228204 300934
rect 227604 265254 228204 300698
rect 227604 265018 227786 265254
rect 228022 265018 228204 265254
rect 227604 264934 228204 265018
rect 227604 264698 227786 264934
rect 228022 264698 228204 264934
rect 227604 229254 228204 264698
rect 227604 229018 227786 229254
rect 228022 229018 228204 229254
rect 227604 228934 228204 229018
rect 227604 228698 227786 228934
rect 228022 228698 228204 228934
rect 227604 193254 228204 228698
rect 227604 193018 227786 193254
rect 228022 193018 228204 193254
rect 227604 192934 228204 193018
rect 227604 192698 227786 192934
rect 228022 192698 228204 192934
rect 227604 157254 228204 192698
rect 227604 157018 227786 157254
rect 228022 157018 228204 157254
rect 227604 156934 228204 157018
rect 227604 156698 227786 156934
rect 228022 156698 228204 156934
rect 227604 121254 228204 156698
rect 227604 121018 227786 121254
rect 228022 121018 228204 121254
rect 227604 120934 228204 121018
rect 227604 120698 227786 120934
rect 228022 120698 228204 120934
rect 227604 85254 228204 120698
rect 227604 85018 227786 85254
rect 228022 85018 228204 85254
rect 227604 84934 228204 85018
rect 227604 84698 227786 84934
rect 228022 84698 228204 84934
rect 227604 49254 228204 84698
rect 227604 49018 227786 49254
rect 228022 49018 228204 49254
rect 227604 48934 228204 49018
rect 227604 48698 227786 48934
rect 228022 48698 228204 48934
rect 227604 13254 228204 48698
rect 227604 13018 227786 13254
rect 228022 13018 228204 13254
rect 227604 12934 228204 13018
rect 227604 12698 227786 12934
rect 228022 12698 228204 12934
rect 209604 -7162 209786 -6926
rect 210022 -7162 210204 -6926
rect 209604 -7246 210204 -7162
rect 209604 -7482 209786 -7246
rect 210022 -7482 210204 -7246
rect 209604 -7504 210204 -7482
rect 227604 -5986 228204 12698
rect 234804 308454 235404 317000
rect 234804 308218 234986 308454
rect 235222 308218 235404 308454
rect 234804 308134 235404 308218
rect 234804 307898 234986 308134
rect 235222 307898 235404 308134
rect 234804 272454 235404 307898
rect 234804 272218 234986 272454
rect 235222 272218 235404 272454
rect 234804 272134 235404 272218
rect 234804 271898 234986 272134
rect 235222 271898 235404 272134
rect 234804 236454 235404 271898
rect 234804 236218 234986 236454
rect 235222 236218 235404 236454
rect 234804 236134 235404 236218
rect 234804 235898 234986 236134
rect 235222 235898 235404 236134
rect 234804 200454 235404 235898
rect 234804 200218 234986 200454
rect 235222 200218 235404 200454
rect 234804 200134 235404 200218
rect 234804 199898 234986 200134
rect 235222 199898 235404 200134
rect 234804 164454 235404 199898
rect 234804 164218 234986 164454
rect 235222 164218 235404 164454
rect 234804 164134 235404 164218
rect 234804 163898 234986 164134
rect 235222 163898 235404 164134
rect 234804 128454 235404 163898
rect 234804 128218 234986 128454
rect 235222 128218 235404 128454
rect 234804 128134 235404 128218
rect 234804 127898 234986 128134
rect 235222 127898 235404 128134
rect 234804 92454 235404 127898
rect 234804 92218 234986 92454
rect 235222 92218 235404 92454
rect 234804 92134 235404 92218
rect 234804 91898 234986 92134
rect 235222 91898 235404 92134
rect 234804 56454 235404 91898
rect 234804 56218 234986 56454
rect 235222 56218 235404 56454
rect 234804 56134 235404 56218
rect 234804 55898 234986 56134
rect 235222 55898 235404 56134
rect 234804 20454 235404 55898
rect 234804 20218 234986 20454
rect 235222 20218 235404 20454
rect 234804 20134 235404 20218
rect 234804 19898 234986 20134
rect 235222 19898 235404 20134
rect 234804 -1286 235404 19898
rect 234804 -1522 234986 -1286
rect 235222 -1522 235404 -1286
rect 234804 -1606 235404 -1522
rect 234804 -1842 234986 -1606
rect 235222 -1842 235404 -1606
rect 234804 -1864 235404 -1842
rect 238404 312054 239004 317000
rect 238404 311818 238586 312054
rect 238822 311818 239004 312054
rect 238404 311734 239004 311818
rect 238404 311498 238586 311734
rect 238822 311498 239004 311734
rect 238404 276054 239004 311498
rect 238404 275818 238586 276054
rect 238822 275818 239004 276054
rect 238404 275734 239004 275818
rect 238404 275498 238586 275734
rect 238822 275498 239004 275734
rect 238404 240054 239004 275498
rect 238404 239818 238586 240054
rect 238822 239818 239004 240054
rect 238404 239734 239004 239818
rect 238404 239498 238586 239734
rect 238822 239498 239004 239734
rect 238404 204054 239004 239498
rect 238404 203818 238586 204054
rect 238822 203818 239004 204054
rect 238404 203734 239004 203818
rect 238404 203498 238586 203734
rect 238822 203498 239004 203734
rect 238404 168054 239004 203498
rect 238404 167818 238586 168054
rect 238822 167818 239004 168054
rect 238404 167734 239004 167818
rect 238404 167498 238586 167734
rect 238822 167498 239004 167734
rect 238404 132054 239004 167498
rect 238404 131818 238586 132054
rect 238822 131818 239004 132054
rect 238404 131734 239004 131818
rect 238404 131498 238586 131734
rect 238822 131498 239004 131734
rect 238404 96054 239004 131498
rect 238404 95818 238586 96054
rect 238822 95818 239004 96054
rect 238404 95734 239004 95818
rect 238404 95498 238586 95734
rect 238822 95498 239004 95734
rect 238404 60054 239004 95498
rect 238404 59818 238586 60054
rect 238822 59818 239004 60054
rect 238404 59734 239004 59818
rect 238404 59498 238586 59734
rect 238822 59498 239004 59734
rect 238404 24054 239004 59498
rect 238404 23818 238586 24054
rect 238822 23818 239004 24054
rect 238404 23734 239004 23818
rect 238404 23498 238586 23734
rect 238822 23498 239004 23734
rect 238404 -3166 239004 23498
rect 238404 -3402 238586 -3166
rect 238822 -3402 239004 -3166
rect 238404 -3486 239004 -3402
rect 238404 -3722 238586 -3486
rect 238822 -3722 239004 -3486
rect 238404 -3744 239004 -3722
rect 242004 315654 242604 317000
rect 242004 315418 242186 315654
rect 242422 315418 242604 315654
rect 242004 315334 242604 315418
rect 242004 315098 242186 315334
rect 242422 315098 242604 315334
rect 242004 279654 242604 315098
rect 242004 279418 242186 279654
rect 242422 279418 242604 279654
rect 242004 279334 242604 279418
rect 242004 279098 242186 279334
rect 242422 279098 242604 279334
rect 242004 243654 242604 279098
rect 242004 243418 242186 243654
rect 242422 243418 242604 243654
rect 242004 243334 242604 243418
rect 242004 243098 242186 243334
rect 242422 243098 242604 243334
rect 242004 207654 242604 243098
rect 242004 207418 242186 207654
rect 242422 207418 242604 207654
rect 242004 207334 242604 207418
rect 242004 207098 242186 207334
rect 242422 207098 242604 207334
rect 242004 171654 242604 207098
rect 242004 171418 242186 171654
rect 242422 171418 242604 171654
rect 242004 171334 242604 171418
rect 242004 171098 242186 171334
rect 242422 171098 242604 171334
rect 242004 135654 242604 171098
rect 242004 135418 242186 135654
rect 242422 135418 242604 135654
rect 242004 135334 242604 135418
rect 242004 135098 242186 135334
rect 242422 135098 242604 135334
rect 242004 99654 242604 135098
rect 242004 99418 242186 99654
rect 242422 99418 242604 99654
rect 242004 99334 242604 99418
rect 242004 99098 242186 99334
rect 242422 99098 242604 99334
rect 242004 63654 242604 99098
rect 242004 63418 242186 63654
rect 242422 63418 242604 63654
rect 242004 63334 242604 63418
rect 242004 63098 242186 63334
rect 242422 63098 242604 63334
rect 242004 27654 242604 63098
rect 242004 27418 242186 27654
rect 242422 27418 242604 27654
rect 242004 27334 242604 27418
rect 242004 27098 242186 27334
rect 242422 27098 242604 27334
rect 242004 -5046 242604 27098
rect 242004 -5282 242186 -5046
rect 242422 -5282 242604 -5046
rect 242004 -5366 242604 -5282
rect 242004 -5602 242186 -5366
rect 242422 -5602 242604 -5366
rect 242004 -5624 242604 -5602
rect 245604 283254 246204 317000
rect 245604 283018 245786 283254
rect 246022 283018 246204 283254
rect 245604 282934 246204 283018
rect 245604 282698 245786 282934
rect 246022 282698 246204 282934
rect 245604 247254 246204 282698
rect 245604 247018 245786 247254
rect 246022 247018 246204 247254
rect 245604 246934 246204 247018
rect 245604 246698 245786 246934
rect 246022 246698 246204 246934
rect 245604 211254 246204 246698
rect 245604 211018 245786 211254
rect 246022 211018 246204 211254
rect 245604 210934 246204 211018
rect 245604 210698 245786 210934
rect 246022 210698 246204 210934
rect 245604 175254 246204 210698
rect 245604 175018 245786 175254
rect 246022 175018 246204 175254
rect 245604 174934 246204 175018
rect 245604 174698 245786 174934
rect 246022 174698 246204 174934
rect 245604 139254 246204 174698
rect 245604 139018 245786 139254
rect 246022 139018 246204 139254
rect 245604 138934 246204 139018
rect 245604 138698 245786 138934
rect 246022 138698 246204 138934
rect 245604 103254 246204 138698
rect 245604 103018 245786 103254
rect 246022 103018 246204 103254
rect 245604 102934 246204 103018
rect 245604 102698 245786 102934
rect 246022 102698 246204 102934
rect 245604 67254 246204 102698
rect 245604 67018 245786 67254
rect 246022 67018 246204 67254
rect 245604 66934 246204 67018
rect 245604 66698 245786 66934
rect 246022 66698 246204 66934
rect 245604 31254 246204 66698
rect 245604 31018 245786 31254
rect 246022 31018 246204 31254
rect 245604 30934 246204 31018
rect 245604 30698 245786 30934
rect 246022 30698 246204 30934
rect 227604 -6222 227786 -5986
rect 228022 -6222 228204 -5986
rect 227604 -6306 228204 -6222
rect 227604 -6542 227786 -6306
rect 228022 -6542 228204 -6306
rect 227604 -7504 228204 -6542
rect 245604 -6926 246204 30698
rect 252804 290454 253404 317000
rect 252804 290218 252986 290454
rect 253222 290218 253404 290454
rect 252804 290134 253404 290218
rect 252804 289898 252986 290134
rect 253222 289898 253404 290134
rect 252804 254454 253404 289898
rect 252804 254218 252986 254454
rect 253222 254218 253404 254454
rect 252804 254134 253404 254218
rect 252804 253898 252986 254134
rect 253222 253898 253404 254134
rect 252804 218454 253404 253898
rect 252804 218218 252986 218454
rect 253222 218218 253404 218454
rect 252804 218134 253404 218218
rect 252804 217898 252986 218134
rect 253222 217898 253404 218134
rect 252804 182454 253404 217898
rect 252804 182218 252986 182454
rect 253222 182218 253404 182454
rect 252804 182134 253404 182218
rect 252804 181898 252986 182134
rect 253222 181898 253404 182134
rect 252804 146454 253404 181898
rect 252804 146218 252986 146454
rect 253222 146218 253404 146454
rect 252804 146134 253404 146218
rect 252804 145898 252986 146134
rect 253222 145898 253404 146134
rect 252804 110454 253404 145898
rect 252804 110218 252986 110454
rect 253222 110218 253404 110454
rect 252804 110134 253404 110218
rect 252804 109898 252986 110134
rect 253222 109898 253404 110134
rect 252804 74454 253404 109898
rect 252804 74218 252986 74454
rect 253222 74218 253404 74454
rect 252804 74134 253404 74218
rect 252804 73898 252986 74134
rect 253222 73898 253404 74134
rect 252804 38454 253404 73898
rect 252804 38218 252986 38454
rect 253222 38218 253404 38454
rect 252804 38134 253404 38218
rect 252804 37898 252986 38134
rect 253222 37898 253404 38134
rect 252804 2454 253404 37898
rect 252804 2218 252986 2454
rect 253222 2218 253404 2454
rect 252804 2134 253404 2218
rect 252804 1898 252986 2134
rect 253222 1898 253404 2134
rect 252804 -346 253404 1898
rect 252804 -582 252986 -346
rect 253222 -582 253404 -346
rect 252804 -666 253404 -582
rect 252804 -902 252986 -666
rect 253222 -902 253404 -666
rect 252804 -1864 253404 -902
rect 256404 294054 257004 317000
rect 256404 293818 256586 294054
rect 256822 293818 257004 294054
rect 256404 293734 257004 293818
rect 256404 293498 256586 293734
rect 256822 293498 257004 293734
rect 256404 258054 257004 293498
rect 256404 257818 256586 258054
rect 256822 257818 257004 258054
rect 256404 257734 257004 257818
rect 256404 257498 256586 257734
rect 256822 257498 257004 257734
rect 256404 222054 257004 257498
rect 256404 221818 256586 222054
rect 256822 221818 257004 222054
rect 256404 221734 257004 221818
rect 256404 221498 256586 221734
rect 256822 221498 257004 221734
rect 256404 186054 257004 221498
rect 256404 185818 256586 186054
rect 256822 185818 257004 186054
rect 256404 185734 257004 185818
rect 256404 185498 256586 185734
rect 256822 185498 257004 185734
rect 256404 150054 257004 185498
rect 256404 149818 256586 150054
rect 256822 149818 257004 150054
rect 256404 149734 257004 149818
rect 256404 149498 256586 149734
rect 256822 149498 257004 149734
rect 256404 114054 257004 149498
rect 256404 113818 256586 114054
rect 256822 113818 257004 114054
rect 256404 113734 257004 113818
rect 256404 113498 256586 113734
rect 256822 113498 257004 113734
rect 256404 78054 257004 113498
rect 256404 77818 256586 78054
rect 256822 77818 257004 78054
rect 256404 77734 257004 77818
rect 256404 77498 256586 77734
rect 256822 77498 257004 77734
rect 256404 42054 257004 77498
rect 256404 41818 256586 42054
rect 256822 41818 257004 42054
rect 256404 41734 257004 41818
rect 256404 41498 256586 41734
rect 256822 41498 257004 41734
rect 256404 6054 257004 41498
rect 256404 5818 256586 6054
rect 256822 5818 257004 6054
rect 256404 5734 257004 5818
rect 256404 5498 256586 5734
rect 256822 5498 257004 5734
rect 256404 -2226 257004 5498
rect 256404 -2462 256586 -2226
rect 256822 -2462 257004 -2226
rect 256404 -2546 257004 -2462
rect 256404 -2782 256586 -2546
rect 256822 -2782 257004 -2546
rect 256404 -3744 257004 -2782
rect 260004 297654 260604 317000
rect 260004 297418 260186 297654
rect 260422 297418 260604 297654
rect 260004 297334 260604 297418
rect 260004 297098 260186 297334
rect 260422 297098 260604 297334
rect 260004 261654 260604 297098
rect 260004 261418 260186 261654
rect 260422 261418 260604 261654
rect 260004 261334 260604 261418
rect 260004 261098 260186 261334
rect 260422 261098 260604 261334
rect 260004 225654 260604 261098
rect 260004 225418 260186 225654
rect 260422 225418 260604 225654
rect 260004 225334 260604 225418
rect 260004 225098 260186 225334
rect 260422 225098 260604 225334
rect 260004 189654 260604 225098
rect 260004 189418 260186 189654
rect 260422 189418 260604 189654
rect 260004 189334 260604 189418
rect 260004 189098 260186 189334
rect 260422 189098 260604 189334
rect 260004 153654 260604 189098
rect 260004 153418 260186 153654
rect 260422 153418 260604 153654
rect 260004 153334 260604 153418
rect 260004 153098 260186 153334
rect 260422 153098 260604 153334
rect 260004 117654 260604 153098
rect 260004 117418 260186 117654
rect 260422 117418 260604 117654
rect 260004 117334 260604 117418
rect 260004 117098 260186 117334
rect 260422 117098 260604 117334
rect 260004 81654 260604 117098
rect 260004 81418 260186 81654
rect 260422 81418 260604 81654
rect 260004 81334 260604 81418
rect 260004 81098 260186 81334
rect 260422 81098 260604 81334
rect 260004 45654 260604 81098
rect 260004 45418 260186 45654
rect 260422 45418 260604 45654
rect 260004 45334 260604 45418
rect 260004 45098 260186 45334
rect 260422 45098 260604 45334
rect 260004 9654 260604 45098
rect 260004 9418 260186 9654
rect 260422 9418 260604 9654
rect 260004 9334 260604 9418
rect 260004 9098 260186 9334
rect 260422 9098 260604 9334
rect 260004 -4106 260604 9098
rect 260004 -4342 260186 -4106
rect 260422 -4342 260604 -4106
rect 260004 -4426 260604 -4342
rect 260004 -4662 260186 -4426
rect 260422 -4662 260604 -4426
rect 260004 -5624 260604 -4662
rect 263604 301254 264204 317000
rect 263604 301018 263786 301254
rect 264022 301018 264204 301254
rect 263604 300934 264204 301018
rect 263604 300698 263786 300934
rect 264022 300698 264204 300934
rect 263604 265254 264204 300698
rect 263604 265018 263786 265254
rect 264022 265018 264204 265254
rect 263604 264934 264204 265018
rect 263604 264698 263786 264934
rect 264022 264698 264204 264934
rect 263604 229254 264204 264698
rect 263604 229018 263786 229254
rect 264022 229018 264204 229254
rect 263604 228934 264204 229018
rect 263604 228698 263786 228934
rect 264022 228698 264204 228934
rect 263604 193254 264204 228698
rect 263604 193018 263786 193254
rect 264022 193018 264204 193254
rect 263604 192934 264204 193018
rect 263604 192698 263786 192934
rect 264022 192698 264204 192934
rect 263604 157254 264204 192698
rect 263604 157018 263786 157254
rect 264022 157018 264204 157254
rect 263604 156934 264204 157018
rect 263604 156698 263786 156934
rect 264022 156698 264204 156934
rect 263604 121254 264204 156698
rect 263604 121018 263786 121254
rect 264022 121018 264204 121254
rect 263604 120934 264204 121018
rect 263604 120698 263786 120934
rect 264022 120698 264204 120934
rect 263604 85254 264204 120698
rect 263604 85018 263786 85254
rect 264022 85018 264204 85254
rect 263604 84934 264204 85018
rect 263604 84698 263786 84934
rect 264022 84698 264204 84934
rect 263604 49254 264204 84698
rect 263604 49018 263786 49254
rect 264022 49018 264204 49254
rect 263604 48934 264204 49018
rect 263604 48698 263786 48934
rect 264022 48698 264204 48934
rect 263604 13254 264204 48698
rect 263604 13018 263786 13254
rect 264022 13018 264204 13254
rect 263604 12934 264204 13018
rect 263604 12698 263786 12934
rect 264022 12698 264204 12934
rect 245604 -7162 245786 -6926
rect 246022 -7162 246204 -6926
rect 245604 -7246 246204 -7162
rect 245604 -7482 245786 -7246
rect 246022 -7482 246204 -7246
rect 245604 -7504 246204 -7482
rect 263604 -5986 264204 12698
rect 270804 308454 271404 317000
rect 270804 308218 270986 308454
rect 271222 308218 271404 308454
rect 270804 308134 271404 308218
rect 270804 307898 270986 308134
rect 271222 307898 271404 308134
rect 270804 272454 271404 307898
rect 270804 272218 270986 272454
rect 271222 272218 271404 272454
rect 270804 272134 271404 272218
rect 270804 271898 270986 272134
rect 271222 271898 271404 272134
rect 270804 236454 271404 271898
rect 270804 236218 270986 236454
rect 271222 236218 271404 236454
rect 270804 236134 271404 236218
rect 270804 235898 270986 236134
rect 271222 235898 271404 236134
rect 270804 200454 271404 235898
rect 270804 200218 270986 200454
rect 271222 200218 271404 200454
rect 270804 200134 271404 200218
rect 270804 199898 270986 200134
rect 271222 199898 271404 200134
rect 270804 164454 271404 199898
rect 270804 164218 270986 164454
rect 271222 164218 271404 164454
rect 270804 164134 271404 164218
rect 270804 163898 270986 164134
rect 271222 163898 271404 164134
rect 270804 128454 271404 163898
rect 270804 128218 270986 128454
rect 271222 128218 271404 128454
rect 270804 128134 271404 128218
rect 270804 127898 270986 128134
rect 271222 127898 271404 128134
rect 270804 92454 271404 127898
rect 270804 92218 270986 92454
rect 271222 92218 271404 92454
rect 270804 92134 271404 92218
rect 270804 91898 270986 92134
rect 271222 91898 271404 92134
rect 270804 56454 271404 91898
rect 270804 56218 270986 56454
rect 271222 56218 271404 56454
rect 270804 56134 271404 56218
rect 270804 55898 270986 56134
rect 271222 55898 271404 56134
rect 270804 20454 271404 55898
rect 270804 20218 270986 20454
rect 271222 20218 271404 20454
rect 270804 20134 271404 20218
rect 270804 19898 270986 20134
rect 271222 19898 271404 20134
rect 270804 -1286 271404 19898
rect 270804 -1522 270986 -1286
rect 271222 -1522 271404 -1286
rect 270804 -1606 271404 -1522
rect 270804 -1842 270986 -1606
rect 271222 -1842 271404 -1606
rect 270804 -1864 271404 -1842
rect 274404 312054 275004 317000
rect 274404 311818 274586 312054
rect 274822 311818 275004 312054
rect 274404 311734 275004 311818
rect 274404 311498 274586 311734
rect 274822 311498 275004 311734
rect 274404 276054 275004 311498
rect 274404 275818 274586 276054
rect 274822 275818 275004 276054
rect 274404 275734 275004 275818
rect 274404 275498 274586 275734
rect 274822 275498 275004 275734
rect 274404 240054 275004 275498
rect 274404 239818 274586 240054
rect 274822 239818 275004 240054
rect 274404 239734 275004 239818
rect 274404 239498 274586 239734
rect 274822 239498 275004 239734
rect 274404 204054 275004 239498
rect 274404 203818 274586 204054
rect 274822 203818 275004 204054
rect 274404 203734 275004 203818
rect 274404 203498 274586 203734
rect 274822 203498 275004 203734
rect 274404 168054 275004 203498
rect 274404 167818 274586 168054
rect 274822 167818 275004 168054
rect 274404 167734 275004 167818
rect 274404 167498 274586 167734
rect 274822 167498 275004 167734
rect 274404 132054 275004 167498
rect 274404 131818 274586 132054
rect 274822 131818 275004 132054
rect 274404 131734 275004 131818
rect 274404 131498 274586 131734
rect 274822 131498 275004 131734
rect 274404 96054 275004 131498
rect 274404 95818 274586 96054
rect 274822 95818 275004 96054
rect 274404 95734 275004 95818
rect 274404 95498 274586 95734
rect 274822 95498 275004 95734
rect 274404 60054 275004 95498
rect 274404 59818 274586 60054
rect 274822 59818 275004 60054
rect 274404 59734 275004 59818
rect 274404 59498 274586 59734
rect 274822 59498 275004 59734
rect 274404 24054 275004 59498
rect 274404 23818 274586 24054
rect 274822 23818 275004 24054
rect 274404 23734 275004 23818
rect 274404 23498 274586 23734
rect 274822 23498 275004 23734
rect 274404 -3166 275004 23498
rect 274404 -3402 274586 -3166
rect 274822 -3402 275004 -3166
rect 274404 -3486 275004 -3402
rect 274404 -3722 274586 -3486
rect 274822 -3722 275004 -3486
rect 274404 -3744 275004 -3722
rect 278004 315654 278604 317000
rect 278004 315418 278186 315654
rect 278422 315418 278604 315654
rect 278004 315334 278604 315418
rect 278004 315098 278186 315334
rect 278422 315098 278604 315334
rect 278004 279654 278604 315098
rect 278004 279418 278186 279654
rect 278422 279418 278604 279654
rect 278004 279334 278604 279418
rect 278004 279098 278186 279334
rect 278422 279098 278604 279334
rect 278004 243654 278604 279098
rect 278004 243418 278186 243654
rect 278422 243418 278604 243654
rect 278004 243334 278604 243418
rect 278004 243098 278186 243334
rect 278422 243098 278604 243334
rect 278004 207654 278604 243098
rect 278004 207418 278186 207654
rect 278422 207418 278604 207654
rect 278004 207334 278604 207418
rect 278004 207098 278186 207334
rect 278422 207098 278604 207334
rect 278004 171654 278604 207098
rect 278004 171418 278186 171654
rect 278422 171418 278604 171654
rect 278004 171334 278604 171418
rect 278004 171098 278186 171334
rect 278422 171098 278604 171334
rect 278004 135654 278604 171098
rect 278004 135418 278186 135654
rect 278422 135418 278604 135654
rect 278004 135334 278604 135418
rect 278004 135098 278186 135334
rect 278422 135098 278604 135334
rect 278004 99654 278604 135098
rect 278004 99418 278186 99654
rect 278422 99418 278604 99654
rect 278004 99334 278604 99418
rect 278004 99098 278186 99334
rect 278422 99098 278604 99334
rect 278004 63654 278604 99098
rect 278004 63418 278186 63654
rect 278422 63418 278604 63654
rect 278004 63334 278604 63418
rect 278004 63098 278186 63334
rect 278422 63098 278604 63334
rect 278004 27654 278604 63098
rect 278004 27418 278186 27654
rect 278422 27418 278604 27654
rect 278004 27334 278604 27418
rect 278004 27098 278186 27334
rect 278422 27098 278604 27334
rect 278004 -5046 278604 27098
rect 278004 -5282 278186 -5046
rect 278422 -5282 278604 -5046
rect 278004 -5366 278604 -5282
rect 278004 -5602 278186 -5366
rect 278422 -5602 278604 -5366
rect 278004 -5624 278604 -5602
rect 281604 283254 282204 317000
rect 281604 283018 281786 283254
rect 282022 283018 282204 283254
rect 281604 282934 282204 283018
rect 281604 282698 281786 282934
rect 282022 282698 282204 282934
rect 281604 247254 282204 282698
rect 281604 247018 281786 247254
rect 282022 247018 282204 247254
rect 281604 246934 282204 247018
rect 281604 246698 281786 246934
rect 282022 246698 282204 246934
rect 281604 211254 282204 246698
rect 281604 211018 281786 211254
rect 282022 211018 282204 211254
rect 281604 210934 282204 211018
rect 281604 210698 281786 210934
rect 282022 210698 282204 210934
rect 281604 175254 282204 210698
rect 281604 175018 281786 175254
rect 282022 175018 282204 175254
rect 281604 174934 282204 175018
rect 281604 174698 281786 174934
rect 282022 174698 282204 174934
rect 281604 139254 282204 174698
rect 281604 139018 281786 139254
rect 282022 139018 282204 139254
rect 281604 138934 282204 139018
rect 281604 138698 281786 138934
rect 282022 138698 282204 138934
rect 281604 103254 282204 138698
rect 281604 103018 281786 103254
rect 282022 103018 282204 103254
rect 281604 102934 282204 103018
rect 281604 102698 281786 102934
rect 282022 102698 282204 102934
rect 281604 67254 282204 102698
rect 281604 67018 281786 67254
rect 282022 67018 282204 67254
rect 281604 66934 282204 67018
rect 281604 66698 281786 66934
rect 282022 66698 282204 66934
rect 281604 31254 282204 66698
rect 281604 31018 281786 31254
rect 282022 31018 282204 31254
rect 281604 30934 282204 31018
rect 281604 30698 281786 30934
rect 282022 30698 282204 30934
rect 263604 -6222 263786 -5986
rect 264022 -6222 264204 -5986
rect 263604 -6306 264204 -6222
rect 263604 -6542 263786 -6306
rect 264022 -6542 264204 -6306
rect 263604 -7504 264204 -6542
rect 281604 -6926 282204 30698
rect 288804 290454 289404 325898
rect 288804 290218 288986 290454
rect 289222 290218 289404 290454
rect 288804 290134 289404 290218
rect 288804 289898 288986 290134
rect 289222 289898 289404 290134
rect 288804 254454 289404 289898
rect 288804 254218 288986 254454
rect 289222 254218 289404 254454
rect 288804 254134 289404 254218
rect 288804 253898 288986 254134
rect 289222 253898 289404 254134
rect 288804 218454 289404 253898
rect 288804 218218 288986 218454
rect 289222 218218 289404 218454
rect 288804 218134 289404 218218
rect 288804 217898 288986 218134
rect 289222 217898 289404 218134
rect 288804 182454 289404 217898
rect 288804 182218 288986 182454
rect 289222 182218 289404 182454
rect 288804 182134 289404 182218
rect 288804 181898 288986 182134
rect 289222 181898 289404 182134
rect 288804 146454 289404 181898
rect 288804 146218 288986 146454
rect 289222 146218 289404 146454
rect 288804 146134 289404 146218
rect 288804 145898 288986 146134
rect 289222 145898 289404 146134
rect 288804 110454 289404 145898
rect 288804 110218 288986 110454
rect 289222 110218 289404 110454
rect 288804 110134 289404 110218
rect 288804 109898 288986 110134
rect 289222 109898 289404 110134
rect 288804 74454 289404 109898
rect 288804 74218 288986 74454
rect 289222 74218 289404 74454
rect 288804 74134 289404 74218
rect 288804 73898 288986 74134
rect 289222 73898 289404 74134
rect 288804 38454 289404 73898
rect 288804 38218 288986 38454
rect 289222 38218 289404 38454
rect 288804 38134 289404 38218
rect 288804 37898 288986 38134
rect 289222 37898 289404 38134
rect 288804 2454 289404 37898
rect 288804 2218 288986 2454
rect 289222 2218 289404 2454
rect 288804 2134 289404 2218
rect 288804 1898 288986 2134
rect 289222 1898 289404 2134
rect 288804 -346 289404 1898
rect 288804 -582 288986 -346
rect 289222 -582 289404 -346
rect 288804 -666 289404 -582
rect 288804 -902 288986 -666
rect 289222 -902 289404 -666
rect 288804 -1864 289404 -902
rect 292404 690054 293004 706162
rect 292404 689818 292586 690054
rect 292822 689818 293004 690054
rect 292404 689734 293004 689818
rect 292404 689498 292586 689734
rect 292822 689498 293004 689734
rect 292404 654054 293004 689498
rect 292404 653818 292586 654054
rect 292822 653818 293004 654054
rect 292404 653734 293004 653818
rect 292404 653498 292586 653734
rect 292822 653498 293004 653734
rect 292404 618054 293004 653498
rect 292404 617818 292586 618054
rect 292822 617818 293004 618054
rect 292404 617734 293004 617818
rect 292404 617498 292586 617734
rect 292822 617498 293004 617734
rect 292404 582054 293004 617498
rect 292404 581818 292586 582054
rect 292822 581818 293004 582054
rect 292404 581734 293004 581818
rect 292404 581498 292586 581734
rect 292822 581498 293004 581734
rect 292404 546054 293004 581498
rect 292404 545818 292586 546054
rect 292822 545818 293004 546054
rect 292404 545734 293004 545818
rect 292404 545498 292586 545734
rect 292822 545498 293004 545734
rect 292404 510054 293004 545498
rect 292404 509818 292586 510054
rect 292822 509818 293004 510054
rect 292404 509734 293004 509818
rect 292404 509498 292586 509734
rect 292822 509498 293004 509734
rect 292404 474054 293004 509498
rect 292404 473818 292586 474054
rect 292822 473818 293004 474054
rect 292404 473734 293004 473818
rect 292404 473498 292586 473734
rect 292822 473498 293004 473734
rect 292404 438054 293004 473498
rect 292404 437818 292586 438054
rect 292822 437818 293004 438054
rect 292404 437734 293004 437818
rect 292404 437498 292586 437734
rect 292822 437498 293004 437734
rect 292404 402054 293004 437498
rect 292404 401818 292586 402054
rect 292822 401818 293004 402054
rect 292404 401734 293004 401818
rect 292404 401498 292586 401734
rect 292822 401498 293004 401734
rect 292404 366054 293004 401498
rect 292404 365818 292586 366054
rect 292822 365818 293004 366054
rect 292404 365734 293004 365818
rect 292404 365498 292586 365734
rect 292822 365498 293004 365734
rect 292404 330054 293004 365498
rect 292404 329818 292586 330054
rect 292822 329818 293004 330054
rect 292404 329734 293004 329818
rect 292404 329498 292586 329734
rect 292822 329498 293004 329734
rect 292404 294054 293004 329498
rect 292404 293818 292586 294054
rect 292822 293818 293004 294054
rect 292404 293734 293004 293818
rect 292404 293498 292586 293734
rect 292822 293498 293004 293734
rect 292404 258054 293004 293498
rect 292404 257818 292586 258054
rect 292822 257818 293004 258054
rect 292404 257734 293004 257818
rect 292404 257498 292586 257734
rect 292822 257498 293004 257734
rect 292404 222054 293004 257498
rect 292404 221818 292586 222054
rect 292822 221818 293004 222054
rect 292404 221734 293004 221818
rect 292404 221498 292586 221734
rect 292822 221498 293004 221734
rect 292404 186054 293004 221498
rect 292404 185818 292586 186054
rect 292822 185818 293004 186054
rect 292404 185734 293004 185818
rect 292404 185498 292586 185734
rect 292822 185498 293004 185734
rect 292404 150054 293004 185498
rect 292404 149818 292586 150054
rect 292822 149818 293004 150054
rect 292404 149734 293004 149818
rect 292404 149498 292586 149734
rect 292822 149498 293004 149734
rect 292404 114054 293004 149498
rect 292404 113818 292586 114054
rect 292822 113818 293004 114054
rect 292404 113734 293004 113818
rect 292404 113498 292586 113734
rect 292822 113498 293004 113734
rect 292404 78054 293004 113498
rect 292404 77818 292586 78054
rect 292822 77818 293004 78054
rect 292404 77734 293004 77818
rect 292404 77498 292586 77734
rect 292822 77498 293004 77734
rect 292404 42054 293004 77498
rect 292404 41818 292586 42054
rect 292822 41818 293004 42054
rect 292404 41734 293004 41818
rect 292404 41498 292586 41734
rect 292822 41498 293004 41734
rect 292404 6054 293004 41498
rect 292404 5818 292586 6054
rect 292822 5818 293004 6054
rect 292404 5734 293004 5818
rect 292404 5498 292586 5734
rect 292822 5498 293004 5734
rect 292404 -2226 293004 5498
rect 292404 -2462 292586 -2226
rect 292822 -2462 293004 -2226
rect 292404 -2546 293004 -2462
rect 292404 -2782 292586 -2546
rect 292822 -2782 293004 -2546
rect 292404 -3744 293004 -2782
rect 296004 693654 296604 708042
rect 296004 693418 296186 693654
rect 296422 693418 296604 693654
rect 296004 693334 296604 693418
rect 296004 693098 296186 693334
rect 296422 693098 296604 693334
rect 296004 657654 296604 693098
rect 296004 657418 296186 657654
rect 296422 657418 296604 657654
rect 296004 657334 296604 657418
rect 296004 657098 296186 657334
rect 296422 657098 296604 657334
rect 296004 621654 296604 657098
rect 296004 621418 296186 621654
rect 296422 621418 296604 621654
rect 296004 621334 296604 621418
rect 296004 621098 296186 621334
rect 296422 621098 296604 621334
rect 296004 585654 296604 621098
rect 296004 585418 296186 585654
rect 296422 585418 296604 585654
rect 296004 585334 296604 585418
rect 296004 585098 296186 585334
rect 296422 585098 296604 585334
rect 296004 549654 296604 585098
rect 296004 549418 296186 549654
rect 296422 549418 296604 549654
rect 296004 549334 296604 549418
rect 296004 549098 296186 549334
rect 296422 549098 296604 549334
rect 296004 513654 296604 549098
rect 296004 513418 296186 513654
rect 296422 513418 296604 513654
rect 296004 513334 296604 513418
rect 296004 513098 296186 513334
rect 296422 513098 296604 513334
rect 296004 477654 296604 513098
rect 296004 477418 296186 477654
rect 296422 477418 296604 477654
rect 296004 477334 296604 477418
rect 296004 477098 296186 477334
rect 296422 477098 296604 477334
rect 296004 441654 296604 477098
rect 296004 441418 296186 441654
rect 296422 441418 296604 441654
rect 296004 441334 296604 441418
rect 296004 441098 296186 441334
rect 296422 441098 296604 441334
rect 296004 405654 296604 441098
rect 296004 405418 296186 405654
rect 296422 405418 296604 405654
rect 296004 405334 296604 405418
rect 296004 405098 296186 405334
rect 296422 405098 296604 405334
rect 296004 369654 296604 405098
rect 296004 369418 296186 369654
rect 296422 369418 296604 369654
rect 296004 369334 296604 369418
rect 296004 369098 296186 369334
rect 296422 369098 296604 369334
rect 296004 333654 296604 369098
rect 296004 333418 296186 333654
rect 296422 333418 296604 333654
rect 296004 333334 296604 333418
rect 296004 333098 296186 333334
rect 296422 333098 296604 333334
rect 296004 297654 296604 333098
rect 296004 297418 296186 297654
rect 296422 297418 296604 297654
rect 296004 297334 296604 297418
rect 296004 297098 296186 297334
rect 296422 297098 296604 297334
rect 296004 261654 296604 297098
rect 296004 261418 296186 261654
rect 296422 261418 296604 261654
rect 296004 261334 296604 261418
rect 296004 261098 296186 261334
rect 296422 261098 296604 261334
rect 296004 225654 296604 261098
rect 296004 225418 296186 225654
rect 296422 225418 296604 225654
rect 296004 225334 296604 225418
rect 296004 225098 296186 225334
rect 296422 225098 296604 225334
rect 296004 189654 296604 225098
rect 296004 189418 296186 189654
rect 296422 189418 296604 189654
rect 296004 189334 296604 189418
rect 296004 189098 296186 189334
rect 296422 189098 296604 189334
rect 296004 153654 296604 189098
rect 296004 153418 296186 153654
rect 296422 153418 296604 153654
rect 296004 153334 296604 153418
rect 296004 153098 296186 153334
rect 296422 153098 296604 153334
rect 296004 117654 296604 153098
rect 296004 117418 296186 117654
rect 296422 117418 296604 117654
rect 296004 117334 296604 117418
rect 296004 117098 296186 117334
rect 296422 117098 296604 117334
rect 296004 81654 296604 117098
rect 296004 81418 296186 81654
rect 296422 81418 296604 81654
rect 296004 81334 296604 81418
rect 296004 81098 296186 81334
rect 296422 81098 296604 81334
rect 296004 45654 296604 81098
rect 296004 45418 296186 45654
rect 296422 45418 296604 45654
rect 296004 45334 296604 45418
rect 296004 45098 296186 45334
rect 296422 45098 296604 45334
rect 296004 9654 296604 45098
rect 296004 9418 296186 9654
rect 296422 9418 296604 9654
rect 296004 9334 296604 9418
rect 296004 9098 296186 9334
rect 296422 9098 296604 9334
rect 296004 -4106 296604 9098
rect 296004 -4342 296186 -4106
rect 296422 -4342 296604 -4106
rect 296004 -4426 296604 -4342
rect 296004 -4662 296186 -4426
rect 296422 -4662 296604 -4426
rect 296004 -5624 296604 -4662
rect 299604 697254 300204 709922
rect 317604 711418 318204 711440
rect 317604 711182 317786 711418
rect 318022 711182 318204 711418
rect 317604 711098 318204 711182
rect 317604 710862 317786 711098
rect 318022 710862 318204 711098
rect 314004 709538 314604 709560
rect 314004 709302 314186 709538
rect 314422 709302 314604 709538
rect 314004 709218 314604 709302
rect 314004 708982 314186 709218
rect 314422 708982 314604 709218
rect 310404 707658 311004 707680
rect 310404 707422 310586 707658
rect 310822 707422 311004 707658
rect 310404 707338 311004 707422
rect 310404 707102 310586 707338
rect 310822 707102 311004 707338
rect 299604 697018 299786 697254
rect 300022 697018 300204 697254
rect 299604 696934 300204 697018
rect 299604 696698 299786 696934
rect 300022 696698 300204 696934
rect 299604 661254 300204 696698
rect 299604 661018 299786 661254
rect 300022 661018 300204 661254
rect 299604 660934 300204 661018
rect 299604 660698 299786 660934
rect 300022 660698 300204 660934
rect 299604 625254 300204 660698
rect 306804 705778 307404 705800
rect 306804 705542 306986 705778
rect 307222 705542 307404 705778
rect 306804 705458 307404 705542
rect 306804 705222 306986 705458
rect 307222 705222 307404 705458
rect 306804 668454 307404 705222
rect 306804 668218 306986 668454
rect 307222 668218 307404 668454
rect 306804 668134 307404 668218
rect 306804 667898 306986 668134
rect 307222 667898 307404 668134
rect 306804 654247 307404 667898
rect 310404 672054 311004 707102
rect 310404 671818 310586 672054
rect 310822 671818 311004 672054
rect 310404 671734 311004 671818
rect 310404 671498 310586 671734
rect 310822 671498 311004 671734
rect 310404 654247 311004 671498
rect 314004 675654 314604 708982
rect 314004 675418 314186 675654
rect 314422 675418 314604 675654
rect 314004 675334 314604 675418
rect 314004 675098 314186 675334
rect 314422 675098 314604 675334
rect 314004 654247 314604 675098
rect 317604 679254 318204 710862
rect 335604 710478 336204 711440
rect 335604 710242 335786 710478
rect 336022 710242 336204 710478
rect 335604 710158 336204 710242
rect 335604 709922 335786 710158
rect 336022 709922 336204 710158
rect 332004 708598 332604 709560
rect 332004 708362 332186 708598
rect 332422 708362 332604 708598
rect 332004 708278 332604 708362
rect 332004 708042 332186 708278
rect 332422 708042 332604 708278
rect 328404 706718 329004 707680
rect 328404 706482 328586 706718
rect 328822 706482 329004 706718
rect 328404 706398 329004 706482
rect 328404 706162 328586 706398
rect 328822 706162 329004 706398
rect 317604 679018 317786 679254
rect 318022 679018 318204 679254
rect 317604 678934 318204 679018
rect 317604 678698 317786 678934
rect 318022 678698 318204 678934
rect 317604 654247 318204 678698
rect 324804 704838 325404 705800
rect 324804 704602 324986 704838
rect 325222 704602 325404 704838
rect 324804 704518 325404 704602
rect 324804 704282 324986 704518
rect 325222 704282 325404 704518
rect 324804 686454 325404 704282
rect 324804 686218 324986 686454
rect 325222 686218 325404 686454
rect 324804 686134 325404 686218
rect 324804 685898 324986 686134
rect 325222 685898 325404 686134
rect 324804 654247 325404 685898
rect 328404 690054 329004 706162
rect 328404 689818 328586 690054
rect 328822 689818 329004 690054
rect 328404 689734 329004 689818
rect 328404 689498 328586 689734
rect 328822 689498 329004 689734
rect 328404 654247 329004 689498
rect 332004 693654 332604 708042
rect 332004 693418 332186 693654
rect 332422 693418 332604 693654
rect 332004 693334 332604 693418
rect 332004 693098 332186 693334
rect 332422 693098 332604 693334
rect 332004 657654 332604 693098
rect 332004 657418 332186 657654
rect 332422 657418 332604 657654
rect 332004 657334 332604 657418
rect 332004 657098 332186 657334
rect 332422 657098 332604 657334
rect 332004 654247 332604 657098
rect 335604 697254 336204 709922
rect 353604 711418 354204 711440
rect 353604 711182 353786 711418
rect 354022 711182 354204 711418
rect 353604 711098 354204 711182
rect 353604 710862 353786 711098
rect 354022 710862 354204 711098
rect 350004 709538 350604 709560
rect 350004 709302 350186 709538
rect 350422 709302 350604 709538
rect 350004 709218 350604 709302
rect 350004 708982 350186 709218
rect 350422 708982 350604 709218
rect 346404 707658 347004 707680
rect 346404 707422 346586 707658
rect 346822 707422 347004 707658
rect 346404 707338 347004 707422
rect 346404 707102 346586 707338
rect 346822 707102 347004 707338
rect 335604 697018 335786 697254
rect 336022 697018 336204 697254
rect 335604 696934 336204 697018
rect 335604 696698 335786 696934
rect 336022 696698 336204 696934
rect 335604 661254 336204 696698
rect 335604 661018 335786 661254
rect 336022 661018 336204 661254
rect 335604 660934 336204 661018
rect 335604 660698 335786 660934
rect 336022 660698 336204 660934
rect 335604 654247 336204 660698
rect 342804 705778 343404 705800
rect 342804 705542 342986 705778
rect 343222 705542 343404 705778
rect 342804 705458 343404 705542
rect 342804 705222 342986 705458
rect 343222 705222 343404 705458
rect 342804 668454 343404 705222
rect 342804 668218 342986 668454
rect 343222 668218 343404 668454
rect 342804 668134 343404 668218
rect 342804 667898 342986 668134
rect 343222 667898 343404 668134
rect 342804 654247 343404 667898
rect 346404 672054 347004 707102
rect 346404 671818 346586 672054
rect 346822 671818 347004 672054
rect 346404 671734 347004 671818
rect 346404 671498 346586 671734
rect 346822 671498 347004 671734
rect 346404 654247 347004 671498
rect 350004 675654 350604 708982
rect 350004 675418 350186 675654
rect 350422 675418 350604 675654
rect 350004 675334 350604 675418
rect 350004 675098 350186 675334
rect 350422 675098 350604 675334
rect 350004 654247 350604 675098
rect 353604 679254 354204 710862
rect 371604 710478 372204 711440
rect 371604 710242 371786 710478
rect 372022 710242 372204 710478
rect 371604 710158 372204 710242
rect 371604 709922 371786 710158
rect 372022 709922 372204 710158
rect 368004 708598 368604 709560
rect 368004 708362 368186 708598
rect 368422 708362 368604 708598
rect 368004 708278 368604 708362
rect 368004 708042 368186 708278
rect 368422 708042 368604 708278
rect 364404 706718 365004 707680
rect 364404 706482 364586 706718
rect 364822 706482 365004 706718
rect 364404 706398 365004 706482
rect 364404 706162 364586 706398
rect 364822 706162 365004 706398
rect 353604 679018 353786 679254
rect 354022 679018 354204 679254
rect 353604 678934 354204 679018
rect 353604 678698 353786 678934
rect 354022 678698 354204 678934
rect 353604 654247 354204 678698
rect 360804 704838 361404 705800
rect 360804 704602 360986 704838
rect 361222 704602 361404 704838
rect 360804 704518 361404 704602
rect 360804 704282 360986 704518
rect 361222 704282 361404 704518
rect 360804 686454 361404 704282
rect 360804 686218 360986 686454
rect 361222 686218 361404 686454
rect 360804 686134 361404 686218
rect 360804 685898 360986 686134
rect 361222 685898 361404 686134
rect 360804 654247 361404 685898
rect 364404 690054 365004 706162
rect 364404 689818 364586 690054
rect 364822 689818 365004 690054
rect 364404 689734 365004 689818
rect 364404 689498 364586 689734
rect 364822 689498 365004 689734
rect 364404 654247 365004 689498
rect 368004 693654 368604 708042
rect 368004 693418 368186 693654
rect 368422 693418 368604 693654
rect 368004 693334 368604 693418
rect 368004 693098 368186 693334
rect 368422 693098 368604 693334
rect 368004 657654 368604 693098
rect 368004 657418 368186 657654
rect 368422 657418 368604 657654
rect 368004 657334 368604 657418
rect 368004 657098 368186 657334
rect 368422 657098 368604 657334
rect 368004 654247 368604 657098
rect 371604 697254 372204 709922
rect 389604 711418 390204 711440
rect 389604 711182 389786 711418
rect 390022 711182 390204 711418
rect 389604 711098 390204 711182
rect 389604 710862 389786 711098
rect 390022 710862 390204 711098
rect 386004 709538 386604 709560
rect 386004 709302 386186 709538
rect 386422 709302 386604 709538
rect 386004 709218 386604 709302
rect 386004 708982 386186 709218
rect 386422 708982 386604 709218
rect 382404 707658 383004 707680
rect 382404 707422 382586 707658
rect 382822 707422 383004 707658
rect 382404 707338 383004 707422
rect 382404 707102 382586 707338
rect 382822 707102 383004 707338
rect 371604 697018 371786 697254
rect 372022 697018 372204 697254
rect 371604 696934 372204 697018
rect 371604 696698 371786 696934
rect 372022 696698 372204 696934
rect 371604 661254 372204 696698
rect 371604 661018 371786 661254
rect 372022 661018 372204 661254
rect 371604 660934 372204 661018
rect 371604 660698 371786 660934
rect 372022 660698 372204 660934
rect 371604 654247 372204 660698
rect 378804 705778 379404 705800
rect 378804 705542 378986 705778
rect 379222 705542 379404 705778
rect 378804 705458 379404 705542
rect 378804 705222 378986 705458
rect 379222 705222 379404 705458
rect 378804 668454 379404 705222
rect 378804 668218 378986 668454
rect 379222 668218 379404 668454
rect 378804 668134 379404 668218
rect 378804 667898 378986 668134
rect 379222 667898 379404 668134
rect 378804 654247 379404 667898
rect 382404 672054 383004 707102
rect 382404 671818 382586 672054
rect 382822 671818 383004 672054
rect 382404 671734 383004 671818
rect 382404 671498 382586 671734
rect 382822 671498 383004 671734
rect 382404 654247 383004 671498
rect 386004 675654 386604 708982
rect 386004 675418 386186 675654
rect 386422 675418 386604 675654
rect 386004 675334 386604 675418
rect 386004 675098 386186 675334
rect 386422 675098 386604 675334
rect 386004 654247 386604 675098
rect 389604 679254 390204 710862
rect 407604 710478 408204 711440
rect 407604 710242 407786 710478
rect 408022 710242 408204 710478
rect 407604 710158 408204 710242
rect 407604 709922 407786 710158
rect 408022 709922 408204 710158
rect 404004 708598 404604 709560
rect 404004 708362 404186 708598
rect 404422 708362 404604 708598
rect 404004 708278 404604 708362
rect 404004 708042 404186 708278
rect 404422 708042 404604 708278
rect 400404 706718 401004 707680
rect 400404 706482 400586 706718
rect 400822 706482 401004 706718
rect 400404 706398 401004 706482
rect 400404 706162 400586 706398
rect 400822 706162 401004 706398
rect 389604 679018 389786 679254
rect 390022 679018 390204 679254
rect 389604 678934 390204 679018
rect 389604 678698 389786 678934
rect 390022 678698 390204 678934
rect 389604 654247 390204 678698
rect 396804 704838 397404 705800
rect 396804 704602 396986 704838
rect 397222 704602 397404 704838
rect 396804 704518 397404 704602
rect 396804 704282 396986 704518
rect 397222 704282 397404 704518
rect 396804 686454 397404 704282
rect 396804 686218 396986 686454
rect 397222 686218 397404 686454
rect 396804 686134 397404 686218
rect 396804 685898 396986 686134
rect 397222 685898 397404 686134
rect 378179 652900 378245 652901
rect 378179 652836 378180 652900
rect 378244 652836 378245 652900
rect 378179 652835 378245 652836
rect 383515 652900 383581 652901
rect 383515 652836 383516 652900
rect 383580 652836 383581 652900
rect 383515 652835 383581 652836
rect 378182 651130 378242 652835
rect 383518 651130 383578 652835
rect 378182 651070 378608 651130
rect 383518 651070 383603 651130
rect 396804 650454 397404 685898
rect 396804 650218 396986 650454
rect 397222 650218 397404 650454
rect 396804 650134 397404 650218
rect 396804 649898 396986 650134
rect 397222 649898 397404 650134
rect 386938 643254 387262 643276
rect 386938 643018 386982 643254
rect 387218 643018 387262 643254
rect 386938 642934 387262 643018
rect 386938 642698 386982 642934
rect 387218 642698 387262 642934
rect 386938 642676 387262 642698
rect 386938 639654 387262 639676
rect 386938 639418 386982 639654
rect 387218 639418 387262 639654
rect 386938 639334 387262 639418
rect 386938 639098 386982 639334
rect 387218 639098 387262 639334
rect 386938 639076 387262 639098
rect 386938 636054 387262 636076
rect 386938 635818 386982 636054
rect 387218 635818 387262 636054
rect 386938 635734 387262 635818
rect 386938 635498 386982 635734
rect 387218 635498 387262 635734
rect 386938 635476 387262 635498
rect 386938 632454 387262 632476
rect 386938 632218 386982 632454
rect 387218 632218 387262 632454
rect 386938 632134 387262 632218
rect 386938 631898 386982 632134
rect 387218 631898 387262 632134
rect 386938 631876 387262 631898
rect 299604 625018 299786 625254
rect 300022 625018 300204 625254
rect 299604 624934 300204 625018
rect 299604 624698 299786 624934
rect 300022 624698 300204 624934
rect 299604 589254 300204 624698
rect 386494 625254 386814 625276
rect 386494 625018 386536 625254
rect 386772 625018 386814 625254
rect 386494 624934 386814 625018
rect 386494 624698 386536 624934
rect 386772 624698 386814 624934
rect 386494 624676 386814 624698
rect 386494 621654 386814 621676
rect 386494 621418 386536 621654
rect 386772 621418 386814 621654
rect 386494 621334 386814 621418
rect 386494 621098 386536 621334
rect 386772 621098 386814 621334
rect 386494 621076 386814 621098
rect 386494 618054 386814 618076
rect 386494 617818 386536 618054
rect 386772 617818 386814 618054
rect 386494 617734 386814 617818
rect 386494 617498 386536 617734
rect 386772 617498 386814 617734
rect 386494 617476 386814 617498
rect 386494 614454 386814 614476
rect 386494 614218 386536 614454
rect 386772 614218 386814 614454
rect 386494 614134 386814 614218
rect 386494 613898 386536 614134
rect 386772 613898 386814 614134
rect 386494 613876 386814 613898
rect 396804 614454 397404 649898
rect 396804 614218 396986 614454
rect 397222 614218 397404 614454
rect 396804 614134 397404 614218
rect 396804 613898 396986 614134
rect 397222 613898 397404 614134
rect 386938 607254 387262 607276
rect 386938 607018 386982 607254
rect 387218 607018 387262 607254
rect 386938 606934 387262 607018
rect 386938 606698 386982 606934
rect 387218 606698 387262 606934
rect 386938 606676 387262 606698
rect 386938 603654 387262 603676
rect 386938 603418 386982 603654
rect 387218 603418 387262 603654
rect 386938 603334 387262 603418
rect 386938 603098 386982 603334
rect 387218 603098 387262 603334
rect 386938 603076 387262 603098
rect 386938 600054 387262 600076
rect 386938 599818 386982 600054
rect 387218 599818 387262 600054
rect 386938 599734 387262 599818
rect 386938 599498 386982 599734
rect 387218 599498 387262 599734
rect 386938 599476 387262 599498
rect 386938 596454 387262 596476
rect 386938 596218 386982 596454
rect 387218 596218 387262 596454
rect 386938 596134 387262 596218
rect 386938 595898 386982 596134
rect 387218 595898 387262 596134
rect 386938 595876 387262 595898
rect 299604 589018 299786 589254
rect 300022 589018 300204 589254
rect 299604 588934 300204 589018
rect 299604 588698 299786 588934
rect 300022 588698 300204 588934
rect 299604 553254 300204 588698
rect 386494 589254 386814 589276
rect 386494 589018 386536 589254
rect 386772 589018 386814 589254
rect 386494 588934 386814 589018
rect 386494 588698 386536 588934
rect 386772 588698 386814 588934
rect 386494 588676 386814 588698
rect 386494 585654 386814 585676
rect 386494 585418 386536 585654
rect 386772 585418 386814 585654
rect 386494 585334 386814 585418
rect 386494 585098 386536 585334
rect 386772 585098 386814 585334
rect 386494 585076 386814 585098
rect 386494 582054 386814 582076
rect 386494 581818 386536 582054
rect 386772 581818 386814 582054
rect 386494 581734 386814 581818
rect 386494 581498 386536 581734
rect 386772 581498 386814 581734
rect 386494 581476 386814 581498
rect 389219 580956 389285 580957
rect 389219 580892 389220 580956
rect 389284 580892 389285 580956
rect 389219 580891 389285 580892
rect 389222 579818 389282 580891
rect 386494 578454 386814 578476
rect 386494 578218 386536 578454
rect 386772 578218 386814 578454
rect 386494 578134 386814 578218
rect 386494 577898 386536 578134
rect 386772 577898 386814 578134
rect 386494 577876 386814 577898
rect 396804 578454 397404 613898
rect 396804 578218 396986 578454
rect 397222 578218 397404 578454
rect 396804 578134 397404 578218
rect 396804 577898 396986 578134
rect 397222 577898 397404 578134
rect 386938 571254 387262 571276
rect 386938 571018 386982 571254
rect 387218 571018 387262 571254
rect 386938 570934 387262 571018
rect 386938 570698 386982 570934
rect 387218 570698 387262 570934
rect 386938 570676 387262 570698
rect 386938 567654 387262 567676
rect 386938 567418 386982 567654
rect 387218 567418 387262 567654
rect 386938 567334 387262 567418
rect 386938 567098 386982 567334
rect 387218 567098 387262 567334
rect 386938 567076 387262 567098
rect 386938 564054 387262 564076
rect 386938 563818 386982 564054
rect 387218 563818 387262 564054
rect 386938 563734 387262 563818
rect 386938 563498 386982 563734
rect 387218 563498 387262 563734
rect 386938 563476 387262 563498
rect 323534 560430 323840 560490
rect 325132 560430 325434 560490
rect 313782 558925 313842 560350
rect 316358 560290 316832 560350
rect 317462 560290 318000 560350
rect 318934 560290 319168 560350
rect 313779 558924 313845 558925
rect 313779 558860 313780 558924
rect 313844 558860 313845 558924
rect 313779 558859 313845 558860
rect 316358 557837 316418 560290
rect 317462 558925 317522 560290
rect 318934 558925 318994 560290
rect 320306 560010 320366 560320
rect 320222 559950 320366 560010
rect 320958 560290 321504 560350
rect 320222 558925 320282 559950
rect 317459 558924 317525 558925
rect 317459 558860 317460 558924
rect 317524 558860 317525 558924
rect 317459 558859 317525 558860
rect 318931 558924 318997 558925
rect 318931 558860 318932 558924
rect 318996 558860 318997 558924
rect 318931 558859 318997 558860
rect 320219 558924 320285 558925
rect 320219 558860 320220 558924
rect 320284 558860 320285 558924
rect 320219 558859 320285 558860
rect 320958 558789 321018 560290
rect 322614 558789 322674 560350
rect 322796 560290 322858 560350
rect 320955 558788 321021 558789
rect 320955 558724 320956 558788
rect 321020 558724 321021 558788
rect 320955 558723 321021 558724
rect 322611 558788 322677 558789
rect 322611 558724 322612 558788
rect 322676 558724 322677 558788
rect 322611 558723 322677 558724
rect 322798 558109 322858 560290
rect 323534 558653 323594 560430
rect 323964 560290 324146 560350
rect 323531 558652 323597 558653
rect 323531 558588 323532 558652
rect 323596 558588 323597 558652
rect 323531 558587 323597 558588
rect 324086 558109 324146 560290
rect 324822 560290 325008 560350
rect 324822 558653 324882 560290
rect 324819 558652 324885 558653
rect 324819 558588 324820 558652
rect 324884 558588 324885 558652
rect 324819 558587 324885 558588
rect 322795 558108 322861 558109
rect 322795 558044 322796 558108
rect 322860 558044 322861 558108
rect 322795 558043 322861 558044
rect 324083 558108 324149 558109
rect 324083 558044 324084 558108
rect 324148 558044 324149 558108
rect 324083 558043 324149 558044
rect 316355 557836 316421 557837
rect 316355 557772 316356 557836
rect 316420 557772 316421 557836
rect 316355 557771 316421 557772
rect 325374 557701 325434 560430
rect 327030 560430 327344 560490
rect 328636 560430 328930 560490
rect 326110 560290 326176 560350
rect 326110 558789 326170 560290
rect 326294 558925 326354 560350
rect 326291 558924 326357 558925
rect 326291 558860 326292 558924
rect 326356 558860 326357 558924
rect 326291 558859 326357 558860
rect 326107 558788 326173 558789
rect 326107 558724 326108 558788
rect 326172 558724 326173 558788
rect 326107 558723 326173 558724
rect 327030 558653 327090 560430
rect 327468 560290 327642 560350
rect 327582 558925 327642 560290
rect 328482 559330 328542 560320
rect 328482 559270 328562 559330
rect 327579 558924 327645 558925
rect 327579 558860 327580 558924
rect 327644 558860 327645 558924
rect 327579 558859 327645 558860
rect 328502 558653 328562 559270
rect 328870 558789 328930 560430
rect 330526 560430 330848 560490
rect 332140 560430 332426 560490
rect 329606 560290 329680 560350
rect 329606 558925 329666 560290
rect 329603 558924 329669 558925
rect 329603 558860 329604 558924
rect 329668 558860 329669 558924
rect 329603 558859 329669 558860
rect 328867 558788 328933 558789
rect 328867 558724 328868 558788
rect 328932 558724 328933 558788
rect 328867 558723 328933 558724
rect 327027 558652 327093 558653
rect 327027 558588 327028 558652
rect 327092 558588 327093 558652
rect 327027 558587 327093 558588
rect 328499 558652 328565 558653
rect 328499 558588 328500 558652
rect 328564 558588 328565 558652
rect 328499 558587 328565 558588
rect 329790 557973 329850 560350
rect 330526 558789 330586 560430
rect 330972 560290 331138 560350
rect 331078 558925 331138 560290
rect 331814 560290 332016 560350
rect 331814 558925 331874 560290
rect 331075 558924 331141 558925
rect 331075 558860 331076 558924
rect 331140 558860 331141 558924
rect 331075 558859 331141 558860
rect 331811 558924 331877 558925
rect 331811 558860 331812 558924
rect 331876 558860 331877 558924
rect 331811 558859 331877 558860
rect 330523 558788 330589 558789
rect 330523 558724 330524 558788
rect 330588 558724 330589 558788
rect 330523 558723 330589 558724
rect 329787 557972 329853 557973
rect 329787 557908 329788 557972
rect 329852 557908 329853 557972
rect 329787 557907 329853 557908
rect 332366 557837 332426 560430
rect 334022 560430 334352 560490
rect 335644 560430 335922 560490
rect 333102 560290 333184 560350
rect 333102 558789 333162 560290
rect 333286 558925 333346 560350
rect 333283 558924 333349 558925
rect 333283 558860 333284 558924
rect 333348 558860 333349 558924
rect 333283 558859 333349 558860
rect 334022 558789 334082 560430
rect 334476 560290 334634 560350
rect 334574 558925 334634 560290
rect 335490 560010 335550 560320
rect 335490 559950 335554 560010
rect 334571 558924 334637 558925
rect 334571 558860 334572 558924
rect 334636 558860 334637 558924
rect 334571 558859 334637 558860
rect 335494 558789 335554 559950
rect 335862 558925 335922 560430
rect 339910 560430 340192 560490
rect 341484 560430 341810 560490
rect 348492 560430 348802 560490
rect 351996 560430 352298 560490
rect 355500 560430 355794 560490
rect 359004 560430 359290 560490
rect 336598 560290 336688 560350
rect 335859 558924 335925 558925
rect 335859 558860 335860 558924
rect 335924 558860 335925 558924
rect 335859 558859 335925 558860
rect 336598 558789 336658 560290
rect 336782 558925 336842 560320
rect 337702 560290 337856 560350
rect 337702 558925 337762 560290
rect 337950 559330 338010 560320
rect 337886 559270 338010 559330
rect 336779 558924 336845 558925
rect 336779 558860 336780 558924
rect 336844 558860 336845 558924
rect 336779 558859 336845 558860
rect 337699 558924 337765 558925
rect 337699 558860 337700 558924
rect 337764 558860 337765 558924
rect 337699 558859 337765 558860
rect 337886 558789 337946 559270
rect 338990 558789 339050 560350
rect 339148 560290 339234 560350
rect 339174 558925 339234 560290
rect 339171 558924 339237 558925
rect 339171 558860 339172 558924
rect 339236 558860 339237 558924
rect 339171 558859 339237 558860
rect 339910 558789 339970 560430
rect 340316 560290 340522 560350
rect 340462 558925 340522 560290
rect 341198 560290 341360 560350
rect 340459 558924 340525 558925
rect 340459 558860 340460 558924
rect 340524 558860 340525 558924
rect 340459 558859 340525 558860
rect 341198 558789 341258 560290
rect 341750 558925 341810 560430
rect 341747 558924 341813 558925
rect 341747 558860 341748 558924
rect 341812 558860 341813 558924
rect 341747 558859 341813 558860
rect 342486 558789 342546 560350
rect 342652 560290 342730 560350
rect 342670 558925 342730 560290
rect 343666 560010 343726 560320
rect 343820 560290 344018 560350
rect 343590 559950 343726 560010
rect 342667 558924 342733 558925
rect 342667 558860 342668 558924
rect 342732 558860 342733 558924
rect 342667 558859 342733 558860
rect 343590 558789 343650 559950
rect 343958 558925 344018 560290
rect 344326 560290 344864 560350
rect 344326 558925 344386 560290
rect 344958 559330 345018 560320
rect 344878 559270 345018 559330
rect 343955 558924 344021 558925
rect 343955 558860 343956 558924
rect 344020 558860 344021 558924
rect 343955 558859 344021 558860
rect 344323 558924 344389 558925
rect 344323 558860 344324 558924
rect 344388 558860 344389 558924
rect 344323 558859 344389 558860
rect 333099 558788 333165 558789
rect 333099 558724 333100 558788
rect 333164 558724 333165 558788
rect 333099 558723 333165 558724
rect 334019 558788 334085 558789
rect 334019 558724 334020 558788
rect 334084 558724 334085 558788
rect 334019 558723 334085 558724
rect 335491 558788 335557 558789
rect 335491 558724 335492 558788
rect 335556 558724 335557 558788
rect 335491 558723 335557 558724
rect 336595 558788 336661 558789
rect 336595 558724 336596 558788
rect 336660 558724 336661 558788
rect 336595 558723 336661 558724
rect 337883 558788 337949 558789
rect 337883 558724 337884 558788
rect 337948 558724 337949 558788
rect 337883 558723 337949 558724
rect 338987 558788 339053 558789
rect 338987 558724 338988 558788
rect 339052 558724 339053 558788
rect 338987 558723 339053 558724
rect 339907 558788 339973 558789
rect 339907 558724 339908 558788
rect 339972 558724 339973 558788
rect 339907 558723 339973 558724
rect 341195 558788 341261 558789
rect 341195 558724 341196 558788
rect 341260 558724 341261 558788
rect 341195 558723 341261 558724
rect 342483 558788 342549 558789
rect 342483 558724 342484 558788
rect 342548 558724 342549 558788
rect 342483 558723 342549 558724
rect 343587 558788 343653 558789
rect 343587 558724 343588 558788
rect 343652 558724 343653 558788
rect 343587 558723 343653 558724
rect 332363 557836 332429 557837
rect 332363 557772 332364 557836
rect 332428 557772 332429 557836
rect 332363 557771 332429 557772
rect 344878 557701 344938 559270
rect 345982 558789 346042 560350
rect 346156 560290 346226 560350
rect 346166 558925 346226 560290
rect 346902 560290 347200 560350
rect 347324 560290 347514 560350
rect 346163 558924 346229 558925
rect 346163 558860 346164 558924
rect 346228 558860 346229 558924
rect 346163 558859 346229 558860
rect 346902 558789 346962 560290
rect 347454 558925 347514 560290
rect 348190 560290 348368 560350
rect 347451 558924 347517 558925
rect 347451 558860 347452 558924
rect 347516 558860 347517 558924
rect 347451 558859 347517 558860
rect 348190 558789 348250 560290
rect 348742 558925 348802 560430
rect 348739 558924 348805 558925
rect 348739 558860 348740 558924
rect 348804 558860 348805 558924
rect 348739 558859 348805 558860
rect 349478 558789 349538 560350
rect 349660 560290 349722 560350
rect 349662 558925 349722 560290
rect 350674 560010 350734 560320
rect 350828 560290 351010 560350
rect 350582 559950 350734 560010
rect 349659 558924 349725 558925
rect 349659 558860 349660 558924
rect 349724 558860 349725 558924
rect 349659 558859 349725 558860
rect 345979 558788 346045 558789
rect 345979 558724 345980 558788
rect 346044 558724 346045 558788
rect 345979 558723 346045 558724
rect 346899 558788 346965 558789
rect 346899 558724 346900 558788
rect 346964 558724 346965 558788
rect 346899 558723 346965 558724
rect 348187 558788 348253 558789
rect 348187 558724 348188 558788
rect 348252 558724 348253 558788
rect 348187 558723 348253 558724
rect 349475 558788 349541 558789
rect 349475 558724 349476 558788
rect 349540 558724 349541 558788
rect 349475 558723 349541 558724
rect 350582 558517 350642 559950
rect 350579 558516 350645 558517
rect 350579 558452 350580 558516
rect 350644 558452 350645 558516
rect 350579 558451 350645 558452
rect 325371 557700 325437 557701
rect 325371 557636 325372 557700
rect 325436 557636 325437 557700
rect 325371 557635 325437 557636
rect 344875 557700 344941 557701
rect 344875 557636 344876 557700
rect 344940 557636 344941 557700
rect 344875 557635 344941 557636
rect 350950 557565 351010 560290
rect 351842 559333 351902 560320
rect 351842 559332 351933 559333
rect 351842 559270 351868 559332
rect 351867 559268 351868 559270
rect 351932 559268 351933 559332
rect 351867 559267 351933 559268
rect 350947 557564 351013 557565
rect 350947 557500 350948 557564
rect 351012 557500 351013 557564
rect 350947 557499 351013 557500
rect 299604 553018 299786 553254
rect 300022 553018 300204 553254
rect 299604 552934 300204 553018
rect 299604 552698 299786 552934
rect 300022 552698 300204 552934
rect 299604 517254 300204 552698
rect 299604 517018 299786 517254
rect 300022 517018 300204 517254
rect 299604 516934 300204 517018
rect 299604 516698 299786 516934
rect 300022 516698 300204 516934
rect 299604 481254 300204 516698
rect 299604 481018 299786 481254
rect 300022 481018 300204 481254
rect 299604 480934 300204 481018
rect 299604 480698 299786 480934
rect 300022 480698 300204 480934
rect 299604 445254 300204 480698
rect 299604 445018 299786 445254
rect 300022 445018 300204 445254
rect 299604 444934 300204 445018
rect 299604 444698 299786 444934
rect 300022 444698 300204 444934
rect 299604 409254 300204 444698
rect 299604 409018 299786 409254
rect 300022 409018 300204 409254
rect 299604 408934 300204 409018
rect 299604 408698 299786 408934
rect 300022 408698 300204 408934
rect 299604 373254 300204 408698
rect 299604 373018 299786 373254
rect 300022 373018 300204 373254
rect 299604 372934 300204 373018
rect 299604 372698 299786 372934
rect 300022 372698 300204 372934
rect 299604 337254 300204 372698
rect 299604 337018 299786 337254
rect 300022 337018 300204 337254
rect 299604 336934 300204 337018
rect 299604 336698 299786 336934
rect 300022 336698 300204 336934
rect 299604 301254 300204 336698
rect 306804 524454 307404 557000
rect 306804 524218 306986 524454
rect 307222 524218 307404 524454
rect 306804 524134 307404 524218
rect 306804 523898 306986 524134
rect 307222 523898 307404 524134
rect 306804 488454 307404 523898
rect 306804 488218 306986 488454
rect 307222 488218 307404 488454
rect 306804 488134 307404 488218
rect 306804 487898 306986 488134
rect 307222 487898 307404 488134
rect 306804 452454 307404 487898
rect 306804 452218 306986 452454
rect 307222 452218 307404 452454
rect 306804 452134 307404 452218
rect 306804 451898 306986 452134
rect 307222 451898 307404 452134
rect 306804 416454 307404 451898
rect 306804 416218 306986 416454
rect 307222 416218 307404 416454
rect 306804 416134 307404 416218
rect 306804 415898 306986 416134
rect 307222 415898 307404 416134
rect 306804 380454 307404 415898
rect 306804 380218 306986 380454
rect 307222 380218 307404 380454
rect 306804 380134 307404 380218
rect 306804 379898 306986 380134
rect 307222 379898 307404 380134
rect 306804 344454 307404 379898
rect 306804 344218 306986 344454
rect 307222 344218 307404 344454
rect 306804 344134 307404 344218
rect 306804 343898 306986 344134
rect 307222 343898 307404 344134
rect 306804 308454 307404 343898
rect 306804 308218 306986 308454
rect 307222 308218 307404 308454
rect 306804 308134 307404 308218
rect 306804 307898 306986 308134
rect 307222 307898 307404 308134
rect 306804 303000 307404 307898
rect 310404 528054 311004 557000
rect 310404 527818 310586 528054
rect 310822 527818 311004 528054
rect 310404 527734 311004 527818
rect 310404 527498 310586 527734
rect 310822 527498 311004 527734
rect 310404 492054 311004 527498
rect 310404 491818 310586 492054
rect 310822 491818 311004 492054
rect 310404 491734 311004 491818
rect 310404 491498 310586 491734
rect 310822 491498 311004 491734
rect 310404 456054 311004 491498
rect 310404 455818 310586 456054
rect 310822 455818 311004 456054
rect 310404 455734 311004 455818
rect 310404 455498 310586 455734
rect 310822 455498 311004 455734
rect 310404 420054 311004 455498
rect 310404 419818 310586 420054
rect 310822 419818 311004 420054
rect 310404 419734 311004 419818
rect 310404 419498 310586 419734
rect 310822 419498 311004 419734
rect 310404 384054 311004 419498
rect 310404 383818 310586 384054
rect 310822 383818 311004 384054
rect 310404 383734 311004 383818
rect 310404 383498 310586 383734
rect 310822 383498 311004 383734
rect 310404 348054 311004 383498
rect 310404 347818 310586 348054
rect 310822 347818 311004 348054
rect 310404 347734 311004 347818
rect 310404 347498 310586 347734
rect 310822 347498 311004 347734
rect 310404 312054 311004 347498
rect 310404 311818 310586 312054
rect 310822 311818 311004 312054
rect 310404 311734 311004 311818
rect 310404 311498 310586 311734
rect 310822 311498 311004 311734
rect 310404 303000 311004 311498
rect 314004 531654 314604 557000
rect 314004 531418 314186 531654
rect 314422 531418 314604 531654
rect 314004 531334 314604 531418
rect 314004 531098 314186 531334
rect 314422 531098 314604 531334
rect 314004 495654 314604 531098
rect 314004 495418 314186 495654
rect 314422 495418 314604 495654
rect 314004 495334 314604 495418
rect 314004 495098 314186 495334
rect 314422 495098 314604 495334
rect 314004 459654 314604 495098
rect 314004 459418 314186 459654
rect 314422 459418 314604 459654
rect 314004 459334 314604 459418
rect 314004 459098 314186 459334
rect 314422 459098 314604 459334
rect 314004 423654 314604 459098
rect 314004 423418 314186 423654
rect 314422 423418 314604 423654
rect 314004 423334 314604 423418
rect 314004 423098 314186 423334
rect 314422 423098 314604 423334
rect 314004 387654 314604 423098
rect 314004 387418 314186 387654
rect 314422 387418 314604 387654
rect 314004 387334 314604 387418
rect 314004 387098 314186 387334
rect 314422 387098 314604 387334
rect 314004 351654 314604 387098
rect 314004 351418 314186 351654
rect 314422 351418 314604 351654
rect 314004 351334 314604 351418
rect 314004 351098 314186 351334
rect 314422 351098 314604 351334
rect 314004 315654 314604 351098
rect 314004 315418 314186 315654
rect 314422 315418 314604 315654
rect 314004 315334 314604 315418
rect 314004 315098 314186 315334
rect 314422 315098 314604 315334
rect 314004 303000 314604 315098
rect 317604 535254 318204 557000
rect 317604 535018 317786 535254
rect 318022 535018 318204 535254
rect 317604 534934 318204 535018
rect 317604 534698 317786 534934
rect 318022 534698 318204 534934
rect 317604 499254 318204 534698
rect 317604 499018 317786 499254
rect 318022 499018 318204 499254
rect 317604 498934 318204 499018
rect 317604 498698 317786 498934
rect 318022 498698 318204 498934
rect 317604 463254 318204 498698
rect 317604 463018 317786 463254
rect 318022 463018 318204 463254
rect 317604 462934 318204 463018
rect 317604 462698 317786 462934
rect 318022 462698 318204 462934
rect 317604 427254 318204 462698
rect 317604 427018 317786 427254
rect 318022 427018 318204 427254
rect 317604 426934 318204 427018
rect 317604 426698 317786 426934
rect 318022 426698 318204 426934
rect 317604 391254 318204 426698
rect 317604 391018 317786 391254
rect 318022 391018 318204 391254
rect 317604 390934 318204 391018
rect 317604 390698 317786 390934
rect 318022 390698 318204 390934
rect 317604 355254 318204 390698
rect 317604 355018 317786 355254
rect 318022 355018 318204 355254
rect 317604 354934 318204 355018
rect 317604 354698 317786 354934
rect 318022 354698 318204 354934
rect 317604 319254 318204 354698
rect 317604 319018 317786 319254
rect 318022 319018 318204 319254
rect 317604 318934 318204 319018
rect 317604 318698 317786 318934
rect 318022 318698 318204 318934
rect 317604 303000 318204 318698
rect 324804 542454 325404 557000
rect 324804 542218 324986 542454
rect 325222 542218 325404 542454
rect 324804 542134 325404 542218
rect 324804 541898 324986 542134
rect 325222 541898 325404 542134
rect 324804 506454 325404 541898
rect 324804 506218 324986 506454
rect 325222 506218 325404 506454
rect 324804 506134 325404 506218
rect 324804 505898 324986 506134
rect 325222 505898 325404 506134
rect 324804 470454 325404 505898
rect 324804 470218 324986 470454
rect 325222 470218 325404 470454
rect 324804 470134 325404 470218
rect 324804 469898 324986 470134
rect 325222 469898 325404 470134
rect 324804 434454 325404 469898
rect 324804 434218 324986 434454
rect 325222 434218 325404 434454
rect 324804 434134 325404 434218
rect 324804 433898 324986 434134
rect 325222 433898 325404 434134
rect 324804 398454 325404 433898
rect 324804 398218 324986 398454
rect 325222 398218 325404 398454
rect 324804 398134 325404 398218
rect 324804 397898 324986 398134
rect 325222 397898 325404 398134
rect 324804 362454 325404 397898
rect 324804 362218 324986 362454
rect 325222 362218 325404 362454
rect 324804 362134 325404 362218
rect 324804 361898 324986 362134
rect 325222 361898 325404 362134
rect 324804 326454 325404 361898
rect 324804 326218 324986 326454
rect 325222 326218 325404 326454
rect 324804 326134 325404 326218
rect 324804 325898 324986 326134
rect 325222 325898 325404 326134
rect 324804 303000 325404 325898
rect 328404 546054 329004 557000
rect 328404 545818 328586 546054
rect 328822 545818 329004 546054
rect 328404 545734 329004 545818
rect 328404 545498 328586 545734
rect 328822 545498 329004 545734
rect 328404 510054 329004 545498
rect 328404 509818 328586 510054
rect 328822 509818 329004 510054
rect 328404 509734 329004 509818
rect 328404 509498 328586 509734
rect 328822 509498 329004 509734
rect 328404 474054 329004 509498
rect 328404 473818 328586 474054
rect 328822 473818 329004 474054
rect 328404 473734 329004 473818
rect 328404 473498 328586 473734
rect 328822 473498 329004 473734
rect 328404 438054 329004 473498
rect 328404 437818 328586 438054
rect 328822 437818 329004 438054
rect 328404 437734 329004 437818
rect 328404 437498 328586 437734
rect 328822 437498 329004 437734
rect 328404 402054 329004 437498
rect 328404 401818 328586 402054
rect 328822 401818 329004 402054
rect 328404 401734 329004 401818
rect 328404 401498 328586 401734
rect 328822 401498 329004 401734
rect 328404 366054 329004 401498
rect 328404 365818 328586 366054
rect 328822 365818 329004 366054
rect 328404 365734 329004 365818
rect 328404 365498 328586 365734
rect 328822 365498 329004 365734
rect 328404 330054 329004 365498
rect 328404 329818 328586 330054
rect 328822 329818 329004 330054
rect 328404 329734 329004 329818
rect 328404 329498 328586 329734
rect 328822 329498 329004 329734
rect 328404 303000 329004 329498
rect 332004 549654 332604 557000
rect 332004 549418 332186 549654
rect 332422 549418 332604 549654
rect 332004 549334 332604 549418
rect 332004 549098 332186 549334
rect 332422 549098 332604 549334
rect 332004 513654 332604 549098
rect 332004 513418 332186 513654
rect 332422 513418 332604 513654
rect 332004 513334 332604 513418
rect 332004 513098 332186 513334
rect 332422 513098 332604 513334
rect 332004 477654 332604 513098
rect 332004 477418 332186 477654
rect 332422 477418 332604 477654
rect 332004 477334 332604 477418
rect 332004 477098 332186 477334
rect 332422 477098 332604 477334
rect 332004 441654 332604 477098
rect 332004 441418 332186 441654
rect 332422 441418 332604 441654
rect 332004 441334 332604 441418
rect 332004 441098 332186 441334
rect 332422 441098 332604 441334
rect 332004 405654 332604 441098
rect 332004 405418 332186 405654
rect 332422 405418 332604 405654
rect 332004 405334 332604 405418
rect 332004 405098 332186 405334
rect 332422 405098 332604 405334
rect 332004 369654 332604 405098
rect 332004 369418 332186 369654
rect 332422 369418 332604 369654
rect 332004 369334 332604 369418
rect 332004 369098 332186 369334
rect 332422 369098 332604 369334
rect 332004 333654 332604 369098
rect 332004 333418 332186 333654
rect 332422 333418 332604 333654
rect 332004 333334 332604 333418
rect 332004 333098 332186 333334
rect 332422 333098 332604 333334
rect 332004 303000 332604 333098
rect 335604 553254 336204 557000
rect 335604 553018 335786 553254
rect 336022 553018 336204 553254
rect 335604 552934 336204 553018
rect 335604 552698 335786 552934
rect 336022 552698 336204 552934
rect 335604 517254 336204 552698
rect 335604 517018 335786 517254
rect 336022 517018 336204 517254
rect 335604 516934 336204 517018
rect 335604 516698 335786 516934
rect 336022 516698 336204 516934
rect 335604 481254 336204 516698
rect 335604 481018 335786 481254
rect 336022 481018 336204 481254
rect 335604 480934 336204 481018
rect 335604 480698 335786 480934
rect 336022 480698 336204 480934
rect 335604 445254 336204 480698
rect 335604 445018 335786 445254
rect 336022 445018 336204 445254
rect 335604 444934 336204 445018
rect 335604 444698 335786 444934
rect 336022 444698 336204 444934
rect 335604 409254 336204 444698
rect 342804 524454 343404 557000
rect 342804 524218 342986 524454
rect 343222 524218 343404 524454
rect 342804 524134 343404 524218
rect 342804 523898 342986 524134
rect 343222 523898 343404 524134
rect 342804 488454 343404 523898
rect 342804 488218 342986 488454
rect 343222 488218 343404 488454
rect 342804 488134 343404 488218
rect 342804 487898 342986 488134
rect 343222 487898 343404 488134
rect 342804 452454 343404 487898
rect 342804 452218 342986 452454
rect 343222 452218 343404 452454
rect 342804 452134 343404 452218
rect 342804 451898 342986 452134
rect 343222 451898 343404 452134
rect 342804 416454 343404 451898
rect 342804 416218 342986 416454
rect 343222 416218 343404 416454
rect 342804 416134 343404 416218
rect 342804 415898 342986 416134
rect 343222 415898 343404 416134
rect 342804 414247 343404 415898
rect 346404 528054 347004 557000
rect 346404 527818 346586 528054
rect 346822 527818 347004 528054
rect 346404 527734 347004 527818
rect 346404 527498 346586 527734
rect 346822 527498 347004 527734
rect 346404 492054 347004 527498
rect 346404 491818 346586 492054
rect 346822 491818 347004 492054
rect 346404 491734 347004 491818
rect 346404 491498 346586 491734
rect 346822 491498 347004 491734
rect 346404 456054 347004 491498
rect 346404 455818 346586 456054
rect 346822 455818 347004 456054
rect 346404 455734 347004 455818
rect 346404 455498 346586 455734
rect 346822 455498 347004 455734
rect 346404 420054 347004 455498
rect 346404 419818 346586 420054
rect 346822 419818 347004 420054
rect 346404 419734 347004 419818
rect 346404 419498 346586 419734
rect 346822 419498 347004 419734
rect 346404 414247 347004 419498
rect 350004 531654 350604 557000
rect 352238 555525 352298 560430
rect 352422 560290 353040 560350
rect 352422 558925 352482 560290
rect 352419 558924 352485 558925
rect 352419 558860 352420 558924
rect 352484 558860 352485 558924
rect 352419 558859 352485 558860
rect 353158 557701 353218 560350
rect 353526 560290 354208 560350
rect 354332 560290 354506 560350
rect 353526 558789 353586 560290
rect 353523 558788 353589 558789
rect 353523 558724 353524 558788
rect 353588 558724 353589 558788
rect 353523 558723 353589 558724
rect 353155 557700 353221 557701
rect 353155 557636 353156 557700
rect 353220 557636 353221 557700
rect 353155 557635 353221 557636
rect 354446 557565 354506 560290
rect 354814 560290 355376 560350
rect 354814 558789 354874 560290
rect 354811 558788 354877 558789
rect 354811 558724 354812 558788
rect 354876 558724 354877 558788
rect 354811 558723 354877 558724
rect 355734 557565 355794 560430
rect 356102 560290 356544 560350
rect 356102 558925 356162 560290
rect 356099 558924 356165 558925
rect 356099 558860 356100 558924
rect 356164 558860 356165 558924
rect 356099 558859 356165 558860
rect 356654 557565 356714 560350
rect 357682 560010 357742 560320
rect 357836 560290 358002 560350
rect 357574 559950 357742 560010
rect 357574 558517 357634 559950
rect 357571 558516 357637 558517
rect 357571 558452 357572 558516
rect 357636 558452 357637 558516
rect 357571 558451 357637 558452
rect 357942 557565 358002 560290
rect 358850 559333 358910 560320
rect 358850 559332 358925 559333
rect 358850 559270 358860 559332
rect 358859 559268 358860 559270
rect 358924 559268 358925 559332
rect 358859 559267 358925 559268
rect 354443 557564 354509 557565
rect 354443 557500 354444 557564
rect 354508 557500 354509 557564
rect 354443 557499 354509 557500
rect 355731 557564 355797 557565
rect 355731 557500 355732 557564
rect 355796 557500 355797 557564
rect 355731 557499 355797 557500
rect 356651 557564 356717 557565
rect 356651 557500 356652 557564
rect 356716 557500 356717 557564
rect 356651 557499 356717 557500
rect 357939 557564 358005 557565
rect 357939 557500 357940 557564
rect 358004 557500 358005 557564
rect 357939 557499 358005 557500
rect 352235 555524 352301 555525
rect 352235 555460 352236 555524
rect 352300 555460 352301 555524
rect 352235 555459 352301 555460
rect 350004 531418 350186 531654
rect 350422 531418 350604 531654
rect 350004 531334 350604 531418
rect 350004 531098 350186 531334
rect 350422 531098 350604 531334
rect 350004 495654 350604 531098
rect 350004 495418 350186 495654
rect 350422 495418 350604 495654
rect 350004 495334 350604 495418
rect 350004 495098 350186 495334
rect 350422 495098 350604 495334
rect 350004 459654 350604 495098
rect 350004 459418 350186 459654
rect 350422 459418 350604 459654
rect 350004 459334 350604 459418
rect 350004 459098 350186 459334
rect 350422 459098 350604 459334
rect 350004 423654 350604 459098
rect 350004 423418 350186 423654
rect 350422 423418 350604 423654
rect 350004 423334 350604 423418
rect 350004 423098 350186 423334
rect 350422 423098 350604 423334
rect 350004 414247 350604 423098
rect 353604 535254 354204 557000
rect 359230 555525 359290 560430
rect 359227 555524 359293 555525
rect 359227 555460 359228 555524
rect 359292 555460 359293 555524
rect 359227 555459 359293 555460
rect 353604 535018 353786 535254
rect 354022 535018 354204 535254
rect 353604 534934 354204 535018
rect 353604 534698 353786 534934
rect 354022 534698 354204 534934
rect 353604 499254 354204 534698
rect 353604 499018 353786 499254
rect 354022 499018 354204 499254
rect 353604 498934 354204 499018
rect 353604 498698 353786 498934
rect 354022 498698 354204 498934
rect 353604 463254 354204 498698
rect 353604 463018 353786 463254
rect 354022 463018 354204 463254
rect 353604 462934 354204 463018
rect 353604 462698 353786 462934
rect 354022 462698 354204 462934
rect 353604 427254 354204 462698
rect 353604 427018 353786 427254
rect 354022 427018 354204 427254
rect 353604 426934 354204 427018
rect 353604 426698 353786 426934
rect 354022 426698 354204 426934
rect 353604 414247 354204 426698
rect 360804 542454 361404 557000
rect 360804 542218 360986 542454
rect 361222 542218 361404 542454
rect 360804 542134 361404 542218
rect 360804 541898 360986 542134
rect 361222 541898 361404 542134
rect 360804 506454 361404 541898
rect 360804 506218 360986 506454
rect 361222 506218 361404 506454
rect 360804 506134 361404 506218
rect 360804 505898 360986 506134
rect 361222 505898 361404 506134
rect 360804 470454 361404 505898
rect 360804 470218 360986 470454
rect 361222 470218 361404 470454
rect 360804 470134 361404 470218
rect 360804 469898 360986 470134
rect 361222 469898 361404 470134
rect 360804 434454 361404 469898
rect 360804 434218 360986 434454
rect 361222 434218 361404 434454
rect 360804 434134 361404 434218
rect 360804 433898 360986 434134
rect 361222 433898 361404 434134
rect 360804 414247 361404 433898
rect 364404 546054 365004 557000
rect 364404 545818 364586 546054
rect 364822 545818 365004 546054
rect 364404 545734 365004 545818
rect 364404 545498 364586 545734
rect 364822 545498 365004 545734
rect 364404 510054 365004 545498
rect 364404 509818 364586 510054
rect 364822 509818 365004 510054
rect 364404 509734 365004 509818
rect 364404 509498 364586 509734
rect 364822 509498 365004 509734
rect 364404 474054 365004 509498
rect 364404 473818 364586 474054
rect 364822 473818 365004 474054
rect 364404 473734 365004 473818
rect 364404 473498 364586 473734
rect 364822 473498 365004 473734
rect 364404 438054 365004 473498
rect 364404 437818 364586 438054
rect 364822 437818 365004 438054
rect 364404 437734 365004 437818
rect 364404 437498 364586 437734
rect 364822 437498 365004 437734
rect 364404 414247 365004 437498
rect 368004 549654 368604 557000
rect 368004 549418 368186 549654
rect 368422 549418 368604 549654
rect 368004 549334 368604 549418
rect 368004 549098 368186 549334
rect 368422 549098 368604 549334
rect 368004 513654 368604 549098
rect 368004 513418 368186 513654
rect 368422 513418 368604 513654
rect 368004 513334 368604 513418
rect 368004 513098 368186 513334
rect 368422 513098 368604 513334
rect 368004 477654 368604 513098
rect 368004 477418 368186 477654
rect 368422 477418 368604 477654
rect 368004 477334 368604 477418
rect 368004 477098 368186 477334
rect 368422 477098 368604 477334
rect 368004 441654 368604 477098
rect 368004 441418 368186 441654
rect 368422 441418 368604 441654
rect 368004 441334 368604 441418
rect 368004 441098 368186 441334
rect 368422 441098 368604 441334
rect 368004 414247 368604 441098
rect 371604 553254 372204 557000
rect 371604 553018 371786 553254
rect 372022 553018 372204 553254
rect 371604 552934 372204 553018
rect 371604 552698 371786 552934
rect 372022 552698 372204 552934
rect 371604 517254 372204 552698
rect 371604 517018 371786 517254
rect 372022 517018 372204 517254
rect 371604 516934 372204 517018
rect 371604 516698 371786 516934
rect 372022 516698 372204 516934
rect 371604 481254 372204 516698
rect 371604 481018 371786 481254
rect 372022 481018 372204 481254
rect 371604 480934 372204 481018
rect 371604 480698 371786 480934
rect 372022 480698 372204 480934
rect 371604 445254 372204 480698
rect 371604 445018 371786 445254
rect 372022 445018 372204 445254
rect 371604 444934 372204 445018
rect 371604 444698 371786 444934
rect 372022 444698 372204 444934
rect 371604 414247 372204 444698
rect 378804 524454 379404 557000
rect 378804 524218 378986 524454
rect 379222 524218 379404 524454
rect 378804 524134 379404 524218
rect 378804 523898 378986 524134
rect 379222 523898 379404 524134
rect 378804 488454 379404 523898
rect 378804 488218 378986 488454
rect 379222 488218 379404 488454
rect 378804 488134 379404 488218
rect 378804 487898 378986 488134
rect 379222 487898 379404 488134
rect 378804 452454 379404 487898
rect 378804 452218 378986 452454
rect 379222 452218 379404 452454
rect 378804 452134 379404 452218
rect 378804 451898 378986 452134
rect 379222 451898 379404 452134
rect 378804 416454 379404 451898
rect 378804 416218 378986 416454
rect 379222 416218 379404 416454
rect 378804 416134 379404 416218
rect 378804 415898 378986 416134
rect 379222 415898 379404 416134
rect 378804 414247 379404 415898
rect 382404 528054 383004 557000
rect 382404 527818 382586 528054
rect 382822 527818 383004 528054
rect 382404 527734 383004 527818
rect 382404 527498 382586 527734
rect 382822 527498 383004 527734
rect 382404 492054 383004 527498
rect 382404 491818 382586 492054
rect 382822 491818 383004 492054
rect 382404 491734 383004 491818
rect 382404 491498 382586 491734
rect 382822 491498 383004 491734
rect 382404 456054 383004 491498
rect 382404 455818 382586 456054
rect 382822 455818 383004 456054
rect 382404 455734 383004 455818
rect 382404 455498 382586 455734
rect 382822 455498 383004 455734
rect 382404 420054 383004 455498
rect 382404 419818 382586 420054
rect 382822 419818 383004 420054
rect 382404 419734 383004 419818
rect 382404 419498 382586 419734
rect 382822 419498 383004 419734
rect 382404 414247 383004 419498
rect 386004 531654 386604 557000
rect 386004 531418 386186 531654
rect 386422 531418 386604 531654
rect 386004 531334 386604 531418
rect 386004 531098 386186 531334
rect 386422 531098 386604 531334
rect 386004 495654 386604 531098
rect 386004 495418 386186 495654
rect 386422 495418 386604 495654
rect 386004 495334 386604 495418
rect 386004 495098 386186 495334
rect 386422 495098 386604 495334
rect 386004 459654 386604 495098
rect 386004 459418 386186 459654
rect 386422 459418 386604 459654
rect 386004 459334 386604 459418
rect 386004 459098 386186 459334
rect 386422 459098 386604 459334
rect 386004 423654 386604 459098
rect 386004 423418 386186 423654
rect 386422 423418 386604 423654
rect 386004 423334 386604 423418
rect 386004 423098 386186 423334
rect 386422 423098 386604 423334
rect 386004 414247 386604 423098
rect 389604 535254 390204 557000
rect 389604 535018 389786 535254
rect 390022 535018 390204 535254
rect 389604 534934 390204 535018
rect 389604 534698 389786 534934
rect 390022 534698 390204 534934
rect 389604 499254 390204 534698
rect 389604 499018 389786 499254
rect 390022 499018 390204 499254
rect 389604 498934 390204 499018
rect 389604 498698 389786 498934
rect 390022 498698 390204 498934
rect 389604 463254 390204 498698
rect 389604 463018 389786 463254
rect 390022 463018 390204 463254
rect 389604 462934 390204 463018
rect 389604 462698 389786 462934
rect 390022 462698 390204 462934
rect 389604 427254 390204 462698
rect 389604 427018 389786 427254
rect 390022 427018 390204 427254
rect 389604 426934 390204 427018
rect 389604 426698 389786 426934
rect 390022 426698 390204 426934
rect 389604 414247 390204 426698
rect 396804 542454 397404 577898
rect 396804 542218 396986 542454
rect 397222 542218 397404 542454
rect 396804 542134 397404 542218
rect 396804 541898 396986 542134
rect 397222 541898 397404 542134
rect 396804 506454 397404 541898
rect 396804 506218 396986 506454
rect 397222 506218 397404 506454
rect 396804 506134 397404 506218
rect 396804 505898 396986 506134
rect 397222 505898 397404 506134
rect 396804 470454 397404 505898
rect 396804 470218 396986 470454
rect 397222 470218 397404 470454
rect 396804 470134 397404 470218
rect 396804 469898 396986 470134
rect 397222 469898 397404 470134
rect 396804 434454 397404 469898
rect 396804 434218 396986 434454
rect 397222 434218 397404 434454
rect 396804 434134 397404 434218
rect 396804 433898 396986 434134
rect 397222 433898 397404 434134
rect 396804 414247 397404 433898
rect 400404 690054 401004 706162
rect 400404 689818 400586 690054
rect 400822 689818 401004 690054
rect 400404 689734 401004 689818
rect 400404 689498 400586 689734
rect 400822 689498 401004 689734
rect 400404 654054 401004 689498
rect 400404 653818 400586 654054
rect 400822 653818 401004 654054
rect 400404 653734 401004 653818
rect 400404 653498 400586 653734
rect 400822 653498 401004 653734
rect 400404 618054 401004 653498
rect 400404 617818 400586 618054
rect 400822 617818 401004 618054
rect 400404 617734 401004 617818
rect 400404 617498 400586 617734
rect 400822 617498 401004 617734
rect 400404 582054 401004 617498
rect 400404 581818 400586 582054
rect 400822 581818 401004 582054
rect 400404 581734 401004 581818
rect 400404 581498 400586 581734
rect 400822 581498 401004 581734
rect 400404 546054 401004 581498
rect 400404 545818 400586 546054
rect 400822 545818 401004 546054
rect 400404 545734 401004 545818
rect 400404 545498 400586 545734
rect 400822 545498 401004 545734
rect 400404 510054 401004 545498
rect 400404 509818 400586 510054
rect 400822 509818 401004 510054
rect 400404 509734 401004 509818
rect 400404 509498 400586 509734
rect 400822 509498 401004 509734
rect 400404 474054 401004 509498
rect 400404 473818 400586 474054
rect 400822 473818 401004 474054
rect 400404 473734 401004 473818
rect 400404 473498 400586 473734
rect 400822 473498 401004 473734
rect 400404 438054 401004 473498
rect 400404 437818 400586 438054
rect 400822 437818 401004 438054
rect 400404 437734 401004 437818
rect 400404 437498 400586 437734
rect 400822 437498 401004 437734
rect 400404 414247 401004 437498
rect 404004 693654 404604 708042
rect 404004 693418 404186 693654
rect 404422 693418 404604 693654
rect 404004 693334 404604 693418
rect 404004 693098 404186 693334
rect 404422 693098 404604 693334
rect 404004 657654 404604 693098
rect 404004 657418 404186 657654
rect 404422 657418 404604 657654
rect 404004 657334 404604 657418
rect 404004 657098 404186 657334
rect 404422 657098 404604 657334
rect 404004 621654 404604 657098
rect 404004 621418 404186 621654
rect 404422 621418 404604 621654
rect 404004 621334 404604 621418
rect 404004 621098 404186 621334
rect 404422 621098 404604 621334
rect 404004 585654 404604 621098
rect 404004 585418 404186 585654
rect 404422 585418 404604 585654
rect 404004 585334 404604 585418
rect 404004 585098 404186 585334
rect 404422 585098 404604 585334
rect 404004 549654 404604 585098
rect 404004 549418 404186 549654
rect 404422 549418 404604 549654
rect 404004 549334 404604 549418
rect 404004 549098 404186 549334
rect 404422 549098 404604 549334
rect 404004 513654 404604 549098
rect 404004 513418 404186 513654
rect 404422 513418 404604 513654
rect 404004 513334 404604 513418
rect 404004 513098 404186 513334
rect 404422 513098 404604 513334
rect 404004 477654 404604 513098
rect 404004 477418 404186 477654
rect 404422 477418 404604 477654
rect 404004 477334 404604 477418
rect 404004 477098 404186 477334
rect 404422 477098 404604 477334
rect 404004 441654 404604 477098
rect 404004 441418 404186 441654
rect 404422 441418 404604 441654
rect 404004 441334 404604 441418
rect 404004 441098 404186 441334
rect 404422 441098 404604 441334
rect 404004 414247 404604 441098
rect 407604 697254 408204 709922
rect 425604 711418 426204 711440
rect 425604 711182 425786 711418
rect 426022 711182 426204 711418
rect 425604 711098 426204 711182
rect 425604 710862 425786 711098
rect 426022 710862 426204 711098
rect 422004 709538 422604 709560
rect 422004 709302 422186 709538
rect 422422 709302 422604 709538
rect 422004 709218 422604 709302
rect 422004 708982 422186 709218
rect 422422 708982 422604 709218
rect 418404 707658 419004 707680
rect 418404 707422 418586 707658
rect 418822 707422 419004 707658
rect 418404 707338 419004 707422
rect 418404 707102 418586 707338
rect 418822 707102 419004 707338
rect 407604 697018 407786 697254
rect 408022 697018 408204 697254
rect 407604 696934 408204 697018
rect 407604 696698 407786 696934
rect 408022 696698 408204 696934
rect 407604 661254 408204 696698
rect 407604 661018 407786 661254
rect 408022 661018 408204 661254
rect 407604 660934 408204 661018
rect 407604 660698 407786 660934
rect 408022 660698 408204 660934
rect 407604 625254 408204 660698
rect 407604 625018 407786 625254
rect 408022 625018 408204 625254
rect 407604 624934 408204 625018
rect 407604 624698 407786 624934
rect 408022 624698 408204 624934
rect 407604 589254 408204 624698
rect 407604 589018 407786 589254
rect 408022 589018 408204 589254
rect 407604 588934 408204 589018
rect 407604 588698 407786 588934
rect 408022 588698 408204 588934
rect 407604 553254 408204 588698
rect 407604 553018 407786 553254
rect 408022 553018 408204 553254
rect 407604 552934 408204 553018
rect 407604 552698 407786 552934
rect 408022 552698 408204 552934
rect 407604 517254 408204 552698
rect 407604 517018 407786 517254
rect 408022 517018 408204 517254
rect 407604 516934 408204 517018
rect 407604 516698 407786 516934
rect 408022 516698 408204 516934
rect 407604 481254 408204 516698
rect 407604 481018 407786 481254
rect 408022 481018 408204 481254
rect 407604 480934 408204 481018
rect 407604 480698 407786 480934
rect 408022 480698 408204 480934
rect 407604 445254 408204 480698
rect 407604 445018 407786 445254
rect 408022 445018 408204 445254
rect 407604 444934 408204 445018
rect 407604 444698 407786 444934
rect 408022 444698 408204 444934
rect 407604 414247 408204 444698
rect 414804 705778 415404 705800
rect 414804 705542 414986 705778
rect 415222 705542 415404 705778
rect 414804 705458 415404 705542
rect 414804 705222 414986 705458
rect 415222 705222 415404 705458
rect 414804 668454 415404 705222
rect 414804 668218 414986 668454
rect 415222 668218 415404 668454
rect 414804 668134 415404 668218
rect 414804 667898 414986 668134
rect 415222 667898 415404 668134
rect 414804 632454 415404 667898
rect 414804 632218 414986 632454
rect 415222 632218 415404 632454
rect 414804 632134 415404 632218
rect 414804 631898 414986 632134
rect 415222 631898 415404 632134
rect 414804 596454 415404 631898
rect 414804 596218 414986 596454
rect 415222 596218 415404 596454
rect 414804 596134 415404 596218
rect 414804 595898 414986 596134
rect 415222 595898 415404 596134
rect 414804 560454 415404 595898
rect 414804 560218 414986 560454
rect 415222 560218 415404 560454
rect 414804 560134 415404 560218
rect 414804 559898 414986 560134
rect 415222 559898 415404 560134
rect 414804 524454 415404 559898
rect 414804 524218 414986 524454
rect 415222 524218 415404 524454
rect 414804 524134 415404 524218
rect 414804 523898 414986 524134
rect 415222 523898 415404 524134
rect 414804 488454 415404 523898
rect 414804 488218 414986 488454
rect 415222 488218 415404 488454
rect 414804 488134 415404 488218
rect 414804 487898 414986 488134
rect 415222 487898 415404 488134
rect 414804 452454 415404 487898
rect 414804 452218 414986 452454
rect 415222 452218 415404 452454
rect 414804 452134 415404 452218
rect 414804 451898 414986 452134
rect 415222 451898 415404 452134
rect 414804 416454 415404 451898
rect 414804 416218 414986 416454
rect 415222 416218 415404 416454
rect 414804 416134 415404 416218
rect 414804 415898 414986 416134
rect 415222 415898 415404 416134
rect 414804 414247 415404 415898
rect 418404 672054 419004 707102
rect 418404 671818 418586 672054
rect 418822 671818 419004 672054
rect 418404 671734 419004 671818
rect 418404 671498 418586 671734
rect 418822 671498 419004 671734
rect 418404 636054 419004 671498
rect 418404 635818 418586 636054
rect 418822 635818 419004 636054
rect 418404 635734 419004 635818
rect 418404 635498 418586 635734
rect 418822 635498 419004 635734
rect 418404 600054 419004 635498
rect 418404 599818 418586 600054
rect 418822 599818 419004 600054
rect 418404 599734 419004 599818
rect 418404 599498 418586 599734
rect 418822 599498 419004 599734
rect 418404 564054 419004 599498
rect 418404 563818 418586 564054
rect 418822 563818 419004 564054
rect 418404 563734 419004 563818
rect 418404 563498 418586 563734
rect 418822 563498 419004 563734
rect 418404 528054 419004 563498
rect 418404 527818 418586 528054
rect 418822 527818 419004 528054
rect 418404 527734 419004 527818
rect 418404 527498 418586 527734
rect 418822 527498 419004 527734
rect 418404 492054 419004 527498
rect 418404 491818 418586 492054
rect 418822 491818 419004 492054
rect 418404 491734 419004 491818
rect 418404 491498 418586 491734
rect 418822 491498 419004 491734
rect 418404 456054 419004 491498
rect 418404 455818 418586 456054
rect 418822 455818 419004 456054
rect 418404 455734 419004 455818
rect 418404 455498 418586 455734
rect 418822 455498 419004 455734
rect 418404 420054 419004 455498
rect 418404 419818 418586 420054
rect 418822 419818 419004 420054
rect 418404 419734 419004 419818
rect 418404 419498 418586 419734
rect 418822 419498 419004 419734
rect 418404 414247 419004 419498
rect 422004 675654 422604 708982
rect 422004 675418 422186 675654
rect 422422 675418 422604 675654
rect 422004 675334 422604 675418
rect 422004 675098 422186 675334
rect 422422 675098 422604 675334
rect 422004 639654 422604 675098
rect 422004 639418 422186 639654
rect 422422 639418 422604 639654
rect 422004 639334 422604 639418
rect 422004 639098 422186 639334
rect 422422 639098 422604 639334
rect 422004 603654 422604 639098
rect 422004 603418 422186 603654
rect 422422 603418 422604 603654
rect 422004 603334 422604 603418
rect 422004 603098 422186 603334
rect 422422 603098 422604 603334
rect 422004 567654 422604 603098
rect 422004 567418 422186 567654
rect 422422 567418 422604 567654
rect 422004 567334 422604 567418
rect 422004 567098 422186 567334
rect 422422 567098 422604 567334
rect 422004 531654 422604 567098
rect 422004 531418 422186 531654
rect 422422 531418 422604 531654
rect 422004 531334 422604 531418
rect 422004 531098 422186 531334
rect 422422 531098 422604 531334
rect 422004 495654 422604 531098
rect 422004 495418 422186 495654
rect 422422 495418 422604 495654
rect 422004 495334 422604 495418
rect 422004 495098 422186 495334
rect 422422 495098 422604 495334
rect 422004 459654 422604 495098
rect 422004 459418 422186 459654
rect 422422 459418 422604 459654
rect 422004 459334 422604 459418
rect 422004 459098 422186 459334
rect 422422 459098 422604 459334
rect 422004 423654 422604 459098
rect 422004 423418 422186 423654
rect 422422 423418 422604 423654
rect 422004 423334 422604 423418
rect 422004 423098 422186 423334
rect 422422 423098 422604 423334
rect 368243 413948 368309 413949
rect 368243 413884 368244 413948
rect 368308 413884 368309 413948
rect 368243 413883 368309 413884
rect 368979 413948 369045 413949
rect 368979 413884 368980 413948
rect 369044 413884 369045 413948
rect 368979 413883 369045 413884
rect 370267 413948 370333 413949
rect 370267 413884 370268 413948
rect 370332 413884 370333 413948
rect 370267 413883 370333 413884
rect 371923 413948 371989 413949
rect 371923 413884 371924 413948
rect 371988 413884 371989 413948
rect 371923 413883 371989 413884
rect 373027 413948 373093 413949
rect 373027 413884 373028 413948
rect 373092 413884 373093 413948
rect 373027 413883 373093 413884
rect 380203 413948 380269 413949
rect 380203 413884 380204 413948
rect 380268 413884 380269 413948
rect 380203 413883 380269 413884
rect 384619 413948 384685 413949
rect 384619 413884 384620 413948
rect 384684 413884 384685 413948
rect 384619 413883 384685 413884
rect 388299 413948 388365 413949
rect 388299 413884 388300 413948
rect 388364 413884 388365 413948
rect 388299 413883 388365 413884
rect 390691 413948 390757 413949
rect 390691 413884 390692 413948
rect 390756 413884 390757 413948
rect 390691 413883 390757 413884
rect 392899 413948 392965 413949
rect 392899 413884 392900 413948
rect 392964 413884 392965 413948
rect 392899 413883 392965 413884
rect 397867 413948 397933 413949
rect 397867 413884 397868 413948
rect 397932 413884 397933 413948
rect 397867 413883 397933 413884
rect 403019 413948 403085 413949
rect 403019 413884 403020 413948
rect 403084 413884 403085 413948
rect 403019 413883 403085 413884
rect 407803 413948 407869 413949
rect 407803 413884 407804 413948
rect 407868 413884 407869 413948
rect 407803 413883 407869 413884
rect 410563 413948 410629 413949
rect 410563 413884 410564 413948
rect 410628 413884 410629 413948
rect 410563 413883 410629 413884
rect 413875 413948 413941 413949
rect 413875 413884 413876 413948
rect 413940 413884 413941 413948
rect 413875 413883 413941 413884
rect 367691 412724 367757 412725
rect 367691 412660 367692 412724
rect 367756 412660 367757 412724
rect 367691 412659 367757 412660
rect 367694 411090 367754 412659
rect 368246 411770 368306 413883
rect 368246 411710 368446 411770
rect 367694 411030 368292 411090
rect 368386 411060 368446 411710
rect 368982 411090 369042 413883
rect 369531 413132 369597 413133
rect 369531 413068 369532 413132
rect 369596 413068 369597 413132
rect 369531 413067 369597 413068
rect 369534 411770 369594 413067
rect 369534 411710 369614 411770
rect 368982 411030 369460 411090
rect 369554 411060 369614 411710
rect 370270 411090 370330 413883
rect 370819 413132 370885 413133
rect 370819 413068 370820 413132
rect 370884 413068 370885 413132
rect 370819 413067 370885 413068
rect 370822 411770 370882 413067
rect 371371 412724 371437 412725
rect 371371 412660 371372 412724
rect 371436 412660 371437 412724
rect 371371 412659 371437 412660
rect 370722 411710 370882 411770
rect 370270 411030 370628 411090
rect 370722 411060 370782 411710
rect 371374 411090 371434 412659
rect 371926 411090 371986 413883
rect 372659 412724 372725 412725
rect 372659 412660 372660 412724
rect 372724 412660 372725 412724
rect 372659 412659 372725 412660
rect 371374 411030 371796 411090
rect 371920 411030 371986 411090
rect 372662 410750 372722 412659
rect 373030 411770 373090 413883
rect 374315 413268 374381 413269
rect 374315 413204 374316 413268
rect 374380 413204 374381 413268
rect 374315 413203 374381 413204
rect 375419 413268 375485 413269
rect 375419 413204 375420 413268
rect 375484 413204 375485 413268
rect 375419 413203 375485 413204
rect 375971 413268 376037 413269
rect 375971 413204 375972 413268
rect 376036 413204 376037 413268
rect 375971 413203 376037 413204
rect 377811 413268 377877 413269
rect 377811 413204 377812 413268
rect 377876 413204 377877 413268
rect 377811 413203 377877 413204
rect 378915 413268 378981 413269
rect 378915 413204 378916 413268
rect 378980 413204 378981 413268
rect 378915 413203 378981 413204
rect 373947 412860 374013 412861
rect 373947 412796 373948 412860
rect 374012 412796 374013 412860
rect 373947 412795 374013 412796
rect 373030 411710 373118 411770
rect 373058 411060 373118 411710
rect 373950 411090 374010 412795
rect 374318 411770 374378 413203
rect 374683 412724 374749 412725
rect 374683 412660 374684 412724
rect 374748 412660 374749 412724
rect 374683 412659 374749 412660
rect 374226 411710 374378 411770
rect 373950 411030 374132 411090
rect 374226 411060 374286 411710
rect 374686 411090 374746 412659
rect 374686 411030 375300 411090
rect 375422 411030 375482 413203
rect 375974 411090 376034 413203
rect 376523 413132 376589 413133
rect 376523 413068 376524 413132
rect 376588 413068 376589 413132
rect 376523 413067 376589 413068
rect 376526 411770 376586 413067
rect 377259 412860 377325 412861
rect 377259 412796 377260 412860
rect 377324 412796 377325 412860
rect 377259 412795 377325 412796
rect 376526 411710 376622 411770
rect 375974 411030 376468 411090
rect 376562 411060 376622 411710
rect 377262 411090 377322 412795
rect 377814 411770 377874 413203
rect 378179 412860 378245 412861
rect 378179 412796 378180 412860
rect 378244 412796 378245 412860
rect 378179 412795 378245 412796
rect 377730 411710 377874 411770
rect 377262 411030 377636 411090
rect 377730 411060 377790 411710
rect 378182 411090 378242 412795
rect 378182 411030 378804 411090
rect 378918 411030 378978 413203
rect 379651 412860 379717 412861
rect 379651 412796 379652 412860
rect 379716 412796 379717 412860
rect 379651 412795 379717 412796
rect 379654 410750 379714 412795
rect 380206 411090 380266 413883
rect 381491 413404 381557 413405
rect 381491 413340 381492 413404
rect 381556 413340 381557 413404
rect 381491 413339 381557 413340
rect 382411 413404 382477 413405
rect 382411 413340 382412 413404
rect 382476 413340 382477 413404
rect 382411 413339 382477 413340
rect 380939 412724 381005 412725
rect 380939 412660 380940 412724
rect 381004 412660 381005 412724
rect 380939 412659 381005 412660
rect 380096 411030 380266 411090
rect 380942 411090 381002 412659
rect 380942 411030 381140 411090
rect 381494 410750 381554 413339
rect 382227 413132 382293 413133
rect 382227 413068 382228 413132
rect 382292 413068 382293 413132
rect 382227 413067 382293 413068
rect 382230 411090 382290 413067
rect 382230 411030 382308 411090
rect 382414 411030 382474 413339
rect 382779 413132 382845 413133
rect 382779 413068 382780 413132
rect 382844 413068 382845 413132
rect 382779 413067 382845 413068
rect 382782 411090 382842 413067
rect 383515 412724 383581 412725
rect 383515 412660 383516 412724
rect 383580 412660 383581 412724
rect 383515 412659 383581 412660
rect 384067 412724 384133 412725
rect 384067 412660 384068 412724
rect 384132 412660 384133 412724
rect 384067 412659 384133 412660
rect 383518 411770 383578 412659
rect 383518 411710 383630 411770
rect 382782 411030 383476 411090
rect 383570 411060 383630 411710
rect 384070 411090 384130 412659
rect 384622 411770 384682 413883
rect 386459 413540 386525 413541
rect 386459 413476 386460 413540
rect 386524 413476 386525 413540
rect 386459 413475 386525 413476
rect 385171 413132 385237 413133
rect 385171 413068 385172 413132
rect 385236 413068 385237 413132
rect 385171 413067 385237 413068
rect 384622 411710 384798 411770
rect 384070 411030 384644 411090
rect 384738 411060 384798 411710
rect 385174 411090 385234 413067
rect 385907 412724 385973 412725
rect 385907 412660 385908 412724
rect 385972 412660 385973 412724
rect 385907 412659 385973 412660
rect 385174 411030 385812 411090
rect 385910 411030 385970 412659
rect 386462 411090 386522 413475
rect 387195 413268 387261 413269
rect 387195 413204 387196 413268
rect 387260 413204 387261 413268
rect 387195 413203 387261 413204
rect 387198 411090 387258 413203
rect 388115 412724 388181 412725
rect 388115 412660 388116 412724
rect 388180 412660 388181 412724
rect 388115 412659 388181 412660
rect 386462 411030 386980 411090
rect 387104 411030 387258 411090
rect 388118 411060 388178 412659
rect 388302 411090 388362 413883
rect 389403 413676 389469 413677
rect 389403 413612 389404 413676
rect 389468 413612 389469 413676
rect 389403 413611 389469 413612
rect 389219 413540 389285 413541
rect 389219 413476 389220 413540
rect 389284 413476 389285 413540
rect 389219 413475 389285 413476
rect 389222 411770 389282 413475
rect 389406 411770 389466 413611
rect 389771 412996 389837 412997
rect 389771 412932 389772 412996
rect 389836 412932 389837 412996
rect 389771 412931 389837 412932
rect 389222 411710 389346 411770
rect 389406 411710 389470 411770
rect 388272 411030 388362 411090
rect 389286 411060 389346 411710
rect 389410 411060 389470 411710
rect 389774 411090 389834 412931
rect 390694 411770 390754 413883
rect 392163 413812 392229 413813
rect 392163 413748 392164 413812
rect 392228 413748 392229 413812
rect 392163 413747 392229 413748
rect 391795 413132 391861 413133
rect 391795 413068 391796 413132
rect 391860 413068 391861 413132
rect 391795 413067 391861 413068
rect 391059 412996 391125 412997
rect 391059 412932 391060 412996
rect 391124 412932 391125 412996
rect 391059 412931 391125 412932
rect 390578 411710 390754 411770
rect 389774 411030 390484 411090
rect 390578 411060 390638 411710
rect 391062 411090 391122 412931
rect 391798 411090 391858 413067
rect 391062 411030 391652 411090
rect 391776 411030 391858 411090
rect 392166 411090 392226 413747
rect 392902 411770 392962 413883
rect 396027 413812 396093 413813
rect 396027 413748 396028 413812
rect 396092 413748 396093 413812
rect 396027 413747 396093 413748
rect 394739 413540 394805 413541
rect 394739 413476 394740 413540
rect 394804 413476 394805 413540
rect 394739 413475 394805 413476
rect 393451 412996 393517 412997
rect 393451 412932 393452 412996
rect 393516 412932 393517 412996
rect 393451 412931 393517 412932
rect 392902 411710 392974 411770
rect 392166 411030 392820 411090
rect 392914 411060 392974 411710
rect 393454 411090 393514 412931
rect 394187 412724 394253 412725
rect 394187 412660 394188 412724
rect 394252 412660 394253 412724
rect 394187 412659 394253 412660
rect 394190 411770 394250 412659
rect 394082 411710 394250 411770
rect 393454 411030 393988 411090
rect 394082 411060 394142 411710
rect 394742 411090 394802 413475
rect 395291 412860 395357 412861
rect 395291 412796 395292 412860
rect 395356 412796 395357 412860
rect 395291 412795 395357 412796
rect 395294 411090 395354 412795
rect 394742 411030 395156 411090
rect 395280 411030 395354 411090
rect 372662 410690 372964 410750
rect 379654 410690 379972 410750
rect 381264 410690 381554 410750
rect 396030 410750 396090 413747
rect 397499 413404 397565 413405
rect 397499 413340 397500 413404
rect 397564 413340 397565 413404
rect 397499 413339 397565 413340
rect 396395 412996 396461 412997
rect 396395 412932 396396 412996
rect 396460 412932 396461 412996
rect 396395 412931 396461 412932
rect 396398 411770 396458 412931
rect 397502 411770 397562 413339
rect 396398 411710 396478 411770
rect 396418 411060 396478 411710
rect 397462 411710 397562 411770
rect 397462 411060 397522 411710
rect 397870 410750 397930 413883
rect 401547 413540 401613 413541
rect 401547 413476 401548 413540
rect 401612 413476 401613 413540
rect 401547 413475 401613 413476
rect 398051 413132 398117 413133
rect 398051 413068 398052 413132
rect 398116 413068 398117 413132
rect 398051 413067 398117 413068
rect 399891 413132 399957 413133
rect 399891 413068 399892 413132
rect 399956 413068 399957 413132
rect 399891 413067 399957 413068
rect 398054 411090 398114 413067
rect 398603 412996 398669 412997
rect 398603 412932 398604 412996
rect 398668 412932 398669 412996
rect 398603 412931 398669 412932
rect 398606 411770 398666 412931
rect 399155 412724 399221 412725
rect 399155 412660 399156 412724
rect 399220 412660 399221 412724
rect 399155 412659 399221 412660
rect 398606 411710 398814 411770
rect 398054 411030 398660 411090
rect 398754 411060 398814 411710
rect 399158 411090 399218 412659
rect 399894 411770 399954 413067
rect 400443 412860 400509 412861
rect 400443 412796 400444 412860
rect 400508 412796 400509 412860
rect 400443 412795 400509 412796
rect 399894 411710 399982 411770
rect 399158 411030 399828 411090
rect 399922 411060 399982 411710
rect 400446 411090 400506 412795
rect 401179 412724 401245 412725
rect 401179 412660 401180 412724
rect 401244 412660 401245 412724
rect 401179 412659 401245 412660
rect 401182 411770 401242 412659
rect 401090 411710 401242 411770
rect 400446 411030 400996 411090
rect 401090 411060 401150 411710
rect 401550 411090 401610 413475
rect 402283 413404 402349 413405
rect 402283 413340 402284 413404
rect 402348 413340 402349 413404
rect 402283 413339 402349 413340
rect 401550 411030 402164 411090
rect 402286 411030 402346 413339
rect 403022 411090 403082 413883
rect 404307 413540 404373 413541
rect 404307 413476 404308 413540
rect 404372 413476 404373 413540
rect 404307 413475 404373 413476
rect 403387 412860 403453 412861
rect 403387 412796 403388 412860
rect 403452 412796 403453 412860
rect 403387 412795 403453 412796
rect 403390 411770 403450 412795
rect 403390 411710 403486 411770
rect 403022 411030 403332 411090
rect 403426 411060 403486 411710
rect 404310 411090 404370 413475
rect 404675 413268 404741 413269
rect 404675 413204 404676 413268
rect 404740 413204 404741 413268
rect 404675 413203 404741 413204
rect 404678 411770 404738 413203
rect 404594 411710 404738 411770
rect 404310 411030 404500 411090
rect 404594 411060 404654 411710
rect 405759 411500 405825 411501
rect 405759 411436 405760 411500
rect 405824 411436 405825 411500
rect 405759 411435 405825 411436
rect 405762 411090 405822 411435
rect 407806 411090 407866 413883
rect 410566 411090 410626 413883
rect 413878 411090 413938 413883
rect 405762 411060 409296 411090
rect 405792 411030 409296 411060
rect 410464 411030 410626 411090
rect 413463 411030 413938 411090
rect 396030 410690 396324 410750
rect 397616 410690 397930 410750
rect 335604 409018 335786 409254
rect 336022 409018 336204 409254
rect 335604 408934 336204 409018
rect 335604 408698 335786 408934
rect 336022 408698 336204 408934
rect 335604 373254 336204 408698
rect 340482 409254 340802 409276
rect 340482 409018 340524 409254
rect 340760 409018 340802 409254
rect 340482 408934 340802 409018
rect 340482 408698 340524 408934
rect 340760 408698 340802 408934
rect 340482 408676 340802 408698
rect 340482 405654 340802 405676
rect 340482 405418 340524 405654
rect 340760 405418 340802 405654
rect 340482 405334 340802 405418
rect 340482 405098 340524 405334
rect 340760 405098 340802 405334
rect 340482 405076 340802 405098
rect 340482 402054 340802 402076
rect 340482 401818 340524 402054
rect 340760 401818 340802 402054
rect 340482 401734 340802 401818
rect 340482 401498 340524 401734
rect 340760 401498 340802 401734
rect 340482 401476 340802 401498
rect 340482 398454 340802 398476
rect 340482 398218 340524 398454
rect 340760 398218 340802 398454
rect 340482 398134 340802 398218
rect 340482 397898 340524 398134
rect 340760 397898 340802 398134
rect 340482 397876 340802 397898
rect 340034 391254 340358 391276
rect 340034 391018 340078 391254
rect 340314 391018 340358 391254
rect 340034 390934 340358 391018
rect 340034 390698 340078 390934
rect 340314 390698 340358 390934
rect 340034 390676 340358 390698
rect 340034 387654 340358 387676
rect 340034 387418 340078 387654
rect 340314 387418 340358 387654
rect 340034 387334 340358 387418
rect 340034 387098 340078 387334
rect 340314 387098 340358 387334
rect 340034 387076 340358 387098
rect 422004 387654 422604 423098
rect 422004 387418 422186 387654
rect 422422 387418 422604 387654
rect 422004 387334 422604 387418
rect 422004 387098 422186 387334
rect 422422 387098 422604 387334
rect 340034 384054 340358 384076
rect 340034 383818 340078 384054
rect 340314 383818 340358 384054
rect 340034 383734 340358 383818
rect 340034 383498 340078 383734
rect 340314 383498 340358 383734
rect 340034 383476 340358 383498
rect 340034 380454 340358 380476
rect 340034 380218 340078 380454
rect 340314 380218 340358 380454
rect 340034 380134 340358 380218
rect 340034 379898 340078 380134
rect 340314 379898 340358 380134
rect 340034 379876 340358 379898
rect 335604 373018 335786 373254
rect 336022 373018 336204 373254
rect 335604 372934 336204 373018
rect 335604 372698 335786 372934
rect 336022 372698 336204 372934
rect 335604 337254 336204 372698
rect 340482 373254 340802 373276
rect 340482 373018 340524 373254
rect 340760 373018 340802 373254
rect 340482 372934 340802 373018
rect 340482 372698 340524 372934
rect 340760 372698 340802 372934
rect 340482 372676 340802 372698
rect 340482 369654 340802 369676
rect 340482 369418 340524 369654
rect 340760 369418 340802 369654
rect 340482 369334 340802 369418
rect 340482 369098 340524 369334
rect 340760 369098 340802 369334
rect 340482 369076 340802 369098
rect 340482 366054 340802 366076
rect 340482 365818 340524 366054
rect 340760 365818 340802 366054
rect 340482 365734 340802 365818
rect 340482 365498 340524 365734
rect 340760 365498 340802 365734
rect 340482 365476 340802 365498
rect 340482 362454 340802 362476
rect 340482 362218 340524 362454
rect 340760 362218 340802 362454
rect 340482 362134 340802 362218
rect 340482 361898 340524 362134
rect 340760 361898 340802 362134
rect 340482 361876 340802 361898
rect 340034 355254 340358 355276
rect 340034 355018 340078 355254
rect 340314 355018 340358 355254
rect 340034 354934 340358 355018
rect 340034 354698 340078 354934
rect 340314 354698 340358 354934
rect 340034 354676 340358 354698
rect 340034 351654 340358 351676
rect 340034 351418 340078 351654
rect 340314 351418 340358 351654
rect 340034 351334 340358 351418
rect 340034 351098 340078 351334
rect 340314 351098 340358 351334
rect 340034 351076 340358 351098
rect 422004 351654 422604 387098
rect 422004 351418 422186 351654
rect 422422 351418 422604 351654
rect 422004 351334 422604 351418
rect 422004 351098 422186 351334
rect 422422 351098 422604 351334
rect 340034 348054 340358 348076
rect 340034 347818 340078 348054
rect 340314 347818 340358 348054
rect 340034 347734 340358 347818
rect 340034 347498 340078 347734
rect 340314 347498 340358 347734
rect 340034 347476 340358 347498
rect 419947 346628 420013 346629
rect 419947 346578 419948 346628
rect 420012 346578 420013 346628
rect 340034 344454 340358 344476
rect 340034 344218 340078 344454
rect 340314 344218 340358 344454
rect 340034 344134 340358 344218
rect 340034 343898 340078 344134
rect 340314 343898 340358 344134
rect 340034 343876 340358 343898
rect 420683 343772 420749 343773
rect 420683 343708 420684 343772
rect 420748 343708 420749 343772
rect 420683 343707 420749 343708
rect 420686 343178 420746 343707
rect 335604 337018 335786 337254
rect 336022 337018 336204 337254
rect 335604 336934 336204 337018
rect 335604 336698 335786 336934
rect 336022 336698 336204 336934
rect 335604 303000 336204 336698
rect 340482 337254 340802 337276
rect 340482 337018 340524 337254
rect 340760 337018 340802 337254
rect 340482 336934 340802 337018
rect 340482 336698 340524 336934
rect 340760 336698 340802 336934
rect 340482 336676 340802 336698
rect 340482 333654 340802 333676
rect 340482 333418 340524 333654
rect 340760 333418 340802 333654
rect 340482 333334 340802 333418
rect 340482 333098 340524 333334
rect 340760 333098 340802 333334
rect 340482 333076 340802 333098
rect 340482 330054 340802 330076
rect 340482 329818 340524 330054
rect 340760 329818 340802 330054
rect 340482 329734 340802 329818
rect 340482 329498 340524 329734
rect 340760 329498 340802 329734
rect 340482 329476 340802 329498
rect 340482 326454 340802 326476
rect 340482 326218 340524 326454
rect 340760 326218 340802 326454
rect 340482 326134 340802 326218
rect 340482 325898 340524 326134
rect 340760 325898 340802 326134
rect 340482 325876 340802 325898
rect 343693 320590 344018 320650
rect 343958 318749 344018 320590
rect 343955 318748 344021 318749
rect 343955 318684 343956 318748
rect 344020 318684 344021 318748
rect 343955 318683 344021 318684
rect 342804 308454 343404 317000
rect 342804 308218 342986 308454
rect 343222 308218 343404 308454
rect 342804 308134 343404 308218
rect 342804 307898 342986 308134
rect 343222 307898 343404 308134
rect 342804 303000 343404 307898
rect 346404 312054 347004 317000
rect 346404 311818 346586 312054
rect 346822 311818 347004 312054
rect 346404 311734 347004 311818
rect 346404 311498 346586 311734
rect 346822 311498 347004 311734
rect 346404 303000 347004 311498
rect 350004 315654 350604 317000
rect 350004 315418 350186 315654
rect 350422 315418 350604 315654
rect 350004 315334 350604 315418
rect 350004 315098 350186 315334
rect 350422 315098 350604 315334
rect 350004 303000 350604 315098
rect 353604 303000 354204 317000
rect 360804 303000 361404 317000
rect 364404 303000 365004 317000
rect 368004 303000 368604 317000
rect 371604 303000 372204 317000
rect 378804 308454 379404 317000
rect 378804 308218 378986 308454
rect 379222 308218 379404 308454
rect 378804 308134 379404 308218
rect 378804 307898 378986 308134
rect 379222 307898 379404 308134
rect 378804 303000 379404 307898
rect 382404 312054 383004 317000
rect 382404 311818 382586 312054
rect 382822 311818 383004 312054
rect 382404 311734 383004 311818
rect 382404 311498 382586 311734
rect 382822 311498 383004 311734
rect 382404 303000 383004 311498
rect 386004 315654 386604 317000
rect 386004 315418 386186 315654
rect 386422 315418 386604 315654
rect 386004 315334 386604 315418
rect 386004 315098 386186 315334
rect 386422 315098 386604 315334
rect 386004 303000 386604 315098
rect 389604 303000 390204 317000
rect 396804 303000 397404 317000
rect 400404 303000 401004 317000
rect 404004 303000 404604 317000
rect 407604 303000 408204 317000
rect 414804 308454 415404 317000
rect 414804 308218 414986 308454
rect 415222 308218 415404 308454
rect 414804 308134 415404 308218
rect 414804 307898 414986 308134
rect 415222 307898 415404 308134
rect 414804 303000 415404 307898
rect 418404 312054 419004 317000
rect 418404 311818 418586 312054
rect 418822 311818 419004 312054
rect 418404 311734 419004 311818
rect 418404 311498 418586 311734
rect 418822 311498 419004 311734
rect 418404 303000 419004 311498
rect 422004 315654 422604 351098
rect 425604 679254 426204 710862
rect 443604 710478 444204 711440
rect 443604 710242 443786 710478
rect 444022 710242 444204 710478
rect 443604 710158 444204 710242
rect 443604 709922 443786 710158
rect 444022 709922 444204 710158
rect 440004 708598 440604 709560
rect 440004 708362 440186 708598
rect 440422 708362 440604 708598
rect 440004 708278 440604 708362
rect 440004 708042 440186 708278
rect 440422 708042 440604 708278
rect 436404 706718 437004 707680
rect 436404 706482 436586 706718
rect 436822 706482 437004 706718
rect 436404 706398 437004 706482
rect 436404 706162 436586 706398
rect 436822 706162 437004 706398
rect 425604 679018 425786 679254
rect 426022 679018 426204 679254
rect 425604 678934 426204 679018
rect 425604 678698 425786 678934
rect 426022 678698 426204 678934
rect 425604 643254 426204 678698
rect 425604 643018 425786 643254
rect 426022 643018 426204 643254
rect 425604 642934 426204 643018
rect 425604 642698 425786 642934
rect 426022 642698 426204 642934
rect 425604 607254 426204 642698
rect 425604 607018 425786 607254
rect 426022 607018 426204 607254
rect 425604 606934 426204 607018
rect 425604 606698 425786 606934
rect 426022 606698 426204 606934
rect 425604 571254 426204 606698
rect 425604 571018 425786 571254
rect 426022 571018 426204 571254
rect 425604 570934 426204 571018
rect 425604 570698 425786 570934
rect 426022 570698 426204 570934
rect 425604 535254 426204 570698
rect 425604 535018 425786 535254
rect 426022 535018 426204 535254
rect 425604 534934 426204 535018
rect 425604 534698 425786 534934
rect 426022 534698 426204 534934
rect 425604 499254 426204 534698
rect 425604 499018 425786 499254
rect 426022 499018 426204 499254
rect 425604 498934 426204 499018
rect 425604 498698 425786 498934
rect 426022 498698 426204 498934
rect 425604 463254 426204 498698
rect 425604 463018 425786 463254
rect 426022 463018 426204 463254
rect 425604 462934 426204 463018
rect 425604 462698 425786 462934
rect 426022 462698 426204 462934
rect 425604 427254 426204 462698
rect 425604 427018 425786 427254
rect 426022 427018 426204 427254
rect 425604 426934 426204 427018
rect 425604 426698 425786 426934
rect 426022 426698 426204 426934
rect 425604 391254 426204 426698
rect 425604 391018 425786 391254
rect 426022 391018 426204 391254
rect 425604 390934 426204 391018
rect 425604 390698 425786 390934
rect 426022 390698 426204 390934
rect 425604 355254 426204 390698
rect 425604 355018 425786 355254
rect 426022 355018 426204 355254
rect 425604 354934 426204 355018
rect 425604 354698 425786 354934
rect 426022 354698 426204 354934
rect 422004 315418 422186 315654
rect 422422 315418 422604 315654
rect 422004 315334 422604 315418
rect 422004 315098 422186 315334
rect 422422 315098 422604 315334
rect 422004 303000 422604 315098
rect 425604 319254 426204 354698
rect 432804 704838 433404 705800
rect 432804 704602 432986 704838
rect 433222 704602 433404 704838
rect 432804 704518 433404 704602
rect 432804 704282 432986 704518
rect 433222 704282 433404 704518
rect 432804 686454 433404 704282
rect 432804 686218 432986 686454
rect 433222 686218 433404 686454
rect 432804 686134 433404 686218
rect 432804 685898 432986 686134
rect 433222 685898 433404 686134
rect 432804 650454 433404 685898
rect 436404 690054 437004 706162
rect 436404 689818 436586 690054
rect 436822 689818 437004 690054
rect 436404 689734 437004 689818
rect 436404 689498 436586 689734
rect 436822 689498 437004 689734
rect 436404 654247 437004 689498
rect 440004 693654 440604 708042
rect 440004 693418 440186 693654
rect 440422 693418 440604 693654
rect 440004 693334 440604 693418
rect 440004 693098 440186 693334
rect 440422 693098 440604 693334
rect 440004 657654 440604 693098
rect 440004 657418 440186 657654
rect 440422 657418 440604 657654
rect 440004 657334 440604 657418
rect 440004 657098 440186 657334
rect 440422 657098 440604 657334
rect 440004 654247 440604 657098
rect 443604 697254 444204 709922
rect 461604 711418 462204 711440
rect 461604 711182 461786 711418
rect 462022 711182 462204 711418
rect 461604 711098 462204 711182
rect 461604 710862 461786 711098
rect 462022 710862 462204 711098
rect 458004 709538 458604 709560
rect 458004 709302 458186 709538
rect 458422 709302 458604 709538
rect 458004 709218 458604 709302
rect 458004 708982 458186 709218
rect 458422 708982 458604 709218
rect 454404 707658 455004 707680
rect 454404 707422 454586 707658
rect 454822 707422 455004 707658
rect 454404 707338 455004 707422
rect 454404 707102 454586 707338
rect 454822 707102 455004 707338
rect 443604 697018 443786 697254
rect 444022 697018 444204 697254
rect 443604 696934 444204 697018
rect 443604 696698 443786 696934
rect 444022 696698 444204 696934
rect 443604 661254 444204 696698
rect 443604 661018 443786 661254
rect 444022 661018 444204 661254
rect 443604 660934 444204 661018
rect 443604 660698 443786 660934
rect 444022 660698 444204 660934
rect 443604 654247 444204 660698
rect 450804 705778 451404 705800
rect 450804 705542 450986 705778
rect 451222 705542 451404 705778
rect 450804 705458 451404 705542
rect 450804 705222 450986 705458
rect 451222 705222 451404 705458
rect 450804 668454 451404 705222
rect 450804 668218 450986 668454
rect 451222 668218 451404 668454
rect 450804 668134 451404 668218
rect 450804 667898 450986 668134
rect 451222 667898 451404 668134
rect 450804 654247 451404 667898
rect 454404 672054 455004 707102
rect 454404 671818 454586 672054
rect 454822 671818 455004 672054
rect 454404 671734 455004 671818
rect 454404 671498 454586 671734
rect 454822 671498 455004 671734
rect 454404 654247 455004 671498
rect 458004 675654 458604 708982
rect 458004 675418 458186 675654
rect 458422 675418 458604 675654
rect 458004 675334 458604 675418
rect 458004 675098 458186 675334
rect 458422 675098 458604 675334
rect 458004 654247 458604 675098
rect 461604 679254 462204 710862
rect 479604 710478 480204 711440
rect 479604 710242 479786 710478
rect 480022 710242 480204 710478
rect 479604 710158 480204 710242
rect 479604 709922 479786 710158
rect 480022 709922 480204 710158
rect 476004 708598 476604 709560
rect 476004 708362 476186 708598
rect 476422 708362 476604 708598
rect 476004 708278 476604 708362
rect 476004 708042 476186 708278
rect 476422 708042 476604 708278
rect 472404 706718 473004 707680
rect 472404 706482 472586 706718
rect 472822 706482 473004 706718
rect 472404 706398 473004 706482
rect 472404 706162 472586 706398
rect 472822 706162 473004 706398
rect 461604 679018 461786 679254
rect 462022 679018 462204 679254
rect 461604 678934 462204 679018
rect 461604 678698 461786 678934
rect 462022 678698 462204 678934
rect 461604 654247 462204 678698
rect 468804 704838 469404 705800
rect 468804 704602 468986 704838
rect 469222 704602 469404 704838
rect 468804 704518 469404 704602
rect 468804 704282 468986 704518
rect 469222 704282 469404 704518
rect 468804 686454 469404 704282
rect 468804 686218 468986 686454
rect 469222 686218 469404 686454
rect 468804 686134 469404 686218
rect 468804 685898 468986 686134
rect 469222 685898 469404 686134
rect 468804 654247 469404 685898
rect 472404 690054 473004 706162
rect 472404 689818 472586 690054
rect 472822 689818 473004 690054
rect 472404 689734 473004 689818
rect 472404 689498 472586 689734
rect 472822 689498 473004 689734
rect 472404 654247 473004 689498
rect 476004 693654 476604 708042
rect 476004 693418 476186 693654
rect 476422 693418 476604 693654
rect 476004 693334 476604 693418
rect 476004 693098 476186 693334
rect 476422 693098 476604 693334
rect 476004 657654 476604 693098
rect 476004 657418 476186 657654
rect 476422 657418 476604 657654
rect 476004 657334 476604 657418
rect 476004 657098 476186 657334
rect 476422 657098 476604 657334
rect 476004 654247 476604 657098
rect 479604 697254 480204 709922
rect 497604 711418 498204 711440
rect 497604 711182 497786 711418
rect 498022 711182 498204 711418
rect 497604 711098 498204 711182
rect 497604 710862 497786 711098
rect 498022 710862 498204 711098
rect 494004 709538 494604 709560
rect 494004 709302 494186 709538
rect 494422 709302 494604 709538
rect 494004 709218 494604 709302
rect 494004 708982 494186 709218
rect 494422 708982 494604 709218
rect 490404 707658 491004 707680
rect 490404 707422 490586 707658
rect 490822 707422 491004 707658
rect 490404 707338 491004 707422
rect 490404 707102 490586 707338
rect 490822 707102 491004 707338
rect 479604 697018 479786 697254
rect 480022 697018 480204 697254
rect 479604 696934 480204 697018
rect 479604 696698 479786 696934
rect 480022 696698 480204 696934
rect 479604 661254 480204 696698
rect 479604 661018 479786 661254
rect 480022 661018 480204 661254
rect 479604 660934 480204 661018
rect 479604 660698 479786 660934
rect 480022 660698 480204 660934
rect 479604 654247 480204 660698
rect 486804 705778 487404 705800
rect 486804 705542 486986 705778
rect 487222 705542 487404 705778
rect 486804 705458 487404 705542
rect 486804 705222 486986 705458
rect 487222 705222 487404 705458
rect 486804 668454 487404 705222
rect 486804 668218 486986 668454
rect 487222 668218 487404 668454
rect 486804 668134 487404 668218
rect 486804 667898 486986 668134
rect 487222 667898 487404 668134
rect 486804 654247 487404 667898
rect 490404 672054 491004 707102
rect 490404 671818 490586 672054
rect 490822 671818 491004 672054
rect 490404 671734 491004 671818
rect 490404 671498 490586 671734
rect 490822 671498 491004 671734
rect 490404 654247 491004 671498
rect 494004 675654 494604 708982
rect 494004 675418 494186 675654
rect 494422 675418 494604 675654
rect 494004 675334 494604 675418
rect 494004 675098 494186 675334
rect 494422 675098 494604 675334
rect 494004 654247 494604 675098
rect 497604 679254 498204 710862
rect 515604 710478 516204 711440
rect 515604 710242 515786 710478
rect 516022 710242 516204 710478
rect 515604 710158 516204 710242
rect 515604 709922 515786 710158
rect 516022 709922 516204 710158
rect 512004 708598 512604 709560
rect 512004 708362 512186 708598
rect 512422 708362 512604 708598
rect 512004 708278 512604 708362
rect 512004 708042 512186 708278
rect 512422 708042 512604 708278
rect 508404 706718 509004 707680
rect 508404 706482 508586 706718
rect 508822 706482 509004 706718
rect 508404 706398 509004 706482
rect 508404 706162 508586 706398
rect 508822 706162 509004 706398
rect 497604 679018 497786 679254
rect 498022 679018 498204 679254
rect 497604 678934 498204 679018
rect 497604 678698 497786 678934
rect 498022 678698 498204 678934
rect 497604 654247 498204 678698
rect 504804 704838 505404 705800
rect 504804 704602 504986 704838
rect 505222 704602 505404 704838
rect 504804 704518 505404 704602
rect 504804 704282 504986 704518
rect 505222 704282 505404 704518
rect 504804 686454 505404 704282
rect 504804 686218 504986 686454
rect 505222 686218 505404 686454
rect 504804 686134 505404 686218
rect 504804 685898 504986 686134
rect 505222 685898 505404 686134
rect 504804 654247 505404 685898
rect 508404 690054 509004 706162
rect 508404 689818 508586 690054
rect 508822 689818 509004 690054
rect 508404 689734 509004 689818
rect 508404 689498 508586 689734
rect 508822 689498 509004 689734
rect 508404 654247 509004 689498
rect 512004 693654 512604 708042
rect 512004 693418 512186 693654
rect 512422 693418 512604 693654
rect 512004 693334 512604 693418
rect 512004 693098 512186 693334
rect 512422 693098 512604 693334
rect 512004 657654 512604 693098
rect 512004 657418 512186 657654
rect 512422 657418 512604 657654
rect 512004 657334 512604 657418
rect 512004 657098 512186 657334
rect 512422 657098 512604 657334
rect 512004 654247 512604 657098
rect 515604 697254 516204 709922
rect 533604 711418 534204 711440
rect 533604 711182 533786 711418
rect 534022 711182 534204 711418
rect 533604 711098 534204 711182
rect 533604 710862 533786 711098
rect 534022 710862 534204 711098
rect 530004 709538 530604 709560
rect 530004 709302 530186 709538
rect 530422 709302 530604 709538
rect 530004 709218 530604 709302
rect 530004 708982 530186 709218
rect 530422 708982 530604 709218
rect 526404 707658 527004 707680
rect 526404 707422 526586 707658
rect 526822 707422 527004 707658
rect 526404 707338 527004 707422
rect 526404 707102 526586 707338
rect 526822 707102 527004 707338
rect 515604 697018 515786 697254
rect 516022 697018 516204 697254
rect 515604 696934 516204 697018
rect 515604 696698 515786 696934
rect 516022 696698 516204 696934
rect 515604 661254 516204 696698
rect 515604 661018 515786 661254
rect 516022 661018 516204 661254
rect 515604 660934 516204 661018
rect 515604 660698 515786 660934
rect 516022 660698 516204 660934
rect 515604 654247 516204 660698
rect 522804 705778 523404 705800
rect 522804 705542 522986 705778
rect 523222 705542 523404 705778
rect 522804 705458 523404 705542
rect 522804 705222 522986 705458
rect 523222 705222 523404 705458
rect 522804 668454 523404 705222
rect 522804 668218 522986 668454
rect 523222 668218 523404 668454
rect 522804 668134 523404 668218
rect 522804 667898 522986 668134
rect 523222 667898 523404 668134
rect 508451 652900 508517 652901
rect 508451 652836 508452 652900
rect 508516 652836 508517 652900
rect 508451 652835 508517 652836
rect 513419 652900 513485 652901
rect 513419 652836 513420 652900
rect 513484 652836 513485 652900
rect 513419 652835 513485 652836
rect 508454 651130 508514 652835
rect 513422 651130 513482 652835
rect 508454 651070 508608 651130
rect 513422 651070 513603 651130
rect 432804 650218 432986 650454
rect 433222 650218 433404 650454
rect 432804 650134 433404 650218
rect 432804 649898 432986 650134
rect 433222 649898 433404 650134
rect 432804 614454 433404 649898
rect 516938 643254 517262 643276
rect 516938 643018 516982 643254
rect 517218 643018 517262 643254
rect 516938 642934 517262 643018
rect 516938 642698 516982 642934
rect 517218 642698 517262 642934
rect 516938 642676 517262 642698
rect 516938 639654 517262 639676
rect 516938 639418 516982 639654
rect 517218 639418 517262 639654
rect 516938 639334 517262 639418
rect 516938 639098 516982 639334
rect 517218 639098 517262 639334
rect 516938 639076 517262 639098
rect 516938 636054 517262 636076
rect 516938 635818 516982 636054
rect 517218 635818 517262 636054
rect 516938 635734 517262 635818
rect 516938 635498 516982 635734
rect 517218 635498 517262 635734
rect 516938 635476 517262 635498
rect 516938 632454 517262 632476
rect 516938 632218 516982 632454
rect 517218 632218 517262 632454
rect 516938 632134 517262 632218
rect 516938 631898 516982 632134
rect 517218 631898 517262 632134
rect 516938 631876 517262 631898
rect 522804 632454 523404 667898
rect 522804 632218 522986 632454
rect 523222 632218 523404 632454
rect 522804 632134 523404 632218
rect 522804 631898 522986 632134
rect 523222 631898 523404 632134
rect 516494 625254 516814 625276
rect 516494 625018 516536 625254
rect 516772 625018 516814 625254
rect 516494 624934 516814 625018
rect 516494 624698 516536 624934
rect 516772 624698 516814 624934
rect 516494 624676 516814 624698
rect 516494 621654 516814 621676
rect 516494 621418 516536 621654
rect 516772 621418 516814 621654
rect 516494 621334 516814 621418
rect 516494 621098 516536 621334
rect 516772 621098 516814 621334
rect 516494 621076 516814 621098
rect 516494 618054 516814 618076
rect 516494 617818 516536 618054
rect 516772 617818 516814 618054
rect 516494 617734 516814 617818
rect 516494 617498 516536 617734
rect 516772 617498 516814 617734
rect 516494 617476 516814 617498
rect 432804 614218 432986 614454
rect 433222 614218 433404 614454
rect 432804 614134 433404 614218
rect 432804 613898 432986 614134
rect 433222 613898 433404 614134
rect 432804 578454 433404 613898
rect 516494 614454 516814 614476
rect 516494 614218 516536 614454
rect 516772 614218 516814 614454
rect 516494 614134 516814 614218
rect 516494 613898 516536 614134
rect 516772 613898 516814 614134
rect 516494 613876 516814 613898
rect 516938 607254 517262 607276
rect 516938 607018 516982 607254
rect 517218 607018 517262 607254
rect 516938 606934 517262 607018
rect 516938 606698 516982 606934
rect 517218 606698 517262 606934
rect 516938 606676 517262 606698
rect 516938 603654 517262 603676
rect 516938 603418 516982 603654
rect 517218 603418 517262 603654
rect 516938 603334 517262 603418
rect 516938 603098 516982 603334
rect 517218 603098 517262 603334
rect 516938 603076 517262 603098
rect 516938 600054 517262 600076
rect 516938 599818 516982 600054
rect 517218 599818 517262 600054
rect 516938 599734 517262 599818
rect 516938 599498 516982 599734
rect 517218 599498 517262 599734
rect 516938 599476 517262 599498
rect 516938 596454 517262 596476
rect 516938 596218 516982 596454
rect 517218 596218 517262 596454
rect 516938 596134 517262 596218
rect 516938 595898 516982 596134
rect 517218 595898 517262 596134
rect 516938 595876 517262 595898
rect 522804 596454 523404 631898
rect 522804 596218 522986 596454
rect 523222 596218 523404 596454
rect 522804 596134 523404 596218
rect 522804 595898 522986 596134
rect 523222 595898 523404 596134
rect 516494 589254 516814 589276
rect 516494 589018 516536 589254
rect 516772 589018 516814 589254
rect 516494 588934 516814 589018
rect 516494 588698 516536 588934
rect 516772 588698 516814 588934
rect 516494 588676 516814 588698
rect 516494 585654 516814 585676
rect 516494 585418 516536 585654
rect 516772 585418 516814 585654
rect 516494 585334 516814 585418
rect 516494 585098 516536 585334
rect 516772 585098 516814 585334
rect 516494 585076 516814 585098
rect 516494 582054 516814 582076
rect 516494 581818 516536 582054
rect 516772 581818 516814 582054
rect 516494 581734 516814 581818
rect 516494 581498 516536 581734
rect 516772 581498 516814 581734
rect 516494 581476 516814 581498
rect 518939 580956 519005 580957
rect 518939 580892 518940 580956
rect 519004 580892 519005 580956
rect 518939 580891 519005 580892
rect 518942 579818 519002 580891
rect 432804 578218 432986 578454
rect 433222 578218 433404 578454
rect 432804 578134 433404 578218
rect 432804 577898 432986 578134
rect 433222 577898 433404 578134
rect 432804 542454 433404 577898
rect 516494 578454 516814 578476
rect 516494 578218 516536 578454
rect 516772 578218 516814 578454
rect 516494 578134 516814 578218
rect 516494 577898 516536 578134
rect 516772 577898 516814 578134
rect 516494 577876 516814 577898
rect 516938 571254 517262 571276
rect 516938 571018 516982 571254
rect 517218 571018 517262 571254
rect 516938 570934 517262 571018
rect 516938 570698 516982 570934
rect 517218 570698 517262 570934
rect 516938 570676 517262 570698
rect 516938 567654 517262 567676
rect 516938 567418 516982 567654
rect 517218 567418 517262 567654
rect 516938 567334 517262 567418
rect 516938 567098 516982 567334
rect 517218 567098 517262 567334
rect 516938 567076 517262 567098
rect 516938 564054 517262 564076
rect 516938 563818 516982 564054
rect 517218 563818 517262 564054
rect 516938 563734 517262 563818
rect 516938 563498 516982 563734
rect 517218 563498 517262 563734
rect 516938 563476 517262 563498
rect 454726 560430 455008 560490
rect 456300 560430 456626 560490
rect 459804 560430 460122 560490
rect 443134 560290 443833 560350
rect 446262 560290 446832 560350
rect 447366 560290 448000 560350
rect 448470 560290 449168 560350
rect 449942 560290 450336 560350
rect 451414 560290 451504 560350
rect 443134 558925 443194 560290
rect 446262 558925 446322 560290
rect 443131 558924 443197 558925
rect 443131 558860 443132 558924
rect 443196 558860 443197 558924
rect 443131 558859 443197 558860
rect 446259 558924 446325 558925
rect 446259 558860 446260 558924
rect 446324 558860 446325 558924
rect 446259 558859 446325 558860
rect 447366 558381 447426 560290
rect 447363 558380 447429 558381
rect 447363 558316 447364 558380
rect 447428 558316 447429 558380
rect 447363 558315 447429 558316
rect 448470 558245 448530 560290
rect 448467 558244 448533 558245
rect 448467 558180 448468 558244
rect 448532 558180 448533 558244
rect 448467 558179 448533 558180
rect 449942 557837 450002 560290
rect 451414 558925 451474 560290
rect 452642 559330 452702 560320
rect 452796 560290 452946 560350
rect 452642 559270 452762 559330
rect 451411 558924 451477 558925
rect 451411 558860 451412 558924
rect 451476 558860 451477 558924
rect 451411 558859 451477 558860
rect 452702 558653 452762 559270
rect 452886 558925 452946 560290
rect 453622 560290 453840 560350
rect 453622 558925 453682 560290
rect 453934 559330 453994 560320
rect 453806 559270 453994 559330
rect 452883 558924 452949 558925
rect 452883 558860 452884 558924
rect 452948 558860 452949 558924
rect 452883 558859 452949 558860
rect 453619 558924 453685 558925
rect 453619 558860 453620 558924
rect 453684 558860 453685 558924
rect 453619 558859 453685 558860
rect 453806 558789 453866 559270
rect 454726 558789 454786 560430
rect 455132 560290 455338 560350
rect 455278 558925 455338 560290
rect 456014 560290 456176 560350
rect 455275 558924 455341 558925
rect 455275 558860 455276 558924
rect 455340 558860 455341 558924
rect 455275 558859 455341 558860
rect 456014 558789 456074 560290
rect 456566 558925 456626 560430
rect 456563 558924 456629 558925
rect 456563 558860 456564 558924
rect 456628 558860 456629 558924
rect 456563 558859 456629 558860
rect 457302 558789 457362 560350
rect 457468 560290 457546 560350
rect 457486 558925 457546 560290
rect 458482 560010 458542 560320
rect 458636 560290 458834 560350
rect 458406 559950 458542 560010
rect 457483 558924 457549 558925
rect 457483 558860 457484 558924
rect 457548 558860 457549 558924
rect 457483 558859 457549 558860
rect 458406 558789 458466 559950
rect 458774 558925 458834 560290
rect 459510 560290 459680 560350
rect 458771 558924 458837 558925
rect 458771 558860 458772 558924
rect 458836 558860 458837 558924
rect 458771 558859 458837 558860
rect 453803 558788 453869 558789
rect 453803 558724 453804 558788
rect 453868 558724 453869 558788
rect 453803 558723 453869 558724
rect 454723 558788 454789 558789
rect 454723 558724 454724 558788
rect 454788 558724 454789 558788
rect 454723 558723 454789 558724
rect 456011 558788 456077 558789
rect 456011 558724 456012 558788
rect 456076 558724 456077 558788
rect 456011 558723 456077 558724
rect 457299 558788 457365 558789
rect 457299 558724 457300 558788
rect 457364 558724 457365 558788
rect 457299 558723 457365 558724
rect 458403 558788 458469 558789
rect 458403 558724 458404 558788
rect 458468 558724 458469 558788
rect 458403 558723 458469 558724
rect 459510 558653 459570 560290
rect 460062 558925 460122 560430
rect 468710 560430 469024 560490
rect 472206 560430 472528 560490
rect 473820 560430 474106 560490
rect 460059 558924 460125 558925
rect 460059 558860 460060 558924
rect 460124 558860 460125 558924
rect 460059 558859 460125 558860
rect 452699 558652 452765 558653
rect 452699 558588 452700 558652
rect 452764 558588 452765 558652
rect 452699 558587 452765 558588
rect 459507 558652 459573 558653
rect 459507 558588 459508 558652
rect 459572 558588 459573 558652
rect 459507 558587 459573 558588
rect 449939 557836 450005 557837
rect 449939 557772 449940 557836
rect 450004 557772 450005 557836
rect 449939 557771 450005 557772
rect 460798 557701 460858 560350
rect 460972 560290 461042 560350
rect 460982 558925 461042 560290
rect 461718 560290 462016 560350
rect 461718 558925 461778 560290
rect 462110 559330 462170 560320
rect 462086 559270 462170 559330
rect 463006 560290 463184 560350
rect 460979 558924 461045 558925
rect 460979 558860 460980 558924
rect 461044 558860 461045 558924
rect 460979 558859 461045 558860
rect 461715 558924 461781 558925
rect 461715 558860 461716 558924
rect 461780 558860 461781 558924
rect 461715 558859 461781 558860
rect 462086 558789 462146 559270
rect 463006 558789 463066 560290
rect 463278 560010 463338 560320
rect 463278 559950 463434 560010
rect 463374 558925 463434 559950
rect 463371 558924 463437 558925
rect 463371 558860 463372 558924
rect 463436 558860 463437 558924
rect 463371 558859 463437 558860
rect 464294 558789 464354 560350
rect 464476 560290 464538 560350
rect 464478 558925 464538 560290
rect 465214 560290 465520 560350
rect 465644 560290 465826 560350
rect 464475 558924 464541 558925
rect 464475 558860 464476 558924
rect 464540 558860 464541 558924
rect 464475 558859 464541 558860
rect 465214 558789 465274 560290
rect 465766 558925 465826 560290
rect 466502 560290 466688 560350
rect 465763 558924 465829 558925
rect 465763 558860 465764 558924
rect 465828 558860 465829 558924
rect 465763 558859 465829 558860
rect 466502 558789 466562 560290
rect 466782 560010 466842 560320
rect 467790 560290 467856 560350
rect 466782 559950 466930 560010
rect 466870 558925 466930 559950
rect 466867 558924 466933 558925
rect 466867 558860 466868 558924
rect 466932 558860 466933 558924
rect 466867 558859 466933 558860
rect 462083 558788 462149 558789
rect 462083 558724 462084 558788
rect 462148 558724 462149 558788
rect 462083 558723 462149 558724
rect 463003 558788 463069 558789
rect 463003 558724 463004 558788
rect 463068 558724 463069 558788
rect 463003 558723 463069 558724
rect 464291 558788 464357 558789
rect 464291 558724 464292 558788
rect 464356 558724 464357 558788
rect 464291 558723 464357 558724
rect 465211 558788 465277 558789
rect 465211 558724 465212 558788
rect 465276 558724 465277 558788
rect 465211 558723 465277 558724
rect 466499 558788 466565 558789
rect 466499 558724 466500 558788
rect 466564 558724 466565 558788
rect 466499 558723 466565 558724
rect 467790 558653 467850 560290
rect 467974 558925 468034 560350
rect 468710 558925 468770 560430
rect 469118 559330 469178 560320
rect 469078 559270 469178 559330
rect 469998 560290 470192 560350
rect 467971 558924 468037 558925
rect 467971 558860 467972 558924
rect 468036 558860 468037 558924
rect 467971 558859 468037 558860
rect 468707 558924 468773 558925
rect 468707 558860 468708 558924
rect 468772 558860 468773 558924
rect 468707 558859 468773 558860
rect 469078 558789 469138 559270
rect 469075 558788 469141 558789
rect 469075 558724 469076 558788
rect 469140 558724 469141 558788
rect 469075 558723 469141 558724
rect 469998 558653 470058 560290
rect 470286 560010 470346 560320
rect 471286 560290 471360 560350
rect 470286 559950 470426 560010
rect 470366 558925 470426 559950
rect 470363 558924 470429 558925
rect 470363 558860 470364 558924
rect 470428 558860 470429 558924
rect 470363 558859 470429 558860
rect 471286 558789 471346 560290
rect 471470 558925 471530 560350
rect 471467 558924 471533 558925
rect 471467 558860 471468 558924
rect 471532 558860 471533 558924
rect 471467 558859 471533 558860
rect 472206 558789 472266 560430
rect 472652 560290 472818 560350
rect 472758 558925 472818 560290
rect 473494 560290 473696 560350
rect 472755 558924 472821 558925
rect 472755 558860 472756 558924
rect 472820 558860 472821 558924
rect 472755 558859 472821 558860
rect 473494 558789 473554 560290
rect 474046 558925 474106 560430
rect 481590 560430 481872 560490
rect 483164 560430 483490 560490
rect 486668 560430 486986 560490
rect 474782 560290 474864 560350
rect 474043 558924 474109 558925
rect 474043 558860 474044 558924
rect 474108 558860 474109 558924
rect 474043 558859 474109 558860
rect 474782 558789 474842 560290
rect 474966 558925 475026 560350
rect 475518 560290 476032 560350
rect 476156 560290 476314 560350
rect 475518 558925 475578 560290
rect 476254 558925 476314 560290
rect 476622 560290 477200 560350
rect 476622 558925 476682 560290
rect 477294 560010 477354 560320
rect 477910 560290 478368 560350
rect 477294 559950 477418 560010
rect 474963 558924 475029 558925
rect 474963 558860 474964 558924
rect 475028 558860 475029 558924
rect 474963 558859 475029 558860
rect 475515 558924 475581 558925
rect 475515 558860 475516 558924
rect 475580 558860 475581 558924
rect 475515 558859 475581 558860
rect 476251 558924 476317 558925
rect 476251 558860 476252 558924
rect 476316 558860 476317 558924
rect 476251 558859 476317 558860
rect 476619 558924 476685 558925
rect 476619 558860 476620 558924
rect 476684 558860 476685 558924
rect 476619 558859 476685 558860
rect 471283 558788 471349 558789
rect 471283 558724 471284 558788
rect 471348 558724 471349 558788
rect 471283 558723 471349 558724
rect 472203 558788 472269 558789
rect 472203 558724 472204 558788
rect 472268 558724 472269 558788
rect 472203 558723 472269 558724
rect 473491 558788 473557 558789
rect 473491 558724 473492 558788
rect 473556 558724 473557 558788
rect 473491 558723 473557 558724
rect 474779 558788 474845 558789
rect 474779 558724 474780 558788
rect 474844 558724 474845 558788
rect 474779 558723 474845 558724
rect 477358 558653 477418 559950
rect 477910 558925 477970 560290
rect 477907 558924 477973 558925
rect 477907 558860 477908 558924
rect 477972 558860 477973 558924
rect 477907 558859 477973 558860
rect 467787 558652 467853 558653
rect 467787 558588 467788 558652
rect 467852 558588 467853 558652
rect 467787 558587 467853 558588
rect 469995 558652 470061 558653
rect 469995 558588 469996 558652
rect 470060 558588 470061 558652
rect 469995 558587 470061 558588
rect 477355 558652 477421 558653
rect 477355 558588 477356 558652
rect 477420 558588 477421 558652
rect 477355 558587 477421 558588
rect 478462 558381 478522 560320
rect 479014 560290 479536 560350
rect 479660 560290 479810 560350
rect 479014 558925 479074 560290
rect 479011 558924 479077 558925
rect 479011 558860 479012 558924
rect 479076 558860 479077 558924
rect 479011 558859 479077 558860
rect 479750 558517 479810 560290
rect 480486 560290 480704 560350
rect 480828 560290 480914 560350
rect 480486 558925 480546 560290
rect 480483 558924 480549 558925
rect 480483 558860 480484 558924
rect 480548 558860 480549 558924
rect 480483 558859 480549 558860
rect 479747 558516 479813 558517
rect 479747 558452 479748 558516
rect 479812 558452 479813 558516
rect 479747 558451 479813 558452
rect 480854 558381 480914 560290
rect 481590 558653 481650 560430
rect 481996 560290 482202 560350
rect 481587 558652 481653 558653
rect 481587 558588 481588 558652
rect 481652 558588 481653 558652
rect 481587 558587 481653 558588
rect 482142 558517 482202 560290
rect 483010 559330 483070 560320
rect 483010 559270 483122 559330
rect 483062 558517 483122 559270
rect 482139 558516 482205 558517
rect 482139 558452 482140 558516
rect 482204 558452 482205 558516
rect 482139 558451 482205 558452
rect 483059 558516 483125 558517
rect 483059 558452 483060 558516
rect 483124 558452 483125 558516
rect 483059 558451 483125 558452
rect 478459 558380 478525 558381
rect 478459 558316 478460 558380
rect 478524 558316 478525 558380
rect 478459 558315 478525 558316
rect 480851 558380 480917 558381
rect 480851 558316 480852 558380
rect 480916 558316 480917 558380
rect 480851 558315 480917 558316
rect 483430 557973 483490 560430
rect 483614 560290 484208 560350
rect 483427 557972 483493 557973
rect 483427 557908 483428 557972
rect 483492 557908 483493 557972
rect 483427 557907 483493 557908
rect 483614 557837 483674 560290
rect 484302 559330 484362 560320
rect 484166 559270 484362 559330
rect 484718 560290 485376 560350
rect 485500 560290 485698 560350
rect 484166 558245 484226 559270
rect 484718 558789 484778 560290
rect 484715 558788 484781 558789
rect 484715 558724 484716 558788
rect 484780 558724 484781 558788
rect 484715 558723 484781 558724
rect 484163 558244 484229 558245
rect 484163 558180 484164 558244
rect 484228 558180 484229 558244
rect 484163 558179 484229 558180
rect 485638 558109 485698 560290
rect 486006 560290 486544 560350
rect 486006 558517 486066 560290
rect 486003 558516 486069 558517
rect 486003 558452 486004 558516
rect 486068 558452 486069 558516
rect 486003 558451 486069 558452
rect 485635 558108 485701 558109
rect 485635 558044 485636 558108
rect 485700 558044 485701 558108
rect 485635 558043 485701 558044
rect 486926 557973 486986 560430
rect 522804 560454 523404 595898
rect 487294 560290 487712 560350
rect 487836 560290 487906 560350
rect 487294 558517 487354 560290
rect 487291 558516 487357 558517
rect 487291 558452 487292 558516
rect 487356 558452 487357 558516
rect 487291 558451 487357 558452
rect 486923 557972 486989 557973
rect 486923 557908 486924 557972
rect 486988 557908 486989 557972
rect 486923 557907 486989 557908
rect 487846 557837 487906 560290
rect 488582 560290 488880 560350
rect 489004 560290 489194 560350
rect 488582 558381 488642 560290
rect 488579 558380 488645 558381
rect 488579 558316 488580 558380
rect 488644 558316 488645 558380
rect 488579 558315 488645 558316
rect 483611 557836 483677 557837
rect 483611 557772 483612 557836
rect 483676 557772 483677 557836
rect 483611 557771 483677 557772
rect 487843 557836 487909 557837
rect 487843 557772 487844 557836
rect 487908 557772 487909 557836
rect 487843 557771 487909 557772
rect 489134 557701 489194 560290
rect 522804 560218 522986 560454
rect 523222 560218 523404 560454
rect 522804 560134 523404 560218
rect 522804 559898 522986 560134
rect 523222 559898 523404 560134
rect 460795 557700 460861 557701
rect 460795 557636 460796 557700
rect 460860 557636 460861 557700
rect 460795 557635 460861 557636
rect 489131 557700 489197 557701
rect 489131 557636 489132 557700
rect 489196 557636 489197 557700
rect 489131 557635 489197 557636
rect 432804 542218 432986 542454
rect 433222 542218 433404 542454
rect 432804 542134 433404 542218
rect 432804 541898 432986 542134
rect 433222 541898 433404 542134
rect 432804 506454 433404 541898
rect 432804 506218 432986 506454
rect 433222 506218 433404 506454
rect 432804 506134 433404 506218
rect 432804 505898 432986 506134
rect 433222 505898 433404 506134
rect 432804 470454 433404 505898
rect 432804 470218 432986 470454
rect 433222 470218 433404 470454
rect 432804 470134 433404 470218
rect 432804 469898 432986 470134
rect 433222 469898 433404 470134
rect 432804 434454 433404 469898
rect 432804 434218 432986 434454
rect 433222 434218 433404 434454
rect 432804 434134 433404 434218
rect 432804 433898 432986 434134
rect 433222 433898 433404 434134
rect 432804 398454 433404 433898
rect 432804 398218 432986 398454
rect 433222 398218 433404 398454
rect 432804 398134 433404 398218
rect 432804 397898 432986 398134
rect 433222 397898 433404 398134
rect 432804 362454 433404 397898
rect 432804 362218 432986 362454
rect 433222 362218 433404 362454
rect 432804 362134 433404 362218
rect 432804 361898 432986 362134
rect 433222 361898 433404 362134
rect 427859 341188 427925 341189
rect 427859 341138 427860 341188
rect 427924 341138 427925 341188
rect 425604 319018 425786 319254
rect 426022 319018 426204 319254
rect 425604 318934 426204 319018
rect 425604 318698 425786 318934
rect 426022 318698 426204 318934
rect 425604 303000 426204 318698
rect 432804 326454 433404 361898
rect 432804 326218 432986 326454
rect 433222 326218 433404 326454
rect 432804 326134 433404 326218
rect 432804 325898 432986 326134
rect 433222 325898 433404 326134
rect 432804 303000 433404 325898
rect 436404 546054 437004 557000
rect 436404 545818 436586 546054
rect 436822 545818 437004 546054
rect 436404 545734 437004 545818
rect 436404 545498 436586 545734
rect 436822 545498 437004 545734
rect 436404 510054 437004 545498
rect 436404 509818 436586 510054
rect 436822 509818 437004 510054
rect 436404 509734 437004 509818
rect 436404 509498 436586 509734
rect 436822 509498 437004 509734
rect 436404 474054 437004 509498
rect 436404 473818 436586 474054
rect 436822 473818 437004 474054
rect 436404 473734 437004 473818
rect 436404 473498 436586 473734
rect 436822 473498 437004 473734
rect 436404 438054 437004 473498
rect 436404 437818 436586 438054
rect 436822 437818 437004 438054
rect 436404 437734 437004 437818
rect 436404 437498 436586 437734
rect 436822 437498 437004 437734
rect 436404 402054 437004 437498
rect 436404 401818 436586 402054
rect 436822 401818 437004 402054
rect 436404 401734 437004 401818
rect 436404 401498 436586 401734
rect 436822 401498 437004 401734
rect 436404 366054 437004 401498
rect 436404 365818 436586 366054
rect 436822 365818 437004 366054
rect 436404 365734 437004 365818
rect 436404 365498 436586 365734
rect 436822 365498 437004 365734
rect 436404 330054 437004 365498
rect 440004 549654 440604 557000
rect 440004 549418 440186 549654
rect 440422 549418 440604 549654
rect 440004 549334 440604 549418
rect 440004 549098 440186 549334
rect 440422 549098 440604 549334
rect 440004 513654 440604 549098
rect 440004 513418 440186 513654
rect 440422 513418 440604 513654
rect 440004 513334 440604 513418
rect 440004 513098 440186 513334
rect 440422 513098 440604 513334
rect 440004 477654 440604 513098
rect 440004 477418 440186 477654
rect 440422 477418 440604 477654
rect 440004 477334 440604 477418
rect 440004 477098 440186 477334
rect 440422 477098 440604 477334
rect 440004 441654 440604 477098
rect 440004 441418 440186 441654
rect 440422 441418 440604 441654
rect 440004 441334 440604 441418
rect 440004 441098 440186 441334
rect 440422 441098 440604 441334
rect 440004 405654 440604 441098
rect 440004 405418 440186 405654
rect 440422 405418 440604 405654
rect 440004 405334 440604 405418
rect 440004 405098 440186 405334
rect 440422 405098 440604 405334
rect 440004 369654 440604 405098
rect 440004 369418 440186 369654
rect 440422 369418 440604 369654
rect 440004 369334 440604 369418
rect 440004 369098 440186 369334
rect 440422 369098 440604 369334
rect 437798 344453 437858 344982
rect 437795 344452 437861 344453
rect 437795 344388 437796 344452
rect 437860 344388 437861 344452
rect 437795 344387 437861 344388
rect 439451 341188 439517 341189
rect 439451 341124 439452 341188
rect 439516 341124 439517 341188
rect 439451 341123 439517 341124
rect 439454 339778 439514 341123
rect 436404 329818 436586 330054
rect 436822 329818 437004 330054
rect 436404 329734 437004 329818
rect 436404 329498 436586 329734
rect 436822 329498 437004 329734
rect 436404 303000 437004 329498
rect 440004 333654 440604 369098
rect 440004 333418 440186 333654
rect 440422 333418 440604 333654
rect 440004 333334 440604 333418
rect 440004 333098 440186 333334
rect 440422 333098 440604 333334
rect 440004 303000 440604 333098
rect 443604 553254 444204 557000
rect 443604 553018 443786 553254
rect 444022 553018 444204 553254
rect 443604 552934 444204 553018
rect 443604 552698 443786 552934
rect 444022 552698 444204 552934
rect 443604 517254 444204 552698
rect 443604 517018 443786 517254
rect 444022 517018 444204 517254
rect 443604 516934 444204 517018
rect 443604 516698 443786 516934
rect 444022 516698 444204 516934
rect 443604 481254 444204 516698
rect 443604 481018 443786 481254
rect 444022 481018 444204 481254
rect 443604 480934 444204 481018
rect 443604 480698 443786 480934
rect 444022 480698 444204 480934
rect 443604 445254 444204 480698
rect 443604 445018 443786 445254
rect 444022 445018 444204 445254
rect 443604 444934 444204 445018
rect 443604 444698 443786 444934
rect 444022 444698 444204 444934
rect 443604 409254 444204 444698
rect 450804 524454 451404 557000
rect 450804 524218 450986 524454
rect 451222 524218 451404 524454
rect 450804 524134 451404 524218
rect 450804 523898 450986 524134
rect 451222 523898 451404 524134
rect 450804 488454 451404 523898
rect 450804 488218 450986 488454
rect 451222 488218 451404 488454
rect 450804 488134 451404 488218
rect 450804 487898 450986 488134
rect 451222 487898 451404 488134
rect 450804 452454 451404 487898
rect 450804 452218 450986 452454
rect 451222 452218 451404 452454
rect 450804 452134 451404 452218
rect 450804 451898 450986 452134
rect 451222 451898 451404 452134
rect 450804 416454 451404 451898
rect 450804 416218 450986 416454
rect 451222 416218 451404 416454
rect 450804 416134 451404 416218
rect 450804 415898 450986 416134
rect 451222 415898 451404 416134
rect 450804 414247 451404 415898
rect 454404 528054 455004 557000
rect 454404 527818 454586 528054
rect 454822 527818 455004 528054
rect 454404 527734 455004 527818
rect 454404 527498 454586 527734
rect 454822 527498 455004 527734
rect 454404 492054 455004 527498
rect 454404 491818 454586 492054
rect 454822 491818 455004 492054
rect 454404 491734 455004 491818
rect 454404 491498 454586 491734
rect 454822 491498 455004 491734
rect 454404 456054 455004 491498
rect 454404 455818 454586 456054
rect 454822 455818 455004 456054
rect 454404 455734 455004 455818
rect 454404 455498 454586 455734
rect 454822 455498 455004 455734
rect 454404 420054 455004 455498
rect 454404 419818 454586 420054
rect 454822 419818 455004 420054
rect 454404 419734 455004 419818
rect 454404 419498 454586 419734
rect 454822 419498 455004 419734
rect 454404 414247 455004 419498
rect 458004 531654 458604 557000
rect 458004 531418 458186 531654
rect 458422 531418 458604 531654
rect 458004 531334 458604 531418
rect 458004 531098 458186 531334
rect 458422 531098 458604 531334
rect 458004 495654 458604 531098
rect 458004 495418 458186 495654
rect 458422 495418 458604 495654
rect 458004 495334 458604 495418
rect 458004 495098 458186 495334
rect 458422 495098 458604 495334
rect 458004 459654 458604 495098
rect 458004 459418 458186 459654
rect 458422 459418 458604 459654
rect 458004 459334 458604 459418
rect 458004 459098 458186 459334
rect 458422 459098 458604 459334
rect 458004 423654 458604 459098
rect 458004 423418 458186 423654
rect 458422 423418 458604 423654
rect 458004 423334 458604 423418
rect 458004 423098 458186 423334
rect 458422 423098 458604 423334
rect 458004 414247 458604 423098
rect 461604 535254 462204 557000
rect 461604 535018 461786 535254
rect 462022 535018 462204 535254
rect 461604 534934 462204 535018
rect 461604 534698 461786 534934
rect 462022 534698 462204 534934
rect 461604 499254 462204 534698
rect 461604 499018 461786 499254
rect 462022 499018 462204 499254
rect 461604 498934 462204 499018
rect 461604 498698 461786 498934
rect 462022 498698 462204 498934
rect 461604 463254 462204 498698
rect 461604 463018 461786 463254
rect 462022 463018 462204 463254
rect 461604 462934 462204 463018
rect 461604 462698 461786 462934
rect 462022 462698 462204 462934
rect 461604 427254 462204 462698
rect 461604 427018 461786 427254
rect 462022 427018 462204 427254
rect 461604 426934 462204 427018
rect 461604 426698 461786 426934
rect 462022 426698 462204 426934
rect 461604 414247 462204 426698
rect 468804 542454 469404 557000
rect 468804 542218 468986 542454
rect 469222 542218 469404 542454
rect 468804 542134 469404 542218
rect 468804 541898 468986 542134
rect 469222 541898 469404 542134
rect 468804 506454 469404 541898
rect 468804 506218 468986 506454
rect 469222 506218 469404 506454
rect 468804 506134 469404 506218
rect 468804 505898 468986 506134
rect 469222 505898 469404 506134
rect 468804 470454 469404 505898
rect 468804 470218 468986 470454
rect 469222 470218 469404 470454
rect 468804 470134 469404 470218
rect 468804 469898 468986 470134
rect 469222 469898 469404 470134
rect 468804 434454 469404 469898
rect 468804 434218 468986 434454
rect 469222 434218 469404 434454
rect 468804 434134 469404 434218
rect 468804 433898 468986 434134
rect 469222 433898 469404 434134
rect 468804 414247 469404 433898
rect 472404 546054 473004 557000
rect 472404 545818 472586 546054
rect 472822 545818 473004 546054
rect 472404 545734 473004 545818
rect 472404 545498 472586 545734
rect 472822 545498 473004 545734
rect 472404 510054 473004 545498
rect 472404 509818 472586 510054
rect 472822 509818 473004 510054
rect 472404 509734 473004 509818
rect 472404 509498 472586 509734
rect 472822 509498 473004 509734
rect 472404 474054 473004 509498
rect 472404 473818 472586 474054
rect 472822 473818 473004 474054
rect 472404 473734 473004 473818
rect 472404 473498 472586 473734
rect 472822 473498 473004 473734
rect 472404 438054 473004 473498
rect 472404 437818 472586 438054
rect 472822 437818 473004 438054
rect 472404 437734 473004 437818
rect 472404 437498 472586 437734
rect 472822 437498 473004 437734
rect 472404 414247 473004 437498
rect 476004 549654 476604 557000
rect 476004 549418 476186 549654
rect 476422 549418 476604 549654
rect 476004 549334 476604 549418
rect 476004 549098 476186 549334
rect 476422 549098 476604 549334
rect 476004 513654 476604 549098
rect 476004 513418 476186 513654
rect 476422 513418 476604 513654
rect 476004 513334 476604 513418
rect 476004 513098 476186 513334
rect 476422 513098 476604 513334
rect 476004 477654 476604 513098
rect 476004 477418 476186 477654
rect 476422 477418 476604 477654
rect 476004 477334 476604 477418
rect 476004 477098 476186 477334
rect 476422 477098 476604 477334
rect 476004 441654 476604 477098
rect 476004 441418 476186 441654
rect 476422 441418 476604 441654
rect 476004 441334 476604 441418
rect 476004 441098 476186 441334
rect 476422 441098 476604 441334
rect 476004 414247 476604 441098
rect 479604 553254 480204 557000
rect 479604 553018 479786 553254
rect 480022 553018 480204 553254
rect 479604 552934 480204 553018
rect 479604 552698 479786 552934
rect 480022 552698 480204 552934
rect 479604 517254 480204 552698
rect 479604 517018 479786 517254
rect 480022 517018 480204 517254
rect 479604 516934 480204 517018
rect 479604 516698 479786 516934
rect 480022 516698 480204 516934
rect 479604 481254 480204 516698
rect 479604 481018 479786 481254
rect 480022 481018 480204 481254
rect 479604 480934 480204 481018
rect 479604 480698 479786 480934
rect 480022 480698 480204 480934
rect 479604 445254 480204 480698
rect 479604 445018 479786 445254
rect 480022 445018 480204 445254
rect 479604 444934 480204 445018
rect 479604 444698 479786 444934
rect 480022 444698 480204 444934
rect 479604 414247 480204 444698
rect 486804 524454 487404 557000
rect 486804 524218 486986 524454
rect 487222 524218 487404 524454
rect 486804 524134 487404 524218
rect 486804 523898 486986 524134
rect 487222 523898 487404 524134
rect 486804 488454 487404 523898
rect 486804 488218 486986 488454
rect 487222 488218 487404 488454
rect 486804 488134 487404 488218
rect 486804 487898 486986 488134
rect 487222 487898 487404 488134
rect 486804 452454 487404 487898
rect 486804 452218 486986 452454
rect 487222 452218 487404 452454
rect 486804 452134 487404 452218
rect 486804 451898 486986 452134
rect 487222 451898 487404 452134
rect 486804 416454 487404 451898
rect 486804 416218 486986 416454
rect 487222 416218 487404 416454
rect 486804 416134 487404 416218
rect 486804 415898 486986 416134
rect 487222 415898 487404 416134
rect 486804 414247 487404 415898
rect 490404 528054 491004 557000
rect 490404 527818 490586 528054
rect 490822 527818 491004 528054
rect 490404 527734 491004 527818
rect 490404 527498 490586 527734
rect 490822 527498 491004 527734
rect 490404 492054 491004 527498
rect 490404 491818 490586 492054
rect 490822 491818 491004 492054
rect 490404 491734 491004 491818
rect 490404 491498 490586 491734
rect 490822 491498 491004 491734
rect 490404 456054 491004 491498
rect 490404 455818 490586 456054
rect 490822 455818 491004 456054
rect 490404 455734 491004 455818
rect 490404 455498 490586 455734
rect 490822 455498 491004 455734
rect 490404 420054 491004 455498
rect 490404 419818 490586 420054
rect 490822 419818 491004 420054
rect 490404 419734 491004 419818
rect 490404 419498 490586 419734
rect 490822 419498 491004 419734
rect 490404 414247 491004 419498
rect 494004 531654 494604 557000
rect 494004 531418 494186 531654
rect 494422 531418 494604 531654
rect 494004 531334 494604 531418
rect 494004 531098 494186 531334
rect 494422 531098 494604 531334
rect 494004 495654 494604 531098
rect 494004 495418 494186 495654
rect 494422 495418 494604 495654
rect 494004 495334 494604 495418
rect 494004 495098 494186 495334
rect 494422 495098 494604 495334
rect 494004 459654 494604 495098
rect 494004 459418 494186 459654
rect 494422 459418 494604 459654
rect 494004 459334 494604 459418
rect 494004 459098 494186 459334
rect 494422 459098 494604 459334
rect 494004 423654 494604 459098
rect 494004 423418 494186 423654
rect 494422 423418 494604 423654
rect 494004 423334 494604 423418
rect 494004 423098 494186 423334
rect 494422 423098 494604 423334
rect 494004 414247 494604 423098
rect 497604 535254 498204 557000
rect 497604 535018 497786 535254
rect 498022 535018 498204 535254
rect 497604 534934 498204 535018
rect 497604 534698 497786 534934
rect 498022 534698 498204 534934
rect 497604 499254 498204 534698
rect 497604 499018 497786 499254
rect 498022 499018 498204 499254
rect 497604 498934 498204 499018
rect 497604 498698 497786 498934
rect 498022 498698 498204 498934
rect 497604 463254 498204 498698
rect 497604 463018 497786 463254
rect 498022 463018 498204 463254
rect 497604 462934 498204 463018
rect 497604 462698 497786 462934
rect 498022 462698 498204 462934
rect 497604 427254 498204 462698
rect 497604 427018 497786 427254
rect 498022 427018 498204 427254
rect 497604 426934 498204 427018
rect 497604 426698 497786 426934
rect 498022 426698 498204 426934
rect 497604 414247 498204 426698
rect 504804 542454 505404 557000
rect 504804 542218 504986 542454
rect 505222 542218 505404 542454
rect 504804 542134 505404 542218
rect 504804 541898 504986 542134
rect 505222 541898 505404 542134
rect 504804 506454 505404 541898
rect 504804 506218 504986 506454
rect 505222 506218 505404 506454
rect 504804 506134 505404 506218
rect 504804 505898 504986 506134
rect 505222 505898 505404 506134
rect 504804 470454 505404 505898
rect 504804 470218 504986 470454
rect 505222 470218 505404 470454
rect 504804 470134 505404 470218
rect 504804 469898 504986 470134
rect 505222 469898 505404 470134
rect 504804 434454 505404 469898
rect 504804 434218 504986 434454
rect 505222 434218 505404 434454
rect 504804 434134 505404 434218
rect 504804 433898 504986 434134
rect 505222 433898 505404 434134
rect 504804 414247 505404 433898
rect 508404 546054 509004 557000
rect 508404 545818 508586 546054
rect 508822 545818 509004 546054
rect 508404 545734 509004 545818
rect 508404 545498 508586 545734
rect 508822 545498 509004 545734
rect 508404 510054 509004 545498
rect 508404 509818 508586 510054
rect 508822 509818 509004 510054
rect 508404 509734 509004 509818
rect 508404 509498 508586 509734
rect 508822 509498 509004 509734
rect 508404 474054 509004 509498
rect 508404 473818 508586 474054
rect 508822 473818 509004 474054
rect 508404 473734 509004 473818
rect 508404 473498 508586 473734
rect 508822 473498 509004 473734
rect 508404 438054 509004 473498
rect 508404 437818 508586 438054
rect 508822 437818 509004 438054
rect 508404 437734 509004 437818
rect 508404 437498 508586 437734
rect 508822 437498 509004 437734
rect 508404 414247 509004 437498
rect 512004 549654 512604 557000
rect 512004 549418 512186 549654
rect 512422 549418 512604 549654
rect 512004 549334 512604 549418
rect 512004 549098 512186 549334
rect 512422 549098 512604 549334
rect 512004 513654 512604 549098
rect 512004 513418 512186 513654
rect 512422 513418 512604 513654
rect 512004 513334 512604 513418
rect 512004 513098 512186 513334
rect 512422 513098 512604 513334
rect 512004 477654 512604 513098
rect 512004 477418 512186 477654
rect 512422 477418 512604 477654
rect 512004 477334 512604 477418
rect 512004 477098 512186 477334
rect 512422 477098 512604 477334
rect 512004 441654 512604 477098
rect 512004 441418 512186 441654
rect 512422 441418 512604 441654
rect 512004 441334 512604 441418
rect 512004 441098 512186 441334
rect 512422 441098 512604 441334
rect 512004 414247 512604 441098
rect 515604 553254 516204 557000
rect 515604 553018 515786 553254
rect 516022 553018 516204 553254
rect 515604 552934 516204 553018
rect 515604 552698 515786 552934
rect 516022 552698 516204 552934
rect 515604 517254 516204 552698
rect 515604 517018 515786 517254
rect 516022 517018 516204 517254
rect 515604 516934 516204 517018
rect 515604 516698 515786 516934
rect 516022 516698 516204 516934
rect 515604 481254 516204 516698
rect 515604 481018 515786 481254
rect 516022 481018 516204 481254
rect 515604 480934 516204 481018
rect 515604 480698 515786 480934
rect 516022 480698 516204 480934
rect 515604 445254 516204 480698
rect 515604 445018 515786 445254
rect 516022 445018 516204 445254
rect 515604 444934 516204 445018
rect 515604 444698 515786 444934
rect 516022 444698 516204 444934
rect 515604 414247 516204 444698
rect 522804 524454 523404 559898
rect 522804 524218 522986 524454
rect 523222 524218 523404 524454
rect 522804 524134 523404 524218
rect 522804 523898 522986 524134
rect 523222 523898 523404 524134
rect 522804 488454 523404 523898
rect 522804 488218 522986 488454
rect 523222 488218 523404 488454
rect 522804 488134 523404 488218
rect 522804 487898 522986 488134
rect 523222 487898 523404 488134
rect 522804 452454 523404 487898
rect 522804 452218 522986 452454
rect 523222 452218 523404 452454
rect 522804 452134 523404 452218
rect 522804 451898 522986 452134
rect 523222 451898 523404 452134
rect 522804 416454 523404 451898
rect 522804 416218 522986 416454
rect 523222 416218 523404 416454
rect 522804 416134 523404 416218
rect 522804 415898 522986 416134
rect 523222 415898 523404 416134
rect 522804 414247 523404 415898
rect 526404 672054 527004 707102
rect 526404 671818 526586 672054
rect 526822 671818 527004 672054
rect 526404 671734 527004 671818
rect 526404 671498 526586 671734
rect 526822 671498 527004 671734
rect 526404 636054 527004 671498
rect 526404 635818 526586 636054
rect 526822 635818 527004 636054
rect 526404 635734 527004 635818
rect 526404 635498 526586 635734
rect 526822 635498 527004 635734
rect 526404 600054 527004 635498
rect 526404 599818 526586 600054
rect 526822 599818 527004 600054
rect 526404 599734 527004 599818
rect 526404 599498 526586 599734
rect 526822 599498 527004 599734
rect 526404 564054 527004 599498
rect 526404 563818 526586 564054
rect 526822 563818 527004 564054
rect 526404 563734 527004 563818
rect 526404 563498 526586 563734
rect 526822 563498 527004 563734
rect 526404 528054 527004 563498
rect 526404 527818 526586 528054
rect 526822 527818 527004 528054
rect 526404 527734 527004 527818
rect 526404 527498 526586 527734
rect 526822 527498 527004 527734
rect 526404 492054 527004 527498
rect 526404 491818 526586 492054
rect 526822 491818 527004 492054
rect 526404 491734 527004 491818
rect 526404 491498 526586 491734
rect 526822 491498 527004 491734
rect 526404 456054 527004 491498
rect 526404 455818 526586 456054
rect 526822 455818 527004 456054
rect 526404 455734 527004 455818
rect 526404 455498 526586 455734
rect 526822 455498 527004 455734
rect 526404 420054 527004 455498
rect 526404 419818 526586 420054
rect 526822 419818 527004 420054
rect 526404 419734 527004 419818
rect 526404 419498 526586 419734
rect 526822 419498 527004 419734
rect 526404 414247 527004 419498
rect 530004 675654 530604 708982
rect 530004 675418 530186 675654
rect 530422 675418 530604 675654
rect 530004 675334 530604 675418
rect 530004 675098 530186 675334
rect 530422 675098 530604 675334
rect 530004 639654 530604 675098
rect 530004 639418 530186 639654
rect 530422 639418 530604 639654
rect 530004 639334 530604 639418
rect 530004 639098 530186 639334
rect 530422 639098 530604 639334
rect 530004 603654 530604 639098
rect 530004 603418 530186 603654
rect 530422 603418 530604 603654
rect 530004 603334 530604 603418
rect 530004 603098 530186 603334
rect 530422 603098 530604 603334
rect 530004 567654 530604 603098
rect 530004 567418 530186 567654
rect 530422 567418 530604 567654
rect 530004 567334 530604 567418
rect 530004 567098 530186 567334
rect 530422 567098 530604 567334
rect 530004 531654 530604 567098
rect 530004 531418 530186 531654
rect 530422 531418 530604 531654
rect 530004 531334 530604 531418
rect 530004 531098 530186 531334
rect 530422 531098 530604 531334
rect 530004 495654 530604 531098
rect 530004 495418 530186 495654
rect 530422 495418 530604 495654
rect 530004 495334 530604 495418
rect 530004 495098 530186 495334
rect 530422 495098 530604 495334
rect 530004 459654 530604 495098
rect 530004 459418 530186 459654
rect 530422 459418 530604 459654
rect 530004 459334 530604 459418
rect 530004 459098 530186 459334
rect 530422 459098 530604 459334
rect 530004 423654 530604 459098
rect 530004 423418 530186 423654
rect 530422 423418 530604 423654
rect 530004 423334 530604 423418
rect 530004 423098 530186 423334
rect 530422 423098 530604 423334
rect 530004 414247 530604 423098
rect 533604 679254 534204 710862
rect 551604 710478 552204 711440
rect 551604 710242 551786 710478
rect 552022 710242 552204 710478
rect 551604 710158 552204 710242
rect 551604 709922 551786 710158
rect 552022 709922 552204 710158
rect 548004 708598 548604 709560
rect 548004 708362 548186 708598
rect 548422 708362 548604 708598
rect 548004 708278 548604 708362
rect 548004 708042 548186 708278
rect 548422 708042 548604 708278
rect 544404 706718 545004 707680
rect 544404 706482 544586 706718
rect 544822 706482 545004 706718
rect 544404 706398 545004 706482
rect 544404 706162 544586 706398
rect 544822 706162 545004 706398
rect 533604 679018 533786 679254
rect 534022 679018 534204 679254
rect 533604 678934 534204 679018
rect 533604 678698 533786 678934
rect 534022 678698 534204 678934
rect 533604 643254 534204 678698
rect 533604 643018 533786 643254
rect 534022 643018 534204 643254
rect 533604 642934 534204 643018
rect 533604 642698 533786 642934
rect 534022 642698 534204 642934
rect 533604 607254 534204 642698
rect 533604 607018 533786 607254
rect 534022 607018 534204 607254
rect 533604 606934 534204 607018
rect 533604 606698 533786 606934
rect 534022 606698 534204 606934
rect 533604 571254 534204 606698
rect 533604 571018 533786 571254
rect 534022 571018 534204 571254
rect 533604 570934 534204 571018
rect 533604 570698 533786 570934
rect 534022 570698 534204 570934
rect 533604 535254 534204 570698
rect 533604 535018 533786 535254
rect 534022 535018 534204 535254
rect 533604 534934 534204 535018
rect 533604 534698 533786 534934
rect 534022 534698 534204 534934
rect 533604 499254 534204 534698
rect 533604 499018 533786 499254
rect 534022 499018 534204 499254
rect 533604 498934 534204 499018
rect 533604 498698 533786 498934
rect 534022 498698 534204 498934
rect 533604 463254 534204 498698
rect 533604 463018 533786 463254
rect 534022 463018 534204 463254
rect 533604 462934 534204 463018
rect 533604 462698 533786 462934
rect 534022 462698 534204 462934
rect 533604 427254 534204 462698
rect 533604 427018 533786 427254
rect 534022 427018 534204 427254
rect 533604 426934 534204 427018
rect 533604 426698 533786 426934
rect 534022 426698 534204 426934
rect 470915 413948 470981 413949
rect 470915 413884 470916 413948
rect 470980 413884 470981 413948
rect 470915 413883 470981 413884
rect 474779 413948 474845 413949
rect 474779 413884 474780 413948
rect 474844 413884 474845 413948
rect 474779 413883 474845 413884
rect 478275 413948 478341 413949
rect 478275 413884 478276 413948
rect 478340 413884 478341 413948
rect 478275 413883 478341 413884
rect 468155 412724 468221 412725
rect 468155 412660 468156 412724
rect 468220 412660 468221 412724
rect 468155 412659 468221 412660
rect 469443 412724 469509 412725
rect 469443 412660 469444 412724
rect 469508 412660 469509 412724
rect 469443 412659 469509 412660
rect 468158 411090 468218 412659
rect 469446 411090 469506 412659
rect 470918 411090 470978 413883
rect 472019 412724 472085 412725
rect 472019 412660 472020 412724
rect 472084 412660 472085 412724
rect 472019 412659 472085 412660
rect 472022 411090 472082 412659
rect 468158 411030 468835 411090
rect 469446 411030 470083 411090
rect 470918 411030 471331 411090
rect 472022 411030 472579 411090
rect 474782 410750 474842 413883
rect 476251 413812 476317 413813
rect 476251 413748 476252 413812
rect 476316 413748 476317 413812
rect 476251 413747 476317 413748
rect 477539 413812 477605 413813
rect 477539 413748 477540 413812
rect 477604 413748 477605 413812
rect 477539 413747 477605 413748
rect 476254 411090 476314 413747
rect 476254 411030 476323 411090
rect 477542 411030 477602 413747
rect 478278 411090 478338 413883
rect 505691 413812 505757 413813
rect 505691 413748 505692 413812
rect 505756 413748 505757 413812
rect 505691 413747 505757 413748
rect 479379 413676 479445 413677
rect 479379 413612 479380 413676
rect 479444 413612 479445 413676
rect 479379 413611 479445 413612
rect 479382 411090 479442 413611
rect 480667 413540 480733 413541
rect 480667 413476 480668 413540
rect 480732 413476 480733 413540
rect 480667 413475 480733 413476
rect 485819 413540 485885 413541
rect 485819 413476 485820 413540
rect 485884 413476 485885 413540
rect 485819 413475 485885 413476
rect 480670 411090 480730 413475
rect 481955 413404 482021 413405
rect 481955 413340 481956 413404
rect 482020 413340 482021 413404
rect 481955 413339 482021 413340
rect 483427 413404 483493 413405
rect 483427 413340 483428 413404
rect 483492 413340 483493 413404
rect 483427 413339 483493 413340
rect 481958 411090 482018 413339
rect 483430 411090 483490 413339
rect 484531 413268 484597 413269
rect 484531 413204 484532 413268
rect 484596 413204 484597 413268
rect 484531 413203 484597 413204
rect 484534 411090 484594 413203
rect 485822 411090 485882 413475
rect 488579 413268 488645 413269
rect 488579 413204 488580 413268
rect 488644 413204 488645 413268
rect 488579 413203 488645 413204
rect 487291 413132 487357 413133
rect 487291 413068 487292 413132
rect 487356 413068 487357 413132
rect 487291 413067 487357 413068
rect 487294 411090 487354 413067
rect 488582 411090 488642 413203
rect 490051 412996 490117 412997
rect 490051 412932 490052 412996
rect 490116 412932 490117 412996
rect 490051 412931 490117 412932
rect 491339 412996 491405 412997
rect 491339 412932 491340 412996
rect 491404 412932 491405 412996
rect 491339 412931 491405 412932
rect 490054 411090 490114 412931
rect 491342 411770 491402 412931
rect 491891 412724 491957 412725
rect 491891 412660 491892 412724
rect 491956 412660 491957 412724
rect 491891 412659 491957 412660
rect 493179 412724 493245 412725
rect 493179 412660 493180 412724
rect 493244 412660 493245 412724
rect 493179 412659 493245 412660
rect 494467 412724 494533 412725
rect 494467 412660 494468 412724
rect 494532 412660 494533 412724
rect 494467 412659 494533 412660
rect 495755 412724 495821 412725
rect 495755 412660 495756 412724
rect 495820 412660 495821 412724
rect 495755 412659 495821 412660
rect 496859 412724 496925 412725
rect 496859 412660 496860 412724
rect 496924 412660 496925 412724
rect 496859 412659 496925 412660
rect 498331 412724 498397 412725
rect 498331 412660 498332 412724
rect 498396 412660 498397 412724
rect 498331 412659 498397 412660
rect 499619 412724 499685 412725
rect 499619 412660 499620 412724
rect 499684 412660 499685 412724
rect 499619 412659 499685 412660
rect 501091 412724 501157 412725
rect 501091 412660 501092 412724
rect 501156 412660 501157 412724
rect 501091 412659 501157 412660
rect 502747 412724 502813 412725
rect 502747 412660 502748 412724
rect 502812 412660 502813 412724
rect 502747 412659 502813 412660
rect 503667 412724 503733 412725
rect 503667 412660 503668 412724
rect 503732 412660 503733 412724
rect 503667 412659 503733 412660
rect 504403 412724 504469 412725
rect 504403 412660 504404 412724
rect 504468 412660 504469 412724
rect 504403 412659 504469 412660
rect 478278 411030 478819 411090
rect 479382 411030 480067 411090
rect 480670 411030 481315 411090
rect 481958 411030 482563 411090
rect 483430 411030 483811 411090
rect 484534 411030 485059 411090
rect 485822 411030 486307 411090
rect 487294 411030 487555 411090
rect 488582 411030 488803 411090
rect 490051 411030 490114 411090
rect 491269 411710 491402 411770
rect 491269 411060 491329 411710
rect 491894 411090 491954 412659
rect 493182 411090 493242 412659
rect 494470 411090 494530 412659
rect 495758 411090 495818 412659
rect 496862 411090 496922 412659
rect 498334 411090 498394 412659
rect 499622 411090 499682 412659
rect 501094 411090 501154 412659
rect 491894 411030 492547 411090
rect 493182 411030 493795 411090
rect 494470 411030 495043 411090
rect 495758 411030 496291 411090
rect 496862 411030 497539 411090
rect 498334 411030 498787 411090
rect 499622 411030 500035 411090
rect 501094 411030 501283 411090
rect 502750 410750 502810 412659
rect 503670 411770 503730 412659
rect 503670 411710 503809 411770
rect 503749 411060 503809 411710
rect 504406 411090 504466 412659
rect 505694 411090 505754 413747
rect 506979 413676 507045 413677
rect 506979 413612 506980 413676
rect 507044 413612 507045 413676
rect 506979 413611 507045 413612
rect 506982 411090 507042 413611
rect 522987 412860 523053 412861
rect 522987 412796 522988 412860
rect 523052 412796 523053 412860
rect 522987 412795 523053 412796
rect 518019 412724 518085 412725
rect 518019 412660 518020 412724
rect 518084 412660 518085 412724
rect 518019 412659 518085 412660
rect 518022 411090 518082 412659
rect 522990 411090 523050 412795
rect 504406 411030 505027 411090
rect 505694 411030 506275 411090
rect 506982 411030 507523 411090
rect 518022 411030 518608 411090
rect 522990 411030 523603 411090
rect 474782 410690 475075 410750
rect 502531 410690 502810 410750
rect 473445 410412 473511 410413
rect 473445 410348 473446 410412
rect 473510 410410 473511 410412
rect 473510 410350 473827 410410
rect 473510 410348 473511 410350
rect 473445 410347 473511 410348
rect 443604 409018 443786 409254
rect 444022 409018 444204 409254
rect 443604 408934 444204 409018
rect 443604 408698 443786 408934
rect 444022 408698 444204 408934
rect 443604 373254 444204 408698
rect 526494 405654 526814 405676
rect 526494 405418 526536 405654
rect 526772 405418 526814 405654
rect 526494 405334 526814 405418
rect 526494 405098 526536 405334
rect 526772 405098 526814 405334
rect 526494 405076 526814 405098
rect 526494 402054 526814 402076
rect 526494 401818 526536 402054
rect 526772 401818 526814 402054
rect 526494 401734 526814 401818
rect 526494 401498 526536 401734
rect 526772 401498 526814 401734
rect 526494 401476 526814 401498
rect 526494 398454 526814 398476
rect 526494 398218 526536 398454
rect 526772 398218 526814 398454
rect 526494 398134 526814 398218
rect 526494 397898 526536 398134
rect 526772 397898 526814 398134
rect 526494 397876 526814 397898
rect 526938 391254 527262 391276
rect 526938 391018 526982 391254
rect 527218 391018 527262 391254
rect 526938 390934 527262 391018
rect 526938 390698 526982 390934
rect 527218 390698 527262 390934
rect 526938 390676 527262 390698
rect 533604 391254 534204 426698
rect 533604 391018 533786 391254
rect 534022 391018 534204 391254
rect 533604 390934 534204 391018
rect 533604 390698 533786 390934
rect 534022 390698 534204 390934
rect 526938 387654 527262 387676
rect 526938 387418 526982 387654
rect 527218 387418 527262 387654
rect 526938 387334 527262 387418
rect 526938 387098 526982 387334
rect 527218 387098 527262 387334
rect 526938 387076 527262 387098
rect 526938 384054 527262 384076
rect 526938 383818 526982 384054
rect 527218 383818 527262 384054
rect 526938 383734 527262 383818
rect 526938 383498 526982 383734
rect 527218 383498 527262 383734
rect 526938 383476 527262 383498
rect 526938 380454 527262 380476
rect 526938 380218 526982 380454
rect 527218 380218 527262 380454
rect 526938 380134 527262 380218
rect 526938 379898 526982 380134
rect 527218 379898 527262 380134
rect 526938 379876 527262 379898
rect 443604 373018 443786 373254
rect 444022 373018 444204 373254
rect 443604 372934 444204 373018
rect 443604 372698 443786 372934
rect 444022 372698 444204 372934
rect 443604 337254 444204 372698
rect 526494 373254 526814 373276
rect 526494 373018 526536 373254
rect 526772 373018 526814 373254
rect 526494 372934 526814 373018
rect 526494 372698 526536 372934
rect 526772 372698 526814 372934
rect 526494 372676 526814 372698
rect 526494 369654 526814 369676
rect 526494 369418 526536 369654
rect 526772 369418 526814 369654
rect 526494 369334 526814 369418
rect 526494 369098 526536 369334
rect 526772 369098 526814 369334
rect 526494 369076 526814 369098
rect 526494 366054 526814 366076
rect 526494 365818 526536 366054
rect 526772 365818 526814 366054
rect 526494 365734 526814 365818
rect 526494 365498 526536 365734
rect 526772 365498 526814 365734
rect 526494 365476 526814 365498
rect 526494 362454 526814 362476
rect 526494 362218 526536 362454
rect 526772 362218 526814 362454
rect 526494 362134 526814 362218
rect 526494 361898 526536 362134
rect 526772 361898 526814 362134
rect 526494 361876 526814 361898
rect 526938 355254 527262 355276
rect 526938 355018 526982 355254
rect 527218 355018 527262 355254
rect 526938 354934 527262 355018
rect 526938 354698 526982 354934
rect 527218 354698 527262 354934
rect 526938 354676 527262 354698
rect 533604 355254 534204 390698
rect 533604 355018 533786 355254
rect 534022 355018 534204 355254
rect 533604 354934 534204 355018
rect 533604 354698 533786 354934
rect 534022 354698 534204 354934
rect 526938 351654 527262 351676
rect 526938 351418 526982 351654
rect 527218 351418 527262 351654
rect 526938 351334 527262 351418
rect 526938 351098 526982 351334
rect 527218 351098 527262 351334
rect 526938 351076 527262 351098
rect 526938 348054 527262 348076
rect 526938 347818 526982 348054
rect 527218 347818 527262 348054
rect 526938 347734 527262 347818
rect 526938 347498 526982 347734
rect 527218 347498 527262 347734
rect 526938 347476 527262 347498
rect 527955 347172 528021 347173
rect 527955 347108 527956 347172
rect 528020 347108 528021 347172
rect 527955 347107 528021 347108
rect 527958 346578 528018 347107
rect 527587 346492 527653 346493
rect 527587 346428 527588 346492
rect 527652 346428 527653 346492
rect 527587 346427 527653 346428
rect 527590 345898 527650 346427
rect 527590 344917 527650 344982
rect 527587 344916 527653 344917
rect 527587 344852 527588 344916
rect 527652 344852 527653 344916
rect 527587 344851 527653 344852
rect 526938 344454 527262 344476
rect 526938 344218 526982 344454
rect 527218 344218 527262 344454
rect 526938 344134 527262 344218
rect 526938 343898 526982 344134
rect 527218 343898 527262 344134
rect 526938 343876 527262 343898
rect 527955 343228 528021 343229
rect 450675 343092 450741 343093
rect 450675 343028 450676 343092
rect 450740 343028 450741 343092
rect 450675 343027 450741 343028
rect 444570 341670 445070 341730
rect 445526 340373 445586 342262
rect 445523 340372 445589 340373
rect 445523 340308 445524 340372
rect 445588 340308 445589 340372
rect 445523 340307 445589 340308
rect 450678 338418 450738 343027
rect 527955 343164 527956 343228
rect 528020 343164 528021 343228
rect 527955 343163 528021 343164
rect 527590 342005 527650 342942
rect 527587 342004 527653 342005
rect 527587 341940 527588 342004
rect 527652 341940 527653 342004
rect 527587 341939 527653 341940
rect 527958 340458 528018 343163
rect 443604 337018 443786 337254
rect 444022 337018 444204 337254
rect 443604 336934 444204 337018
rect 443604 336698 443786 336934
rect 444022 336698 444204 336934
rect 443604 303000 444204 336698
rect 526494 337254 526814 337276
rect 526494 337018 526536 337254
rect 526772 337018 526814 337254
rect 526494 336934 526814 337018
rect 526494 336698 526536 336934
rect 526772 336698 526814 336934
rect 526494 336676 526814 336698
rect 526494 333654 526814 333676
rect 526494 333418 526536 333654
rect 526772 333418 526814 333654
rect 526494 333334 526814 333418
rect 526494 333098 526536 333334
rect 526772 333098 526814 333334
rect 526494 333076 526814 333098
rect 526494 330054 526814 330076
rect 526494 329818 526536 330054
rect 526772 329818 526814 330054
rect 526494 329734 526814 329818
rect 526494 329498 526536 329734
rect 526772 329498 526814 329734
rect 526494 329476 526814 329498
rect 526494 326454 526814 326476
rect 526494 326218 526536 326454
rect 526772 326218 526814 326454
rect 526494 326134 526814 326218
rect 526494 325898 526536 326134
rect 526772 325898 526814 326134
rect 526494 325876 526814 325898
rect 453254 320250 453833 320310
rect 453254 318749 453314 320250
rect 533604 319254 534204 354698
rect 533604 319018 533786 319254
rect 534022 319018 534204 319254
rect 533604 318934 534204 319018
rect 453251 318748 453317 318749
rect 453251 318684 453252 318748
rect 453316 318684 453317 318748
rect 453251 318683 453317 318684
rect 533604 318698 533786 318934
rect 534022 318698 534204 318934
rect 450804 308454 451404 317000
rect 450804 308218 450986 308454
rect 451222 308218 451404 308454
rect 450804 308134 451404 308218
rect 450804 307898 450986 308134
rect 451222 307898 451404 308134
rect 450804 303000 451404 307898
rect 454404 312054 455004 317000
rect 454404 311818 454586 312054
rect 454822 311818 455004 312054
rect 454404 311734 455004 311818
rect 454404 311498 454586 311734
rect 454822 311498 455004 311734
rect 454404 303000 455004 311498
rect 458004 315654 458604 317000
rect 458004 315418 458186 315654
rect 458422 315418 458604 315654
rect 458004 315334 458604 315418
rect 458004 315098 458186 315334
rect 458422 315098 458604 315334
rect 458004 303000 458604 315098
rect 461604 303000 462204 317000
rect 468804 303000 469404 317000
rect 472404 303000 473004 317000
rect 476004 303000 476604 317000
rect 479604 303000 480204 317000
rect 486804 308454 487404 317000
rect 486804 308218 486986 308454
rect 487222 308218 487404 308454
rect 486804 308134 487404 308218
rect 486804 307898 486986 308134
rect 487222 307898 487404 308134
rect 486804 303000 487404 307898
rect 490404 312054 491004 317000
rect 490404 311818 490586 312054
rect 490822 311818 491004 312054
rect 490404 311734 491004 311818
rect 490404 311498 490586 311734
rect 490822 311498 491004 311734
rect 490404 303000 491004 311498
rect 494004 315654 494604 317000
rect 494004 315418 494186 315654
rect 494422 315418 494604 315654
rect 494004 315334 494604 315418
rect 494004 315098 494186 315334
rect 494422 315098 494604 315334
rect 494004 303000 494604 315098
rect 497604 303000 498204 317000
rect 504804 303000 505404 317000
rect 508404 303000 509004 317000
rect 512004 303000 512604 317000
rect 515604 303000 516204 317000
rect 522804 308454 523404 317000
rect 522804 308218 522986 308454
rect 523222 308218 523404 308454
rect 522804 308134 523404 308218
rect 522804 307898 522986 308134
rect 523222 307898 523404 308134
rect 522804 303000 523404 307898
rect 526404 312054 527004 317000
rect 526404 311818 526586 312054
rect 526822 311818 527004 312054
rect 526404 311734 527004 311818
rect 526404 311498 526586 311734
rect 526822 311498 527004 311734
rect 526404 303000 527004 311498
rect 530004 315654 530604 317000
rect 530004 315418 530186 315654
rect 530422 315418 530604 315654
rect 530004 315334 530604 315418
rect 530004 315098 530186 315334
rect 530422 315098 530604 315334
rect 530004 303000 530604 315098
rect 299604 301018 299786 301254
rect 300022 301018 300204 301254
rect 299604 300934 300204 301018
rect 299604 300698 299786 300934
rect 300022 300698 300204 300934
rect 299604 265254 300204 300698
rect 314208 294054 314528 294076
rect 314208 293818 314250 294054
rect 314486 293818 314528 294054
rect 314208 293734 314528 293818
rect 314208 293498 314250 293734
rect 314486 293498 314528 293734
rect 314208 293476 314528 293498
rect 314208 290454 314528 290476
rect 314208 290218 314250 290454
rect 314486 290218 314528 290454
rect 314208 290134 314528 290218
rect 314208 289898 314250 290134
rect 314486 289898 314528 290134
rect 314208 289876 314528 289898
rect 329568 283254 329888 283276
rect 329568 283018 329610 283254
rect 329846 283018 329888 283254
rect 329568 282934 329888 283018
rect 329568 282698 329610 282934
rect 329846 282698 329888 282934
rect 329568 282676 329888 282698
rect 533604 283254 534204 318698
rect 533604 283018 533786 283254
rect 534022 283018 534204 283254
rect 533604 282934 534204 283018
rect 533604 282698 533786 282934
rect 534022 282698 534204 282934
rect 329568 279654 329888 279676
rect 329568 279418 329610 279654
rect 329846 279418 329888 279654
rect 329568 279334 329888 279418
rect 329568 279098 329610 279334
rect 329846 279098 329888 279334
rect 329568 279076 329888 279098
rect 329568 276054 329888 276076
rect 329568 275818 329610 276054
rect 329846 275818 329888 276054
rect 329568 275734 329888 275818
rect 329568 275498 329610 275734
rect 329846 275498 329888 275734
rect 329568 275476 329888 275498
rect 329568 272454 329888 272476
rect 329568 272218 329610 272454
rect 329846 272218 329888 272454
rect 329568 272134 329888 272218
rect 329568 271898 329610 272134
rect 329846 271898 329888 272134
rect 329568 271876 329888 271898
rect 299604 265018 299786 265254
rect 300022 265018 300204 265254
rect 299604 264934 300204 265018
rect 299604 264698 299786 264934
rect 300022 264698 300204 264934
rect 299604 229254 300204 264698
rect 314208 265254 314528 265276
rect 314208 265018 314250 265254
rect 314486 265018 314528 265254
rect 314208 264934 314528 265018
rect 314208 264698 314250 264934
rect 314486 264698 314528 264934
rect 314208 264676 314528 264698
rect 314208 261654 314528 261676
rect 314208 261418 314250 261654
rect 314486 261418 314528 261654
rect 314208 261334 314528 261418
rect 314208 261098 314250 261334
rect 314486 261098 314528 261334
rect 314208 261076 314528 261098
rect 314208 258054 314528 258076
rect 314208 257818 314250 258054
rect 314486 257818 314528 258054
rect 314208 257734 314528 257818
rect 314208 257498 314250 257734
rect 314486 257498 314528 257734
rect 314208 257476 314528 257498
rect 314208 254454 314528 254476
rect 314208 254218 314250 254454
rect 314486 254218 314528 254454
rect 314208 254134 314528 254218
rect 314208 253898 314250 254134
rect 314486 253898 314528 254134
rect 314208 253876 314528 253898
rect 329568 247254 329888 247276
rect 329568 247018 329610 247254
rect 329846 247018 329888 247254
rect 329568 246934 329888 247018
rect 329568 246698 329610 246934
rect 329846 246698 329888 246934
rect 329568 246676 329888 246698
rect 533604 247254 534204 282698
rect 533604 247018 533786 247254
rect 534022 247018 534204 247254
rect 533604 246934 534204 247018
rect 533604 246698 533786 246934
rect 534022 246698 534204 246934
rect 329568 243654 329888 243676
rect 329568 243418 329610 243654
rect 329846 243418 329888 243654
rect 329568 243334 329888 243418
rect 329568 243098 329610 243334
rect 329846 243098 329888 243334
rect 329568 243076 329888 243098
rect 329568 240054 329888 240076
rect 329568 239818 329610 240054
rect 329846 239818 329888 240054
rect 329568 239734 329888 239818
rect 329568 239498 329610 239734
rect 329846 239498 329888 239734
rect 329568 239476 329888 239498
rect 329568 236454 329888 236476
rect 329568 236218 329610 236454
rect 329846 236218 329888 236454
rect 329568 236134 329888 236218
rect 329568 235898 329610 236134
rect 329846 235898 329888 236134
rect 329568 235876 329888 235898
rect 299604 229018 299786 229254
rect 300022 229018 300204 229254
rect 299604 228934 300204 229018
rect 299604 228698 299786 228934
rect 300022 228698 300204 228934
rect 299604 193254 300204 228698
rect 314208 229254 314528 229276
rect 314208 229018 314250 229254
rect 314486 229018 314528 229254
rect 314208 228934 314528 229018
rect 314208 228698 314250 228934
rect 314486 228698 314528 228934
rect 314208 228676 314528 228698
rect 314208 225654 314528 225676
rect 314208 225418 314250 225654
rect 314486 225418 314528 225654
rect 314208 225334 314528 225418
rect 314208 225098 314250 225334
rect 314486 225098 314528 225334
rect 314208 225076 314528 225098
rect 314208 222054 314528 222076
rect 314208 221818 314250 222054
rect 314486 221818 314528 222054
rect 314208 221734 314528 221818
rect 314208 221498 314250 221734
rect 314486 221498 314528 221734
rect 314208 221476 314528 221498
rect 314208 218454 314528 218476
rect 314208 218218 314250 218454
rect 314486 218218 314528 218454
rect 314208 218134 314528 218218
rect 314208 217898 314250 218134
rect 314486 217898 314528 218134
rect 314208 217876 314528 217898
rect 329568 211254 329888 211276
rect 329568 211018 329610 211254
rect 329846 211018 329888 211254
rect 329568 210934 329888 211018
rect 329568 210698 329610 210934
rect 329846 210698 329888 210934
rect 329568 210676 329888 210698
rect 533604 211254 534204 246698
rect 533604 211018 533786 211254
rect 534022 211018 534204 211254
rect 533604 210934 534204 211018
rect 533604 210698 533786 210934
rect 534022 210698 534204 210934
rect 329568 207654 329888 207676
rect 329568 207418 329610 207654
rect 329846 207418 329888 207654
rect 329568 207334 329888 207418
rect 329568 207098 329610 207334
rect 329846 207098 329888 207334
rect 329568 207076 329888 207098
rect 329568 204054 329888 204076
rect 329568 203818 329610 204054
rect 329846 203818 329888 204054
rect 329568 203734 329888 203818
rect 329568 203498 329610 203734
rect 329846 203498 329888 203734
rect 329568 203476 329888 203498
rect 329568 200454 329888 200476
rect 329568 200218 329610 200454
rect 329846 200218 329888 200454
rect 329568 200134 329888 200218
rect 329568 199898 329610 200134
rect 329846 199898 329888 200134
rect 329568 199876 329888 199898
rect 299604 193018 299786 193254
rect 300022 193018 300204 193254
rect 299604 192934 300204 193018
rect 299604 192698 299786 192934
rect 300022 192698 300204 192934
rect 299604 157254 300204 192698
rect 314208 193254 314528 193276
rect 314208 193018 314250 193254
rect 314486 193018 314528 193254
rect 314208 192934 314528 193018
rect 314208 192698 314250 192934
rect 314486 192698 314528 192934
rect 314208 192676 314528 192698
rect 314208 189654 314528 189676
rect 314208 189418 314250 189654
rect 314486 189418 314528 189654
rect 314208 189334 314528 189418
rect 314208 189098 314250 189334
rect 314486 189098 314528 189334
rect 314208 189076 314528 189098
rect 314208 186054 314528 186076
rect 314208 185818 314250 186054
rect 314486 185818 314528 186054
rect 314208 185734 314528 185818
rect 314208 185498 314250 185734
rect 314486 185498 314528 185734
rect 314208 185476 314528 185498
rect 314208 182454 314528 182476
rect 314208 182218 314250 182454
rect 314486 182218 314528 182454
rect 314208 182134 314528 182218
rect 314208 181898 314250 182134
rect 314486 181898 314528 182134
rect 314208 181876 314528 181898
rect 329568 175254 329888 175276
rect 329568 175018 329610 175254
rect 329846 175018 329888 175254
rect 329568 174934 329888 175018
rect 329568 174698 329610 174934
rect 329846 174698 329888 174934
rect 329568 174676 329888 174698
rect 533604 175254 534204 210698
rect 533604 175018 533786 175254
rect 534022 175018 534204 175254
rect 533604 174934 534204 175018
rect 533604 174698 533786 174934
rect 534022 174698 534204 174934
rect 329568 171654 329888 171676
rect 329568 171418 329610 171654
rect 329846 171418 329888 171654
rect 329568 171334 329888 171418
rect 329568 171098 329610 171334
rect 329846 171098 329888 171334
rect 329568 171076 329888 171098
rect 329568 168054 329888 168076
rect 329568 167818 329610 168054
rect 329846 167818 329888 168054
rect 329568 167734 329888 167818
rect 329568 167498 329610 167734
rect 329846 167498 329888 167734
rect 329568 167476 329888 167498
rect 329568 164454 329888 164476
rect 329568 164218 329610 164454
rect 329846 164218 329888 164454
rect 329568 164134 329888 164218
rect 329568 163898 329610 164134
rect 329846 163898 329888 164134
rect 329568 163876 329888 163898
rect 299604 157018 299786 157254
rect 300022 157018 300204 157254
rect 299604 156934 300204 157018
rect 299604 156698 299786 156934
rect 300022 156698 300204 156934
rect 299604 121254 300204 156698
rect 314208 157254 314528 157276
rect 314208 157018 314250 157254
rect 314486 157018 314528 157254
rect 314208 156934 314528 157018
rect 314208 156698 314250 156934
rect 314486 156698 314528 156934
rect 314208 156676 314528 156698
rect 314208 153654 314528 153676
rect 314208 153418 314250 153654
rect 314486 153418 314528 153654
rect 314208 153334 314528 153418
rect 314208 153098 314250 153334
rect 314486 153098 314528 153334
rect 314208 153076 314528 153098
rect 314208 150054 314528 150076
rect 314208 149818 314250 150054
rect 314486 149818 314528 150054
rect 314208 149734 314528 149818
rect 314208 149498 314250 149734
rect 314486 149498 314528 149734
rect 314208 149476 314528 149498
rect 314208 146454 314528 146476
rect 314208 146218 314250 146454
rect 314486 146218 314528 146454
rect 314208 146134 314528 146218
rect 314208 145898 314250 146134
rect 314486 145898 314528 146134
rect 314208 145876 314528 145898
rect 329568 139254 329888 139276
rect 329568 139018 329610 139254
rect 329846 139018 329888 139254
rect 329568 138934 329888 139018
rect 329568 138698 329610 138934
rect 329846 138698 329888 138934
rect 329568 138676 329888 138698
rect 533604 139254 534204 174698
rect 533604 139018 533786 139254
rect 534022 139018 534204 139254
rect 533604 138934 534204 139018
rect 533604 138698 533786 138934
rect 534022 138698 534204 138934
rect 329568 135654 329888 135676
rect 329568 135418 329610 135654
rect 329846 135418 329888 135654
rect 329568 135334 329888 135418
rect 329568 135098 329610 135334
rect 329846 135098 329888 135334
rect 329568 135076 329888 135098
rect 329568 132054 329888 132076
rect 329568 131818 329610 132054
rect 329846 131818 329888 132054
rect 329568 131734 329888 131818
rect 329568 131498 329610 131734
rect 329846 131498 329888 131734
rect 329568 131476 329888 131498
rect 329568 128454 329888 128476
rect 329568 128218 329610 128454
rect 329846 128218 329888 128454
rect 329568 128134 329888 128218
rect 329568 127898 329610 128134
rect 329846 127898 329888 128134
rect 329568 127876 329888 127898
rect 299604 121018 299786 121254
rect 300022 121018 300204 121254
rect 299604 120934 300204 121018
rect 299604 120698 299786 120934
rect 300022 120698 300204 120934
rect 299604 85254 300204 120698
rect 314208 121254 314528 121276
rect 314208 121018 314250 121254
rect 314486 121018 314528 121254
rect 314208 120934 314528 121018
rect 314208 120698 314250 120934
rect 314486 120698 314528 120934
rect 314208 120676 314528 120698
rect 314208 117654 314528 117676
rect 314208 117418 314250 117654
rect 314486 117418 314528 117654
rect 314208 117334 314528 117418
rect 314208 117098 314250 117334
rect 314486 117098 314528 117334
rect 314208 117076 314528 117098
rect 314208 114054 314528 114076
rect 314208 113818 314250 114054
rect 314486 113818 314528 114054
rect 314208 113734 314528 113818
rect 314208 113498 314250 113734
rect 314486 113498 314528 113734
rect 314208 113476 314528 113498
rect 314208 110454 314528 110476
rect 314208 110218 314250 110454
rect 314486 110218 314528 110454
rect 314208 110134 314528 110218
rect 314208 109898 314250 110134
rect 314486 109898 314528 110134
rect 314208 109876 314528 109898
rect 329568 103254 329888 103276
rect 329568 103018 329610 103254
rect 329846 103018 329888 103254
rect 329568 102934 329888 103018
rect 329568 102698 329610 102934
rect 329846 102698 329888 102934
rect 329568 102676 329888 102698
rect 533604 103254 534204 138698
rect 533604 103018 533786 103254
rect 534022 103018 534204 103254
rect 533604 102934 534204 103018
rect 533604 102698 533786 102934
rect 534022 102698 534204 102934
rect 329568 99654 329888 99676
rect 329568 99418 329610 99654
rect 329846 99418 329888 99654
rect 329568 99334 329888 99418
rect 329568 99098 329610 99334
rect 329846 99098 329888 99334
rect 329568 99076 329888 99098
rect 329568 96054 329888 96076
rect 329568 95818 329610 96054
rect 329846 95818 329888 96054
rect 329568 95734 329888 95818
rect 329568 95498 329610 95734
rect 329846 95498 329888 95734
rect 329568 95476 329888 95498
rect 329568 92454 329888 92476
rect 329568 92218 329610 92454
rect 329846 92218 329888 92454
rect 329568 92134 329888 92218
rect 329568 91898 329610 92134
rect 329846 91898 329888 92134
rect 329568 91876 329888 91898
rect 299604 85018 299786 85254
rect 300022 85018 300204 85254
rect 299604 84934 300204 85018
rect 299604 84698 299786 84934
rect 300022 84698 300204 84934
rect 299604 49254 300204 84698
rect 314208 85254 314528 85276
rect 314208 85018 314250 85254
rect 314486 85018 314528 85254
rect 314208 84934 314528 85018
rect 314208 84698 314250 84934
rect 314486 84698 314528 84934
rect 314208 84676 314528 84698
rect 299604 49018 299786 49254
rect 300022 49018 300204 49254
rect 299604 48934 300204 49018
rect 299604 48698 299786 48934
rect 300022 48698 300204 48934
rect 299604 13254 300204 48698
rect 299604 13018 299786 13254
rect 300022 13018 300204 13254
rect 299604 12934 300204 13018
rect 299604 12698 299786 12934
rect 300022 12698 300204 12934
rect 281604 -7162 281786 -6926
rect 282022 -7162 282204 -6926
rect 281604 -7246 282204 -7162
rect 281604 -7482 281786 -7246
rect 282022 -7482 282204 -7246
rect 281604 -7504 282204 -7482
rect 299604 -5986 300204 12698
rect 306804 56454 307404 77000
rect 306804 56218 306986 56454
rect 307222 56218 307404 56454
rect 306804 56134 307404 56218
rect 306804 55898 306986 56134
rect 307222 55898 307404 56134
rect 306804 20454 307404 55898
rect 306804 20218 306986 20454
rect 307222 20218 307404 20454
rect 306804 20134 307404 20218
rect 306804 19898 306986 20134
rect 307222 19898 307404 20134
rect 306804 -1286 307404 19898
rect 306804 -1522 306986 -1286
rect 307222 -1522 307404 -1286
rect 306804 -1606 307404 -1522
rect 306804 -1842 306986 -1606
rect 307222 -1842 307404 -1606
rect 306804 -1864 307404 -1842
rect 310404 60054 311004 77000
rect 310404 59818 310586 60054
rect 310822 59818 311004 60054
rect 310404 59734 311004 59818
rect 310404 59498 310586 59734
rect 310822 59498 311004 59734
rect 310404 24054 311004 59498
rect 310404 23818 310586 24054
rect 310822 23818 311004 24054
rect 310404 23734 311004 23818
rect 310404 23498 310586 23734
rect 310822 23498 311004 23734
rect 310404 -3166 311004 23498
rect 310404 -3402 310586 -3166
rect 310822 -3402 311004 -3166
rect 310404 -3486 311004 -3402
rect 310404 -3722 310586 -3486
rect 310822 -3722 311004 -3486
rect 310404 -3744 311004 -3722
rect 314004 63654 314604 77000
rect 314004 63418 314186 63654
rect 314422 63418 314604 63654
rect 314004 63334 314604 63418
rect 314004 63098 314186 63334
rect 314422 63098 314604 63334
rect 314004 27654 314604 63098
rect 314004 27418 314186 27654
rect 314422 27418 314604 27654
rect 314004 27334 314604 27418
rect 314004 27098 314186 27334
rect 314422 27098 314604 27334
rect 314004 -5046 314604 27098
rect 314004 -5282 314186 -5046
rect 314422 -5282 314604 -5046
rect 314004 -5366 314604 -5282
rect 314004 -5602 314186 -5366
rect 314422 -5602 314604 -5366
rect 314004 -5624 314604 -5602
rect 317604 67254 318204 77000
rect 317604 67018 317786 67254
rect 318022 67018 318204 67254
rect 317604 66934 318204 67018
rect 317604 66698 317786 66934
rect 318022 66698 318204 66934
rect 317604 31254 318204 66698
rect 317604 31018 317786 31254
rect 318022 31018 318204 31254
rect 317604 30934 318204 31018
rect 317604 30698 317786 30934
rect 318022 30698 318204 30934
rect 299604 -6222 299786 -5986
rect 300022 -6222 300204 -5986
rect 299604 -6306 300204 -6222
rect 299604 -6542 299786 -6306
rect 300022 -6542 300204 -6306
rect 299604 -7504 300204 -6542
rect 317604 -6926 318204 30698
rect 324804 74454 325404 77000
rect 324804 74218 324986 74454
rect 325222 74218 325404 74454
rect 324804 74134 325404 74218
rect 324804 73898 324986 74134
rect 325222 73898 325404 74134
rect 324804 38454 325404 73898
rect 324804 38218 324986 38454
rect 325222 38218 325404 38454
rect 324804 38134 325404 38218
rect 324804 37898 324986 38134
rect 325222 37898 325404 38134
rect 324804 2454 325404 37898
rect 324804 2218 324986 2454
rect 325222 2218 325404 2454
rect 324804 2134 325404 2218
rect 324804 1898 324986 2134
rect 325222 1898 325404 2134
rect 324804 -346 325404 1898
rect 324804 -582 324986 -346
rect 325222 -582 325404 -346
rect 324804 -666 325404 -582
rect 324804 -902 324986 -666
rect 325222 -902 325404 -666
rect 324804 -1864 325404 -902
rect 328404 42054 329004 77000
rect 328404 41818 328586 42054
rect 328822 41818 329004 42054
rect 328404 41734 329004 41818
rect 328404 41498 328586 41734
rect 328822 41498 329004 41734
rect 328404 6054 329004 41498
rect 328404 5818 328586 6054
rect 328822 5818 329004 6054
rect 328404 5734 329004 5818
rect 328404 5498 328586 5734
rect 328822 5498 329004 5734
rect 328404 -2226 329004 5498
rect 328404 -2462 328586 -2226
rect 328822 -2462 329004 -2226
rect 328404 -2546 329004 -2462
rect 328404 -2782 328586 -2546
rect 328822 -2782 329004 -2546
rect 328404 -3744 329004 -2782
rect 332004 45654 332604 77000
rect 332004 45418 332186 45654
rect 332422 45418 332604 45654
rect 332004 45334 332604 45418
rect 332004 45098 332186 45334
rect 332422 45098 332604 45334
rect 332004 9654 332604 45098
rect 332004 9418 332186 9654
rect 332422 9418 332604 9654
rect 332004 9334 332604 9418
rect 332004 9098 332186 9334
rect 332422 9098 332604 9334
rect 332004 -4106 332604 9098
rect 332004 -4342 332186 -4106
rect 332422 -4342 332604 -4106
rect 332004 -4426 332604 -4342
rect 332004 -4662 332186 -4426
rect 332422 -4662 332604 -4426
rect 332004 -5624 332604 -4662
rect 335604 49254 336204 77000
rect 335604 49018 335786 49254
rect 336022 49018 336204 49254
rect 335604 48934 336204 49018
rect 335604 48698 335786 48934
rect 336022 48698 336204 48934
rect 335604 13254 336204 48698
rect 335604 13018 335786 13254
rect 336022 13018 336204 13254
rect 335604 12934 336204 13018
rect 335604 12698 335786 12934
rect 336022 12698 336204 12934
rect 317604 -7162 317786 -6926
rect 318022 -7162 318204 -6926
rect 317604 -7246 318204 -7162
rect 317604 -7482 317786 -7246
rect 318022 -7482 318204 -7246
rect 317604 -7504 318204 -7482
rect 335604 -5986 336204 12698
rect 342804 56454 343404 77000
rect 342804 56218 342986 56454
rect 343222 56218 343404 56454
rect 342804 56134 343404 56218
rect 342804 55898 342986 56134
rect 343222 55898 343404 56134
rect 342804 20454 343404 55898
rect 342804 20218 342986 20454
rect 343222 20218 343404 20454
rect 342804 20134 343404 20218
rect 342804 19898 342986 20134
rect 343222 19898 343404 20134
rect 342804 -1286 343404 19898
rect 342804 -1522 342986 -1286
rect 343222 -1522 343404 -1286
rect 342804 -1606 343404 -1522
rect 342804 -1842 342986 -1606
rect 343222 -1842 343404 -1606
rect 342804 -1864 343404 -1842
rect 346404 60054 347004 77000
rect 346404 59818 346586 60054
rect 346822 59818 347004 60054
rect 346404 59734 347004 59818
rect 346404 59498 346586 59734
rect 346822 59498 347004 59734
rect 346404 24054 347004 59498
rect 346404 23818 346586 24054
rect 346822 23818 347004 24054
rect 346404 23734 347004 23818
rect 346404 23498 346586 23734
rect 346822 23498 347004 23734
rect 346404 -3166 347004 23498
rect 346404 -3402 346586 -3166
rect 346822 -3402 347004 -3166
rect 346404 -3486 347004 -3402
rect 346404 -3722 346586 -3486
rect 346822 -3722 347004 -3486
rect 346404 -3744 347004 -3722
rect 350004 63654 350604 77000
rect 350004 63418 350186 63654
rect 350422 63418 350604 63654
rect 350004 63334 350604 63418
rect 350004 63098 350186 63334
rect 350422 63098 350604 63334
rect 350004 27654 350604 63098
rect 350004 27418 350186 27654
rect 350422 27418 350604 27654
rect 350004 27334 350604 27418
rect 350004 27098 350186 27334
rect 350422 27098 350604 27334
rect 350004 -5046 350604 27098
rect 350004 -5282 350186 -5046
rect 350422 -5282 350604 -5046
rect 350004 -5366 350604 -5282
rect 350004 -5602 350186 -5366
rect 350422 -5602 350604 -5366
rect 350004 -5624 350604 -5602
rect 353604 67254 354204 77000
rect 353604 67018 353786 67254
rect 354022 67018 354204 67254
rect 353604 66934 354204 67018
rect 353604 66698 353786 66934
rect 354022 66698 354204 66934
rect 353604 31254 354204 66698
rect 353604 31018 353786 31254
rect 354022 31018 354204 31254
rect 353604 30934 354204 31018
rect 353604 30698 353786 30934
rect 354022 30698 354204 30934
rect 335604 -6222 335786 -5986
rect 336022 -6222 336204 -5986
rect 335604 -6306 336204 -6222
rect 335604 -6542 335786 -6306
rect 336022 -6542 336204 -6306
rect 335604 -7504 336204 -6542
rect 353604 -6926 354204 30698
rect 360804 74454 361404 77000
rect 360804 74218 360986 74454
rect 361222 74218 361404 74454
rect 360804 74134 361404 74218
rect 360804 73898 360986 74134
rect 361222 73898 361404 74134
rect 360804 38454 361404 73898
rect 360804 38218 360986 38454
rect 361222 38218 361404 38454
rect 360804 38134 361404 38218
rect 360804 37898 360986 38134
rect 361222 37898 361404 38134
rect 360804 2454 361404 37898
rect 360804 2218 360986 2454
rect 361222 2218 361404 2454
rect 360804 2134 361404 2218
rect 360804 1898 360986 2134
rect 361222 1898 361404 2134
rect 360804 -346 361404 1898
rect 360804 -582 360986 -346
rect 361222 -582 361404 -346
rect 360804 -666 361404 -582
rect 360804 -902 360986 -666
rect 361222 -902 361404 -666
rect 360804 -1864 361404 -902
rect 364404 42054 365004 77000
rect 364404 41818 364586 42054
rect 364822 41818 365004 42054
rect 364404 41734 365004 41818
rect 364404 41498 364586 41734
rect 364822 41498 365004 41734
rect 364404 6054 365004 41498
rect 364404 5818 364586 6054
rect 364822 5818 365004 6054
rect 364404 5734 365004 5818
rect 364404 5498 364586 5734
rect 364822 5498 365004 5734
rect 364404 -2226 365004 5498
rect 364404 -2462 364586 -2226
rect 364822 -2462 365004 -2226
rect 364404 -2546 365004 -2462
rect 364404 -2782 364586 -2546
rect 364822 -2782 365004 -2546
rect 364404 -3744 365004 -2782
rect 368004 45654 368604 77000
rect 368004 45418 368186 45654
rect 368422 45418 368604 45654
rect 368004 45334 368604 45418
rect 368004 45098 368186 45334
rect 368422 45098 368604 45334
rect 368004 9654 368604 45098
rect 368004 9418 368186 9654
rect 368422 9418 368604 9654
rect 368004 9334 368604 9418
rect 368004 9098 368186 9334
rect 368422 9098 368604 9334
rect 368004 -4106 368604 9098
rect 368004 -4342 368186 -4106
rect 368422 -4342 368604 -4106
rect 368004 -4426 368604 -4342
rect 368004 -4662 368186 -4426
rect 368422 -4662 368604 -4426
rect 368004 -5624 368604 -4662
rect 371604 49254 372204 77000
rect 371604 49018 371786 49254
rect 372022 49018 372204 49254
rect 371604 48934 372204 49018
rect 371604 48698 371786 48934
rect 372022 48698 372204 48934
rect 371604 13254 372204 48698
rect 371604 13018 371786 13254
rect 372022 13018 372204 13254
rect 371604 12934 372204 13018
rect 371604 12698 371786 12934
rect 372022 12698 372204 12934
rect 353604 -7162 353786 -6926
rect 354022 -7162 354204 -6926
rect 353604 -7246 354204 -7162
rect 353604 -7482 353786 -7246
rect 354022 -7482 354204 -7246
rect 353604 -7504 354204 -7482
rect 371604 -5986 372204 12698
rect 378804 56454 379404 77000
rect 378804 56218 378986 56454
rect 379222 56218 379404 56454
rect 378804 56134 379404 56218
rect 378804 55898 378986 56134
rect 379222 55898 379404 56134
rect 378804 20454 379404 55898
rect 378804 20218 378986 20454
rect 379222 20218 379404 20454
rect 378804 20134 379404 20218
rect 378804 19898 378986 20134
rect 379222 19898 379404 20134
rect 378804 -1286 379404 19898
rect 378804 -1522 378986 -1286
rect 379222 -1522 379404 -1286
rect 378804 -1606 379404 -1522
rect 378804 -1842 378986 -1606
rect 379222 -1842 379404 -1606
rect 378804 -1864 379404 -1842
rect 382404 60054 383004 77000
rect 382404 59818 382586 60054
rect 382822 59818 383004 60054
rect 382404 59734 383004 59818
rect 382404 59498 382586 59734
rect 382822 59498 383004 59734
rect 382404 24054 383004 59498
rect 382404 23818 382586 24054
rect 382822 23818 383004 24054
rect 382404 23734 383004 23818
rect 382404 23498 382586 23734
rect 382822 23498 383004 23734
rect 382404 -3166 383004 23498
rect 382404 -3402 382586 -3166
rect 382822 -3402 383004 -3166
rect 382404 -3486 383004 -3402
rect 382404 -3722 382586 -3486
rect 382822 -3722 383004 -3486
rect 382404 -3744 383004 -3722
rect 386004 63654 386604 77000
rect 386004 63418 386186 63654
rect 386422 63418 386604 63654
rect 386004 63334 386604 63418
rect 386004 63098 386186 63334
rect 386422 63098 386604 63334
rect 386004 27654 386604 63098
rect 386004 27418 386186 27654
rect 386422 27418 386604 27654
rect 386004 27334 386604 27418
rect 386004 27098 386186 27334
rect 386422 27098 386604 27334
rect 386004 -5046 386604 27098
rect 386004 -5282 386186 -5046
rect 386422 -5282 386604 -5046
rect 386004 -5366 386604 -5282
rect 386004 -5602 386186 -5366
rect 386422 -5602 386604 -5366
rect 386004 -5624 386604 -5602
rect 389604 67254 390204 77000
rect 389604 67018 389786 67254
rect 390022 67018 390204 67254
rect 389604 66934 390204 67018
rect 389604 66698 389786 66934
rect 390022 66698 390204 66934
rect 389604 31254 390204 66698
rect 389604 31018 389786 31254
rect 390022 31018 390204 31254
rect 389604 30934 390204 31018
rect 389604 30698 389786 30934
rect 390022 30698 390204 30934
rect 371604 -6222 371786 -5986
rect 372022 -6222 372204 -5986
rect 371604 -6306 372204 -6222
rect 371604 -6542 371786 -6306
rect 372022 -6542 372204 -6306
rect 371604 -7504 372204 -6542
rect 389604 -6926 390204 30698
rect 396804 74454 397404 77000
rect 396804 74218 396986 74454
rect 397222 74218 397404 74454
rect 396804 74134 397404 74218
rect 396804 73898 396986 74134
rect 397222 73898 397404 74134
rect 396804 38454 397404 73898
rect 396804 38218 396986 38454
rect 397222 38218 397404 38454
rect 396804 38134 397404 38218
rect 396804 37898 396986 38134
rect 397222 37898 397404 38134
rect 396804 2454 397404 37898
rect 396804 2218 396986 2454
rect 397222 2218 397404 2454
rect 396804 2134 397404 2218
rect 396804 1898 396986 2134
rect 397222 1898 397404 2134
rect 396804 -346 397404 1898
rect 396804 -582 396986 -346
rect 397222 -582 397404 -346
rect 396804 -666 397404 -582
rect 396804 -902 396986 -666
rect 397222 -902 397404 -666
rect 396804 -1864 397404 -902
rect 400404 42054 401004 77000
rect 400404 41818 400586 42054
rect 400822 41818 401004 42054
rect 400404 41734 401004 41818
rect 400404 41498 400586 41734
rect 400822 41498 401004 41734
rect 400404 6054 401004 41498
rect 400404 5818 400586 6054
rect 400822 5818 401004 6054
rect 400404 5734 401004 5818
rect 400404 5498 400586 5734
rect 400822 5498 401004 5734
rect 400404 -2226 401004 5498
rect 400404 -2462 400586 -2226
rect 400822 -2462 401004 -2226
rect 400404 -2546 401004 -2462
rect 400404 -2782 400586 -2546
rect 400822 -2782 401004 -2546
rect 400404 -3744 401004 -2782
rect 404004 45654 404604 77000
rect 404004 45418 404186 45654
rect 404422 45418 404604 45654
rect 404004 45334 404604 45418
rect 404004 45098 404186 45334
rect 404422 45098 404604 45334
rect 404004 9654 404604 45098
rect 404004 9418 404186 9654
rect 404422 9418 404604 9654
rect 404004 9334 404604 9418
rect 404004 9098 404186 9334
rect 404422 9098 404604 9334
rect 404004 -4106 404604 9098
rect 404004 -4342 404186 -4106
rect 404422 -4342 404604 -4106
rect 404004 -4426 404604 -4342
rect 404004 -4662 404186 -4426
rect 404422 -4662 404604 -4426
rect 404004 -5624 404604 -4662
rect 407604 49254 408204 77000
rect 407604 49018 407786 49254
rect 408022 49018 408204 49254
rect 407604 48934 408204 49018
rect 407604 48698 407786 48934
rect 408022 48698 408204 48934
rect 407604 13254 408204 48698
rect 407604 13018 407786 13254
rect 408022 13018 408204 13254
rect 407604 12934 408204 13018
rect 407604 12698 407786 12934
rect 408022 12698 408204 12934
rect 389604 -7162 389786 -6926
rect 390022 -7162 390204 -6926
rect 389604 -7246 390204 -7162
rect 389604 -7482 389786 -7246
rect 390022 -7482 390204 -7246
rect 389604 -7504 390204 -7482
rect 407604 -5986 408204 12698
rect 414804 56454 415404 77000
rect 414804 56218 414986 56454
rect 415222 56218 415404 56454
rect 414804 56134 415404 56218
rect 414804 55898 414986 56134
rect 415222 55898 415404 56134
rect 414804 20454 415404 55898
rect 414804 20218 414986 20454
rect 415222 20218 415404 20454
rect 414804 20134 415404 20218
rect 414804 19898 414986 20134
rect 415222 19898 415404 20134
rect 414804 -1286 415404 19898
rect 414804 -1522 414986 -1286
rect 415222 -1522 415404 -1286
rect 414804 -1606 415404 -1522
rect 414804 -1842 414986 -1606
rect 415222 -1842 415404 -1606
rect 414804 -1864 415404 -1842
rect 418404 60054 419004 77000
rect 418404 59818 418586 60054
rect 418822 59818 419004 60054
rect 418404 59734 419004 59818
rect 418404 59498 418586 59734
rect 418822 59498 419004 59734
rect 418404 24054 419004 59498
rect 418404 23818 418586 24054
rect 418822 23818 419004 24054
rect 418404 23734 419004 23818
rect 418404 23498 418586 23734
rect 418822 23498 419004 23734
rect 418404 -3166 419004 23498
rect 418404 -3402 418586 -3166
rect 418822 -3402 419004 -3166
rect 418404 -3486 419004 -3402
rect 418404 -3722 418586 -3486
rect 418822 -3722 419004 -3486
rect 418404 -3744 419004 -3722
rect 422004 63654 422604 77000
rect 422004 63418 422186 63654
rect 422422 63418 422604 63654
rect 422004 63334 422604 63418
rect 422004 63098 422186 63334
rect 422422 63098 422604 63334
rect 422004 27654 422604 63098
rect 422004 27418 422186 27654
rect 422422 27418 422604 27654
rect 422004 27334 422604 27418
rect 422004 27098 422186 27334
rect 422422 27098 422604 27334
rect 422004 -5046 422604 27098
rect 422004 -5282 422186 -5046
rect 422422 -5282 422604 -5046
rect 422004 -5366 422604 -5282
rect 422004 -5602 422186 -5366
rect 422422 -5602 422604 -5366
rect 422004 -5624 422604 -5602
rect 425604 67254 426204 77000
rect 425604 67018 425786 67254
rect 426022 67018 426204 67254
rect 425604 66934 426204 67018
rect 425604 66698 425786 66934
rect 426022 66698 426204 66934
rect 425604 31254 426204 66698
rect 425604 31018 425786 31254
rect 426022 31018 426204 31254
rect 425604 30934 426204 31018
rect 425604 30698 425786 30934
rect 426022 30698 426204 30934
rect 407604 -6222 407786 -5986
rect 408022 -6222 408204 -5986
rect 407604 -6306 408204 -6222
rect 407604 -6542 407786 -6306
rect 408022 -6542 408204 -6306
rect 407604 -7504 408204 -6542
rect 425604 -6926 426204 30698
rect 432804 74454 433404 77000
rect 432804 74218 432986 74454
rect 433222 74218 433404 74454
rect 432804 74134 433404 74218
rect 432804 73898 432986 74134
rect 433222 73898 433404 74134
rect 432804 38454 433404 73898
rect 432804 38218 432986 38454
rect 433222 38218 433404 38454
rect 432804 38134 433404 38218
rect 432804 37898 432986 38134
rect 433222 37898 433404 38134
rect 432804 2454 433404 37898
rect 432804 2218 432986 2454
rect 433222 2218 433404 2454
rect 432804 2134 433404 2218
rect 432804 1898 432986 2134
rect 433222 1898 433404 2134
rect 432804 -346 433404 1898
rect 432804 -582 432986 -346
rect 433222 -582 433404 -346
rect 432804 -666 433404 -582
rect 432804 -902 432986 -666
rect 433222 -902 433404 -666
rect 432804 -1864 433404 -902
rect 436404 42054 437004 77000
rect 436404 41818 436586 42054
rect 436822 41818 437004 42054
rect 436404 41734 437004 41818
rect 436404 41498 436586 41734
rect 436822 41498 437004 41734
rect 436404 6054 437004 41498
rect 436404 5818 436586 6054
rect 436822 5818 437004 6054
rect 436404 5734 437004 5818
rect 436404 5498 436586 5734
rect 436822 5498 437004 5734
rect 436404 -2226 437004 5498
rect 436404 -2462 436586 -2226
rect 436822 -2462 437004 -2226
rect 436404 -2546 437004 -2462
rect 436404 -2782 436586 -2546
rect 436822 -2782 437004 -2546
rect 436404 -3744 437004 -2782
rect 440004 45654 440604 77000
rect 440004 45418 440186 45654
rect 440422 45418 440604 45654
rect 440004 45334 440604 45418
rect 440004 45098 440186 45334
rect 440422 45098 440604 45334
rect 440004 9654 440604 45098
rect 440004 9418 440186 9654
rect 440422 9418 440604 9654
rect 440004 9334 440604 9418
rect 440004 9098 440186 9334
rect 440422 9098 440604 9334
rect 440004 -4106 440604 9098
rect 440004 -4342 440186 -4106
rect 440422 -4342 440604 -4106
rect 440004 -4426 440604 -4342
rect 440004 -4662 440186 -4426
rect 440422 -4662 440604 -4426
rect 440004 -5624 440604 -4662
rect 443604 49254 444204 77000
rect 443604 49018 443786 49254
rect 444022 49018 444204 49254
rect 443604 48934 444204 49018
rect 443604 48698 443786 48934
rect 444022 48698 444204 48934
rect 443604 13254 444204 48698
rect 443604 13018 443786 13254
rect 444022 13018 444204 13254
rect 443604 12934 444204 13018
rect 443604 12698 443786 12934
rect 444022 12698 444204 12934
rect 425604 -7162 425786 -6926
rect 426022 -7162 426204 -6926
rect 425604 -7246 426204 -7162
rect 425604 -7482 425786 -7246
rect 426022 -7482 426204 -7246
rect 425604 -7504 426204 -7482
rect 443604 -5986 444204 12698
rect 450804 56454 451404 77000
rect 450804 56218 450986 56454
rect 451222 56218 451404 56454
rect 450804 56134 451404 56218
rect 450804 55898 450986 56134
rect 451222 55898 451404 56134
rect 450804 20454 451404 55898
rect 450804 20218 450986 20454
rect 451222 20218 451404 20454
rect 450804 20134 451404 20218
rect 450804 19898 450986 20134
rect 451222 19898 451404 20134
rect 450804 -1286 451404 19898
rect 450804 -1522 450986 -1286
rect 451222 -1522 451404 -1286
rect 450804 -1606 451404 -1522
rect 450804 -1842 450986 -1606
rect 451222 -1842 451404 -1606
rect 450804 -1864 451404 -1842
rect 454404 60054 455004 77000
rect 454404 59818 454586 60054
rect 454822 59818 455004 60054
rect 454404 59734 455004 59818
rect 454404 59498 454586 59734
rect 454822 59498 455004 59734
rect 454404 24054 455004 59498
rect 454404 23818 454586 24054
rect 454822 23818 455004 24054
rect 454404 23734 455004 23818
rect 454404 23498 454586 23734
rect 454822 23498 455004 23734
rect 454404 -3166 455004 23498
rect 454404 -3402 454586 -3166
rect 454822 -3402 455004 -3166
rect 454404 -3486 455004 -3402
rect 454404 -3722 454586 -3486
rect 454822 -3722 455004 -3486
rect 454404 -3744 455004 -3722
rect 458004 63654 458604 77000
rect 458004 63418 458186 63654
rect 458422 63418 458604 63654
rect 458004 63334 458604 63418
rect 458004 63098 458186 63334
rect 458422 63098 458604 63334
rect 458004 27654 458604 63098
rect 458004 27418 458186 27654
rect 458422 27418 458604 27654
rect 458004 27334 458604 27418
rect 458004 27098 458186 27334
rect 458422 27098 458604 27334
rect 458004 -5046 458604 27098
rect 458004 -5282 458186 -5046
rect 458422 -5282 458604 -5046
rect 458004 -5366 458604 -5282
rect 458004 -5602 458186 -5366
rect 458422 -5602 458604 -5366
rect 458004 -5624 458604 -5602
rect 461604 67254 462204 77000
rect 461604 67018 461786 67254
rect 462022 67018 462204 67254
rect 461604 66934 462204 67018
rect 461604 66698 461786 66934
rect 462022 66698 462204 66934
rect 461604 31254 462204 66698
rect 461604 31018 461786 31254
rect 462022 31018 462204 31254
rect 461604 30934 462204 31018
rect 461604 30698 461786 30934
rect 462022 30698 462204 30934
rect 443604 -6222 443786 -5986
rect 444022 -6222 444204 -5986
rect 443604 -6306 444204 -6222
rect 443604 -6542 443786 -6306
rect 444022 -6542 444204 -6306
rect 443604 -7504 444204 -6542
rect 461604 -6926 462204 30698
rect 468804 74454 469404 77000
rect 468804 74218 468986 74454
rect 469222 74218 469404 74454
rect 468804 74134 469404 74218
rect 468804 73898 468986 74134
rect 469222 73898 469404 74134
rect 468804 38454 469404 73898
rect 468804 38218 468986 38454
rect 469222 38218 469404 38454
rect 468804 38134 469404 38218
rect 468804 37898 468986 38134
rect 469222 37898 469404 38134
rect 468804 2454 469404 37898
rect 468804 2218 468986 2454
rect 469222 2218 469404 2454
rect 468804 2134 469404 2218
rect 468804 1898 468986 2134
rect 469222 1898 469404 2134
rect 468804 -346 469404 1898
rect 468804 -582 468986 -346
rect 469222 -582 469404 -346
rect 468804 -666 469404 -582
rect 468804 -902 468986 -666
rect 469222 -902 469404 -666
rect 468804 -1864 469404 -902
rect 472404 42054 473004 77000
rect 472404 41818 472586 42054
rect 472822 41818 473004 42054
rect 472404 41734 473004 41818
rect 472404 41498 472586 41734
rect 472822 41498 473004 41734
rect 472404 6054 473004 41498
rect 472404 5818 472586 6054
rect 472822 5818 473004 6054
rect 472404 5734 473004 5818
rect 472404 5498 472586 5734
rect 472822 5498 473004 5734
rect 472404 -2226 473004 5498
rect 472404 -2462 472586 -2226
rect 472822 -2462 473004 -2226
rect 472404 -2546 473004 -2462
rect 472404 -2782 472586 -2546
rect 472822 -2782 473004 -2546
rect 472404 -3744 473004 -2782
rect 476004 45654 476604 77000
rect 476004 45418 476186 45654
rect 476422 45418 476604 45654
rect 476004 45334 476604 45418
rect 476004 45098 476186 45334
rect 476422 45098 476604 45334
rect 476004 9654 476604 45098
rect 476004 9418 476186 9654
rect 476422 9418 476604 9654
rect 476004 9334 476604 9418
rect 476004 9098 476186 9334
rect 476422 9098 476604 9334
rect 476004 -4106 476604 9098
rect 476004 -4342 476186 -4106
rect 476422 -4342 476604 -4106
rect 476004 -4426 476604 -4342
rect 476004 -4662 476186 -4426
rect 476422 -4662 476604 -4426
rect 476004 -5624 476604 -4662
rect 479604 49254 480204 77000
rect 479604 49018 479786 49254
rect 480022 49018 480204 49254
rect 479604 48934 480204 49018
rect 479604 48698 479786 48934
rect 480022 48698 480204 48934
rect 479604 13254 480204 48698
rect 479604 13018 479786 13254
rect 480022 13018 480204 13254
rect 479604 12934 480204 13018
rect 479604 12698 479786 12934
rect 480022 12698 480204 12934
rect 461604 -7162 461786 -6926
rect 462022 -7162 462204 -6926
rect 461604 -7246 462204 -7162
rect 461604 -7482 461786 -7246
rect 462022 -7482 462204 -7246
rect 461604 -7504 462204 -7482
rect 479604 -5986 480204 12698
rect 486804 56454 487404 77000
rect 486804 56218 486986 56454
rect 487222 56218 487404 56454
rect 486804 56134 487404 56218
rect 486804 55898 486986 56134
rect 487222 55898 487404 56134
rect 486804 20454 487404 55898
rect 486804 20218 486986 20454
rect 487222 20218 487404 20454
rect 486804 20134 487404 20218
rect 486804 19898 486986 20134
rect 487222 19898 487404 20134
rect 486804 -1286 487404 19898
rect 486804 -1522 486986 -1286
rect 487222 -1522 487404 -1286
rect 486804 -1606 487404 -1522
rect 486804 -1842 486986 -1606
rect 487222 -1842 487404 -1606
rect 486804 -1864 487404 -1842
rect 490404 60054 491004 77000
rect 490404 59818 490586 60054
rect 490822 59818 491004 60054
rect 490404 59734 491004 59818
rect 490404 59498 490586 59734
rect 490822 59498 491004 59734
rect 490404 24054 491004 59498
rect 490404 23818 490586 24054
rect 490822 23818 491004 24054
rect 490404 23734 491004 23818
rect 490404 23498 490586 23734
rect 490822 23498 491004 23734
rect 490404 -3166 491004 23498
rect 490404 -3402 490586 -3166
rect 490822 -3402 491004 -3166
rect 490404 -3486 491004 -3402
rect 490404 -3722 490586 -3486
rect 490822 -3722 491004 -3486
rect 490404 -3744 491004 -3722
rect 494004 63654 494604 77000
rect 494004 63418 494186 63654
rect 494422 63418 494604 63654
rect 494004 63334 494604 63418
rect 494004 63098 494186 63334
rect 494422 63098 494604 63334
rect 494004 27654 494604 63098
rect 494004 27418 494186 27654
rect 494422 27418 494604 27654
rect 494004 27334 494604 27418
rect 494004 27098 494186 27334
rect 494422 27098 494604 27334
rect 494004 -5046 494604 27098
rect 494004 -5282 494186 -5046
rect 494422 -5282 494604 -5046
rect 494004 -5366 494604 -5282
rect 494004 -5602 494186 -5366
rect 494422 -5602 494604 -5366
rect 494004 -5624 494604 -5602
rect 497604 67254 498204 77000
rect 497604 67018 497786 67254
rect 498022 67018 498204 67254
rect 497604 66934 498204 67018
rect 497604 66698 497786 66934
rect 498022 66698 498204 66934
rect 497604 31254 498204 66698
rect 497604 31018 497786 31254
rect 498022 31018 498204 31254
rect 497604 30934 498204 31018
rect 497604 30698 497786 30934
rect 498022 30698 498204 30934
rect 479604 -6222 479786 -5986
rect 480022 -6222 480204 -5986
rect 479604 -6306 480204 -6222
rect 479604 -6542 479786 -6306
rect 480022 -6542 480204 -6306
rect 479604 -7504 480204 -6542
rect 497604 -6926 498204 30698
rect 504804 74454 505404 77000
rect 504804 74218 504986 74454
rect 505222 74218 505404 74454
rect 504804 74134 505404 74218
rect 504804 73898 504986 74134
rect 505222 73898 505404 74134
rect 504804 38454 505404 73898
rect 504804 38218 504986 38454
rect 505222 38218 505404 38454
rect 504804 38134 505404 38218
rect 504804 37898 504986 38134
rect 505222 37898 505404 38134
rect 504804 2454 505404 37898
rect 504804 2218 504986 2454
rect 505222 2218 505404 2454
rect 504804 2134 505404 2218
rect 504804 1898 504986 2134
rect 505222 1898 505404 2134
rect 504804 -346 505404 1898
rect 504804 -582 504986 -346
rect 505222 -582 505404 -346
rect 504804 -666 505404 -582
rect 504804 -902 504986 -666
rect 505222 -902 505404 -666
rect 504804 -1864 505404 -902
rect 508404 42054 509004 77000
rect 508404 41818 508586 42054
rect 508822 41818 509004 42054
rect 508404 41734 509004 41818
rect 508404 41498 508586 41734
rect 508822 41498 509004 41734
rect 508404 6054 509004 41498
rect 508404 5818 508586 6054
rect 508822 5818 509004 6054
rect 508404 5734 509004 5818
rect 508404 5498 508586 5734
rect 508822 5498 509004 5734
rect 508404 -2226 509004 5498
rect 508404 -2462 508586 -2226
rect 508822 -2462 509004 -2226
rect 508404 -2546 509004 -2462
rect 508404 -2782 508586 -2546
rect 508822 -2782 509004 -2546
rect 508404 -3744 509004 -2782
rect 512004 45654 512604 77000
rect 512004 45418 512186 45654
rect 512422 45418 512604 45654
rect 512004 45334 512604 45418
rect 512004 45098 512186 45334
rect 512422 45098 512604 45334
rect 512004 9654 512604 45098
rect 512004 9418 512186 9654
rect 512422 9418 512604 9654
rect 512004 9334 512604 9418
rect 512004 9098 512186 9334
rect 512422 9098 512604 9334
rect 512004 -4106 512604 9098
rect 512004 -4342 512186 -4106
rect 512422 -4342 512604 -4106
rect 512004 -4426 512604 -4342
rect 512004 -4662 512186 -4426
rect 512422 -4662 512604 -4426
rect 512004 -5624 512604 -4662
rect 515604 49254 516204 77000
rect 515604 49018 515786 49254
rect 516022 49018 516204 49254
rect 515604 48934 516204 49018
rect 515604 48698 515786 48934
rect 516022 48698 516204 48934
rect 515604 13254 516204 48698
rect 515604 13018 515786 13254
rect 516022 13018 516204 13254
rect 515604 12934 516204 13018
rect 515604 12698 515786 12934
rect 516022 12698 516204 12934
rect 497604 -7162 497786 -6926
rect 498022 -7162 498204 -6926
rect 497604 -7246 498204 -7162
rect 497604 -7482 497786 -7246
rect 498022 -7482 498204 -7246
rect 497604 -7504 498204 -7482
rect 515604 -5986 516204 12698
rect 522804 56454 523404 77000
rect 522804 56218 522986 56454
rect 523222 56218 523404 56454
rect 522804 56134 523404 56218
rect 522804 55898 522986 56134
rect 523222 55898 523404 56134
rect 522804 20454 523404 55898
rect 522804 20218 522986 20454
rect 523222 20218 523404 20454
rect 522804 20134 523404 20218
rect 522804 19898 522986 20134
rect 523222 19898 523404 20134
rect 522804 -1286 523404 19898
rect 522804 -1522 522986 -1286
rect 523222 -1522 523404 -1286
rect 522804 -1606 523404 -1522
rect 522804 -1842 522986 -1606
rect 523222 -1842 523404 -1606
rect 522804 -1864 523404 -1842
rect 526404 60054 527004 77000
rect 526404 59818 526586 60054
rect 526822 59818 527004 60054
rect 526404 59734 527004 59818
rect 526404 59498 526586 59734
rect 526822 59498 527004 59734
rect 526404 24054 527004 59498
rect 526404 23818 526586 24054
rect 526822 23818 527004 24054
rect 526404 23734 527004 23818
rect 526404 23498 526586 23734
rect 526822 23498 527004 23734
rect 526404 -3166 527004 23498
rect 526404 -3402 526586 -3166
rect 526822 -3402 527004 -3166
rect 526404 -3486 527004 -3402
rect 526404 -3722 526586 -3486
rect 526822 -3722 527004 -3486
rect 526404 -3744 527004 -3722
rect 530004 63654 530604 77000
rect 530004 63418 530186 63654
rect 530422 63418 530604 63654
rect 530004 63334 530604 63418
rect 530004 63098 530186 63334
rect 530422 63098 530604 63334
rect 530004 27654 530604 63098
rect 530004 27418 530186 27654
rect 530422 27418 530604 27654
rect 530004 27334 530604 27418
rect 530004 27098 530186 27334
rect 530422 27098 530604 27334
rect 530004 -5046 530604 27098
rect 530004 -5282 530186 -5046
rect 530422 -5282 530604 -5046
rect 530004 -5366 530604 -5282
rect 530004 -5602 530186 -5366
rect 530422 -5602 530604 -5366
rect 530004 -5624 530604 -5602
rect 533604 67254 534204 102698
rect 533604 67018 533786 67254
rect 534022 67018 534204 67254
rect 533604 66934 534204 67018
rect 533604 66698 533786 66934
rect 534022 66698 534204 66934
rect 533604 31254 534204 66698
rect 533604 31018 533786 31254
rect 534022 31018 534204 31254
rect 533604 30934 534204 31018
rect 533604 30698 533786 30934
rect 534022 30698 534204 30934
rect 515604 -6222 515786 -5986
rect 516022 -6222 516204 -5986
rect 515604 -6306 516204 -6222
rect 515604 -6542 515786 -6306
rect 516022 -6542 516204 -6306
rect 515604 -7504 516204 -6542
rect 533604 -6926 534204 30698
rect 540804 704838 541404 705800
rect 540804 704602 540986 704838
rect 541222 704602 541404 704838
rect 540804 704518 541404 704602
rect 540804 704282 540986 704518
rect 541222 704282 541404 704518
rect 540804 686454 541404 704282
rect 540804 686218 540986 686454
rect 541222 686218 541404 686454
rect 540804 686134 541404 686218
rect 540804 685898 540986 686134
rect 541222 685898 541404 686134
rect 540804 650454 541404 685898
rect 540804 650218 540986 650454
rect 541222 650218 541404 650454
rect 540804 650134 541404 650218
rect 540804 649898 540986 650134
rect 541222 649898 541404 650134
rect 540804 614454 541404 649898
rect 540804 614218 540986 614454
rect 541222 614218 541404 614454
rect 540804 614134 541404 614218
rect 540804 613898 540986 614134
rect 541222 613898 541404 614134
rect 540804 578454 541404 613898
rect 540804 578218 540986 578454
rect 541222 578218 541404 578454
rect 540804 578134 541404 578218
rect 540804 577898 540986 578134
rect 541222 577898 541404 578134
rect 540804 542454 541404 577898
rect 540804 542218 540986 542454
rect 541222 542218 541404 542454
rect 540804 542134 541404 542218
rect 540804 541898 540986 542134
rect 541222 541898 541404 542134
rect 540804 506454 541404 541898
rect 540804 506218 540986 506454
rect 541222 506218 541404 506454
rect 540804 506134 541404 506218
rect 540804 505898 540986 506134
rect 541222 505898 541404 506134
rect 540804 470454 541404 505898
rect 540804 470218 540986 470454
rect 541222 470218 541404 470454
rect 540804 470134 541404 470218
rect 540804 469898 540986 470134
rect 541222 469898 541404 470134
rect 540804 434454 541404 469898
rect 540804 434218 540986 434454
rect 541222 434218 541404 434454
rect 540804 434134 541404 434218
rect 540804 433898 540986 434134
rect 541222 433898 541404 434134
rect 540804 398454 541404 433898
rect 540804 398218 540986 398454
rect 541222 398218 541404 398454
rect 540804 398134 541404 398218
rect 540804 397898 540986 398134
rect 541222 397898 541404 398134
rect 540804 362454 541404 397898
rect 540804 362218 540986 362454
rect 541222 362218 541404 362454
rect 540804 362134 541404 362218
rect 540804 361898 540986 362134
rect 541222 361898 541404 362134
rect 540804 326454 541404 361898
rect 540804 326218 540986 326454
rect 541222 326218 541404 326454
rect 540804 326134 541404 326218
rect 540804 325898 540986 326134
rect 541222 325898 541404 326134
rect 540804 290454 541404 325898
rect 540804 290218 540986 290454
rect 541222 290218 541404 290454
rect 540804 290134 541404 290218
rect 540804 289898 540986 290134
rect 541222 289898 541404 290134
rect 540804 254454 541404 289898
rect 540804 254218 540986 254454
rect 541222 254218 541404 254454
rect 540804 254134 541404 254218
rect 540804 253898 540986 254134
rect 541222 253898 541404 254134
rect 540804 218454 541404 253898
rect 540804 218218 540986 218454
rect 541222 218218 541404 218454
rect 540804 218134 541404 218218
rect 540804 217898 540986 218134
rect 541222 217898 541404 218134
rect 540804 182454 541404 217898
rect 540804 182218 540986 182454
rect 541222 182218 541404 182454
rect 540804 182134 541404 182218
rect 540804 181898 540986 182134
rect 541222 181898 541404 182134
rect 540804 146454 541404 181898
rect 540804 146218 540986 146454
rect 541222 146218 541404 146454
rect 540804 146134 541404 146218
rect 540804 145898 540986 146134
rect 541222 145898 541404 146134
rect 540804 110454 541404 145898
rect 540804 110218 540986 110454
rect 541222 110218 541404 110454
rect 540804 110134 541404 110218
rect 540804 109898 540986 110134
rect 541222 109898 541404 110134
rect 540804 74454 541404 109898
rect 540804 74218 540986 74454
rect 541222 74218 541404 74454
rect 540804 74134 541404 74218
rect 540804 73898 540986 74134
rect 541222 73898 541404 74134
rect 540804 38454 541404 73898
rect 540804 38218 540986 38454
rect 541222 38218 541404 38454
rect 540804 38134 541404 38218
rect 540804 37898 540986 38134
rect 541222 37898 541404 38134
rect 540804 2454 541404 37898
rect 540804 2218 540986 2454
rect 541222 2218 541404 2454
rect 540804 2134 541404 2218
rect 540804 1898 540986 2134
rect 541222 1898 541404 2134
rect 540804 -346 541404 1898
rect 540804 -582 540986 -346
rect 541222 -582 541404 -346
rect 540804 -666 541404 -582
rect 540804 -902 540986 -666
rect 541222 -902 541404 -666
rect 540804 -1864 541404 -902
rect 544404 690054 545004 706162
rect 544404 689818 544586 690054
rect 544822 689818 545004 690054
rect 544404 689734 545004 689818
rect 544404 689498 544586 689734
rect 544822 689498 545004 689734
rect 544404 654054 545004 689498
rect 544404 653818 544586 654054
rect 544822 653818 545004 654054
rect 544404 653734 545004 653818
rect 544404 653498 544586 653734
rect 544822 653498 545004 653734
rect 544404 618054 545004 653498
rect 544404 617818 544586 618054
rect 544822 617818 545004 618054
rect 544404 617734 545004 617818
rect 544404 617498 544586 617734
rect 544822 617498 545004 617734
rect 544404 582054 545004 617498
rect 544404 581818 544586 582054
rect 544822 581818 545004 582054
rect 544404 581734 545004 581818
rect 544404 581498 544586 581734
rect 544822 581498 545004 581734
rect 544404 546054 545004 581498
rect 544404 545818 544586 546054
rect 544822 545818 545004 546054
rect 544404 545734 545004 545818
rect 544404 545498 544586 545734
rect 544822 545498 545004 545734
rect 544404 510054 545004 545498
rect 544404 509818 544586 510054
rect 544822 509818 545004 510054
rect 544404 509734 545004 509818
rect 544404 509498 544586 509734
rect 544822 509498 545004 509734
rect 544404 474054 545004 509498
rect 544404 473818 544586 474054
rect 544822 473818 545004 474054
rect 544404 473734 545004 473818
rect 544404 473498 544586 473734
rect 544822 473498 545004 473734
rect 544404 438054 545004 473498
rect 544404 437818 544586 438054
rect 544822 437818 545004 438054
rect 544404 437734 545004 437818
rect 544404 437498 544586 437734
rect 544822 437498 545004 437734
rect 544404 402054 545004 437498
rect 544404 401818 544586 402054
rect 544822 401818 545004 402054
rect 544404 401734 545004 401818
rect 544404 401498 544586 401734
rect 544822 401498 545004 401734
rect 544404 366054 545004 401498
rect 544404 365818 544586 366054
rect 544822 365818 545004 366054
rect 544404 365734 545004 365818
rect 544404 365498 544586 365734
rect 544822 365498 545004 365734
rect 544404 330054 545004 365498
rect 544404 329818 544586 330054
rect 544822 329818 545004 330054
rect 544404 329734 545004 329818
rect 544404 329498 544586 329734
rect 544822 329498 545004 329734
rect 544404 294054 545004 329498
rect 544404 293818 544586 294054
rect 544822 293818 545004 294054
rect 544404 293734 545004 293818
rect 544404 293498 544586 293734
rect 544822 293498 545004 293734
rect 544404 258054 545004 293498
rect 544404 257818 544586 258054
rect 544822 257818 545004 258054
rect 544404 257734 545004 257818
rect 544404 257498 544586 257734
rect 544822 257498 545004 257734
rect 544404 222054 545004 257498
rect 544404 221818 544586 222054
rect 544822 221818 545004 222054
rect 544404 221734 545004 221818
rect 544404 221498 544586 221734
rect 544822 221498 545004 221734
rect 544404 186054 545004 221498
rect 544404 185818 544586 186054
rect 544822 185818 545004 186054
rect 544404 185734 545004 185818
rect 544404 185498 544586 185734
rect 544822 185498 545004 185734
rect 544404 150054 545004 185498
rect 544404 149818 544586 150054
rect 544822 149818 545004 150054
rect 544404 149734 545004 149818
rect 544404 149498 544586 149734
rect 544822 149498 545004 149734
rect 544404 114054 545004 149498
rect 544404 113818 544586 114054
rect 544822 113818 545004 114054
rect 544404 113734 545004 113818
rect 544404 113498 544586 113734
rect 544822 113498 545004 113734
rect 544404 78054 545004 113498
rect 544404 77818 544586 78054
rect 544822 77818 545004 78054
rect 544404 77734 545004 77818
rect 544404 77498 544586 77734
rect 544822 77498 545004 77734
rect 544404 42054 545004 77498
rect 544404 41818 544586 42054
rect 544822 41818 545004 42054
rect 544404 41734 545004 41818
rect 544404 41498 544586 41734
rect 544822 41498 545004 41734
rect 544404 6054 545004 41498
rect 544404 5818 544586 6054
rect 544822 5818 545004 6054
rect 544404 5734 545004 5818
rect 544404 5498 544586 5734
rect 544822 5498 545004 5734
rect 544404 -2226 545004 5498
rect 544404 -2462 544586 -2226
rect 544822 -2462 545004 -2226
rect 544404 -2546 545004 -2462
rect 544404 -2782 544586 -2546
rect 544822 -2782 545004 -2546
rect 544404 -3744 545004 -2782
rect 548004 693654 548604 708042
rect 548004 693418 548186 693654
rect 548422 693418 548604 693654
rect 548004 693334 548604 693418
rect 548004 693098 548186 693334
rect 548422 693098 548604 693334
rect 548004 657654 548604 693098
rect 548004 657418 548186 657654
rect 548422 657418 548604 657654
rect 548004 657334 548604 657418
rect 548004 657098 548186 657334
rect 548422 657098 548604 657334
rect 548004 621654 548604 657098
rect 548004 621418 548186 621654
rect 548422 621418 548604 621654
rect 548004 621334 548604 621418
rect 548004 621098 548186 621334
rect 548422 621098 548604 621334
rect 548004 585654 548604 621098
rect 548004 585418 548186 585654
rect 548422 585418 548604 585654
rect 548004 585334 548604 585418
rect 548004 585098 548186 585334
rect 548422 585098 548604 585334
rect 548004 549654 548604 585098
rect 548004 549418 548186 549654
rect 548422 549418 548604 549654
rect 548004 549334 548604 549418
rect 548004 549098 548186 549334
rect 548422 549098 548604 549334
rect 548004 513654 548604 549098
rect 548004 513418 548186 513654
rect 548422 513418 548604 513654
rect 548004 513334 548604 513418
rect 548004 513098 548186 513334
rect 548422 513098 548604 513334
rect 548004 477654 548604 513098
rect 548004 477418 548186 477654
rect 548422 477418 548604 477654
rect 548004 477334 548604 477418
rect 548004 477098 548186 477334
rect 548422 477098 548604 477334
rect 548004 441654 548604 477098
rect 548004 441418 548186 441654
rect 548422 441418 548604 441654
rect 548004 441334 548604 441418
rect 548004 441098 548186 441334
rect 548422 441098 548604 441334
rect 548004 405654 548604 441098
rect 548004 405418 548186 405654
rect 548422 405418 548604 405654
rect 548004 405334 548604 405418
rect 548004 405098 548186 405334
rect 548422 405098 548604 405334
rect 548004 369654 548604 405098
rect 548004 369418 548186 369654
rect 548422 369418 548604 369654
rect 548004 369334 548604 369418
rect 548004 369098 548186 369334
rect 548422 369098 548604 369334
rect 548004 333654 548604 369098
rect 548004 333418 548186 333654
rect 548422 333418 548604 333654
rect 548004 333334 548604 333418
rect 548004 333098 548186 333334
rect 548422 333098 548604 333334
rect 548004 297654 548604 333098
rect 548004 297418 548186 297654
rect 548422 297418 548604 297654
rect 548004 297334 548604 297418
rect 548004 297098 548186 297334
rect 548422 297098 548604 297334
rect 548004 261654 548604 297098
rect 548004 261418 548186 261654
rect 548422 261418 548604 261654
rect 548004 261334 548604 261418
rect 548004 261098 548186 261334
rect 548422 261098 548604 261334
rect 548004 225654 548604 261098
rect 548004 225418 548186 225654
rect 548422 225418 548604 225654
rect 548004 225334 548604 225418
rect 548004 225098 548186 225334
rect 548422 225098 548604 225334
rect 548004 189654 548604 225098
rect 548004 189418 548186 189654
rect 548422 189418 548604 189654
rect 548004 189334 548604 189418
rect 548004 189098 548186 189334
rect 548422 189098 548604 189334
rect 548004 153654 548604 189098
rect 548004 153418 548186 153654
rect 548422 153418 548604 153654
rect 548004 153334 548604 153418
rect 548004 153098 548186 153334
rect 548422 153098 548604 153334
rect 548004 117654 548604 153098
rect 548004 117418 548186 117654
rect 548422 117418 548604 117654
rect 548004 117334 548604 117418
rect 548004 117098 548186 117334
rect 548422 117098 548604 117334
rect 548004 81654 548604 117098
rect 548004 81418 548186 81654
rect 548422 81418 548604 81654
rect 548004 81334 548604 81418
rect 548004 81098 548186 81334
rect 548422 81098 548604 81334
rect 548004 45654 548604 81098
rect 548004 45418 548186 45654
rect 548422 45418 548604 45654
rect 548004 45334 548604 45418
rect 548004 45098 548186 45334
rect 548422 45098 548604 45334
rect 548004 9654 548604 45098
rect 548004 9418 548186 9654
rect 548422 9418 548604 9654
rect 548004 9334 548604 9418
rect 548004 9098 548186 9334
rect 548422 9098 548604 9334
rect 548004 -4106 548604 9098
rect 548004 -4342 548186 -4106
rect 548422 -4342 548604 -4106
rect 548004 -4426 548604 -4342
rect 548004 -4662 548186 -4426
rect 548422 -4662 548604 -4426
rect 548004 -5624 548604 -4662
rect 551604 697254 552204 709922
rect 569604 711418 570204 711440
rect 569604 711182 569786 711418
rect 570022 711182 570204 711418
rect 569604 711098 570204 711182
rect 569604 710862 569786 711098
rect 570022 710862 570204 711098
rect 566004 709538 566604 709560
rect 566004 709302 566186 709538
rect 566422 709302 566604 709538
rect 566004 709218 566604 709302
rect 566004 708982 566186 709218
rect 566422 708982 566604 709218
rect 562404 707658 563004 707680
rect 562404 707422 562586 707658
rect 562822 707422 563004 707658
rect 562404 707338 563004 707422
rect 562404 707102 562586 707338
rect 562822 707102 563004 707338
rect 551604 697018 551786 697254
rect 552022 697018 552204 697254
rect 551604 696934 552204 697018
rect 551604 696698 551786 696934
rect 552022 696698 552204 696934
rect 551604 661254 552204 696698
rect 551604 661018 551786 661254
rect 552022 661018 552204 661254
rect 551604 660934 552204 661018
rect 551604 660698 551786 660934
rect 552022 660698 552204 660934
rect 551604 625254 552204 660698
rect 551604 625018 551786 625254
rect 552022 625018 552204 625254
rect 551604 624934 552204 625018
rect 551604 624698 551786 624934
rect 552022 624698 552204 624934
rect 551604 589254 552204 624698
rect 551604 589018 551786 589254
rect 552022 589018 552204 589254
rect 551604 588934 552204 589018
rect 551604 588698 551786 588934
rect 552022 588698 552204 588934
rect 551604 553254 552204 588698
rect 551604 553018 551786 553254
rect 552022 553018 552204 553254
rect 551604 552934 552204 553018
rect 551604 552698 551786 552934
rect 552022 552698 552204 552934
rect 551604 517254 552204 552698
rect 551604 517018 551786 517254
rect 552022 517018 552204 517254
rect 551604 516934 552204 517018
rect 551604 516698 551786 516934
rect 552022 516698 552204 516934
rect 551604 481254 552204 516698
rect 551604 481018 551786 481254
rect 552022 481018 552204 481254
rect 551604 480934 552204 481018
rect 551604 480698 551786 480934
rect 552022 480698 552204 480934
rect 551604 445254 552204 480698
rect 551604 445018 551786 445254
rect 552022 445018 552204 445254
rect 551604 444934 552204 445018
rect 551604 444698 551786 444934
rect 552022 444698 552204 444934
rect 551604 409254 552204 444698
rect 551604 409018 551786 409254
rect 552022 409018 552204 409254
rect 551604 408934 552204 409018
rect 551604 408698 551786 408934
rect 552022 408698 552204 408934
rect 551604 373254 552204 408698
rect 551604 373018 551786 373254
rect 552022 373018 552204 373254
rect 551604 372934 552204 373018
rect 551604 372698 551786 372934
rect 552022 372698 552204 372934
rect 551604 337254 552204 372698
rect 551604 337018 551786 337254
rect 552022 337018 552204 337254
rect 551604 336934 552204 337018
rect 551604 336698 551786 336934
rect 552022 336698 552204 336934
rect 551604 301254 552204 336698
rect 551604 301018 551786 301254
rect 552022 301018 552204 301254
rect 551604 300934 552204 301018
rect 551604 300698 551786 300934
rect 552022 300698 552204 300934
rect 551604 265254 552204 300698
rect 551604 265018 551786 265254
rect 552022 265018 552204 265254
rect 551604 264934 552204 265018
rect 551604 264698 551786 264934
rect 552022 264698 552204 264934
rect 551604 229254 552204 264698
rect 551604 229018 551786 229254
rect 552022 229018 552204 229254
rect 551604 228934 552204 229018
rect 551604 228698 551786 228934
rect 552022 228698 552204 228934
rect 551604 193254 552204 228698
rect 551604 193018 551786 193254
rect 552022 193018 552204 193254
rect 551604 192934 552204 193018
rect 551604 192698 551786 192934
rect 552022 192698 552204 192934
rect 551604 157254 552204 192698
rect 551604 157018 551786 157254
rect 552022 157018 552204 157254
rect 551604 156934 552204 157018
rect 551604 156698 551786 156934
rect 552022 156698 552204 156934
rect 551604 121254 552204 156698
rect 551604 121018 551786 121254
rect 552022 121018 552204 121254
rect 551604 120934 552204 121018
rect 551604 120698 551786 120934
rect 552022 120698 552204 120934
rect 551604 85254 552204 120698
rect 551604 85018 551786 85254
rect 552022 85018 552204 85254
rect 551604 84934 552204 85018
rect 551604 84698 551786 84934
rect 552022 84698 552204 84934
rect 551604 49254 552204 84698
rect 551604 49018 551786 49254
rect 552022 49018 552204 49254
rect 551604 48934 552204 49018
rect 551604 48698 551786 48934
rect 552022 48698 552204 48934
rect 551604 13254 552204 48698
rect 551604 13018 551786 13254
rect 552022 13018 552204 13254
rect 551604 12934 552204 13018
rect 551604 12698 551786 12934
rect 552022 12698 552204 12934
rect 533604 -7162 533786 -6926
rect 534022 -7162 534204 -6926
rect 533604 -7246 534204 -7162
rect 533604 -7482 533786 -7246
rect 534022 -7482 534204 -7246
rect 533604 -7504 534204 -7482
rect 551604 -5986 552204 12698
rect 558804 705778 559404 705800
rect 558804 705542 558986 705778
rect 559222 705542 559404 705778
rect 558804 705458 559404 705542
rect 558804 705222 558986 705458
rect 559222 705222 559404 705458
rect 558804 668454 559404 705222
rect 558804 668218 558986 668454
rect 559222 668218 559404 668454
rect 558804 668134 559404 668218
rect 558804 667898 558986 668134
rect 559222 667898 559404 668134
rect 558804 632454 559404 667898
rect 558804 632218 558986 632454
rect 559222 632218 559404 632454
rect 558804 632134 559404 632218
rect 558804 631898 558986 632134
rect 559222 631898 559404 632134
rect 558804 596454 559404 631898
rect 558804 596218 558986 596454
rect 559222 596218 559404 596454
rect 558804 596134 559404 596218
rect 558804 595898 558986 596134
rect 559222 595898 559404 596134
rect 558804 560454 559404 595898
rect 558804 560218 558986 560454
rect 559222 560218 559404 560454
rect 558804 560134 559404 560218
rect 558804 559898 558986 560134
rect 559222 559898 559404 560134
rect 558804 524454 559404 559898
rect 558804 524218 558986 524454
rect 559222 524218 559404 524454
rect 558804 524134 559404 524218
rect 558804 523898 558986 524134
rect 559222 523898 559404 524134
rect 558804 488454 559404 523898
rect 558804 488218 558986 488454
rect 559222 488218 559404 488454
rect 558804 488134 559404 488218
rect 558804 487898 558986 488134
rect 559222 487898 559404 488134
rect 558804 452454 559404 487898
rect 558804 452218 558986 452454
rect 559222 452218 559404 452454
rect 558804 452134 559404 452218
rect 558804 451898 558986 452134
rect 559222 451898 559404 452134
rect 558804 416454 559404 451898
rect 558804 416218 558986 416454
rect 559222 416218 559404 416454
rect 558804 416134 559404 416218
rect 558804 415898 558986 416134
rect 559222 415898 559404 416134
rect 558804 380454 559404 415898
rect 558804 380218 558986 380454
rect 559222 380218 559404 380454
rect 558804 380134 559404 380218
rect 558804 379898 558986 380134
rect 559222 379898 559404 380134
rect 558804 344454 559404 379898
rect 558804 344218 558986 344454
rect 559222 344218 559404 344454
rect 558804 344134 559404 344218
rect 558804 343898 558986 344134
rect 559222 343898 559404 344134
rect 558804 308454 559404 343898
rect 558804 308218 558986 308454
rect 559222 308218 559404 308454
rect 558804 308134 559404 308218
rect 558804 307898 558986 308134
rect 559222 307898 559404 308134
rect 558804 272454 559404 307898
rect 558804 272218 558986 272454
rect 559222 272218 559404 272454
rect 558804 272134 559404 272218
rect 558804 271898 558986 272134
rect 559222 271898 559404 272134
rect 558804 236454 559404 271898
rect 558804 236218 558986 236454
rect 559222 236218 559404 236454
rect 558804 236134 559404 236218
rect 558804 235898 558986 236134
rect 559222 235898 559404 236134
rect 558804 200454 559404 235898
rect 558804 200218 558986 200454
rect 559222 200218 559404 200454
rect 558804 200134 559404 200218
rect 558804 199898 558986 200134
rect 559222 199898 559404 200134
rect 558804 164454 559404 199898
rect 558804 164218 558986 164454
rect 559222 164218 559404 164454
rect 558804 164134 559404 164218
rect 558804 163898 558986 164134
rect 559222 163898 559404 164134
rect 558804 128454 559404 163898
rect 558804 128218 558986 128454
rect 559222 128218 559404 128454
rect 558804 128134 559404 128218
rect 558804 127898 558986 128134
rect 559222 127898 559404 128134
rect 558804 92454 559404 127898
rect 558804 92218 558986 92454
rect 559222 92218 559404 92454
rect 558804 92134 559404 92218
rect 558804 91898 558986 92134
rect 559222 91898 559404 92134
rect 558804 56454 559404 91898
rect 558804 56218 558986 56454
rect 559222 56218 559404 56454
rect 558804 56134 559404 56218
rect 558804 55898 558986 56134
rect 559222 55898 559404 56134
rect 558804 20454 559404 55898
rect 558804 20218 558986 20454
rect 559222 20218 559404 20454
rect 558804 20134 559404 20218
rect 558804 19898 558986 20134
rect 559222 19898 559404 20134
rect 558804 -1286 559404 19898
rect 558804 -1522 558986 -1286
rect 559222 -1522 559404 -1286
rect 558804 -1606 559404 -1522
rect 558804 -1842 558986 -1606
rect 559222 -1842 559404 -1606
rect 558804 -1864 559404 -1842
rect 562404 672054 563004 707102
rect 562404 671818 562586 672054
rect 562822 671818 563004 672054
rect 562404 671734 563004 671818
rect 562404 671498 562586 671734
rect 562822 671498 563004 671734
rect 562404 636054 563004 671498
rect 562404 635818 562586 636054
rect 562822 635818 563004 636054
rect 562404 635734 563004 635818
rect 562404 635498 562586 635734
rect 562822 635498 563004 635734
rect 562404 600054 563004 635498
rect 562404 599818 562586 600054
rect 562822 599818 563004 600054
rect 562404 599734 563004 599818
rect 562404 599498 562586 599734
rect 562822 599498 563004 599734
rect 562404 564054 563004 599498
rect 562404 563818 562586 564054
rect 562822 563818 563004 564054
rect 562404 563734 563004 563818
rect 562404 563498 562586 563734
rect 562822 563498 563004 563734
rect 562404 528054 563004 563498
rect 562404 527818 562586 528054
rect 562822 527818 563004 528054
rect 562404 527734 563004 527818
rect 562404 527498 562586 527734
rect 562822 527498 563004 527734
rect 562404 492054 563004 527498
rect 562404 491818 562586 492054
rect 562822 491818 563004 492054
rect 562404 491734 563004 491818
rect 562404 491498 562586 491734
rect 562822 491498 563004 491734
rect 562404 456054 563004 491498
rect 562404 455818 562586 456054
rect 562822 455818 563004 456054
rect 562404 455734 563004 455818
rect 562404 455498 562586 455734
rect 562822 455498 563004 455734
rect 562404 420054 563004 455498
rect 562404 419818 562586 420054
rect 562822 419818 563004 420054
rect 562404 419734 563004 419818
rect 562404 419498 562586 419734
rect 562822 419498 563004 419734
rect 562404 384054 563004 419498
rect 562404 383818 562586 384054
rect 562822 383818 563004 384054
rect 562404 383734 563004 383818
rect 562404 383498 562586 383734
rect 562822 383498 563004 383734
rect 562404 348054 563004 383498
rect 562404 347818 562586 348054
rect 562822 347818 563004 348054
rect 562404 347734 563004 347818
rect 562404 347498 562586 347734
rect 562822 347498 563004 347734
rect 562404 312054 563004 347498
rect 562404 311818 562586 312054
rect 562822 311818 563004 312054
rect 562404 311734 563004 311818
rect 562404 311498 562586 311734
rect 562822 311498 563004 311734
rect 562404 276054 563004 311498
rect 562404 275818 562586 276054
rect 562822 275818 563004 276054
rect 562404 275734 563004 275818
rect 562404 275498 562586 275734
rect 562822 275498 563004 275734
rect 562404 240054 563004 275498
rect 562404 239818 562586 240054
rect 562822 239818 563004 240054
rect 562404 239734 563004 239818
rect 562404 239498 562586 239734
rect 562822 239498 563004 239734
rect 562404 204054 563004 239498
rect 562404 203818 562586 204054
rect 562822 203818 563004 204054
rect 562404 203734 563004 203818
rect 562404 203498 562586 203734
rect 562822 203498 563004 203734
rect 562404 168054 563004 203498
rect 562404 167818 562586 168054
rect 562822 167818 563004 168054
rect 562404 167734 563004 167818
rect 562404 167498 562586 167734
rect 562822 167498 563004 167734
rect 562404 132054 563004 167498
rect 562404 131818 562586 132054
rect 562822 131818 563004 132054
rect 562404 131734 563004 131818
rect 562404 131498 562586 131734
rect 562822 131498 563004 131734
rect 562404 96054 563004 131498
rect 562404 95818 562586 96054
rect 562822 95818 563004 96054
rect 562404 95734 563004 95818
rect 562404 95498 562586 95734
rect 562822 95498 563004 95734
rect 562404 60054 563004 95498
rect 562404 59818 562586 60054
rect 562822 59818 563004 60054
rect 562404 59734 563004 59818
rect 562404 59498 562586 59734
rect 562822 59498 563004 59734
rect 562404 24054 563004 59498
rect 562404 23818 562586 24054
rect 562822 23818 563004 24054
rect 562404 23734 563004 23818
rect 562404 23498 562586 23734
rect 562822 23498 563004 23734
rect 562404 -3166 563004 23498
rect 562404 -3402 562586 -3166
rect 562822 -3402 563004 -3166
rect 562404 -3486 563004 -3402
rect 562404 -3722 562586 -3486
rect 562822 -3722 563004 -3486
rect 562404 -3744 563004 -3722
rect 566004 675654 566604 708982
rect 566004 675418 566186 675654
rect 566422 675418 566604 675654
rect 566004 675334 566604 675418
rect 566004 675098 566186 675334
rect 566422 675098 566604 675334
rect 566004 639654 566604 675098
rect 566004 639418 566186 639654
rect 566422 639418 566604 639654
rect 566004 639334 566604 639418
rect 566004 639098 566186 639334
rect 566422 639098 566604 639334
rect 566004 603654 566604 639098
rect 566004 603418 566186 603654
rect 566422 603418 566604 603654
rect 566004 603334 566604 603418
rect 566004 603098 566186 603334
rect 566422 603098 566604 603334
rect 566004 567654 566604 603098
rect 566004 567418 566186 567654
rect 566422 567418 566604 567654
rect 566004 567334 566604 567418
rect 566004 567098 566186 567334
rect 566422 567098 566604 567334
rect 566004 531654 566604 567098
rect 566004 531418 566186 531654
rect 566422 531418 566604 531654
rect 566004 531334 566604 531418
rect 566004 531098 566186 531334
rect 566422 531098 566604 531334
rect 566004 495654 566604 531098
rect 566004 495418 566186 495654
rect 566422 495418 566604 495654
rect 566004 495334 566604 495418
rect 566004 495098 566186 495334
rect 566422 495098 566604 495334
rect 566004 459654 566604 495098
rect 566004 459418 566186 459654
rect 566422 459418 566604 459654
rect 566004 459334 566604 459418
rect 566004 459098 566186 459334
rect 566422 459098 566604 459334
rect 566004 423654 566604 459098
rect 566004 423418 566186 423654
rect 566422 423418 566604 423654
rect 566004 423334 566604 423418
rect 566004 423098 566186 423334
rect 566422 423098 566604 423334
rect 566004 387654 566604 423098
rect 566004 387418 566186 387654
rect 566422 387418 566604 387654
rect 566004 387334 566604 387418
rect 566004 387098 566186 387334
rect 566422 387098 566604 387334
rect 566004 351654 566604 387098
rect 566004 351418 566186 351654
rect 566422 351418 566604 351654
rect 566004 351334 566604 351418
rect 566004 351098 566186 351334
rect 566422 351098 566604 351334
rect 566004 315654 566604 351098
rect 566004 315418 566186 315654
rect 566422 315418 566604 315654
rect 566004 315334 566604 315418
rect 566004 315098 566186 315334
rect 566422 315098 566604 315334
rect 566004 279654 566604 315098
rect 566004 279418 566186 279654
rect 566422 279418 566604 279654
rect 566004 279334 566604 279418
rect 566004 279098 566186 279334
rect 566422 279098 566604 279334
rect 566004 243654 566604 279098
rect 566004 243418 566186 243654
rect 566422 243418 566604 243654
rect 566004 243334 566604 243418
rect 566004 243098 566186 243334
rect 566422 243098 566604 243334
rect 566004 207654 566604 243098
rect 566004 207418 566186 207654
rect 566422 207418 566604 207654
rect 566004 207334 566604 207418
rect 566004 207098 566186 207334
rect 566422 207098 566604 207334
rect 566004 171654 566604 207098
rect 566004 171418 566186 171654
rect 566422 171418 566604 171654
rect 566004 171334 566604 171418
rect 566004 171098 566186 171334
rect 566422 171098 566604 171334
rect 566004 135654 566604 171098
rect 566004 135418 566186 135654
rect 566422 135418 566604 135654
rect 566004 135334 566604 135418
rect 566004 135098 566186 135334
rect 566422 135098 566604 135334
rect 566004 99654 566604 135098
rect 566004 99418 566186 99654
rect 566422 99418 566604 99654
rect 566004 99334 566604 99418
rect 566004 99098 566186 99334
rect 566422 99098 566604 99334
rect 566004 63654 566604 99098
rect 566004 63418 566186 63654
rect 566422 63418 566604 63654
rect 566004 63334 566604 63418
rect 566004 63098 566186 63334
rect 566422 63098 566604 63334
rect 566004 27654 566604 63098
rect 566004 27418 566186 27654
rect 566422 27418 566604 27654
rect 566004 27334 566604 27418
rect 566004 27098 566186 27334
rect 566422 27098 566604 27334
rect 566004 -5046 566604 27098
rect 566004 -5282 566186 -5046
rect 566422 -5282 566604 -5046
rect 566004 -5366 566604 -5282
rect 566004 -5602 566186 -5366
rect 566422 -5602 566604 -5366
rect 566004 -5624 566604 -5602
rect 569604 679254 570204 710862
rect 591900 711418 592500 711440
rect 591900 711182 592082 711418
rect 592318 711182 592500 711418
rect 591900 711098 592500 711182
rect 591900 710862 592082 711098
rect 592318 710862 592500 711098
rect 590960 710478 591560 710500
rect 590960 710242 591142 710478
rect 591378 710242 591560 710478
rect 590960 710158 591560 710242
rect 590960 709922 591142 710158
rect 591378 709922 591560 710158
rect 590020 709538 590620 709560
rect 590020 709302 590202 709538
rect 590438 709302 590620 709538
rect 590020 709218 590620 709302
rect 590020 708982 590202 709218
rect 590438 708982 590620 709218
rect 589080 708598 589680 708620
rect 589080 708362 589262 708598
rect 589498 708362 589680 708598
rect 589080 708278 589680 708362
rect 589080 708042 589262 708278
rect 589498 708042 589680 708278
rect 580404 706718 581004 707680
rect 588140 707658 588740 707680
rect 588140 707422 588322 707658
rect 588558 707422 588740 707658
rect 588140 707338 588740 707422
rect 588140 707102 588322 707338
rect 588558 707102 588740 707338
rect 580404 706482 580586 706718
rect 580822 706482 581004 706718
rect 580404 706398 581004 706482
rect 580404 706162 580586 706398
rect 580822 706162 581004 706398
rect 569604 679018 569786 679254
rect 570022 679018 570204 679254
rect 569604 678934 570204 679018
rect 569604 678698 569786 678934
rect 570022 678698 570204 678934
rect 569604 643254 570204 678698
rect 569604 643018 569786 643254
rect 570022 643018 570204 643254
rect 569604 642934 570204 643018
rect 569604 642698 569786 642934
rect 570022 642698 570204 642934
rect 569604 607254 570204 642698
rect 569604 607018 569786 607254
rect 570022 607018 570204 607254
rect 569604 606934 570204 607018
rect 569604 606698 569786 606934
rect 570022 606698 570204 606934
rect 569604 571254 570204 606698
rect 569604 571018 569786 571254
rect 570022 571018 570204 571254
rect 569604 570934 570204 571018
rect 569604 570698 569786 570934
rect 570022 570698 570204 570934
rect 569604 535254 570204 570698
rect 569604 535018 569786 535254
rect 570022 535018 570204 535254
rect 569604 534934 570204 535018
rect 569604 534698 569786 534934
rect 570022 534698 570204 534934
rect 569604 499254 570204 534698
rect 569604 499018 569786 499254
rect 570022 499018 570204 499254
rect 569604 498934 570204 499018
rect 569604 498698 569786 498934
rect 570022 498698 570204 498934
rect 569604 463254 570204 498698
rect 569604 463018 569786 463254
rect 570022 463018 570204 463254
rect 569604 462934 570204 463018
rect 569604 462698 569786 462934
rect 570022 462698 570204 462934
rect 569604 427254 570204 462698
rect 569604 427018 569786 427254
rect 570022 427018 570204 427254
rect 569604 426934 570204 427018
rect 569604 426698 569786 426934
rect 570022 426698 570204 426934
rect 569604 391254 570204 426698
rect 569604 391018 569786 391254
rect 570022 391018 570204 391254
rect 569604 390934 570204 391018
rect 569604 390698 569786 390934
rect 570022 390698 570204 390934
rect 569604 355254 570204 390698
rect 569604 355018 569786 355254
rect 570022 355018 570204 355254
rect 569604 354934 570204 355018
rect 569604 354698 569786 354934
rect 570022 354698 570204 354934
rect 569604 319254 570204 354698
rect 569604 319018 569786 319254
rect 570022 319018 570204 319254
rect 569604 318934 570204 319018
rect 569604 318698 569786 318934
rect 570022 318698 570204 318934
rect 569604 283254 570204 318698
rect 569604 283018 569786 283254
rect 570022 283018 570204 283254
rect 569604 282934 570204 283018
rect 569604 282698 569786 282934
rect 570022 282698 570204 282934
rect 569604 247254 570204 282698
rect 569604 247018 569786 247254
rect 570022 247018 570204 247254
rect 569604 246934 570204 247018
rect 569604 246698 569786 246934
rect 570022 246698 570204 246934
rect 569604 211254 570204 246698
rect 569604 211018 569786 211254
rect 570022 211018 570204 211254
rect 569604 210934 570204 211018
rect 569604 210698 569786 210934
rect 570022 210698 570204 210934
rect 569604 175254 570204 210698
rect 569604 175018 569786 175254
rect 570022 175018 570204 175254
rect 569604 174934 570204 175018
rect 569604 174698 569786 174934
rect 570022 174698 570204 174934
rect 569604 139254 570204 174698
rect 569604 139018 569786 139254
rect 570022 139018 570204 139254
rect 569604 138934 570204 139018
rect 569604 138698 569786 138934
rect 570022 138698 570204 138934
rect 569604 103254 570204 138698
rect 569604 103018 569786 103254
rect 570022 103018 570204 103254
rect 569604 102934 570204 103018
rect 569604 102698 569786 102934
rect 570022 102698 570204 102934
rect 569604 67254 570204 102698
rect 569604 67018 569786 67254
rect 570022 67018 570204 67254
rect 569604 66934 570204 67018
rect 569604 66698 569786 66934
rect 570022 66698 570204 66934
rect 569604 31254 570204 66698
rect 569604 31018 569786 31254
rect 570022 31018 570204 31254
rect 569604 30934 570204 31018
rect 569604 30698 569786 30934
rect 570022 30698 570204 30934
rect 551604 -6222 551786 -5986
rect 552022 -6222 552204 -5986
rect 551604 -6306 552204 -6222
rect 551604 -6542 551786 -6306
rect 552022 -6542 552204 -6306
rect 551604 -7504 552204 -6542
rect 569604 -6926 570204 30698
rect 576804 704838 577404 705800
rect 576804 704602 576986 704838
rect 577222 704602 577404 704838
rect 576804 704518 577404 704602
rect 576804 704282 576986 704518
rect 577222 704282 577404 704518
rect 576804 686454 577404 704282
rect 576804 686218 576986 686454
rect 577222 686218 577404 686454
rect 576804 686134 577404 686218
rect 576804 685898 576986 686134
rect 577222 685898 577404 686134
rect 576804 650454 577404 685898
rect 576804 650218 576986 650454
rect 577222 650218 577404 650454
rect 576804 650134 577404 650218
rect 576804 649898 576986 650134
rect 577222 649898 577404 650134
rect 576804 614454 577404 649898
rect 576804 614218 576986 614454
rect 577222 614218 577404 614454
rect 576804 614134 577404 614218
rect 576804 613898 576986 614134
rect 577222 613898 577404 614134
rect 576804 578454 577404 613898
rect 576804 578218 576986 578454
rect 577222 578218 577404 578454
rect 576804 578134 577404 578218
rect 576804 577898 576986 578134
rect 577222 577898 577404 578134
rect 576804 542454 577404 577898
rect 576804 542218 576986 542454
rect 577222 542218 577404 542454
rect 576804 542134 577404 542218
rect 576804 541898 576986 542134
rect 577222 541898 577404 542134
rect 576804 506454 577404 541898
rect 576804 506218 576986 506454
rect 577222 506218 577404 506454
rect 576804 506134 577404 506218
rect 576804 505898 576986 506134
rect 577222 505898 577404 506134
rect 576804 470454 577404 505898
rect 576804 470218 576986 470454
rect 577222 470218 577404 470454
rect 576804 470134 577404 470218
rect 576804 469898 576986 470134
rect 577222 469898 577404 470134
rect 576804 434454 577404 469898
rect 576804 434218 576986 434454
rect 577222 434218 577404 434454
rect 576804 434134 577404 434218
rect 576804 433898 576986 434134
rect 577222 433898 577404 434134
rect 576804 398454 577404 433898
rect 576804 398218 576986 398454
rect 577222 398218 577404 398454
rect 576804 398134 577404 398218
rect 576804 397898 576986 398134
rect 577222 397898 577404 398134
rect 576804 362454 577404 397898
rect 576804 362218 576986 362454
rect 577222 362218 577404 362454
rect 576804 362134 577404 362218
rect 576804 361898 576986 362134
rect 577222 361898 577404 362134
rect 576804 326454 577404 361898
rect 576804 326218 576986 326454
rect 577222 326218 577404 326454
rect 576804 326134 577404 326218
rect 576804 325898 576986 326134
rect 577222 325898 577404 326134
rect 576804 290454 577404 325898
rect 576804 290218 576986 290454
rect 577222 290218 577404 290454
rect 576804 290134 577404 290218
rect 576804 289898 576986 290134
rect 577222 289898 577404 290134
rect 576804 254454 577404 289898
rect 576804 254218 576986 254454
rect 577222 254218 577404 254454
rect 576804 254134 577404 254218
rect 576804 253898 576986 254134
rect 577222 253898 577404 254134
rect 576804 218454 577404 253898
rect 576804 218218 576986 218454
rect 577222 218218 577404 218454
rect 576804 218134 577404 218218
rect 576804 217898 576986 218134
rect 577222 217898 577404 218134
rect 576804 182454 577404 217898
rect 576804 182218 576986 182454
rect 577222 182218 577404 182454
rect 576804 182134 577404 182218
rect 576804 181898 576986 182134
rect 577222 181898 577404 182134
rect 576804 146454 577404 181898
rect 576804 146218 576986 146454
rect 577222 146218 577404 146454
rect 576804 146134 577404 146218
rect 576804 145898 576986 146134
rect 577222 145898 577404 146134
rect 576804 110454 577404 145898
rect 576804 110218 576986 110454
rect 577222 110218 577404 110454
rect 576804 110134 577404 110218
rect 576804 109898 576986 110134
rect 577222 109898 577404 110134
rect 576804 74454 577404 109898
rect 576804 74218 576986 74454
rect 577222 74218 577404 74454
rect 576804 74134 577404 74218
rect 576804 73898 576986 74134
rect 577222 73898 577404 74134
rect 576804 38454 577404 73898
rect 576804 38218 576986 38454
rect 577222 38218 577404 38454
rect 576804 38134 577404 38218
rect 576804 37898 576986 38134
rect 577222 37898 577404 38134
rect 576804 2454 577404 37898
rect 576804 2218 576986 2454
rect 577222 2218 577404 2454
rect 576804 2134 577404 2218
rect 576804 1898 576986 2134
rect 577222 1898 577404 2134
rect 576804 -346 577404 1898
rect 576804 -582 576986 -346
rect 577222 -582 577404 -346
rect 576804 -666 577404 -582
rect 576804 -902 576986 -666
rect 577222 -902 577404 -666
rect 576804 -1864 577404 -902
rect 580404 690054 581004 706162
rect 587200 706718 587800 706740
rect 587200 706482 587382 706718
rect 587618 706482 587800 706718
rect 587200 706398 587800 706482
rect 587200 706162 587382 706398
rect 587618 706162 587800 706398
rect 586260 705778 586860 705800
rect 586260 705542 586442 705778
rect 586678 705542 586860 705778
rect 586260 705458 586860 705542
rect 586260 705222 586442 705458
rect 586678 705222 586860 705458
rect 580404 689818 580586 690054
rect 580822 689818 581004 690054
rect 580404 689734 581004 689818
rect 580404 689498 580586 689734
rect 580822 689498 581004 689734
rect 580404 654054 581004 689498
rect 580404 653818 580586 654054
rect 580822 653818 581004 654054
rect 580404 653734 581004 653818
rect 580404 653498 580586 653734
rect 580822 653498 581004 653734
rect 580404 618054 581004 653498
rect 580404 617818 580586 618054
rect 580822 617818 581004 618054
rect 580404 617734 581004 617818
rect 580404 617498 580586 617734
rect 580822 617498 581004 617734
rect 580404 582054 581004 617498
rect 580404 581818 580586 582054
rect 580822 581818 581004 582054
rect 580404 581734 581004 581818
rect 580404 581498 580586 581734
rect 580822 581498 581004 581734
rect 580404 546054 581004 581498
rect 580404 545818 580586 546054
rect 580822 545818 581004 546054
rect 580404 545734 581004 545818
rect 580404 545498 580586 545734
rect 580822 545498 581004 545734
rect 580404 510054 581004 545498
rect 580404 509818 580586 510054
rect 580822 509818 581004 510054
rect 580404 509734 581004 509818
rect 580404 509498 580586 509734
rect 580822 509498 581004 509734
rect 580404 474054 581004 509498
rect 580404 473818 580586 474054
rect 580822 473818 581004 474054
rect 580404 473734 581004 473818
rect 580404 473498 580586 473734
rect 580822 473498 581004 473734
rect 580404 438054 581004 473498
rect 580404 437818 580586 438054
rect 580822 437818 581004 438054
rect 580404 437734 581004 437818
rect 580404 437498 580586 437734
rect 580822 437498 581004 437734
rect 580404 402054 581004 437498
rect 580404 401818 580586 402054
rect 580822 401818 581004 402054
rect 580404 401734 581004 401818
rect 580404 401498 580586 401734
rect 580822 401498 581004 401734
rect 580404 366054 581004 401498
rect 580404 365818 580586 366054
rect 580822 365818 581004 366054
rect 580404 365734 581004 365818
rect 580404 365498 580586 365734
rect 580822 365498 581004 365734
rect 580404 330054 581004 365498
rect 580404 329818 580586 330054
rect 580822 329818 581004 330054
rect 580404 329734 581004 329818
rect 580404 329498 580586 329734
rect 580822 329498 581004 329734
rect 580404 294054 581004 329498
rect 580404 293818 580586 294054
rect 580822 293818 581004 294054
rect 580404 293734 581004 293818
rect 580404 293498 580586 293734
rect 580822 293498 581004 293734
rect 580404 258054 581004 293498
rect 580404 257818 580586 258054
rect 580822 257818 581004 258054
rect 580404 257734 581004 257818
rect 580404 257498 580586 257734
rect 580822 257498 581004 257734
rect 580404 222054 581004 257498
rect 580404 221818 580586 222054
rect 580822 221818 581004 222054
rect 580404 221734 581004 221818
rect 580404 221498 580586 221734
rect 580822 221498 581004 221734
rect 580404 186054 581004 221498
rect 580404 185818 580586 186054
rect 580822 185818 581004 186054
rect 580404 185734 581004 185818
rect 580404 185498 580586 185734
rect 580822 185498 581004 185734
rect 580404 150054 581004 185498
rect 580404 149818 580586 150054
rect 580822 149818 581004 150054
rect 580404 149734 581004 149818
rect 580404 149498 580586 149734
rect 580822 149498 581004 149734
rect 580404 114054 581004 149498
rect 580404 113818 580586 114054
rect 580822 113818 581004 114054
rect 580404 113734 581004 113818
rect 580404 113498 580586 113734
rect 580822 113498 581004 113734
rect 580404 78054 581004 113498
rect 580404 77818 580586 78054
rect 580822 77818 581004 78054
rect 580404 77734 581004 77818
rect 580404 77498 580586 77734
rect 580822 77498 581004 77734
rect 580404 42054 581004 77498
rect 580404 41818 580586 42054
rect 580822 41818 581004 42054
rect 580404 41734 581004 41818
rect 580404 41498 580586 41734
rect 580822 41498 581004 41734
rect 580404 6054 581004 41498
rect 580404 5818 580586 6054
rect 580822 5818 581004 6054
rect 580404 5734 581004 5818
rect 580404 5498 580586 5734
rect 580822 5498 581004 5734
rect 580404 -2226 581004 5498
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 585320 686454 585920 704282
rect 585320 686218 585502 686454
rect 585738 686218 585920 686454
rect 585320 686134 585920 686218
rect 585320 685898 585502 686134
rect 585738 685898 585920 686134
rect 585320 650454 585920 685898
rect 585320 650218 585502 650454
rect 585738 650218 585920 650454
rect 585320 650134 585920 650218
rect 585320 649898 585502 650134
rect 585738 649898 585920 650134
rect 585320 614454 585920 649898
rect 585320 614218 585502 614454
rect 585738 614218 585920 614454
rect 585320 614134 585920 614218
rect 585320 613898 585502 614134
rect 585738 613898 585920 614134
rect 585320 578454 585920 613898
rect 585320 578218 585502 578454
rect 585738 578218 585920 578454
rect 585320 578134 585920 578218
rect 585320 577898 585502 578134
rect 585738 577898 585920 578134
rect 585320 542454 585920 577898
rect 585320 542218 585502 542454
rect 585738 542218 585920 542454
rect 585320 542134 585920 542218
rect 585320 541898 585502 542134
rect 585738 541898 585920 542134
rect 585320 506454 585920 541898
rect 585320 506218 585502 506454
rect 585738 506218 585920 506454
rect 585320 506134 585920 506218
rect 585320 505898 585502 506134
rect 585738 505898 585920 506134
rect 585320 470454 585920 505898
rect 585320 470218 585502 470454
rect 585738 470218 585920 470454
rect 585320 470134 585920 470218
rect 585320 469898 585502 470134
rect 585738 469898 585920 470134
rect 585320 434454 585920 469898
rect 585320 434218 585502 434454
rect 585738 434218 585920 434454
rect 585320 434134 585920 434218
rect 585320 433898 585502 434134
rect 585738 433898 585920 434134
rect 585320 398454 585920 433898
rect 585320 398218 585502 398454
rect 585738 398218 585920 398454
rect 585320 398134 585920 398218
rect 585320 397898 585502 398134
rect 585738 397898 585920 398134
rect 585320 362454 585920 397898
rect 585320 362218 585502 362454
rect 585738 362218 585920 362454
rect 585320 362134 585920 362218
rect 585320 361898 585502 362134
rect 585738 361898 585920 362134
rect 585320 326454 585920 361898
rect 585320 326218 585502 326454
rect 585738 326218 585920 326454
rect 585320 326134 585920 326218
rect 585320 325898 585502 326134
rect 585738 325898 585920 326134
rect 585320 290454 585920 325898
rect 585320 290218 585502 290454
rect 585738 290218 585920 290454
rect 585320 290134 585920 290218
rect 585320 289898 585502 290134
rect 585738 289898 585920 290134
rect 585320 254454 585920 289898
rect 585320 254218 585502 254454
rect 585738 254218 585920 254454
rect 585320 254134 585920 254218
rect 585320 253898 585502 254134
rect 585738 253898 585920 254134
rect 585320 218454 585920 253898
rect 585320 218218 585502 218454
rect 585738 218218 585920 218454
rect 585320 218134 585920 218218
rect 585320 217898 585502 218134
rect 585738 217898 585920 218134
rect 585320 182454 585920 217898
rect 585320 182218 585502 182454
rect 585738 182218 585920 182454
rect 585320 182134 585920 182218
rect 585320 181898 585502 182134
rect 585738 181898 585920 182134
rect 585320 146454 585920 181898
rect 585320 146218 585502 146454
rect 585738 146218 585920 146454
rect 585320 146134 585920 146218
rect 585320 145898 585502 146134
rect 585738 145898 585920 146134
rect 585320 110454 585920 145898
rect 585320 110218 585502 110454
rect 585738 110218 585920 110454
rect 585320 110134 585920 110218
rect 585320 109898 585502 110134
rect 585738 109898 585920 110134
rect 585320 74454 585920 109898
rect 585320 74218 585502 74454
rect 585738 74218 585920 74454
rect 585320 74134 585920 74218
rect 585320 73898 585502 74134
rect 585738 73898 585920 74134
rect 585320 38454 585920 73898
rect 585320 38218 585502 38454
rect 585738 38218 585920 38454
rect 585320 38134 585920 38218
rect 585320 37898 585502 38134
rect 585738 37898 585920 38134
rect 585320 2454 585920 37898
rect 585320 2218 585502 2454
rect 585738 2218 585920 2454
rect 585320 2134 585920 2218
rect 585320 1898 585502 2134
rect 585738 1898 585920 2134
rect 585320 -346 585920 1898
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586260 668454 586860 705222
rect 586260 668218 586442 668454
rect 586678 668218 586860 668454
rect 586260 668134 586860 668218
rect 586260 667898 586442 668134
rect 586678 667898 586860 668134
rect 586260 632454 586860 667898
rect 586260 632218 586442 632454
rect 586678 632218 586860 632454
rect 586260 632134 586860 632218
rect 586260 631898 586442 632134
rect 586678 631898 586860 632134
rect 586260 596454 586860 631898
rect 586260 596218 586442 596454
rect 586678 596218 586860 596454
rect 586260 596134 586860 596218
rect 586260 595898 586442 596134
rect 586678 595898 586860 596134
rect 586260 560454 586860 595898
rect 586260 560218 586442 560454
rect 586678 560218 586860 560454
rect 586260 560134 586860 560218
rect 586260 559898 586442 560134
rect 586678 559898 586860 560134
rect 586260 524454 586860 559898
rect 586260 524218 586442 524454
rect 586678 524218 586860 524454
rect 586260 524134 586860 524218
rect 586260 523898 586442 524134
rect 586678 523898 586860 524134
rect 586260 488454 586860 523898
rect 586260 488218 586442 488454
rect 586678 488218 586860 488454
rect 586260 488134 586860 488218
rect 586260 487898 586442 488134
rect 586678 487898 586860 488134
rect 586260 452454 586860 487898
rect 586260 452218 586442 452454
rect 586678 452218 586860 452454
rect 586260 452134 586860 452218
rect 586260 451898 586442 452134
rect 586678 451898 586860 452134
rect 586260 416454 586860 451898
rect 586260 416218 586442 416454
rect 586678 416218 586860 416454
rect 586260 416134 586860 416218
rect 586260 415898 586442 416134
rect 586678 415898 586860 416134
rect 586260 380454 586860 415898
rect 586260 380218 586442 380454
rect 586678 380218 586860 380454
rect 586260 380134 586860 380218
rect 586260 379898 586442 380134
rect 586678 379898 586860 380134
rect 586260 344454 586860 379898
rect 586260 344218 586442 344454
rect 586678 344218 586860 344454
rect 586260 344134 586860 344218
rect 586260 343898 586442 344134
rect 586678 343898 586860 344134
rect 586260 308454 586860 343898
rect 586260 308218 586442 308454
rect 586678 308218 586860 308454
rect 586260 308134 586860 308218
rect 586260 307898 586442 308134
rect 586678 307898 586860 308134
rect 586260 272454 586860 307898
rect 586260 272218 586442 272454
rect 586678 272218 586860 272454
rect 586260 272134 586860 272218
rect 586260 271898 586442 272134
rect 586678 271898 586860 272134
rect 586260 236454 586860 271898
rect 586260 236218 586442 236454
rect 586678 236218 586860 236454
rect 586260 236134 586860 236218
rect 586260 235898 586442 236134
rect 586678 235898 586860 236134
rect 586260 200454 586860 235898
rect 586260 200218 586442 200454
rect 586678 200218 586860 200454
rect 586260 200134 586860 200218
rect 586260 199898 586442 200134
rect 586678 199898 586860 200134
rect 586260 164454 586860 199898
rect 586260 164218 586442 164454
rect 586678 164218 586860 164454
rect 586260 164134 586860 164218
rect 586260 163898 586442 164134
rect 586678 163898 586860 164134
rect 586260 128454 586860 163898
rect 586260 128218 586442 128454
rect 586678 128218 586860 128454
rect 586260 128134 586860 128218
rect 586260 127898 586442 128134
rect 586678 127898 586860 128134
rect 586260 92454 586860 127898
rect 586260 92218 586442 92454
rect 586678 92218 586860 92454
rect 586260 92134 586860 92218
rect 586260 91898 586442 92134
rect 586678 91898 586860 92134
rect 586260 56454 586860 91898
rect 586260 56218 586442 56454
rect 586678 56218 586860 56454
rect 586260 56134 586860 56218
rect 586260 55898 586442 56134
rect 586678 55898 586860 56134
rect 586260 20454 586860 55898
rect 586260 20218 586442 20454
rect 586678 20218 586860 20454
rect 586260 20134 586860 20218
rect 586260 19898 586442 20134
rect 586678 19898 586860 20134
rect 586260 -1286 586860 19898
rect 586260 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect 586260 -1606 586860 -1522
rect 586260 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect 586260 -1864 586860 -1842
rect 587200 690054 587800 706162
rect 587200 689818 587382 690054
rect 587618 689818 587800 690054
rect 587200 689734 587800 689818
rect 587200 689498 587382 689734
rect 587618 689498 587800 689734
rect 587200 654054 587800 689498
rect 587200 653818 587382 654054
rect 587618 653818 587800 654054
rect 587200 653734 587800 653818
rect 587200 653498 587382 653734
rect 587618 653498 587800 653734
rect 587200 618054 587800 653498
rect 587200 617818 587382 618054
rect 587618 617818 587800 618054
rect 587200 617734 587800 617818
rect 587200 617498 587382 617734
rect 587618 617498 587800 617734
rect 587200 582054 587800 617498
rect 587200 581818 587382 582054
rect 587618 581818 587800 582054
rect 587200 581734 587800 581818
rect 587200 581498 587382 581734
rect 587618 581498 587800 581734
rect 587200 546054 587800 581498
rect 587200 545818 587382 546054
rect 587618 545818 587800 546054
rect 587200 545734 587800 545818
rect 587200 545498 587382 545734
rect 587618 545498 587800 545734
rect 587200 510054 587800 545498
rect 587200 509818 587382 510054
rect 587618 509818 587800 510054
rect 587200 509734 587800 509818
rect 587200 509498 587382 509734
rect 587618 509498 587800 509734
rect 587200 474054 587800 509498
rect 587200 473818 587382 474054
rect 587618 473818 587800 474054
rect 587200 473734 587800 473818
rect 587200 473498 587382 473734
rect 587618 473498 587800 473734
rect 587200 438054 587800 473498
rect 587200 437818 587382 438054
rect 587618 437818 587800 438054
rect 587200 437734 587800 437818
rect 587200 437498 587382 437734
rect 587618 437498 587800 437734
rect 587200 402054 587800 437498
rect 587200 401818 587382 402054
rect 587618 401818 587800 402054
rect 587200 401734 587800 401818
rect 587200 401498 587382 401734
rect 587618 401498 587800 401734
rect 587200 366054 587800 401498
rect 587200 365818 587382 366054
rect 587618 365818 587800 366054
rect 587200 365734 587800 365818
rect 587200 365498 587382 365734
rect 587618 365498 587800 365734
rect 587200 330054 587800 365498
rect 587200 329818 587382 330054
rect 587618 329818 587800 330054
rect 587200 329734 587800 329818
rect 587200 329498 587382 329734
rect 587618 329498 587800 329734
rect 587200 294054 587800 329498
rect 587200 293818 587382 294054
rect 587618 293818 587800 294054
rect 587200 293734 587800 293818
rect 587200 293498 587382 293734
rect 587618 293498 587800 293734
rect 587200 258054 587800 293498
rect 587200 257818 587382 258054
rect 587618 257818 587800 258054
rect 587200 257734 587800 257818
rect 587200 257498 587382 257734
rect 587618 257498 587800 257734
rect 587200 222054 587800 257498
rect 587200 221818 587382 222054
rect 587618 221818 587800 222054
rect 587200 221734 587800 221818
rect 587200 221498 587382 221734
rect 587618 221498 587800 221734
rect 587200 186054 587800 221498
rect 587200 185818 587382 186054
rect 587618 185818 587800 186054
rect 587200 185734 587800 185818
rect 587200 185498 587382 185734
rect 587618 185498 587800 185734
rect 587200 150054 587800 185498
rect 587200 149818 587382 150054
rect 587618 149818 587800 150054
rect 587200 149734 587800 149818
rect 587200 149498 587382 149734
rect 587618 149498 587800 149734
rect 587200 114054 587800 149498
rect 587200 113818 587382 114054
rect 587618 113818 587800 114054
rect 587200 113734 587800 113818
rect 587200 113498 587382 113734
rect 587618 113498 587800 113734
rect 587200 78054 587800 113498
rect 587200 77818 587382 78054
rect 587618 77818 587800 78054
rect 587200 77734 587800 77818
rect 587200 77498 587382 77734
rect 587618 77498 587800 77734
rect 587200 42054 587800 77498
rect 587200 41818 587382 42054
rect 587618 41818 587800 42054
rect 587200 41734 587800 41818
rect 587200 41498 587382 41734
rect 587618 41498 587800 41734
rect 587200 6054 587800 41498
rect 587200 5818 587382 6054
rect 587618 5818 587800 6054
rect 587200 5734 587800 5818
rect 587200 5498 587382 5734
rect 587618 5498 587800 5734
rect 580404 -2462 580586 -2226
rect 580822 -2462 581004 -2226
rect 580404 -2546 581004 -2462
rect 580404 -2782 580586 -2546
rect 580822 -2782 581004 -2546
rect 580404 -3744 581004 -2782
rect 587200 -2226 587800 5498
rect 587200 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect 587200 -2546 587800 -2462
rect 587200 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect 587200 -2804 587800 -2782
rect 588140 672054 588740 707102
rect 588140 671818 588322 672054
rect 588558 671818 588740 672054
rect 588140 671734 588740 671818
rect 588140 671498 588322 671734
rect 588558 671498 588740 671734
rect 588140 636054 588740 671498
rect 588140 635818 588322 636054
rect 588558 635818 588740 636054
rect 588140 635734 588740 635818
rect 588140 635498 588322 635734
rect 588558 635498 588740 635734
rect 588140 600054 588740 635498
rect 588140 599818 588322 600054
rect 588558 599818 588740 600054
rect 588140 599734 588740 599818
rect 588140 599498 588322 599734
rect 588558 599498 588740 599734
rect 588140 564054 588740 599498
rect 588140 563818 588322 564054
rect 588558 563818 588740 564054
rect 588140 563734 588740 563818
rect 588140 563498 588322 563734
rect 588558 563498 588740 563734
rect 588140 528054 588740 563498
rect 588140 527818 588322 528054
rect 588558 527818 588740 528054
rect 588140 527734 588740 527818
rect 588140 527498 588322 527734
rect 588558 527498 588740 527734
rect 588140 492054 588740 527498
rect 588140 491818 588322 492054
rect 588558 491818 588740 492054
rect 588140 491734 588740 491818
rect 588140 491498 588322 491734
rect 588558 491498 588740 491734
rect 588140 456054 588740 491498
rect 588140 455818 588322 456054
rect 588558 455818 588740 456054
rect 588140 455734 588740 455818
rect 588140 455498 588322 455734
rect 588558 455498 588740 455734
rect 588140 420054 588740 455498
rect 588140 419818 588322 420054
rect 588558 419818 588740 420054
rect 588140 419734 588740 419818
rect 588140 419498 588322 419734
rect 588558 419498 588740 419734
rect 588140 384054 588740 419498
rect 588140 383818 588322 384054
rect 588558 383818 588740 384054
rect 588140 383734 588740 383818
rect 588140 383498 588322 383734
rect 588558 383498 588740 383734
rect 588140 348054 588740 383498
rect 588140 347818 588322 348054
rect 588558 347818 588740 348054
rect 588140 347734 588740 347818
rect 588140 347498 588322 347734
rect 588558 347498 588740 347734
rect 588140 312054 588740 347498
rect 588140 311818 588322 312054
rect 588558 311818 588740 312054
rect 588140 311734 588740 311818
rect 588140 311498 588322 311734
rect 588558 311498 588740 311734
rect 588140 276054 588740 311498
rect 588140 275818 588322 276054
rect 588558 275818 588740 276054
rect 588140 275734 588740 275818
rect 588140 275498 588322 275734
rect 588558 275498 588740 275734
rect 588140 240054 588740 275498
rect 588140 239818 588322 240054
rect 588558 239818 588740 240054
rect 588140 239734 588740 239818
rect 588140 239498 588322 239734
rect 588558 239498 588740 239734
rect 588140 204054 588740 239498
rect 588140 203818 588322 204054
rect 588558 203818 588740 204054
rect 588140 203734 588740 203818
rect 588140 203498 588322 203734
rect 588558 203498 588740 203734
rect 588140 168054 588740 203498
rect 588140 167818 588322 168054
rect 588558 167818 588740 168054
rect 588140 167734 588740 167818
rect 588140 167498 588322 167734
rect 588558 167498 588740 167734
rect 588140 132054 588740 167498
rect 588140 131818 588322 132054
rect 588558 131818 588740 132054
rect 588140 131734 588740 131818
rect 588140 131498 588322 131734
rect 588558 131498 588740 131734
rect 588140 96054 588740 131498
rect 588140 95818 588322 96054
rect 588558 95818 588740 96054
rect 588140 95734 588740 95818
rect 588140 95498 588322 95734
rect 588558 95498 588740 95734
rect 588140 60054 588740 95498
rect 588140 59818 588322 60054
rect 588558 59818 588740 60054
rect 588140 59734 588740 59818
rect 588140 59498 588322 59734
rect 588558 59498 588740 59734
rect 588140 24054 588740 59498
rect 588140 23818 588322 24054
rect 588558 23818 588740 24054
rect 588140 23734 588740 23818
rect 588140 23498 588322 23734
rect 588558 23498 588740 23734
rect 588140 -3166 588740 23498
rect 588140 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect 588140 -3486 588740 -3402
rect 588140 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect 588140 -3744 588740 -3722
rect 589080 693654 589680 708042
rect 589080 693418 589262 693654
rect 589498 693418 589680 693654
rect 589080 693334 589680 693418
rect 589080 693098 589262 693334
rect 589498 693098 589680 693334
rect 589080 657654 589680 693098
rect 589080 657418 589262 657654
rect 589498 657418 589680 657654
rect 589080 657334 589680 657418
rect 589080 657098 589262 657334
rect 589498 657098 589680 657334
rect 589080 621654 589680 657098
rect 589080 621418 589262 621654
rect 589498 621418 589680 621654
rect 589080 621334 589680 621418
rect 589080 621098 589262 621334
rect 589498 621098 589680 621334
rect 589080 585654 589680 621098
rect 589080 585418 589262 585654
rect 589498 585418 589680 585654
rect 589080 585334 589680 585418
rect 589080 585098 589262 585334
rect 589498 585098 589680 585334
rect 589080 549654 589680 585098
rect 589080 549418 589262 549654
rect 589498 549418 589680 549654
rect 589080 549334 589680 549418
rect 589080 549098 589262 549334
rect 589498 549098 589680 549334
rect 589080 513654 589680 549098
rect 589080 513418 589262 513654
rect 589498 513418 589680 513654
rect 589080 513334 589680 513418
rect 589080 513098 589262 513334
rect 589498 513098 589680 513334
rect 589080 477654 589680 513098
rect 589080 477418 589262 477654
rect 589498 477418 589680 477654
rect 589080 477334 589680 477418
rect 589080 477098 589262 477334
rect 589498 477098 589680 477334
rect 589080 441654 589680 477098
rect 589080 441418 589262 441654
rect 589498 441418 589680 441654
rect 589080 441334 589680 441418
rect 589080 441098 589262 441334
rect 589498 441098 589680 441334
rect 589080 405654 589680 441098
rect 589080 405418 589262 405654
rect 589498 405418 589680 405654
rect 589080 405334 589680 405418
rect 589080 405098 589262 405334
rect 589498 405098 589680 405334
rect 589080 369654 589680 405098
rect 589080 369418 589262 369654
rect 589498 369418 589680 369654
rect 589080 369334 589680 369418
rect 589080 369098 589262 369334
rect 589498 369098 589680 369334
rect 589080 333654 589680 369098
rect 589080 333418 589262 333654
rect 589498 333418 589680 333654
rect 589080 333334 589680 333418
rect 589080 333098 589262 333334
rect 589498 333098 589680 333334
rect 589080 297654 589680 333098
rect 589080 297418 589262 297654
rect 589498 297418 589680 297654
rect 589080 297334 589680 297418
rect 589080 297098 589262 297334
rect 589498 297098 589680 297334
rect 589080 261654 589680 297098
rect 589080 261418 589262 261654
rect 589498 261418 589680 261654
rect 589080 261334 589680 261418
rect 589080 261098 589262 261334
rect 589498 261098 589680 261334
rect 589080 225654 589680 261098
rect 589080 225418 589262 225654
rect 589498 225418 589680 225654
rect 589080 225334 589680 225418
rect 589080 225098 589262 225334
rect 589498 225098 589680 225334
rect 589080 189654 589680 225098
rect 589080 189418 589262 189654
rect 589498 189418 589680 189654
rect 589080 189334 589680 189418
rect 589080 189098 589262 189334
rect 589498 189098 589680 189334
rect 589080 153654 589680 189098
rect 589080 153418 589262 153654
rect 589498 153418 589680 153654
rect 589080 153334 589680 153418
rect 589080 153098 589262 153334
rect 589498 153098 589680 153334
rect 589080 117654 589680 153098
rect 589080 117418 589262 117654
rect 589498 117418 589680 117654
rect 589080 117334 589680 117418
rect 589080 117098 589262 117334
rect 589498 117098 589680 117334
rect 589080 81654 589680 117098
rect 589080 81418 589262 81654
rect 589498 81418 589680 81654
rect 589080 81334 589680 81418
rect 589080 81098 589262 81334
rect 589498 81098 589680 81334
rect 589080 45654 589680 81098
rect 589080 45418 589262 45654
rect 589498 45418 589680 45654
rect 589080 45334 589680 45418
rect 589080 45098 589262 45334
rect 589498 45098 589680 45334
rect 589080 9654 589680 45098
rect 589080 9418 589262 9654
rect 589498 9418 589680 9654
rect 589080 9334 589680 9418
rect 589080 9098 589262 9334
rect 589498 9098 589680 9334
rect 589080 -4106 589680 9098
rect 589080 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect 589080 -4426 589680 -4342
rect 589080 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect 589080 -4684 589680 -4662
rect 590020 675654 590620 708982
rect 590020 675418 590202 675654
rect 590438 675418 590620 675654
rect 590020 675334 590620 675418
rect 590020 675098 590202 675334
rect 590438 675098 590620 675334
rect 590020 639654 590620 675098
rect 590020 639418 590202 639654
rect 590438 639418 590620 639654
rect 590020 639334 590620 639418
rect 590020 639098 590202 639334
rect 590438 639098 590620 639334
rect 590020 603654 590620 639098
rect 590020 603418 590202 603654
rect 590438 603418 590620 603654
rect 590020 603334 590620 603418
rect 590020 603098 590202 603334
rect 590438 603098 590620 603334
rect 590020 567654 590620 603098
rect 590020 567418 590202 567654
rect 590438 567418 590620 567654
rect 590020 567334 590620 567418
rect 590020 567098 590202 567334
rect 590438 567098 590620 567334
rect 590020 531654 590620 567098
rect 590020 531418 590202 531654
rect 590438 531418 590620 531654
rect 590020 531334 590620 531418
rect 590020 531098 590202 531334
rect 590438 531098 590620 531334
rect 590020 495654 590620 531098
rect 590020 495418 590202 495654
rect 590438 495418 590620 495654
rect 590020 495334 590620 495418
rect 590020 495098 590202 495334
rect 590438 495098 590620 495334
rect 590020 459654 590620 495098
rect 590020 459418 590202 459654
rect 590438 459418 590620 459654
rect 590020 459334 590620 459418
rect 590020 459098 590202 459334
rect 590438 459098 590620 459334
rect 590020 423654 590620 459098
rect 590020 423418 590202 423654
rect 590438 423418 590620 423654
rect 590020 423334 590620 423418
rect 590020 423098 590202 423334
rect 590438 423098 590620 423334
rect 590020 387654 590620 423098
rect 590020 387418 590202 387654
rect 590438 387418 590620 387654
rect 590020 387334 590620 387418
rect 590020 387098 590202 387334
rect 590438 387098 590620 387334
rect 590020 351654 590620 387098
rect 590020 351418 590202 351654
rect 590438 351418 590620 351654
rect 590020 351334 590620 351418
rect 590020 351098 590202 351334
rect 590438 351098 590620 351334
rect 590020 315654 590620 351098
rect 590020 315418 590202 315654
rect 590438 315418 590620 315654
rect 590020 315334 590620 315418
rect 590020 315098 590202 315334
rect 590438 315098 590620 315334
rect 590020 279654 590620 315098
rect 590020 279418 590202 279654
rect 590438 279418 590620 279654
rect 590020 279334 590620 279418
rect 590020 279098 590202 279334
rect 590438 279098 590620 279334
rect 590020 243654 590620 279098
rect 590020 243418 590202 243654
rect 590438 243418 590620 243654
rect 590020 243334 590620 243418
rect 590020 243098 590202 243334
rect 590438 243098 590620 243334
rect 590020 207654 590620 243098
rect 590020 207418 590202 207654
rect 590438 207418 590620 207654
rect 590020 207334 590620 207418
rect 590020 207098 590202 207334
rect 590438 207098 590620 207334
rect 590020 171654 590620 207098
rect 590020 171418 590202 171654
rect 590438 171418 590620 171654
rect 590020 171334 590620 171418
rect 590020 171098 590202 171334
rect 590438 171098 590620 171334
rect 590020 135654 590620 171098
rect 590020 135418 590202 135654
rect 590438 135418 590620 135654
rect 590020 135334 590620 135418
rect 590020 135098 590202 135334
rect 590438 135098 590620 135334
rect 590020 99654 590620 135098
rect 590020 99418 590202 99654
rect 590438 99418 590620 99654
rect 590020 99334 590620 99418
rect 590020 99098 590202 99334
rect 590438 99098 590620 99334
rect 590020 63654 590620 99098
rect 590020 63418 590202 63654
rect 590438 63418 590620 63654
rect 590020 63334 590620 63418
rect 590020 63098 590202 63334
rect 590438 63098 590620 63334
rect 590020 27654 590620 63098
rect 590020 27418 590202 27654
rect 590438 27418 590620 27654
rect 590020 27334 590620 27418
rect 590020 27098 590202 27334
rect 590438 27098 590620 27334
rect 590020 -5046 590620 27098
rect 590020 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect 590020 -5366 590620 -5282
rect 590020 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect 590020 -5624 590620 -5602
rect 590960 697254 591560 709922
rect 590960 697018 591142 697254
rect 591378 697018 591560 697254
rect 590960 696934 591560 697018
rect 590960 696698 591142 696934
rect 591378 696698 591560 696934
rect 590960 661254 591560 696698
rect 590960 661018 591142 661254
rect 591378 661018 591560 661254
rect 590960 660934 591560 661018
rect 590960 660698 591142 660934
rect 591378 660698 591560 660934
rect 590960 625254 591560 660698
rect 590960 625018 591142 625254
rect 591378 625018 591560 625254
rect 590960 624934 591560 625018
rect 590960 624698 591142 624934
rect 591378 624698 591560 624934
rect 590960 589254 591560 624698
rect 590960 589018 591142 589254
rect 591378 589018 591560 589254
rect 590960 588934 591560 589018
rect 590960 588698 591142 588934
rect 591378 588698 591560 588934
rect 590960 553254 591560 588698
rect 590960 553018 591142 553254
rect 591378 553018 591560 553254
rect 590960 552934 591560 553018
rect 590960 552698 591142 552934
rect 591378 552698 591560 552934
rect 590960 517254 591560 552698
rect 590960 517018 591142 517254
rect 591378 517018 591560 517254
rect 590960 516934 591560 517018
rect 590960 516698 591142 516934
rect 591378 516698 591560 516934
rect 590960 481254 591560 516698
rect 590960 481018 591142 481254
rect 591378 481018 591560 481254
rect 590960 480934 591560 481018
rect 590960 480698 591142 480934
rect 591378 480698 591560 480934
rect 590960 445254 591560 480698
rect 590960 445018 591142 445254
rect 591378 445018 591560 445254
rect 590960 444934 591560 445018
rect 590960 444698 591142 444934
rect 591378 444698 591560 444934
rect 590960 409254 591560 444698
rect 590960 409018 591142 409254
rect 591378 409018 591560 409254
rect 590960 408934 591560 409018
rect 590960 408698 591142 408934
rect 591378 408698 591560 408934
rect 590960 373254 591560 408698
rect 590960 373018 591142 373254
rect 591378 373018 591560 373254
rect 590960 372934 591560 373018
rect 590960 372698 591142 372934
rect 591378 372698 591560 372934
rect 590960 337254 591560 372698
rect 590960 337018 591142 337254
rect 591378 337018 591560 337254
rect 590960 336934 591560 337018
rect 590960 336698 591142 336934
rect 591378 336698 591560 336934
rect 590960 301254 591560 336698
rect 590960 301018 591142 301254
rect 591378 301018 591560 301254
rect 590960 300934 591560 301018
rect 590960 300698 591142 300934
rect 591378 300698 591560 300934
rect 590960 265254 591560 300698
rect 590960 265018 591142 265254
rect 591378 265018 591560 265254
rect 590960 264934 591560 265018
rect 590960 264698 591142 264934
rect 591378 264698 591560 264934
rect 590960 229254 591560 264698
rect 590960 229018 591142 229254
rect 591378 229018 591560 229254
rect 590960 228934 591560 229018
rect 590960 228698 591142 228934
rect 591378 228698 591560 228934
rect 590960 193254 591560 228698
rect 590960 193018 591142 193254
rect 591378 193018 591560 193254
rect 590960 192934 591560 193018
rect 590960 192698 591142 192934
rect 591378 192698 591560 192934
rect 590960 157254 591560 192698
rect 590960 157018 591142 157254
rect 591378 157018 591560 157254
rect 590960 156934 591560 157018
rect 590960 156698 591142 156934
rect 591378 156698 591560 156934
rect 590960 121254 591560 156698
rect 590960 121018 591142 121254
rect 591378 121018 591560 121254
rect 590960 120934 591560 121018
rect 590960 120698 591142 120934
rect 591378 120698 591560 120934
rect 590960 85254 591560 120698
rect 590960 85018 591142 85254
rect 591378 85018 591560 85254
rect 590960 84934 591560 85018
rect 590960 84698 591142 84934
rect 591378 84698 591560 84934
rect 590960 49254 591560 84698
rect 590960 49018 591142 49254
rect 591378 49018 591560 49254
rect 590960 48934 591560 49018
rect 590960 48698 591142 48934
rect 591378 48698 591560 48934
rect 590960 13254 591560 48698
rect 590960 13018 591142 13254
rect 591378 13018 591560 13254
rect 590960 12934 591560 13018
rect 590960 12698 591142 12934
rect 591378 12698 591560 12934
rect 590960 -5986 591560 12698
rect 590960 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect 590960 -6306 591560 -6222
rect 590960 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect 590960 -6564 591560 -6542
rect 591900 679254 592500 710862
rect 591900 679018 592082 679254
rect 592318 679018 592500 679254
rect 591900 678934 592500 679018
rect 591900 678698 592082 678934
rect 592318 678698 592500 678934
rect 591900 643254 592500 678698
rect 591900 643018 592082 643254
rect 592318 643018 592500 643254
rect 591900 642934 592500 643018
rect 591900 642698 592082 642934
rect 592318 642698 592500 642934
rect 591900 607254 592500 642698
rect 591900 607018 592082 607254
rect 592318 607018 592500 607254
rect 591900 606934 592500 607018
rect 591900 606698 592082 606934
rect 592318 606698 592500 606934
rect 591900 571254 592500 606698
rect 591900 571018 592082 571254
rect 592318 571018 592500 571254
rect 591900 570934 592500 571018
rect 591900 570698 592082 570934
rect 592318 570698 592500 570934
rect 591900 535254 592500 570698
rect 591900 535018 592082 535254
rect 592318 535018 592500 535254
rect 591900 534934 592500 535018
rect 591900 534698 592082 534934
rect 592318 534698 592500 534934
rect 591900 499254 592500 534698
rect 591900 499018 592082 499254
rect 592318 499018 592500 499254
rect 591900 498934 592500 499018
rect 591900 498698 592082 498934
rect 592318 498698 592500 498934
rect 591900 463254 592500 498698
rect 591900 463018 592082 463254
rect 592318 463018 592500 463254
rect 591900 462934 592500 463018
rect 591900 462698 592082 462934
rect 592318 462698 592500 462934
rect 591900 427254 592500 462698
rect 591900 427018 592082 427254
rect 592318 427018 592500 427254
rect 591900 426934 592500 427018
rect 591900 426698 592082 426934
rect 592318 426698 592500 426934
rect 591900 391254 592500 426698
rect 591900 391018 592082 391254
rect 592318 391018 592500 391254
rect 591900 390934 592500 391018
rect 591900 390698 592082 390934
rect 592318 390698 592500 390934
rect 591900 355254 592500 390698
rect 591900 355018 592082 355254
rect 592318 355018 592500 355254
rect 591900 354934 592500 355018
rect 591900 354698 592082 354934
rect 592318 354698 592500 354934
rect 591900 319254 592500 354698
rect 591900 319018 592082 319254
rect 592318 319018 592500 319254
rect 591900 318934 592500 319018
rect 591900 318698 592082 318934
rect 592318 318698 592500 318934
rect 591900 283254 592500 318698
rect 591900 283018 592082 283254
rect 592318 283018 592500 283254
rect 591900 282934 592500 283018
rect 591900 282698 592082 282934
rect 592318 282698 592500 282934
rect 591900 247254 592500 282698
rect 591900 247018 592082 247254
rect 592318 247018 592500 247254
rect 591900 246934 592500 247018
rect 591900 246698 592082 246934
rect 592318 246698 592500 246934
rect 591900 211254 592500 246698
rect 591900 211018 592082 211254
rect 592318 211018 592500 211254
rect 591900 210934 592500 211018
rect 591900 210698 592082 210934
rect 592318 210698 592500 210934
rect 591900 175254 592500 210698
rect 591900 175018 592082 175254
rect 592318 175018 592500 175254
rect 591900 174934 592500 175018
rect 591900 174698 592082 174934
rect 592318 174698 592500 174934
rect 591900 139254 592500 174698
rect 591900 139018 592082 139254
rect 592318 139018 592500 139254
rect 591900 138934 592500 139018
rect 591900 138698 592082 138934
rect 592318 138698 592500 138934
rect 591900 103254 592500 138698
rect 591900 103018 592082 103254
rect 592318 103018 592500 103254
rect 591900 102934 592500 103018
rect 591900 102698 592082 102934
rect 592318 102698 592500 102934
rect 591900 67254 592500 102698
rect 591900 67018 592082 67254
rect 592318 67018 592500 67254
rect 591900 66934 592500 67018
rect 591900 66698 592082 66934
rect 592318 66698 592500 66934
rect 591900 31254 592500 66698
rect 591900 31018 592082 31254
rect 592318 31018 592500 31254
rect 591900 30934 592500 31018
rect 591900 30698 592082 30934
rect 592318 30698 592500 30934
rect 569604 -7162 569786 -6926
rect 570022 -7162 570204 -6926
rect 569604 -7246 570204 -7162
rect 569604 -7482 569786 -7246
rect 570022 -7482 570204 -7246
rect 569604 -7504 570204 -7482
rect 591900 -6926 592500 30698
rect 591900 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect 591900 -7246 592500 -7162
rect 591900 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect 591900 -7504 592500 -7482
<< via4 >>
rect -8394 711182 -8158 711418
rect -8394 710862 -8158 711098
rect -8394 679018 -8158 679254
rect -8394 678698 -8158 678934
rect -8394 643018 -8158 643254
rect -8394 642698 -8158 642934
rect -8394 607018 -8158 607254
rect -8394 606698 -8158 606934
rect -8394 571018 -8158 571254
rect -8394 570698 -8158 570934
rect -8394 535018 -8158 535254
rect -8394 534698 -8158 534934
rect -8394 499018 -8158 499254
rect -8394 498698 -8158 498934
rect -8394 463018 -8158 463254
rect -8394 462698 -8158 462934
rect -8394 427018 -8158 427254
rect -8394 426698 -8158 426934
rect -8394 391018 -8158 391254
rect -8394 390698 -8158 390934
rect -8394 355018 -8158 355254
rect -8394 354698 -8158 354934
rect -8394 319018 -8158 319254
rect -8394 318698 -8158 318934
rect -8394 283018 -8158 283254
rect -8394 282698 -8158 282934
rect -8394 247018 -8158 247254
rect -8394 246698 -8158 246934
rect -8394 211018 -8158 211254
rect -8394 210698 -8158 210934
rect -8394 175018 -8158 175254
rect -8394 174698 -8158 174934
rect -8394 139018 -8158 139254
rect -8394 138698 -8158 138934
rect -8394 103018 -8158 103254
rect -8394 102698 -8158 102934
rect -8394 67018 -8158 67254
rect -8394 66698 -8158 66934
rect -8394 31018 -8158 31254
rect -8394 30698 -8158 30934
rect -7454 710242 -7218 710478
rect -7454 709922 -7218 710158
rect 11786 710242 12022 710478
rect 11786 709922 12022 710158
rect -7454 697018 -7218 697254
rect -7454 696698 -7218 696934
rect -7454 661018 -7218 661254
rect -7454 660698 -7218 660934
rect -7454 625018 -7218 625254
rect -7454 624698 -7218 624934
rect -7454 589018 -7218 589254
rect -7454 588698 -7218 588934
rect -7454 553018 -7218 553254
rect -7454 552698 -7218 552934
rect -7454 517018 -7218 517254
rect -7454 516698 -7218 516934
rect -7454 481018 -7218 481254
rect -7454 480698 -7218 480934
rect -7454 445018 -7218 445254
rect -7454 444698 -7218 444934
rect -7454 409018 -7218 409254
rect -7454 408698 -7218 408934
rect -7454 373018 -7218 373254
rect -7454 372698 -7218 372934
rect -7454 337018 -7218 337254
rect -7454 336698 -7218 336934
rect -7454 301018 -7218 301254
rect -7454 300698 -7218 300934
rect -7454 265018 -7218 265254
rect -7454 264698 -7218 264934
rect -7454 229018 -7218 229254
rect -7454 228698 -7218 228934
rect -7454 193018 -7218 193254
rect -7454 192698 -7218 192934
rect -7454 157018 -7218 157254
rect -7454 156698 -7218 156934
rect -7454 121018 -7218 121254
rect -7454 120698 -7218 120934
rect -7454 85018 -7218 85254
rect -7454 84698 -7218 84934
rect -7454 49018 -7218 49254
rect -7454 48698 -7218 48934
rect -7454 13018 -7218 13254
rect -7454 12698 -7218 12934
rect -6514 709302 -6278 709538
rect -6514 708982 -6278 709218
rect -6514 675418 -6278 675654
rect -6514 675098 -6278 675334
rect -6514 639418 -6278 639654
rect -6514 639098 -6278 639334
rect -6514 603418 -6278 603654
rect -6514 603098 -6278 603334
rect -6514 567418 -6278 567654
rect -6514 567098 -6278 567334
rect -6514 531418 -6278 531654
rect -6514 531098 -6278 531334
rect -6514 495418 -6278 495654
rect -6514 495098 -6278 495334
rect -6514 459418 -6278 459654
rect -6514 459098 -6278 459334
rect -6514 423418 -6278 423654
rect -6514 423098 -6278 423334
rect -6514 387418 -6278 387654
rect -6514 387098 -6278 387334
rect -6514 351418 -6278 351654
rect -6514 351098 -6278 351334
rect -6514 315418 -6278 315654
rect -6514 315098 -6278 315334
rect -6514 279418 -6278 279654
rect -6514 279098 -6278 279334
rect -6514 243418 -6278 243654
rect -6514 243098 -6278 243334
rect -6514 207418 -6278 207654
rect -6514 207098 -6278 207334
rect -6514 171418 -6278 171654
rect -6514 171098 -6278 171334
rect -6514 135418 -6278 135654
rect -6514 135098 -6278 135334
rect -6514 99418 -6278 99654
rect -6514 99098 -6278 99334
rect -6514 63418 -6278 63654
rect -6514 63098 -6278 63334
rect -6514 27418 -6278 27654
rect -6514 27098 -6278 27334
rect -5574 708362 -5338 708598
rect -5574 708042 -5338 708278
rect 8186 708362 8422 708598
rect 8186 708042 8422 708278
rect -5574 693418 -5338 693654
rect -5574 693098 -5338 693334
rect -5574 657418 -5338 657654
rect -5574 657098 -5338 657334
rect -5574 621418 -5338 621654
rect -5574 621098 -5338 621334
rect -5574 585418 -5338 585654
rect -5574 585098 -5338 585334
rect -5574 549418 -5338 549654
rect -5574 549098 -5338 549334
rect -5574 513418 -5338 513654
rect -5574 513098 -5338 513334
rect -5574 477418 -5338 477654
rect -5574 477098 -5338 477334
rect -5574 441418 -5338 441654
rect -5574 441098 -5338 441334
rect -5574 405418 -5338 405654
rect -5574 405098 -5338 405334
rect -5574 369418 -5338 369654
rect -5574 369098 -5338 369334
rect -5574 333418 -5338 333654
rect -5574 333098 -5338 333334
rect -5574 297418 -5338 297654
rect -5574 297098 -5338 297334
rect -5574 261418 -5338 261654
rect -5574 261098 -5338 261334
rect -5574 225418 -5338 225654
rect -5574 225098 -5338 225334
rect -5574 189418 -5338 189654
rect -5574 189098 -5338 189334
rect -5574 153418 -5338 153654
rect -5574 153098 -5338 153334
rect -5574 117418 -5338 117654
rect -5574 117098 -5338 117334
rect -5574 81418 -5338 81654
rect -5574 81098 -5338 81334
rect -5574 45418 -5338 45654
rect -5574 45098 -5338 45334
rect -5574 9418 -5338 9654
rect -5574 9098 -5338 9334
rect -4634 707422 -4398 707658
rect -4634 707102 -4398 707338
rect -4634 671818 -4398 672054
rect -4634 671498 -4398 671734
rect -4634 635818 -4398 636054
rect -4634 635498 -4398 635734
rect -4634 599818 -4398 600054
rect -4634 599498 -4398 599734
rect -4634 563818 -4398 564054
rect -4634 563498 -4398 563734
rect -4634 527818 -4398 528054
rect -4634 527498 -4398 527734
rect -4634 491818 -4398 492054
rect -4634 491498 -4398 491734
rect -4634 455818 -4398 456054
rect -4634 455498 -4398 455734
rect -4634 419818 -4398 420054
rect -4634 419498 -4398 419734
rect -4634 383818 -4398 384054
rect -4634 383498 -4398 383734
rect -4634 347818 -4398 348054
rect -4634 347498 -4398 347734
rect -4634 311818 -4398 312054
rect -4634 311498 -4398 311734
rect -4634 275818 -4398 276054
rect -4634 275498 -4398 275734
rect -4634 239818 -4398 240054
rect -4634 239498 -4398 239734
rect -4634 203818 -4398 204054
rect -4634 203498 -4398 203734
rect -4634 167818 -4398 168054
rect -4634 167498 -4398 167734
rect -4634 131818 -4398 132054
rect -4634 131498 -4398 131734
rect -4634 95818 -4398 96054
rect -4634 95498 -4398 95734
rect -4634 59818 -4398 60054
rect -4634 59498 -4398 59734
rect -4634 23818 -4398 24054
rect -4634 23498 -4398 23734
rect -3694 706482 -3458 706718
rect -3694 706162 -3458 706398
rect 4586 706482 4822 706718
rect 4586 706162 4822 706398
rect -3694 689818 -3458 690054
rect -3694 689498 -3458 689734
rect -3694 653818 -3458 654054
rect -3694 653498 -3458 653734
rect -3694 617818 -3458 618054
rect -3694 617498 -3458 617734
rect -3694 581818 -3458 582054
rect -3694 581498 -3458 581734
rect -3694 545818 -3458 546054
rect -3694 545498 -3458 545734
rect -3694 509818 -3458 510054
rect -3694 509498 -3458 509734
rect -3694 473818 -3458 474054
rect -3694 473498 -3458 473734
rect -3694 437818 -3458 438054
rect -3694 437498 -3458 437734
rect -3694 401818 -3458 402054
rect -3694 401498 -3458 401734
rect -3694 365818 -3458 366054
rect -3694 365498 -3458 365734
rect -3694 329818 -3458 330054
rect -3694 329498 -3458 329734
rect -3694 293818 -3458 294054
rect -3694 293498 -3458 293734
rect -3694 257818 -3458 258054
rect -3694 257498 -3458 257734
rect -3694 221818 -3458 222054
rect -3694 221498 -3458 221734
rect -3694 185818 -3458 186054
rect -3694 185498 -3458 185734
rect -3694 149818 -3458 150054
rect -3694 149498 -3458 149734
rect -3694 113818 -3458 114054
rect -3694 113498 -3458 113734
rect -3694 77818 -3458 78054
rect -3694 77498 -3458 77734
rect -3694 41818 -3458 42054
rect -3694 41498 -3458 41734
rect -3694 5818 -3458 6054
rect -3694 5498 -3458 5734
rect -2754 705542 -2518 705778
rect -2754 705222 -2518 705458
rect -2754 668218 -2518 668454
rect -2754 667898 -2518 668134
rect -2754 632218 -2518 632454
rect -2754 631898 -2518 632134
rect -2754 596218 -2518 596454
rect -2754 595898 -2518 596134
rect -2754 560218 -2518 560454
rect -2754 559898 -2518 560134
rect -2754 524218 -2518 524454
rect -2754 523898 -2518 524134
rect -2754 488218 -2518 488454
rect -2754 487898 -2518 488134
rect -2754 452218 -2518 452454
rect -2754 451898 -2518 452134
rect -2754 416218 -2518 416454
rect -2754 415898 -2518 416134
rect -2754 380218 -2518 380454
rect -2754 379898 -2518 380134
rect -2754 344218 -2518 344454
rect -2754 343898 -2518 344134
rect -2754 308218 -2518 308454
rect -2754 307898 -2518 308134
rect -2754 272218 -2518 272454
rect -2754 271898 -2518 272134
rect -2754 236218 -2518 236454
rect -2754 235898 -2518 236134
rect -2754 200218 -2518 200454
rect -2754 199898 -2518 200134
rect -2754 164218 -2518 164454
rect -2754 163898 -2518 164134
rect -2754 128218 -2518 128454
rect -2754 127898 -2518 128134
rect -2754 92218 -2518 92454
rect -2754 91898 -2518 92134
rect -2754 56218 -2518 56454
rect -2754 55898 -2518 56134
rect -2754 20218 -2518 20454
rect -2754 19898 -2518 20134
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect -1814 686218 -1578 686454
rect -1814 685898 -1578 686134
rect -1814 650218 -1578 650454
rect -1814 649898 -1578 650134
rect -1814 614218 -1578 614454
rect -1814 613898 -1578 614134
rect -1814 578218 -1578 578454
rect -1814 577898 -1578 578134
rect -1814 542218 -1578 542454
rect -1814 541898 -1578 542134
rect -1814 506218 -1578 506454
rect -1814 505898 -1578 506134
rect -1814 470218 -1578 470454
rect -1814 469898 -1578 470134
rect -1814 434218 -1578 434454
rect -1814 433898 -1578 434134
rect -1814 398218 -1578 398454
rect -1814 397898 -1578 398134
rect -1814 362218 -1578 362454
rect -1814 361898 -1578 362134
rect -1814 326218 -1578 326454
rect -1814 325898 -1578 326134
rect -1814 290218 -1578 290454
rect -1814 289898 -1578 290134
rect -1814 254218 -1578 254454
rect -1814 253898 -1578 254134
rect -1814 218218 -1578 218454
rect -1814 217898 -1578 218134
rect -1814 182218 -1578 182454
rect -1814 181898 -1578 182134
rect -1814 146218 -1578 146454
rect -1814 145898 -1578 146134
rect -1814 110218 -1578 110454
rect -1814 109898 -1578 110134
rect -1814 74218 -1578 74454
rect -1814 73898 -1578 74134
rect -1814 38218 -1578 38454
rect -1814 37898 -1578 38134
rect -1814 2218 -1578 2454
rect -1814 1898 -1578 2134
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 986 704602 1222 704838
rect 986 704282 1222 704518
rect 986 686218 1222 686454
rect 986 685898 1222 686134
rect 986 650218 1222 650454
rect 986 649898 1222 650134
rect 986 614218 1222 614454
rect 986 613898 1222 614134
rect 986 578218 1222 578454
rect 986 577898 1222 578134
rect 986 542218 1222 542454
rect 986 541898 1222 542134
rect 986 506218 1222 506454
rect 986 505898 1222 506134
rect 986 470218 1222 470454
rect 986 469898 1222 470134
rect 986 434218 1222 434454
rect 986 433898 1222 434134
rect 986 398218 1222 398454
rect 986 397898 1222 398134
rect 986 362218 1222 362454
rect 986 361898 1222 362134
rect 986 326218 1222 326454
rect 986 325898 1222 326134
rect 986 290218 1222 290454
rect 986 289898 1222 290134
rect 986 254218 1222 254454
rect 986 253898 1222 254134
rect 986 218218 1222 218454
rect 986 217898 1222 218134
rect 986 182218 1222 182454
rect 986 181898 1222 182134
rect 986 146218 1222 146454
rect 986 145898 1222 146134
rect 986 110218 1222 110454
rect 986 109898 1222 110134
rect 986 74218 1222 74454
rect 986 73898 1222 74134
rect 986 38218 1222 38454
rect 986 37898 1222 38134
rect 986 2218 1222 2454
rect 986 1898 1222 2134
rect 986 -582 1222 -346
rect 986 -902 1222 -666
rect -2754 -1522 -2518 -1286
rect -2754 -1842 -2518 -1606
rect 4586 689818 4822 690054
rect 4586 689498 4822 689734
rect 4586 653818 4822 654054
rect 4586 653498 4822 653734
rect 4586 617818 4822 618054
rect 4586 617498 4822 617734
rect 4586 581818 4822 582054
rect 4586 581498 4822 581734
rect 4586 545818 4822 546054
rect 4586 545498 4822 545734
rect 4586 509818 4822 510054
rect 4586 509498 4822 509734
rect 4586 473818 4822 474054
rect 4586 473498 4822 473734
rect 4586 437818 4822 438054
rect 4586 437498 4822 437734
rect 4586 401818 4822 402054
rect 4586 401498 4822 401734
rect 4586 365818 4822 366054
rect 4586 365498 4822 365734
rect 4586 329818 4822 330054
rect 4586 329498 4822 329734
rect 4586 293818 4822 294054
rect 4586 293498 4822 293734
rect 4586 257818 4822 258054
rect 4586 257498 4822 257734
rect 4586 221818 4822 222054
rect 4586 221498 4822 221734
rect 4586 185818 4822 186054
rect 4586 185498 4822 185734
rect 4586 149818 4822 150054
rect 4586 149498 4822 149734
rect 4586 113818 4822 114054
rect 4586 113498 4822 113734
rect 4586 77818 4822 78054
rect 4586 77498 4822 77734
rect 4586 41818 4822 42054
rect 4586 41498 4822 41734
rect 4586 5818 4822 6054
rect 4586 5498 4822 5734
rect -3694 -2462 -3458 -2226
rect -3694 -2782 -3458 -2546
rect 4586 -2462 4822 -2226
rect 4586 -2782 4822 -2546
rect -4634 -3402 -4398 -3166
rect -4634 -3722 -4398 -3486
rect 8186 693418 8422 693654
rect 8186 693098 8422 693334
rect 8186 657418 8422 657654
rect 8186 657098 8422 657334
rect 8186 621418 8422 621654
rect 8186 621098 8422 621334
rect 8186 585418 8422 585654
rect 8186 585098 8422 585334
rect 8186 549418 8422 549654
rect 8186 549098 8422 549334
rect 8186 513418 8422 513654
rect 8186 513098 8422 513334
rect 8186 477418 8422 477654
rect 8186 477098 8422 477334
rect 8186 441418 8422 441654
rect 8186 441098 8422 441334
rect 8186 405418 8422 405654
rect 8186 405098 8422 405334
rect 8186 369418 8422 369654
rect 8186 369098 8422 369334
rect 8186 333418 8422 333654
rect 8186 333098 8422 333334
rect 8186 297418 8422 297654
rect 8186 297098 8422 297334
rect 8186 261418 8422 261654
rect 8186 261098 8422 261334
rect 8186 225418 8422 225654
rect 8186 225098 8422 225334
rect 8186 189418 8422 189654
rect 8186 189098 8422 189334
rect 8186 153418 8422 153654
rect 8186 153098 8422 153334
rect 8186 117418 8422 117654
rect 8186 117098 8422 117334
rect 8186 81418 8422 81654
rect 8186 81098 8422 81334
rect 8186 45418 8422 45654
rect 8186 45098 8422 45334
rect 8186 9418 8422 9654
rect 8186 9098 8422 9334
rect -5574 -4342 -5338 -4106
rect -5574 -4662 -5338 -4426
rect 8186 -4342 8422 -4106
rect 8186 -4662 8422 -4426
rect -6514 -5282 -6278 -5046
rect -6514 -5602 -6278 -5366
rect 29786 711182 30022 711418
rect 29786 710862 30022 711098
rect 26186 709302 26422 709538
rect 26186 708982 26422 709218
rect 22586 707422 22822 707658
rect 22586 707102 22822 707338
rect 11786 697018 12022 697254
rect 11786 696698 12022 696934
rect 11786 661018 12022 661254
rect 11786 660698 12022 660934
rect 11786 625018 12022 625254
rect 11786 624698 12022 624934
rect 11786 589018 12022 589254
rect 11786 588698 12022 588934
rect 11786 553018 12022 553254
rect 11786 552698 12022 552934
rect 11786 517018 12022 517254
rect 11786 516698 12022 516934
rect 11786 481018 12022 481254
rect 11786 480698 12022 480934
rect 11786 445018 12022 445254
rect 11786 444698 12022 444934
rect 11786 409018 12022 409254
rect 11786 408698 12022 408934
rect 11786 373018 12022 373254
rect 11786 372698 12022 372934
rect 11786 337018 12022 337254
rect 11786 336698 12022 336934
rect 11786 301018 12022 301254
rect 11786 300698 12022 300934
rect 11786 265018 12022 265254
rect 11786 264698 12022 264934
rect 11786 229018 12022 229254
rect 11786 228698 12022 228934
rect 11786 193018 12022 193254
rect 11786 192698 12022 192934
rect 11786 157018 12022 157254
rect 11786 156698 12022 156934
rect 11786 121018 12022 121254
rect 11786 120698 12022 120934
rect 11786 85018 12022 85254
rect 11786 84698 12022 84934
rect 11786 49018 12022 49254
rect 11786 48698 12022 48934
rect 11786 13018 12022 13254
rect 11786 12698 12022 12934
rect -7454 -6222 -7218 -5986
rect -7454 -6542 -7218 -6306
rect 18986 705542 19222 705778
rect 18986 705222 19222 705458
rect 18986 668218 19222 668454
rect 18986 667898 19222 668134
rect 18986 632218 19222 632454
rect 18986 631898 19222 632134
rect 18986 596218 19222 596454
rect 18986 595898 19222 596134
rect 18986 560218 19222 560454
rect 18986 559898 19222 560134
rect 18986 524218 19222 524454
rect 18986 523898 19222 524134
rect 18986 488218 19222 488454
rect 18986 487898 19222 488134
rect 18986 452218 19222 452454
rect 18986 451898 19222 452134
rect 18986 416218 19222 416454
rect 18986 415898 19222 416134
rect 18986 380218 19222 380454
rect 18986 379898 19222 380134
rect 18986 344218 19222 344454
rect 18986 343898 19222 344134
rect 18986 308218 19222 308454
rect 18986 307898 19222 308134
rect 18986 272218 19222 272454
rect 18986 271898 19222 272134
rect 18986 236218 19222 236454
rect 18986 235898 19222 236134
rect 18986 200218 19222 200454
rect 18986 199898 19222 200134
rect 18986 164218 19222 164454
rect 18986 163898 19222 164134
rect 18986 128218 19222 128454
rect 18986 127898 19222 128134
rect 18986 92218 19222 92454
rect 18986 91898 19222 92134
rect 18986 56218 19222 56454
rect 18986 55898 19222 56134
rect 18986 20218 19222 20454
rect 18986 19898 19222 20134
rect 18986 -1522 19222 -1286
rect 18986 -1842 19222 -1606
rect 22586 671818 22822 672054
rect 22586 671498 22822 671734
rect 22586 635818 22822 636054
rect 22586 635498 22822 635734
rect 22586 599818 22822 600054
rect 22586 599498 22822 599734
rect 22586 563818 22822 564054
rect 22586 563498 22822 563734
rect 22586 527818 22822 528054
rect 22586 527498 22822 527734
rect 22586 491818 22822 492054
rect 22586 491498 22822 491734
rect 22586 455818 22822 456054
rect 22586 455498 22822 455734
rect 22586 419818 22822 420054
rect 22586 419498 22822 419734
rect 22586 383818 22822 384054
rect 22586 383498 22822 383734
rect 22586 347818 22822 348054
rect 22586 347498 22822 347734
rect 22586 311818 22822 312054
rect 22586 311498 22822 311734
rect 22586 275818 22822 276054
rect 22586 275498 22822 275734
rect 22586 239818 22822 240054
rect 22586 239498 22822 239734
rect 22586 203818 22822 204054
rect 22586 203498 22822 203734
rect 22586 167818 22822 168054
rect 22586 167498 22822 167734
rect 22586 131818 22822 132054
rect 22586 131498 22822 131734
rect 22586 95818 22822 96054
rect 22586 95498 22822 95734
rect 22586 59818 22822 60054
rect 22586 59498 22822 59734
rect 22586 23818 22822 24054
rect 22586 23498 22822 23734
rect 22586 -3402 22822 -3166
rect 22586 -3722 22822 -3486
rect 26186 675418 26422 675654
rect 26186 675098 26422 675334
rect 26186 639418 26422 639654
rect 26186 639098 26422 639334
rect 26186 603418 26422 603654
rect 26186 603098 26422 603334
rect 26186 567418 26422 567654
rect 26186 567098 26422 567334
rect 26186 531418 26422 531654
rect 26186 531098 26422 531334
rect 26186 495418 26422 495654
rect 26186 495098 26422 495334
rect 26186 459418 26422 459654
rect 26186 459098 26422 459334
rect 26186 423418 26422 423654
rect 26186 423098 26422 423334
rect 26186 387418 26422 387654
rect 26186 387098 26422 387334
rect 26186 351418 26422 351654
rect 26186 351098 26422 351334
rect 26186 315418 26422 315654
rect 26186 315098 26422 315334
rect 26186 279418 26422 279654
rect 26186 279098 26422 279334
rect 26186 243418 26422 243654
rect 26186 243098 26422 243334
rect 26186 207418 26422 207654
rect 26186 207098 26422 207334
rect 26186 171418 26422 171654
rect 26186 171098 26422 171334
rect 26186 135418 26422 135654
rect 26186 135098 26422 135334
rect 26186 99418 26422 99654
rect 26186 99098 26422 99334
rect 26186 63418 26422 63654
rect 26186 63098 26422 63334
rect 26186 27418 26422 27654
rect 26186 27098 26422 27334
rect 26186 -5282 26422 -5046
rect 26186 -5602 26422 -5366
rect 47786 710242 48022 710478
rect 47786 709922 48022 710158
rect 44186 708362 44422 708598
rect 44186 708042 44422 708278
rect 40586 706482 40822 706718
rect 40586 706162 40822 706398
rect 29786 679018 30022 679254
rect 29786 678698 30022 678934
rect 29786 643018 30022 643254
rect 29786 642698 30022 642934
rect 29786 607018 30022 607254
rect 29786 606698 30022 606934
rect 29786 571018 30022 571254
rect 29786 570698 30022 570934
rect 29786 535018 30022 535254
rect 29786 534698 30022 534934
rect 29786 499018 30022 499254
rect 29786 498698 30022 498934
rect 29786 463018 30022 463254
rect 29786 462698 30022 462934
rect 29786 427018 30022 427254
rect 29786 426698 30022 426934
rect 29786 391018 30022 391254
rect 29786 390698 30022 390934
rect 29786 355018 30022 355254
rect 29786 354698 30022 354934
rect 29786 319018 30022 319254
rect 29786 318698 30022 318934
rect 29786 283018 30022 283254
rect 29786 282698 30022 282934
rect 29786 247018 30022 247254
rect 29786 246698 30022 246934
rect 29786 211018 30022 211254
rect 29786 210698 30022 210934
rect 29786 175018 30022 175254
rect 29786 174698 30022 174934
rect 29786 139018 30022 139254
rect 29786 138698 30022 138934
rect 29786 103018 30022 103254
rect 29786 102698 30022 102934
rect 29786 67018 30022 67254
rect 29786 66698 30022 66934
rect 29786 31018 30022 31254
rect 29786 30698 30022 30934
rect 11786 -6222 12022 -5986
rect 11786 -6542 12022 -6306
rect -8394 -7162 -8158 -6926
rect -8394 -7482 -8158 -7246
rect 36986 704602 37222 704838
rect 36986 704282 37222 704518
rect 36986 686218 37222 686454
rect 36986 685898 37222 686134
rect 36986 650218 37222 650454
rect 36986 649898 37222 650134
rect 36986 614218 37222 614454
rect 36986 613898 37222 614134
rect 36986 578218 37222 578454
rect 36986 577898 37222 578134
rect 36986 542218 37222 542454
rect 36986 541898 37222 542134
rect 36986 506218 37222 506454
rect 36986 505898 37222 506134
rect 36986 470218 37222 470454
rect 36986 469898 37222 470134
rect 36986 434218 37222 434454
rect 36986 433898 37222 434134
rect 36986 398218 37222 398454
rect 36986 397898 37222 398134
rect 36986 362218 37222 362454
rect 36986 361898 37222 362134
rect 36986 326218 37222 326454
rect 36986 325898 37222 326134
rect 36986 290218 37222 290454
rect 36986 289898 37222 290134
rect 36986 254218 37222 254454
rect 36986 253898 37222 254134
rect 36986 218218 37222 218454
rect 36986 217898 37222 218134
rect 36986 182218 37222 182454
rect 36986 181898 37222 182134
rect 36986 146218 37222 146454
rect 36986 145898 37222 146134
rect 36986 110218 37222 110454
rect 36986 109898 37222 110134
rect 36986 74218 37222 74454
rect 36986 73898 37222 74134
rect 36986 38218 37222 38454
rect 36986 37898 37222 38134
rect 36986 2218 37222 2454
rect 36986 1898 37222 2134
rect 36986 -582 37222 -346
rect 36986 -902 37222 -666
rect 40586 689818 40822 690054
rect 40586 689498 40822 689734
rect 40586 653818 40822 654054
rect 40586 653498 40822 653734
rect 40586 617818 40822 618054
rect 40586 617498 40822 617734
rect 40586 581818 40822 582054
rect 40586 581498 40822 581734
rect 40586 545818 40822 546054
rect 40586 545498 40822 545734
rect 40586 509818 40822 510054
rect 40586 509498 40822 509734
rect 40586 473818 40822 474054
rect 40586 473498 40822 473734
rect 40586 437818 40822 438054
rect 40586 437498 40822 437734
rect 40586 401818 40822 402054
rect 40586 401498 40822 401734
rect 40586 365818 40822 366054
rect 40586 365498 40822 365734
rect 40586 329818 40822 330054
rect 40586 329498 40822 329734
rect 40586 293818 40822 294054
rect 40586 293498 40822 293734
rect 40586 257818 40822 258054
rect 40586 257498 40822 257734
rect 40586 221818 40822 222054
rect 40586 221498 40822 221734
rect 40586 185818 40822 186054
rect 40586 185498 40822 185734
rect 40586 149818 40822 150054
rect 40586 149498 40822 149734
rect 40586 113818 40822 114054
rect 40586 113498 40822 113734
rect 40586 77818 40822 78054
rect 40586 77498 40822 77734
rect 40586 41818 40822 42054
rect 40586 41498 40822 41734
rect 40586 5818 40822 6054
rect 40586 5498 40822 5734
rect 40586 -2462 40822 -2226
rect 40586 -2782 40822 -2546
rect 44186 693418 44422 693654
rect 44186 693098 44422 693334
rect 44186 657418 44422 657654
rect 44186 657098 44422 657334
rect 44186 621418 44422 621654
rect 44186 621098 44422 621334
rect 44186 585418 44422 585654
rect 44186 585098 44422 585334
rect 44186 549418 44422 549654
rect 44186 549098 44422 549334
rect 44186 513418 44422 513654
rect 44186 513098 44422 513334
rect 44186 477418 44422 477654
rect 44186 477098 44422 477334
rect 44186 441418 44422 441654
rect 44186 441098 44422 441334
rect 44186 405418 44422 405654
rect 44186 405098 44422 405334
rect 44186 369418 44422 369654
rect 44186 369098 44422 369334
rect 44186 333418 44422 333654
rect 44186 333098 44422 333334
rect 44186 297418 44422 297654
rect 44186 297098 44422 297334
rect 44186 261418 44422 261654
rect 44186 261098 44422 261334
rect 44186 225418 44422 225654
rect 44186 225098 44422 225334
rect 44186 189418 44422 189654
rect 44186 189098 44422 189334
rect 44186 153418 44422 153654
rect 44186 153098 44422 153334
rect 44186 117418 44422 117654
rect 44186 117098 44422 117334
rect 44186 81418 44422 81654
rect 44186 81098 44422 81334
rect 44186 45418 44422 45654
rect 44186 45098 44422 45334
rect 44186 9418 44422 9654
rect 44186 9098 44422 9334
rect 44186 -4342 44422 -4106
rect 44186 -4662 44422 -4426
rect 65786 711182 66022 711418
rect 65786 710862 66022 711098
rect 62186 709302 62422 709538
rect 62186 708982 62422 709218
rect 58586 707422 58822 707658
rect 58586 707102 58822 707338
rect 47786 697018 48022 697254
rect 47786 696698 48022 696934
rect 47786 661018 48022 661254
rect 47786 660698 48022 660934
rect 47786 625018 48022 625254
rect 47786 624698 48022 624934
rect 47786 589018 48022 589254
rect 47786 588698 48022 588934
rect 47786 553018 48022 553254
rect 47786 552698 48022 552934
rect 47786 517018 48022 517254
rect 47786 516698 48022 516934
rect 47786 481018 48022 481254
rect 47786 480698 48022 480934
rect 47786 445018 48022 445254
rect 47786 444698 48022 444934
rect 47786 409018 48022 409254
rect 47786 408698 48022 408934
rect 47786 373018 48022 373254
rect 47786 372698 48022 372934
rect 47786 337018 48022 337254
rect 47786 336698 48022 336934
rect 47786 301018 48022 301254
rect 47786 300698 48022 300934
rect 47786 265018 48022 265254
rect 47786 264698 48022 264934
rect 47786 229018 48022 229254
rect 47786 228698 48022 228934
rect 47786 193018 48022 193254
rect 47786 192698 48022 192934
rect 47786 157018 48022 157254
rect 47786 156698 48022 156934
rect 47786 121018 48022 121254
rect 47786 120698 48022 120934
rect 47786 85018 48022 85254
rect 47786 84698 48022 84934
rect 47786 49018 48022 49254
rect 47786 48698 48022 48934
rect 47786 13018 48022 13254
rect 47786 12698 48022 12934
rect 29786 -7162 30022 -6926
rect 29786 -7482 30022 -7246
rect 54986 705542 55222 705778
rect 54986 705222 55222 705458
rect 54986 668218 55222 668454
rect 54986 667898 55222 668134
rect 58586 671818 58822 672054
rect 58586 671498 58822 671734
rect 62186 675418 62422 675654
rect 62186 675098 62422 675334
rect 83786 710242 84022 710478
rect 83786 709922 84022 710158
rect 80186 708362 80422 708598
rect 80186 708042 80422 708278
rect 76586 706482 76822 706718
rect 76586 706162 76822 706398
rect 65786 679018 66022 679254
rect 65786 678698 66022 678934
rect 72986 704602 73222 704838
rect 72986 704282 73222 704518
rect 72986 686218 73222 686454
rect 72986 685898 73222 686134
rect 76586 689818 76822 690054
rect 76586 689498 76822 689734
rect 80186 693418 80422 693654
rect 80186 693098 80422 693334
rect 80186 657418 80422 657654
rect 80186 657098 80422 657334
rect 101786 711182 102022 711418
rect 101786 710862 102022 711098
rect 98186 709302 98422 709538
rect 98186 708982 98422 709218
rect 94586 707422 94822 707658
rect 94586 707102 94822 707338
rect 83786 697018 84022 697254
rect 83786 696698 84022 696934
rect 83786 661018 84022 661254
rect 83786 660698 84022 660934
rect 90986 705542 91222 705778
rect 90986 705222 91222 705458
rect 90986 668218 91222 668454
rect 90986 667898 91222 668134
rect 94586 671818 94822 672054
rect 94586 671498 94822 671734
rect 98186 675418 98422 675654
rect 98186 675098 98422 675334
rect 119786 710242 120022 710478
rect 119786 709922 120022 710158
rect 116186 708362 116422 708598
rect 116186 708042 116422 708278
rect 112586 706482 112822 706718
rect 112586 706162 112822 706398
rect 101786 679018 102022 679254
rect 101786 678698 102022 678934
rect 108986 704602 109222 704838
rect 108986 704282 109222 704518
rect 108986 686218 109222 686454
rect 108986 685898 109222 686134
rect 112586 689818 112822 690054
rect 112586 689498 112822 689734
rect 116186 693418 116422 693654
rect 116186 693098 116422 693334
rect 116186 657418 116422 657654
rect 116186 657098 116422 657334
rect 137786 711182 138022 711418
rect 137786 710862 138022 711098
rect 134186 709302 134422 709538
rect 134186 708982 134422 709218
rect 130586 707422 130822 707658
rect 130586 707102 130822 707338
rect 119786 697018 120022 697254
rect 119786 696698 120022 696934
rect 119786 661018 120022 661254
rect 119786 660698 120022 660934
rect 126986 705542 127222 705778
rect 126986 705222 127222 705458
rect 126986 668218 127222 668454
rect 126986 667898 127222 668134
rect 130586 671818 130822 672054
rect 130586 671498 130822 671734
rect 134186 675418 134422 675654
rect 134186 675098 134422 675334
rect 155786 710242 156022 710478
rect 155786 709922 156022 710158
rect 152186 708362 152422 708598
rect 152186 708042 152422 708278
rect 148586 706482 148822 706718
rect 148586 706162 148822 706398
rect 137786 679018 138022 679254
rect 137786 678698 138022 678934
rect 144986 704602 145222 704838
rect 144986 704282 145222 704518
rect 144986 686218 145222 686454
rect 144986 685898 145222 686134
rect 144986 650218 145222 650454
rect 144986 649898 145222 650134
rect 136982 643018 137218 643254
rect 136982 642698 137218 642934
rect 136982 639418 137218 639654
rect 136982 639098 137218 639334
rect 136982 635818 137218 636054
rect 136982 635498 137218 635734
rect 54986 632218 55222 632454
rect 54986 631898 55222 632134
rect 136982 632218 137218 632454
rect 136982 631898 137218 632134
rect 136536 625018 136772 625254
rect 136536 624698 136772 624934
rect 136536 621418 136772 621654
rect 136536 621098 136772 621334
rect 136536 617818 136772 618054
rect 136536 617498 136772 617734
rect 136536 614218 136772 614454
rect 136536 613898 136772 614134
rect 144986 614218 145222 614454
rect 144986 613898 145222 614134
rect 136982 607018 137218 607254
rect 136982 606698 137218 606934
rect 136982 603418 137218 603654
rect 136982 603098 137218 603334
rect 136982 599818 137218 600054
rect 136982 599498 137218 599734
rect 54986 596218 55222 596454
rect 54986 595898 55222 596134
rect 136982 596218 137218 596454
rect 136982 595898 137218 596134
rect 136536 589018 136772 589254
rect 136536 588698 136772 588934
rect 136536 585418 136772 585654
rect 136536 585098 136772 585334
rect 136536 581818 136772 582054
rect 136536 581498 136772 581734
rect 60510 579052 60746 579138
rect 60510 578988 60596 579052
rect 60596 578988 60660 579052
rect 60660 578988 60746 579052
rect 60510 578902 60746 578988
rect 136536 578218 136772 578454
rect 136536 577898 136772 578134
rect 144986 578218 145222 578454
rect 144986 577898 145222 578134
rect 136982 571018 137218 571254
rect 136982 570698 137218 570934
rect 136982 567418 137218 567654
rect 136982 567098 137218 567334
rect 136982 563818 137218 564054
rect 136982 563498 137218 563734
rect 54986 560218 55222 560454
rect 54986 559898 55222 560134
rect 76586 545818 76822 546054
rect 76586 545498 76822 545734
rect 80186 549418 80422 549654
rect 80186 549098 80422 549334
rect 83786 553018 84022 553254
rect 83786 552698 84022 552934
rect 112586 545818 112822 546054
rect 112586 545498 112822 545734
rect 116186 549418 116422 549654
rect 116186 549098 116422 549334
rect 119786 553018 120022 553254
rect 119786 552698 120022 552934
rect 148586 689818 148822 690054
rect 148586 689498 148822 689734
rect 148586 653818 148822 654054
rect 148586 653498 148822 653734
rect 148586 617818 148822 618054
rect 148586 617498 148822 617734
rect 148586 581818 148822 582054
rect 148586 581498 148822 581734
rect 148586 545818 148822 546054
rect 148586 545498 148822 545734
rect 152186 693418 152422 693654
rect 152186 693098 152422 693334
rect 152186 657418 152422 657654
rect 152186 657098 152422 657334
rect 152186 621418 152422 621654
rect 152186 621098 152422 621334
rect 152186 585418 152422 585654
rect 152186 585098 152422 585334
rect 152186 549418 152422 549654
rect 152186 549098 152422 549334
rect 173786 711182 174022 711418
rect 173786 710862 174022 711098
rect 170186 709302 170422 709538
rect 170186 708982 170422 709218
rect 166586 707422 166822 707658
rect 166586 707102 166822 707338
rect 155786 697018 156022 697254
rect 155786 696698 156022 696934
rect 155786 661018 156022 661254
rect 155786 660698 156022 660934
rect 155786 625018 156022 625254
rect 155786 624698 156022 624934
rect 155786 589018 156022 589254
rect 155786 588698 156022 588934
rect 155786 553018 156022 553254
rect 155786 552698 156022 552934
rect 162986 705542 163222 705778
rect 162986 705222 163222 705458
rect 162986 668218 163222 668454
rect 162986 667898 163222 668134
rect 162986 632218 163222 632454
rect 162986 631898 163222 632134
rect 162986 596218 163222 596454
rect 162986 595898 163222 596134
rect 162986 560218 163222 560454
rect 162986 559898 163222 560134
rect 166586 671818 166822 672054
rect 166586 671498 166822 671734
rect 166586 635818 166822 636054
rect 166586 635498 166822 635734
rect 166586 599818 166822 600054
rect 166586 599498 166822 599734
rect 166586 563818 166822 564054
rect 166586 563498 166822 563734
rect 170186 675418 170422 675654
rect 170186 675098 170422 675334
rect 170186 639418 170422 639654
rect 170186 639098 170422 639334
rect 170186 603418 170422 603654
rect 170186 603098 170422 603334
rect 170186 567418 170422 567654
rect 170186 567098 170422 567334
rect 191786 710242 192022 710478
rect 191786 709922 192022 710158
rect 188186 708362 188422 708598
rect 188186 708042 188422 708278
rect 184586 706482 184822 706718
rect 184586 706162 184822 706398
rect 173786 679018 174022 679254
rect 173786 678698 174022 678934
rect 173786 643018 174022 643254
rect 173786 642698 174022 642934
rect 173786 607018 174022 607254
rect 173786 606698 174022 606934
rect 173786 571018 174022 571254
rect 173786 570698 174022 570934
rect 180986 704602 181222 704838
rect 180986 704282 181222 704518
rect 180986 686218 181222 686454
rect 180986 685898 181222 686134
rect 180986 650218 181222 650454
rect 180986 649898 181222 650134
rect 180986 614218 181222 614454
rect 180986 613898 181222 614134
rect 180986 578218 181222 578454
rect 180986 577898 181222 578134
rect 184586 689818 184822 690054
rect 184586 689498 184822 689734
rect 188186 693418 188422 693654
rect 188186 693098 188422 693334
rect 188186 657418 188422 657654
rect 188186 657098 188422 657334
rect 209786 711182 210022 711418
rect 209786 710862 210022 711098
rect 206186 709302 206422 709538
rect 206186 708982 206422 709218
rect 202586 707422 202822 707658
rect 202586 707102 202822 707338
rect 191786 697018 192022 697254
rect 191786 696698 192022 696934
rect 191786 661018 192022 661254
rect 191786 660698 192022 660934
rect 198986 705542 199222 705778
rect 198986 705222 199222 705458
rect 198986 668218 199222 668454
rect 198986 667898 199222 668134
rect 202586 671818 202822 672054
rect 202586 671498 202822 671734
rect 206186 675418 206422 675654
rect 206186 675098 206422 675334
rect 227786 710242 228022 710478
rect 227786 709922 228022 710158
rect 224186 708362 224422 708598
rect 224186 708042 224422 708278
rect 220586 706482 220822 706718
rect 220586 706162 220822 706398
rect 209786 679018 210022 679254
rect 209786 678698 210022 678934
rect 216986 704602 217222 704838
rect 216986 704282 217222 704518
rect 216986 686218 217222 686454
rect 216986 685898 217222 686134
rect 220586 689818 220822 690054
rect 220586 689498 220822 689734
rect 224186 693418 224422 693654
rect 224186 693098 224422 693334
rect 224186 657418 224422 657654
rect 224186 657098 224422 657334
rect 245786 711182 246022 711418
rect 245786 710862 246022 711098
rect 242186 709302 242422 709538
rect 242186 708982 242422 709218
rect 238586 707422 238822 707658
rect 238586 707102 238822 707338
rect 227786 697018 228022 697254
rect 227786 696698 228022 696934
rect 227786 661018 228022 661254
rect 227786 660698 228022 660934
rect 234986 705542 235222 705778
rect 234986 705222 235222 705458
rect 234986 668218 235222 668454
rect 234986 667898 235222 668134
rect 238586 671818 238822 672054
rect 238586 671498 238822 671734
rect 242186 675418 242422 675654
rect 242186 675098 242422 675334
rect 263786 710242 264022 710478
rect 263786 709922 264022 710158
rect 260186 708362 260422 708598
rect 260186 708042 260422 708278
rect 256586 706482 256822 706718
rect 256586 706162 256822 706398
rect 245786 679018 246022 679254
rect 245786 678698 246022 678934
rect 252986 704602 253222 704838
rect 252986 704282 253222 704518
rect 252986 686218 253222 686454
rect 252986 685898 253222 686134
rect 256586 689818 256822 690054
rect 256586 689498 256822 689734
rect 260186 693418 260422 693654
rect 260186 693098 260422 693334
rect 260186 657418 260422 657654
rect 260186 657098 260422 657334
rect 281786 711182 282022 711418
rect 281786 710862 282022 711098
rect 278186 709302 278422 709538
rect 278186 708982 278422 709218
rect 274586 707422 274822 707658
rect 274586 707102 274822 707338
rect 263786 697018 264022 697254
rect 263786 696698 264022 696934
rect 263786 661018 264022 661254
rect 263786 660698 264022 660934
rect 270986 705542 271222 705778
rect 270986 705222 271222 705458
rect 270986 668218 271222 668454
rect 270986 667898 271222 668134
rect 184586 653818 184822 654054
rect 184586 653498 184822 653734
rect 266982 643018 267218 643254
rect 266982 642698 267218 642934
rect 266982 639418 267218 639654
rect 266982 639098 267218 639334
rect 266982 635818 267218 636054
rect 266982 635498 267218 635734
rect 266982 632218 267218 632454
rect 266982 631898 267218 632134
rect 270986 632218 271222 632454
rect 270986 631898 271222 632134
rect 266536 625018 266772 625254
rect 266536 624698 266772 624934
rect 266536 621418 266772 621654
rect 266536 621098 266772 621334
rect 184586 617818 184822 618054
rect 184586 617498 184822 617734
rect 266536 617818 266772 618054
rect 266536 617498 266772 617734
rect 266536 614218 266772 614454
rect 266536 613898 266772 614134
rect 266982 607018 267218 607254
rect 266982 606698 267218 606934
rect 266982 603418 267218 603654
rect 266982 603098 267218 603334
rect 266982 599818 267218 600054
rect 266982 599498 267218 599734
rect 266982 596218 267218 596454
rect 266982 595898 267218 596134
rect 270986 596218 271222 596454
rect 270986 595898 271222 596134
rect 266536 589018 266772 589254
rect 266536 588698 266772 588934
rect 270270 587212 270506 587298
rect 270270 587148 270356 587212
rect 270356 587148 270420 587212
rect 270420 587148 270506 587212
rect 270270 587062 270506 587148
rect 266536 585418 266772 585654
rect 266536 585098 266772 585334
rect 184586 581818 184822 582054
rect 184586 581498 184822 581734
rect 266536 581818 266772 582054
rect 266536 581498 266772 581734
rect 188758 579052 188994 579138
rect 188758 578988 188844 579052
rect 188844 578988 188908 579052
rect 188908 578988 188994 579052
rect 188758 578902 188994 578988
rect 266536 578218 266772 578454
rect 266536 577898 266772 578134
rect 266982 571018 267218 571254
rect 266982 570698 267218 570934
rect 266982 567418 267218 567654
rect 266982 567098 267218 567334
rect 266982 563818 267218 564054
rect 266982 563498 267218 563734
rect 270986 560218 271222 560454
rect 270986 559898 271222 560134
rect 184586 545818 184822 546054
rect 184586 545498 184822 545734
rect 188186 549418 188422 549654
rect 188186 549098 188422 549334
rect 191786 553018 192022 553254
rect 191786 552698 192022 552934
rect 220586 545818 220822 546054
rect 220586 545498 220822 545734
rect 224186 549418 224422 549654
rect 224186 549098 224422 549334
rect 227786 553018 228022 553254
rect 227786 552698 228022 552934
rect 256586 545818 256822 546054
rect 256586 545498 256822 545734
rect 260186 549418 260422 549654
rect 260186 549098 260422 549334
rect 263786 553018 264022 553254
rect 263786 552698 264022 552934
rect 274586 671818 274822 672054
rect 274586 671498 274822 671734
rect 274586 635818 274822 636054
rect 274586 635498 274822 635734
rect 274586 599818 274822 600054
rect 274586 599498 274822 599734
rect 274586 563818 274822 564054
rect 274586 563498 274822 563734
rect 278186 675418 278422 675654
rect 278186 675098 278422 675334
rect 278186 639418 278422 639654
rect 278186 639098 278422 639334
rect 278186 603418 278422 603654
rect 278186 603098 278422 603334
rect 278186 567418 278422 567654
rect 278186 567098 278422 567334
rect 299786 710242 300022 710478
rect 299786 709922 300022 710158
rect 296186 708362 296422 708598
rect 296186 708042 296422 708278
rect 292586 706482 292822 706718
rect 292586 706162 292822 706398
rect 281786 679018 282022 679254
rect 281786 678698 282022 678934
rect 281786 643018 282022 643254
rect 281786 642698 282022 642934
rect 281786 607018 282022 607254
rect 281786 606698 282022 606934
rect 288986 704602 289222 704838
rect 288986 704282 289222 704518
rect 288986 686218 289222 686454
rect 288986 685898 289222 686134
rect 288986 650218 289222 650454
rect 288986 649898 289222 650134
rect 288986 614218 289222 614454
rect 288986 613898 289222 614134
rect 282414 579052 282650 579138
rect 282414 578988 282500 579052
rect 282500 578988 282564 579052
rect 282564 578988 282650 579052
rect 282414 578902 282650 578988
rect 281786 571018 282022 571254
rect 281786 570698 282022 570934
rect 288986 578218 289222 578454
rect 288986 577898 289222 578134
rect 79610 535018 79846 535254
rect 79610 534698 79846 534934
rect 79610 531418 79846 531654
rect 79610 531098 79846 531334
rect 79610 527818 79846 528054
rect 79610 527498 79846 527734
rect 54986 524218 55222 524454
rect 54986 523898 55222 524134
rect 79610 524218 79846 524454
rect 79610 523898 79846 524134
rect 64250 517018 64486 517254
rect 64250 516698 64486 516934
rect 64250 513418 64486 513654
rect 64250 513098 64486 513334
rect 64250 509818 64486 510054
rect 64250 509498 64486 509734
rect 64250 506218 64486 506454
rect 64250 505898 64486 506134
rect 79610 499018 79846 499254
rect 79610 498698 79846 498934
rect 79610 495418 79846 495654
rect 79610 495098 79846 495334
rect 79610 491818 79846 492054
rect 79610 491498 79846 491734
rect 54986 488218 55222 488454
rect 54986 487898 55222 488134
rect 79610 488218 79846 488454
rect 79610 487898 79846 488134
rect 64250 481018 64486 481254
rect 64250 480698 64486 480934
rect 64250 477418 64486 477654
rect 64250 477098 64486 477334
rect 64250 473818 64486 474054
rect 64250 473498 64486 473734
rect 64250 470218 64486 470454
rect 64250 469898 64486 470134
rect 79610 463018 79846 463254
rect 79610 462698 79846 462934
rect 79610 459418 79846 459654
rect 79610 459098 79846 459334
rect 79610 455818 79846 456054
rect 79610 455498 79846 455734
rect 54986 452218 55222 452454
rect 54986 451898 55222 452134
rect 79610 452218 79846 452454
rect 79610 451898 79846 452134
rect 64250 445018 64486 445254
rect 64250 444698 64486 444934
rect 64250 441418 64486 441654
rect 64250 441098 64486 441334
rect 64250 437818 64486 438054
rect 64250 437498 64486 437734
rect 64250 434218 64486 434454
rect 64250 433898 64486 434134
rect 79610 427018 79846 427254
rect 79610 426698 79846 426934
rect 79610 423418 79846 423654
rect 79610 423098 79846 423334
rect 79610 419818 79846 420054
rect 79610 419498 79846 419734
rect 54986 416218 55222 416454
rect 54986 415898 55222 416134
rect 79610 416218 79846 416454
rect 79610 415898 79846 416134
rect 64250 409018 64486 409254
rect 64250 408698 64486 408934
rect 64250 405418 64486 405654
rect 64250 405098 64486 405334
rect 64250 401818 64486 402054
rect 64250 401498 64486 401734
rect 64250 398218 64486 398454
rect 64250 397898 64486 398134
rect 79610 391018 79846 391254
rect 79610 390698 79846 390934
rect 79610 387418 79846 387654
rect 79610 387098 79846 387334
rect 79610 383818 79846 384054
rect 79610 383498 79846 383734
rect 54986 380218 55222 380454
rect 54986 379898 55222 380134
rect 79610 380218 79846 380454
rect 79610 379898 79846 380134
rect 64250 373018 64486 373254
rect 64250 372698 64486 372934
rect 64250 369418 64486 369654
rect 64250 369098 64486 369334
rect 64250 365818 64486 366054
rect 64250 365498 64486 365734
rect 64250 362218 64486 362454
rect 64250 361898 64486 362134
rect 79610 355018 79846 355254
rect 79610 354698 79846 354934
rect 79610 351418 79846 351654
rect 79610 351098 79846 351334
rect 79610 347818 79846 348054
rect 79610 347498 79846 347734
rect 54986 344218 55222 344454
rect 54986 343898 55222 344134
rect 79610 344218 79846 344454
rect 79610 343898 79846 344134
rect 64250 337018 64486 337254
rect 64250 336698 64486 336934
rect 64250 333418 64486 333654
rect 64250 333098 64486 333334
rect 64250 329818 64486 330054
rect 64250 329498 64486 329734
rect 64250 326218 64486 326454
rect 64250 325898 64486 326134
rect 288986 542218 289222 542454
rect 288986 541898 289222 542134
rect 288986 506218 289222 506454
rect 288986 505898 289222 506134
rect 288986 470218 289222 470454
rect 288986 469898 289222 470134
rect 288986 434218 289222 434454
rect 288986 433898 289222 434134
rect 288986 398218 289222 398454
rect 288986 397898 289222 398134
rect 288986 362218 289222 362454
rect 288986 361898 289222 362134
rect 288986 326218 289222 326454
rect 288986 325898 289222 326134
rect 54986 308218 55222 308454
rect 54986 307898 55222 308134
rect 54986 272218 55222 272454
rect 54986 271898 55222 272134
rect 54986 236218 55222 236454
rect 54986 235898 55222 236134
rect 54986 200218 55222 200454
rect 54986 199898 55222 200134
rect 54986 164218 55222 164454
rect 54986 163898 55222 164134
rect 54986 128218 55222 128454
rect 54986 127898 55222 128134
rect 54986 92218 55222 92454
rect 54986 91898 55222 92134
rect 54986 56218 55222 56454
rect 54986 55898 55222 56134
rect 54986 20218 55222 20454
rect 54986 19898 55222 20134
rect 54986 -1522 55222 -1286
rect 54986 -1842 55222 -1606
rect 58586 311818 58822 312054
rect 58586 311498 58822 311734
rect 58586 275818 58822 276054
rect 58586 275498 58822 275734
rect 58586 239818 58822 240054
rect 58586 239498 58822 239734
rect 58586 203818 58822 204054
rect 58586 203498 58822 203734
rect 58586 167818 58822 168054
rect 58586 167498 58822 167734
rect 58586 131818 58822 132054
rect 58586 131498 58822 131734
rect 58586 95818 58822 96054
rect 58586 95498 58822 95734
rect 58586 59818 58822 60054
rect 58586 59498 58822 59734
rect 58586 23818 58822 24054
rect 58586 23498 58822 23734
rect 58586 -3402 58822 -3166
rect 58586 -3722 58822 -3486
rect 62186 315418 62422 315654
rect 62186 315098 62422 315334
rect 62186 279418 62422 279654
rect 62186 279098 62422 279334
rect 62186 243418 62422 243654
rect 62186 243098 62422 243334
rect 62186 207418 62422 207654
rect 62186 207098 62422 207334
rect 62186 171418 62422 171654
rect 62186 171098 62422 171334
rect 62186 135418 62422 135654
rect 62186 135098 62422 135334
rect 62186 99418 62422 99654
rect 62186 99098 62422 99334
rect 62186 63418 62422 63654
rect 62186 63098 62422 63334
rect 62186 27418 62422 27654
rect 62186 27098 62422 27334
rect 62186 -5282 62422 -5046
rect 62186 -5602 62422 -5366
rect 65786 283018 66022 283254
rect 65786 282698 66022 282934
rect 65786 247018 66022 247254
rect 65786 246698 66022 246934
rect 65786 211018 66022 211254
rect 65786 210698 66022 210934
rect 65786 175018 66022 175254
rect 65786 174698 66022 174934
rect 65786 139018 66022 139254
rect 65786 138698 66022 138934
rect 65786 103018 66022 103254
rect 65786 102698 66022 102934
rect 65786 67018 66022 67254
rect 65786 66698 66022 66934
rect 65786 31018 66022 31254
rect 65786 30698 66022 30934
rect 47786 -6222 48022 -5986
rect 47786 -6542 48022 -6306
rect 72986 290218 73222 290454
rect 72986 289898 73222 290134
rect 72986 254218 73222 254454
rect 72986 253898 73222 254134
rect 72986 218218 73222 218454
rect 72986 217898 73222 218134
rect 72986 182218 73222 182454
rect 72986 181898 73222 182134
rect 72986 146218 73222 146454
rect 72986 145898 73222 146134
rect 72986 110218 73222 110454
rect 72986 109898 73222 110134
rect 72986 74218 73222 74454
rect 72986 73898 73222 74134
rect 72986 38218 73222 38454
rect 72986 37898 73222 38134
rect 72986 2218 73222 2454
rect 72986 1898 73222 2134
rect 72986 -582 73222 -346
rect 72986 -902 73222 -666
rect 76586 293818 76822 294054
rect 76586 293498 76822 293734
rect 76586 257818 76822 258054
rect 76586 257498 76822 257734
rect 76586 221818 76822 222054
rect 76586 221498 76822 221734
rect 76586 185818 76822 186054
rect 76586 185498 76822 185734
rect 76586 149818 76822 150054
rect 76586 149498 76822 149734
rect 76586 113818 76822 114054
rect 76586 113498 76822 113734
rect 76586 77818 76822 78054
rect 76586 77498 76822 77734
rect 76586 41818 76822 42054
rect 76586 41498 76822 41734
rect 76586 5818 76822 6054
rect 76586 5498 76822 5734
rect 76586 -2462 76822 -2226
rect 76586 -2782 76822 -2546
rect 80186 297418 80422 297654
rect 80186 297098 80422 297334
rect 80186 261418 80422 261654
rect 80186 261098 80422 261334
rect 80186 225418 80422 225654
rect 80186 225098 80422 225334
rect 80186 189418 80422 189654
rect 80186 189098 80422 189334
rect 80186 153418 80422 153654
rect 80186 153098 80422 153334
rect 80186 117418 80422 117654
rect 80186 117098 80422 117334
rect 80186 81418 80422 81654
rect 80186 81098 80422 81334
rect 80186 45418 80422 45654
rect 80186 45098 80422 45334
rect 80186 9418 80422 9654
rect 80186 9098 80422 9334
rect 80186 -4342 80422 -4106
rect 80186 -4662 80422 -4426
rect 83786 301018 84022 301254
rect 83786 300698 84022 300934
rect 83786 265018 84022 265254
rect 83786 264698 84022 264934
rect 83786 229018 84022 229254
rect 83786 228698 84022 228934
rect 83786 193018 84022 193254
rect 83786 192698 84022 192934
rect 83786 157018 84022 157254
rect 83786 156698 84022 156934
rect 83786 121018 84022 121254
rect 83786 120698 84022 120934
rect 83786 85018 84022 85254
rect 83786 84698 84022 84934
rect 83786 49018 84022 49254
rect 83786 48698 84022 48934
rect 83786 13018 84022 13254
rect 83786 12698 84022 12934
rect 65786 -7162 66022 -6926
rect 65786 -7482 66022 -7246
rect 90986 308218 91222 308454
rect 90986 307898 91222 308134
rect 90986 272218 91222 272454
rect 90986 271898 91222 272134
rect 90986 236218 91222 236454
rect 90986 235898 91222 236134
rect 90986 200218 91222 200454
rect 90986 199898 91222 200134
rect 90986 164218 91222 164454
rect 90986 163898 91222 164134
rect 90986 128218 91222 128454
rect 90986 127898 91222 128134
rect 90986 92218 91222 92454
rect 90986 91898 91222 92134
rect 90986 56218 91222 56454
rect 90986 55898 91222 56134
rect 90986 20218 91222 20454
rect 90986 19898 91222 20134
rect 90986 -1522 91222 -1286
rect 90986 -1842 91222 -1606
rect 94586 311818 94822 312054
rect 94586 311498 94822 311734
rect 94586 275818 94822 276054
rect 94586 275498 94822 275734
rect 94586 239818 94822 240054
rect 94586 239498 94822 239734
rect 94586 203818 94822 204054
rect 94586 203498 94822 203734
rect 94586 167818 94822 168054
rect 94586 167498 94822 167734
rect 94586 131818 94822 132054
rect 94586 131498 94822 131734
rect 94586 95818 94822 96054
rect 94586 95498 94822 95734
rect 94586 59818 94822 60054
rect 94586 59498 94822 59734
rect 94586 23818 94822 24054
rect 94586 23498 94822 23734
rect 94586 -3402 94822 -3166
rect 94586 -3722 94822 -3486
rect 98186 315418 98422 315654
rect 98186 315098 98422 315334
rect 98186 279418 98422 279654
rect 98186 279098 98422 279334
rect 98186 243418 98422 243654
rect 98186 243098 98422 243334
rect 98186 207418 98422 207654
rect 98186 207098 98422 207334
rect 98186 171418 98422 171654
rect 98186 171098 98422 171334
rect 98186 135418 98422 135654
rect 98186 135098 98422 135334
rect 98186 99418 98422 99654
rect 98186 99098 98422 99334
rect 98186 63418 98422 63654
rect 98186 63098 98422 63334
rect 98186 27418 98422 27654
rect 98186 27098 98422 27334
rect 98186 -5282 98422 -5046
rect 98186 -5602 98422 -5366
rect 101786 283018 102022 283254
rect 101786 282698 102022 282934
rect 101786 247018 102022 247254
rect 101786 246698 102022 246934
rect 101786 211018 102022 211254
rect 101786 210698 102022 210934
rect 101786 175018 102022 175254
rect 101786 174698 102022 174934
rect 101786 139018 102022 139254
rect 101786 138698 102022 138934
rect 101786 103018 102022 103254
rect 101786 102698 102022 102934
rect 101786 67018 102022 67254
rect 101786 66698 102022 66934
rect 101786 31018 102022 31254
rect 101786 30698 102022 30934
rect 83786 -6222 84022 -5986
rect 83786 -6542 84022 -6306
rect 108986 290218 109222 290454
rect 108986 289898 109222 290134
rect 108986 254218 109222 254454
rect 108986 253898 109222 254134
rect 108986 218218 109222 218454
rect 108986 217898 109222 218134
rect 108986 182218 109222 182454
rect 108986 181898 109222 182134
rect 108986 146218 109222 146454
rect 108986 145898 109222 146134
rect 108986 110218 109222 110454
rect 108986 109898 109222 110134
rect 108986 74218 109222 74454
rect 108986 73898 109222 74134
rect 108986 38218 109222 38454
rect 108986 37898 109222 38134
rect 108986 2218 109222 2454
rect 108986 1898 109222 2134
rect 108986 -582 109222 -346
rect 108986 -902 109222 -666
rect 112586 293818 112822 294054
rect 112586 293498 112822 293734
rect 112586 257818 112822 258054
rect 112586 257498 112822 257734
rect 112586 221818 112822 222054
rect 112586 221498 112822 221734
rect 112586 185818 112822 186054
rect 112586 185498 112822 185734
rect 112586 149818 112822 150054
rect 112586 149498 112822 149734
rect 112586 113818 112822 114054
rect 112586 113498 112822 113734
rect 112586 77818 112822 78054
rect 112586 77498 112822 77734
rect 112586 41818 112822 42054
rect 112586 41498 112822 41734
rect 112586 5818 112822 6054
rect 112586 5498 112822 5734
rect 112586 -2462 112822 -2226
rect 112586 -2782 112822 -2546
rect 116186 297418 116422 297654
rect 116186 297098 116422 297334
rect 116186 261418 116422 261654
rect 116186 261098 116422 261334
rect 116186 225418 116422 225654
rect 116186 225098 116422 225334
rect 116186 189418 116422 189654
rect 116186 189098 116422 189334
rect 116186 153418 116422 153654
rect 116186 153098 116422 153334
rect 116186 117418 116422 117654
rect 116186 117098 116422 117334
rect 116186 81418 116422 81654
rect 116186 81098 116422 81334
rect 116186 45418 116422 45654
rect 116186 45098 116422 45334
rect 116186 9418 116422 9654
rect 116186 9098 116422 9334
rect 116186 -4342 116422 -4106
rect 116186 -4662 116422 -4426
rect 119786 301018 120022 301254
rect 119786 300698 120022 300934
rect 119786 265018 120022 265254
rect 119786 264698 120022 264934
rect 119786 229018 120022 229254
rect 119786 228698 120022 228934
rect 119786 193018 120022 193254
rect 119786 192698 120022 192934
rect 119786 157018 120022 157254
rect 119786 156698 120022 156934
rect 119786 121018 120022 121254
rect 119786 120698 120022 120934
rect 119786 85018 120022 85254
rect 119786 84698 120022 84934
rect 119786 49018 120022 49254
rect 119786 48698 120022 48934
rect 119786 13018 120022 13254
rect 119786 12698 120022 12934
rect 101786 -7162 102022 -6926
rect 101786 -7482 102022 -7246
rect 126986 308218 127222 308454
rect 126986 307898 127222 308134
rect 126986 272218 127222 272454
rect 126986 271898 127222 272134
rect 126986 236218 127222 236454
rect 126986 235898 127222 236134
rect 126986 200218 127222 200454
rect 126986 199898 127222 200134
rect 126986 164218 127222 164454
rect 126986 163898 127222 164134
rect 126986 128218 127222 128454
rect 126986 127898 127222 128134
rect 126986 92218 127222 92454
rect 126986 91898 127222 92134
rect 126986 56218 127222 56454
rect 126986 55898 127222 56134
rect 126986 20218 127222 20454
rect 126986 19898 127222 20134
rect 126986 -1522 127222 -1286
rect 126986 -1842 127222 -1606
rect 130586 311818 130822 312054
rect 130586 311498 130822 311734
rect 130586 275818 130822 276054
rect 130586 275498 130822 275734
rect 130586 239818 130822 240054
rect 130586 239498 130822 239734
rect 130586 203818 130822 204054
rect 130586 203498 130822 203734
rect 130586 167818 130822 168054
rect 130586 167498 130822 167734
rect 130586 131818 130822 132054
rect 130586 131498 130822 131734
rect 130586 95818 130822 96054
rect 130586 95498 130822 95734
rect 130586 59818 130822 60054
rect 130586 59498 130822 59734
rect 130586 23818 130822 24054
rect 130586 23498 130822 23734
rect 130586 -3402 130822 -3166
rect 130586 -3722 130822 -3486
rect 134186 315418 134422 315654
rect 134186 315098 134422 315334
rect 134186 279418 134422 279654
rect 134186 279098 134422 279334
rect 134186 243418 134422 243654
rect 134186 243098 134422 243334
rect 134186 207418 134422 207654
rect 134186 207098 134422 207334
rect 134186 171418 134422 171654
rect 134186 171098 134422 171334
rect 134186 135418 134422 135654
rect 134186 135098 134422 135334
rect 134186 99418 134422 99654
rect 134186 99098 134422 99334
rect 134186 63418 134422 63654
rect 134186 63098 134422 63334
rect 134186 27418 134422 27654
rect 134186 27098 134422 27334
rect 134186 -5282 134422 -5046
rect 134186 -5602 134422 -5366
rect 137786 283018 138022 283254
rect 137786 282698 138022 282934
rect 137786 247018 138022 247254
rect 137786 246698 138022 246934
rect 137786 211018 138022 211254
rect 137786 210698 138022 210934
rect 137786 175018 138022 175254
rect 137786 174698 138022 174934
rect 137786 139018 138022 139254
rect 137786 138698 138022 138934
rect 137786 103018 138022 103254
rect 137786 102698 138022 102934
rect 137786 67018 138022 67254
rect 137786 66698 138022 66934
rect 137786 31018 138022 31254
rect 137786 30698 138022 30934
rect 119786 -6222 120022 -5986
rect 119786 -6542 120022 -6306
rect 144986 290218 145222 290454
rect 144986 289898 145222 290134
rect 144986 254218 145222 254454
rect 144986 253898 145222 254134
rect 144986 218218 145222 218454
rect 144986 217898 145222 218134
rect 144986 182218 145222 182454
rect 144986 181898 145222 182134
rect 144986 146218 145222 146454
rect 144986 145898 145222 146134
rect 144986 110218 145222 110454
rect 144986 109898 145222 110134
rect 144986 74218 145222 74454
rect 144986 73898 145222 74134
rect 144986 38218 145222 38454
rect 144986 37898 145222 38134
rect 144986 2218 145222 2454
rect 144986 1898 145222 2134
rect 144986 -582 145222 -346
rect 144986 -902 145222 -666
rect 148586 293818 148822 294054
rect 148586 293498 148822 293734
rect 148586 257818 148822 258054
rect 148586 257498 148822 257734
rect 148586 221818 148822 222054
rect 148586 221498 148822 221734
rect 148586 185818 148822 186054
rect 148586 185498 148822 185734
rect 148586 149818 148822 150054
rect 148586 149498 148822 149734
rect 148586 113818 148822 114054
rect 148586 113498 148822 113734
rect 148586 77818 148822 78054
rect 148586 77498 148822 77734
rect 148586 41818 148822 42054
rect 148586 41498 148822 41734
rect 148586 5818 148822 6054
rect 148586 5498 148822 5734
rect 148586 -2462 148822 -2226
rect 148586 -2782 148822 -2546
rect 152186 297418 152422 297654
rect 152186 297098 152422 297334
rect 152186 261418 152422 261654
rect 152186 261098 152422 261334
rect 152186 225418 152422 225654
rect 152186 225098 152422 225334
rect 152186 189418 152422 189654
rect 152186 189098 152422 189334
rect 152186 153418 152422 153654
rect 152186 153098 152422 153334
rect 152186 117418 152422 117654
rect 152186 117098 152422 117334
rect 152186 81418 152422 81654
rect 152186 81098 152422 81334
rect 152186 45418 152422 45654
rect 152186 45098 152422 45334
rect 152186 9418 152422 9654
rect 152186 9098 152422 9334
rect 152186 -4342 152422 -4106
rect 152186 -4662 152422 -4426
rect 155786 301018 156022 301254
rect 155786 300698 156022 300934
rect 155786 265018 156022 265254
rect 155786 264698 156022 264934
rect 155786 229018 156022 229254
rect 155786 228698 156022 228934
rect 155786 193018 156022 193254
rect 155786 192698 156022 192934
rect 155786 157018 156022 157254
rect 155786 156698 156022 156934
rect 155786 121018 156022 121254
rect 155786 120698 156022 120934
rect 155786 85018 156022 85254
rect 155786 84698 156022 84934
rect 155786 49018 156022 49254
rect 155786 48698 156022 48934
rect 155786 13018 156022 13254
rect 155786 12698 156022 12934
rect 137786 -7162 138022 -6926
rect 137786 -7482 138022 -7246
rect 162986 308218 163222 308454
rect 162986 307898 163222 308134
rect 162986 272218 163222 272454
rect 162986 271898 163222 272134
rect 162986 236218 163222 236454
rect 162986 235898 163222 236134
rect 162986 200218 163222 200454
rect 162986 199898 163222 200134
rect 162986 164218 163222 164454
rect 162986 163898 163222 164134
rect 162986 128218 163222 128454
rect 162986 127898 163222 128134
rect 162986 92218 163222 92454
rect 162986 91898 163222 92134
rect 162986 56218 163222 56454
rect 162986 55898 163222 56134
rect 162986 20218 163222 20454
rect 162986 19898 163222 20134
rect 162986 -1522 163222 -1286
rect 162986 -1842 163222 -1606
rect 166586 311818 166822 312054
rect 166586 311498 166822 311734
rect 166586 275818 166822 276054
rect 166586 275498 166822 275734
rect 166586 239818 166822 240054
rect 166586 239498 166822 239734
rect 166586 203818 166822 204054
rect 166586 203498 166822 203734
rect 166586 167818 166822 168054
rect 166586 167498 166822 167734
rect 166586 131818 166822 132054
rect 166586 131498 166822 131734
rect 166586 95818 166822 96054
rect 166586 95498 166822 95734
rect 166586 59818 166822 60054
rect 166586 59498 166822 59734
rect 166586 23818 166822 24054
rect 166586 23498 166822 23734
rect 166586 -3402 166822 -3166
rect 166586 -3722 166822 -3486
rect 170186 315418 170422 315654
rect 170186 315098 170422 315334
rect 170186 279418 170422 279654
rect 170186 279098 170422 279334
rect 170186 243418 170422 243654
rect 170186 243098 170422 243334
rect 170186 207418 170422 207654
rect 170186 207098 170422 207334
rect 170186 171418 170422 171654
rect 170186 171098 170422 171334
rect 170186 135418 170422 135654
rect 170186 135098 170422 135334
rect 170186 99418 170422 99654
rect 170186 99098 170422 99334
rect 170186 63418 170422 63654
rect 170186 63098 170422 63334
rect 170186 27418 170422 27654
rect 170186 27098 170422 27334
rect 170186 -5282 170422 -5046
rect 170186 -5602 170422 -5366
rect 173786 283018 174022 283254
rect 173786 282698 174022 282934
rect 173786 247018 174022 247254
rect 173786 246698 174022 246934
rect 173786 211018 174022 211254
rect 173786 210698 174022 210934
rect 173786 175018 174022 175254
rect 173786 174698 174022 174934
rect 173786 139018 174022 139254
rect 173786 138698 174022 138934
rect 173786 103018 174022 103254
rect 173786 102698 174022 102934
rect 173786 67018 174022 67254
rect 173786 66698 174022 66934
rect 173786 31018 174022 31254
rect 173786 30698 174022 30934
rect 155786 -6222 156022 -5986
rect 155786 -6542 156022 -6306
rect 180986 290218 181222 290454
rect 180986 289898 181222 290134
rect 180986 254218 181222 254454
rect 180986 253898 181222 254134
rect 180986 218218 181222 218454
rect 180986 217898 181222 218134
rect 180986 182218 181222 182454
rect 180986 181898 181222 182134
rect 180986 146218 181222 146454
rect 180986 145898 181222 146134
rect 180986 110218 181222 110454
rect 180986 109898 181222 110134
rect 180986 74218 181222 74454
rect 180986 73898 181222 74134
rect 180986 38218 181222 38454
rect 180986 37898 181222 38134
rect 180986 2218 181222 2454
rect 180986 1898 181222 2134
rect 180986 -582 181222 -346
rect 180986 -902 181222 -666
rect 184586 293818 184822 294054
rect 184586 293498 184822 293734
rect 184586 257818 184822 258054
rect 184586 257498 184822 257734
rect 184586 221818 184822 222054
rect 184586 221498 184822 221734
rect 184586 185818 184822 186054
rect 184586 185498 184822 185734
rect 184586 149818 184822 150054
rect 184586 149498 184822 149734
rect 184586 113818 184822 114054
rect 184586 113498 184822 113734
rect 184586 77818 184822 78054
rect 184586 77498 184822 77734
rect 184586 41818 184822 42054
rect 184586 41498 184822 41734
rect 184586 5818 184822 6054
rect 184586 5498 184822 5734
rect 184586 -2462 184822 -2226
rect 184586 -2782 184822 -2546
rect 188186 297418 188422 297654
rect 188186 297098 188422 297334
rect 188186 261418 188422 261654
rect 188186 261098 188422 261334
rect 188186 225418 188422 225654
rect 188186 225098 188422 225334
rect 188186 189418 188422 189654
rect 188186 189098 188422 189334
rect 188186 153418 188422 153654
rect 188186 153098 188422 153334
rect 188186 117418 188422 117654
rect 188186 117098 188422 117334
rect 188186 81418 188422 81654
rect 188186 81098 188422 81334
rect 188186 45418 188422 45654
rect 188186 45098 188422 45334
rect 188186 9418 188422 9654
rect 188186 9098 188422 9334
rect 188186 -4342 188422 -4106
rect 188186 -4662 188422 -4426
rect 191786 301018 192022 301254
rect 191786 300698 192022 300934
rect 191786 265018 192022 265254
rect 191786 264698 192022 264934
rect 191786 229018 192022 229254
rect 191786 228698 192022 228934
rect 191786 193018 192022 193254
rect 191786 192698 192022 192934
rect 191786 157018 192022 157254
rect 191786 156698 192022 156934
rect 191786 121018 192022 121254
rect 191786 120698 192022 120934
rect 191786 85018 192022 85254
rect 191786 84698 192022 84934
rect 191786 49018 192022 49254
rect 191786 48698 192022 48934
rect 191786 13018 192022 13254
rect 191786 12698 192022 12934
rect 173786 -7162 174022 -6926
rect 173786 -7482 174022 -7246
rect 198986 308218 199222 308454
rect 198986 307898 199222 308134
rect 198986 272218 199222 272454
rect 198986 271898 199222 272134
rect 198986 236218 199222 236454
rect 198986 235898 199222 236134
rect 198986 200218 199222 200454
rect 198986 199898 199222 200134
rect 198986 164218 199222 164454
rect 198986 163898 199222 164134
rect 198986 128218 199222 128454
rect 198986 127898 199222 128134
rect 198986 92218 199222 92454
rect 198986 91898 199222 92134
rect 198986 56218 199222 56454
rect 198986 55898 199222 56134
rect 198986 20218 199222 20454
rect 198986 19898 199222 20134
rect 198986 -1522 199222 -1286
rect 198986 -1842 199222 -1606
rect 202586 311818 202822 312054
rect 202586 311498 202822 311734
rect 202586 275818 202822 276054
rect 202586 275498 202822 275734
rect 202586 239818 202822 240054
rect 202586 239498 202822 239734
rect 202586 203818 202822 204054
rect 202586 203498 202822 203734
rect 202586 167818 202822 168054
rect 202586 167498 202822 167734
rect 202586 131818 202822 132054
rect 202586 131498 202822 131734
rect 202586 95818 202822 96054
rect 202586 95498 202822 95734
rect 202586 59818 202822 60054
rect 202586 59498 202822 59734
rect 202586 23818 202822 24054
rect 202586 23498 202822 23734
rect 202586 -3402 202822 -3166
rect 202586 -3722 202822 -3486
rect 206186 315418 206422 315654
rect 206186 315098 206422 315334
rect 206186 279418 206422 279654
rect 206186 279098 206422 279334
rect 206186 243418 206422 243654
rect 206186 243098 206422 243334
rect 206186 207418 206422 207654
rect 206186 207098 206422 207334
rect 206186 171418 206422 171654
rect 206186 171098 206422 171334
rect 206186 135418 206422 135654
rect 206186 135098 206422 135334
rect 206186 99418 206422 99654
rect 206186 99098 206422 99334
rect 206186 63418 206422 63654
rect 206186 63098 206422 63334
rect 206186 27418 206422 27654
rect 206186 27098 206422 27334
rect 206186 -5282 206422 -5046
rect 206186 -5602 206422 -5366
rect 209786 283018 210022 283254
rect 209786 282698 210022 282934
rect 209786 247018 210022 247254
rect 209786 246698 210022 246934
rect 209786 211018 210022 211254
rect 209786 210698 210022 210934
rect 209786 175018 210022 175254
rect 209786 174698 210022 174934
rect 209786 139018 210022 139254
rect 209786 138698 210022 138934
rect 209786 103018 210022 103254
rect 209786 102698 210022 102934
rect 209786 67018 210022 67254
rect 209786 66698 210022 66934
rect 209786 31018 210022 31254
rect 209786 30698 210022 30934
rect 191786 -6222 192022 -5986
rect 191786 -6542 192022 -6306
rect 216986 290218 217222 290454
rect 216986 289898 217222 290134
rect 216986 254218 217222 254454
rect 216986 253898 217222 254134
rect 216986 218218 217222 218454
rect 216986 217898 217222 218134
rect 216986 182218 217222 182454
rect 216986 181898 217222 182134
rect 216986 146218 217222 146454
rect 216986 145898 217222 146134
rect 216986 110218 217222 110454
rect 216986 109898 217222 110134
rect 216986 74218 217222 74454
rect 216986 73898 217222 74134
rect 216986 38218 217222 38454
rect 216986 37898 217222 38134
rect 216986 2218 217222 2454
rect 216986 1898 217222 2134
rect 216986 -582 217222 -346
rect 216986 -902 217222 -666
rect 220586 293818 220822 294054
rect 220586 293498 220822 293734
rect 220586 257818 220822 258054
rect 220586 257498 220822 257734
rect 220586 221818 220822 222054
rect 220586 221498 220822 221734
rect 220586 185818 220822 186054
rect 220586 185498 220822 185734
rect 220586 149818 220822 150054
rect 220586 149498 220822 149734
rect 220586 113818 220822 114054
rect 220586 113498 220822 113734
rect 220586 77818 220822 78054
rect 220586 77498 220822 77734
rect 220586 41818 220822 42054
rect 220586 41498 220822 41734
rect 220586 5818 220822 6054
rect 220586 5498 220822 5734
rect 220586 -2462 220822 -2226
rect 220586 -2782 220822 -2546
rect 224186 297418 224422 297654
rect 224186 297098 224422 297334
rect 224186 261418 224422 261654
rect 224186 261098 224422 261334
rect 224186 225418 224422 225654
rect 224186 225098 224422 225334
rect 224186 189418 224422 189654
rect 224186 189098 224422 189334
rect 224186 153418 224422 153654
rect 224186 153098 224422 153334
rect 224186 117418 224422 117654
rect 224186 117098 224422 117334
rect 224186 81418 224422 81654
rect 224186 81098 224422 81334
rect 224186 45418 224422 45654
rect 224186 45098 224422 45334
rect 224186 9418 224422 9654
rect 224186 9098 224422 9334
rect 224186 -4342 224422 -4106
rect 224186 -4662 224422 -4426
rect 227786 301018 228022 301254
rect 227786 300698 228022 300934
rect 227786 265018 228022 265254
rect 227786 264698 228022 264934
rect 227786 229018 228022 229254
rect 227786 228698 228022 228934
rect 227786 193018 228022 193254
rect 227786 192698 228022 192934
rect 227786 157018 228022 157254
rect 227786 156698 228022 156934
rect 227786 121018 228022 121254
rect 227786 120698 228022 120934
rect 227786 85018 228022 85254
rect 227786 84698 228022 84934
rect 227786 49018 228022 49254
rect 227786 48698 228022 48934
rect 227786 13018 228022 13254
rect 227786 12698 228022 12934
rect 209786 -7162 210022 -6926
rect 209786 -7482 210022 -7246
rect 234986 308218 235222 308454
rect 234986 307898 235222 308134
rect 234986 272218 235222 272454
rect 234986 271898 235222 272134
rect 234986 236218 235222 236454
rect 234986 235898 235222 236134
rect 234986 200218 235222 200454
rect 234986 199898 235222 200134
rect 234986 164218 235222 164454
rect 234986 163898 235222 164134
rect 234986 128218 235222 128454
rect 234986 127898 235222 128134
rect 234986 92218 235222 92454
rect 234986 91898 235222 92134
rect 234986 56218 235222 56454
rect 234986 55898 235222 56134
rect 234986 20218 235222 20454
rect 234986 19898 235222 20134
rect 234986 -1522 235222 -1286
rect 234986 -1842 235222 -1606
rect 238586 311818 238822 312054
rect 238586 311498 238822 311734
rect 238586 275818 238822 276054
rect 238586 275498 238822 275734
rect 238586 239818 238822 240054
rect 238586 239498 238822 239734
rect 238586 203818 238822 204054
rect 238586 203498 238822 203734
rect 238586 167818 238822 168054
rect 238586 167498 238822 167734
rect 238586 131818 238822 132054
rect 238586 131498 238822 131734
rect 238586 95818 238822 96054
rect 238586 95498 238822 95734
rect 238586 59818 238822 60054
rect 238586 59498 238822 59734
rect 238586 23818 238822 24054
rect 238586 23498 238822 23734
rect 238586 -3402 238822 -3166
rect 238586 -3722 238822 -3486
rect 242186 315418 242422 315654
rect 242186 315098 242422 315334
rect 242186 279418 242422 279654
rect 242186 279098 242422 279334
rect 242186 243418 242422 243654
rect 242186 243098 242422 243334
rect 242186 207418 242422 207654
rect 242186 207098 242422 207334
rect 242186 171418 242422 171654
rect 242186 171098 242422 171334
rect 242186 135418 242422 135654
rect 242186 135098 242422 135334
rect 242186 99418 242422 99654
rect 242186 99098 242422 99334
rect 242186 63418 242422 63654
rect 242186 63098 242422 63334
rect 242186 27418 242422 27654
rect 242186 27098 242422 27334
rect 242186 -5282 242422 -5046
rect 242186 -5602 242422 -5366
rect 245786 283018 246022 283254
rect 245786 282698 246022 282934
rect 245786 247018 246022 247254
rect 245786 246698 246022 246934
rect 245786 211018 246022 211254
rect 245786 210698 246022 210934
rect 245786 175018 246022 175254
rect 245786 174698 246022 174934
rect 245786 139018 246022 139254
rect 245786 138698 246022 138934
rect 245786 103018 246022 103254
rect 245786 102698 246022 102934
rect 245786 67018 246022 67254
rect 245786 66698 246022 66934
rect 245786 31018 246022 31254
rect 245786 30698 246022 30934
rect 227786 -6222 228022 -5986
rect 227786 -6542 228022 -6306
rect 252986 290218 253222 290454
rect 252986 289898 253222 290134
rect 252986 254218 253222 254454
rect 252986 253898 253222 254134
rect 252986 218218 253222 218454
rect 252986 217898 253222 218134
rect 252986 182218 253222 182454
rect 252986 181898 253222 182134
rect 252986 146218 253222 146454
rect 252986 145898 253222 146134
rect 252986 110218 253222 110454
rect 252986 109898 253222 110134
rect 252986 74218 253222 74454
rect 252986 73898 253222 74134
rect 252986 38218 253222 38454
rect 252986 37898 253222 38134
rect 252986 2218 253222 2454
rect 252986 1898 253222 2134
rect 252986 -582 253222 -346
rect 252986 -902 253222 -666
rect 256586 293818 256822 294054
rect 256586 293498 256822 293734
rect 256586 257818 256822 258054
rect 256586 257498 256822 257734
rect 256586 221818 256822 222054
rect 256586 221498 256822 221734
rect 256586 185818 256822 186054
rect 256586 185498 256822 185734
rect 256586 149818 256822 150054
rect 256586 149498 256822 149734
rect 256586 113818 256822 114054
rect 256586 113498 256822 113734
rect 256586 77818 256822 78054
rect 256586 77498 256822 77734
rect 256586 41818 256822 42054
rect 256586 41498 256822 41734
rect 256586 5818 256822 6054
rect 256586 5498 256822 5734
rect 256586 -2462 256822 -2226
rect 256586 -2782 256822 -2546
rect 260186 297418 260422 297654
rect 260186 297098 260422 297334
rect 260186 261418 260422 261654
rect 260186 261098 260422 261334
rect 260186 225418 260422 225654
rect 260186 225098 260422 225334
rect 260186 189418 260422 189654
rect 260186 189098 260422 189334
rect 260186 153418 260422 153654
rect 260186 153098 260422 153334
rect 260186 117418 260422 117654
rect 260186 117098 260422 117334
rect 260186 81418 260422 81654
rect 260186 81098 260422 81334
rect 260186 45418 260422 45654
rect 260186 45098 260422 45334
rect 260186 9418 260422 9654
rect 260186 9098 260422 9334
rect 260186 -4342 260422 -4106
rect 260186 -4662 260422 -4426
rect 263786 301018 264022 301254
rect 263786 300698 264022 300934
rect 263786 265018 264022 265254
rect 263786 264698 264022 264934
rect 263786 229018 264022 229254
rect 263786 228698 264022 228934
rect 263786 193018 264022 193254
rect 263786 192698 264022 192934
rect 263786 157018 264022 157254
rect 263786 156698 264022 156934
rect 263786 121018 264022 121254
rect 263786 120698 264022 120934
rect 263786 85018 264022 85254
rect 263786 84698 264022 84934
rect 263786 49018 264022 49254
rect 263786 48698 264022 48934
rect 263786 13018 264022 13254
rect 263786 12698 264022 12934
rect 245786 -7162 246022 -6926
rect 245786 -7482 246022 -7246
rect 270986 308218 271222 308454
rect 270986 307898 271222 308134
rect 270986 272218 271222 272454
rect 270986 271898 271222 272134
rect 270986 236218 271222 236454
rect 270986 235898 271222 236134
rect 270986 200218 271222 200454
rect 270986 199898 271222 200134
rect 270986 164218 271222 164454
rect 270986 163898 271222 164134
rect 270986 128218 271222 128454
rect 270986 127898 271222 128134
rect 270986 92218 271222 92454
rect 270986 91898 271222 92134
rect 270986 56218 271222 56454
rect 270986 55898 271222 56134
rect 270986 20218 271222 20454
rect 270986 19898 271222 20134
rect 270986 -1522 271222 -1286
rect 270986 -1842 271222 -1606
rect 274586 311818 274822 312054
rect 274586 311498 274822 311734
rect 274586 275818 274822 276054
rect 274586 275498 274822 275734
rect 274586 239818 274822 240054
rect 274586 239498 274822 239734
rect 274586 203818 274822 204054
rect 274586 203498 274822 203734
rect 274586 167818 274822 168054
rect 274586 167498 274822 167734
rect 274586 131818 274822 132054
rect 274586 131498 274822 131734
rect 274586 95818 274822 96054
rect 274586 95498 274822 95734
rect 274586 59818 274822 60054
rect 274586 59498 274822 59734
rect 274586 23818 274822 24054
rect 274586 23498 274822 23734
rect 274586 -3402 274822 -3166
rect 274586 -3722 274822 -3486
rect 278186 315418 278422 315654
rect 278186 315098 278422 315334
rect 278186 279418 278422 279654
rect 278186 279098 278422 279334
rect 278186 243418 278422 243654
rect 278186 243098 278422 243334
rect 278186 207418 278422 207654
rect 278186 207098 278422 207334
rect 278186 171418 278422 171654
rect 278186 171098 278422 171334
rect 278186 135418 278422 135654
rect 278186 135098 278422 135334
rect 278186 99418 278422 99654
rect 278186 99098 278422 99334
rect 278186 63418 278422 63654
rect 278186 63098 278422 63334
rect 278186 27418 278422 27654
rect 278186 27098 278422 27334
rect 278186 -5282 278422 -5046
rect 278186 -5602 278422 -5366
rect 281786 283018 282022 283254
rect 281786 282698 282022 282934
rect 281786 247018 282022 247254
rect 281786 246698 282022 246934
rect 281786 211018 282022 211254
rect 281786 210698 282022 210934
rect 281786 175018 282022 175254
rect 281786 174698 282022 174934
rect 281786 139018 282022 139254
rect 281786 138698 282022 138934
rect 281786 103018 282022 103254
rect 281786 102698 282022 102934
rect 281786 67018 282022 67254
rect 281786 66698 282022 66934
rect 281786 31018 282022 31254
rect 281786 30698 282022 30934
rect 263786 -6222 264022 -5986
rect 263786 -6542 264022 -6306
rect 288986 290218 289222 290454
rect 288986 289898 289222 290134
rect 288986 254218 289222 254454
rect 288986 253898 289222 254134
rect 288986 218218 289222 218454
rect 288986 217898 289222 218134
rect 288986 182218 289222 182454
rect 288986 181898 289222 182134
rect 288986 146218 289222 146454
rect 288986 145898 289222 146134
rect 288986 110218 289222 110454
rect 288986 109898 289222 110134
rect 288986 74218 289222 74454
rect 288986 73898 289222 74134
rect 288986 38218 289222 38454
rect 288986 37898 289222 38134
rect 288986 2218 289222 2454
rect 288986 1898 289222 2134
rect 288986 -582 289222 -346
rect 288986 -902 289222 -666
rect 292586 689818 292822 690054
rect 292586 689498 292822 689734
rect 292586 653818 292822 654054
rect 292586 653498 292822 653734
rect 292586 617818 292822 618054
rect 292586 617498 292822 617734
rect 292586 581818 292822 582054
rect 292586 581498 292822 581734
rect 292586 545818 292822 546054
rect 292586 545498 292822 545734
rect 292586 509818 292822 510054
rect 292586 509498 292822 509734
rect 292586 473818 292822 474054
rect 292586 473498 292822 473734
rect 292586 437818 292822 438054
rect 292586 437498 292822 437734
rect 292586 401818 292822 402054
rect 292586 401498 292822 401734
rect 292586 365818 292822 366054
rect 292586 365498 292822 365734
rect 292586 329818 292822 330054
rect 292586 329498 292822 329734
rect 292586 293818 292822 294054
rect 292586 293498 292822 293734
rect 292586 257818 292822 258054
rect 292586 257498 292822 257734
rect 292586 221818 292822 222054
rect 292586 221498 292822 221734
rect 292586 185818 292822 186054
rect 292586 185498 292822 185734
rect 292586 149818 292822 150054
rect 292586 149498 292822 149734
rect 292586 113818 292822 114054
rect 292586 113498 292822 113734
rect 292586 77818 292822 78054
rect 292586 77498 292822 77734
rect 292586 41818 292822 42054
rect 292586 41498 292822 41734
rect 292586 5818 292822 6054
rect 292586 5498 292822 5734
rect 292586 -2462 292822 -2226
rect 292586 -2782 292822 -2546
rect 296186 693418 296422 693654
rect 296186 693098 296422 693334
rect 296186 657418 296422 657654
rect 296186 657098 296422 657334
rect 296186 621418 296422 621654
rect 296186 621098 296422 621334
rect 296186 585418 296422 585654
rect 296186 585098 296422 585334
rect 296186 549418 296422 549654
rect 296186 549098 296422 549334
rect 296186 513418 296422 513654
rect 296186 513098 296422 513334
rect 296186 477418 296422 477654
rect 296186 477098 296422 477334
rect 296186 441418 296422 441654
rect 296186 441098 296422 441334
rect 296186 405418 296422 405654
rect 296186 405098 296422 405334
rect 296186 369418 296422 369654
rect 296186 369098 296422 369334
rect 296186 333418 296422 333654
rect 296186 333098 296422 333334
rect 296186 297418 296422 297654
rect 296186 297098 296422 297334
rect 296186 261418 296422 261654
rect 296186 261098 296422 261334
rect 296186 225418 296422 225654
rect 296186 225098 296422 225334
rect 296186 189418 296422 189654
rect 296186 189098 296422 189334
rect 296186 153418 296422 153654
rect 296186 153098 296422 153334
rect 296186 117418 296422 117654
rect 296186 117098 296422 117334
rect 296186 81418 296422 81654
rect 296186 81098 296422 81334
rect 296186 45418 296422 45654
rect 296186 45098 296422 45334
rect 296186 9418 296422 9654
rect 296186 9098 296422 9334
rect 296186 -4342 296422 -4106
rect 296186 -4662 296422 -4426
rect 317786 711182 318022 711418
rect 317786 710862 318022 711098
rect 314186 709302 314422 709538
rect 314186 708982 314422 709218
rect 310586 707422 310822 707658
rect 310586 707102 310822 707338
rect 299786 697018 300022 697254
rect 299786 696698 300022 696934
rect 299786 661018 300022 661254
rect 299786 660698 300022 660934
rect 306986 705542 307222 705778
rect 306986 705222 307222 705458
rect 306986 668218 307222 668454
rect 306986 667898 307222 668134
rect 310586 671818 310822 672054
rect 310586 671498 310822 671734
rect 314186 675418 314422 675654
rect 314186 675098 314422 675334
rect 335786 710242 336022 710478
rect 335786 709922 336022 710158
rect 332186 708362 332422 708598
rect 332186 708042 332422 708278
rect 328586 706482 328822 706718
rect 328586 706162 328822 706398
rect 317786 679018 318022 679254
rect 317786 678698 318022 678934
rect 324986 704602 325222 704838
rect 324986 704282 325222 704518
rect 324986 686218 325222 686454
rect 324986 685898 325222 686134
rect 328586 689818 328822 690054
rect 328586 689498 328822 689734
rect 332186 693418 332422 693654
rect 332186 693098 332422 693334
rect 332186 657418 332422 657654
rect 332186 657098 332422 657334
rect 353786 711182 354022 711418
rect 353786 710862 354022 711098
rect 350186 709302 350422 709538
rect 350186 708982 350422 709218
rect 346586 707422 346822 707658
rect 346586 707102 346822 707338
rect 335786 697018 336022 697254
rect 335786 696698 336022 696934
rect 335786 661018 336022 661254
rect 335786 660698 336022 660934
rect 342986 705542 343222 705778
rect 342986 705222 343222 705458
rect 342986 668218 343222 668454
rect 342986 667898 343222 668134
rect 346586 671818 346822 672054
rect 346586 671498 346822 671734
rect 350186 675418 350422 675654
rect 350186 675098 350422 675334
rect 371786 710242 372022 710478
rect 371786 709922 372022 710158
rect 368186 708362 368422 708598
rect 368186 708042 368422 708278
rect 364586 706482 364822 706718
rect 364586 706162 364822 706398
rect 353786 679018 354022 679254
rect 353786 678698 354022 678934
rect 360986 704602 361222 704838
rect 360986 704282 361222 704518
rect 360986 686218 361222 686454
rect 360986 685898 361222 686134
rect 364586 689818 364822 690054
rect 364586 689498 364822 689734
rect 368186 693418 368422 693654
rect 368186 693098 368422 693334
rect 368186 657418 368422 657654
rect 368186 657098 368422 657334
rect 389786 711182 390022 711418
rect 389786 710862 390022 711098
rect 386186 709302 386422 709538
rect 386186 708982 386422 709218
rect 382586 707422 382822 707658
rect 382586 707102 382822 707338
rect 371786 697018 372022 697254
rect 371786 696698 372022 696934
rect 371786 661018 372022 661254
rect 371786 660698 372022 660934
rect 378986 705542 379222 705778
rect 378986 705222 379222 705458
rect 378986 668218 379222 668454
rect 378986 667898 379222 668134
rect 382586 671818 382822 672054
rect 382586 671498 382822 671734
rect 386186 675418 386422 675654
rect 386186 675098 386422 675334
rect 407786 710242 408022 710478
rect 407786 709922 408022 710158
rect 404186 708362 404422 708598
rect 404186 708042 404422 708278
rect 400586 706482 400822 706718
rect 400586 706162 400822 706398
rect 389786 679018 390022 679254
rect 389786 678698 390022 678934
rect 396986 704602 397222 704838
rect 396986 704282 397222 704518
rect 396986 686218 397222 686454
rect 396986 685898 397222 686134
rect 396986 650218 397222 650454
rect 396986 649898 397222 650134
rect 386982 643018 387218 643254
rect 386982 642698 387218 642934
rect 386982 639418 387218 639654
rect 386982 639098 387218 639334
rect 386982 635818 387218 636054
rect 386982 635498 387218 635734
rect 386982 632218 387218 632454
rect 386982 631898 387218 632134
rect 299786 625018 300022 625254
rect 299786 624698 300022 624934
rect 386536 625018 386772 625254
rect 386536 624698 386772 624934
rect 386536 621418 386772 621654
rect 386536 621098 386772 621334
rect 386536 617818 386772 618054
rect 386536 617498 386772 617734
rect 386536 614218 386772 614454
rect 386536 613898 386772 614134
rect 396986 614218 397222 614454
rect 396986 613898 397222 614134
rect 386982 607018 387218 607254
rect 386982 606698 387218 606934
rect 386982 603418 387218 603654
rect 386982 603098 387218 603334
rect 386982 599818 387218 600054
rect 386982 599498 387218 599734
rect 386982 596218 387218 596454
rect 386982 595898 387218 596134
rect 299786 589018 300022 589254
rect 299786 588698 300022 588934
rect 386536 589018 386772 589254
rect 386536 588698 386772 588934
rect 387478 587212 387714 587298
rect 387478 587148 387564 587212
rect 387564 587148 387628 587212
rect 387628 587148 387714 587212
rect 387478 587062 387714 587148
rect 386536 585418 386772 585654
rect 386536 585098 386772 585334
rect 386536 581818 386772 582054
rect 386536 581498 386772 581734
rect 389134 579582 389370 579818
rect 310198 579052 310434 579138
rect 310198 578988 310284 579052
rect 310284 578988 310348 579052
rect 310348 578988 310434 579052
rect 310198 578902 310434 578988
rect 386536 578218 386772 578454
rect 386536 577898 386772 578134
rect 396986 578218 397222 578454
rect 396986 577898 397222 578134
rect 386982 571018 387218 571254
rect 386982 570698 387218 570934
rect 386982 567418 387218 567654
rect 386982 567098 387218 567334
rect 386982 563818 387218 564054
rect 386982 563498 387218 563734
rect 299786 553018 300022 553254
rect 299786 552698 300022 552934
rect 299786 517018 300022 517254
rect 299786 516698 300022 516934
rect 299786 481018 300022 481254
rect 299786 480698 300022 480934
rect 299786 445018 300022 445254
rect 299786 444698 300022 444934
rect 299786 409018 300022 409254
rect 299786 408698 300022 408934
rect 299786 373018 300022 373254
rect 299786 372698 300022 372934
rect 299786 337018 300022 337254
rect 299786 336698 300022 336934
rect 306986 524218 307222 524454
rect 306986 523898 307222 524134
rect 306986 488218 307222 488454
rect 306986 487898 307222 488134
rect 306986 452218 307222 452454
rect 306986 451898 307222 452134
rect 306986 416218 307222 416454
rect 306986 415898 307222 416134
rect 306986 380218 307222 380454
rect 306986 379898 307222 380134
rect 306986 344218 307222 344454
rect 306986 343898 307222 344134
rect 306986 308218 307222 308454
rect 306986 307898 307222 308134
rect 310586 527818 310822 528054
rect 310586 527498 310822 527734
rect 310586 491818 310822 492054
rect 310586 491498 310822 491734
rect 310586 455818 310822 456054
rect 310586 455498 310822 455734
rect 310586 419818 310822 420054
rect 310586 419498 310822 419734
rect 310586 383818 310822 384054
rect 310586 383498 310822 383734
rect 310586 347818 310822 348054
rect 310586 347498 310822 347734
rect 310586 311818 310822 312054
rect 310586 311498 310822 311734
rect 314186 531418 314422 531654
rect 314186 531098 314422 531334
rect 314186 495418 314422 495654
rect 314186 495098 314422 495334
rect 314186 459418 314422 459654
rect 314186 459098 314422 459334
rect 314186 423418 314422 423654
rect 314186 423098 314422 423334
rect 314186 387418 314422 387654
rect 314186 387098 314422 387334
rect 314186 351418 314422 351654
rect 314186 351098 314422 351334
rect 314186 315418 314422 315654
rect 314186 315098 314422 315334
rect 317786 535018 318022 535254
rect 317786 534698 318022 534934
rect 317786 499018 318022 499254
rect 317786 498698 318022 498934
rect 317786 463018 318022 463254
rect 317786 462698 318022 462934
rect 317786 427018 318022 427254
rect 317786 426698 318022 426934
rect 317786 391018 318022 391254
rect 317786 390698 318022 390934
rect 317786 355018 318022 355254
rect 317786 354698 318022 354934
rect 317786 319018 318022 319254
rect 317786 318698 318022 318934
rect 324986 542218 325222 542454
rect 324986 541898 325222 542134
rect 324986 506218 325222 506454
rect 324986 505898 325222 506134
rect 324986 470218 325222 470454
rect 324986 469898 325222 470134
rect 324986 434218 325222 434454
rect 324986 433898 325222 434134
rect 324986 398218 325222 398454
rect 324986 397898 325222 398134
rect 324986 362218 325222 362454
rect 324986 361898 325222 362134
rect 324986 326218 325222 326454
rect 324986 325898 325222 326134
rect 328586 545818 328822 546054
rect 328586 545498 328822 545734
rect 328586 509818 328822 510054
rect 328586 509498 328822 509734
rect 328586 473818 328822 474054
rect 328586 473498 328822 473734
rect 328586 437818 328822 438054
rect 328586 437498 328822 437734
rect 328586 401818 328822 402054
rect 328586 401498 328822 401734
rect 328586 365818 328822 366054
rect 328586 365498 328822 365734
rect 328586 329818 328822 330054
rect 328586 329498 328822 329734
rect 332186 549418 332422 549654
rect 332186 549098 332422 549334
rect 332186 513418 332422 513654
rect 332186 513098 332422 513334
rect 332186 477418 332422 477654
rect 332186 477098 332422 477334
rect 332186 441418 332422 441654
rect 332186 441098 332422 441334
rect 332186 405418 332422 405654
rect 332186 405098 332422 405334
rect 332186 369418 332422 369654
rect 332186 369098 332422 369334
rect 332186 333418 332422 333654
rect 332186 333098 332422 333334
rect 335786 553018 336022 553254
rect 335786 552698 336022 552934
rect 335786 517018 336022 517254
rect 335786 516698 336022 516934
rect 335786 481018 336022 481254
rect 335786 480698 336022 480934
rect 335786 445018 336022 445254
rect 335786 444698 336022 444934
rect 342986 524218 343222 524454
rect 342986 523898 343222 524134
rect 342986 488218 343222 488454
rect 342986 487898 343222 488134
rect 342986 452218 343222 452454
rect 342986 451898 343222 452134
rect 342986 416218 343222 416454
rect 342986 415898 343222 416134
rect 346586 527818 346822 528054
rect 346586 527498 346822 527734
rect 346586 491818 346822 492054
rect 346586 491498 346822 491734
rect 346586 455818 346822 456054
rect 346586 455498 346822 455734
rect 346586 419818 346822 420054
rect 346586 419498 346822 419734
rect 350186 531418 350422 531654
rect 350186 531098 350422 531334
rect 350186 495418 350422 495654
rect 350186 495098 350422 495334
rect 350186 459418 350422 459654
rect 350186 459098 350422 459334
rect 350186 423418 350422 423654
rect 350186 423098 350422 423334
rect 353786 535018 354022 535254
rect 353786 534698 354022 534934
rect 353786 499018 354022 499254
rect 353786 498698 354022 498934
rect 353786 463018 354022 463254
rect 353786 462698 354022 462934
rect 353786 427018 354022 427254
rect 353786 426698 354022 426934
rect 360986 542218 361222 542454
rect 360986 541898 361222 542134
rect 360986 506218 361222 506454
rect 360986 505898 361222 506134
rect 360986 470218 361222 470454
rect 360986 469898 361222 470134
rect 360986 434218 361222 434454
rect 360986 433898 361222 434134
rect 364586 545818 364822 546054
rect 364586 545498 364822 545734
rect 364586 509818 364822 510054
rect 364586 509498 364822 509734
rect 364586 473818 364822 474054
rect 364586 473498 364822 473734
rect 364586 437818 364822 438054
rect 364586 437498 364822 437734
rect 368186 549418 368422 549654
rect 368186 549098 368422 549334
rect 368186 513418 368422 513654
rect 368186 513098 368422 513334
rect 368186 477418 368422 477654
rect 368186 477098 368422 477334
rect 368186 441418 368422 441654
rect 368186 441098 368422 441334
rect 371786 553018 372022 553254
rect 371786 552698 372022 552934
rect 371786 517018 372022 517254
rect 371786 516698 372022 516934
rect 371786 481018 372022 481254
rect 371786 480698 372022 480934
rect 371786 445018 372022 445254
rect 371786 444698 372022 444934
rect 378986 524218 379222 524454
rect 378986 523898 379222 524134
rect 378986 488218 379222 488454
rect 378986 487898 379222 488134
rect 378986 452218 379222 452454
rect 378986 451898 379222 452134
rect 378986 416218 379222 416454
rect 378986 415898 379222 416134
rect 382586 527818 382822 528054
rect 382586 527498 382822 527734
rect 382586 491818 382822 492054
rect 382586 491498 382822 491734
rect 382586 455818 382822 456054
rect 382586 455498 382822 455734
rect 382586 419818 382822 420054
rect 382586 419498 382822 419734
rect 386186 531418 386422 531654
rect 386186 531098 386422 531334
rect 386186 495418 386422 495654
rect 386186 495098 386422 495334
rect 386186 459418 386422 459654
rect 386186 459098 386422 459334
rect 386186 423418 386422 423654
rect 386186 423098 386422 423334
rect 389786 535018 390022 535254
rect 389786 534698 390022 534934
rect 389786 499018 390022 499254
rect 389786 498698 390022 498934
rect 389786 463018 390022 463254
rect 389786 462698 390022 462934
rect 389786 427018 390022 427254
rect 389786 426698 390022 426934
rect 396986 542218 397222 542454
rect 396986 541898 397222 542134
rect 396986 506218 397222 506454
rect 396986 505898 397222 506134
rect 396986 470218 397222 470454
rect 396986 469898 397222 470134
rect 396986 434218 397222 434454
rect 396986 433898 397222 434134
rect 400586 689818 400822 690054
rect 400586 689498 400822 689734
rect 400586 653818 400822 654054
rect 400586 653498 400822 653734
rect 400586 617818 400822 618054
rect 400586 617498 400822 617734
rect 400586 581818 400822 582054
rect 400586 581498 400822 581734
rect 400586 545818 400822 546054
rect 400586 545498 400822 545734
rect 400586 509818 400822 510054
rect 400586 509498 400822 509734
rect 400586 473818 400822 474054
rect 400586 473498 400822 473734
rect 400586 437818 400822 438054
rect 400586 437498 400822 437734
rect 404186 693418 404422 693654
rect 404186 693098 404422 693334
rect 404186 657418 404422 657654
rect 404186 657098 404422 657334
rect 404186 621418 404422 621654
rect 404186 621098 404422 621334
rect 404186 585418 404422 585654
rect 404186 585098 404422 585334
rect 404186 549418 404422 549654
rect 404186 549098 404422 549334
rect 404186 513418 404422 513654
rect 404186 513098 404422 513334
rect 404186 477418 404422 477654
rect 404186 477098 404422 477334
rect 404186 441418 404422 441654
rect 404186 441098 404422 441334
rect 425786 711182 426022 711418
rect 425786 710862 426022 711098
rect 422186 709302 422422 709538
rect 422186 708982 422422 709218
rect 418586 707422 418822 707658
rect 418586 707102 418822 707338
rect 407786 697018 408022 697254
rect 407786 696698 408022 696934
rect 407786 661018 408022 661254
rect 407786 660698 408022 660934
rect 407786 625018 408022 625254
rect 407786 624698 408022 624934
rect 407786 589018 408022 589254
rect 407786 588698 408022 588934
rect 407786 553018 408022 553254
rect 407786 552698 408022 552934
rect 407786 517018 408022 517254
rect 407786 516698 408022 516934
rect 407786 481018 408022 481254
rect 407786 480698 408022 480934
rect 407786 445018 408022 445254
rect 407786 444698 408022 444934
rect 414986 705542 415222 705778
rect 414986 705222 415222 705458
rect 414986 668218 415222 668454
rect 414986 667898 415222 668134
rect 414986 632218 415222 632454
rect 414986 631898 415222 632134
rect 414986 596218 415222 596454
rect 414986 595898 415222 596134
rect 414986 560218 415222 560454
rect 414986 559898 415222 560134
rect 414986 524218 415222 524454
rect 414986 523898 415222 524134
rect 414986 488218 415222 488454
rect 414986 487898 415222 488134
rect 414986 452218 415222 452454
rect 414986 451898 415222 452134
rect 414986 416218 415222 416454
rect 414986 415898 415222 416134
rect 418586 671818 418822 672054
rect 418586 671498 418822 671734
rect 418586 635818 418822 636054
rect 418586 635498 418822 635734
rect 418586 599818 418822 600054
rect 418586 599498 418822 599734
rect 418586 563818 418822 564054
rect 418586 563498 418822 563734
rect 418586 527818 418822 528054
rect 418586 527498 418822 527734
rect 418586 491818 418822 492054
rect 418586 491498 418822 491734
rect 418586 455818 418822 456054
rect 418586 455498 418822 455734
rect 418586 419818 418822 420054
rect 418586 419498 418822 419734
rect 422186 675418 422422 675654
rect 422186 675098 422422 675334
rect 422186 639418 422422 639654
rect 422186 639098 422422 639334
rect 422186 603418 422422 603654
rect 422186 603098 422422 603334
rect 422186 567418 422422 567654
rect 422186 567098 422422 567334
rect 422186 531418 422422 531654
rect 422186 531098 422422 531334
rect 422186 495418 422422 495654
rect 422186 495098 422422 495334
rect 422186 459418 422422 459654
rect 422186 459098 422422 459334
rect 422186 423418 422422 423654
rect 422186 423098 422422 423334
rect 335786 409018 336022 409254
rect 335786 408698 336022 408934
rect 340524 409018 340760 409254
rect 340524 408698 340760 408934
rect 340524 405418 340760 405654
rect 340524 405098 340760 405334
rect 340524 401818 340760 402054
rect 340524 401498 340760 401734
rect 340524 398218 340760 398454
rect 340524 397898 340760 398134
rect 340078 391018 340314 391254
rect 340078 390698 340314 390934
rect 340078 387418 340314 387654
rect 340078 387098 340314 387334
rect 422186 387418 422422 387654
rect 422186 387098 422422 387334
rect 340078 383818 340314 384054
rect 340078 383498 340314 383734
rect 340078 380218 340314 380454
rect 340078 379898 340314 380134
rect 335786 373018 336022 373254
rect 335786 372698 336022 372934
rect 340524 373018 340760 373254
rect 340524 372698 340760 372934
rect 340524 369418 340760 369654
rect 340524 369098 340760 369334
rect 340524 365818 340760 366054
rect 340524 365498 340760 365734
rect 340524 362218 340760 362454
rect 340524 361898 340760 362134
rect 340078 355018 340314 355254
rect 340078 354698 340314 354934
rect 340078 351418 340314 351654
rect 340078 351098 340314 351334
rect 422186 351418 422422 351654
rect 422186 351098 422422 351334
rect 420598 349212 420834 349298
rect 420598 349148 420684 349212
rect 420684 349148 420748 349212
rect 420748 349148 420834 349212
rect 420598 349062 420834 349148
rect 340078 347818 340314 348054
rect 340078 347498 340314 347734
rect 419862 346564 419948 346578
rect 419948 346564 420012 346578
rect 420012 346564 420098 346578
rect 419862 346342 420098 346564
rect 420598 346492 420834 346578
rect 420598 346428 420684 346492
rect 420684 346428 420748 346492
rect 420748 346428 420834 346492
rect 420598 346342 420834 346428
rect 340078 344218 340314 344454
rect 340078 343898 340314 344134
rect 420598 342942 420834 343178
rect 420414 341732 420650 341818
rect 420414 341668 420500 341732
rect 420500 341668 420564 341732
rect 420564 341668 420650 341732
rect 420414 341582 420650 341668
rect 420414 341052 420650 341138
rect 420414 340988 420500 341052
rect 420500 340988 420564 341052
rect 420564 340988 420650 341052
rect 420414 340902 420650 340988
rect 335786 337018 336022 337254
rect 335786 336698 336022 336934
rect 340524 337018 340760 337254
rect 340524 336698 340760 336934
rect 340524 333418 340760 333654
rect 340524 333098 340760 333334
rect 340524 329818 340760 330054
rect 340524 329498 340760 329734
rect 340524 326218 340760 326454
rect 340524 325898 340760 326134
rect 342986 308218 343222 308454
rect 342986 307898 343222 308134
rect 346586 311818 346822 312054
rect 346586 311498 346822 311734
rect 350186 315418 350422 315654
rect 350186 315098 350422 315334
rect 378986 308218 379222 308454
rect 378986 307898 379222 308134
rect 382586 311818 382822 312054
rect 382586 311498 382822 311734
rect 386186 315418 386422 315654
rect 386186 315098 386422 315334
rect 414986 308218 415222 308454
rect 414986 307898 415222 308134
rect 418586 311818 418822 312054
rect 418586 311498 418822 311734
rect 443786 710242 444022 710478
rect 443786 709922 444022 710158
rect 440186 708362 440422 708598
rect 440186 708042 440422 708278
rect 436586 706482 436822 706718
rect 436586 706162 436822 706398
rect 425786 679018 426022 679254
rect 425786 678698 426022 678934
rect 425786 643018 426022 643254
rect 425786 642698 426022 642934
rect 425786 607018 426022 607254
rect 425786 606698 426022 606934
rect 425786 571018 426022 571254
rect 425786 570698 426022 570934
rect 425786 535018 426022 535254
rect 425786 534698 426022 534934
rect 425786 499018 426022 499254
rect 425786 498698 426022 498934
rect 425786 463018 426022 463254
rect 425786 462698 426022 462934
rect 425786 427018 426022 427254
rect 425786 426698 426022 426934
rect 425786 391018 426022 391254
rect 425786 390698 426022 390934
rect 425786 355018 426022 355254
rect 425786 354698 426022 354934
rect 422806 346492 423042 346578
rect 422806 346428 422892 346492
rect 422892 346428 422956 346492
rect 422956 346428 423042 346492
rect 422806 346342 423042 346428
rect 422186 315418 422422 315654
rect 422186 315098 422422 315334
rect 432986 704602 433222 704838
rect 432986 704282 433222 704518
rect 432986 686218 433222 686454
rect 432986 685898 433222 686134
rect 436586 689818 436822 690054
rect 436586 689498 436822 689734
rect 440186 693418 440422 693654
rect 440186 693098 440422 693334
rect 440186 657418 440422 657654
rect 440186 657098 440422 657334
rect 461786 711182 462022 711418
rect 461786 710862 462022 711098
rect 458186 709302 458422 709538
rect 458186 708982 458422 709218
rect 454586 707422 454822 707658
rect 454586 707102 454822 707338
rect 443786 697018 444022 697254
rect 443786 696698 444022 696934
rect 443786 661018 444022 661254
rect 443786 660698 444022 660934
rect 450986 705542 451222 705778
rect 450986 705222 451222 705458
rect 450986 668218 451222 668454
rect 450986 667898 451222 668134
rect 454586 671818 454822 672054
rect 454586 671498 454822 671734
rect 458186 675418 458422 675654
rect 458186 675098 458422 675334
rect 479786 710242 480022 710478
rect 479786 709922 480022 710158
rect 476186 708362 476422 708598
rect 476186 708042 476422 708278
rect 472586 706482 472822 706718
rect 472586 706162 472822 706398
rect 461786 679018 462022 679254
rect 461786 678698 462022 678934
rect 468986 704602 469222 704838
rect 468986 704282 469222 704518
rect 468986 686218 469222 686454
rect 468986 685898 469222 686134
rect 472586 689818 472822 690054
rect 472586 689498 472822 689734
rect 476186 693418 476422 693654
rect 476186 693098 476422 693334
rect 476186 657418 476422 657654
rect 476186 657098 476422 657334
rect 497786 711182 498022 711418
rect 497786 710862 498022 711098
rect 494186 709302 494422 709538
rect 494186 708982 494422 709218
rect 490586 707422 490822 707658
rect 490586 707102 490822 707338
rect 479786 697018 480022 697254
rect 479786 696698 480022 696934
rect 479786 661018 480022 661254
rect 479786 660698 480022 660934
rect 486986 705542 487222 705778
rect 486986 705222 487222 705458
rect 486986 668218 487222 668454
rect 486986 667898 487222 668134
rect 490586 671818 490822 672054
rect 490586 671498 490822 671734
rect 494186 675418 494422 675654
rect 494186 675098 494422 675334
rect 515786 710242 516022 710478
rect 515786 709922 516022 710158
rect 512186 708362 512422 708598
rect 512186 708042 512422 708278
rect 508586 706482 508822 706718
rect 508586 706162 508822 706398
rect 497786 679018 498022 679254
rect 497786 678698 498022 678934
rect 504986 704602 505222 704838
rect 504986 704282 505222 704518
rect 504986 686218 505222 686454
rect 504986 685898 505222 686134
rect 508586 689818 508822 690054
rect 508586 689498 508822 689734
rect 512186 693418 512422 693654
rect 512186 693098 512422 693334
rect 512186 657418 512422 657654
rect 512186 657098 512422 657334
rect 533786 711182 534022 711418
rect 533786 710862 534022 711098
rect 530186 709302 530422 709538
rect 530186 708982 530422 709218
rect 526586 707422 526822 707658
rect 526586 707102 526822 707338
rect 515786 697018 516022 697254
rect 515786 696698 516022 696934
rect 515786 661018 516022 661254
rect 515786 660698 516022 660934
rect 522986 705542 523222 705778
rect 522986 705222 523222 705458
rect 522986 668218 523222 668454
rect 522986 667898 523222 668134
rect 432986 650218 433222 650454
rect 432986 649898 433222 650134
rect 516982 643018 517218 643254
rect 516982 642698 517218 642934
rect 516982 639418 517218 639654
rect 516982 639098 517218 639334
rect 516982 635818 517218 636054
rect 516982 635498 517218 635734
rect 516982 632218 517218 632454
rect 516982 631898 517218 632134
rect 522986 632218 523222 632454
rect 522986 631898 523222 632134
rect 516536 625018 516772 625254
rect 516536 624698 516772 624934
rect 516536 621418 516772 621654
rect 516536 621098 516772 621334
rect 516536 617818 516772 618054
rect 516536 617498 516772 617734
rect 432986 614218 433222 614454
rect 432986 613898 433222 614134
rect 516536 614218 516772 614454
rect 516536 613898 516772 614134
rect 516982 607018 517218 607254
rect 516982 606698 517218 606934
rect 516982 603418 517218 603654
rect 516982 603098 517218 603334
rect 516982 599818 517218 600054
rect 516982 599498 517218 599734
rect 516982 596218 517218 596454
rect 516982 595898 517218 596134
rect 522986 596218 523222 596454
rect 522986 595898 523222 596134
rect 516536 589018 516772 589254
rect 516536 588698 516772 588934
rect 516536 585418 516772 585654
rect 516536 585098 516772 585334
rect 516536 581818 516772 582054
rect 516536 581498 516772 581734
rect 518854 579582 519090 579818
rect 437342 579052 437578 579138
rect 437342 578988 437428 579052
rect 437428 578988 437492 579052
rect 437492 578988 437578 579052
rect 437342 578902 437578 578988
rect 432986 578218 433222 578454
rect 432986 577898 433222 578134
rect 516536 578218 516772 578454
rect 516536 577898 516772 578134
rect 516982 571018 517218 571254
rect 516982 570698 517218 570934
rect 516982 567418 517218 567654
rect 516982 567098 517218 567334
rect 516982 563818 517218 564054
rect 516982 563498 517218 563734
rect 522986 560218 523222 560454
rect 522986 559898 523222 560134
rect 432986 542218 433222 542454
rect 432986 541898 433222 542134
rect 432986 506218 433222 506454
rect 432986 505898 433222 506134
rect 432986 470218 433222 470454
rect 432986 469898 433222 470134
rect 432986 434218 433222 434454
rect 432986 433898 433222 434134
rect 432986 398218 433222 398454
rect 432986 397898 433222 398134
rect 432986 362218 433222 362454
rect 432986 361898 433222 362134
rect 427774 346492 428010 346578
rect 427774 346428 427860 346492
rect 427860 346428 427924 346492
rect 427924 346428 428010 346492
rect 427774 346342 428010 346428
rect 427774 341124 427860 341138
rect 427860 341124 427924 341138
rect 427924 341124 428010 341138
rect 427774 340902 428010 341124
rect 425786 319018 426022 319254
rect 425786 318698 426022 318934
rect 432986 326218 433222 326454
rect 432986 325898 433222 326134
rect 436586 545818 436822 546054
rect 436586 545498 436822 545734
rect 436586 509818 436822 510054
rect 436586 509498 436822 509734
rect 436586 473818 436822 474054
rect 436586 473498 436822 473734
rect 436586 437818 436822 438054
rect 436586 437498 436822 437734
rect 436586 401818 436822 402054
rect 436586 401498 436822 401734
rect 436586 365818 436822 366054
rect 436586 365498 436822 365734
rect 440186 549418 440422 549654
rect 440186 549098 440422 549334
rect 440186 513418 440422 513654
rect 440186 513098 440422 513334
rect 440186 477418 440422 477654
rect 440186 477098 440422 477334
rect 440186 441418 440422 441654
rect 440186 441098 440422 441334
rect 440186 405418 440422 405654
rect 440186 405098 440422 405334
rect 440186 369418 440422 369654
rect 440186 369098 440422 369334
rect 437894 345812 438130 345898
rect 437894 345748 437980 345812
rect 437980 345748 438044 345812
rect 438044 345748 438130 345812
rect 437894 345662 438130 345748
rect 437710 344982 437946 345218
rect 437526 343092 437762 343178
rect 437526 343028 437612 343092
rect 437612 343028 437676 343092
rect 437676 343028 437762 343092
rect 437526 342942 437762 343028
rect 439366 339542 439602 339778
rect 436586 329818 436822 330054
rect 436586 329498 436822 329734
rect 440186 333418 440422 333654
rect 440186 333098 440422 333334
rect 443786 553018 444022 553254
rect 443786 552698 444022 552934
rect 443786 517018 444022 517254
rect 443786 516698 444022 516934
rect 443786 481018 444022 481254
rect 443786 480698 444022 480934
rect 443786 445018 444022 445254
rect 443786 444698 444022 444934
rect 450986 524218 451222 524454
rect 450986 523898 451222 524134
rect 450986 488218 451222 488454
rect 450986 487898 451222 488134
rect 450986 452218 451222 452454
rect 450986 451898 451222 452134
rect 450986 416218 451222 416454
rect 450986 415898 451222 416134
rect 454586 527818 454822 528054
rect 454586 527498 454822 527734
rect 454586 491818 454822 492054
rect 454586 491498 454822 491734
rect 454586 455818 454822 456054
rect 454586 455498 454822 455734
rect 454586 419818 454822 420054
rect 454586 419498 454822 419734
rect 458186 531418 458422 531654
rect 458186 531098 458422 531334
rect 458186 495418 458422 495654
rect 458186 495098 458422 495334
rect 458186 459418 458422 459654
rect 458186 459098 458422 459334
rect 458186 423418 458422 423654
rect 458186 423098 458422 423334
rect 461786 535018 462022 535254
rect 461786 534698 462022 534934
rect 461786 499018 462022 499254
rect 461786 498698 462022 498934
rect 461786 463018 462022 463254
rect 461786 462698 462022 462934
rect 461786 427018 462022 427254
rect 461786 426698 462022 426934
rect 468986 542218 469222 542454
rect 468986 541898 469222 542134
rect 468986 506218 469222 506454
rect 468986 505898 469222 506134
rect 468986 470218 469222 470454
rect 468986 469898 469222 470134
rect 468986 434218 469222 434454
rect 468986 433898 469222 434134
rect 472586 545818 472822 546054
rect 472586 545498 472822 545734
rect 472586 509818 472822 510054
rect 472586 509498 472822 509734
rect 472586 473818 472822 474054
rect 472586 473498 472822 473734
rect 472586 437818 472822 438054
rect 472586 437498 472822 437734
rect 476186 549418 476422 549654
rect 476186 549098 476422 549334
rect 476186 513418 476422 513654
rect 476186 513098 476422 513334
rect 476186 477418 476422 477654
rect 476186 477098 476422 477334
rect 476186 441418 476422 441654
rect 476186 441098 476422 441334
rect 479786 553018 480022 553254
rect 479786 552698 480022 552934
rect 479786 517018 480022 517254
rect 479786 516698 480022 516934
rect 479786 481018 480022 481254
rect 479786 480698 480022 480934
rect 479786 445018 480022 445254
rect 479786 444698 480022 444934
rect 486986 524218 487222 524454
rect 486986 523898 487222 524134
rect 486986 488218 487222 488454
rect 486986 487898 487222 488134
rect 486986 452218 487222 452454
rect 486986 451898 487222 452134
rect 486986 416218 487222 416454
rect 486986 415898 487222 416134
rect 490586 527818 490822 528054
rect 490586 527498 490822 527734
rect 490586 491818 490822 492054
rect 490586 491498 490822 491734
rect 490586 455818 490822 456054
rect 490586 455498 490822 455734
rect 490586 419818 490822 420054
rect 490586 419498 490822 419734
rect 494186 531418 494422 531654
rect 494186 531098 494422 531334
rect 494186 495418 494422 495654
rect 494186 495098 494422 495334
rect 494186 459418 494422 459654
rect 494186 459098 494422 459334
rect 494186 423418 494422 423654
rect 494186 423098 494422 423334
rect 497786 535018 498022 535254
rect 497786 534698 498022 534934
rect 497786 499018 498022 499254
rect 497786 498698 498022 498934
rect 497786 463018 498022 463254
rect 497786 462698 498022 462934
rect 497786 427018 498022 427254
rect 497786 426698 498022 426934
rect 504986 542218 505222 542454
rect 504986 541898 505222 542134
rect 504986 506218 505222 506454
rect 504986 505898 505222 506134
rect 504986 470218 505222 470454
rect 504986 469898 505222 470134
rect 504986 434218 505222 434454
rect 504986 433898 505222 434134
rect 508586 545818 508822 546054
rect 508586 545498 508822 545734
rect 508586 509818 508822 510054
rect 508586 509498 508822 509734
rect 508586 473818 508822 474054
rect 508586 473498 508822 473734
rect 508586 437818 508822 438054
rect 508586 437498 508822 437734
rect 512186 549418 512422 549654
rect 512186 549098 512422 549334
rect 512186 513418 512422 513654
rect 512186 513098 512422 513334
rect 512186 477418 512422 477654
rect 512186 477098 512422 477334
rect 512186 441418 512422 441654
rect 512186 441098 512422 441334
rect 515786 553018 516022 553254
rect 515786 552698 516022 552934
rect 515786 517018 516022 517254
rect 515786 516698 516022 516934
rect 515786 481018 516022 481254
rect 515786 480698 516022 480934
rect 515786 445018 516022 445254
rect 515786 444698 516022 444934
rect 522986 524218 523222 524454
rect 522986 523898 523222 524134
rect 522986 488218 523222 488454
rect 522986 487898 523222 488134
rect 522986 452218 523222 452454
rect 522986 451898 523222 452134
rect 522986 416218 523222 416454
rect 522986 415898 523222 416134
rect 526586 671818 526822 672054
rect 526586 671498 526822 671734
rect 526586 635818 526822 636054
rect 526586 635498 526822 635734
rect 526586 599818 526822 600054
rect 526586 599498 526822 599734
rect 526586 563818 526822 564054
rect 526586 563498 526822 563734
rect 526586 527818 526822 528054
rect 526586 527498 526822 527734
rect 526586 491818 526822 492054
rect 526586 491498 526822 491734
rect 526586 455818 526822 456054
rect 526586 455498 526822 455734
rect 526586 419818 526822 420054
rect 526586 419498 526822 419734
rect 530186 675418 530422 675654
rect 530186 675098 530422 675334
rect 530186 639418 530422 639654
rect 530186 639098 530422 639334
rect 530186 603418 530422 603654
rect 530186 603098 530422 603334
rect 530186 567418 530422 567654
rect 530186 567098 530422 567334
rect 530186 531418 530422 531654
rect 530186 531098 530422 531334
rect 530186 495418 530422 495654
rect 530186 495098 530422 495334
rect 530186 459418 530422 459654
rect 530186 459098 530422 459334
rect 530186 423418 530422 423654
rect 530186 423098 530422 423334
rect 551786 710242 552022 710478
rect 551786 709922 552022 710158
rect 548186 708362 548422 708598
rect 548186 708042 548422 708278
rect 544586 706482 544822 706718
rect 544586 706162 544822 706398
rect 533786 679018 534022 679254
rect 533786 678698 534022 678934
rect 533786 643018 534022 643254
rect 533786 642698 534022 642934
rect 533786 607018 534022 607254
rect 533786 606698 534022 606934
rect 533786 571018 534022 571254
rect 533786 570698 534022 570934
rect 533786 535018 534022 535254
rect 533786 534698 534022 534934
rect 533786 499018 534022 499254
rect 533786 498698 534022 498934
rect 533786 463018 534022 463254
rect 533786 462698 534022 462934
rect 533786 427018 534022 427254
rect 533786 426698 534022 426934
rect 443786 409018 444022 409254
rect 443786 408698 444022 408934
rect 526536 405418 526772 405654
rect 526536 405098 526772 405334
rect 526536 401818 526772 402054
rect 526536 401498 526772 401734
rect 526536 398218 526772 398454
rect 526536 397898 526772 398134
rect 526982 391018 527218 391254
rect 526982 390698 527218 390934
rect 533786 391018 534022 391254
rect 533786 390698 534022 390934
rect 526982 387418 527218 387654
rect 526982 387098 527218 387334
rect 526982 383818 527218 384054
rect 526982 383498 527218 383734
rect 526982 380218 527218 380454
rect 526982 379898 527218 380134
rect 443786 373018 444022 373254
rect 443786 372698 444022 372934
rect 526536 373018 526772 373254
rect 526536 372698 526772 372934
rect 526536 369418 526772 369654
rect 526536 369098 526772 369334
rect 526536 365818 526772 366054
rect 526536 365498 526772 365734
rect 526536 362218 526772 362454
rect 526536 361898 526772 362134
rect 526982 355018 527218 355254
rect 526982 354698 527218 354934
rect 533786 355018 534022 355254
rect 533786 354698 534022 354934
rect 526982 351418 527218 351654
rect 526982 351098 527218 351334
rect 527502 349212 527738 349298
rect 527502 349148 527588 349212
rect 527588 349148 527652 349212
rect 527652 349148 527738 349212
rect 527502 349062 527738 349148
rect 526982 347818 527218 348054
rect 526982 347498 527218 347734
rect 446726 346492 446962 346578
rect 446726 346428 446812 346492
rect 446812 346428 446876 346492
rect 446876 346428 446962 346492
rect 446726 346342 446962 346428
rect 447646 346492 447882 346578
rect 447646 346428 447732 346492
rect 447732 346428 447796 346492
rect 447796 346428 447882 346492
rect 447646 346342 447882 346428
rect 527870 346342 528106 346578
rect 447094 345812 447330 345898
rect 447094 345748 447180 345812
rect 447180 345748 447244 345812
rect 447244 345748 447330 345812
rect 447094 345662 447330 345748
rect 527502 345662 527738 345898
rect 527502 344982 527738 345218
rect 526982 344218 527218 344454
rect 526982 343898 527218 344134
rect 448014 343092 448250 343178
rect 448014 343028 448100 343092
rect 448100 343028 448164 343092
rect 448164 343028 448250 343092
rect 448014 342942 448250 343028
rect 449486 343092 449722 343178
rect 449486 343028 449572 343092
rect 449572 343028 449636 343092
rect 449636 343028 449722 343092
rect 449486 342942 449722 343028
rect 445438 342262 445674 342498
rect 444334 341582 444570 341818
rect 445070 341582 445306 341818
rect 444334 340372 444570 340458
rect 444334 340308 444420 340372
rect 444420 340308 444484 340372
rect 444484 340308 444570 340372
rect 444334 340222 444570 340308
rect 527502 342942 527738 343178
rect 527502 341732 527738 341818
rect 527502 341668 527588 341732
rect 527588 341668 527652 341732
rect 527652 341668 527738 341732
rect 527502 341582 527738 341668
rect 527870 340222 528106 340458
rect 450590 338182 450826 338418
rect 443786 337018 444022 337254
rect 443786 336698 444022 336934
rect 526536 337018 526772 337254
rect 526536 336698 526772 336934
rect 526536 333418 526772 333654
rect 526536 333098 526772 333334
rect 526536 329818 526772 330054
rect 526536 329498 526772 329734
rect 526536 326218 526772 326454
rect 526536 325898 526772 326134
rect 533786 319018 534022 319254
rect 533786 318698 534022 318934
rect 450986 308218 451222 308454
rect 450986 307898 451222 308134
rect 454586 311818 454822 312054
rect 454586 311498 454822 311734
rect 458186 315418 458422 315654
rect 458186 315098 458422 315334
rect 486986 308218 487222 308454
rect 486986 307898 487222 308134
rect 490586 311818 490822 312054
rect 490586 311498 490822 311734
rect 494186 315418 494422 315654
rect 494186 315098 494422 315334
rect 522986 308218 523222 308454
rect 522986 307898 523222 308134
rect 526586 311818 526822 312054
rect 526586 311498 526822 311734
rect 530186 315418 530422 315654
rect 530186 315098 530422 315334
rect 299786 301018 300022 301254
rect 299786 300698 300022 300934
rect 314250 293818 314486 294054
rect 314250 293498 314486 293734
rect 314250 290218 314486 290454
rect 314250 289898 314486 290134
rect 329610 283018 329846 283254
rect 329610 282698 329846 282934
rect 533786 283018 534022 283254
rect 533786 282698 534022 282934
rect 329610 279418 329846 279654
rect 329610 279098 329846 279334
rect 329610 275818 329846 276054
rect 329610 275498 329846 275734
rect 329610 272218 329846 272454
rect 329610 271898 329846 272134
rect 299786 265018 300022 265254
rect 299786 264698 300022 264934
rect 314250 265018 314486 265254
rect 314250 264698 314486 264934
rect 314250 261418 314486 261654
rect 314250 261098 314486 261334
rect 314250 257818 314486 258054
rect 314250 257498 314486 257734
rect 314250 254218 314486 254454
rect 314250 253898 314486 254134
rect 329610 247018 329846 247254
rect 329610 246698 329846 246934
rect 533786 247018 534022 247254
rect 533786 246698 534022 246934
rect 329610 243418 329846 243654
rect 329610 243098 329846 243334
rect 329610 239818 329846 240054
rect 329610 239498 329846 239734
rect 329610 236218 329846 236454
rect 329610 235898 329846 236134
rect 299786 229018 300022 229254
rect 299786 228698 300022 228934
rect 314250 229018 314486 229254
rect 314250 228698 314486 228934
rect 314250 225418 314486 225654
rect 314250 225098 314486 225334
rect 314250 221818 314486 222054
rect 314250 221498 314486 221734
rect 314250 218218 314486 218454
rect 314250 217898 314486 218134
rect 329610 211018 329846 211254
rect 329610 210698 329846 210934
rect 533786 211018 534022 211254
rect 533786 210698 534022 210934
rect 329610 207418 329846 207654
rect 329610 207098 329846 207334
rect 329610 203818 329846 204054
rect 329610 203498 329846 203734
rect 329610 200218 329846 200454
rect 329610 199898 329846 200134
rect 299786 193018 300022 193254
rect 299786 192698 300022 192934
rect 314250 193018 314486 193254
rect 314250 192698 314486 192934
rect 314250 189418 314486 189654
rect 314250 189098 314486 189334
rect 314250 185818 314486 186054
rect 314250 185498 314486 185734
rect 314250 182218 314486 182454
rect 314250 181898 314486 182134
rect 329610 175018 329846 175254
rect 329610 174698 329846 174934
rect 533786 175018 534022 175254
rect 533786 174698 534022 174934
rect 329610 171418 329846 171654
rect 329610 171098 329846 171334
rect 329610 167818 329846 168054
rect 329610 167498 329846 167734
rect 329610 164218 329846 164454
rect 329610 163898 329846 164134
rect 299786 157018 300022 157254
rect 299786 156698 300022 156934
rect 314250 157018 314486 157254
rect 314250 156698 314486 156934
rect 314250 153418 314486 153654
rect 314250 153098 314486 153334
rect 314250 149818 314486 150054
rect 314250 149498 314486 149734
rect 314250 146218 314486 146454
rect 314250 145898 314486 146134
rect 329610 139018 329846 139254
rect 329610 138698 329846 138934
rect 533786 139018 534022 139254
rect 533786 138698 534022 138934
rect 329610 135418 329846 135654
rect 329610 135098 329846 135334
rect 329610 131818 329846 132054
rect 329610 131498 329846 131734
rect 329610 128218 329846 128454
rect 329610 127898 329846 128134
rect 299786 121018 300022 121254
rect 299786 120698 300022 120934
rect 314250 121018 314486 121254
rect 314250 120698 314486 120934
rect 314250 117418 314486 117654
rect 314250 117098 314486 117334
rect 314250 113818 314486 114054
rect 314250 113498 314486 113734
rect 314250 110218 314486 110454
rect 314250 109898 314486 110134
rect 329610 103018 329846 103254
rect 329610 102698 329846 102934
rect 533786 103018 534022 103254
rect 533786 102698 534022 102934
rect 329610 99418 329846 99654
rect 329610 99098 329846 99334
rect 329610 95818 329846 96054
rect 329610 95498 329846 95734
rect 329610 92218 329846 92454
rect 329610 91898 329846 92134
rect 299786 85018 300022 85254
rect 299786 84698 300022 84934
rect 314250 85018 314486 85254
rect 314250 84698 314486 84934
rect 299786 49018 300022 49254
rect 299786 48698 300022 48934
rect 299786 13018 300022 13254
rect 299786 12698 300022 12934
rect 281786 -7162 282022 -6926
rect 281786 -7482 282022 -7246
rect 306986 56218 307222 56454
rect 306986 55898 307222 56134
rect 306986 20218 307222 20454
rect 306986 19898 307222 20134
rect 306986 -1522 307222 -1286
rect 306986 -1842 307222 -1606
rect 310586 59818 310822 60054
rect 310586 59498 310822 59734
rect 310586 23818 310822 24054
rect 310586 23498 310822 23734
rect 310586 -3402 310822 -3166
rect 310586 -3722 310822 -3486
rect 314186 63418 314422 63654
rect 314186 63098 314422 63334
rect 314186 27418 314422 27654
rect 314186 27098 314422 27334
rect 314186 -5282 314422 -5046
rect 314186 -5602 314422 -5366
rect 317786 67018 318022 67254
rect 317786 66698 318022 66934
rect 317786 31018 318022 31254
rect 317786 30698 318022 30934
rect 299786 -6222 300022 -5986
rect 299786 -6542 300022 -6306
rect 324986 74218 325222 74454
rect 324986 73898 325222 74134
rect 324986 38218 325222 38454
rect 324986 37898 325222 38134
rect 324986 2218 325222 2454
rect 324986 1898 325222 2134
rect 324986 -582 325222 -346
rect 324986 -902 325222 -666
rect 328586 41818 328822 42054
rect 328586 41498 328822 41734
rect 328586 5818 328822 6054
rect 328586 5498 328822 5734
rect 328586 -2462 328822 -2226
rect 328586 -2782 328822 -2546
rect 332186 45418 332422 45654
rect 332186 45098 332422 45334
rect 332186 9418 332422 9654
rect 332186 9098 332422 9334
rect 332186 -4342 332422 -4106
rect 332186 -4662 332422 -4426
rect 335786 49018 336022 49254
rect 335786 48698 336022 48934
rect 335786 13018 336022 13254
rect 335786 12698 336022 12934
rect 317786 -7162 318022 -6926
rect 317786 -7482 318022 -7246
rect 342986 56218 343222 56454
rect 342986 55898 343222 56134
rect 342986 20218 343222 20454
rect 342986 19898 343222 20134
rect 342986 -1522 343222 -1286
rect 342986 -1842 343222 -1606
rect 346586 59818 346822 60054
rect 346586 59498 346822 59734
rect 346586 23818 346822 24054
rect 346586 23498 346822 23734
rect 346586 -3402 346822 -3166
rect 346586 -3722 346822 -3486
rect 350186 63418 350422 63654
rect 350186 63098 350422 63334
rect 350186 27418 350422 27654
rect 350186 27098 350422 27334
rect 350186 -5282 350422 -5046
rect 350186 -5602 350422 -5366
rect 353786 67018 354022 67254
rect 353786 66698 354022 66934
rect 353786 31018 354022 31254
rect 353786 30698 354022 30934
rect 335786 -6222 336022 -5986
rect 335786 -6542 336022 -6306
rect 360986 74218 361222 74454
rect 360986 73898 361222 74134
rect 360986 38218 361222 38454
rect 360986 37898 361222 38134
rect 360986 2218 361222 2454
rect 360986 1898 361222 2134
rect 360986 -582 361222 -346
rect 360986 -902 361222 -666
rect 364586 41818 364822 42054
rect 364586 41498 364822 41734
rect 364586 5818 364822 6054
rect 364586 5498 364822 5734
rect 364586 -2462 364822 -2226
rect 364586 -2782 364822 -2546
rect 368186 45418 368422 45654
rect 368186 45098 368422 45334
rect 368186 9418 368422 9654
rect 368186 9098 368422 9334
rect 368186 -4342 368422 -4106
rect 368186 -4662 368422 -4426
rect 371786 49018 372022 49254
rect 371786 48698 372022 48934
rect 371786 13018 372022 13254
rect 371786 12698 372022 12934
rect 353786 -7162 354022 -6926
rect 353786 -7482 354022 -7246
rect 378986 56218 379222 56454
rect 378986 55898 379222 56134
rect 378986 20218 379222 20454
rect 378986 19898 379222 20134
rect 378986 -1522 379222 -1286
rect 378986 -1842 379222 -1606
rect 382586 59818 382822 60054
rect 382586 59498 382822 59734
rect 382586 23818 382822 24054
rect 382586 23498 382822 23734
rect 382586 -3402 382822 -3166
rect 382586 -3722 382822 -3486
rect 386186 63418 386422 63654
rect 386186 63098 386422 63334
rect 386186 27418 386422 27654
rect 386186 27098 386422 27334
rect 386186 -5282 386422 -5046
rect 386186 -5602 386422 -5366
rect 389786 67018 390022 67254
rect 389786 66698 390022 66934
rect 389786 31018 390022 31254
rect 389786 30698 390022 30934
rect 371786 -6222 372022 -5986
rect 371786 -6542 372022 -6306
rect 396986 74218 397222 74454
rect 396986 73898 397222 74134
rect 396986 38218 397222 38454
rect 396986 37898 397222 38134
rect 396986 2218 397222 2454
rect 396986 1898 397222 2134
rect 396986 -582 397222 -346
rect 396986 -902 397222 -666
rect 400586 41818 400822 42054
rect 400586 41498 400822 41734
rect 400586 5818 400822 6054
rect 400586 5498 400822 5734
rect 400586 -2462 400822 -2226
rect 400586 -2782 400822 -2546
rect 404186 45418 404422 45654
rect 404186 45098 404422 45334
rect 404186 9418 404422 9654
rect 404186 9098 404422 9334
rect 404186 -4342 404422 -4106
rect 404186 -4662 404422 -4426
rect 407786 49018 408022 49254
rect 407786 48698 408022 48934
rect 407786 13018 408022 13254
rect 407786 12698 408022 12934
rect 389786 -7162 390022 -6926
rect 389786 -7482 390022 -7246
rect 414986 56218 415222 56454
rect 414986 55898 415222 56134
rect 414986 20218 415222 20454
rect 414986 19898 415222 20134
rect 414986 -1522 415222 -1286
rect 414986 -1842 415222 -1606
rect 418586 59818 418822 60054
rect 418586 59498 418822 59734
rect 418586 23818 418822 24054
rect 418586 23498 418822 23734
rect 418586 -3402 418822 -3166
rect 418586 -3722 418822 -3486
rect 422186 63418 422422 63654
rect 422186 63098 422422 63334
rect 422186 27418 422422 27654
rect 422186 27098 422422 27334
rect 422186 -5282 422422 -5046
rect 422186 -5602 422422 -5366
rect 425786 67018 426022 67254
rect 425786 66698 426022 66934
rect 425786 31018 426022 31254
rect 425786 30698 426022 30934
rect 407786 -6222 408022 -5986
rect 407786 -6542 408022 -6306
rect 432986 74218 433222 74454
rect 432986 73898 433222 74134
rect 432986 38218 433222 38454
rect 432986 37898 433222 38134
rect 432986 2218 433222 2454
rect 432986 1898 433222 2134
rect 432986 -582 433222 -346
rect 432986 -902 433222 -666
rect 436586 41818 436822 42054
rect 436586 41498 436822 41734
rect 436586 5818 436822 6054
rect 436586 5498 436822 5734
rect 436586 -2462 436822 -2226
rect 436586 -2782 436822 -2546
rect 440186 45418 440422 45654
rect 440186 45098 440422 45334
rect 440186 9418 440422 9654
rect 440186 9098 440422 9334
rect 440186 -4342 440422 -4106
rect 440186 -4662 440422 -4426
rect 443786 49018 444022 49254
rect 443786 48698 444022 48934
rect 443786 13018 444022 13254
rect 443786 12698 444022 12934
rect 425786 -7162 426022 -6926
rect 425786 -7482 426022 -7246
rect 450986 56218 451222 56454
rect 450986 55898 451222 56134
rect 450986 20218 451222 20454
rect 450986 19898 451222 20134
rect 450986 -1522 451222 -1286
rect 450986 -1842 451222 -1606
rect 454586 59818 454822 60054
rect 454586 59498 454822 59734
rect 454586 23818 454822 24054
rect 454586 23498 454822 23734
rect 454586 -3402 454822 -3166
rect 454586 -3722 454822 -3486
rect 458186 63418 458422 63654
rect 458186 63098 458422 63334
rect 458186 27418 458422 27654
rect 458186 27098 458422 27334
rect 458186 -5282 458422 -5046
rect 458186 -5602 458422 -5366
rect 461786 67018 462022 67254
rect 461786 66698 462022 66934
rect 461786 31018 462022 31254
rect 461786 30698 462022 30934
rect 443786 -6222 444022 -5986
rect 443786 -6542 444022 -6306
rect 468986 74218 469222 74454
rect 468986 73898 469222 74134
rect 468986 38218 469222 38454
rect 468986 37898 469222 38134
rect 468986 2218 469222 2454
rect 468986 1898 469222 2134
rect 468986 -582 469222 -346
rect 468986 -902 469222 -666
rect 472586 41818 472822 42054
rect 472586 41498 472822 41734
rect 472586 5818 472822 6054
rect 472586 5498 472822 5734
rect 472586 -2462 472822 -2226
rect 472586 -2782 472822 -2546
rect 476186 45418 476422 45654
rect 476186 45098 476422 45334
rect 476186 9418 476422 9654
rect 476186 9098 476422 9334
rect 476186 -4342 476422 -4106
rect 476186 -4662 476422 -4426
rect 479786 49018 480022 49254
rect 479786 48698 480022 48934
rect 479786 13018 480022 13254
rect 479786 12698 480022 12934
rect 461786 -7162 462022 -6926
rect 461786 -7482 462022 -7246
rect 486986 56218 487222 56454
rect 486986 55898 487222 56134
rect 486986 20218 487222 20454
rect 486986 19898 487222 20134
rect 486986 -1522 487222 -1286
rect 486986 -1842 487222 -1606
rect 490586 59818 490822 60054
rect 490586 59498 490822 59734
rect 490586 23818 490822 24054
rect 490586 23498 490822 23734
rect 490586 -3402 490822 -3166
rect 490586 -3722 490822 -3486
rect 494186 63418 494422 63654
rect 494186 63098 494422 63334
rect 494186 27418 494422 27654
rect 494186 27098 494422 27334
rect 494186 -5282 494422 -5046
rect 494186 -5602 494422 -5366
rect 497786 67018 498022 67254
rect 497786 66698 498022 66934
rect 497786 31018 498022 31254
rect 497786 30698 498022 30934
rect 479786 -6222 480022 -5986
rect 479786 -6542 480022 -6306
rect 504986 74218 505222 74454
rect 504986 73898 505222 74134
rect 504986 38218 505222 38454
rect 504986 37898 505222 38134
rect 504986 2218 505222 2454
rect 504986 1898 505222 2134
rect 504986 -582 505222 -346
rect 504986 -902 505222 -666
rect 508586 41818 508822 42054
rect 508586 41498 508822 41734
rect 508586 5818 508822 6054
rect 508586 5498 508822 5734
rect 508586 -2462 508822 -2226
rect 508586 -2782 508822 -2546
rect 512186 45418 512422 45654
rect 512186 45098 512422 45334
rect 512186 9418 512422 9654
rect 512186 9098 512422 9334
rect 512186 -4342 512422 -4106
rect 512186 -4662 512422 -4426
rect 515786 49018 516022 49254
rect 515786 48698 516022 48934
rect 515786 13018 516022 13254
rect 515786 12698 516022 12934
rect 497786 -7162 498022 -6926
rect 497786 -7482 498022 -7246
rect 522986 56218 523222 56454
rect 522986 55898 523222 56134
rect 522986 20218 523222 20454
rect 522986 19898 523222 20134
rect 522986 -1522 523222 -1286
rect 522986 -1842 523222 -1606
rect 526586 59818 526822 60054
rect 526586 59498 526822 59734
rect 526586 23818 526822 24054
rect 526586 23498 526822 23734
rect 526586 -3402 526822 -3166
rect 526586 -3722 526822 -3486
rect 530186 63418 530422 63654
rect 530186 63098 530422 63334
rect 530186 27418 530422 27654
rect 530186 27098 530422 27334
rect 530186 -5282 530422 -5046
rect 530186 -5602 530422 -5366
rect 533786 67018 534022 67254
rect 533786 66698 534022 66934
rect 533786 31018 534022 31254
rect 533786 30698 534022 30934
rect 515786 -6222 516022 -5986
rect 515786 -6542 516022 -6306
rect 540986 704602 541222 704838
rect 540986 704282 541222 704518
rect 540986 686218 541222 686454
rect 540986 685898 541222 686134
rect 540986 650218 541222 650454
rect 540986 649898 541222 650134
rect 540986 614218 541222 614454
rect 540986 613898 541222 614134
rect 540986 578218 541222 578454
rect 540986 577898 541222 578134
rect 540986 542218 541222 542454
rect 540986 541898 541222 542134
rect 540986 506218 541222 506454
rect 540986 505898 541222 506134
rect 540986 470218 541222 470454
rect 540986 469898 541222 470134
rect 540986 434218 541222 434454
rect 540986 433898 541222 434134
rect 540986 398218 541222 398454
rect 540986 397898 541222 398134
rect 540986 362218 541222 362454
rect 540986 361898 541222 362134
rect 540986 326218 541222 326454
rect 540986 325898 541222 326134
rect 540986 290218 541222 290454
rect 540986 289898 541222 290134
rect 540986 254218 541222 254454
rect 540986 253898 541222 254134
rect 540986 218218 541222 218454
rect 540986 217898 541222 218134
rect 540986 182218 541222 182454
rect 540986 181898 541222 182134
rect 540986 146218 541222 146454
rect 540986 145898 541222 146134
rect 540986 110218 541222 110454
rect 540986 109898 541222 110134
rect 540986 74218 541222 74454
rect 540986 73898 541222 74134
rect 540986 38218 541222 38454
rect 540986 37898 541222 38134
rect 540986 2218 541222 2454
rect 540986 1898 541222 2134
rect 540986 -582 541222 -346
rect 540986 -902 541222 -666
rect 544586 689818 544822 690054
rect 544586 689498 544822 689734
rect 544586 653818 544822 654054
rect 544586 653498 544822 653734
rect 544586 617818 544822 618054
rect 544586 617498 544822 617734
rect 544586 581818 544822 582054
rect 544586 581498 544822 581734
rect 544586 545818 544822 546054
rect 544586 545498 544822 545734
rect 544586 509818 544822 510054
rect 544586 509498 544822 509734
rect 544586 473818 544822 474054
rect 544586 473498 544822 473734
rect 544586 437818 544822 438054
rect 544586 437498 544822 437734
rect 544586 401818 544822 402054
rect 544586 401498 544822 401734
rect 544586 365818 544822 366054
rect 544586 365498 544822 365734
rect 544586 329818 544822 330054
rect 544586 329498 544822 329734
rect 544586 293818 544822 294054
rect 544586 293498 544822 293734
rect 544586 257818 544822 258054
rect 544586 257498 544822 257734
rect 544586 221818 544822 222054
rect 544586 221498 544822 221734
rect 544586 185818 544822 186054
rect 544586 185498 544822 185734
rect 544586 149818 544822 150054
rect 544586 149498 544822 149734
rect 544586 113818 544822 114054
rect 544586 113498 544822 113734
rect 544586 77818 544822 78054
rect 544586 77498 544822 77734
rect 544586 41818 544822 42054
rect 544586 41498 544822 41734
rect 544586 5818 544822 6054
rect 544586 5498 544822 5734
rect 544586 -2462 544822 -2226
rect 544586 -2782 544822 -2546
rect 548186 693418 548422 693654
rect 548186 693098 548422 693334
rect 548186 657418 548422 657654
rect 548186 657098 548422 657334
rect 548186 621418 548422 621654
rect 548186 621098 548422 621334
rect 548186 585418 548422 585654
rect 548186 585098 548422 585334
rect 548186 549418 548422 549654
rect 548186 549098 548422 549334
rect 548186 513418 548422 513654
rect 548186 513098 548422 513334
rect 548186 477418 548422 477654
rect 548186 477098 548422 477334
rect 548186 441418 548422 441654
rect 548186 441098 548422 441334
rect 548186 405418 548422 405654
rect 548186 405098 548422 405334
rect 548186 369418 548422 369654
rect 548186 369098 548422 369334
rect 548186 333418 548422 333654
rect 548186 333098 548422 333334
rect 548186 297418 548422 297654
rect 548186 297098 548422 297334
rect 548186 261418 548422 261654
rect 548186 261098 548422 261334
rect 548186 225418 548422 225654
rect 548186 225098 548422 225334
rect 548186 189418 548422 189654
rect 548186 189098 548422 189334
rect 548186 153418 548422 153654
rect 548186 153098 548422 153334
rect 548186 117418 548422 117654
rect 548186 117098 548422 117334
rect 548186 81418 548422 81654
rect 548186 81098 548422 81334
rect 548186 45418 548422 45654
rect 548186 45098 548422 45334
rect 548186 9418 548422 9654
rect 548186 9098 548422 9334
rect 548186 -4342 548422 -4106
rect 548186 -4662 548422 -4426
rect 569786 711182 570022 711418
rect 569786 710862 570022 711098
rect 566186 709302 566422 709538
rect 566186 708982 566422 709218
rect 562586 707422 562822 707658
rect 562586 707102 562822 707338
rect 551786 697018 552022 697254
rect 551786 696698 552022 696934
rect 551786 661018 552022 661254
rect 551786 660698 552022 660934
rect 551786 625018 552022 625254
rect 551786 624698 552022 624934
rect 551786 589018 552022 589254
rect 551786 588698 552022 588934
rect 551786 553018 552022 553254
rect 551786 552698 552022 552934
rect 551786 517018 552022 517254
rect 551786 516698 552022 516934
rect 551786 481018 552022 481254
rect 551786 480698 552022 480934
rect 551786 445018 552022 445254
rect 551786 444698 552022 444934
rect 551786 409018 552022 409254
rect 551786 408698 552022 408934
rect 551786 373018 552022 373254
rect 551786 372698 552022 372934
rect 551786 337018 552022 337254
rect 551786 336698 552022 336934
rect 551786 301018 552022 301254
rect 551786 300698 552022 300934
rect 551786 265018 552022 265254
rect 551786 264698 552022 264934
rect 551786 229018 552022 229254
rect 551786 228698 552022 228934
rect 551786 193018 552022 193254
rect 551786 192698 552022 192934
rect 551786 157018 552022 157254
rect 551786 156698 552022 156934
rect 551786 121018 552022 121254
rect 551786 120698 552022 120934
rect 551786 85018 552022 85254
rect 551786 84698 552022 84934
rect 551786 49018 552022 49254
rect 551786 48698 552022 48934
rect 551786 13018 552022 13254
rect 551786 12698 552022 12934
rect 533786 -7162 534022 -6926
rect 533786 -7482 534022 -7246
rect 558986 705542 559222 705778
rect 558986 705222 559222 705458
rect 558986 668218 559222 668454
rect 558986 667898 559222 668134
rect 558986 632218 559222 632454
rect 558986 631898 559222 632134
rect 558986 596218 559222 596454
rect 558986 595898 559222 596134
rect 558986 560218 559222 560454
rect 558986 559898 559222 560134
rect 558986 524218 559222 524454
rect 558986 523898 559222 524134
rect 558986 488218 559222 488454
rect 558986 487898 559222 488134
rect 558986 452218 559222 452454
rect 558986 451898 559222 452134
rect 558986 416218 559222 416454
rect 558986 415898 559222 416134
rect 558986 380218 559222 380454
rect 558986 379898 559222 380134
rect 558986 344218 559222 344454
rect 558986 343898 559222 344134
rect 558986 308218 559222 308454
rect 558986 307898 559222 308134
rect 558986 272218 559222 272454
rect 558986 271898 559222 272134
rect 558986 236218 559222 236454
rect 558986 235898 559222 236134
rect 558986 200218 559222 200454
rect 558986 199898 559222 200134
rect 558986 164218 559222 164454
rect 558986 163898 559222 164134
rect 558986 128218 559222 128454
rect 558986 127898 559222 128134
rect 558986 92218 559222 92454
rect 558986 91898 559222 92134
rect 558986 56218 559222 56454
rect 558986 55898 559222 56134
rect 558986 20218 559222 20454
rect 558986 19898 559222 20134
rect 558986 -1522 559222 -1286
rect 558986 -1842 559222 -1606
rect 562586 671818 562822 672054
rect 562586 671498 562822 671734
rect 562586 635818 562822 636054
rect 562586 635498 562822 635734
rect 562586 599818 562822 600054
rect 562586 599498 562822 599734
rect 562586 563818 562822 564054
rect 562586 563498 562822 563734
rect 562586 527818 562822 528054
rect 562586 527498 562822 527734
rect 562586 491818 562822 492054
rect 562586 491498 562822 491734
rect 562586 455818 562822 456054
rect 562586 455498 562822 455734
rect 562586 419818 562822 420054
rect 562586 419498 562822 419734
rect 562586 383818 562822 384054
rect 562586 383498 562822 383734
rect 562586 347818 562822 348054
rect 562586 347498 562822 347734
rect 562586 311818 562822 312054
rect 562586 311498 562822 311734
rect 562586 275818 562822 276054
rect 562586 275498 562822 275734
rect 562586 239818 562822 240054
rect 562586 239498 562822 239734
rect 562586 203818 562822 204054
rect 562586 203498 562822 203734
rect 562586 167818 562822 168054
rect 562586 167498 562822 167734
rect 562586 131818 562822 132054
rect 562586 131498 562822 131734
rect 562586 95818 562822 96054
rect 562586 95498 562822 95734
rect 562586 59818 562822 60054
rect 562586 59498 562822 59734
rect 562586 23818 562822 24054
rect 562586 23498 562822 23734
rect 562586 -3402 562822 -3166
rect 562586 -3722 562822 -3486
rect 566186 675418 566422 675654
rect 566186 675098 566422 675334
rect 566186 639418 566422 639654
rect 566186 639098 566422 639334
rect 566186 603418 566422 603654
rect 566186 603098 566422 603334
rect 566186 567418 566422 567654
rect 566186 567098 566422 567334
rect 566186 531418 566422 531654
rect 566186 531098 566422 531334
rect 566186 495418 566422 495654
rect 566186 495098 566422 495334
rect 566186 459418 566422 459654
rect 566186 459098 566422 459334
rect 566186 423418 566422 423654
rect 566186 423098 566422 423334
rect 566186 387418 566422 387654
rect 566186 387098 566422 387334
rect 566186 351418 566422 351654
rect 566186 351098 566422 351334
rect 566186 315418 566422 315654
rect 566186 315098 566422 315334
rect 566186 279418 566422 279654
rect 566186 279098 566422 279334
rect 566186 243418 566422 243654
rect 566186 243098 566422 243334
rect 566186 207418 566422 207654
rect 566186 207098 566422 207334
rect 566186 171418 566422 171654
rect 566186 171098 566422 171334
rect 566186 135418 566422 135654
rect 566186 135098 566422 135334
rect 566186 99418 566422 99654
rect 566186 99098 566422 99334
rect 566186 63418 566422 63654
rect 566186 63098 566422 63334
rect 566186 27418 566422 27654
rect 566186 27098 566422 27334
rect 566186 -5282 566422 -5046
rect 566186 -5602 566422 -5366
rect 592082 711182 592318 711418
rect 592082 710862 592318 711098
rect 591142 710242 591378 710478
rect 591142 709922 591378 710158
rect 590202 709302 590438 709538
rect 590202 708982 590438 709218
rect 589262 708362 589498 708598
rect 589262 708042 589498 708278
rect 588322 707422 588558 707658
rect 588322 707102 588558 707338
rect 580586 706482 580822 706718
rect 580586 706162 580822 706398
rect 569786 679018 570022 679254
rect 569786 678698 570022 678934
rect 569786 643018 570022 643254
rect 569786 642698 570022 642934
rect 569786 607018 570022 607254
rect 569786 606698 570022 606934
rect 569786 571018 570022 571254
rect 569786 570698 570022 570934
rect 569786 535018 570022 535254
rect 569786 534698 570022 534934
rect 569786 499018 570022 499254
rect 569786 498698 570022 498934
rect 569786 463018 570022 463254
rect 569786 462698 570022 462934
rect 569786 427018 570022 427254
rect 569786 426698 570022 426934
rect 569786 391018 570022 391254
rect 569786 390698 570022 390934
rect 569786 355018 570022 355254
rect 569786 354698 570022 354934
rect 569786 319018 570022 319254
rect 569786 318698 570022 318934
rect 569786 283018 570022 283254
rect 569786 282698 570022 282934
rect 569786 247018 570022 247254
rect 569786 246698 570022 246934
rect 569786 211018 570022 211254
rect 569786 210698 570022 210934
rect 569786 175018 570022 175254
rect 569786 174698 570022 174934
rect 569786 139018 570022 139254
rect 569786 138698 570022 138934
rect 569786 103018 570022 103254
rect 569786 102698 570022 102934
rect 569786 67018 570022 67254
rect 569786 66698 570022 66934
rect 569786 31018 570022 31254
rect 569786 30698 570022 30934
rect 551786 -6222 552022 -5986
rect 551786 -6542 552022 -6306
rect 576986 704602 577222 704838
rect 576986 704282 577222 704518
rect 576986 686218 577222 686454
rect 576986 685898 577222 686134
rect 576986 650218 577222 650454
rect 576986 649898 577222 650134
rect 576986 614218 577222 614454
rect 576986 613898 577222 614134
rect 576986 578218 577222 578454
rect 576986 577898 577222 578134
rect 576986 542218 577222 542454
rect 576986 541898 577222 542134
rect 576986 506218 577222 506454
rect 576986 505898 577222 506134
rect 576986 470218 577222 470454
rect 576986 469898 577222 470134
rect 576986 434218 577222 434454
rect 576986 433898 577222 434134
rect 576986 398218 577222 398454
rect 576986 397898 577222 398134
rect 576986 362218 577222 362454
rect 576986 361898 577222 362134
rect 576986 326218 577222 326454
rect 576986 325898 577222 326134
rect 576986 290218 577222 290454
rect 576986 289898 577222 290134
rect 576986 254218 577222 254454
rect 576986 253898 577222 254134
rect 576986 218218 577222 218454
rect 576986 217898 577222 218134
rect 576986 182218 577222 182454
rect 576986 181898 577222 182134
rect 576986 146218 577222 146454
rect 576986 145898 577222 146134
rect 576986 110218 577222 110454
rect 576986 109898 577222 110134
rect 576986 74218 577222 74454
rect 576986 73898 577222 74134
rect 576986 38218 577222 38454
rect 576986 37898 577222 38134
rect 576986 2218 577222 2454
rect 576986 1898 577222 2134
rect 576986 -582 577222 -346
rect 576986 -902 577222 -666
rect 587382 706482 587618 706718
rect 587382 706162 587618 706398
rect 586442 705542 586678 705778
rect 586442 705222 586678 705458
rect 580586 689818 580822 690054
rect 580586 689498 580822 689734
rect 580586 653818 580822 654054
rect 580586 653498 580822 653734
rect 580586 617818 580822 618054
rect 580586 617498 580822 617734
rect 580586 581818 580822 582054
rect 580586 581498 580822 581734
rect 580586 545818 580822 546054
rect 580586 545498 580822 545734
rect 580586 509818 580822 510054
rect 580586 509498 580822 509734
rect 580586 473818 580822 474054
rect 580586 473498 580822 473734
rect 580586 437818 580822 438054
rect 580586 437498 580822 437734
rect 580586 401818 580822 402054
rect 580586 401498 580822 401734
rect 580586 365818 580822 366054
rect 580586 365498 580822 365734
rect 580586 329818 580822 330054
rect 580586 329498 580822 329734
rect 580586 293818 580822 294054
rect 580586 293498 580822 293734
rect 580586 257818 580822 258054
rect 580586 257498 580822 257734
rect 580586 221818 580822 222054
rect 580586 221498 580822 221734
rect 580586 185818 580822 186054
rect 580586 185498 580822 185734
rect 580586 149818 580822 150054
rect 580586 149498 580822 149734
rect 580586 113818 580822 114054
rect 580586 113498 580822 113734
rect 580586 77818 580822 78054
rect 580586 77498 580822 77734
rect 580586 41818 580822 42054
rect 580586 41498 580822 41734
rect 580586 5818 580822 6054
rect 580586 5498 580822 5734
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 686218 585738 686454
rect 585502 685898 585738 686134
rect 585502 650218 585738 650454
rect 585502 649898 585738 650134
rect 585502 614218 585738 614454
rect 585502 613898 585738 614134
rect 585502 578218 585738 578454
rect 585502 577898 585738 578134
rect 585502 542218 585738 542454
rect 585502 541898 585738 542134
rect 585502 506218 585738 506454
rect 585502 505898 585738 506134
rect 585502 470218 585738 470454
rect 585502 469898 585738 470134
rect 585502 434218 585738 434454
rect 585502 433898 585738 434134
rect 585502 398218 585738 398454
rect 585502 397898 585738 398134
rect 585502 362218 585738 362454
rect 585502 361898 585738 362134
rect 585502 326218 585738 326454
rect 585502 325898 585738 326134
rect 585502 290218 585738 290454
rect 585502 289898 585738 290134
rect 585502 254218 585738 254454
rect 585502 253898 585738 254134
rect 585502 218218 585738 218454
rect 585502 217898 585738 218134
rect 585502 182218 585738 182454
rect 585502 181898 585738 182134
rect 585502 146218 585738 146454
rect 585502 145898 585738 146134
rect 585502 110218 585738 110454
rect 585502 109898 585738 110134
rect 585502 74218 585738 74454
rect 585502 73898 585738 74134
rect 585502 38218 585738 38454
rect 585502 37898 585738 38134
rect 585502 2218 585738 2454
rect 585502 1898 585738 2134
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586442 668218 586678 668454
rect 586442 667898 586678 668134
rect 586442 632218 586678 632454
rect 586442 631898 586678 632134
rect 586442 596218 586678 596454
rect 586442 595898 586678 596134
rect 586442 560218 586678 560454
rect 586442 559898 586678 560134
rect 586442 524218 586678 524454
rect 586442 523898 586678 524134
rect 586442 488218 586678 488454
rect 586442 487898 586678 488134
rect 586442 452218 586678 452454
rect 586442 451898 586678 452134
rect 586442 416218 586678 416454
rect 586442 415898 586678 416134
rect 586442 380218 586678 380454
rect 586442 379898 586678 380134
rect 586442 344218 586678 344454
rect 586442 343898 586678 344134
rect 586442 308218 586678 308454
rect 586442 307898 586678 308134
rect 586442 272218 586678 272454
rect 586442 271898 586678 272134
rect 586442 236218 586678 236454
rect 586442 235898 586678 236134
rect 586442 200218 586678 200454
rect 586442 199898 586678 200134
rect 586442 164218 586678 164454
rect 586442 163898 586678 164134
rect 586442 128218 586678 128454
rect 586442 127898 586678 128134
rect 586442 92218 586678 92454
rect 586442 91898 586678 92134
rect 586442 56218 586678 56454
rect 586442 55898 586678 56134
rect 586442 20218 586678 20454
rect 586442 19898 586678 20134
rect 586442 -1522 586678 -1286
rect 586442 -1842 586678 -1606
rect 587382 689818 587618 690054
rect 587382 689498 587618 689734
rect 587382 653818 587618 654054
rect 587382 653498 587618 653734
rect 587382 617818 587618 618054
rect 587382 617498 587618 617734
rect 587382 581818 587618 582054
rect 587382 581498 587618 581734
rect 587382 545818 587618 546054
rect 587382 545498 587618 545734
rect 587382 509818 587618 510054
rect 587382 509498 587618 509734
rect 587382 473818 587618 474054
rect 587382 473498 587618 473734
rect 587382 437818 587618 438054
rect 587382 437498 587618 437734
rect 587382 401818 587618 402054
rect 587382 401498 587618 401734
rect 587382 365818 587618 366054
rect 587382 365498 587618 365734
rect 587382 329818 587618 330054
rect 587382 329498 587618 329734
rect 587382 293818 587618 294054
rect 587382 293498 587618 293734
rect 587382 257818 587618 258054
rect 587382 257498 587618 257734
rect 587382 221818 587618 222054
rect 587382 221498 587618 221734
rect 587382 185818 587618 186054
rect 587382 185498 587618 185734
rect 587382 149818 587618 150054
rect 587382 149498 587618 149734
rect 587382 113818 587618 114054
rect 587382 113498 587618 113734
rect 587382 77818 587618 78054
rect 587382 77498 587618 77734
rect 587382 41818 587618 42054
rect 587382 41498 587618 41734
rect 587382 5818 587618 6054
rect 587382 5498 587618 5734
rect 580586 -2462 580822 -2226
rect 580586 -2782 580822 -2546
rect 587382 -2462 587618 -2226
rect 587382 -2782 587618 -2546
rect 588322 671818 588558 672054
rect 588322 671498 588558 671734
rect 588322 635818 588558 636054
rect 588322 635498 588558 635734
rect 588322 599818 588558 600054
rect 588322 599498 588558 599734
rect 588322 563818 588558 564054
rect 588322 563498 588558 563734
rect 588322 527818 588558 528054
rect 588322 527498 588558 527734
rect 588322 491818 588558 492054
rect 588322 491498 588558 491734
rect 588322 455818 588558 456054
rect 588322 455498 588558 455734
rect 588322 419818 588558 420054
rect 588322 419498 588558 419734
rect 588322 383818 588558 384054
rect 588322 383498 588558 383734
rect 588322 347818 588558 348054
rect 588322 347498 588558 347734
rect 588322 311818 588558 312054
rect 588322 311498 588558 311734
rect 588322 275818 588558 276054
rect 588322 275498 588558 275734
rect 588322 239818 588558 240054
rect 588322 239498 588558 239734
rect 588322 203818 588558 204054
rect 588322 203498 588558 203734
rect 588322 167818 588558 168054
rect 588322 167498 588558 167734
rect 588322 131818 588558 132054
rect 588322 131498 588558 131734
rect 588322 95818 588558 96054
rect 588322 95498 588558 95734
rect 588322 59818 588558 60054
rect 588322 59498 588558 59734
rect 588322 23818 588558 24054
rect 588322 23498 588558 23734
rect 588322 -3402 588558 -3166
rect 588322 -3722 588558 -3486
rect 589262 693418 589498 693654
rect 589262 693098 589498 693334
rect 589262 657418 589498 657654
rect 589262 657098 589498 657334
rect 589262 621418 589498 621654
rect 589262 621098 589498 621334
rect 589262 585418 589498 585654
rect 589262 585098 589498 585334
rect 589262 549418 589498 549654
rect 589262 549098 589498 549334
rect 589262 513418 589498 513654
rect 589262 513098 589498 513334
rect 589262 477418 589498 477654
rect 589262 477098 589498 477334
rect 589262 441418 589498 441654
rect 589262 441098 589498 441334
rect 589262 405418 589498 405654
rect 589262 405098 589498 405334
rect 589262 369418 589498 369654
rect 589262 369098 589498 369334
rect 589262 333418 589498 333654
rect 589262 333098 589498 333334
rect 589262 297418 589498 297654
rect 589262 297098 589498 297334
rect 589262 261418 589498 261654
rect 589262 261098 589498 261334
rect 589262 225418 589498 225654
rect 589262 225098 589498 225334
rect 589262 189418 589498 189654
rect 589262 189098 589498 189334
rect 589262 153418 589498 153654
rect 589262 153098 589498 153334
rect 589262 117418 589498 117654
rect 589262 117098 589498 117334
rect 589262 81418 589498 81654
rect 589262 81098 589498 81334
rect 589262 45418 589498 45654
rect 589262 45098 589498 45334
rect 589262 9418 589498 9654
rect 589262 9098 589498 9334
rect 589262 -4342 589498 -4106
rect 589262 -4662 589498 -4426
rect 590202 675418 590438 675654
rect 590202 675098 590438 675334
rect 590202 639418 590438 639654
rect 590202 639098 590438 639334
rect 590202 603418 590438 603654
rect 590202 603098 590438 603334
rect 590202 567418 590438 567654
rect 590202 567098 590438 567334
rect 590202 531418 590438 531654
rect 590202 531098 590438 531334
rect 590202 495418 590438 495654
rect 590202 495098 590438 495334
rect 590202 459418 590438 459654
rect 590202 459098 590438 459334
rect 590202 423418 590438 423654
rect 590202 423098 590438 423334
rect 590202 387418 590438 387654
rect 590202 387098 590438 387334
rect 590202 351418 590438 351654
rect 590202 351098 590438 351334
rect 590202 315418 590438 315654
rect 590202 315098 590438 315334
rect 590202 279418 590438 279654
rect 590202 279098 590438 279334
rect 590202 243418 590438 243654
rect 590202 243098 590438 243334
rect 590202 207418 590438 207654
rect 590202 207098 590438 207334
rect 590202 171418 590438 171654
rect 590202 171098 590438 171334
rect 590202 135418 590438 135654
rect 590202 135098 590438 135334
rect 590202 99418 590438 99654
rect 590202 99098 590438 99334
rect 590202 63418 590438 63654
rect 590202 63098 590438 63334
rect 590202 27418 590438 27654
rect 590202 27098 590438 27334
rect 590202 -5282 590438 -5046
rect 590202 -5602 590438 -5366
rect 591142 697018 591378 697254
rect 591142 696698 591378 696934
rect 591142 661018 591378 661254
rect 591142 660698 591378 660934
rect 591142 625018 591378 625254
rect 591142 624698 591378 624934
rect 591142 589018 591378 589254
rect 591142 588698 591378 588934
rect 591142 553018 591378 553254
rect 591142 552698 591378 552934
rect 591142 517018 591378 517254
rect 591142 516698 591378 516934
rect 591142 481018 591378 481254
rect 591142 480698 591378 480934
rect 591142 445018 591378 445254
rect 591142 444698 591378 444934
rect 591142 409018 591378 409254
rect 591142 408698 591378 408934
rect 591142 373018 591378 373254
rect 591142 372698 591378 372934
rect 591142 337018 591378 337254
rect 591142 336698 591378 336934
rect 591142 301018 591378 301254
rect 591142 300698 591378 300934
rect 591142 265018 591378 265254
rect 591142 264698 591378 264934
rect 591142 229018 591378 229254
rect 591142 228698 591378 228934
rect 591142 193018 591378 193254
rect 591142 192698 591378 192934
rect 591142 157018 591378 157254
rect 591142 156698 591378 156934
rect 591142 121018 591378 121254
rect 591142 120698 591378 120934
rect 591142 85018 591378 85254
rect 591142 84698 591378 84934
rect 591142 49018 591378 49254
rect 591142 48698 591378 48934
rect 591142 13018 591378 13254
rect 591142 12698 591378 12934
rect 591142 -6222 591378 -5986
rect 591142 -6542 591378 -6306
rect 592082 679018 592318 679254
rect 592082 678698 592318 678934
rect 592082 643018 592318 643254
rect 592082 642698 592318 642934
rect 592082 607018 592318 607254
rect 592082 606698 592318 606934
rect 592082 571018 592318 571254
rect 592082 570698 592318 570934
rect 592082 535018 592318 535254
rect 592082 534698 592318 534934
rect 592082 499018 592318 499254
rect 592082 498698 592318 498934
rect 592082 463018 592318 463254
rect 592082 462698 592318 462934
rect 592082 427018 592318 427254
rect 592082 426698 592318 426934
rect 592082 391018 592318 391254
rect 592082 390698 592318 390934
rect 592082 355018 592318 355254
rect 592082 354698 592318 354934
rect 592082 319018 592318 319254
rect 592082 318698 592318 318934
rect 592082 283018 592318 283254
rect 592082 282698 592318 282934
rect 592082 247018 592318 247254
rect 592082 246698 592318 246934
rect 592082 211018 592318 211254
rect 592082 210698 592318 210934
rect 592082 175018 592318 175254
rect 592082 174698 592318 174934
rect 592082 139018 592318 139254
rect 592082 138698 592318 138934
rect 592082 103018 592318 103254
rect 592082 102698 592318 102934
rect 592082 67018 592318 67254
rect 592082 66698 592318 66934
rect 592082 31018 592318 31254
rect 592082 30698 592318 30934
rect 569786 -7162 570022 -6926
rect 569786 -7482 570022 -7246
rect 592082 -7162 592318 -6926
rect 592082 -7482 592318 -7246
<< metal5 >>
rect -8576 711440 -7976 711442
rect 29604 711440 30204 711442
rect 65604 711440 66204 711442
rect 101604 711440 102204 711442
rect 137604 711440 138204 711442
rect 173604 711440 174204 711442
rect 209604 711440 210204 711442
rect 245604 711440 246204 711442
rect 281604 711440 282204 711442
rect 317604 711440 318204 711442
rect 353604 711440 354204 711442
rect 389604 711440 390204 711442
rect 425604 711440 426204 711442
rect 461604 711440 462204 711442
rect 497604 711440 498204 711442
rect 533604 711440 534204 711442
rect 569604 711440 570204 711442
rect 591900 711440 592500 711442
rect -8576 711418 592500 711440
rect -8576 711182 -8394 711418
rect -8158 711182 29786 711418
rect 30022 711182 65786 711418
rect 66022 711182 101786 711418
rect 102022 711182 137786 711418
rect 138022 711182 173786 711418
rect 174022 711182 209786 711418
rect 210022 711182 245786 711418
rect 246022 711182 281786 711418
rect 282022 711182 317786 711418
rect 318022 711182 353786 711418
rect 354022 711182 389786 711418
rect 390022 711182 425786 711418
rect 426022 711182 461786 711418
rect 462022 711182 497786 711418
rect 498022 711182 533786 711418
rect 534022 711182 569786 711418
rect 570022 711182 592082 711418
rect 592318 711182 592500 711418
rect -8576 711098 592500 711182
rect -8576 710862 -8394 711098
rect -8158 710862 29786 711098
rect 30022 710862 65786 711098
rect 66022 710862 101786 711098
rect 102022 710862 137786 711098
rect 138022 710862 173786 711098
rect 174022 710862 209786 711098
rect 210022 710862 245786 711098
rect 246022 710862 281786 711098
rect 282022 710862 317786 711098
rect 318022 710862 353786 711098
rect 354022 710862 389786 711098
rect 390022 710862 425786 711098
rect 426022 710862 461786 711098
rect 462022 710862 497786 711098
rect 498022 710862 533786 711098
rect 534022 710862 569786 711098
rect 570022 710862 592082 711098
rect 592318 710862 592500 711098
rect -8576 710840 592500 710862
rect -8576 710838 -7976 710840
rect 29604 710838 30204 710840
rect 65604 710838 66204 710840
rect 101604 710838 102204 710840
rect 137604 710838 138204 710840
rect 173604 710838 174204 710840
rect 209604 710838 210204 710840
rect 245604 710838 246204 710840
rect 281604 710838 282204 710840
rect 317604 710838 318204 710840
rect 353604 710838 354204 710840
rect 389604 710838 390204 710840
rect 425604 710838 426204 710840
rect 461604 710838 462204 710840
rect 497604 710838 498204 710840
rect 533604 710838 534204 710840
rect 569604 710838 570204 710840
rect 591900 710838 592500 710840
rect -7636 710500 -7036 710502
rect 11604 710500 12204 710502
rect 47604 710500 48204 710502
rect 83604 710500 84204 710502
rect 119604 710500 120204 710502
rect 155604 710500 156204 710502
rect 191604 710500 192204 710502
rect 227604 710500 228204 710502
rect 263604 710500 264204 710502
rect 299604 710500 300204 710502
rect 335604 710500 336204 710502
rect 371604 710500 372204 710502
rect 407604 710500 408204 710502
rect 443604 710500 444204 710502
rect 479604 710500 480204 710502
rect 515604 710500 516204 710502
rect 551604 710500 552204 710502
rect 590960 710500 591560 710502
rect -7636 710478 591560 710500
rect -7636 710242 -7454 710478
rect -7218 710242 11786 710478
rect 12022 710242 47786 710478
rect 48022 710242 83786 710478
rect 84022 710242 119786 710478
rect 120022 710242 155786 710478
rect 156022 710242 191786 710478
rect 192022 710242 227786 710478
rect 228022 710242 263786 710478
rect 264022 710242 299786 710478
rect 300022 710242 335786 710478
rect 336022 710242 371786 710478
rect 372022 710242 407786 710478
rect 408022 710242 443786 710478
rect 444022 710242 479786 710478
rect 480022 710242 515786 710478
rect 516022 710242 551786 710478
rect 552022 710242 591142 710478
rect 591378 710242 591560 710478
rect -7636 710158 591560 710242
rect -7636 709922 -7454 710158
rect -7218 709922 11786 710158
rect 12022 709922 47786 710158
rect 48022 709922 83786 710158
rect 84022 709922 119786 710158
rect 120022 709922 155786 710158
rect 156022 709922 191786 710158
rect 192022 709922 227786 710158
rect 228022 709922 263786 710158
rect 264022 709922 299786 710158
rect 300022 709922 335786 710158
rect 336022 709922 371786 710158
rect 372022 709922 407786 710158
rect 408022 709922 443786 710158
rect 444022 709922 479786 710158
rect 480022 709922 515786 710158
rect 516022 709922 551786 710158
rect 552022 709922 591142 710158
rect 591378 709922 591560 710158
rect -7636 709900 591560 709922
rect -7636 709898 -7036 709900
rect 11604 709898 12204 709900
rect 47604 709898 48204 709900
rect 83604 709898 84204 709900
rect 119604 709898 120204 709900
rect 155604 709898 156204 709900
rect 191604 709898 192204 709900
rect 227604 709898 228204 709900
rect 263604 709898 264204 709900
rect 299604 709898 300204 709900
rect 335604 709898 336204 709900
rect 371604 709898 372204 709900
rect 407604 709898 408204 709900
rect 443604 709898 444204 709900
rect 479604 709898 480204 709900
rect 515604 709898 516204 709900
rect 551604 709898 552204 709900
rect 590960 709898 591560 709900
rect -6696 709560 -6096 709562
rect 26004 709560 26604 709562
rect 62004 709560 62604 709562
rect 98004 709560 98604 709562
rect 134004 709560 134604 709562
rect 170004 709560 170604 709562
rect 206004 709560 206604 709562
rect 242004 709560 242604 709562
rect 278004 709560 278604 709562
rect 314004 709560 314604 709562
rect 350004 709560 350604 709562
rect 386004 709560 386604 709562
rect 422004 709560 422604 709562
rect 458004 709560 458604 709562
rect 494004 709560 494604 709562
rect 530004 709560 530604 709562
rect 566004 709560 566604 709562
rect 590020 709560 590620 709562
rect -6696 709538 590620 709560
rect -6696 709302 -6514 709538
rect -6278 709302 26186 709538
rect 26422 709302 62186 709538
rect 62422 709302 98186 709538
rect 98422 709302 134186 709538
rect 134422 709302 170186 709538
rect 170422 709302 206186 709538
rect 206422 709302 242186 709538
rect 242422 709302 278186 709538
rect 278422 709302 314186 709538
rect 314422 709302 350186 709538
rect 350422 709302 386186 709538
rect 386422 709302 422186 709538
rect 422422 709302 458186 709538
rect 458422 709302 494186 709538
rect 494422 709302 530186 709538
rect 530422 709302 566186 709538
rect 566422 709302 590202 709538
rect 590438 709302 590620 709538
rect -6696 709218 590620 709302
rect -6696 708982 -6514 709218
rect -6278 708982 26186 709218
rect 26422 708982 62186 709218
rect 62422 708982 98186 709218
rect 98422 708982 134186 709218
rect 134422 708982 170186 709218
rect 170422 708982 206186 709218
rect 206422 708982 242186 709218
rect 242422 708982 278186 709218
rect 278422 708982 314186 709218
rect 314422 708982 350186 709218
rect 350422 708982 386186 709218
rect 386422 708982 422186 709218
rect 422422 708982 458186 709218
rect 458422 708982 494186 709218
rect 494422 708982 530186 709218
rect 530422 708982 566186 709218
rect 566422 708982 590202 709218
rect 590438 708982 590620 709218
rect -6696 708960 590620 708982
rect -6696 708958 -6096 708960
rect 26004 708958 26604 708960
rect 62004 708958 62604 708960
rect 98004 708958 98604 708960
rect 134004 708958 134604 708960
rect 170004 708958 170604 708960
rect 206004 708958 206604 708960
rect 242004 708958 242604 708960
rect 278004 708958 278604 708960
rect 314004 708958 314604 708960
rect 350004 708958 350604 708960
rect 386004 708958 386604 708960
rect 422004 708958 422604 708960
rect 458004 708958 458604 708960
rect 494004 708958 494604 708960
rect 530004 708958 530604 708960
rect 566004 708958 566604 708960
rect 590020 708958 590620 708960
rect -5756 708620 -5156 708622
rect 8004 708620 8604 708622
rect 44004 708620 44604 708622
rect 80004 708620 80604 708622
rect 116004 708620 116604 708622
rect 152004 708620 152604 708622
rect 188004 708620 188604 708622
rect 224004 708620 224604 708622
rect 260004 708620 260604 708622
rect 296004 708620 296604 708622
rect 332004 708620 332604 708622
rect 368004 708620 368604 708622
rect 404004 708620 404604 708622
rect 440004 708620 440604 708622
rect 476004 708620 476604 708622
rect 512004 708620 512604 708622
rect 548004 708620 548604 708622
rect 589080 708620 589680 708622
rect -5756 708598 589680 708620
rect -5756 708362 -5574 708598
rect -5338 708362 8186 708598
rect 8422 708362 44186 708598
rect 44422 708362 80186 708598
rect 80422 708362 116186 708598
rect 116422 708362 152186 708598
rect 152422 708362 188186 708598
rect 188422 708362 224186 708598
rect 224422 708362 260186 708598
rect 260422 708362 296186 708598
rect 296422 708362 332186 708598
rect 332422 708362 368186 708598
rect 368422 708362 404186 708598
rect 404422 708362 440186 708598
rect 440422 708362 476186 708598
rect 476422 708362 512186 708598
rect 512422 708362 548186 708598
rect 548422 708362 589262 708598
rect 589498 708362 589680 708598
rect -5756 708278 589680 708362
rect -5756 708042 -5574 708278
rect -5338 708042 8186 708278
rect 8422 708042 44186 708278
rect 44422 708042 80186 708278
rect 80422 708042 116186 708278
rect 116422 708042 152186 708278
rect 152422 708042 188186 708278
rect 188422 708042 224186 708278
rect 224422 708042 260186 708278
rect 260422 708042 296186 708278
rect 296422 708042 332186 708278
rect 332422 708042 368186 708278
rect 368422 708042 404186 708278
rect 404422 708042 440186 708278
rect 440422 708042 476186 708278
rect 476422 708042 512186 708278
rect 512422 708042 548186 708278
rect 548422 708042 589262 708278
rect 589498 708042 589680 708278
rect -5756 708020 589680 708042
rect -5756 708018 -5156 708020
rect 8004 708018 8604 708020
rect 44004 708018 44604 708020
rect 80004 708018 80604 708020
rect 116004 708018 116604 708020
rect 152004 708018 152604 708020
rect 188004 708018 188604 708020
rect 224004 708018 224604 708020
rect 260004 708018 260604 708020
rect 296004 708018 296604 708020
rect 332004 708018 332604 708020
rect 368004 708018 368604 708020
rect 404004 708018 404604 708020
rect 440004 708018 440604 708020
rect 476004 708018 476604 708020
rect 512004 708018 512604 708020
rect 548004 708018 548604 708020
rect 589080 708018 589680 708020
rect -4816 707680 -4216 707682
rect 22404 707680 23004 707682
rect 58404 707680 59004 707682
rect 94404 707680 95004 707682
rect 130404 707680 131004 707682
rect 166404 707680 167004 707682
rect 202404 707680 203004 707682
rect 238404 707680 239004 707682
rect 274404 707680 275004 707682
rect 310404 707680 311004 707682
rect 346404 707680 347004 707682
rect 382404 707680 383004 707682
rect 418404 707680 419004 707682
rect 454404 707680 455004 707682
rect 490404 707680 491004 707682
rect 526404 707680 527004 707682
rect 562404 707680 563004 707682
rect 588140 707680 588740 707682
rect -4816 707658 588740 707680
rect -4816 707422 -4634 707658
rect -4398 707422 22586 707658
rect 22822 707422 58586 707658
rect 58822 707422 94586 707658
rect 94822 707422 130586 707658
rect 130822 707422 166586 707658
rect 166822 707422 202586 707658
rect 202822 707422 238586 707658
rect 238822 707422 274586 707658
rect 274822 707422 310586 707658
rect 310822 707422 346586 707658
rect 346822 707422 382586 707658
rect 382822 707422 418586 707658
rect 418822 707422 454586 707658
rect 454822 707422 490586 707658
rect 490822 707422 526586 707658
rect 526822 707422 562586 707658
rect 562822 707422 588322 707658
rect 588558 707422 588740 707658
rect -4816 707338 588740 707422
rect -4816 707102 -4634 707338
rect -4398 707102 22586 707338
rect 22822 707102 58586 707338
rect 58822 707102 94586 707338
rect 94822 707102 130586 707338
rect 130822 707102 166586 707338
rect 166822 707102 202586 707338
rect 202822 707102 238586 707338
rect 238822 707102 274586 707338
rect 274822 707102 310586 707338
rect 310822 707102 346586 707338
rect 346822 707102 382586 707338
rect 382822 707102 418586 707338
rect 418822 707102 454586 707338
rect 454822 707102 490586 707338
rect 490822 707102 526586 707338
rect 526822 707102 562586 707338
rect 562822 707102 588322 707338
rect 588558 707102 588740 707338
rect -4816 707080 588740 707102
rect -4816 707078 -4216 707080
rect 22404 707078 23004 707080
rect 58404 707078 59004 707080
rect 94404 707078 95004 707080
rect 130404 707078 131004 707080
rect 166404 707078 167004 707080
rect 202404 707078 203004 707080
rect 238404 707078 239004 707080
rect 274404 707078 275004 707080
rect 310404 707078 311004 707080
rect 346404 707078 347004 707080
rect 382404 707078 383004 707080
rect 418404 707078 419004 707080
rect 454404 707078 455004 707080
rect 490404 707078 491004 707080
rect 526404 707078 527004 707080
rect 562404 707078 563004 707080
rect 588140 707078 588740 707080
rect -3876 706740 -3276 706742
rect 4404 706740 5004 706742
rect 40404 706740 41004 706742
rect 76404 706740 77004 706742
rect 112404 706740 113004 706742
rect 148404 706740 149004 706742
rect 184404 706740 185004 706742
rect 220404 706740 221004 706742
rect 256404 706740 257004 706742
rect 292404 706740 293004 706742
rect 328404 706740 329004 706742
rect 364404 706740 365004 706742
rect 400404 706740 401004 706742
rect 436404 706740 437004 706742
rect 472404 706740 473004 706742
rect 508404 706740 509004 706742
rect 544404 706740 545004 706742
rect 580404 706740 581004 706742
rect 587200 706740 587800 706742
rect -3876 706718 587800 706740
rect -3876 706482 -3694 706718
rect -3458 706482 4586 706718
rect 4822 706482 40586 706718
rect 40822 706482 76586 706718
rect 76822 706482 112586 706718
rect 112822 706482 148586 706718
rect 148822 706482 184586 706718
rect 184822 706482 220586 706718
rect 220822 706482 256586 706718
rect 256822 706482 292586 706718
rect 292822 706482 328586 706718
rect 328822 706482 364586 706718
rect 364822 706482 400586 706718
rect 400822 706482 436586 706718
rect 436822 706482 472586 706718
rect 472822 706482 508586 706718
rect 508822 706482 544586 706718
rect 544822 706482 580586 706718
rect 580822 706482 587382 706718
rect 587618 706482 587800 706718
rect -3876 706398 587800 706482
rect -3876 706162 -3694 706398
rect -3458 706162 4586 706398
rect 4822 706162 40586 706398
rect 40822 706162 76586 706398
rect 76822 706162 112586 706398
rect 112822 706162 148586 706398
rect 148822 706162 184586 706398
rect 184822 706162 220586 706398
rect 220822 706162 256586 706398
rect 256822 706162 292586 706398
rect 292822 706162 328586 706398
rect 328822 706162 364586 706398
rect 364822 706162 400586 706398
rect 400822 706162 436586 706398
rect 436822 706162 472586 706398
rect 472822 706162 508586 706398
rect 508822 706162 544586 706398
rect 544822 706162 580586 706398
rect 580822 706162 587382 706398
rect 587618 706162 587800 706398
rect -3876 706140 587800 706162
rect -3876 706138 -3276 706140
rect 4404 706138 5004 706140
rect 40404 706138 41004 706140
rect 76404 706138 77004 706140
rect 112404 706138 113004 706140
rect 148404 706138 149004 706140
rect 184404 706138 185004 706140
rect 220404 706138 221004 706140
rect 256404 706138 257004 706140
rect 292404 706138 293004 706140
rect 328404 706138 329004 706140
rect 364404 706138 365004 706140
rect 400404 706138 401004 706140
rect 436404 706138 437004 706140
rect 472404 706138 473004 706140
rect 508404 706138 509004 706140
rect 544404 706138 545004 706140
rect 580404 706138 581004 706140
rect 587200 706138 587800 706140
rect -2936 705800 -2336 705802
rect 18804 705800 19404 705802
rect 54804 705800 55404 705802
rect 90804 705800 91404 705802
rect 126804 705800 127404 705802
rect 162804 705800 163404 705802
rect 198804 705800 199404 705802
rect 234804 705800 235404 705802
rect 270804 705800 271404 705802
rect 306804 705800 307404 705802
rect 342804 705800 343404 705802
rect 378804 705800 379404 705802
rect 414804 705800 415404 705802
rect 450804 705800 451404 705802
rect 486804 705800 487404 705802
rect 522804 705800 523404 705802
rect 558804 705800 559404 705802
rect 586260 705800 586860 705802
rect -2936 705778 586860 705800
rect -2936 705542 -2754 705778
rect -2518 705542 18986 705778
rect 19222 705542 54986 705778
rect 55222 705542 90986 705778
rect 91222 705542 126986 705778
rect 127222 705542 162986 705778
rect 163222 705542 198986 705778
rect 199222 705542 234986 705778
rect 235222 705542 270986 705778
rect 271222 705542 306986 705778
rect 307222 705542 342986 705778
rect 343222 705542 378986 705778
rect 379222 705542 414986 705778
rect 415222 705542 450986 705778
rect 451222 705542 486986 705778
rect 487222 705542 522986 705778
rect 523222 705542 558986 705778
rect 559222 705542 586442 705778
rect 586678 705542 586860 705778
rect -2936 705458 586860 705542
rect -2936 705222 -2754 705458
rect -2518 705222 18986 705458
rect 19222 705222 54986 705458
rect 55222 705222 90986 705458
rect 91222 705222 126986 705458
rect 127222 705222 162986 705458
rect 163222 705222 198986 705458
rect 199222 705222 234986 705458
rect 235222 705222 270986 705458
rect 271222 705222 306986 705458
rect 307222 705222 342986 705458
rect 343222 705222 378986 705458
rect 379222 705222 414986 705458
rect 415222 705222 450986 705458
rect 451222 705222 486986 705458
rect 487222 705222 522986 705458
rect 523222 705222 558986 705458
rect 559222 705222 586442 705458
rect 586678 705222 586860 705458
rect -2936 705200 586860 705222
rect -2936 705198 -2336 705200
rect 18804 705198 19404 705200
rect 54804 705198 55404 705200
rect 90804 705198 91404 705200
rect 126804 705198 127404 705200
rect 162804 705198 163404 705200
rect 198804 705198 199404 705200
rect 234804 705198 235404 705200
rect 270804 705198 271404 705200
rect 306804 705198 307404 705200
rect 342804 705198 343404 705200
rect 378804 705198 379404 705200
rect 414804 705198 415404 705200
rect 450804 705198 451404 705200
rect 486804 705198 487404 705200
rect 522804 705198 523404 705200
rect 558804 705198 559404 705200
rect 586260 705198 586860 705200
rect -1996 704860 -1396 704862
rect 804 704860 1404 704862
rect 36804 704860 37404 704862
rect 72804 704860 73404 704862
rect 108804 704860 109404 704862
rect 144804 704860 145404 704862
rect 180804 704860 181404 704862
rect 216804 704860 217404 704862
rect 252804 704860 253404 704862
rect 288804 704860 289404 704862
rect 324804 704860 325404 704862
rect 360804 704860 361404 704862
rect 396804 704860 397404 704862
rect 432804 704860 433404 704862
rect 468804 704860 469404 704862
rect 504804 704860 505404 704862
rect 540804 704860 541404 704862
rect 576804 704860 577404 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 986 704838
rect 1222 704602 36986 704838
rect 37222 704602 72986 704838
rect 73222 704602 108986 704838
rect 109222 704602 144986 704838
rect 145222 704602 180986 704838
rect 181222 704602 216986 704838
rect 217222 704602 252986 704838
rect 253222 704602 288986 704838
rect 289222 704602 324986 704838
rect 325222 704602 360986 704838
rect 361222 704602 396986 704838
rect 397222 704602 432986 704838
rect 433222 704602 468986 704838
rect 469222 704602 504986 704838
rect 505222 704602 540986 704838
rect 541222 704602 576986 704838
rect 577222 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 986 704518
rect 1222 704282 36986 704518
rect 37222 704282 72986 704518
rect 73222 704282 108986 704518
rect 109222 704282 144986 704518
rect 145222 704282 180986 704518
rect 181222 704282 216986 704518
rect 217222 704282 252986 704518
rect 253222 704282 288986 704518
rect 289222 704282 324986 704518
rect 325222 704282 360986 704518
rect 361222 704282 396986 704518
rect 397222 704282 432986 704518
rect 433222 704282 468986 704518
rect 469222 704282 504986 704518
rect 505222 704282 540986 704518
rect 541222 704282 576986 704518
rect 577222 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 804 704258 1404 704260
rect 36804 704258 37404 704260
rect 72804 704258 73404 704260
rect 108804 704258 109404 704260
rect 144804 704258 145404 704260
rect 180804 704258 181404 704260
rect 216804 704258 217404 704260
rect 252804 704258 253404 704260
rect 288804 704258 289404 704260
rect 324804 704258 325404 704260
rect 360804 704258 361404 704260
rect 396804 704258 397404 704260
rect 432804 704258 433404 704260
rect 468804 704258 469404 704260
rect 504804 704258 505404 704260
rect 540804 704258 541404 704260
rect 576804 704258 577404 704260
rect 585320 704258 585920 704260
rect -7636 697276 -7036 697278
rect 11604 697276 12204 697278
rect 47604 697276 48204 697278
rect 83604 697276 84204 697278
rect 119604 697276 120204 697278
rect 155604 697276 156204 697278
rect 191604 697276 192204 697278
rect 227604 697276 228204 697278
rect 263604 697276 264204 697278
rect 299604 697276 300204 697278
rect 335604 697276 336204 697278
rect 371604 697276 372204 697278
rect 407604 697276 408204 697278
rect 443604 697276 444204 697278
rect 479604 697276 480204 697278
rect 515604 697276 516204 697278
rect 551604 697276 552204 697278
rect 590960 697276 591560 697278
rect -8576 697254 592500 697276
rect -8576 697018 -7454 697254
rect -7218 697018 11786 697254
rect 12022 697018 47786 697254
rect 48022 697018 83786 697254
rect 84022 697018 119786 697254
rect 120022 697018 155786 697254
rect 156022 697018 191786 697254
rect 192022 697018 227786 697254
rect 228022 697018 263786 697254
rect 264022 697018 299786 697254
rect 300022 697018 335786 697254
rect 336022 697018 371786 697254
rect 372022 697018 407786 697254
rect 408022 697018 443786 697254
rect 444022 697018 479786 697254
rect 480022 697018 515786 697254
rect 516022 697018 551786 697254
rect 552022 697018 591142 697254
rect 591378 697018 592500 697254
rect -8576 696934 592500 697018
rect -8576 696698 -7454 696934
rect -7218 696698 11786 696934
rect 12022 696698 47786 696934
rect 48022 696698 83786 696934
rect 84022 696698 119786 696934
rect 120022 696698 155786 696934
rect 156022 696698 191786 696934
rect 192022 696698 227786 696934
rect 228022 696698 263786 696934
rect 264022 696698 299786 696934
rect 300022 696698 335786 696934
rect 336022 696698 371786 696934
rect 372022 696698 407786 696934
rect 408022 696698 443786 696934
rect 444022 696698 479786 696934
rect 480022 696698 515786 696934
rect 516022 696698 551786 696934
rect 552022 696698 591142 696934
rect 591378 696698 592500 696934
rect -8576 696676 592500 696698
rect -7636 696674 -7036 696676
rect 11604 696674 12204 696676
rect 47604 696674 48204 696676
rect 83604 696674 84204 696676
rect 119604 696674 120204 696676
rect 155604 696674 156204 696676
rect 191604 696674 192204 696676
rect 227604 696674 228204 696676
rect 263604 696674 264204 696676
rect 299604 696674 300204 696676
rect 335604 696674 336204 696676
rect 371604 696674 372204 696676
rect 407604 696674 408204 696676
rect 443604 696674 444204 696676
rect 479604 696674 480204 696676
rect 515604 696674 516204 696676
rect 551604 696674 552204 696676
rect 590960 696674 591560 696676
rect -5756 693676 -5156 693678
rect 8004 693676 8604 693678
rect 44004 693676 44604 693678
rect 80004 693676 80604 693678
rect 116004 693676 116604 693678
rect 152004 693676 152604 693678
rect 188004 693676 188604 693678
rect 224004 693676 224604 693678
rect 260004 693676 260604 693678
rect 296004 693676 296604 693678
rect 332004 693676 332604 693678
rect 368004 693676 368604 693678
rect 404004 693676 404604 693678
rect 440004 693676 440604 693678
rect 476004 693676 476604 693678
rect 512004 693676 512604 693678
rect 548004 693676 548604 693678
rect 589080 693676 589680 693678
rect -6696 693654 590620 693676
rect -6696 693418 -5574 693654
rect -5338 693418 8186 693654
rect 8422 693418 44186 693654
rect 44422 693418 80186 693654
rect 80422 693418 116186 693654
rect 116422 693418 152186 693654
rect 152422 693418 188186 693654
rect 188422 693418 224186 693654
rect 224422 693418 260186 693654
rect 260422 693418 296186 693654
rect 296422 693418 332186 693654
rect 332422 693418 368186 693654
rect 368422 693418 404186 693654
rect 404422 693418 440186 693654
rect 440422 693418 476186 693654
rect 476422 693418 512186 693654
rect 512422 693418 548186 693654
rect 548422 693418 589262 693654
rect 589498 693418 590620 693654
rect -6696 693334 590620 693418
rect -6696 693098 -5574 693334
rect -5338 693098 8186 693334
rect 8422 693098 44186 693334
rect 44422 693098 80186 693334
rect 80422 693098 116186 693334
rect 116422 693098 152186 693334
rect 152422 693098 188186 693334
rect 188422 693098 224186 693334
rect 224422 693098 260186 693334
rect 260422 693098 296186 693334
rect 296422 693098 332186 693334
rect 332422 693098 368186 693334
rect 368422 693098 404186 693334
rect 404422 693098 440186 693334
rect 440422 693098 476186 693334
rect 476422 693098 512186 693334
rect 512422 693098 548186 693334
rect 548422 693098 589262 693334
rect 589498 693098 590620 693334
rect -6696 693076 590620 693098
rect -5756 693074 -5156 693076
rect 8004 693074 8604 693076
rect 44004 693074 44604 693076
rect 80004 693074 80604 693076
rect 116004 693074 116604 693076
rect 152004 693074 152604 693076
rect 188004 693074 188604 693076
rect 224004 693074 224604 693076
rect 260004 693074 260604 693076
rect 296004 693074 296604 693076
rect 332004 693074 332604 693076
rect 368004 693074 368604 693076
rect 404004 693074 404604 693076
rect 440004 693074 440604 693076
rect 476004 693074 476604 693076
rect 512004 693074 512604 693076
rect 548004 693074 548604 693076
rect 589080 693074 589680 693076
rect -3876 690076 -3276 690078
rect 4404 690076 5004 690078
rect 40404 690076 41004 690078
rect 76404 690076 77004 690078
rect 112404 690076 113004 690078
rect 148404 690076 149004 690078
rect 184404 690076 185004 690078
rect 220404 690076 221004 690078
rect 256404 690076 257004 690078
rect 292404 690076 293004 690078
rect 328404 690076 329004 690078
rect 364404 690076 365004 690078
rect 400404 690076 401004 690078
rect 436404 690076 437004 690078
rect 472404 690076 473004 690078
rect 508404 690076 509004 690078
rect 544404 690076 545004 690078
rect 580404 690076 581004 690078
rect 587200 690076 587800 690078
rect -4816 690054 588740 690076
rect -4816 689818 -3694 690054
rect -3458 689818 4586 690054
rect 4822 689818 40586 690054
rect 40822 689818 76586 690054
rect 76822 689818 112586 690054
rect 112822 689818 148586 690054
rect 148822 689818 184586 690054
rect 184822 689818 220586 690054
rect 220822 689818 256586 690054
rect 256822 689818 292586 690054
rect 292822 689818 328586 690054
rect 328822 689818 364586 690054
rect 364822 689818 400586 690054
rect 400822 689818 436586 690054
rect 436822 689818 472586 690054
rect 472822 689818 508586 690054
rect 508822 689818 544586 690054
rect 544822 689818 580586 690054
rect 580822 689818 587382 690054
rect 587618 689818 588740 690054
rect -4816 689734 588740 689818
rect -4816 689498 -3694 689734
rect -3458 689498 4586 689734
rect 4822 689498 40586 689734
rect 40822 689498 76586 689734
rect 76822 689498 112586 689734
rect 112822 689498 148586 689734
rect 148822 689498 184586 689734
rect 184822 689498 220586 689734
rect 220822 689498 256586 689734
rect 256822 689498 292586 689734
rect 292822 689498 328586 689734
rect 328822 689498 364586 689734
rect 364822 689498 400586 689734
rect 400822 689498 436586 689734
rect 436822 689498 472586 689734
rect 472822 689498 508586 689734
rect 508822 689498 544586 689734
rect 544822 689498 580586 689734
rect 580822 689498 587382 689734
rect 587618 689498 588740 689734
rect -4816 689476 588740 689498
rect -3876 689474 -3276 689476
rect 4404 689474 5004 689476
rect 40404 689474 41004 689476
rect 76404 689474 77004 689476
rect 112404 689474 113004 689476
rect 148404 689474 149004 689476
rect 184404 689474 185004 689476
rect 220404 689474 221004 689476
rect 256404 689474 257004 689476
rect 292404 689474 293004 689476
rect 328404 689474 329004 689476
rect 364404 689474 365004 689476
rect 400404 689474 401004 689476
rect 436404 689474 437004 689476
rect 472404 689474 473004 689476
rect 508404 689474 509004 689476
rect 544404 689474 545004 689476
rect 580404 689474 581004 689476
rect 587200 689474 587800 689476
rect -1996 686476 -1396 686478
rect 804 686476 1404 686478
rect 36804 686476 37404 686478
rect 72804 686476 73404 686478
rect 108804 686476 109404 686478
rect 144804 686476 145404 686478
rect 180804 686476 181404 686478
rect 216804 686476 217404 686478
rect 252804 686476 253404 686478
rect 288804 686476 289404 686478
rect 324804 686476 325404 686478
rect 360804 686476 361404 686478
rect 396804 686476 397404 686478
rect 432804 686476 433404 686478
rect 468804 686476 469404 686478
rect 504804 686476 505404 686478
rect 540804 686476 541404 686478
rect 576804 686476 577404 686478
rect 585320 686476 585920 686478
rect -2936 686454 586860 686476
rect -2936 686218 -1814 686454
rect -1578 686218 986 686454
rect 1222 686218 36986 686454
rect 37222 686218 72986 686454
rect 73222 686218 108986 686454
rect 109222 686218 144986 686454
rect 145222 686218 180986 686454
rect 181222 686218 216986 686454
rect 217222 686218 252986 686454
rect 253222 686218 288986 686454
rect 289222 686218 324986 686454
rect 325222 686218 360986 686454
rect 361222 686218 396986 686454
rect 397222 686218 432986 686454
rect 433222 686218 468986 686454
rect 469222 686218 504986 686454
rect 505222 686218 540986 686454
rect 541222 686218 576986 686454
rect 577222 686218 585502 686454
rect 585738 686218 586860 686454
rect -2936 686134 586860 686218
rect -2936 685898 -1814 686134
rect -1578 685898 986 686134
rect 1222 685898 36986 686134
rect 37222 685898 72986 686134
rect 73222 685898 108986 686134
rect 109222 685898 144986 686134
rect 145222 685898 180986 686134
rect 181222 685898 216986 686134
rect 217222 685898 252986 686134
rect 253222 685898 288986 686134
rect 289222 685898 324986 686134
rect 325222 685898 360986 686134
rect 361222 685898 396986 686134
rect 397222 685898 432986 686134
rect 433222 685898 468986 686134
rect 469222 685898 504986 686134
rect 505222 685898 540986 686134
rect 541222 685898 576986 686134
rect 577222 685898 585502 686134
rect 585738 685898 586860 686134
rect -2936 685876 586860 685898
rect -1996 685874 -1396 685876
rect 804 685874 1404 685876
rect 36804 685874 37404 685876
rect 72804 685874 73404 685876
rect 108804 685874 109404 685876
rect 144804 685874 145404 685876
rect 180804 685874 181404 685876
rect 216804 685874 217404 685876
rect 252804 685874 253404 685876
rect 288804 685874 289404 685876
rect 324804 685874 325404 685876
rect 360804 685874 361404 685876
rect 396804 685874 397404 685876
rect 432804 685874 433404 685876
rect 468804 685874 469404 685876
rect 504804 685874 505404 685876
rect 540804 685874 541404 685876
rect 576804 685874 577404 685876
rect 585320 685874 585920 685876
rect -8576 679276 -7976 679278
rect 29604 679276 30204 679278
rect 65604 679276 66204 679278
rect 101604 679276 102204 679278
rect 137604 679276 138204 679278
rect 173604 679276 174204 679278
rect 209604 679276 210204 679278
rect 245604 679276 246204 679278
rect 281604 679276 282204 679278
rect 317604 679276 318204 679278
rect 353604 679276 354204 679278
rect 389604 679276 390204 679278
rect 425604 679276 426204 679278
rect 461604 679276 462204 679278
rect 497604 679276 498204 679278
rect 533604 679276 534204 679278
rect 569604 679276 570204 679278
rect 591900 679276 592500 679278
rect -8576 679254 592500 679276
rect -8576 679018 -8394 679254
rect -8158 679018 29786 679254
rect 30022 679018 65786 679254
rect 66022 679018 101786 679254
rect 102022 679018 137786 679254
rect 138022 679018 173786 679254
rect 174022 679018 209786 679254
rect 210022 679018 245786 679254
rect 246022 679018 281786 679254
rect 282022 679018 317786 679254
rect 318022 679018 353786 679254
rect 354022 679018 389786 679254
rect 390022 679018 425786 679254
rect 426022 679018 461786 679254
rect 462022 679018 497786 679254
rect 498022 679018 533786 679254
rect 534022 679018 569786 679254
rect 570022 679018 592082 679254
rect 592318 679018 592500 679254
rect -8576 678934 592500 679018
rect -8576 678698 -8394 678934
rect -8158 678698 29786 678934
rect 30022 678698 65786 678934
rect 66022 678698 101786 678934
rect 102022 678698 137786 678934
rect 138022 678698 173786 678934
rect 174022 678698 209786 678934
rect 210022 678698 245786 678934
rect 246022 678698 281786 678934
rect 282022 678698 317786 678934
rect 318022 678698 353786 678934
rect 354022 678698 389786 678934
rect 390022 678698 425786 678934
rect 426022 678698 461786 678934
rect 462022 678698 497786 678934
rect 498022 678698 533786 678934
rect 534022 678698 569786 678934
rect 570022 678698 592082 678934
rect 592318 678698 592500 678934
rect -8576 678676 592500 678698
rect -8576 678674 -7976 678676
rect 29604 678674 30204 678676
rect 65604 678674 66204 678676
rect 101604 678674 102204 678676
rect 137604 678674 138204 678676
rect 173604 678674 174204 678676
rect 209604 678674 210204 678676
rect 245604 678674 246204 678676
rect 281604 678674 282204 678676
rect 317604 678674 318204 678676
rect 353604 678674 354204 678676
rect 389604 678674 390204 678676
rect 425604 678674 426204 678676
rect 461604 678674 462204 678676
rect 497604 678674 498204 678676
rect 533604 678674 534204 678676
rect 569604 678674 570204 678676
rect 591900 678674 592500 678676
rect -6696 675676 -6096 675678
rect 26004 675676 26604 675678
rect 62004 675676 62604 675678
rect 98004 675676 98604 675678
rect 134004 675676 134604 675678
rect 170004 675676 170604 675678
rect 206004 675676 206604 675678
rect 242004 675676 242604 675678
rect 278004 675676 278604 675678
rect 314004 675676 314604 675678
rect 350004 675676 350604 675678
rect 386004 675676 386604 675678
rect 422004 675676 422604 675678
rect 458004 675676 458604 675678
rect 494004 675676 494604 675678
rect 530004 675676 530604 675678
rect 566004 675676 566604 675678
rect 590020 675676 590620 675678
rect -6696 675654 590620 675676
rect -6696 675418 -6514 675654
rect -6278 675418 26186 675654
rect 26422 675418 62186 675654
rect 62422 675418 98186 675654
rect 98422 675418 134186 675654
rect 134422 675418 170186 675654
rect 170422 675418 206186 675654
rect 206422 675418 242186 675654
rect 242422 675418 278186 675654
rect 278422 675418 314186 675654
rect 314422 675418 350186 675654
rect 350422 675418 386186 675654
rect 386422 675418 422186 675654
rect 422422 675418 458186 675654
rect 458422 675418 494186 675654
rect 494422 675418 530186 675654
rect 530422 675418 566186 675654
rect 566422 675418 590202 675654
rect 590438 675418 590620 675654
rect -6696 675334 590620 675418
rect -6696 675098 -6514 675334
rect -6278 675098 26186 675334
rect 26422 675098 62186 675334
rect 62422 675098 98186 675334
rect 98422 675098 134186 675334
rect 134422 675098 170186 675334
rect 170422 675098 206186 675334
rect 206422 675098 242186 675334
rect 242422 675098 278186 675334
rect 278422 675098 314186 675334
rect 314422 675098 350186 675334
rect 350422 675098 386186 675334
rect 386422 675098 422186 675334
rect 422422 675098 458186 675334
rect 458422 675098 494186 675334
rect 494422 675098 530186 675334
rect 530422 675098 566186 675334
rect 566422 675098 590202 675334
rect 590438 675098 590620 675334
rect -6696 675076 590620 675098
rect -6696 675074 -6096 675076
rect 26004 675074 26604 675076
rect 62004 675074 62604 675076
rect 98004 675074 98604 675076
rect 134004 675074 134604 675076
rect 170004 675074 170604 675076
rect 206004 675074 206604 675076
rect 242004 675074 242604 675076
rect 278004 675074 278604 675076
rect 314004 675074 314604 675076
rect 350004 675074 350604 675076
rect 386004 675074 386604 675076
rect 422004 675074 422604 675076
rect 458004 675074 458604 675076
rect 494004 675074 494604 675076
rect 530004 675074 530604 675076
rect 566004 675074 566604 675076
rect 590020 675074 590620 675076
rect -4816 672076 -4216 672078
rect 22404 672076 23004 672078
rect 58404 672076 59004 672078
rect 94404 672076 95004 672078
rect 130404 672076 131004 672078
rect 166404 672076 167004 672078
rect 202404 672076 203004 672078
rect 238404 672076 239004 672078
rect 274404 672076 275004 672078
rect 310404 672076 311004 672078
rect 346404 672076 347004 672078
rect 382404 672076 383004 672078
rect 418404 672076 419004 672078
rect 454404 672076 455004 672078
rect 490404 672076 491004 672078
rect 526404 672076 527004 672078
rect 562404 672076 563004 672078
rect 588140 672076 588740 672078
rect -4816 672054 588740 672076
rect -4816 671818 -4634 672054
rect -4398 671818 22586 672054
rect 22822 671818 58586 672054
rect 58822 671818 94586 672054
rect 94822 671818 130586 672054
rect 130822 671818 166586 672054
rect 166822 671818 202586 672054
rect 202822 671818 238586 672054
rect 238822 671818 274586 672054
rect 274822 671818 310586 672054
rect 310822 671818 346586 672054
rect 346822 671818 382586 672054
rect 382822 671818 418586 672054
rect 418822 671818 454586 672054
rect 454822 671818 490586 672054
rect 490822 671818 526586 672054
rect 526822 671818 562586 672054
rect 562822 671818 588322 672054
rect 588558 671818 588740 672054
rect -4816 671734 588740 671818
rect -4816 671498 -4634 671734
rect -4398 671498 22586 671734
rect 22822 671498 58586 671734
rect 58822 671498 94586 671734
rect 94822 671498 130586 671734
rect 130822 671498 166586 671734
rect 166822 671498 202586 671734
rect 202822 671498 238586 671734
rect 238822 671498 274586 671734
rect 274822 671498 310586 671734
rect 310822 671498 346586 671734
rect 346822 671498 382586 671734
rect 382822 671498 418586 671734
rect 418822 671498 454586 671734
rect 454822 671498 490586 671734
rect 490822 671498 526586 671734
rect 526822 671498 562586 671734
rect 562822 671498 588322 671734
rect 588558 671498 588740 671734
rect -4816 671476 588740 671498
rect -4816 671474 -4216 671476
rect 22404 671474 23004 671476
rect 58404 671474 59004 671476
rect 94404 671474 95004 671476
rect 130404 671474 131004 671476
rect 166404 671474 167004 671476
rect 202404 671474 203004 671476
rect 238404 671474 239004 671476
rect 274404 671474 275004 671476
rect 310404 671474 311004 671476
rect 346404 671474 347004 671476
rect 382404 671474 383004 671476
rect 418404 671474 419004 671476
rect 454404 671474 455004 671476
rect 490404 671474 491004 671476
rect 526404 671474 527004 671476
rect 562404 671474 563004 671476
rect 588140 671474 588740 671476
rect -2936 668476 -2336 668478
rect 18804 668476 19404 668478
rect 54804 668476 55404 668478
rect 90804 668476 91404 668478
rect 126804 668476 127404 668478
rect 162804 668476 163404 668478
rect 198804 668476 199404 668478
rect 234804 668476 235404 668478
rect 270804 668476 271404 668478
rect 306804 668476 307404 668478
rect 342804 668476 343404 668478
rect 378804 668476 379404 668478
rect 414804 668476 415404 668478
rect 450804 668476 451404 668478
rect 486804 668476 487404 668478
rect 522804 668476 523404 668478
rect 558804 668476 559404 668478
rect 586260 668476 586860 668478
rect -2936 668454 586860 668476
rect -2936 668218 -2754 668454
rect -2518 668218 18986 668454
rect 19222 668218 54986 668454
rect 55222 668218 90986 668454
rect 91222 668218 126986 668454
rect 127222 668218 162986 668454
rect 163222 668218 198986 668454
rect 199222 668218 234986 668454
rect 235222 668218 270986 668454
rect 271222 668218 306986 668454
rect 307222 668218 342986 668454
rect 343222 668218 378986 668454
rect 379222 668218 414986 668454
rect 415222 668218 450986 668454
rect 451222 668218 486986 668454
rect 487222 668218 522986 668454
rect 523222 668218 558986 668454
rect 559222 668218 586442 668454
rect 586678 668218 586860 668454
rect -2936 668134 586860 668218
rect -2936 667898 -2754 668134
rect -2518 667898 18986 668134
rect 19222 667898 54986 668134
rect 55222 667898 90986 668134
rect 91222 667898 126986 668134
rect 127222 667898 162986 668134
rect 163222 667898 198986 668134
rect 199222 667898 234986 668134
rect 235222 667898 270986 668134
rect 271222 667898 306986 668134
rect 307222 667898 342986 668134
rect 343222 667898 378986 668134
rect 379222 667898 414986 668134
rect 415222 667898 450986 668134
rect 451222 667898 486986 668134
rect 487222 667898 522986 668134
rect 523222 667898 558986 668134
rect 559222 667898 586442 668134
rect 586678 667898 586860 668134
rect -2936 667876 586860 667898
rect -2936 667874 -2336 667876
rect 18804 667874 19404 667876
rect 54804 667874 55404 667876
rect 90804 667874 91404 667876
rect 126804 667874 127404 667876
rect 162804 667874 163404 667876
rect 198804 667874 199404 667876
rect 234804 667874 235404 667876
rect 270804 667874 271404 667876
rect 306804 667874 307404 667876
rect 342804 667874 343404 667876
rect 378804 667874 379404 667876
rect 414804 667874 415404 667876
rect 450804 667874 451404 667876
rect 486804 667874 487404 667876
rect 522804 667874 523404 667876
rect 558804 667874 559404 667876
rect 586260 667874 586860 667876
rect -7636 661276 -7036 661278
rect 11604 661276 12204 661278
rect 47604 661276 48204 661278
rect 83604 661276 84204 661278
rect 119604 661276 120204 661278
rect 155604 661276 156204 661278
rect 191604 661276 192204 661278
rect 227604 661276 228204 661278
rect 263604 661276 264204 661278
rect 299604 661276 300204 661278
rect 335604 661276 336204 661278
rect 371604 661276 372204 661278
rect 407604 661276 408204 661278
rect 443604 661276 444204 661278
rect 479604 661276 480204 661278
rect 515604 661276 516204 661278
rect 551604 661276 552204 661278
rect 590960 661276 591560 661278
rect -8576 661254 592500 661276
rect -8576 661018 -7454 661254
rect -7218 661018 11786 661254
rect 12022 661018 47786 661254
rect 48022 661018 83786 661254
rect 84022 661018 119786 661254
rect 120022 661018 155786 661254
rect 156022 661018 191786 661254
rect 192022 661018 227786 661254
rect 228022 661018 263786 661254
rect 264022 661018 299786 661254
rect 300022 661018 335786 661254
rect 336022 661018 371786 661254
rect 372022 661018 407786 661254
rect 408022 661018 443786 661254
rect 444022 661018 479786 661254
rect 480022 661018 515786 661254
rect 516022 661018 551786 661254
rect 552022 661018 591142 661254
rect 591378 661018 592500 661254
rect -8576 660934 592500 661018
rect -8576 660698 -7454 660934
rect -7218 660698 11786 660934
rect 12022 660698 47786 660934
rect 48022 660698 83786 660934
rect 84022 660698 119786 660934
rect 120022 660698 155786 660934
rect 156022 660698 191786 660934
rect 192022 660698 227786 660934
rect 228022 660698 263786 660934
rect 264022 660698 299786 660934
rect 300022 660698 335786 660934
rect 336022 660698 371786 660934
rect 372022 660698 407786 660934
rect 408022 660698 443786 660934
rect 444022 660698 479786 660934
rect 480022 660698 515786 660934
rect 516022 660698 551786 660934
rect 552022 660698 591142 660934
rect 591378 660698 592500 660934
rect -8576 660676 592500 660698
rect -7636 660674 -7036 660676
rect 11604 660674 12204 660676
rect 47604 660674 48204 660676
rect 83604 660674 84204 660676
rect 119604 660674 120204 660676
rect 155604 660674 156204 660676
rect 191604 660674 192204 660676
rect 227604 660674 228204 660676
rect 263604 660674 264204 660676
rect 299604 660674 300204 660676
rect 335604 660674 336204 660676
rect 371604 660674 372204 660676
rect 407604 660674 408204 660676
rect 443604 660674 444204 660676
rect 479604 660674 480204 660676
rect 515604 660674 516204 660676
rect 551604 660674 552204 660676
rect 590960 660674 591560 660676
rect -5756 657676 -5156 657678
rect 8004 657676 8604 657678
rect 44004 657676 44604 657678
rect 80004 657676 80604 657678
rect 116004 657676 116604 657678
rect 152004 657676 152604 657678
rect 188004 657676 188604 657678
rect 224004 657676 224604 657678
rect 260004 657676 260604 657678
rect 296004 657676 296604 657678
rect 332004 657676 332604 657678
rect 368004 657676 368604 657678
rect 404004 657676 404604 657678
rect 440004 657676 440604 657678
rect 476004 657676 476604 657678
rect 512004 657676 512604 657678
rect 548004 657676 548604 657678
rect 589080 657676 589680 657678
rect -6696 657654 590620 657676
rect -6696 657418 -5574 657654
rect -5338 657418 8186 657654
rect 8422 657418 44186 657654
rect 44422 657418 80186 657654
rect 80422 657418 116186 657654
rect 116422 657418 152186 657654
rect 152422 657418 188186 657654
rect 188422 657418 224186 657654
rect 224422 657418 260186 657654
rect 260422 657418 296186 657654
rect 296422 657418 332186 657654
rect 332422 657418 368186 657654
rect 368422 657418 404186 657654
rect 404422 657418 440186 657654
rect 440422 657418 476186 657654
rect 476422 657418 512186 657654
rect 512422 657418 548186 657654
rect 548422 657418 589262 657654
rect 589498 657418 590620 657654
rect -6696 657334 590620 657418
rect -6696 657098 -5574 657334
rect -5338 657098 8186 657334
rect 8422 657098 44186 657334
rect 44422 657098 80186 657334
rect 80422 657098 116186 657334
rect 116422 657098 152186 657334
rect 152422 657098 188186 657334
rect 188422 657098 224186 657334
rect 224422 657098 260186 657334
rect 260422 657098 296186 657334
rect 296422 657098 332186 657334
rect 332422 657098 368186 657334
rect 368422 657098 404186 657334
rect 404422 657098 440186 657334
rect 440422 657098 476186 657334
rect 476422 657098 512186 657334
rect 512422 657098 548186 657334
rect 548422 657098 589262 657334
rect 589498 657098 590620 657334
rect -6696 657076 590620 657098
rect -5756 657074 -5156 657076
rect 8004 657074 8604 657076
rect 44004 657074 44604 657076
rect 80004 657074 80604 657076
rect 116004 657074 116604 657076
rect 152004 657074 152604 657076
rect 188004 657074 188604 657076
rect 224004 657074 224604 657076
rect 260004 657074 260604 657076
rect 296004 657074 296604 657076
rect 332004 657074 332604 657076
rect 368004 657074 368604 657076
rect 404004 657074 404604 657076
rect 440004 657074 440604 657076
rect 476004 657074 476604 657076
rect 512004 657074 512604 657076
rect 548004 657074 548604 657076
rect 589080 657074 589680 657076
rect -3876 654076 -3276 654078
rect 4404 654076 5004 654078
rect 40404 654076 41004 654078
rect 148404 654076 149004 654078
rect 184404 654076 185004 654078
rect 292404 654076 293004 654078
rect 400404 654076 401004 654078
rect 544404 654076 545004 654078
rect 580404 654076 581004 654078
rect 587200 654076 587800 654078
rect -4816 654054 588740 654076
rect -4816 653818 -3694 654054
rect -3458 653818 4586 654054
rect 4822 653818 40586 654054
rect 40822 653818 148586 654054
rect 148822 653818 184586 654054
rect 184822 653818 292586 654054
rect 292822 653818 400586 654054
rect 400822 653818 544586 654054
rect 544822 653818 580586 654054
rect 580822 653818 587382 654054
rect 587618 653818 588740 654054
rect -4816 653734 588740 653818
rect -4816 653498 -3694 653734
rect -3458 653498 4586 653734
rect 4822 653498 40586 653734
rect 40822 653498 148586 653734
rect 148822 653498 184586 653734
rect 184822 653498 292586 653734
rect 292822 653498 400586 653734
rect 400822 653498 544586 653734
rect 544822 653498 580586 653734
rect 580822 653498 587382 653734
rect 587618 653498 588740 653734
rect -4816 653476 588740 653498
rect -3876 653474 -3276 653476
rect 4404 653474 5004 653476
rect 40404 653474 41004 653476
rect 148404 653474 149004 653476
rect 184404 653474 185004 653476
rect 292404 653474 293004 653476
rect 400404 653474 401004 653476
rect 544404 653474 545004 653476
rect 580404 653474 581004 653476
rect 587200 653474 587800 653476
rect -1996 650476 -1396 650478
rect 804 650476 1404 650478
rect 36804 650476 37404 650478
rect 144804 650476 145404 650478
rect 180804 650476 181404 650478
rect 288804 650476 289404 650478
rect 396804 650476 397404 650478
rect 432804 650476 433404 650478
rect 540804 650476 541404 650478
rect 576804 650476 577404 650478
rect 585320 650476 585920 650478
rect -2936 650454 586860 650476
rect -2936 650218 -1814 650454
rect -1578 650218 986 650454
rect 1222 650218 36986 650454
rect 37222 650218 144986 650454
rect 145222 650218 180986 650454
rect 181222 650218 288986 650454
rect 289222 650218 396986 650454
rect 397222 650218 432986 650454
rect 433222 650218 540986 650454
rect 541222 650218 576986 650454
rect 577222 650218 585502 650454
rect 585738 650218 586860 650454
rect -2936 650134 586860 650218
rect -2936 649898 -1814 650134
rect -1578 649898 986 650134
rect 1222 649898 36986 650134
rect 37222 649898 144986 650134
rect 145222 649898 180986 650134
rect 181222 649898 288986 650134
rect 289222 649898 396986 650134
rect 397222 649898 432986 650134
rect 433222 649898 540986 650134
rect 541222 649898 576986 650134
rect 577222 649898 585502 650134
rect 585738 649898 586860 650134
rect -2936 649876 586860 649898
rect -1996 649874 -1396 649876
rect 804 649874 1404 649876
rect 36804 649874 37404 649876
rect 144804 649874 145404 649876
rect 180804 649874 181404 649876
rect 288804 649874 289404 649876
rect 396804 649874 397404 649876
rect 432804 649874 433404 649876
rect 540804 649874 541404 649876
rect 576804 649874 577404 649876
rect 585320 649874 585920 649876
rect -8576 643276 -7976 643278
rect 29604 643276 30204 643278
rect 136938 643276 137262 643278
rect 173604 643276 174204 643278
rect 266938 643276 267262 643278
rect 281604 643276 282204 643278
rect 386938 643276 387262 643278
rect 425604 643276 426204 643278
rect 516938 643276 517262 643278
rect 533604 643276 534204 643278
rect 569604 643276 570204 643278
rect 591900 643276 592500 643278
rect -8576 643254 592500 643276
rect -8576 643018 -8394 643254
rect -8158 643018 29786 643254
rect 30022 643018 136982 643254
rect 137218 643018 173786 643254
rect 174022 643018 266982 643254
rect 267218 643018 281786 643254
rect 282022 643018 386982 643254
rect 387218 643018 425786 643254
rect 426022 643018 516982 643254
rect 517218 643018 533786 643254
rect 534022 643018 569786 643254
rect 570022 643018 592082 643254
rect 592318 643018 592500 643254
rect -8576 642934 592500 643018
rect -8576 642698 -8394 642934
rect -8158 642698 29786 642934
rect 30022 642698 136982 642934
rect 137218 642698 173786 642934
rect 174022 642698 266982 642934
rect 267218 642698 281786 642934
rect 282022 642698 386982 642934
rect 387218 642698 425786 642934
rect 426022 642698 516982 642934
rect 517218 642698 533786 642934
rect 534022 642698 569786 642934
rect 570022 642698 592082 642934
rect 592318 642698 592500 642934
rect -8576 642676 592500 642698
rect -8576 642674 -7976 642676
rect 29604 642674 30204 642676
rect 136938 642674 137262 642676
rect 173604 642674 174204 642676
rect 266938 642674 267262 642676
rect 281604 642674 282204 642676
rect 386938 642674 387262 642676
rect 425604 642674 426204 642676
rect 516938 642674 517262 642676
rect 533604 642674 534204 642676
rect 569604 642674 570204 642676
rect 591900 642674 592500 642676
rect -6696 639676 -6096 639678
rect 26004 639676 26604 639678
rect 136938 639676 137262 639678
rect 170004 639676 170604 639678
rect 266938 639676 267262 639678
rect 278004 639676 278604 639678
rect 386938 639676 387262 639678
rect 422004 639676 422604 639678
rect 516938 639676 517262 639678
rect 530004 639676 530604 639678
rect 566004 639676 566604 639678
rect 590020 639676 590620 639678
rect -6696 639654 590620 639676
rect -6696 639418 -6514 639654
rect -6278 639418 26186 639654
rect 26422 639418 136982 639654
rect 137218 639418 170186 639654
rect 170422 639418 266982 639654
rect 267218 639418 278186 639654
rect 278422 639418 386982 639654
rect 387218 639418 422186 639654
rect 422422 639418 516982 639654
rect 517218 639418 530186 639654
rect 530422 639418 566186 639654
rect 566422 639418 590202 639654
rect 590438 639418 590620 639654
rect -6696 639334 590620 639418
rect -6696 639098 -6514 639334
rect -6278 639098 26186 639334
rect 26422 639098 136982 639334
rect 137218 639098 170186 639334
rect 170422 639098 266982 639334
rect 267218 639098 278186 639334
rect 278422 639098 386982 639334
rect 387218 639098 422186 639334
rect 422422 639098 516982 639334
rect 517218 639098 530186 639334
rect 530422 639098 566186 639334
rect 566422 639098 590202 639334
rect 590438 639098 590620 639334
rect -6696 639076 590620 639098
rect -6696 639074 -6096 639076
rect 26004 639074 26604 639076
rect 136938 639074 137262 639076
rect 170004 639074 170604 639076
rect 266938 639074 267262 639076
rect 278004 639074 278604 639076
rect 386938 639074 387262 639076
rect 422004 639074 422604 639076
rect 516938 639074 517262 639076
rect 530004 639074 530604 639076
rect 566004 639074 566604 639076
rect 590020 639074 590620 639076
rect -4816 636076 -4216 636078
rect 22404 636076 23004 636078
rect 136938 636076 137262 636078
rect 166404 636076 167004 636078
rect 266938 636076 267262 636078
rect 274404 636076 275004 636078
rect 386938 636076 387262 636078
rect 418404 636076 419004 636078
rect 516938 636076 517262 636078
rect 526404 636076 527004 636078
rect 562404 636076 563004 636078
rect 588140 636076 588740 636078
rect -4816 636054 588740 636076
rect -4816 635818 -4634 636054
rect -4398 635818 22586 636054
rect 22822 635818 136982 636054
rect 137218 635818 166586 636054
rect 166822 635818 266982 636054
rect 267218 635818 274586 636054
rect 274822 635818 386982 636054
rect 387218 635818 418586 636054
rect 418822 635818 516982 636054
rect 517218 635818 526586 636054
rect 526822 635818 562586 636054
rect 562822 635818 588322 636054
rect 588558 635818 588740 636054
rect -4816 635734 588740 635818
rect -4816 635498 -4634 635734
rect -4398 635498 22586 635734
rect 22822 635498 136982 635734
rect 137218 635498 166586 635734
rect 166822 635498 266982 635734
rect 267218 635498 274586 635734
rect 274822 635498 386982 635734
rect 387218 635498 418586 635734
rect 418822 635498 516982 635734
rect 517218 635498 526586 635734
rect 526822 635498 562586 635734
rect 562822 635498 588322 635734
rect 588558 635498 588740 635734
rect -4816 635476 588740 635498
rect -4816 635474 -4216 635476
rect 22404 635474 23004 635476
rect 136938 635474 137262 635476
rect 166404 635474 167004 635476
rect 266938 635474 267262 635476
rect 274404 635474 275004 635476
rect 386938 635474 387262 635476
rect 418404 635474 419004 635476
rect 516938 635474 517262 635476
rect 526404 635474 527004 635476
rect 562404 635474 563004 635476
rect 588140 635474 588740 635476
rect -2936 632476 -2336 632478
rect 18804 632476 19404 632478
rect 54804 632476 55404 632478
rect 136938 632476 137262 632478
rect 162804 632476 163404 632478
rect 266938 632476 267262 632478
rect 270804 632476 271404 632478
rect 386938 632476 387262 632478
rect 414804 632476 415404 632478
rect 516938 632476 517262 632478
rect 522804 632476 523404 632478
rect 558804 632476 559404 632478
rect 586260 632476 586860 632478
rect -2936 632454 586860 632476
rect -2936 632218 -2754 632454
rect -2518 632218 18986 632454
rect 19222 632218 54986 632454
rect 55222 632218 136982 632454
rect 137218 632218 162986 632454
rect 163222 632218 266982 632454
rect 267218 632218 270986 632454
rect 271222 632218 386982 632454
rect 387218 632218 414986 632454
rect 415222 632218 516982 632454
rect 517218 632218 522986 632454
rect 523222 632218 558986 632454
rect 559222 632218 586442 632454
rect 586678 632218 586860 632454
rect -2936 632134 586860 632218
rect -2936 631898 -2754 632134
rect -2518 631898 18986 632134
rect 19222 631898 54986 632134
rect 55222 631898 136982 632134
rect 137218 631898 162986 632134
rect 163222 631898 266982 632134
rect 267218 631898 270986 632134
rect 271222 631898 386982 632134
rect 387218 631898 414986 632134
rect 415222 631898 516982 632134
rect 517218 631898 522986 632134
rect 523222 631898 558986 632134
rect 559222 631898 586442 632134
rect 586678 631898 586860 632134
rect -2936 631876 586860 631898
rect -2936 631874 -2336 631876
rect 18804 631874 19404 631876
rect 54804 631874 55404 631876
rect 136938 631874 137262 631876
rect 162804 631874 163404 631876
rect 266938 631874 267262 631876
rect 270804 631874 271404 631876
rect 386938 631874 387262 631876
rect 414804 631874 415404 631876
rect 516938 631874 517262 631876
rect 522804 631874 523404 631876
rect 558804 631874 559404 631876
rect 586260 631874 586860 631876
rect -7636 625276 -7036 625278
rect 11604 625276 12204 625278
rect 47604 625276 48204 625278
rect 136494 625276 136814 625278
rect 155604 625276 156204 625278
rect 266494 625276 266814 625278
rect 299604 625276 300204 625278
rect 386494 625276 386814 625278
rect 407604 625276 408204 625278
rect 516494 625276 516814 625278
rect 551604 625276 552204 625278
rect 590960 625276 591560 625278
rect -8576 625254 592500 625276
rect -8576 625018 -7454 625254
rect -7218 625018 11786 625254
rect 12022 625018 47786 625254
rect 48022 625018 136536 625254
rect 136772 625018 155786 625254
rect 156022 625018 266536 625254
rect 266772 625018 299786 625254
rect 300022 625018 386536 625254
rect 386772 625018 407786 625254
rect 408022 625018 516536 625254
rect 516772 625018 551786 625254
rect 552022 625018 591142 625254
rect 591378 625018 592500 625254
rect -8576 624934 592500 625018
rect -8576 624698 -7454 624934
rect -7218 624698 11786 624934
rect 12022 624698 47786 624934
rect 48022 624698 136536 624934
rect 136772 624698 155786 624934
rect 156022 624698 266536 624934
rect 266772 624698 299786 624934
rect 300022 624698 386536 624934
rect 386772 624698 407786 624934
rect 408022 624698 516536 624934
rect 516772 624698 551786 624934
rect 552022 624698 591142 624934
rect 591378 624698 592500 624934
rect -8576 624676 592500 624698
rect -7636 624674 -7036 624676
rect 11604 624674 12204 624676
rect 47604 624674 48204 624676
rect 136494 624674 136814 624676
rect 155604 624674 156204 624676
rect 266494 624674 266814 624676
rect 299604 624674 300204 624676
rect 386494 624674 386814 624676
rect 407604 624674 408204 624676
rect 516494 624674 516814 624676
rect 551604 624674 552204 624676
rect 590960 624674 591560 624676
rect -5756 621676 -5156 621678
rect 8004 621676 8604 621678
rect 44004 621676 44604 621678
rect 136494 621676 136814 621678
rect 152004 621676 152604 621678
rect 266494 621676 266814 621678
rect 296004 621676 296604 621678
rect 386494 621676 386814 621678
rect 404004 621676 404604 621678
rect 516494 621676 516814 621678
rect 548004 621676 548604 621678
rect 589080 621676 589680 621678
rect -6696 621654 590620 621676
rect -6696 621418 -5574 621654
rect -5338 621418 8186 621654
rect 8422 621418 44186 621654
rect 44422 621418 136536 621654
rect 136772 621418 152186 621654
rect 152422 621418 266536 621654
rect 266772 621418 296186 621654
rect 296422 621418 386536 621654
rect 386772 621418 404186 621654
rect 404422 621418 516536 621654
rect 516772 621418 548186 621654
rect 548422 621418 589262 621654
rect 589498 621418 590620 621654
rect -6696 621334 590620 621418
rect -6696 621098 -5574 621334
rect -5338 621098 8186 621334
rect 8422 621098 44186 621334
rect 44422 621098 136536 621334
rect 136772 621098 152186 621334
rect 152422 621098 266536 621334
rect 266772 621098 296186 621334
rect 296422 621098 386536 621334
rect 386772 621098 404186 621334
rect 404422 621098 516536 621334
rect 516772 621098 548186 621334
rect 548422 621098 589262 621334
rect 589498 621098 590620 621334
rect -6696 621076 590620 621098
rect -5756 621074 -5156 621076
rect 8004 621074 8604 621076
rect 44004 621074 44604 621076
rect 136494 621074 136814 621076
rect 152004 621074 152604 621076
rect 266494 621074 266814 621076
rect 296004 621074 296604 621076
rect 386494 621074 386814 621076
rect 404004 621074 404604 621076
rect 516494 621074 516814 621076
rect 548004 621074 548604 621076
rect 589080 621074 589680 621076
rect -3876 618076 -3276 618078
rect 4404 618076 5004 618078
rect 40404 618076 41004 618078
rect 136494 618076 136814 618078
rect 148404 618076 149004 618078
rect 184404 618076 185004 618078
rect 266494 618076 266814 618078
rect 292404 618076 293004 618078
rect 386494 618076 386814 618078
rect 400404 618076 401004 618078
rect 516494 618076 516814 618078
rect 544404 618076 545004 618078
rect 580404 618076 581004 618078
rect 587200 618076 587800 618078
rect -4816 618054 588740 618076
rect -4816 617818 -3694 618054
rect -3458 617818 4586 618054
rect 4822 617818 40586 618054
rect 40822 617818 136536 618054
rect 136772 617818 148586 618054
rect 148822 617818 184586 618054
rect 184822 617818 266536 618054
rect 266772 617818 292586 618054
rect 292822 617818 386536 618054
rect 386772 617818 400586 618054
rect 400822 617818 516536 618054
rect 516772 617818 544586 618054
rect 544822 617818 580586 618054
rect 580822 617818 587382 618054
rect 587618 617818 588740 618054
rect -4816 617734 588740 617818
rect -4816 617498 -3694 617734
rect -3458 617498 4586 617734
rect 4822 617498 40586 617734
rect 40822 617498 136536 617734
rect 136772 617498 148586 617734
rect 148822 617498 184586 617734
rect 184822 617498 266536 617734
rect 266772 617498 292586 617734
rect 292822 617498 386536 617734
rect 386772 617498 400586 617734
rect 400822 617498 516536 617734
rect 516772 617498 544586 617734
rect 544822 617498 580586 617734
rect 580822 617498 587382 617734
rect 587618 617498 588740 617734
rect -4816 617476 588740 617498
rect -3876 617474 -3276 617476
rect 4404 617474 5004 617476
rect 40404 617474 41004 617476
rect 136494 617474 136814 617476
rect 148404 617474 149004 617476
rect 184404 617474 185004 617476
rect 266494 617474 266814 617476
rect 292404 617474 293004 617476
rect 386494 617474 386814 617476
rect 400404 617474 401004 617476
rect 516494 617474 516814 617476
rect 544404 617474 545004 617476
rect 580404 617474 581004 617476
rect 587200 617474 587800 617476
rect -1996 614476 -1396 614478
rect 804 614476 1404 614478
rect 36804 614476 37404 614478
rect 136494 614476 136814 614478
rect 144804 614476 145404 614478
rect 180804 614476 181404 614478
rect 266494 614476 266814 614478
rect 288804 614476 289404 614478
rect 386494 614476 386814 614478
rect 396804 614476 397404 614478
rect 432804 614476 433404 614478
rect 516494 614476 516814 614478
rect 540804 614476 541404 614478
rect 576804 614476 577404 614478
rect 585320 614476 585920 614478
rect -2936 614454 586860 614476
rect -2936 614218 -1814 614454
rect -1578 614218 986 614454
rect 1222 614218 36986 614454
rect 37222 614218 136536 614454
rect 136772 614218 144986 614454
rect 145222 614218 180986 614454
rect 181222 614218 266536 614454
rect 266772 614218 288986 614454
rect 289222 614218 386536 614454
rect 386772 614218 396986 614454
rect 397222 614218 432986 614454
rect 433222 614218 516536 614454
rect 516772 614218 540986 614454
rect 541222 614218 576986 614454
rect 577222 614218 585502 614454
rect 585738 614218 586860 614454
rect -2936 614134 586860 614218
rect -2936 613898 -1814 614134
rect -1578 613898 986 614134
rect 1222 613898 36986 614134
rect 37222 613898 136536 614134
rect 136772 613898 144986 614134
rect 145222 613898 180986 614134
rect 181222 613898 266536 614134
rect 266772 613898 288986 614134
rect 289222 613898 386536 614134
rect 386772 613898 396986 614134
rect 397222 613898 432986 614134
rect 433222 613898 516536 614134
rect 516772 613898 540986 614134
rect 541222 613898 576986 614134
rect 577222 613898 585502 614134
rect 585738 613898 586860 614134
rect -2936 613876 586860 613898
rect -1996 613874 -1396 613876
rect 804 613874 1404 613876
rect 36804 613874 37404 613876
rect 136494 613874 136814 613876
rect 144804 613874 145404 613876
rect 180804 613874 181404 613876
rect 266494 613874 266814 613876
rect 288804 613874 289404 613876
rect 386494 613874 386814 613876
rect 396804 613874 397404 613876
rect 432804 613874 433404 613876
rect 516494 613874 516814 613876
rect 540804 613874 541404 613876
rect 576804 613874 577404 613876
rect 585320 613874 585920 613876
rect -8576 607276 -7976 607278
rect 29604 607276 30204 607278
rect 136938 607276 137262 607278
rect 173604 607276 174204 607278
rect 266938 607276 267262 607278
rect 281604 607276 282204 607278
rect 386938 607276 387262 607278
rect 425604 607276 426204 607278
rect 516938 607276 517262 607278
rect 533604 607276 534204 607278
rect 569604 607276 570204 607278
rect 591900 607276 592500 607278
rect -8576 607254 592500 607276
rect -8576 607018 -8394 607254
rect -8158 607018 29786 607254
rect 30022 607018 136982 607254
rect 137218 607018 173786 607254
rect 174022 607018 266982 607254
rect 267218 607018 281786 607254
rect 282022 607018 386982 607254
rect 387218 607018 425786 607254
rect 426022 607018 516982 607254
rect 517218 607018 533786 607254
rect 534022 607018 569786 607254
rect 570022 607018 592082 607254
rect 592318 607018 592500 607254
rect -8576 606934 592500 607018
rect -8576 606698 -8394 606934
rect -8158 606698 29786 606934
rect 30022 606698 136982 606934
rect 137218 606698 173786 606934
rect 174022 606698 266982 606934
rect 267218 606698 281786 606934
rect 282022 606698 386982 606934
rect 387218 606698 425786 606934
rect 426022 606698 516982 606934
rect 517218 606698 533786 606934
rect 534022 606698 569786 606934
rect 570022 606698 592082 606934
rect 592318 606698 592500 606934
rect -8576 606676 592500 606698
rect -8576 606674 -7976 606676
rect 29604 606674 30204 606676
rect 136938 606674 137262 606676
rect 173604 606674 174204 606676
rect 266938 606674 267262 606676
rect 281604 606674 282204 606676
rect 386938 606674 387262 606676
rect 425604 606674 426204 606676
rect 516938 606674 517262 606676
rect 533604 606674 534204 606676
rect 569604 606674 570204 606676
rect 591900 606674 592500 606676
rect -6696 603676 -6096 603678
rect 26004 603676 26604 603678
rect 136938 603676 137262 603678
rect 170004 603676 170604 603678
rect 266938 603676 267262 603678
rect 278004 603676 278604 603678
rect 386938 603676 387262 603678
rect 422004 603676 422604 603678
rect 516938 603676 517262 603678
rect 530004 603676 530604 603678
rect 566004 603676 566604 603678
rect 590020 603676 590620 603678
rect -6696 603654 590620 603676
rect -6696 603418 -6514 603654
rect -6278 603418 26186 603654
rect 26422 603418 136982 603654
rect 137218 603418 170186 603654
rect 170422 603418 266982 603654
rect 267218 603418 278186 603654
rect 278422 603418 386982 603654
rect 387218 603418 422186 603654
rect 422422 603418 516982 603654
rect 517218 603418 530186 603654
rect 530422 603418 566186 603654
rect 566422 603418 590202 603654
rect 590438 603418 590620 603654
rect -6696 603334 590620 603418
rect -6696 603098 -6514 603334
rect -6278 603098 26186 603334
rect 26422 603098 136982 603334
rect 137218 603098 170186 603334
rect 170422 603098 266982 603334
rect 267218 603098 278186 603334
rect 278422 603098 386982 603334
rect 387218 603098 422186 603334
rect 422422 603098 516982 603334
rect 517218 603098 530186 603334
rect 530422 603098 566186 603334
rect 566422 603098 590202 603334
rect 590438 603098 590620 603334
rect -6696 603076 590620 603098
rect -6696 603074 -6096 603076
rect 26004 603074 26604 603076
rect 136938 603074 137262 603076
rect 170004 603074 170604 603076
rect 266938 603074 267262 603076
rect 278004 603074 278604 603076
rect 386938 603074 387262 603076
rect 422004 603074 422604 603076
rect 516938 603074 517262 603076
rect 530004 603074 530604 603076
rect 566004 603074 566604 603076
rect 590020 603074 590620 603076
rect -4816 600076 -4216 600078
rect 22404 600076 23004 600078
rect 136938 600076 137262 600078
rect 166404 600076 167004 600078
rect 266938 600076 267262 600078
rect 274404 600076 275004 600078
rect 386938 600076 387262 600078
rect 418404 600076 419004 600078
rect 516938 600076 517262 600078
rect 526404 600076 527004 600078
rect 562404 600076 563004 600078
rect 588140 600076 588740 600078
rect -4816 600054 588740 600076
rect -4816 599818 -4634 600054
rect -4398 599818 22586 600054
rect 22822 599818 136982 600054
rect 137218 599818 166586 600054
rect 166822 599818 266982 600054
rect 267218 599818 274586 600054
rect 274822 599818 386982 600054
rect 387218 599818 418586 600054
rect 418822 599818 516982 600054
rect 517218 599818 526586 600054
rect 526822 599818 562586 600054
rect 562822 599818 588322 600054
rect 588558 599818 588740 600054
rect -4816 599734 588740 599818
rect -4816 599498 -4634 599734
rect -4398 599498 22586 599734
rect 22822 599498 136982 599734
rect 137218 599498 166586 599734
rect 166822 599498 266982 599734
rect 267218 599498 274586 599734
rect 274822 599498 386982 599734
rect 387218 599498 418586 599734
rect 418822 599498 516982 599734
rect 517218 599498 526586 599734
rect 526822 599498 562586 599734
rect 562822 599498 588322 599734
rect 588558 599498 588740 599734
rect -4816 599476 588740 599498
rect -4816 599474 -4216 599476
rect 22404 599474 23004 599476
rect 136938 599474 137262 599476
rect 166404 599474 167004 599476
rect 266938 599474 267262 599476
rect 274404 599474 275004 599476
rect 386938 599474 387262 599476
rect 418404 599474 419004 599476
rect 516938 599474 517262 599476
rect 526404 599474 527004 599476
rect 562404 599474 563004 599476
rect 588140 599474 588740 599476
rect -2936 596476 -2336 596478
rect 18804 596476 19404 596478
rect 54804 596476 55404 596478
rect 136938 596476 137262 596478
rect 162804 596476 163404 596478
rect 266938 596476 267262 596478
rect 270804 596476 271404 596478
rect 386938 596476 387262 596478
rect 414804 596476 415404 596478
rect 516938 596476 517262 596478
rect 522804 596476 523404 596478
rect 558804 596476 559404 596478
rect 586260 596476 586860 596478
rect -2936 596454 586860 596476
rect -2936 596218 -2754 596454
rect -2518 596218 18986 596454
rect 19222 596218 54986 596454
rect 55222 596218 136982 596454
rect 137218 596218 162986 596454
rect 163222 596218 266982 596454
rect 267218 596218 270986 596454
rect 271222 596218 386982 596454
rect 387218 596218 414986 596454
rect 415222 596218 516982 596454
rect 517218 596218 522986 596454
rect 523222 596218 558986 596454
rect 559222 596218 586442 596454
rect 586678 596218 586860 596454
rect -2936 596134 586860 596218
rect -2936 595898 -2754 596134
rect -2518 595898 18986 596134
rect 19222 595898 54986 596134
rect 55222 595898 136982 596134
rect 137218 595898 162986 596134
rect 163222 595898 266982 596134
rect 267218 595898 270986 596134
rect 271222 595898 386982 596134
rect 387218 595898 414986 596134
rect 415222 595898 516982 596134
rect 517218 595898 522986 596134
rect 523222 595898 558986 596134
rect 559222 595898 586442 596134
rect 586678 595898 586860 596134
rect -2936 595876 586860 595898
rect -2936 595874 -2336 595876
rect 18804 595874 19404 595876
rect 54804 595874 55404 595876
rect 136938 595874 137262 595876
rect 162804 595874 163404 595876
rect 266938 595874 267262 595876
rect 270804 595874 271404 595876
rect 386938 595874 387262 595876
rect 414804 595874 415404 595876
rect 516938 595874 517262 595876
rect 522804 595874 523404 595876
rect 558804 595874 559404 595876
rect 586260 595874 586860 595876
rect -7636 589276 -7036 589278
rect 11604 589276 12204 589278
rect 47604 589276 48204 589278
rect 136494 589276 136814 589278
rect 155604 589276 156204 589278
rect 266494 589276 266814 589278
rect 299604 589276 300204 589278
rect 386494 589276 386814 589278
rect 407604 589276 408204 589278
rect 516494 589276 516814 589278
rect 551604 589276 552204 589278
rect 590960 589276 591560 589278
rect -8576 589254 592500 589276
rect -8576 589018 -7454 589254
rect -7218 589018 11786 589254
rect 12022 589018 47786 589254
rect 48022 589018 136536 589254
rect 136772 589018 155786 589254
rect 156022 589018 266536 589254
rect 266772 589018 299786 589254
rect 300022 589018 386536 589254
rect 386772 589018 407786 589254
rect 408022 589018 516536 589254
rect 516772 589018 551786 589254
rect 552022 589018 591142 589254
rect 591378 589018 592500 589254
rect -8576 588934 592500 589018
rect -8576 588698 -7454 588934
rect -7218 588698 11786 588934
rect 12022 588698 47786 588934
rect 48022 588698 136536 588934
rect 136772 588698 155786 588934
rect 156022 588698 266536 588934
rect 266772 588698 299786 588934
rect 300022 588698 386536 588934
rect 386772 588698 407786 588934
rect 408022 588698 516536 588934
rect 516772 588698 551786 588934
rect 552022 588698 591142 588934
rect 591378 588698 592500 588934
rect -8576 588676 592500 588698
rect -7636 588674 -7036 588676
rect 11604 588674 12204 588676
rect 47604 588674 48204 588676
rect 136494 588674 136814 588676
rect 155604 588674 156204 588676
rect 266494 588674 266814 588676
rect 299604 588674 300204 588676
rect 386494 588674 386814 588676
rect 407604 588674 408204 588676
rect 516494 588674 516814 588676
rect 551604 588674 552204 588676
rect 590960 588674 591560 588676
rect 270228 587298 387756 587340
rect 270228 587062 270270 587298
rect 270506 587062 387478 587298
rect 387714 587062 387756 587298
rect 270228 587020 387756 587062
rect -5756 585676 -5156 585678
rect 8004 585676 8604 585678
rect 44004 585676 44604 585678
rect 136494 585676 136814 585678
rect 152004 585676 152604 585678
rect 266494 585676 266814 585678
rect 296004 585676 296604 585678
rect 386494 585676 386814 585678
rect 404004 585676 404604 585678
rect 516494 585676 516814 585678
rect 548004 585676 548604 585678
rect 589080 585676 589680 585678
rect -6696 585654 590620 585676
rect -6696 585418 -5574 585654
rect -5338 585418 8186 585654
rect 8422 585418 44186 585654
rect 44422 585418 136536 585654
rect 136772 585418 152186 585654
rect 152422 585418 266536 585654
rect 266772 585418 296186 585654
rect 296422 585418 386536 585654
rect 386772 585418 404186 585654
rect 404422 585418 516536 585654
rect 516772 585418 548186 585654
rect 548422 585418 589262 585654
rect 589498 585418 590620 585654
rect -6696 585334 590620 585418
rect -6696 585098 -5574 585334
rect -5338 585098 8186 585334
rect 8422 585098 44186 585334
rect 44422 585098 136536 585334
rect 136772 585098 152186 585334
rect 152422 585098 266536 585334
rect 266772 585098 296186 585334
rect 296422 585098 386536 585334
rect 386772 585098 404186 585334
rect 404422 585098 516536 585334
rect 516772 585098 548186 585334
rect 548422 585098 589262 585334
rect 589498 585098 590620 585334
rect -6696 585076 590620 585098
rect -5756 585074 -5156 585076
rect 8004 585074 8604 585076
rect 44004 585074 44604 585076
rect 136494 585074 136814 585076
rect 152004 585074 152604 585076
rect 266494 585074 266814 585076
rect 296004 585074 296604 585076
rect 386494 585074 386814 585076
rect 404004 585074 404604 585076
rect 516494 585074 516814 585076
rect 548004 585074 548604 585076
rect 589080 585074 589680 585076
rect -3876 582076 -3276 582078
rect 4404 582076 5004 582078
rect 40404 582076 41004 582078
rect 136494 582076 136814 582078
rect 148404 582076 149004 582078
rect 184404 582076 185004 582078
rect 266494 582076 266814 582078
rect 292404 582076 293004 582078
rect 386494 582076 386814 582078
rect 400404 582076 401004 582078
rect 516494 582076 516814 582078
rect 544404 582076 545004 582078
rect 580404 582076 581004 582078
rect 587200 582076 587800 582078
rect -4816 582054 588740 582076
rect -4816 581818 -3694 582054
rect -3458 581818 4586 582054
rect 4822 581818 40586 582054
rect 40822 581818 136536 582054
rect 136772 581818 148586 582054
rect 148822 581818 184586 582054
rect 184822 581818 266536 582054
rect 266772 581818 292586 582054
rect 292822 581818 386536 582054
rect 386772 581818 400586 582054
rect 400822 581818 516536 582054
rect 516772 581818 544586 582054
rect 544822 581818 580586 582054
rect 580822 581818 587382 582054
rect 587618 581818 588740 582054
rect -4816 581734 588740 581818
rect -4816 581498 -3694 581734
rect -3458 581498 4586 581734
rect 4822 581498 40586 581734
rect 40822 581498 136536 581734
rect 136772 581498 148586 581734
rect 148822 581498 184586 581734
rect 184822 581498 266536 581734
rect 266772 581498 292586 581734
rect 292822 581498 386536 581734
rect 386772 581498 400586 581734
rect 400822 581498 516536 581734
rect 516772 581498 544586 581734
rect 544822 581498 580586 581734
rect 580822 581498 587382 581734
rect 587618 581498 588740 581734
rect -4816 581476 588740 581498
rect -3876 581474 -3276 581476
rect 4404 581474 5004 581476
rect 40404 581474 41004 581476
rect 136494 581474 136814 581476
rect 148404 581474 149004 581476
rect 184404 581474 185004 581476
rect 266494 581474 266814 581476
rect 292404 581474 293004 581476
rect 386494 581474 386814 581476
rect 400404 581474 401004 581476
rect 516494 581474 516814 581476
rect 544404 581474 545004 581476
rect 580404 581474 581004 581476
rect 587200 581474 587800 581476
rect 389092 579818 519132 579860
rect 389092 579582 389134 579818
rect 389370 579582 518854 579818
rect 519090 579582 519132 579818
rect 389092 579540 519132 579582
rect 60468 579138 437620 579180
rect 60468 578902 60510 579138
rect 60746 578902 188758 579138
rect 188994 578902 282414 579138
rect 282650 578902 310198 579138
rect 310434 578902 437342 579138
rect 437578 578902 437620 579138
rect 60468 578860 437620 578902
rect -1996 578476 -1396 578478
rect 804 578476 1404 578478
rect 36804 578476 37404 578478
rect 136494 578476 136814 578478
rect 144804 578476 145404 578478
rect 180804 578476 181404 578478
rect 266494 578476 266814 578478
rect 288804 578476 289404 578478
rect 386494 578476 386814 578478
rect 396804 578476 397404 578478
rect 432804 578476 433404 578478
rect 516494 578476 516814 578478
rect 540804 578476 541404 578478
rect 576804 578476 577404 578478
rect 585320 578476 585920 578478
rect -2936 578454 586860 578476
rect -2936 578218 -1814 578454
rect -1578 578218 986 578454
rect 1222 578218 36986 578454
rect 37222 578218 136536 578454
rect 136772 578218 144986 578454
rect 145222 578218 180986 578454
rect 181222 578218 266536 578454
rect 266772 578218 288986 578454
rect 289222 578218 386536 578454
rect 386772 578218 396986 578454
rect 397222 578218 432986 578454
rect 433222 578218 516536 578454
rect 516772 578218 540986 578454
rect 541222 578218 576986 578454
rect 577222 578218 585502 578454
rect 585738 578218 586860 578454
rect -2936 578134 586860 578218
rect -2936 577898 -1814 578134
rect -1578 577898 986 578134
rect 1222 577898 36986 578134
rect 37222 577898 136536 578134
rect 136772 577898 144986 578134
rect 145222 577898 180986 578134
rect 181222 577898 266536 578134
rect 266772 577898 288986 578134
rect 289222 577898 386536 578134
rect 386772 577898 396986 578134
rect 397222 577898 432986 578134
rect 433222 577898 516536 578134
rect 516772 577898 540986 578134
rect 541222 577898 576986 578134
rect 577222 577898 585502 578134
rect 585738 577898 586860 578134
rect -2936 577876 586860 577898
rect -1996 577874 -1396 577876
rect 804 577874 1404 577876
rect 36804 577874 37404 577876
rect 136494 577874 136814 577876
rect 144804 577874 145404 577876
rect 180804 577874 181404 577876
rect 266494 577874 266814 577876
rect 288804 577874 289404 577876
rect 386494 577874 386814 577876
rect 396804 577874 397404 577876
rect 432804 577874 433404 577876
rect 516494 577874 516814 577876
rect 540804 577874 541404 577876
rect 576804 577874 577404 577876
rect 585320 577874 585920 577876
rect -8576 571276 -7976 571278
rect 29604 571276 30204 571278
rect 136938 571276 137262 571278
rect 173604 571276 174204 571278
rect 266938 571276 267262 571278
rect 281604 571276 282204 571278
rect 386938 571276 387262 571278
rect 425604 571276 426204 571278
rect 516938 571276 517262 571278
rect 533604 571276 534204 571278
rect 569604 571276 570204 571278
rect 591900 571276 592500 571278
rect -8576 571254 592500 571276
rect -8576 571018 -8394 571254
rect -8158 571018 29786 571254
rect 30022 571018 136982 571254
rect 137218 571018 173786 571254
rect 174022 571018 266982 571254
rect 267218 571018 281786 571254
rect 282022 571018 386982 571254
rect 387218 571018 425786 571254
rect 426022 571018 516982 571254
rect 517218 571018 533786 571254
rect 534022 571018 569786 571254
rect 570022 571018 592082 571254
rect 592318 571018 592500 571254
rect -8576 570934 592500 571018
rect -8576 570698 -8394 570934
rect -8158 570698 29786 570934
rect 30022 570698 136982 570934
rect 137218 570698 173786 570934
rect 174022 570698 266982 570934
rect 267218 570698 281786 570934
rect 282022 570698 386982 570934
rect 387218 570698 425786 570934
rect 426022 570698 516982 570934
rect 517218 570698 533786 570934
rect 534022 570698 569786 570934
rect 570022 570698 592082 570934
rect 592318 570698 592500 570934
rect -8576 570676 592500 570698
rect -8576 570674 -7976 570676
rect 29604 570674 30204 570676
rect 136938 570674 137262 570676
rect 173604 570674 174204 570676
rect 266938 570674 267262 570676
rect 281604 570674 282204 570676
rect 386938 570674 387262 570676
rect 425604 570674 426204 570676
rect 516938 570674 517262 570676
rect 533604 570674 534204 570676
rect 569604 570674 570204 570676
rect 591900 570674 592500 570676
rect -6696 567676 -6096 567678
rect 26004 567676 26604 567678
rect 136938 567676 137262 567678
rect 170004 567676 170604 567678
rect 266938 567676 267262 567678
rect 278004 567676 278604 567678
rect 386938 567676 387262 567678
rect 422004 567676 422604 567678
rect 516938 567676 517262 567678
rect 530004 567676 530604 567678
rect 566004 567676 566604 567678
rect 590020 567676 590620 567678
rect -6696 567654 590620 567676
rect -6696 567418 -6514 567654
rect -6278 567418 26186 567654
rect 26422 567418 136982 567654
rect 137218 567418 170186 567654
rect 170422 567418 266982 567654
rect 267218 567418 278186 567654
rect 278422 567418 386982 567654
rect 387218 567418 422186 567654
rect 422422 567418 516982 567654
rect 517218 567418 530186 567654
rect 530422 567418 566186 567654
rect 566422 567418 590202 567654
rect 590438 567418 590620 567654
rect -6696 567334 590620 567418
rect -6696 567098 -6514 567334
rect -6278 567098 26186 567334
rect 26422 567098 136982 567334
rect 137218 567098 170186 567334
rect 170422 567098 266982 567334
rect 267218 567098 278186 567334
rect 278422 567098 386982 567334
rect 387218 567098 422186 567334
rect 422422 567098 516982 567334
rect 517218 567098 530186 567334
rect 530422 567098 566186 567334
rect 566422 567098 590202 567334
rect 590438 567098 590620 567334
rect -6696 567076 590620 567098
rect -6696 567074 -6096 567076
rect 26004 567074 26604 567076
rect 136938 567074 137262 567076
rect 170004 567074 170604 567076
rect 266938 567074 267262 567076
rect 278004 567074 278604 567076
rect 386938 567074 387262 567076
rect 422004 567074 422604 567076
rect 516938 567074 517262 567076
rect 530004 567074 530604 567076
rect 566004 567074 566604 567076
rect 590020 567074 590620 567076
rect -4816 564076 -4216 564078
rect 22404 564076 23004 564078
rect 136938 564076 137262 564078
rect 166404 564076 167004 564078
rect 266938 564076 267262 564078
rect 274404 564076 275004 564078
rect 386938 564076 387262 564078
rect 418404 564076 419004 564078
rect 516938 564076 517262 564078
rect 526404 564076 527004 564078
rect 562404 564076 563004 564078
rect 588140 564076 588740 564078
rect -4816 564054 588740 564076
rect -4816 563818 -4634 564054
rect -4398 563818 22586 564054
rect 22822 563818 136982 564054
rect 137218 563818 166586 564054
rect 166822 563818 266982 564054
rect 267218 563818 274586 564054
rect 274822 563818 386982 564054
rect 387218 563818 418586 564054
rect 418822 563818 516982 564054
rect 517218 563818 526586 564054
rect 526822 563818 562586 564054
rect 562822 563818 588322 564054
rect 588558 563818 588740 564054
rect -4816 563734 588740 563818
rect -4816 563498 -4634 563734
rect -4398 563498 22586 563734
rect 22822 563498 136982 563734
rect 137218 563498 166586 563734
rect 166822 563498 266982 563734
rect 267218 563498 274586 563734
rect 274822 563498 386982 563734
rect 387218 563498 418586 563734
rect 418822 563498 516982 563734
rect 517218 563498 526586 563734
rect 526822 563498 562586 563734
rect 562822 563498 588322 563734
rect 588558 563498 588740 563734
rect -4816 563476 588740 563498
rect -4816 563474 -4216 563476
rect 22404 563474 23004 563476
rect 136938 563474 137262 563476
rect 166404 563474 167004 563476
rect 266938 563474 267262 563476
rect 274404 563474 275004 563476
rect 386938 563474 387262 563476
rect 418404 563474 419004 563476
rect 516938 563474 517262 563476
rect 526404 563474 527004 563476
rect 562404 563474 563004 563476
rect 588140 563474 588740 563476
rect -2936 560476 -2336 560478
rect 18804 560476 19404 560478
rect 54804 560476 55404 560478
rect 162804 560476 163404 560478
rect 270804 560476 271404 560478
rect 414804 560476 415404 560478
rect 522804 560476 523404 560478
rect 558804 560476 559404 560478
rect 586260 560476 586860 560478
rect -2936 560454 586860 560476
rect -2936 560218 -2754 560454
rect -2518 560218 18986 560454
rect 19222 560218 54986 560454
rect 55222 560218 162986 560454
rect 163222 560218 270986 560454
rect 271222 560218 414986 560454
rect 415222 560218 522986 560454
rect 523222 560218 558986 560454
rect 559222 560218 586442 560454
rect 586678 560218 586860 560454
rect -2936 560134 586860 560218
rect -2936 559898 -2754 560134
rect -2518 559898 18986 560134
rect 19222 559898 54986 560134
rect 55222 559898 162986 560134
rect 163222 559898 270986 560134
rect 271222 559898 414986 560134
rect 415222 559898 522986 560134
rect 523222 559898 558986 560134
rect 559222 559898 586442 560134
rect 586678 559898 586860 560134
rect -2936 559876 586860 559898
rect -2936 559874 -2336 559876
rect 18804 559874 19404 559876
rect 54804 559874 55404 559876
rect 162804 559874 163404 559876
rect 270804 559874 271404 559876
rect 414804 559874 415404 559876
rect 522804 559874 523404 559876
rect 558804 559874 559404 559876
rect 586260 559874 586860 559876
rect -7636 553276 -7036 553278
rect 11604 553276 12204 553278
rect 47604 553276 48204 553278
rect 83604 553276 84204 553278
rect 119604 553276 120204 553278
rect 155604 553276 156204 553278
rect 191604 553276 192204 553278
rect 227604 553276 228204 553278
rect 263604 553276 264204 553278
rect 299604 553276 300204 553278
rect 335604 553276 336204 553278
rect 371604 553276 372204 553278
rect 407604 553276 408204 553278
rect 443604 553276 444204 553278
rect 479604 553276 480204 553278
rect 515604 553276 516204 553278
rect 551604 553276 552204 553278
rect 590960 553276 591560 553278
rect -8576 553254 592500 553276
rect -8576 553018 -7454 553254
rect -7218 553018 11786 553254
rect 12022 553018 47786 553254
rect 48022 553018 83786 553254
rect 84022 553018 119786 553254
rect 120022 553018 155786 553254
rect 156022 553018 191786 553254
rect 192022 553018 227786 553254
rect 228022 553018 263786 553254
rect 264022 553018 299786 553254
rect 300022 553018 335786 553254
rect 336022 553018 371786 553254
rect 372022 553018 407786 553254
rect 408022 553018 443786 553254
rect 444022 553018 479786 553254
rect 480022 553018 515786 553254
rect 516022 553018 551786 553254
rect 552022 553018 591142 553254
rect 591378 553018 592500 553254
rect -8576 552934 592500 553018
rect -8576 552698 -7454 552934
rect -7218 552698 11786 552934
rect 12022 552698 47786 552934
rect 48022 552698 83786 552934
rect 84022 552698 119786 552934
rect 120022 552698 155786 552934
rect 156022 552698 191786 552934
rect 192022 552698 227786 552934
rect 228022 552698 263786 552934
rect 264022 552698 299786 552934
rect 300022 552698 335786 552934
rect 336022 552698 371786 552934
rect 372022 552698 407786 552934
rect 408022 552698 443786 552934
rect 444022 552698 479786 552934
rect 480022 552698 515786 552934
rect 516022 552698 551786 552934
rect 552022 552698 591142 552934
rect 591378 552698 592500 552934
rect -8576 552676 592500 552698
rect -7636 552674 -7036 552676
rect 11604 552674 12204 552676
rect 47604 552674 48204 552676
rect 83604 552674 84204 552676
rect 119604 552674 120204 552676
rect 155604 552674 156204 552676
rect 191604 552674 192204 552676
rect 227604 552674 228204 552676
rect 263604 552674 264204 552676
rect 299604 552674 300204 552676
rect 335604 552674 336204 552676
rect 371604 552674 372204 552676
rect 407604 552674 408204 552676
rect 443604 552674 444204 552676
rect 479604 552674 480204 552676
rect 515604 552674 516204 552676
rect 551604 552674 552204 552676
rect 590960 552674 591560 552676
rect -5756 549676 -5156 549678
rect 8004 549676 8604 549678
rect 44004 549676 44604 549678
rect 80004 549676 80604 549678
rect 116004 549676 116604 549678
rect 152004 549676 152604 549678
rect 188004 549676 188604 549678
rect 224004 549676 224604 549678
rect 260004 549676 260604 549678
rect 296004 549676 296604 549678
rect 332004 549676 332604 549678
rect 368004 549676 368604 549678
rect 404004 549676 404604 549678
rect 440004 549676 440604 549678
rect 476004 549676 476604 549678
rect 512004 549676 512604 549678
rect 548004 549676 548604 549678
rect 589080 549676 589680 549678
rect -6696 549654 590620 549676
rect -6696 549418 -5574 549654
rect -5338 549418 8186 549654
rect 8422 549418 44186 549654
rect 44422 549418 80186 549654
rect 80422 549418 116186 549654
rect 116422 549418 152186 549654
rect 152422 549418 188186 549654
rect 188422 549418 224186 549654
rect 224422 549418 260186 549654
rect 260422 549418 296186 549654
rect 296422 549418 332186 549654
rect 332422 549418 368186 549654
rect 368422 549418 404186 549654
rect 404422 549418 440186 549654
rect 440422 549418 476186 549654
rect 476422 549418 512186 549654
rect 512422 549418 548186 549654
rect 548422 549418 589262 549654
rect 589498 549418 590620 549654
rect -6696 549334 590620 549418
rect -6696 549098 -5574 549334
rect -5338 549098 8186 549334
rect 8422 549098 44186 549334
rect 44422 549098 80186 549334
rect 80422 549098 116186 549334
rect 116422 549098 152186 549334
rect 152422 549098 188186 549334
rect 188422 549098 224186 549334
rect 224422 549098 260186 549334
rect 260422 549098 296186 549334
rect 296422 549098 332186 549334
rect 332422 549098 368186 549334
rect 368422 549098 404186 549334
rect 404422 549098 440186 549334
rect 440422 549098 476186 549334
rect 476422 549098 512186 549334
rect 512422 549098 548186 549334
rect 548422 549098 589262 549334
rect 589498 549098 590620 549334
rect -6696 549076 590620 549098
rect -5756 549074 -5156 549076
rect 8004 549074 8604 549076
rect 44004 549074 44604 549076
rect 80004 549074 80604 549076
rect 116004 549074 116604 549076
rect 152004 549074 152604 549076
rect 188004 549074 188604 549076
rect 224004 549074 224604 549076
rect 260004 549074 260604 549076
rect 296004 549074 296604 549076
rect 332004 549074 332604 549076
rect 368004 549074 368604 549076
rect 404004 549074 404604 549076
rect 440004 549074 440604 549076
rect 476004 549074 476604 549076
rect 512004 549074 512604 549076
rect 548004 549074 548604 549076
rect 589080 549074 589680 549076
rect -3876 546076 -3276 546078
rect 4404 546076 5004 546078
rect 40404 546076 41004 546078
rect 76404 546076 77004 546078
rect 112404 546076 113004 546078
rect 148404 546076 149004 546078
rect 184404 546076 185004 546078
rect 220404 546076 221004 546078
rect 256404 546076 257004 546078
rect 292404 546076 293004 546078
rect 328404 546076 329004 546078
rect 364404 546076 365004 546078
rect 400404 546076 401004 546078
rect 436404 546076 437004 546078
rect 472404 546076 473004 546078
rect 508404 546076 509004 546078
rect 544404 546076 545004 546078
rect 580404 546076 581004 546078
rect 587200 546076 587800 546078
rect -4816 546054 588740 546076
rect -4816 545818 -3694 546054
rect -3458 545818 4586 546054
rect 4822 545818 40586 546054
rect 40822 545818 76586 546054
rect 76822 545818 112586 546054
rect 112822 545818 148586 546054
rect 148822 545818 184586 546054
rect 184822 545818 220586 546054
rect 220822 545818 256586 546054
rect 256822 545818 292586 546054
rect 292822 545818 328586 546054
rect 328822 545818 364586 546054
rect 364822 545818 400586 546054
rect 400822 545818 436586 546054
rect 436822 545818 472586 546054
rect 472822 545818 508586 546054
rect 508822 545818 544586 546054
rect 544822 545818 580586 546054
rect 580822 545818 587382 546054
rect 587618 545818 588740 546054
rect -4816 545734 588740 545818
rect -4816 545498 -3694 545734
rect -3458 545498 4586 545734
rect 4822 545498 40586 545734
rect 40822 545498 76586 545734
rect 76822 545498 112586 545734
rect 112822 545498 148586 545734
rect 148822 545498 184586 545734
rect 184822 545498 220586 545734
rect 220822 545498 256586 545734
rect 256822 545498 292586 545734
rect 292822 545498 328586 545734
rect 328822 545498 364586 545734
rect 364822 545498 400586 545734
rect 400822 545498 436586 545734
rect 436822 545498 472586 545734
rect 472822 545498 508586 545734
rect 508822 545498 544586 545734
rect 544822 545498 580586 545734
rect 580822 545498 587382 545734
rect 587618 545498 588740 545734
rect -4816 545476 588740 545498
rect -3876 545474 -3276 545476
rect 4404 545474 5004 545476
rect 40404 545474 41004 545476
rect 76404 545474 77004 545476
rect 112404 545474 113004 545476
rect 148404 545474 149004 545476
rect 184404 545474 185004 545476
rect 220404 545474 221004 545476
rect 256404 545474 257004 545476
rect 292404 545474 293004 545476
rect 328404 545474 329004 545476
rect 364404 545474 365004 545476
rect 400404 545474 401004 545476
rect 436404 545474 437004 545476
rect 472404 545474 473004 545476
rect 508404 545474 509004 545476
rect 544404 545474 545004 545476
rect 580404 545474 581004 545476
rect 587200 545474 587800 545476
rect -1996 542476 -1396 542478
rect 804 542476 1404 542478
rect 36804 542476 37404 542478
rect 288804 542476 289404 542478
rect 324804 542476 325404 542478
rect 360804 542476 361404 542478
rect 396804 542476 397404 542478
rect 432804 542476 433404 542478
rect 468804 542476 469404 542478
rect 504804 542476 505404 542478
rect 540804 542476 541404 542478
rect 576804 542476 577404 542478
rect 585320 542476 585920 542478
rect -2936 542454 586860 542476
rect -2936 542218 -1814 542454
rect -1578 542218 986 542454
rect 1222 542218 36986 542454
rect 37222 542218 288986 542454
rect 289222 542218 324986 542454
rect 325222 542218 360986 542454
rect 361222 542218 396986 542454
rect 397222 542218 432986 542454
rect 433222 542218 468986 542454
rect 469222 542218 504986 542454
rect 505222 542218 540986 542454
rect 541222 542218 576986 542454
rect 577222 542218 585502 542454
rect 585738 542218 586860 542454
rect -2936 542134 586860 542218
rect -2936 541898 -1814 542134
rect -1578 541898 986 542134
rect 1222 541898 36986 542134
rect 37222 541898 288986 542134
rect 289222 541898 324986 542134
rect 325222 541898 360986 542134
rect 361222 541898 396986 542134
rect 397222 541898 432986 542134
rect 433222 541898 468986 542134
rect 469222 541898 504986 542134
rect 505222 541898 540986 542134
rect 541222 541898 576986 542134
rect 577222 541898 585502 542134
rect 585738 541898 586860 542134
rect -2936 541876 586860 541898
rect -1996 541874 -1396 541876
rect 804 541874 1404 541876
rect 36804 541874 37404 541876
rect 288804 541874 289404 541876
rect 324804 541874 325404 541876
rect 360804 541874 361404 541876
rect 396804 541874 397404 541876
rect 432804 541874 433404 541876
rect 468804 541874 469404 541876
rect 504804 541874 505404 541876
rect 540804 541874 541404 541876
rect 576804 541874 577404 541876
rect 585320 541874 585920 541876
rect -8576 535276 -7976 535278
rect 29604 535276 30204 535278
rect 79568 535276 79888 535278
rect 317604 535276 318204 535278
rect 353604 535276 354204 535278
rect 389604 535276 390204 535278
rect 425604 535276 426204 535278
rect 461604 535276 462204 535278
rect 497604 535276 498204 535278
rect 533604 535276 534204 535278
rect 569604 535276 570204 535278
rect 591900 535276 592500 535278
rect -8576 535254 592500 535276
rect -8576 535018 -8394 535254
rect -8158 535018 29786 535254
rect 30022 535018 79610 535254
rect 79846 535018 317786 535254
rect 318022 535018 353786 535254
rect 354022 535018 389786 535254
rect 390022 535018 425786 535254
rect 426022 535018 461786 535254
rect 462022 535018 497786 535254
rect 498022 535018 533786 535254
rect 534022 535018 569786 535254
rect 570022 535018 592082 535254
rect 592318 535018 592500 535254
rect -8576 534934 592500 535018
rect -8576 534698 -8394 534934
rect -8158 534698 29786 534934
rect 30022 534698 79610 534934
rect 79846 534698 317786 534934
rect 318022 534698 353786 534934
rect 354022 534698 389786 534934
rect 390022 534698 425786 534934
rect 426022 534698 461786 534934
rect 462022 534698 497786 534934
rect 498022 534698 533786 534934
rect 534022 534698 569786 534934
rect 570022 534698 592082 534934
rect 592318 534698 592500 534934
rect -8576 534676 592500 534698
rect -8576 534674 -7976 534676
rect 29604 534674 30204 534676
rect 79568 534674 79888 534676
rect 317604 534674 318204 534676
rect 353604 534674 354204 534676
rect 389604 534674 390204 534676
rect 425604 534674 426204 534676
rect 461604 534674 462204 534676
rect 497604 534674 498204 534676
rect 533604 534674 534204 534676
rect 569604 534674 570204 534676
rect 591900 534674 592500 534676
rect -6696 531676 -6096 531678
rect 26004 531676 26604 531678
rect 79568 531676 79888 531678
rect 314004 531676 314604 531678
rect 350004 531676 350604 531678
rect 386004 531676 386604 531678
rect 422004 531676 422604 531678
rect 458004 531676 458604 531678
rect 494004 531676 494604 531678
rect 530004 531676 530604 531678
rect 566004 531676 566604 531678
rect 590020 531676 590620 531678
rect -6696 531654 590620 531676
rect -6696 531418 -6514 531654
rect -6278 531418 26186 531654
rect 26422 531418 79610 531654
rect 79846 531418 314186 531654
rect 314422 531418 350186 531654
rect 350422 531418 386186 531654
rect 386422 531418 422186 531654
rect 422422 531418 458186 531654
rect 458422 531418 494186 531654
rect 494422 531418 530186 531654
rect 530422 531418 566186 531654
rect 566422 531418 590202 531654
rect 590438 531418 590620 531654
rect -6696 531334 590620 531418
rect -6696 531098 -6514 531334
rect -6278 531098 26186 531334
rect 26422 531098 79610 531334
rect 79846 531098 314186 531334
rect 314422 531098 350186 531334
rect 350422 531098 386186 531334
rect 386422 531098 422186 531334
rect 422422 531098 458186 531334
rect 458422 531098 494186 531334
rect 494422 531098 530186 531334
rect 530422 531098 566186 531334
rect 566422 531098 590202 531334
rect 590438 531098 590620 531334
rect -6696 531076 590620 531098
rect -6696 531074 -6096 531076
rect 26004 531074 26604 531076
rect 79568 531074 79888 531076
rect 314004 531074 314604 531076
rect 350004 531074 350604 531076
rect 386004 531074 386604 531076
rect 422004 531074 422604 531076
rect 458004 531074 458604 531076
rect 494004 531074 494604 531076
rect 530004 531074 530604 531076
rect 566004 531074 566604 531076
rect 590020 531074 590620 531076
rect -4816 528076 -4216 528078
rect 22404 528076 23004 528078
rect 79568 528076 79888 528078
rect 310404 528076 311004 528078
rect 346404 528076 347004 528078
rect 382404 528076 383004 528078
rect 418404 528076 419004 528078
rect 454404 528076 455004 528078
rect 490404 528076 491004 528078
rect 526404 528076 527004 528078
rect 562404 528076 563004 528078
rect 588140 528076 588740 528078
rect -4816 528054 588740 528076
rect -4816 527818 -4634 528054
rect -4398 527818 22586 528054
rect 22822 527818 79610 528054
rect 79846 527818 310586 528054
rect 310822 527818 346586 528054
rect 346822 527818 382586 528054
rect 382822 527818 418586 528054
rect 418822 527818 454586 528054
rect 454822 527818 490586 528054
rect 490822 527818 526586 528054
rect 526822 527818 562586 528054
rect 562822 527818 588322 528054
rect 588558 527818 588740 528054
rect -4816 527734 588740 527818
rect -4816 527498 -4634 527734
rect -4398 527498 22586 527734
rect 22822 527498 79610 527734
rect 79846 527498 310586 527734
rect 310822 527498 346586 527734
rect 346822 527498 382586 527734
rect 382822 527498 418586 527734
rect 418822 527498 454586 527734
rect 454822 527498 490586 527734
rect 490822 527498 526586 527734
rect 526822 527498 562586 527734
rect 562822 527498 588322 527734
rect 588558 527498 588740 527734
rect -4816 527476 588740 527498
rect -4816 527474 -4216 527476
rect 22404 527474 23004 527476
rect 79568 527474 79888 527476
rect 310404 527474 311004 527476
rect 346404 527474 347004 527476
rect 382404 527474 383004 527476
rect 418404 527474 419004 527476
rect 454404 527474 455004 527476
rect 490404 527474 491004 527476
rect 526404 527474 527004 527476
rect 562404 527474 563004 527476
rect 588140 527474 588740 527476
rect -2936 524476 -2336 524478
rect 18804 524476 19404 524478
rect 54804 524476 55404 524478
rect 79568 524476 79888 524478
rect 306804 524476 307404 524478
rect 342804 524476 343404 524478
rect 378804 524476 379404 524478
rect 414804 524476 415404 524478
rect 450804 524476 451404 524478
rect 486804 524476 487404 524478
rect 522804 524476 523404 524478
rect 558804 524476 559404 524478
rect 586260 524476 586860 524478
rect -2936 524454 586860 524476
rect -2936 524218 -2754 524454
rect -2518 524218 18986 524454
rect 19222 524218 54986 524454
rect 55222 524218 79610 524454
rect 79846 524218 306986 524454
rect 307222 524218 342986 524454
rect 343222 524218 378986 524454
rect 379222 524218 414986 524454
rect 415222 524218 450986 524454
rect 451222 524218 486986 524454
rect 487222 524218 522986 524454
rect 523222 524218 558986 524454
rect 559222 524218 586442 524454
rect 586678 524218 586860 524454
rect -2936 524134 586860 524218
rect -2936 523898 -2754 524134
rect -2518 523898 18986 524134
rect 19222 523898 54986 524134
rect 55222 523898 79610 524134
rect 79846 523898 306986 524134
rect 307222 523898 342986 524134
rect 343222 523898 378986 524134
rect 379222 523898 414986 524134
rect 415222 523898 450986 524134
rect 451222 523898 486986 524134
rect 487222 523898 522986 524134
rect 523222 523898 558986 524134
rect 559222 523898 586442 524134
rect 586678 523898 586860 524134
rect -2936 523876 586860 523898
rect -2936 523874 -2336 523876
rect 18804 523874 19404 523876
rect 54804 523874 55404 523876
rect 79568 523874 79888 523876
rect 306804 523874 307404 523876
rect 342804 523874 343404 523876
rect 378804 523874 379404 523876
rect 414804 523874 415404 523876
rect 450804 523874 451404 523876
rect 486804 523874 487404 523876
rect 522804 523874 523404 523876
rect 558804 523874 559404 523876
rect 586260 523874 586860 523876
rect -7636 517276 -7036 517278
rect 11604 517276 12204 517278
rect 47604 517276 48204 517278
rect 64208 517276 64528 517278
rect 299604 517276 300204 517278
rect 335604 517276 336204 517278
rect 371604 517276 372204 517278
rect 407604 517276 408204 517278
rect 443604 517276 444204 517278
rect 479604 517276 480204 517278
rect 515604 517276 516204 517278
rect 551604 517276 552204 517278
rect 590960 517276 591560 517278
rect -8576 517254 592500 517276
rect -8576 517018 -7454 517254
rect -7218 517018 11786 517254
rect 12022 517018 47786 517254
rect 48022 517018 64250 517254
rect 64486 517018 299786 517254
rect 300022 517018 335786 517254
rect 336022 517018 371786 517254
rect 372022 517018 407786 517254
rect 408022 517018 443786 517254
rect 444022 517018 479786 517254
rect 480022 517018 515786 517254
rect 516022 517018 551786 517254
rect 552022 517018 591142 517254
rect 591378 517018 592500 517254
rect -8576 516934 592500 517018
rect -8576 516698 -7454 516934
rect -7218 516698 11786 516934
rect 12022 516698 47786 516934
rect 48022 516698 64250 516934
rect 64486 516698 299786 516934
rect 300022 516698 335786 516934
rect 336022 516698 371786 516934
rect 372022 516698 407786 516934
rect 408022 516698 443786 516934
rect 444022 516698 479786 516934
rect 480022 516698 515786 516934
rect 516022 516698 551786 516934
rect 552022 516698 591142 516934
rect 591378 516698 592500 516934
rect -8576 516676 592500 516698
rect -7636 516674 -7036 516676
rect 11604 516674 12204 516676
rect 47604 516674 48204 516676
rect 64208 516674 64528 516676
rect 299604 516674 300204 516676
rect 335604 516674 336204 516676
rect 371604 516674 372204 516676
rect 407604 516674 408204 516676
rect 443604 516674 444204 516676
rect 479604 516674 480204 516676
rect 515604 516674 516204 516676
rect 551604 516674 552204 516676
rect 590960 516674 591560 516676
rect -5756 513676 -5156 513678
rect 8004 513676 8604 513678
rect 44004 513676 44604 513678
rect 64208 513676 64528 513678
rect 296004 513676 296604 513678
rect 332004 513676 332604 513678
rect 368004 513676 368604 513678
rect 404004 513676 404604 513678
rect 440004 513676 440604 513678
rect 476004 513676 476604 513678
rect 512004 513676 512604 513678
rect 548004 513676 548604 513678
rect 589080 513676 589680 513678
rect -6696 513654 590620 513676
rect -6696 513418 -5574 513654
rect -5338 513418 8186 513654
rect 8422 513418 44186 513654
rect 44422 513418 64250 513654
rect 64486 513418 296186 513654
rect 296422 513418 332186 513654
rect 332422 513418 368186 513654
rect 368422 513418 404186 513654
rect 404422 513418 440186 513654
rect 440422 513418 476186 513654
rect 476422 513418 512186 513654
rect 512422 513418 548186 513654
rect 548422 513418 589262 513654
rect 589498 513418 590620 513654
rect -6696 513334 590620 513418
rect -6696 513098 -5574 513334
rect -5338 513098 8186 513334
rect 8422 513098 44186 513334
rect 44422 513098 64250 513334
rect 64486 513098 296186 513334
rect 296422 513098 332186 513334
rect 332422 513098 368186 513334
rect 368422 513098 404186 513334
rect 404422 513098 440186 513334
rect 440422 513098 476186 513334
rect 476422 513098 512186 513334
rect 512422 513098 548186 513334
rect 548422 513098 589262 513334
rect 589498 513098 590620 513334
rect -6696 513076 590620 513098
rect -5756 513074 -5156 513076
rect 8004 513074 8604 513076
rect 44004 513074 44604 513076
rect 64208 513074 64528 513076
rect 296004 513074 296604 513076
rect 332004 513074 332604 513076
rect 368004 513074 368604 513076
rect 404004 513074 404604 513076
rect 440004 513074 440604 513076
rect 476004 513074 476604 513076
rect 512004 513074 512604 513076
rect 548004 513074 548604 513076
rect 589080 513074 589680 513076
rect -3876 510076 -3276 510078
rect 4404 510076 5004 510078
rect 40404 510076 41004 510078
rect 64208 510076 64528 510078
rect 292404 510076 293004 510078
rect 328404 510076 329004 510078
rect 364404 510076 365004 510078
rect 400404 510076 401004 510078
rect 436404 510076 437004 510078
rect 472404 510076 473004 510078
rect 508404 510076 509004 510078
rect 544404 510076 545004 510078
rect 580404 510076 581004 510078
rect 587200 510076 587800 510078
rect -4816 510054 588740 510076
rect -4816 509818 -3694 510054
rect -3458 509818 4586 510054
rect 4822 509818 40586 510054
rect 40822 509818 64250 510054
rect 64486 509818 292586 510054
rect 292822 509818 328586 510054
rect 328822 509818 364586 510054
rect 364822 509818 400586 510054
rect 400822 509818 436586 510054
rect 436822 509818 472586 510054
rect 472822 509818 508586 510054
rect 508822 509818 544586 510054
rect 544822 509818 580586 510054
rect 580822 509818 587382 510054
rect 587618 509818 588740 510054
rect -4816 509734 588740 509818
rect -4816 509498 -3694 509734
rect -3458 509498 4586 509734
rect 4822 509498 40586 509734
rect 40822 509498 64250 509734
rect 64486 509498 292586 509734
rect 292822 509498 328586 509734
rect 328822 509498 364586 509734
rect 364822 509498 400586 509734
rect 400822 509498 436586 509734
rect 436822 509498 472586 509734
rect 472822 509498 508586 509734
rect 508822 509498 544586 509734
rect 544822 509498 580586 509734
rect 580822 509498 587382 509734
rect 587618 509498 588740 509734
rect -4816 509476 588740 509498
rect -3876 509474 -3276 509476
rect 4404 509474 5004 509476
rect 40404 509474 41004 509476
rect 64208 509474 64528 509476
rect 292404 509474 293004 509476
rect 328404 509474 329004 509476
rect 364404 509474 365004 509476
rect 400404 509474 401004 509476
rect 436404 509474 437004 509476
rect 472404 509474 473004 509476
rect 508404 509474 509004 509476
rect 544404 509474 545004 509476
rect 580404 509474 581004 509476
rect 587200 509474 587800 509476
rect -1996 506476 -1396 506478
rect 804 506476 1404 506478
rect 36804 506476 37404 506478
rect 64208 506476 64528 506478
rect 288804 506476 289404 506478
rect 324804 506476 325404 506478
rect 360804 506476 361404 506478
rect 396804 506476 397404 506478
rect 432804 506476 433404 506478
rect 468804 506476 469404 506478
rect 504804 506476 505404 506478
rect 540804 506476 541404 506478
rect 576804 506476 577404 506478
rect 585320 506476 585920 506478
rect -2936 506454 586860 506476
rect -2936 506218 -1814 506454
rect -1578 506218 986 506454
rect 1222 506218 36986 506454
rect 37222 506218 64250 506454
rect 64486 506218 288986 506454
rect 289222 506218 324986 506454
rect 325222 506218 360986 506454
rect 361222 506218 396986 506454
rect 397222 506218 432986 506454
rect 433222 506218 468986 506454
rect 469222 506218 504986 506454
rect 505222 506218 540986 506454
rect 541222 506218 576986 506454
rect 577222 506218 585502 506454
rect 585738 506218 586860 506454
rect -2936 506134 586860 506218
rect -2936 505898 -1814 506134
rect -1578 505898 986 506134
rect 1222 505898 36986 506134
rect 37222 505898 64250 506134
rect 64486 505898 288986 506134
rect 289222 505898 324986 506134
rect 325222 505898 360986 506134
rect 361222 505898 396986 506134
rect 397222 505898 432986 506134
rect 433222 505898 468986 506134
rect 469222 505898 504986 506134
rect 505222 505898 540986 506134
rect 541222 505898 576986 506134
rect 577222 505898 585502 506134
rect 585738 505898 586860 506134
rect -2936 505876 586860 505898
rect -1996 505874 -1396 505876
rect 804 505874 1404 505876
rect 36804 505874 37404 505876
rect 64208 505874 64528 505876
rect 288804 505874 289404 505876
rect 324804 505874 325404 505876
rect 360804 505874 361404 505876
rect 396804 505874 397404 505876
rect 432804 505874 433404 505876
rect 468804 505874 469404 505876
rect 504804 505874 505404 505876
rect 540804 505874 541404 505876
rect 576804 505874 577404 505876
rect 585320 505874 585920 505876
rect -8576 499276 -7976 499278
rect 29604 499276 30204 499278
rect 79568 499276 79888 499278
rect 317604 499276 318204 499278
rect 353604 499276 354204 499278
rect 389604 499276 390204 499278
rect 425604 499276 426204 499278
rect 461604 499276 462204 499278
rect 497604 499276 498204 499278
rect 533604 499276 534204 499278
rect 569604 499276 570204 499278
rect 591900 499276 592500 499278
rect -8576 499254 592500 499276
rect -8576 499018 -8394 499254
rect -8158 499018 29786 499254
rect 30022 499018 79610 499254
rect 79846 499018 317786 499254
rect 318022 499018 353786 499254
rect 354022 499018 389786 499254
rect 390022 499018 425786 499254
rect 426022 499018 461786 499254
rect 462022 499018 497786 499254
rect 498022 499018 533786 499254
rect 534022 499018 569786 499254
rect 570022 499018 592082 499254
rect 592318 499018 592500 499254
rect -8576 498934 592500 499018
rect -8576 498698 -8394 498934
rect -8158 498698 29786 498934
rect 30022 498698 79610 498934
rect 79846 498698 317786 498934
rect 318022 498698 353786 498934
rect 354022 498698 389786 498934
rect 390022 498698 425786 498934
rect 426022 498698 461786 498934
rect 462022 498698 497786 498934
rect 498022 498698 533786 498934
rect 534022 498698 569786 498934
rect 570022 498698 592082 498934
rect 592318 498698 592500 498934
rect -8576 498676 592500 498698
rect -8576 498674 -7976 498676
rect 29604 498674 30204 498676
rect 79568 498674 79888 498676
rect 317604 498674 318204 498676
rect 353604 498674 354204 498676
rect 389604 498674 390204 498676
rect 425604 498674 426204 498676
rect 461604 498674 462204 498676
rect 497604 498674 498204 498676
rect 533604 498674 534204 498676
rect 569604 498674 570204 498676
rect 591900 498674 592500 498676
rect -6696 495676 -6096 495678
rect 26004 495676 26604 495678
rect 79568 495676 79888 495678
rect 314004 495676 314604 495678
rect 350004 495676 350604 495678
rect 386004 495676 386604 495678
rect 422004 495676 422604 495678
rect 458004 495676 458604 495678
rect 494004 495676 494604 495678
rect 530004 495676 530604 495678
rect 566004 495676 566604 495678
rect 590020 495676 590620 495678
rect -6696 495654 590620 495676
rect -6696 495418 -6514 495654
rect -6278 495418 26186 495654
rect 26422 495418 79610 495654
rect 79846 495418 314186 495654
rect 314422 495418 350186 495654
rect 350422 495418 386186 495654
rect 386422 495418 422186 495654
rect 422422 495418 458186 495654
rect 458422 495418 494186 495654
rect 494422 495418 530186 495654
rect 530422 495418 566186 495654
rect 566422 495418 590202 495654
rect 590438 495418 590620 495654
rect -6696 495334 590620 495418
rect -6696 495098 -6514 495334
rect -6278 495098 26186 495334
rect 26422 495098 79610 495334
rect 79846 495098 314186 495334
rect 314422 495098 350186 495334
rect 350422 495098 386186 495334
rect 386422 495098 422186 495334
rect 422422 495098 458186 495334
rect 458422 495098 494186 495334
rect 494422 495098 530186 495334
rect 530422 495098 566186 495334
rect 566422 495098 590202 495334
rect 590438 495098 590620 495334
rect -6696 495076 590620 495098
rect -6696 495074 -6096 495076
rect 26004 495074 26604 495076
rect 79568 495074 79888 495076
rect 314004 495074 314604 495076
rect 350004 495074 350604 495076
rect 386004 495074 386604 495076
rect 422004 495074 422604 495076
rect 458004 495074 458604 495076
rect 494004 495074 494604 495076
rect 530004 495074 530604 495076
rect 566004 495074 566604 495076
rect 590020 495074 590620 495076
rect -4816 492076 -4216 492078
rect 22404 492076 23004 492078
rect 79568 492076 79888 492078
rect 310404 492076 311004 492078
rect 346404 492076 347004 492078
rect 382404 492076 383004 492078
rect 418404 492076 419004 492078
rect 454404 492076 455004 492078
rect 490404 492076 491004 492078
rect 526404 492076 527004 492078
rect 562404 492076 563004 492078
rect 588140 492076 588740 492078
rect -4816 492054 588740 492076
rect -4816 491818 -4634 492054
rect -4398 491818 22586 492054
rect 22822 491818 79610 492054
rect 79846 491818 310586 492054
rect 310822 491818 346586 492054
rect 346822 491818 382586 492054
rect 382822 491818 418586 492054
rect 418822 491818 454586 492054
rect 454822 491818 490586 492054
rect 490822 491818 526586 492054
rect 526822 491818 562586 492054
rect 562822 491818 588322 492054
rect 588558 491818 588740 492054
rect -4816 491734 588740 491818
rect -4816 491498 -4634 491734
rect -4398 491498 22586 491734
rect 22822 491498 79610 491734
rect 79846 491498 310586 491734
rect 310822 491498 346586 491734
rect 346822 491498 382586 491734
rect 382822 491498 418586 491734
rect 418822 491498 454586 491734
rect 454822 491498 490586 491734
rect 490822 491498 526586 491734
rect 526822 491498 562586 491734
rect 562822 491498 588322 491734
rect 588558 491498 588740 491734
rect -4816 491476 588740 491498
rect -4816 491474 -4216 491476
rect 22404 491474 23004 491476
rect 79568 491474 79888 491476
rect 310404 491474 311004 491476
rect 346404 491474 347004 491476
rect 382404 491474 383004 491476
rect 418404 491474 419004 491476
rect 454404 491474 455004 491476
rect 490404 491474 491004 491476
rect 526404 491474 527004 491476
rect 562404 491474 563004 491476
rect 588140 491474 588740 491476
rect -2936 488476 -2336 488478
rect 18804 488476 19404 488478
rect 54804 488476 55404 488478
rect 79568 488476 79888 488478
rect 306804 488476 307404 488478
rect 342804 488476 343404 488478
rect 378804 488476 379404 488478
rect 414804 488476 415404 488478
rect 450804 488476 451404 488478
rect 486804 488476 487404 488478
rect 522804 488476 523404 488478
rect 558804 488476 559404 488478
rect 586260 488476 586860 488478
rect -2936 488454 586860 488476
rect -2936 488218 -2754 488454
rect -2518 488218 18986 488454
rect 19222 488218 54986 488454
rect 55222 488218 79610 488454
rect 79846 488218 306986 488454
rect 307222 488218 342986 488454
rect 343222 488218 378986 488454
rect 379222 488218 414986 488454
rect 415222 488218 450986 488454
rect 451222 488218 486986 488454
rect 487222 488218 522986 488454
rect 523222 488218 558986 488454
rect 559222 488218 586442 488454
rect 586678 488218 586860 488454
rect -2936 488134 586860 488218
rect -2936 487898 -2754 488134
rect -2518 487898 18986 488134
rect 19222 487898 54986 488134
rect 55222 487898 79610 488134
rect 79846 487898 306986 488134
rect 307222 487898 342986 488134
rect 343222 487898 378986 488134
rect 379222 487898 414986 488134
rect 415222 487898 450986 488134
rect 451222 487898 486986 488134
rect 487222 487898 522986 488134
rect 523222 487898 558986 488134
rect 559222 487898 586442 488134
rect 586678 487898 586860 488134
rect -2936 487876 586860 487898
rect -2936 487874 -2336 487876
rect 18804 487874 19404 487876
rect 54804 487874 55404 487876
rect 79568 487874 79888 487876
rect 306804 487874 307404 487876
rect 342804 487874 343404 487876
rect 378804 487874 379404 487876
rect 414804 487874 415404 487876
rect 450804 487874 451404 487876
rect 486804 487874 487404 487876
rect 522804 487874 523404 487876
rect 558804 487874 559404 487876
rect 586260 487874 586860 487876
rect -7636 481276 -7036 481278
rect 11604 481276 12204 481278
rect 47604 481276 48204 481278
rect 64208 481276 64528 481278
rect 299604 481276 300204 481278
rect 335604 481276 336204 481278
rect 371604 481276 372204 481278
rect 407604 481276 408204 481278
rect 443604 481276 444204 481278
rect 479604 481276 480204 481278
rect 515604 481276 516204 481278
rect 551604 481276 552204 481278
rect 590960 481276 591560 481278
rect -8576 481254 592500 481276
rect -8576 481018 -7454 481254
rect -7218 481018 11786 481254
rect 12022 481018 47786 481254
rect 48022 481018 64250 481254
rect 64486 481018 299786 481254
rect 300022 481018 335786 481254
rect 336022 481018 371786 481254
rect 372022 481018 407786 481254
rect 408022 481018 443786 481254
rect 444022 481018 479786 481254
rect 480022 481018 515786 481254
rect 516022 481018 551786 481254
rect 552022 481018 591142 481254
rect 591378 481018 592500 481254
rect -8576 480934 592500 481018
rect -8576 480698 -7454 480934
rect -7218 480698 11786 480934
rect 12022 480698 47786 480934
rect 48022 480698 64250 480934
rect 64486 480698 299786 480934
rect 300022 480698 335786 480934
rect 336022 480698 371786 480934
rect 372022 480698 407786 480934
rect 408022 480698 443786 480934
rect 444022 480698 479786 480934
rect 480022 480698 515786 480934
rect 516022 480698 551786 480934
rect 552022 480698 591142 480934
rect 591378 480698 592500 480934
rect -8576 480676 592500 480698
rect -7636 480674 -7036 480676
rect 11604 480674 12204 480676
rect 47604 480674 48204 480676
rect 64208 480674 64528 480676
rect 299604 480674 300204 480676
rect 335604 480674 336204 480676
rect 371604 480674 372204 480676
rect 407604 480674 408204 480676
rect 443604 480674 444204 480676
rect 479604 480674 480204 480676
rect 515604 480674 516204 480676
rect 551604 480674 552204 480676
rect 590960 480674 591560 480676
rect -5756 477676 -5156 477678
rect 8004 477676 8604 477678
rect 44004 477676 44604 477678
rect 64208 477676 64528 477678
rect 296004 477676 296604 477678
rect 332004 477676 332604 477678
rect 368004 477676 368604 477678
rect 404004 477676 404604 477678
rect 440004 477676 440604 477678
rect 476004 477676 476604 477678
rect 512004 477676 512604 477678
rect 548004 477676 548604 477678
rect 589080 477676 589680 477678
rect -6696 477654 590620 477676
rect -6696 477418 -5574 477654
rect -5338 477418 8186 477654
rect 8422 477418 44186 477654
rect 44422 477418 64250 477654
rect 64486 477418 296186 477654
rect 296422 477418 332186 477654
rect 332422 477418 368186 477654
rect 368422 477418 404186 477654
rect 404422 477418 440186 477654
rect 440422 477418 476186 477654
rect 476422 477418 512186 477654
rect 512422 477418 548186 477654
rect 548422 477418 589262 477654
rect 589498 477418 590620 477654
rect -6696 477334 590620 477418
rect -6696 477098 -5574 477334
rect -5338 477098 8186 477334
rect 8422 477098 44186 477334
rect 44422 477098 64250 477334
rect 64486 477098 296186 477334
rect 296422 477098 332186 477334
rect 332422 477098 368186 477334
rect 368422 477098 404186 477334
rect 404422 477098 440186 477334
rect 440422 477098 476186 477334
rect 476422 477098 512186 477334
rect 512422 477098 548186 477334
rect 548422 477098 589262 477334
rect 589498 477098 590620 477334
rect -6696 477076 590620 477098
rect -5756 477074 -5156 477076
rect 8004 477074 8604 477076
rect 44004 477074 44604 477076
rect 64208 477074 64528 477076
rect 296004 477074 296604 477076
rect 332004 477074 332604 477076
rect 368004 477074 368604 477076
rect 404004 477074 404604 477076
rect 440004 477074 440604 477076
rect 476004 477074 476604 477076
rect 512004 477074 512604 477076
rect 548004 477074 548604 477076
rect 589080 477074 589680 477076
rect -3876 474076 -3276 474078
rect 4404 474076 5004 474078
rect 40404 474076 41004 474078
rect 64208 474076 64528 474078
rect 292404 474076 293004 474078
rect 328404 474076 329004 474078
rect 364404 474076 365004 474078
rect 400404 474076 401004 474078
rect 436404 474076 437004 474078
rect 472404 474076 473004 474078
rect 508404 474076 509004 474078
rect 544404 474076 545004 474078
rect 580404 474076 581004 474078
rect 587200 474076 587800 474078
rect -4816 474054 588740 474076
rect -4816 473818 -3694 474054
rect -3458 473818 4586 474054
rect 4822 473818 40586 474054
rect 40822 473818 64250 474054
rect 64486 473818 292586 474054
rect 292822 473818 328586 474054
rect 328822 473818 364586 474054
rect 364822 473818 400586 474054
rect 400822 473818 436586 474054
rect 436822 473818 472586 474054
rect 472822 473818 508586 474054
rect 508822 473818 544586 474054
rect 544822 473818 580586 474054
rect 580822 473818 587382 474054
rect 587618 473818 588740 474054
rect -4816 473734 588740 473818
rect -4816 473498 -3694 473734
rect -3458 473498 4586 473734
rect 4822 473498 40586 473734
rect 40822 473498 64250 473734
rect 64486 473498 292586 473734
rect 292822 473498 328586 473734
rect 328822 473498 364586 473734
rect 364822 473498 400586 473734
rect 400822 473498 436586 473734
rect 436822 473498 472586 473734
rect 472822 473498 508586 473734
rect 508822 473498 544586 473734
rect 544822 473498 580586 473734
rect 580822 473498 587382 473734
rect 587618 473498 588740 473734
rect -4816 473476 588740 473498
rect -3876 473474 -3276 473476
rect 4404 473474 5004 473476
rect 40404 473474 41004 473476
rect 64208 473474 64528 473476
rect 292404 473474 293004 473476
rect 328404 473474 329004 473476
rect 364404 473474 365004 473476
rect 400404 473474 401004 473476
rect 436404 473474 437004 473476
rect 472404 473474 473004 473476
rect 508404 473474 509004 473476
rect 544404 473474 545004 473476
rect 580404 473474 581004 473476
rect 587200 473474 587800 473476
rect -1996 470476 -1396 470478
rect 804 470476 1404 470478
rect 36804 470476 37404 470478
rect 64208 470476 64528 470478
rect 288804 470476 289404 470478
rect 324804 470476 325404 470478
rect 360804 470476 361404 470478
rect 396804 470476 397404 470478
rect 432804 470476 433404 470478
rect 468804 470476 469404 470478
rect 504804 470476 505404 470478
rect 540804 470476 541404 470478
rect 576804 470476 577404 470478
rect 585320 470476 585920 470478
rect -2936 470454 586860 470476
rect -2936 470218 -1814 470454
rect -1578 470218 986 470454
rect 1222 470218 36986 470454
rect 37222 470218 64250 470454
rect 64486 470218 288986 470454
rect 289222 470218 324986 470454
rect 325222 470218 360986 470454
rect 361222 470218 396986 470454
rect 397222 470218 432986 470454
rect 433222 470218 468986 470454
rect 469222 470218 504986 470454
rect 505222 470218 540986 470454
rect 541222 470218 576986 470454
rect 577222 470218 585502 470454
rect 585738 470218 586860 470454
rect -2936 470134 586860 470218
rect -2936 469898 -1814 470134
rect -1578 469898 986 470134
rect 1222 469898 36986 470134
rect 37222 469898 64250 470134
rect 64486 469898 288986 470134
rect 289222 469898 324986 470134
rect 325222 469898 360986 470134
rect 361222 469898 396986 470134
rect 397222 469898 432986 470134
rect 433222 469898 468986 470134
rect 469222 469898 504986 470134
rect 505222 469898 540986 470134
rect 541222 469898 576986 470134
rect 577222 469898 585502 470134
rect 585738 469898 586860 470134
rect -2936 469876 586860 469898
rect -1996 469874 -1396 469876
rect 804 469874 1404 469876
rect 36804 469874 37404 469876
rect 64208 469874 64528 469876
rect 288804 469874 289404 469876
rect 324804 469874 325404 469876
rect 360804 469874 361404 469876
rect 396804 469874 397404 469876
rect 432804 469874 433404 469876
rect 468804 469874 469404 469876
rect 504804 469874 505404 469876
rect 540804 469874 541404 469876
rect 576804 469874 577404 469876
rect 585320 469874 585920 469876
rect -8576 463276 -7976 463278
rect 29604 463276 30204 463278
rect 79568 463276 79888 463278
rect 317604 463276 318204 463278
rect 353604 463276 354204 463278
rect 389604 463276 390204 463278
rect 425604 463276 426204 463278
rect 461604 463276 462204 463278
rect 497604 463276 498204 463278
rect 533604 463276 534204 463278
rect 569604 463276 570204 463278
rect 591900 463276 592500 463278
rect -8576 463254 592500 463276
rect -8576 463018 -8394 463254
rect -8158 463018 29786 463254
rect 30022 463018 79610 463254
rect 79846 463018 317786 463254
rect 318022 463018 353786 463254
rect 354022 463018 389786 463254
rect 390022 463018 425786 463254
rect 426022 463018 461786 463254
rect 462022 463018 497786 463254
rect 498022 463018 533786 463254
rect 534022 463018 569786 463254
rect 570022 463018 592082 463254
rect 592318 463018 592500 463254
rect -8576 462934 592500 463018
rect -8576 462698 -8394 462934
rect -8158 462698 29786 462934
rect 30022 462698 79610 462934
rect 79846 462698 317786 462934
rect 318022 462698 353786 462934
rect 354022 462698 389786 462934
rect 390022 462698 425786 462934
rect 426022 462698 461786 462934
rect 462022 462698 497786 462934
rect 498022 462698 533786 462934
rect 534022 462698 569786 462934
rect 570022 462698 592082 462934
rect 592318 462698 592500 462934
rect -8576 462676 592500 462698
rect -8576 462674 -7976 462676
rect 29604 462674 30204 462676
rect 79568 462674 79888 462676
rect 317604 462674 318204 462676
rect 353604 462674 354204 462676
rect 389604 462674 390204 462676
rect 425604 462674 426204 462676
rect 461604 462674 462204 462676
rect 497604 462674 498204 462676
rect 533604 462674 534204 462676
rect 569604 462674 570204 462676
rect 591900 462674 592500 462676
rect -6696 459676 -6096 459678
rect 26004 459676 26604 459678
rect 79568 459676 79888 459678
rect 314004 459676 314604 459678
rect 350004 459676 350604 459678
rect 386004 459676 386604 459678
rect 422004 459676 422604 459678
rect 458004 459676 458604 459678
rect 494004 459676 494604 459678
rect 530004 459676 530604 459678
rect 566004 459676 566604 459678
rect 590020 459676 590620 459678
rect -6696 459654 590620 459676
rect -6696 459418 -6514 459654
rect -6278 459418 26186 459654
rect 26422 459418 79610 459654
rect 79846 459418 314186 459654
rect 314422 459418 350186 459654
rect 350422 459418 386186 459654
rect 386422 459418 422186 459654
rect 422422 459418 458186 459654
rect 458422 459418 494186 459654
rect 494422 459418 530186 459654
rect 530422 459418 566186 459654
rect 566422 459418 590202 459654
rect 590438 459418 590620 459654
rect -6696 459334 590620 459418
rect -6696 459098 -6514 459334
rect -6278 459098 26186 459334
rect 26422 459098 79610 459334
rect 79846 459098 314186 459334
rect 314422 459098 350186 459334
rect 350422 459098 386186 459334
rect 386422 459098 422186 459334
rect 422422 459098 458186 459334
rect 458422 459098 494186 459334
rect 494422 459098 530186 459334
rect 530422 459098 566186 459334
rect 566422 459098 590202 459334
rect 590438 459098 590620 459334
rect -6696 459076 590620 459098
rect -6696 459074 -6096 459076
rect 26004 459074 26604 459076
rect 79568 459074 79888 459076
rect 314004 459074 314604 459076
rect 350004 459074 350604 459076
rect 386004 459074 386604 459076
rect 422004 459074 422604 459076
rect 458004 459074 458604 459076
rect 494004 459074 494604 459076
rect 530004 459074 530604 459076
rect 566004 459074 566604 459076
rect 590020 459074 590620 459076
rect -4816 456076 -4216 456078
rect 22404 456076 23004 456078
rect 79568 456076 79888 456078
rect 310404 456076 311004 456078
rect 346404 456076 347004 456078
rect 382404 456076 383004 456078
rect 418404 456076 419004 456078
rect 454404 456076 455004 456078
rect 490404 456076 491004 456078
rect 526404 456076 527004 456078
rect 562404 456076 563004 456078
rect 588140 456076 588740 456078
rect -4816 456054 588740 456076
rect -4816 455818 -4634 456054
rect -4398 455818 22586 456054
rect 22822 455818 79610 456054
rect 79846 455818 310586 456054
rect 310822 455818 346586 456054
rect 346822 455818 382586 456054
rect 382822 455818 418586 456054
rect 418822 455818 454586 456054
rect 454822 455818 490586 456054
rect 490822 455818 526586 456054
rect 526822 455818 562586 456054
rect 562822 455818 588322 456054
rect 588558 455818 588740 456054
rect -4816 455734 588740 455818
rect -4816 455498 -4634 455734
rect -4398 455498 22586 455734
rect 22822 455498 79610 455734
rect 79846 455498 310586 455734
rect 310822 455498 346586 455734
rect 346822 455498 382586 455734
rect 382822 455498 418586 455734
rect 418822 455498 454586 455734
rect 454822 455498 490586 455734
rect 490822 455498 526586 455734
rect 526822 455498 562586 455734
rect 562822 455498 588322 455734
rect 588558 455498 588740 455734
rect -4816 455476 588740 455498
rect -4816 455474 -4216 455476
rect 22404 455474 23004 455476
rect 79568 455474 79888 455476
rect 310404 455474 311004 455476
rect 346404 455474 347004 455476
rect 382404 455474 383004 455476
rect 418404 455474 419004 455476
rect 454404 455474 455004 455476
rect 490404 455474 491004 455476
rect 526404 455474 527004 455476
rect 562404 455474 563004 455476
rect 588140 455474 588740 455476
rect -2936 452476 -2336 452478
rect 18804 452476 19404 452478
rect 54804 452476 55404 452478
rect 79568 452476 79888 452478
rect 306804 452476 307404 452478
rect 342804 452476 343404 452478
rect 378804 452476 379404 452478
rect 414804 452476 415404 452478
rect 450804 452476 451404 452478
rect 486804 452476 487404 452478
rect 522804 452476 523404 452478
rect 558804 452476 559404 452478
rect 586260 452476 586860 452478
rect -2936 452454 586860 452476
rect -2936 452218 -2754 452454
rect -2518 452218 18986 452454
rect 19222 452218 54986 452454
rect 55222 452218 79610 452454
rect 79846 452218 306986 452454
rect 307222 452218 342986 452454
rect 343222 452218 378986 452454
rect 379222 452218 414986 452454
rect 415222 452218 450986 452454
rect 451222 452218 486986 452454
rect 487222 452218 522986 452454
rect 523222 452218 558986 452454
rect 559222 452218 586442 452454
rect 586678 452218 586860 452454
rect -2936 452134 586860 452218
rect -2936 451898 -2754 452134
rect -2518 451898 18986 452134
rect 19222 451898 54986 452134
rect 55222 451898 79610 452134
rect 79846 451898 306986 452134
rect 307222 451898 342986 452134
rect 343222 451898 378986 452134
rect 379222 451898 414986 452134
rect 415222 451898 450986 452134
rect 451222 451898 486986 452134
rect 487222 451898 522986 452134
rect 523222 451898 558986 452134
rect 559222 451898 586442 452134
rect 586678 451898 586860 452134
rect -2936 451876 586860 451898
rect -2936 451874 -2336 451876
rect 18804 451874 19404 451876
rect 54804 451874 55404 451876
rect 79568 451874 79888 451876
rect 306804 451874 307404 451876
rect 342804 451874 343404 451876
rect 378804 451874 379404 451876
rect 414804 451874 415404 451876
rect 450804 451874 451404 451876
rect 486804 451874 487404 451876
rect 522804 451874 523404 451876
rect 558804 451874 559404 451876
rect 586260 451874 586860 451876
rect -7636 445276 -7036 445278
rect 11604 445276 12204 445278
rect 47604 445276 48204 445278
rect 64208 445276 64528 445278
rect 299604 445276 300204 445278
rect 335604 445276 336204 445278
rect 371604 445276 372204 445278
rect 407604 445276 408204 445278
rect 443604 445276 444204 445278
rect 479604 445276 480204 445278
rect 515604 445276 516204 445278
rect 551604 445276 552204 445278
rect 590960 445276 591560 445278
rect -8576 445254 592500 445276
rect -8576 445018 -7454 445254
rect -7218 445018 11786 445254
rect 12022 445018 47786 445254
rect 48022 445018 64250 445254
rect 64486 445018 299786 445254
rect 300022 445018 335786 445254
rect 336022 445018 371786 445254
rect 372022 445018 407786 445254
rect 408022 445018 443786 445254
rect 444022 445018 479786 445254
rect 480022 445018 515786 445254
rect 516022 445018 551786 445254
rect 552022 445018 591142 445254
rect 591378 445018 592500 445254
rect -8576 444934 592500 445018
rect -8576 444698 -7454 444934
rect -7218 444698 11786 444934
rect 12022 444698 47786 444934
rect 48022 444698 64250 444934
rect 64486 444698 299786 444934
rect 300022 444698 335786 444934
rect 336022 444698 371786 444934
rect 372022 444698 407786 444934
rect 408022 444698 443786 444934
rect 444022 444698 479786 444934
rect 480022 444698 515786 444934
rect 516022 444698 551786 444934
rect 552022 444698 591142 444934
rect 591378 444698 592500 444934
rect -8576 444676 592500 444698
rect -7636 444674 -7036 444676
rect 11604 444674 12204 444676
rect 47604 444674 48204 444676
rect 64208 444674 64528 444676
rect 299604 444674 300204 444676
rect 335604 444674 336204 444676
rect 371604 444674 372204 444676
rect 407604 444674 408204 444676
rect 443604 444674 444204 444676
rect 479604 444674 480204 444676
rect 515604 444674 516204 444676
rect 551604 444674 552204 444676
rect 590960 444674 591560 444676
rect -5756 441676 -5156 441678
rect 8004 441676 8604 441678
rect 44004 441676 44604 441678
rect 64208 441676 64528 441678
rect 296004 441676 296604 441678
rect 332004 441676 332604 441678
rect 368004 441676 368604 441678
rect 404004 441676 404604 441678
rect 440004 441676 440604 441678
rect 476004 441676 476604 441678
rect 512004 441676 512604 441678
rect 548004 441676 548604 441678
rect 589080 441676 589680 441678
rect -6696 441654 590620 441676
rect -6696 441418 -5574 441654
rect -5338 441418 8186 441654
rect 8422 441418 44186 441654
rect 44422 441418 64250 441654
rect 64486 441418 296186 441654
rect 296422 441418 332186 441654
rect 332422 441418 368186 441654
rect 368422 441418 404186 441654
rect 404422 441418 440186 441654
rect 440422 441418 476186 441654
rect 476422 441418 512186 441654
rect 512422 441418 548186 441654
rect 548422 441418 589262 441654
rect 589498 441418 590620 441654
rect -6696 441334 590620 441418
rect -6696 441098 -5574 441334
rect -5338 441098 8186 441334
rect 8422 441098 44186 441334
rect 44422 441098 64250 441334
rect 64486 441098 296186 441334
rect 296422 441098 332186 441334
rect 332422 441098 368186 441334
rect 368422 441098 404186 441334
rect 404422 441098 440186 441334
rect 440422 441098 476186 441334
rect 476422 441098 512186 441334
rect 512422 441098 548186 441334
rect 548422 441098 589262 441334
rect 589498 441098 590620 441334
rect -6696 441076 590620 441098
rect -5756 441074 -5156 441076
rect 8004 441074 8604 441076
rect 44004 441074 44604 441076
rect 64208 441074 64528 441076
rect 296004 441074 296604 441076
rect 332004 441074 332604 441076
rect 368004 441074 368604 441076
rect 404004 441074 404604 441076
rect 440004 441074 440604 441076
rect 476004 441074 476604 441076
rect 512004 441074 512604 441076
rect 548004 441074 548604 441076
rect 589080 441074 589680 441076
rect -3876 438076 -3276 438078
rect 4404 438076 5004 438078
rect 40404 438076 41004 438078
rect 64208 438076 64528 438078
rect 292404 438076 293004 438078
rect 328404 438076 329004 438078
rect 364404 438076 365004 438078
rect 400404 438076 401004 438078
rect 436404 438076 437004 438078
rect 472404 438076 473004 438078
rect 508404 438076 509004 438078
rect 544404 438076 545004 438078
rect 580404 438076 581004 438078
rect 587200 438076 587800 438078
rect -4816 438054 588740 438076
rect -4816 437818 -3694 438054
rect -3458 437818 4586 438054
rect 4822 437818 40586 438054
rect 40822 437818 64250 438054
rect 64486 437818 292586 438054
rect 292822 437818 328586 438054
rect 328822 437818 364586 438054
rect 364822 437818 400586 438054
rect 400822 437818 436586 438054
rect 436822 437818 472586 438054
rect 472822 437818 508586 438054
rect 508822 437818 544586 438054
rect 544822 437818 580586 438054
rect 580822 437818 587382 438054
rect 587618 437818 588740 438054
rect -4816 437734 588740 437818
rect -4816 437498 -3694 437734
rect -3458 437498 4586 437734
rect 4822 437498 40586 437734
rect 40822 437498 64250 437734
rect 64486 437498 292586 437734
rect 292822 437498 328586 437734
rect 328822 437498 364586 437734
rect 364822 437498 400586 437734
rect 400822 437498 436586 437734
rect 436822 437498 472586 437734
rect 472822 437498 508586 437734
rect 508822 437498 544586 437734
rect 544822 437498 580586 437734
rect 580822 437498 587382 437734
rect 587618 437498 588740 437734
rect -4816 437476 588740 437498
rect -3876 437474 -3276 437476
rect 4404 437474 5004 437476
rect 40404 437474 41004 437476
rect 64208 437474 64528 437476
rect 292404 437474 293004 437476
rect 328404 437474 329004 437476
rect 364404 437474 365004 437476
rect 400404 437474 401004 437476
rect 436404 437474 437004 437476
rect 472404 437474 473004 437476
rect 508404 437474 509004 437476
rect 544404 437474 545004 437476
rect 580404 437474 581004 437476
rect 587200 437474 587800 437476
rect -1996 434476 -1396 434478
rect 804 434476 1404 434478
rect 36804 434476 37404 434478
rect 64208 434476 64528 434478
rect 288804 434476 289404 434478
rect 324804 434476 325404 434478
rect 360804 434476 361404 434478
rect 396804 434476 397404 434478
rect 432804 434476 433404 434478
rect 468804 434476 469404 434478
rect 504804 434476 505404 434478
rect 540804 434476 541404 434478
rect 576804 434476 577404 434478
rect 585320 434476 585920 434478
rect -2936 434454 586860 434476
rect -2936 434218 -1814 434454
rect -1578 434218 986 434454
rect 1222 434218 36986 434454
rect 37222 434218 64250 434454
rect 64486 434218 288986 434454
rect 289222 434218 324986 434454
rect 325222 434218 360986 434454
rect 361222 434218 396986 434454
rect 397222 434218 432986 434454
rect 433222 434218 468986 434454
rect 469222 434218 504986 434454
rect 505222 434218 540986 434454
rect 541222 434218 576986 434454
rect 577222 434218 585502 434454
rect 585738 434218 586860 434454
rect -2936 434134 586860 434218
rect -2936 433898 -1814 434134
rect -1578 433898 986 434134
rect 1222 433898 36986 434134
rect 37222 433898 64250 434134
rect 64486 433898 288986 434134
rect 289222 433898 324986 434134
rect 325222 433898 360986 434134
rect 361222 433898 396986 434134
rect 397222 433898 432986 434134
rect 433222 433898 468986 434134
rect 469222 433898 504986 434134
rect 505222 433898 540986 434134
rect 541222 433898 576986 434134
rect 577222 433898 585502 434134
rect 585738 433898 586860 434134
rect -2936 433876 586860 433898
rect -1996 433874 -1396 433876
rect 804 433874 1404 433876
rect 36804 433874 37404 433876
rect 64208 433874 64528 433876
rect 288804 433874 289404 433876
rect 324804 433874 325404 433876
rect 360804 433874 361404 433876
rect 396804 433874 397404 433876
rect 432804 433874 433404 433876
rect 468804 433874 469404 433876
rect 504804 433874 505404 433876
rect 540804 433874 541404 433876
rect 576804 433874 577404 433876
rect 585320 433874 585920 433876
rect -8576 427276 -7976 427278
rect 29604 427276 30204 427278
rect 79568 427276 79888 427278
rect 317604 427276 318204 427278
rect 353604 427276 354204 427278
rect 389604 427276 390204 427278
rect 425604 427276 426204 427278
rect 461604 427276 462204 427278
rect 497604 427276 498204 427278
rect 533604 427276 534204 427278
rect 569604 427276 570204 427278
rect 591900 427276 592500 427278
rect -8576 427254 592500 427276
rect -8576 427018 -8394 427254
rect -8158 427018 29786 427254
rect 30022 427018 79610 427254
rect 79846 427018 317786 427254
rect 318022 427018 353786 427254
rect 354022 427018 389786 427254
rect 390022 427018 425786 427254
rect 426022 427018 461786 427254
rect 462022 427018 497786 427254
rect 498022 427018 533786 427254
rect 534022 427018 569786 427254
rect 570022 427018 592082 427254
rect 592318 427018 592500 427254
rect -8576 426934 592500 427018
rect -8576 426698 -8394 426934
rect -8158 426698 29786 426934
rect 30022 426698 79610 426934
rect 79846 426698 317786 426934
rect 318022 426698 353786 426934
rect 354022 426698 389786 426934
rect 390022 426698 425786 426934
rect 426022 426698 461786 426934
rect 462022 426698 497786 426934
rect 498022 426698 533786 426934
rect 534022 426698 569786 426934
rect 570022 426698 592082 426934
rect 592318 426698 592500 426934
rect -8576 426676 592500 426698
rect -8576 426674 -7976 426676
rect 29604 426674 30204 426676
rect 79568 426674 79888 426676
rect 317604 426674 318204 426676
rect 353604 426674 354204 426676
rect 389604 426674 390204 426676
rect 425604 426674 426204 426676
rect 461604 426674 462204 426676
rect 497604 426674 498204 426676
rect 533604 426674 534204 426676
rect 569604 426674 570204 426676
rect 591900 426674 592500 426676
rect -6696 423676 -6096 423678
rect 26004 423676 26604 423678
rect 79568 423676 79888 423678
rect 314004 423676 314604 423678
rect 350004 423676 350604 423678
rect 386004 423676 386604 423678
rect 422004 423676 422604 423678
rect 458004 423676 458604 423678
rect 494004 423676 494604 423678
rect 530004 423676 530604 423678
rect 566004 423676 566604 423678
rect 590020 423676 590620 423678
rect -6696 423654 590620 423676
rect -6696 423418 -6514 423654
rect -6278 423418 26186 423654
rect 26422 423418 79610 423654
rect 79846 423418 314186 423654
rect 314422 423418 350186 423654
rect 350422 423418 386186 423654
rect 386422 423418 422186 423654
rect 422422 423418 458186 423654
rect 458422 423418 494186 423654
rect 494422 423418 530186 423654
rect 530422 423418 566186 423654
rect 566422 423418 590202 423654
rect 590438 423418 590620 423654
rect -6696 423334 590620 423418
rect -6696 423098 -6514 423334
rect -6278 423098 26186 423334
rect 26422 423098 79610 423334
rect 79846 423098 314186 423334
rect 314422 423098 350186 423334
rect 350422 423098 386186 423334
rect 386422 423098 422186 423334
rect 422422 423098 458186 423334
rect 458422 423098 494186 423334
rect 494422 423098 530186 423334
rect 530422 423098 566186 423334
rect 566422 423098 590202 423334
rect 590438 423098 590620 423334
rect -6696 423076 590620 423098
rect -6696 423074 -6096 423076
rect 26004 423074 26604 423076
rect 79568 423074 79888 423076
rect 314004 423074 314604 423076
rect 350004 423074 350604 423076
rect 386004 423074 386604 423076
rect 422004 423074 422604 423076
rect 458004 423074 458604 423076
rect 494004 423074 494604 423076
rect 530004 423074 530604 423076
rect 566004 423074 566604 423076
rect 590020 423074 590620 423076
rect -4816 420076 -4216 420078
rect 22404 420076 23004 420078
rect 79568 420076 79888 420078
rect 310404 420076 311004 420078
rect 346404 420076 347004 420078
rect 382404 420076 383004 420078
rect 418404 420076 419004 420078
rect 454404 420076 455004 420078
rect 490404 420076 491004 420078
rect 526404 420076 527004 420078
rect 562404 420076 563004 420078
rect 588140 420076 588740 420078
rect -4816 420054 588740 420076
rect -4816 419818 -4634 420054
rect -4398 419818 22586 420054
rect 22822 419818 79610 420054
rect 79846 419818 310586 420054
rect 310822 419818 346586 420054
rect 346822 419818 382586 420054
rect 382822 419818 418586 420054
rect 418822 419818 454586 420054
rect 454822 419818 490586 420054
rect 490822 419818 526586 420054
rect 526822 419818 562586 420054
rect 562822 419818 588322 420054
rect 588558 419818 588740 420054
rect -4816 419734 588740 419818
rect -4816 419498 -4634 419734
rect -4398 419498 22586 419734
rect 22822 419498 79610 419734
rect 79846 419498 310586 419734
rect 310822 419498 346586 419734
rect 346822 419498 382586 419734
rect 382822 419498 418586 419734
rect 418822 419498 454586 419734
rect 454822 419498 490586 419734
rect 490822 419498 526586 419734
rect 526822 419498 562586 419734
rect 562822 419498 588322 419734
rect 588558 419498 588740 419734
rect -4816 419476 588740 419498
rect -4816 419474 -4216 419476
rect 22404 419474 23004 419476
rect 79568 419474 79888 419476
rect 310404 419474 311004 419476
rect 346404 419474 347004 419476
rect 382404 419474 383004 419476
rect 418404 419474 419004 419476
rect 454404 419474 455004 419476
rect 490404 419474 491004 419476
rect 526404 419474 527004 419476
rect 562404 419474 563004 419476
rect 588140 419474 588740 419476
rect -2936 416476 -2336 416478
rect 18804 416476 19404 416478
rect 54804 416476 55404 416478
rect 79568 416476 79888 416478
rect 306804 416476 307404 416478
rect 342804 416476 343404 416478
rect 378804 416476 379404 416478
rect 414804 416476 415404 416478
rect 450804 416476 451404 416478
rect 486804 416476 487404 416478
rect 522804 416476 523404 416478
rect 558804 416476 559404 416478
rect 586260 416476 586860 416478
rect -2936 416454 586860 416476
rect -2936 416218 -2754 416454
rect -2518 416218 18986 416454
rect 19222 416218 54986 416454
rect 55222 416218 79610 416454
rect 79846 416218 306986 416454
rect 307222 416218 342986 416454
rect 343222 416218 378986 416454
rect 379222 416218 414986 416454
rect 415222 416218 450986 416454
rect 451222 416218 486986 416454
rect 487222 416218 522986 416454
rect 523222 416218 558986 416454
rect 559222 416218 586442 416454
rect 586678 416218 586860 416454
rect -2936 416134 586860 416218
rect -2936 415898 -2754 416134
rect -2518 415898 18986 416134
rect 19222 415898 54986 416134
rect 55222 415898 79610 416134
rect 79846 415898 306986 416134
rect 307222 415898 342986 416134
rect 343222 415898 378986 416134
rect 379222 415898 414986 416134
rect 415222 415898 450986 416134
rect 451222 415898 486986 416134
rect 487222 415898 522986 416134
rect 523222 415898 558986 416134
rect 559222 415898 586442 416134
rect 586678 415898 586860 416134
rect -2936 415876 586860 415898
rect -2936 415874 -2336 415876
rect 18804 415874 19404 415876
rect 54804 415874 55404 415876
rect 79568 415874 79888 415876
rect 306804 415874 307404 415876
rect 342804 415874 343404 415876
rect 378804 415874 379404 415876
rect 414804 415874 415404 415876
rect 450804 415874 451404 415876
rect 486804 415874 487404 415876
rect 522804 415874 523404 415876
rect 558804 415874 559404 415876
rect 586260 415874 586860 415876
rect -7636 409276 -7036 409278
rect 11604 409276 12204 409278
rect 47604 409276 48204 409278
rect 64208 409276 64528 409278
rect 299604 409276 300204 409278
rect 335604 409276 336204 409278
rect 340482 409276 340802 409278
rect 443604 409276 444204 409278
rect 551604 409276 552204 409278
rect 590960 409276 591560 409278
rect -8576 409254 592500 409276
rect -8576 409018 -7454 409254
rect -7218 409018 11786 409254
rect 12022 409018 47786 409254
rect 48022 409018 64250 409254
rect 64486 409018 299786 409254
rect 300022 409018 335786 409254
rect 336022 409018 340524 409254
rect 340760 409018 443786 409254
rect 444022 409018 551786 409254
rect 552022 409018 591142 409254
rect 591378 409018 592500 409254
rect -8576 408934 592500 409018
rect -8576 408698 -7454 408934
rect -7218 408698 11786 408934
rect 12022 408698 47786 408934
rect 48022 408698 64250 408934
rect 64486 408698 299786 408934
rect 300022 408698 335786 408934
rect 336022 408698 340524 408934
rect 340760 408698 443786 408934
rect 444022 408698 551786 408934
rect 552022 408698 591142 408934
rect 591378 408698 592500 408934
rect -8576 408676 592500 408698
rect -7636 408674 -7036 408676
rect 11604 408674 12204 408676
rect 47604 408674 48204 408676
rect 64208 408674 64528 408676
rect 299604 408674 300204 408676
rect 335604 408674 336204 408676
rect 340482 408674 340802 408676
rect 443604 408674 444204 408676
rect 551604 408674 552204 408676
rect 590960 408674 591560 408676
rect -5756 405676 -5156 405678
rect 8004 405676 8604 405678
rect 44004 405676 44604 405678
rect 64208 405676 64528 405678
rect 296004 405676 296604 405678
rect 332004 405676 332604 405678
rect 340482 405676 340802 405678
rect 440004 405676 440604 405678
rect 526494 405676 526814 405678
rect 548004 405676 548604 405678
rect 589080 405676 589680 405678
rect -6696 405654 590620 405676
rect -6696 405418 -5574 405654
rect -5338 405418 8186 405654
rect 8422 405418 44186 405654
rect 44422 405418 64250 405654
rect 64486 405418 296186 405654
rect 296422 405418 332186 405654
rect 332422 405418 340524 405654
rect 340760 405418 440186 405654
rect 440422 405418 526536 405654
rect 526772 405418 548186 405654
rect 548422 405418 589262 405654
rect 589498 405418 590620 405654
rect -6696 405334 590620 405418
rect -6696 405098 -5574 405334
rect -5338 405098 8186 405334
rect 8422 405098 44186 405334
rect 44422 405098 64250 405334
rect 64486 405098 296186 405334
rect 296422 405098 332186 405334
rect 332422 405098 340524 405334
rect 340760 405098 440186 405334
rect 440422 405098 526536 405334
rect 526772 405098 548186 405334
rect 548422 405098 589262 405334
rect 589498 405098 590620 405334
rect -6696 405076 590620 405098
rect -5756 405074 -5156 405076
rect 8004 405074 8604 405076
rect 44004 405074 44604 405076
rect 64208 405074 64528 405076
rect 296004 405074 296604 405076
rect 332004 405074 332604 405076
rect 340482 405074 340802 405076
rect 440004 405074 440604 405076
rect 526494 405074 526814 405076
rect 548004 405074 548604 405076
rect 589080 405074 589680 405076
rect -3876 402076 -3276 402078
rect 4404 402076 5004 402078
rect 40404 402076 41004 402078
rect 64208 402076 64528 402078
rect 292404 402076 293004 402078
rect 328404 402076 329004 402078
rect 340482 402076 340802 402078
rect 436404 402076 437004 402078
rect 526494 402076 526814 402078
rect 544404 402076 545004 402078
rect 580404 402076 581004 402078
rect 587200 402076 587800 402078
rect -4816 402054 588740 402076
rect -4816 401818 -3694 402054
rect -3458 401818 4586 402054
rect 4822 401818 40586 402054
rect 40822 401818 64250 402054
rect 64486 401818 292586 402054
rect 292822 401818 328586 402054
rect 328822 401818 340524 402054
rect 340760 401818 436586 402054
rect 436822 401818 526536 402054
rect 526772 401818 544586 402054
rect 544822 401818 580586 402054
rect 580822 401818 587382 402054
rect 587618 401818 588740 402054
rect -4816 401734 588740 401818
rect -4816 401498 -3694 401734
rect -3458 401498 4586 401734
rect 4822 401498 40586 401734
rect 40822 401498 64250 401734
rect 64486 401498 292586 401734
rect 292822 401498 328586 401734
rect 328822 401498 340524 401734
rect 340760 401498 436586 401734
rect 436822 401498 526536 401734
rect 526772 401498 544586 401734
rect 544822 401498 580586 401734
rect 580822 401498 587382 401734
rect 587618 401498 588740 401734
rect -4816 401476 588740 401498
rect -3876 401474 -3276 401476
rect 4404 401474 5004 401476
rect 40404 401474 41004 401476
rect 64208 401474 64528 401476
rect 292404 401474 293004 401476
rect 328404 401474 329004 401476
rect 340482 401474 340802 401476
rect 436404 401474 437004 401476
rect 526494 401474 526814 401476
rect 544404 401474 545004 401476
rect 580404 401474 581004 401476
rect 587200 401474 587800 401476
rect -1996 398476 -1396 398478
rect 804 398476 1404 398478
rect 36804 398476 37404 398478
rect 64208 398476 64528 398478
rect 288804 398476 289404 398478
rect 324804 398476 325404 398478
rect 340482 398476 340802 398478
rect 432804 398476 433404 398478
rect 526494 398476 526814 398478
rect 540804 398476 541404 398478
rect 576804 398476 577404 398478
rect 585320 398476 585920 398478
rect -2936 398454 586860 398476
rect -2936 398218 -1814 398454
rect -1578 398218 986 398454
rect 1222 398218 36986 398454
rect 37222 398218 64250 398454
rect 64486 398218 288986 398454
rect 289222 398218 324986 398454
rect 325222 398218 340524 398454
rect 340760 398218 432986 398454
rect 433222 398218 526536 398454
rect 526772 398218 540986 398454
rect 541222 398218 576986 398454
rect 577222 398218 585502 398454
rect 585738 398218 586860 398454
rect -2936 398134 586860 398218
rect -2936 397898 -1814 398134
rect -1578 397898 986 398134
rect 1222 397898 36986 398134
rect 37222 397898 64250 398134
rect 64486 397898 288986 398134
rect 289222 397898 324986 398134
rect 325222 397898 340524 398134
rect 340760 397898 432986 398134
rect 433222 397898 526536 398134
rect 526772 397898 540986 398134
rect 541222 397898 576986 398134
rect 577222 397898 585502 398134
rect 585738 397898 586860 398134
rect -2936 397876 586860 397898
rect -1996 397874 -1396 397876
rect 804 397874 1404 397876
rect 36804 397874 37404 397876
rect 64208 397874 64528 397876
rect 288804 397874 289404 397876
rect 324804 397874 325404 397876
rect 340482 397874 340802 397876
rect 432804 397874 433404 397876
rect 526494 397874 526814 397876
rect 540804 397874 541404 397876
rect 576804 397874 577404 397876
rect 585320 397874 585920 397876
rect -8576 391276 -7976 391278
rect 29604 391276 30204 391278
rect 79568 391276 79888 391278
rect 317604 391276 318204 391278
rect 340034 391276 340358 391278
rect 425604 391276 426204 391278
rect 526938 391276 527262 391278
rect 533604 391276 534204 391278
rect 569604 391276 570204 391278
rect 591900 391276 592500 391278
rect -8576 391254 592500 391276
rect -8576 391018 -8394 391254
rect -8158 391018 29786 391254
rect 30022 391018 79610 391254
rect 79846 391018 317786 391254
rect 318022 391018 340078 391254
rect 340314 391018 425786 391254
rect 426022 391018 526982 391254
rect 527218 391018 533786 391254
rect 534022 391018 569786 391254
rect 570022 391018 592082 391254
rect 592318 391018 592500 391254
rect -8576 390934 592500 391018
rect -8576 390698 -8394 390934
rect -8158 390698 29786 390934
rect 30022 390698 79610 390934
rect 79846 390698 317786 390934
rect 318022 390698 340078 390934
rect 340314 390698 425786 390934
rect 426022 390698 526982 390934
rect 527218 390698 533786 390934
rect 534022 390698 569786 390934
rect 570022 390698 592082 390934
rect 592318 390698 592500 390934
rect -8576 390676 592500 390698
rect -8576 390674 -7976 390676
rect 29604 390674 30204 390676
rect 79568 390674 79888 390676
rect 317604 390674 318204 390676
rect 340034 390674 340358 390676
rect 425604 390674 426204 390676
rect 526938 390674 527262 390676
rect 533604 390674 534204 390676
rect 569604 390674 570204 390676
rect 591900 390674 592500 390676
rect -6696 387676 -6096 387678
rect 26004 387676 26604 387678
rect 79568 387676 79888 387678
rect 314004 387676 314604 387678
rect 340034 387676 340358 387678
rect 422004 387676 422604 387678
rect 526938 387676 527262 387678
rect 566004 387676 566604 387678
rect 590020 387676 590620 387678
rect -6696 387654 590620 387676
rect -6696 387418 -6514 387654
rect -6278 387418 26186 387654
rect 26422 387418 79610 387654
rect 79846 387418 314186 387654
rect 314422 387418 340078 387654
rect 340314 387418 422186 387654
rect 422422 387418 526982 387654
rect 527218 387418 566186 387654
rect 566422 387418 590202 387654
rect 590438 387418 590620 387654
rect -6696 387334 590620 387418
rect -6696 387098 -6514 387334
rect -6278 387098 26186 387334
rect 26422 387098 79610 387334
rect 79846 387098 314186 387334
rect 314422 387098 340078 387334
rect 340314 387098 422186 387334
rect 422422 387098 526982 387334
rect 527218 387098 566186 387334
rect 566422 387098 590202 387334
rect 590438 387098 590620 387334
rect -6696 387076 590620 387098
rect -6696 387074 -6096 387076
rect 26004 387074 26604 387076
rect 79568 387074 79888 387076
rect 314004 387074 314604 387076
rect 340034 387074 340358 387076
rect 422004 387074 422604 387076
rect 526938 387074 527262 387076
rect 566004 387074 566604 387076
rect 590020 387074 590620 387076
rect -4816 384076 -4216 384078
rect 22404 384076 23004 384078
rect 79568 384076 79888 384078
rect 310404 384076 311004 384078
rect 340034 384076 340358 384078
rect 526938 384076 527262 384078
rect 562404 384076 563004 384078
rect 588140 384076 588740 384078
rect -4816 384054 588740 384076
rect -4816 383818 -4634 384054
rect -4398 383818 22586 384054
rect 22822 383818 79610 384054
rect 79846 383818 310586 384054
rect 310822 383818 340078 384054
rect 340314 383818 526982 384054
rect 527218 383818 562586 384054
rect 562822 383818 588322 384054
rect 588558 383818 588740 384054
rect -4816 383734 588740 383818
rect -4816 383498 -4634 383734
rect -4398 383498 22586 383734
rect 22822 383498 79610 383734
rect 79846 383498 310586 383734
rect 310822 383498 340078 383734
rect 340314 383498 526982 383734
rect 527218 383498 562586 383734
rect 562822 383498 588322 383734
rect 588558 383498 588740 383734
rect -4816 383476 588740 383498
rect -4816 383474 -4216 383476
rect 22404 383474 23004 383476
rect 79568 383474 79888 383476
rect 310404 383474 311004 383476
rect 340034 383474 340358 383476
rect 526938 383474 527262 383476
rect 562404 383474 563004 383476
rect 588140 383474 588740 383476
rect -2936 380476 -2336 380478
rect 18804 380476 19404 380478
rect 54804 380476 55404 380478
rect 79568 380476 79888 380478
rect 306804 380476 307404 380478
rect 340034 380476 340358 380478
rect 526938 380476 527262 380478
rect 558804 380476 559404 380478
rect 586260 380476 586860 380478
rect -2936 380454 586860 380476
rect -2936 380218 -2754 380454
rect -2518 380218 18986 380454
rect 19222 380218 54986 380454
rect 55222 380218 79610 380454
rect 79846 380218 306986 380454
rect 307222 380218 340078 380454
rect 340314 380218 526982 380454
rect 527218 380218 558986 380454
rect 559222 380218 586442 380454
rect 586678 380218 586860 380454
rect -2936 380134 586860 380218
rect -2936 379898 -2754 380134
rect -2518 379898 18986 380134
rect 19222 379898 54986 380134
rect 55222 379898 79610 380134
rect 79846 379898 306986 380134
rect 307222 379898 340078 380134
rect 340314 379898 526982 380134
rect 527218 379898 558986 380134
rect 559222 379898 586442 380134
rect 586678 379898 586860 380134
rect -2936 379876 586860 379898
rect -2936 379874 -2336 379876
rect 18804 379874 19404 379876
rect 54804 379874 55404 379876
rect 79568 379874 79888 379876
rect 306804 379874 307404 379876
rect 340034 379874 340358 379876
rect 526938 379874 527262 379876
rect 558804 379874 559404 379876
rect 586260 379874 586860 379876
rect -7636 373276 -7036 373278
rect 11604 373276 12204 373278
rect 47604 373276 48204 373278
rect 64208 373276 64528 373278
rect 299604 373276 300204 373278
rect 335604 373276 336204 373278
rect 340482 373276 340802 373278
rect 443604 373276 444204 373278
rect 526494 373276 526814 373278
rect 551604 373276 552204 373278
rect 590960 373276 591560 373278
rect -8576 373254 592500 373276
rect -8576 373018 -7454 373254
rect -7218 373018 11786 373254
rect 12022 373018 47786 373254
rect 48022 373018 64250 373254
rect 64486 373018 299786 373254
rect 300022 373018 335786 373254
rect 336022 373018 340524 373254
rect 340760 373018 443786 373254
rect 444022 373018 526536 373254
rect 526772 373018 551786 373254
rect 552022 373018 591142 373254
rect 591378 373018 592500 373254
rect -8576 372934 592500 373018
rect -8576 372698 -7454 372934
rect -7218 372698 11786 372934
rect 12022 372698 47786 372934
rect 48022 372698 64250 372934
rect 64486 372698 299786 372934
rect 300022 372698 335786 372934
rect 336022 372698 340524 372934
rect 340760 372698 443786 372934
rect 444022 372698 526536 372934
rect 526772 372698 551786 372934
rect 552022 372698 591142 372934
rect 591378 372698 592500 372934
rect -8576 372676 592500 372698
rect -7636 372674 -7036 372676
rect 11604 372674 12204 372676
rect 47604 372674 48204 372676
rect 64208 372674 64528 372676
rect 299604 372674 300204 372676
rect 335604 372674 336204 372676
rect 340482 372674 340802 372676
rect 443604 372674 444204 372676
rect 526494 372674 526814 372676
rect 551604 372674 552204 372676
rect 590960 372674 591560 372676
rect -5756 369676 -5156 369678
rect 8004 369676 8604 369678
rect 44004 369676 44604 369678
rect 64208 369676 64528 369678
rect 296004 369676 296604 369678
rect 332004 369676 332604 369678
rect 340482 369676 340802 369678
rect 440004 369676 440604 369678
rect 526494 369676 526814 369678
rect 548004 369676 548604 369678
rect 589080 369676 589680 369678
rect -6696 369654 590620 369676
rect -6696 369418 -5574 369654
rect -5338 369418 8186 369654
rect 8422 369418 44186 369654
rect 44422 369418 64250 369654
rect 64486 369418 296186 369654
rect 296422 369418 332186 369654
rect 332422 369418 340524 369654
rect 340760 369418 440186 369654
rect 440422 369418 526536 369654
rect 526772 369418 548186 369654
rect 548422 369418 589262 369654
rect 589498 369418 590620 369654
rect -6696 369334 590620 369418
rect -6696 369098 -5574 369334
rect -5338 369098 8186 369334
rect 8422 369098 44186 369334
rect 44422 369098 64250 369334
rect 64486 369098 296186 369334
rect 296422 369098 332186 369334
rect 332422 369098 340524 369334
rect 340760 369098 440186 369334
rect 440422 369098 526536 369334
rect 526772 369098 548186 369334
rect 548422 369098 589262 369334
rect 589498 369098 590620 369334
rect -6696 369076 590620 369098
rect -5756 369074 -5156 369076
rect 8004 369074 8604 369076
rect 44004 369074 44604 369076
rect 64208 369074 64528 369076
rect 296004 369074 296604 369076
rect 332004 369074 332604 369076
rect 340482 369074 340802 369076
rect 440004 369074 440604 369076
rect 526494 369074 526814 369076
rect 548004 369074 548604 369076
rect 589080 369074 589680 369076
rect -3876 366076 -3276 366078
rect 4404 366076 5004 366078
rect 40404 366076 41004 366078
rect 64208 366076 64528 366078
rect 292404 366076 293004 366078
rect 328404 366076 329004 366078
rect 340482 366076 340802 366078
rect 436404 366076 437004 366078
rect 526494 366076 526814 366078
rect 544404 366076 545004 366078
rect 580404 366076 581004 366078
rect 587200 366076 587800 366078
rect -4816 366054 588740 366076
rect -4816 365818 -3694 366054
rect -3458 365818 4586 366054
rect 4822 365818 40586 366054
rect 40822 365818 64250 366054
rect 64486 365818 292586 366054
rect 292822 365818 328586 366054
rect 328822 365818 340524 366054
rect 340760 365818 436586 366054
rect 436822 365818 526536 366054
rect 526772 365818 544586 366054
rect 544822 365818 580586 366054
rect 580822 365818 587382 366054
rect 587618 365818 588740 366054
rect -4816 365734 588740 365818
rect -4816 365498 -3694 365734
rect -3458 365498 4586 365734
rect 4822 365498 40586 365734
rect 40822 365498 64250 365734
rect 64486 365498 292586 365734
rect 292822 365498 328586 365734
rect 328822 365498 340524 365734
rect 340760 365498 436586 365734
rect 436822 365498 526536 365734
rect 526772 365498 544586 365734
rect 544822 365498 580586 365734
rect 580822 365498 587382 365734
rect 587618 365498 588740 365734
rect -4816 365476 588740 365498
rect -3876 365474 -3276 365476
rect 4404 365474 5004 365476
rect 40404 365474 41004 365476
rect 64208 365474 64528 365476
rect 292404 365474 293004 365476
rect 328404 365474 329004 365476
rect 340482 365474 340802 365476
rect 436404 365474 437004 365476
rect 526494 365474 526814 365476
rect 544404 365474 545004 365476
rect 580404 365474 581004 365476
rect 587200 365474 587800 365476
rect -1996 362476 -1396 362478
rect 804 362476 1404 362478
rect 36804 362476 37404 362478
rect 64208 362476 64528 362478
rect 288804 362476 289404 362478
rect 324804 362476 325404 362478
rect 340482 362476 340802 362478
rect 432804 362476 433404 362478
rect 526494 362476 526814 362478
rect 540804 362476 541404 362478
rect 576804 362476 577404 362478
rect 585320 362476 585920 362478
rect -2936 362454 586860 362476
rect -2936 362218 -1814 362454
rect -1578 362218 986 362454
rect 1222 362218 36986 362454
rect 37222 362218 64250 362454
rect 64486 362218 288986 362454
rect 289222 362218 324986 362454
rect 325222 362218 340524 362454
rect 340760 362218 432986 362454
rect 433222 362218 526536 362454
rect 526772 362218 540986 362454
rect 541222 362218 576986 362454
rect 577222 362218 585502 362454
rect 585738 362218 586860 362454
rect -2936 362134 586860 362218
rect -2936 361898 -1814 362134
rect -1578 361898 986 362134
rect 1222 361898 36986 362134
rect 37222 361898 64250 362134
rect 64486 361898 288986 362134
rect 289222 361898 324986 362134
rect 325222 361898 340524 362134
rect 340760 361898 432986 362134
rect 433222 361898 526536 362134
rect 526772 361898 540986 362134
rect 541222 361898 576986 362134
rect 577222 361898 585502 362134
rect 585738 361898 586860 362134
rect -2936 361876 586860 361898
rect -1996 361874 -1396 361876
rect 804 361874 1404 361876
rect 36804 361874 37404 361876
rect 64208 361874 64528 361876
rect 288804 361874 289404 361876
rect 324804 361874 325404 361876
rect 340482 361874 340802 361876
rect 432804 361874 433404 361876
rect 526494 361874 526814 361876
rect 540804 361874 541404 361876
rect 576804 361874 577404 361876
rect 585320 361874 585920 361876
rect -8576 355276 -7976 355278
rect 29604 355276 30204 355278
rect 79568 355276 79888 355278
rect 317604 355276 318204 355278
rect 340034 355276 340358 355278
rect 425604 355276 426204 355278
rect 526938 355276 527262 355278
rect 533604 355276 534204 355278
rect 569604 355276 570204 355278
rect 591900 355276 592500 355278
rect -8576 355254 592500 355276
rect -8576 355018 -8394 355254
rect -8158 355018 29786 355254
rect 30022 355018 79610 355254
rect 79846 355018 317786 355254
rect 318022 355018 340078 355254
rect 340314 355018 425786 355254
rect 426022 355018 526982 355254
rect 527218 355018 533786 355254
rect 534022 355018 569786 355254
rect 570022 355018 592082 355254
rect 592318 355018 592500 355254
rect -8576 354934 592500 355018
rect -8576 354698 -8394 354934
rect -8158 354698 29786 354934
rect 30022 354698 79610 354934
rect 79846 354698 317786 354934
rect 318022 354698 340078 354934
rect 340314 354698 425786 354934
rect 426022 354698 526982 354934
rect 527218 354698 533786 354934
rect 534022 354698 569786 354934
rect 570022 354698 592082 354934
rect 592318 354698 592500 354934
rect -8576 354676 592500 354698
rect -8576 354674 -7976 354676
rect 29604 354674 30204 354676
rect 79568 354674 79888 354676
rect 317604 354674 318204 354676
rect 340034 354674 340358 354676
rect 425604 354674 426204 354676
rect 526938 354674 527262 354676
rect 533604 354674 534204 354676
rect 569604 354674 570204 354676
rect 591900 354674 592500 354676
rect -6696 351676 -6096 351678
rect 26004 351676 26604 351678
rect 79568 351676 79888 351678
rect 314004 351676 314604 351678
rect 340034 351676 340358 351678
rect 422004 351676 422604 351678
rect 526938 351676 527262 351678
rect 566004 351676 566604 351678
rect 590020 351676 590620 351678
rect -6696 351654 590620 351676
rect -6696 351418 -6514 351654
rect -6278 351418 26186 351654
rect 26422 351418 79610 351654
rect 79846 351418 314186 351654
rect 314422 351418 340078 351654
rect 340314 351418 422186 351654
rect 422422 351418 526982 351654
rect 527218 351418 566186 351654
rect 566422 351418 590202 351654
rect 590438 351418 590620 351654
rect -6696 351334 590620 351418
rect -6696 351098 -6514 351334
rect -6278 351098 26186 351334
rect 26422 351098 79610 351334
rect 79846 351098 314186 351334
rect 314422 351098 340078 351334
rect 340314 351098 422186 351334
rect 422422 351098 526982 351334
rect 527218 351098 566186 351334
rect 566422 351098 590202 351334
rect 590438 351098 590620 351334
rect -6696 351076 590620 351098
rect -6696 351074 -6096 351076
rect 26004 351074 26604 351076
rect 79568 351074 79888 351076
rect 314004 351074 314604 351076
rect 340034 351074 340358 351076
rect 422004 351074 422604 351076
rect 526938 351074 527262 351076
rect 566004 351074 566604 351076
rect 590020 351074 590620 351076
rect 420556 349298 527780 349340
rect 420556 349062 420598 349298
rect 420834 349062 527502 349298
rect 527738 349062 527780 349298
rect 420556 349020 527780 349062
rect -4816 348076 -4216 348078
rect 22404 348076 23004 348078
rect 79568 348076 79888 348078
rect 310404 348076 311004 348078
rect 340034 348076 340358 348078
rect 526938 348076 527262 348078
rect 562404 348076 563004 348078
rect 588140 348076 588740 348078
rect -4816 348054 588740 348076
rect -4816 347818 -4634 348054
rect -4398 347818 22586 348054
rect 22822 347818 79610 348054
rect 79846 347818 310586 348054
rect 310822 347818 340078 348054
rect 340314 347818 526982 348054
rect 527218 347818 562586 348054
rect 562822 347818 588322 348054
rect 588558 347818 588740 348054
rect -4816 347734 588740 347818
rect -4816 347498 -4634 347734
rect -4398 347498 22586 347734
rect 22822 347498 79610 347734
rect 79846 347498 310586 347734
rect 310822 347498 340078 347734
rect 340314 347498 526982 347734
rect 527218 347498 562586 347734
rect 562822 347498 588322 347734
rect 588558 347498 588740 347734
rect -4816 347476 588740 347498
rect -4816 347474 -4216 347476
rect 22404 347474 23004 347476
rect 79568 347474 79888 347476
rect 310404 347474 311004 347476
rect 340034 347474 340358 347476
rect 526938 347474 527262 347476
rect 562404 347474 563004 347476
rect 588140 347474 588740 347476
rect 419820 346578 420140 346620
rect 419820 346342 419862 346578
rect 420098 346342 420140 346578
rect 419820 345940 420140 346342
rect 420556 346578 423084 346620
rect 420556 346342 420598 346578
rect 420834 346342 422806 346578
rect 423042 346342 423084 346578
rect 420556 346300 423084 346342
rect 427732 346578 447004 346620
rect 427732 346342 427774 346578
rect 428010 346342 446726 346578
rect 446962 346342 447004 346578
rect 427732 346300 447004 346342
rect 447604 346578 528148 346620
rect 447604 346342 447646 346578
rect 447882 346342 527870 346578
rect 528106 346342 528148 346578
rect 447604 346300 528148 346342
rect 419820 345898 438172 345940
rect 419820 345662 437894 345898
rect 438130 345662 438172 345898
rect 419820 345620 438172 345662
rect 447052 345898 527780 345940
rect 447052 345662 447094 345898
rect 447330 345662 527502 345898
rect 527738 345662 527780 345898
rect 447052 345620 527780 345662
rect 437668 345218 527780 345260
rect 437668 344982 437710 345218
rect 437946 344982 527502 345218
rect 527738 344982 527780 345218
rect 437668 344940 527780 344982
rect -2936 344476 -2336 344478
rect 18804 344476 19404 344478
rect 54804 344476 55404 344478
rect 79568 344476 79888 344478
rect 306804 344476 307404 344478
rect 340034 344476 340358 344478
rect 526938 344476 527262 344478
rect 558804 344476 559404 344478
rect 586260 344476 586860 344478
rect -2936 344454 586860 344476
rect -2936 344218 -2754 344454
rect -2518 344218 18986 344454
rect 19222 344218 54986 344454
rect 55222 344218 79610 344454
rect 79846 344218 306986 344454
rect 307222 344218 340078 344454
rect 340314 344218 526982 344454
rect 527218 344218 558986 344454
rect 559222 344218 586442 344454
rect 586678 344218 586860 344454
rect -2936 344134 586860 344218
rect -2936 343898 -2754 344134
rect -2518 343898 18986 344134
rect 19222 343898 54986 344134
rect 55222 343898 79610 344134
rect 79846 343898 306986 344134
rect 307222 343898 340078 344134
rect 340314 343898 526982 344134
rect 527218 343898 558986 344134
rect 559222 343898 586442 344134
rect 586678 343898 586860 344134
rect -2936 343876 586860 343898
rect -2936 343874 -2336 343876
rect 18804 343874 19404 343876
rect 54804 343874 55404 343876
rect 79568 343874 79888 343876
rect 306804 343874 307404 343876
rect 340034 343874 340358 343876
rect 526938 343874 527262 343876
rect 558804 343874 559404 343876
rect 586260 343874 586860 343876
rect 420556 343178 437804 343220
rect 420556 342942 420598 343178
rect 420834 342942 437526 343178
rect 437762 342942 437804 343178
rect 420556 342900 437804 342942
rect 447972 343178 449764 343220
rect 447972 342942 448014 343178
rect 448250 342942 449486 343178
rect 449722 342942 449764 343178
rect 447972 342900 449764 342942
rect 453492 342900 469820 343220
rect 453492 342540 453812 342900
rect 445396 342498 453812 342540
rect 445396 342262 445438 342498
rect 445674 342262 453812 342498
rect 445396 342220 453812 342262
rect 469500 342540 469820 342900
rect 478884 342900 486012 343220
rect 478884 342540 479204 342900
rect 469500 342220 471292 342540
rect 470972 341860 471292 342220
rect 471892 342220 479204 342540
rect 485692 342540 486012 342900
rect 488636 342900 502572 343220
rect 488636 342540 488956 342900
rect 502252 342540 502572 342900
rect 521388 343178 527780 343220
rect 521388 342942 527502 343178
rect 527738 342942 527780 343178
rect 521388 342900 527780 342942
rect 485692 342220 488956 342540
rect 495076 342220 498156 342540
rect 502252 342220 515452 342540
rect 471892 341860 472212 342220
rect 420372 341818 444612 341860
rect 420372 341582 420414 341818
rect 420650 341582 444334 341818
rect 444570 341582 444612 341818
rect 420372 341540 444612 341582
rect 445028 341818 450132 341860
rect 445028 341582 445070 341818
rect 445306 341582 450132 341818
rect 445028 341540 450132 341582
rect 449812 341180 450132 341540
rect 460300 341540 470556 341860
rect 470972 341540 472212 341860
rect 472628 341540 477732 341860
rect 460300 341180 460620 341540
rect 420372 341138 428052 341180
rect 420372 340902 420414 341138
rect 420650 340902 427774 341138
rect 428010 340902 428052 341138
rect 420372 340860 428052 340902
rect 444108 340458 444612 341180
rect 449812 340860 459516 341180
rect 444108 340222 444334 340458
rect 444570 340222 444612 340458
rect 444108 340180 444612 340222
rect 459196 340500 459516 340860
rect 460116 340860 460620 341180
rect 470236 341180 470556 341540
rect 472628 341180 472948 341540
rect 470236 340860 472948 341180
rect 460116 340500 460436 340860
rect 477412 340500 477732 341540
rect 495076 341180 495396 342220
rect 497836 341860 498156 342220
rect 515132 341860 515452 342220
rect 521388 341860 521708 342900
rect 497836 341540 508092 341860
rect 515132 341540 521708 341860
rect 522124 341818 527780 341860
rect 522124 341582 527502 341818
rect 527738 341582 527780 341818
rect 522124 341540 527780 341582
rect 486244 340860 495396 341180
rect 486244 340500 486564 340860
rect 459196 340180 460436 340500
rect 467844 340180 469820 340500
rect 477412 340180 486564 340500
rect 507772 340500 508092 341540
rect 522124 341180 522444 341540
rect 521940 340860 522444 341180
rect 507772 340180 514900 340500
rect 444108 339820 444428 340180
rect 439324 339778 444428 339820
rect 439324 339542 439366 339778
rect 439602 339542 444428 339778
rect 439324 339500 444428 339542
rect 459196 338820 459700 340180
rect 467844 339820 468164 340180
rect 464164 339500 468164 339820
rect 464164 338460 464484 339500
rect 469500 339140 469820 340180
rect 514580 339820 514900 340180
rect 521940 339820 522260 340860
rect 486980 339500 497420 339820
rect 486980 339140 487300 339500
rect 469500 338820 470004 339140
rect 450548 338418 464484 338460
rect 450548 338182 450590 338418
rect 450826 338182 464484 338418
rect 450548 338140 464484 338182
rect 469684 338460 470004 338820
rect 478148 338820 487300 339140
rect 478148 338460 478468 338820
rect 469684 338140 478468 338460
rect 497100 338460 497420 339500
rect 497836 339500 506988 339820
rect 514580 339500 522260 339820
rect 522860 340458 528148 340500
rect 522860 340222 527870 340458
rect 528106 340222 528148 340458
rect 522860 340180 528148 340222
rect 497836 338460 498156 339500
rect 506668 339140 506988 339500
rect 506668 338820 507540 339140
rect 497100 338140 498156 338460
rect 507220 338460 507540 338820
rect 507956 338820 509932 339140
rect 507956 338460 508276 338820
rect 507220 338140 508276 338460
rect 509612 338460 509932 338820
rect 522860 338460 523180 340180
rect 509612 338140 523180 338460
rect -7636 337276 -7036 337278
rect 11604 337276 12204 337278
rect 47604 337276 48204 337278
rect 64208 337276 64528 337278
rect 299604 337276 300204 337278
rect 335604 337276 336204 337278
rect 340482 337276 340802 337278
rect 443604 337276 444204 337278
rect 526494 337276 526814 337278
rect 551604 337276 552204 337278
rect 590960 337276 591560 337278
rect -8576 337254 592500 337276
rect -8576 337018 -7454 337254
rect -7218 337018 11786 337254
rect 12022 337018 47786 337254
rect 48022 337018 64250 337254
rect 64486 337018 299786 337254
rect 300022 337018 335786 337254
rect 336022 337018 340524 337254
rect 340760 337018 443786 337254
rect 444022 337018 526536 337254
rect 526772 337018 551786 337254
rect 552022 337018 591142 337254
rect 591378 337018 592500 337254
rect -8576 336934 592500 337018
rect -8576 336698 -7454 336934
rect -7218 336698 11786 336934
rect 12022 336698 47786 336934
rect 48022 336698 64250 336934
rect 64486 336698 299786 336934
rect 300022 336698 335786 336934
rect 336022 336698 340524 336934
rect 340760 336698 443786 336934
rect 444022 336698 526536 336934
rect 526772 336698 551786 336934
rect 552022 336698 591142 336934
rect 591378 336698 592500 336934
rect -8576 336676 592500 336698
rect -7636 336674 -7036 336676
rect 11604 336674 12204 336676
rect 47604 336674 48204 336676
rect 64208 336674 64528 336676
rect 299604 336674 300204 336676
rect 335604 336674 336204 336676
rect 340482 336674 340802 336676
rect 443604 336674 444204 336676
rect 526494 336674 526814 336676
rect 551604 336674 552204 336676
rect 590960 336674 591560 336676
rect -5756 333676 -5156 333678
rect 8004 333676 8604 333678
rect 44004 333676 44604 333678
rect 64208 333676 64528 333678
rect 296004 333676 296604 333678
rect 332004 333676 332604 333678
rect 340482 333676 340802 333678
rect 440004 333676 440604 333678
rect 526494 333676 526814 333678
rect 548004 333676 548604 333678
rect 589080 333676 589680 333678
rect -6696 333654 590620 333676
rect -6696 333418 -5574 333654
rect -5338 333418 8186 333654
rect 8422 333418 44186 333654
rect 44422 333418 64250 333654
rect 64486 333418 296186 333654
rect 296422 333418 332186 333654
rect 332422 333418 340524 333654
rect 340760 333418 440186 333654
rect 440422 333418 526536 333654
rect 526772 333418 548186 333654
rect 548422 333418 589262 333654
rect 589498 333418 590620 333654
rect -6696 333334 590620 333418
rect -6696 333098 -5574 333334
rect -5338 333098 8186 333334
rect 8422 333098 44186 333334
rect 44422 333098 64250 333334
rect 64486 333098 296186 333334
rect 296422 333098 332186 333334
rect 332422 333098 340524 333334
rect 340760 333098 440186 333334
rect 440422 333098 526536 333334
rect 526772 333098 548186 333334
rect 548422 333098 589262 333334
rect 589498 333098 590620 333334
rect -6696 333076 590620 333098
rect -5756 333074 -5156 333076
rect 8004 333074 8604 333076
rect 44004 333074 44604 333076
rect 64208 333074 64528 333076
rect 296004 333074 296604 333076
rect 332004 333074 332604 333076
rect 340482 333074 340802 333076
rect 440004 333074 440604 333076
rect 526494 333074 526814 333076
rect 548004 333074 548604 333076
rect 589080 333074 589680 333076
rect -3876 330076 -3276 330078
rect 4404 330076 5004 330078
rect 40404 330076 41004 330078
rect 64208 330076 64528 330078
rect 292404 330076 293004 330078
rect 328404 330076 329004 330078
rect 340482 330076 340802 330078
rect 436404 330076 437004 330078
rect 526494 330076 526814 330078
rect 544404 330076 545004 330078
rect 580404 330076 581004 330078
rect 587200 330076 587800 330078
rect -4816 330054 588740 330076
rect -4816 329818 -3694 330054
rect -3458 329818 4586 330054
rect 4822 329818 40586 330054
rect 40822 329818 64250 330054
rect 64486 329818 292586 330054
rect 292822 329818 328586 330054
rect 328822 329818 340524 330054
rect 340760 329818 436586 330054
rect 436822 329818 526536 330054
rect 526772 329818 544586 330054
rect 544822 329818 580586 330054
rect 580822 329818 587382 330054
rect 587618 329818 588740 330054
rect -4816 329734 588740 329818
rect -4816 329498 -3694 329734
rect -3458 329498 4586 329734
rect 4822 329498 40586 329734
rect 40822 329498 64250 329734
rect 64486 329498 292586 329734
rect 292822 329498 328586 329734
rect 328822 329498 340524 329734
rect 340760 329498 436586 329734
rect 436822 329498 526536 329734
rect 526772 329498 544586 329734
rect 544822 329498 580586 329734
rect 580822 329498 587382 329734
rect 587618 329498 588740 329734
rect -4816 329476 588740 329498
rect -3876 329474 -3276 329476
rect 4404 329474 5004 329476
rect 40404 329474 41004 329476
rect 64208 329474 64528 329476
rect 292404 329474 293004 329476
rect 328404 329474 329004 329476
rect 340482 329474 340802 329476
rect 436404 329474 437004 329476
rect 526494 329474 526814 329476
rect 544404 329474 545004 329476
rect 580404 329474 581004 329476
rect 587200 329474 587800 329476
rect -1996 326476 -1396 326478
rect 804 326476 1404 326478
rect 36804 326476 37404 326478
rect 64208 326476 64528 326478
rect 288804 326476 289404 326478
rect 324804 326476 325404 326478
rect 340482 326476 340802 326478
rect 432804 326476 433404 326478
rect 526494 326476 526814 326478
rect 540804 326476 541404 326478
rect 576804 326476 577404 326478
rect 585320 326476 585920 326478
rect -2936 326454 586860 326476
rect -2936 326218 -1814 326454
rect -1578 326218 986 326454
rect 1222 326218 36986 326454
rect 37222 326218 64250 326454
rect 64486 326218 288986 326454
rect 289222 326218 324986 326454
rect 325222 326218 340524 326454
rect 340760 326218 432986 326454
rect 433222 326218 526536 326454
rect 526772 326218 540986 326454
rect 541222 326218 576986 326454
rect 577222 326218 585502 326454
rect 585738 326218 586860 326454
rect -2936 326134 586860 326218
rect -2936 325898 -1814 326134
rect -1578 325898 986 326134
rect 1222 325898 36986 326134
rect 37222 325898 64250 326134
rect 64486 325898 288986 326134
rect 289222 325898 324986 326134
rect 325222 325898 340524 326134
rect 340760 325898 432986 326134
rect 433222 325898 526536 326134
rect 526772 325898 540986 326134
rect 541222 325898 576986 326134
rect 577222 325898 585502 326134
rect 585738 325898 586860 326134
rect -2936 325876 586860 325898
rect -1996 325874 -1396 325876
rect 804 325874 1404 325876
rect 36804 325874 37404 325876
rect 64208 325874 64528 325876
rect 288804 325874 289404 325876
rect 324804 325874 325404 325876
rect 340482 325874 340802 325876
rect 432804 325874 433404 325876
rect 526494 325874 526814 325876
rect 540804 325874 541404 325876
rect 576804 325874 577404 325876
rect 585320 325874 585920 325876
rect -8576 319276 -7976 319278
rect 29604 319276 30204 319278
rect 317604 319276 318204 319278
rect 425604 319276 426204 319278
rect 533604 319276 534204 319278
rect 569604 319276 570204 319278
rect 591900 319276 592500 319278
rect -8576 319254 592500 319276
rect -8576 319018 -8394 319254
rect -8158 319018 29786 319254
rect 30022 319018 317786 319254
rect 318022 319018 425786 319254
rect 426022 319018 533786 319254
rect 534022 319018 569786 319254
rect 570022 319018 592082 319254
rect 592318 319018 592500 319254
rect -8576 318934 592500 319018
rect -8576 318698 -8394 318934
rect -8158 318698 29786 318934
rect 30022 318698 317786 318934
rect 318022 318698 425786 318934
rect 426022 318698 533786 318934
rect 534022 318698 569786 318934
rect 570022 318698 592082 318934
rect 592318 318698 592500 318934
rect -8576 318676 592500 318698
rect -8576 318674 -7976 318676
rect 29604 318674 30204 318676
rect 317604 318674 318204 318676
rect 425604 318674 426204 318676
rect 533604 318674 534204 318676
rect 569604 318674 570204 318676
rect 591900 318674 592500 318676
rect -6696 315676 -6096 315678
rect 26004 315676 26604 315678
rect 62004 315676 62604 315678
rect 98004 315676 98604 315678
rect 134004 315676 134604 315678
rect 170004 315676 170604 315678
rect 206004 315676 206604 315678
rect 242004 315676 242604 315678
rect 278004 315676 278604 315678
rect 314004 315676 314604 315678
rect 350004 315676 350604 315678
rect 386004 315676 386604 315678
rect 422004 315676 422604 315678
rect 458004 315676 458604 315678
rect 494004 315676 494604 315678
rect 530004 315676 530604 315678
rect 566004 315676 566604 315678
rect 590020 315676 590620 315678
rect -6696 315654 590620 315676
rect -6696 315418 -6514 315654
rect -6278 315418 26186 315654
rect 26422 315418 62186 315654
rect 62422 315418 98186 315654
rect 98422 315418 134186 315654
rect 134422 315418 170186 315654
rect 170422 315418 206186 315654
rect 206422 315418 242186 315654
rect 242422 315418 278186 315654
rect 278422 315418 314186 315654
rect 314422 315418 350186 315654
rect 350422 315418 386186 315654
rect 386422 315418 422186 315654
rect 422422 315418 458186 315654
rect 458422 315418 494186 315654
rect 494422 315418 530186 315654
rect 530422 315418 566186 315654
rect 566422 315418 590202 315654
rect 590438 315418 590620 315654
rect -6696 315334 590620 315418
rect -6696 315098 -6514 315334
rect -6278 315098 26186 315334
rect 26422 315098 62186 315334
rect 62422 315098 98186 315334
rect 98422 315098 134186 315334
rect 134422 315098 170186 315334
rect 170422 315098 206186 315334
rect 206422 315098 242186 315334
rect 242422 315098 278186 315334
rect 278422 315098 314186 315334
rect 314422 315098 350186 315334
rect 350422 315098 386186 315334
rect 386422 315098 422186 315334
rect 422422 315098 458186 315334
rect 458422 315098 494186 315334
rect 494422 315098 530186 315334
rect 530422 315098 566186 315334
rect 566422 315098 590202 315334
rect 590438 315098 590620 315334
rect -6696 315076 590620 315098
rect -6696 315074 -6096 315076
rect 26004 315074 26604 315076
rect 62004 315074 62604 315076
rect 98004 315074 98604 315076
rect 134004 315074 134604 315076
rect 170004 315074 170604 315076
rect 206004 315074 206604 315076
rect 242004 315074 242604 315076
rect 278004 315074 278604 315076
rect 314004 315074 314604 315076
rect 350004 315074 350604 315076
rect 386004 315074 386604 315076
rect 422004 315074 422604 315076
rect 458004 315074 458604 315076
rect 494004 315074 494604 315076
rect 530004 315074 530604 315076
rect 566004 315074 566604 315076
rect 590020 315074 590620 315076
rect -4816 312076 -4216 312078
rect 22404 312076 23004 312078
rect 58404 312076 59004 312078
rect 94404 312076 95004 312078
rect 130404 312076 131004 312078
rect 166404 312076 167004 312078
rect 202404 312076 203004 312078
rect 238404 312076 239004 312078
rect 274404 312076 275004 312078
rect 310404 312076 311004 312078
rect 346404 312076 347004 312078
rect 382404 312076 383004 312078
rect 418404 312076 419004 312078
rect 454404 312076 455004 312078
rect 490404 312076 491004 312078
rect 526404 312076 527004 312078
rect 562404 312076 563004 312078
rect 588140 312076 588740 312078
rect -4816 312054 588740 312076
rect -4816 311818 -4634 312054
rect -4398 311818 22586 312054
rect 22822 311818 58586 312054
rect 58822 311818 94586 312054
rect 94822 311818 130586 312054
rect 130822 311818 166586 312054
rect 166822 311818 202586 312054
rect 202822 311818 238586 312054
rect 238822 311818 274586 312054
rect 274822 311818 310586 312054
rect 310822 311818 346586 312054
rect 346822 311818 382586 312054
rect 382822 311818 418586 312054
rect 418822 311818 454586 312054
rect 454822 311818 490586 312054
rect 490822 311818 526586 312054
rect 526822 311818 562586 312054
rect 562822 311818 588322 312054
rect 588558 311818 588740 312054
rect -4816 311734 588740 311818
rect -4816 311498 -4634 311734
rect -4398 311498 22586 311734
rect 22822 311498 58586 311734
rect 58822 311498 94586 311734
rect 94822 311498 130586 311734
rect 130822 311498 166586 311734
rect 166822 311498 202586 311734
rect 202822 311498 238586 311734
rect 238822 311498 274586 311734
rect 274822 311498 310586 311734
rect 310822 311498 346586 311734
rect 346822 311498 382586 311734
rect 382822 311498 418586 311734
rect 418822 311498 454586 311734
rect 454822 311498 490586 311734
rect 490822 311498 526586 311734
rect 526822 311498 562586 311734
rect 562822 311498 588322 311734
rect 588558 311498 588740 311734
rect -4816 311476 588740 311498
rect -4816 311474 -4216 311476
rect 22404 311474 23004 311476
rect 58404 311474 59004 311476
rect 94404 311474 95004 311476
rect 130404 311474 131004 311476
rect 166404 311474 167004 311476
rect 202404 311474 203004 311476
rect 238404 311474 239004 311476
rect 274404 311474 275004 311476
rect 310404 311474 311004 311476
rect 346404 311474 347004 311476
rect 382404 311474 383004 311476
rect 418404 311474 419004 311476
rect 454404 311474 455004 311476
rect 490404 311474 491004 311476
rect 526404 311474 527004 311476
rect 562404 311474 563004 311476
rect 588140 311474 588740 311476
rect -2936 308476 -2336 308478
rect 18804 308476 19404 308478
rect 54804 308476 55404 308478
rect 90804 308476 91404 308478
rect 126804 308476 127404 308478
rect 162804 308476 163404 308478
rect 198804 308476 199404 308478
rect 234804 308476 235404 308478
rect 270804 308476 271404 308478
rect 306804 308476 307404 308478
rect 342804 308476 343404 308478
rect 378804 308476 379404 308478
rect 414804 308476 415404 308478
rect 450804 308476 451404 308478
rect 486804 308476 487404 308478
rect 522804 308476 523404 308478
rect 558804 308476 559404 308478
rect 586260 308476 586860 308478
rect -2936 308454 586860 308476
rect -2936 308218 -2754 308454
rect -2518 308218 18986 308454
rect 19222 308218 54986 308454
rect 55222 308218 90986 308454
rect 91222 308218 126986 308454
rect 127222 308218 162986 308454
rect 163222 308218 198986 308454
rect 199222 308218 234986 308454
rect 235222 308218 270986 308454
rect 271222 308218 306986 308454
rect 307222 308218 342986 308454
rect 343222 308218 378986 308454
rect 379222 308218 414986 308454
rect 415222 308218 450986 308454
rect 451222 308218 486986 308454
rect 487222 308218 522986 308454
rect 523222 308218 558986 308454
rect 559222 308218 586442 308454
rect 586678 308218 586860 308454
rect -2936 308134 586860 308218
rect -2936 307898 -2754 308134
rect -2518 307898 18986 308134
rect 19222 307898 54986 308134
rect 55222 307898 90986 308134
rect 91222 307898 126986 308134
rect 127222 307898 162986 308134
rect 163222 307898 198986 308134
rect 199222 307898 234986 308134
rect 235222 307898 270986 308134
rect 271222 307898 306986 308134
rect 307222 307898 342986 308134
rect 343222 307898 378986 308134
rect 379222 307898 414986 308134
rect 415222 307898 450986 308134
rect 451222 307898 486986 308134
rect 487222 307898 522986 308134
rect 523222 307898 558986 308134
rect 559222 307898 586442 308134
rect 586678 307898 586860 308134
rect -2936 307876 586860 307898
rect -2936 307874 -2336 307876
rect 18804 307874 19404 307876
rect 54804 307874 55404 307876
rect 90804 307874 91404 307876
rect 126804 307874 127404 307876
rect 162804 307874 163404 307876
rect 198804 307874 199404 307876
rect 234804 307874 235404 307876
rect 270804 307874 271404 307876
rect 306804 307874 307404 307876
rect 342804 307874 343404 307876
rect 378804 307874 379404 307876
rect 414804 307874 415404 307876
rect 450804 307874 451404 307876
rect 486804 307874 487404 307876
rect 522804 307874 523404 307876
rect 558804 307874 559404 307876
rect 586260 307874 586860 307876
rect -7636 301276 -7036 301278
rect 11604 301276 12204 301278
rect 47604 301276 48204 301278
rect 83604 301276 84204 301278
rect 119604 301276 120204 301278
rect 155604 301276 156204 301278
rect 191604 301276 192204 301278
rect 227604 301276 228204 301278
rect 263604 301276 264204 301278
rect 299604 301276 300204 301278
rect 551604 301276 552204 301278
rect 590960 301276 591560 301278
rect -8576 301254 592500 301276
rect -8576 301018 -7454 301254
rect -7218 301018 11786 301254
rect 12022 301018 47786 301254
rect 48022 301018 83786 301254
rect 84022 301018 119786 301254
rect 120022 301018 155786 301254
rect 156022 301018 191786 301254
rect 192022 301018 227786 301254
rect 228022 301018 263786 301254
rect 264022 301018 299786 301254
rect 300022 301018 551786 301254
rect 552022 301018 591142 301254
rect 591378 301018 592500 301254
rect -8576 300934 592500 301018
rect -8576 300698 -7454 300934
rect -7218 300698 11786 300934
rect 12022 300698 47786 300934
rect 48022 300698 83786 300934
rect 84022 300698 119786 300934
rect 120022 300698 155786 300934
rect 156022 300698 191786 300934
rect 192022 300698 227786 300934
rect 228022 300698 263786 300934
rect 264022 300698 299786 300934
rect 300022 300698 551786 300934
rect 552022 300698 591142 300934
rect 591378 300698 592500 300934
rect -8576 300676 592500 300698
rect -7636 300674 -7036 300676
rect 11604 300674 12204 300676
rect 47604 300674 48204 300676
rect 83604 300674 84204 300676
rect 119604 300674 120204 300676
rect 155604 300674 156204 300676
rect 191604 300674 192204 300676
rect 227604 300674 228204 300676
rect 263604 300674 264204 300676
rect 299604 300674 300204 300676
rect 551604 300674 552204 300676
rect 590960 300674 591560 300676
rect -5756 297676 -5156 297678
rect 8004 297676 8604 297678
rect 44004 297676 44604 297678
rect 80004 297676 80604 297678
rect 116004 297676 116604 297678
rect 152004 297676 152604 297678
rect 188004 297676 188604 297678
rect 224004 297676 224604 297678
rect 260004 297676 260604 297678
rect 296004 297676 296604 297678
rect 548004 297676 548604 297678
rect 589080 297676 589680 297678
rect -6696 297654 590620 297676
rect -6696 297418 -5574 297654
rect -5338 297418 8186 297654
rect 8422 297418 44186 297654
rect 44422 297418 80186 297654
rect 80422 297418 116186 297654
rect 116422 297418 152186 297654
rect 152422 297418 188186 297654
rect 188422 297418 224186 297654
rect 224422 297418 260186 297654
rect 260422 297418 296186 297654
rect 296422 297418 548186 297654
rect 548422 297418 589262 297654
rect 589498 297418 590620 297654
rect -6696 297334 590620 297418
rect -6696 297098 -5574 297334
rect -5338 297098 8186 297334
rect 8422 297098 44186 297334
rect 44422 297098 80186 297334
rect 80422 297098 116186 297334
rect 116422 297098 152186 297334
rect 152422 297098 188186 297334
rect 188422 297098 224186 297334
rect 224422 297098 260186 297334
rect 260422 297098 296186 297334
rect 296422 297098 548186 297334
rect 548422 297098 589262 297334
rect 589498 297098 590620 297334
rect -6696 297076 590620 297098
rect -5756 297074 -5156 297076
rect 8004 297074 8604 297076
rect 44004 297074 44604 297076
rect 80004 297074 80604 297076
rect 116004 297074 116604 297076
rect 152004 297074 152604 297076
rect 188004 297074 188604 297076
rect 224004 297074 224604 297076
rect 260004 297074 260604 297076
rect 296004 297074 296604 297076
rect 548004 297074 548604 297076
rect 589080 297074 589680 297076
rect -3876 294076 -3276 294078
rect 4404 294076 5004 294078
rect 40404 294076 41004 294078
rect 76404 294076 77004 294078
rect 112404 294076 113004 294078
rect 148404 294076 149004 294078
rect 184404 294076 185004 294078
rect 220404 294076 221004 294078
rect 256404 294076 257004 294078
rect 292404 294076 293004 294078
rect 314208 294076 314528 294078
rect 544404 294076 545004 294078
rect 580404 294076 581004 294078
rect 587200 294076 587800 294078
rect -4816 294054 588740 294076
rect -4816 293818 -3694 294054
rect -3458 293818 4586 294054
rect 4822 293818 40586 294054
rect 40822 293818 76586 294054
rect 76822 293818 112586 294054
rect 112822 293818 148586 294054
rect 148822 293818 184586 294054
rect 184822 293818 220586 294054
rect 220822 293818 256586 294054
rect 256822 293818 292586 294054
rect 292822 293818 314250 294054
rect 314486 293818 544586 294054
rect 544822 293818 580586 294054
rect 580822 293818 587382 294054
rect 587618 293818 588740 294054
rect -4816 293734 588740 293818
rect -4816 293498 -3694 293734
rect -3458 293498 4586 293734
rect 4822 293498 40586 293734
rect 40822 293498 76586 293734
rect 76822 293498 112586 293734
rect 112822 293498 148586 293734
rect 148822 293498 184586 293734
rect 184822 293498 220586 293734
rect 220822 293498 256586 293734
rect 256822 293498 292586 293734
rect 292822 293498 314250 293734
rect 314486 293498 544586 293734
rect 544822 293498 580586 293734
rect 580822 293498 587382 293734
rect 587618 293498 588740 293734
rect -4816 293476 588740 293498
rect -3876 293474 -3276 293476
rect 4404 293474 5004 293476
rect 40404 293474 41004 293476
rect 76404 293474 77004 293476
rect 112404 293474 113004 293476
rect 148404 293474 149004 293476
rect 184404 293474 185004 293476
rect 220404 293474 221004 293476
rect 256404 293474 257004 293476
rect 292404 293474 293004 293476
rect 314208 293474 314528 293476
rect 544404 293474 545004 293476
rect 580404 293474 581004 293476
rect 587200 293474 587800 293476
rect -1996 290476 -1396 290478
rect 804 290476 1404 290478
rect 36804 290476 37404 290478
rect 72804 290476 73404 290478
rect 108804 290476 109404 290478
rect 144804 290476 145404 290478
rect 180804 290476 181404 290478
rect 216804 290476 217404 290478
rect 252804 290476 253404 290478
rect 288804 290476 289404 290478
rect 314208 290476 314528 290478
rect 540804 290476 541404 290478
rect 576804 290476 577404 290478
rect 585320 290476 585920 290478
rect -2936 290454 586860 290476
rect -2936 290218 -1814 290454
rect -1578 290218 986 290454
rect 1222 290218 36986 290454
rect 37222 290218 72986 290454
rect 73222 290218 108986 290454
rect 109222 290218 144986 290454
rect 145222 290218 180986 290454
rect 181222 290218 216986 290454
rect 217222 290218 252986 290454
rect 253222 290218 288986 290454
rect 289222 290218 314250 290454
rect 314486 290218 540986 290454
rect 541222 290218 576986 290454
rect 577222 290218 585502 290454
rect 585738 290218 586860 290454
rect -2936 290134 586860 290218
rect -2936 289898 -1814 290134
rect -1578 289898 986 290134
rect 1222 289898 36986 290134
rect 37222 289898 72986 290134
rect 73222 289898 108986 290134
rect 109222 289898 144986 290134
rect 145222 289898 180986 290134
rect 181222 289898 216986 290134
rect 217222 289898 252986 290134
rect 253222 289898 288986 290134
rect 289222 289898 314250 290134
rect 314486 289898 540986 290134
rect 541222 289898 576986 290134
rect 577222 289898 585502 290134
rect 585738 289898 586860 290134
rect -2936 289876 586860 289898
rect -1996 289874 -1396 289876
rect 804 289874 1404 289876
rect 36804 289874 37404 289876
rect 72804 289874 73404 289876
rect 108804 289874 109404 289876
rect 144804 289874 145404 289876
rect 180804 289874 181404 289876
rect 216804 289874 217404 289876
rect 252804 289874 253404 289876
rect 288804 289874 289404 289876
rect 314208 289874 314528 289876
rect 540804 289874 541404 289876
rect 576804 289874 577404 289876
rect 585320 289874 585920 289876
rect -8576 283276 -7976 283278
rect 29604 283276 30204 283278
rect 65604 283276 66204 283278
rect 101604 283276 102204 283278
rect 137604 283276 138204 283278
rect 173604 283276 174204 283278
rect 209604 283276 210204 283278
rect 245604 283276 246204 283278
rect 281604 283276 282204 283278
rect 329568 283276 329888 283278
rect 533604 283276 534204 283278
rect 569604 283276 570204 283278
rect 591900 283276 592500 283278
rect -8576 283254 592500 283276
rect -8576 283018 -8394 283254
rect -8158 283018 29786 283254
rect 30022 283018 65786 283254
rect 66022 283018 101786 283254
rect 102022 283018 137786 283254
rect 138022 283018 173786 283254
rect 174022 283018 209786 283254
rect 210022 283018 245786 283254
rect 246022 283018 281786 283254
rect 282022 283018 329610 283254
rect 329846 283018 533786 283254
rect 534022 283018 569786 283254
rect 570022 283018 592082 283254
rect 592318 283018 592500 283254
rect -8576 282934 592500 283018
rect -8576 282698 -8394 282934
rect -8158 282698 29786 282934
rect 30022 282698 65786 282934
rect 66022 282698 101786 282934
rect 102022 282698 137786 282934
rect 138022 282698 173786 282934
rect 174022 282698 209786 282934
rect 210022 282698 245786 282934
rect 246022 282698 281786 282934
rect 282022 282698 329610 282934
rect 329846 282698 533786 282934
rect 534022 282698 569786 282934
rect 570022 282698 592082 282934
rect 592318 282698 592500 282934
rect -8576 282676 592500 282698
rect -8576 282674 -7976 282676
rect 29604 282674 30204 282676
rect 65604 282674 66204 282676
rect 101604 282674 102204 282676
rect 137604 282674 138204 282676
rect 173604 282674 174204 282676
rect 209604 282674 210204 282676
rect 245604 282674 246204 282676
rect 281604 282674 282204 282676
rect 329568 282674 329888 282676
rect 533604 282674 534204 282676
rect 569604 282674 570204 282676
rect 591900 282674 592500 282676
rect -6696 279676 -6096 279678
rect 26004 279676 26604 279678
rect 62004 279676 62604 279678
rect 98004 279676 98604 279678
rect 134004 279676 134604 279678
rect 170004 279676 170604 279678
rect 206004 279676 206604 279678
rect 242004 279676 242604 279678
rect 278004 279676 278604 279678
rect 329568 279676 329888 279678
rect 566004 279676 566604 279678
rect 590020 279676 590620 279678
rect -6696 279654 590620 279676
rect -6696 279418 -6514 279654
rect -6278 279418 26186 279654
rect 26422 279418 62186 279654
rect 62422 279418 98186 279654
rect 98422 279418 134186 279654
rect 134422 279418 170186 279654
rect 170422 279418 206186 279654
rect 206422 279418 242186 279654
rect 242422 279418 278186 279654
rect 278422 279418 329610 279654
rect 329846 279418 566186 279654
rect 566422 279418 590202 279654
rect 590438 279418 590620 279654
rect -6696 279334 590620 279418
rect -6696 279098 -6514 279334
rect -6278 279098 26186 279334
rect 26422 279098 62186 279334
rect 62422 279098 98186 279334
rect 98422 279098 134186 279334
rect 134422 279098 170186 279334
rect 170422 279098 206186 279334
rect 206422 279098 242186 279334
rect 242422 279098 278186 279334
rect 278422 279098 329610 279334
rect 329846 279098 566186 279334
rect 566422 279098 590202 279334
rect 590438 279098 590620 279334
rect -6696 279076 590620 279098
rect -6696 279074 -6096 279076
rect 26004 279074 26604 279076
rect 62004 279074 62604 279076
rect 98004 279074 98604 279076
rect 134004 279074 134604 279076
rect 170004 279074 170604 279076
rect 206004 279074 206604 279076
rect 242004 279074 242604 279076
rect 278004 279074 278604 279076
rect 329568 279074 329888 279076
rect 566004 279074 566604 279076
rect 590020 279074 590620 279076
rect -4816 276076 -4216 276078
rect 22404 276076 23004 276078
rect 58404 276076 59004 276078
rect 94404 276076 95004 276078
rect 130404 276076 131004 276078
rect 166404 276076 167004 276078
rect 202404 276076 203004 276078
rect 238404 276076 239004 276078
rect 274404 276076 275004 276078
rect 329568 276076 329888 276078
rect 562404 276076 563004 276078
rect 588140 276076 588740 276078
rect -4816 276054 588740 276076
rect -4816 275818 -4634 276054
rect -4398 275818 22586 276054
rect 22822 275818 58586 276054
rect 58822 275818 94586 276054
rect 94822 275818 130586 276054
rect 130822 275818 166586 276054
rect 166822 275818 202586 276054
rect 202822 275818 238586 276054
rect 238822 275818 274586 276054
rect 274822 275818 329610 276054
rect 329846 275818 562586 276054
rect 562822 275818 588322 276054
rect 588558 275818 588740 276054
rect -4816 275734 588740 275818
rect -4816 275498 -4634 275734
rect -4398 275498 22586 275734
rect 22822 275498 58586 275734
rect 58822 275498 94586 275734
rect 94822 275498 130586 275734
rect 130822 275498 166586 275734
rect 166822 275498 202586 275734
rect 202822 275498 238586 275734
rect 238822 275498 274586 275734
rect 274822 275498 329610 275734
rect 329846 275498 562586 275734
rect 562822 275498 588322 275734
rect 588558 275498 588740 275734
rect -4816 275476 588740 275498
rect -4816 275474 -4216 275476
rect 22404 275474 23004 275476
rect 58404 275474 59004 275476
rect 94404 275474 95004 275476
rect 130404 275474 131004 275476
rect 166404 275474 167004 275476
rect 202404 275474 203004 275476
rect 238404 275474 239004 275476
rect 274404 275474 275004 275476
rect 329568 275474 329888 275476
rect 562404 275474 563004 275476
rect 588140 275474 588740 275476
rect -2936 272476 -2336 272478
rect 18804 272476 19404 272478
rect 54804 272476 55404 272478
rect 90804 272476 91404 272478
rect 126804 272476 127404 272478
rect 162804 272476 163404 272478
rect 198804 272476 199404 272478
rect 234804 272476 235404 272478
rect 270804 272476 271404 272478
rect 329568 272476 329888 272478
rect 558804 272476 559404 272478
rect 586260 272476 586860 272478
rect -2936 272454 586860 272476
rect -2936 272218 -2754 272454
rect -2518 272218 18986 272454
rect 19222 272218 54986 272454
rect 55222 272218 90986 272454
rect 91222 272218 126986 272454
rect 127222 272218 162986 272454
rect 163222 272218 198986 272454
rect 199222 272218 234986 272454
rect 235222 272218 270986 272454
rect 271222 272218 329610 272454
rect 329846 272218 558986 272454
rect 559222 272218 586442 272454
rect 586678 272218 586860 272454
rect -2936 272134 586860 272218
rect -2936 271898 -2754 272134
rect -2518 271898 18986 272134
rect 19222 271898 54986 272134
rect 55222 271898 90986 272134
rect 91222 271898 126986 272134
rect 127222 271898 162986 272134
rect 163222 271898 198986 272134
rect 199222 271898 234986 272134
rect 235222 271898 270986 272134
rect 271222 271898 329610 272134
rect 329846 271898 558986 272134
rect 559222 271898 586442 272134
rect 586678 271898 586860 272134
rect -2936 271876 586860 271898
rect -2936 271874 -2336 271876
rect 18804 271874 19404 271876
rect 54804 271874 55404 271876
rect 90804 271874 91404 271876
rect 126804 271874 127404 271876
rect 162804 271874 163404 271876
rect 198804 271874 199404 271876
rect 234804 271874 235404 271876
rect 270804 271874 271404 271876
rect 329568 271874 329888 271876
rect 558804 271874 559404 271876
rect 586260 271874 586860 271876
rect -7636 265276 -7036 265278
rect 11604 265276 12204 265278
rect 47604 265276 48204 265278
rect 83604 265276 84204 265278
rect 119604 265276 120204 265278
rect 155604 265276 156204 265278
rect 191604 265276 192204 265278
rect 227604 265276 228204 265278
rect 263604 265276 264204 265278
rect 299604 265276 300204 265278
rect 314208 265276 314528 265278
rect 551604 265276 552204 265278
rect 590960 265276 591560 265278
rect -8576 265254 592500 265276
rect -8576 265018 -7454 265254
rect -7218 265018 11786 265254
rect 12022 265018 47786 265254
rect 48022 265018 83786 265254
rect 84022 265018 119786 265254
rect 120022 265018 155786 265254
rect 156022 265018 191786 265254
rect 192022 265018 227786 265254
rect 228022 265018 263786 265254
rect 264022 265018 299786 265254
rect 300022 265018 314250 265254
rect 314486 265018 551786 265254
rect 552022 265018 591142 265254
rect 591378 265018 592500 265254
rect -8576 264934 592500 265018
rect -8576 264698 -7454 264934
rect -7218 264698 11786 264934
rect 12022 264698 47786 264934
rect 48022 264698 83786 264934
rect 84022 264698 119786 264934
rect 120022 264698 155786 264934
rect 156022 264698 191786 264934
rect 192022 264698 227786 264934
rect 228022 264698 263786 264934
rect 264022 264698 299786 264934
rect 300022 264698 314250 264934
rect 314486 264698 551786 264934
rect 552022 264698 591142 264934
rect 591378 264698 592500 264934
rect -8576 264676 592500 264698
rect -7636 264674 -7036 264676
rect 11604 264674 12204 264676
rect 47604 264674 48204 264676
rect 83604 264674 84204 264676
rect 119604 264674 120204 264676
rect 155604 264674 156204 264676
rect 191604 264674 192204 264676
rect 227604 264674 228204 264676
rect 263604 264674 264204 264676
rect 299604 264674 300204 264676
rect 314208 264674 314528 264676
rect 551604 264674 552204 264676
rect 590960 264674 591560 264676
rect -5756 261676 -5156 261678
rect 8004 261676 8604 261678
rect 44004 261676 44604 261678
rect 80004 261676 80604 261678
rect 116004 261676 116604 261678
rect 152004 261676 152604 261678
rect 188004 261676 188604 261678
rect 224004 261676 224604 261678
rect 260004 261676 260604 261678
rect 296004 261676 296604 261678
rect 314208 261676 314528 261678
rect 548004 261676 548604 261678
rect 589080 261676 589680 261678
rect -6696 261654 590620 261676
rect -6696 261418 -5574 261654
rect -5338 261418 8186 261654
rect 8422 261418 44186 261654
rect 44422 261418 80186 261654
rect 80422 261418 116186 261654
rect 116422 261418 152186 261654
rect 152422 261418 188186 261654
rect 188422 261418 224186 261654
rect 224422 261418 260186 261654
rect 260422 261418 296186 261654
rect 296422 261418 314250 261654
rect 314486 261418 548186 261654
rect 548422 261418 589262 261654
rect 589498 261418 590620 261654
rect -6696 261334 590620 261418
rect -6696 261098 -5574 261334
rect -5338 261098 8186 261334
rect 8422 261098 44186 261334
rect 44422 261098 80186 261334
rect 80422 261098 116186 261334
rect 116422 261098 152186 261334
rect 152422 261098 188186 261334
rect 188422 261098 224186 261334
rect 224422 261098 260186 261334
rect 260422 261098 296186 261334
rect 296422 261098 314250 261334
rect 314486 261098 548186 261334
rect 548422 261098 589262 261334
rect 589498 261098 590620 261334
rect -6696 261076 590620 261098
rect -5756 261074 -5156 261076
rect 8004 261074 8604 261076
rect 44004 261074 44604 261076
rect 80004 261074 80604 261076
rect 116004 261074 116604 261076
rect 152004 261074 152604 261076
rect 188004 261074 188604 261076
rect 224004 261074 224604 261076
rect 260004 261074 260604 261076
rect 296004 261074 296604 261076
rect 314208 261074 314528 261076
rect 548004 261074 548604 261076
rect 589080 261074 589680 261076
rect -3876 258076 -3276 258078
rect 4404 258076 5004 258078
rect 40404 258076 41004 258078
rect 76404 258076 77004 258078
rect 112404 258076 113004 258078
rect 148404 258076 149004 258078
rect 184404 258076 185004 258078
rect 220404 258076 221004 258078
rect 256404 258076 257004 258078
rect 292404 258076 293004 258078
rect 314208 258076 314528 258078
rect 544404 258076 545004 258078
rect 580404 258076 581004 258078
rect 587200 258076 587800 258078
rect -4816 258054 588740 258076
rect -4816 257818 -3694 258054
rect -3458 257818 4586 258054
rect 4822 257818 40586 258054
rect 40822 257818 76586 258054
rect 76822 257818 112586 258054
rect 112822 257818 148586 258054
rect 148822 257818 184586 258054
rect 184822 257818 220586 258054
rect 220822 257818 256586 258054
rect 256822 257818 292586 258054
rect 292822 257818 314250 258054
rect 314486 257818 544586 258054
rect 544822 257818 580586 258054
rect 580822 257818 587382 258054
rect 587618 257818 588740 258054
rect -4816 257734 588740 257818
rect -4816 257498 -3694 257734
rect -3458 257498 4586 257734
rect 4822 257498 40586 257734
rect 40822 257498 76586 257734
rect 76822 257498 112586 257734
rect 112822 257498 148586 257734
rect 148822 257498 184586 257734
rect 184822 257498 220586 257734
rect 220822 257498 256586 257734
rect 256822 257498 292586 257734
rect 292822 257498 314250 257734
rect 314486 257498 544586 257734
rect 544822 257498 580586 257734
rect 580822 257498 587382 257734
rect 587618 257498 588740 257734
rect -4816 257476 588740 257498
rect -3876 257474 -3276 257476
rect 4404 257474 5004 257476
rect 40404 257474 41004 257476
rect 76404 257474 77004 257476
rect 112404 257474 113004 257476
rect 148404 257474 149004 257476
rect 184404 257474 185004 257476
rect 220404 257474 221004 257476
rect 256404 257474 257004 257476
rect 292404 257474 293004 257476
rect 314208 257474 314528 257476
rect 544404 257474 545004 257476
rect 580404 257474 581004 257476
rect 587200 257474 587800 257476
rect -1996 254476 -1396 254478
rect 804 254476 1404 254478
rect 36804 254476 37404 254478
rect 72804 254476 73404 254478
rect 108804 254476 109404 254478
rect 144804 254476 145404 254478
rect 180804 254476 181404 254478
rect 216804 254476 217404 254478
rect 252804 254476 253404 254478
rect 288804 254476 289404 254478
rect 314208 254476 314528 254478
rect 540804 254476 541404 254478
rect 576804 254476 577404 254478
rect 585320 254476 585920 254478
rect -2936 254454 586860 254476
rect -2936 254218 -1814 254454
rect -1578 254218 986 254454
rect 1222 254218 36986 254454
rect 37222 254218 72986 254454
rect 73222 254218 108986 254454
rect 109222 254218 144986 254454
rect 145222 254218 180986 254454
rect 181222 254218 216986 254454
rect 217222 254218 252986 254454
rect 253222 254218 288986 254454
rect 289222 254218 314250 254454
rect 314486 254218 540986 254454
rect 541222 254218 576986 254454
rect 577222 254218 585502 254454
rect 585738 254218 586860 254454
rect -2936 254134 586860 254218
rect -2936 253898 -1814 254134
rect -1578 253898 986 254134
rect 1222 253898 36986 254134
rect 37222 253898 72986 254134
rect 73222 253898 108986 254134
rect 109222 253898 144986 254134
rect 145222 253898 180986 254134
rect 181222 253898 216986 254134
rect 217222 253898 252986 254134
rect 253222 253898 288986 254134
rect 289222 253898 314250 254134
rect 314486 253898 540986 254134
rect 541222 253898 576986 254134
rect 577222 253898 585502 254134
rect 585738 253898 586860 254134
rect -2936 253876 586860 253898
rect -1996 253874 -1396 253876
rect 804 253874 1404 253876
rect 36804 253874 37404 253876
rect 72804 253874 73404 253876
rect 108804 253874 109404 253876
rect 144804 253874 145404 253876
rect 180804 253874 181404 253876
rect 216804 253874 217404 253876
rect 252804 253874 253404 253876
rect 288804 253874 289404 253876
rect 314208 253874 314528 253876
rect 540804 253874 541404 253876
rect 576804 253874 577404 253876
rect 585320 253874 585920 253876
rect -8576 247276 -7976 247278
rect 29604 247276 30204 247278
rect 65604 247276 66204 247278
rect 101604 247276 102204 247278
rect 137604 247276 138204 247278
rect 173604 247276 174204 247278
rect 209604 247276 210204 247278
rect 245604 247276 246204 247278
rect 281604 247276 282204 247278
rect 329568 247276 329888 247278
rect 533604 247276 534204 247278
rect 569604 247276 570204 247278
rect 591900 247276 592500 247278
rect -8576 247254 592500 247276
rect -8576 247018 -8394 247254
rect -8158 247018 29786 247254
rect 30022 247018 65786 247254
rect 66022 247018 101786 247254
rect 102022 247018 137786 247254
rect 138022 247018 173786 247254
rect 174022 247018 209786 247254
rect 210022 247018 245786 247254
rect 246022 247018 281786 247254
rect 282022 247018 329610 247254
rect 329846 247018 533786 247254
rect 534022 247018 569786 247254
rect 570022 247018 592082 247254
rect 592318 247018 592500 247254
rect -8576 246934 592500 247018
rect -8576 246698 -8394 246934
rect -8158 246698 29786 246934
rect 30022 246698 65786 246934
rect 66022 246698 101786 246934
rect 102022 246698 137786 246934
rect 138022 246698 173786 246934
rect 174022 246698 209786 246934
rect 210022 246698 245786 246934
rect 246022 246698 281786 246934
rect 282022 246698 329610 246934
rect 329846 246698 533786 246934
rect 534022 246698 569786 246934
rect 570022 246698 592082 246934
rect 592318 246698 592500 246934
rect -8576 246676 592500 246698
rect -8576 246674 -7976 246676
rect 29604 246674 30204 246676
rect 65604 246674 66204 246676
rect 101604 246674 102204 246676
rect 137604 246674 138204 246676
rect 173604 246674 174204 246676
rect 209604 246674 210204 246676
rect 245604 246674 246204 246676
rect 281604 246674 282204 246676
rect 329568 246674 329888 246676
rect 533604 246674 534204 246676
rect 569604 246674 570204 246676
rect 591900 246674 592500 246676
rect -6696 243676 -6096 243678
rect 26004 243676 26604 243678
rect 62004 243676 62604 243678
rect 98004 243676 98604 243678
rect 134004 243676 134604 243678
rect 170004 243676 170604 243678
rect 206004 243676 206604 243678
rect 242004 243676 242604 243678
rect 278004 243676 278604 243678
rect 329568 243676 329888 243678
rect 566004 243676 566604 243678
rect 590020 243676 590620 243678
rect -6696 243654 590620 243676
rect -6696 243418 -6514 243654
rect -6278 243418 26186 243654
rect 26422 243418 62186 243654
rect 62422 243418 98186 243654
rect 98422 243418 134186 243654
rect 134422 243418 170186 243654
rect 170422 243418 206186 243654
rect 206422 243418 242186 243654
rect 242422 243418 278186 243654
rect 278422 243418 329610 243654
rect 329846 243418 566186 243654
rect 566422 243418 590202 243654
rect 590438 243418 590620 243654
rect -6696 243334 590620 243418
rect -6696 243098 -6514 243334
rect -6278 243098 26186 243334
rect 26422 243098 62186 243334
rect 62422 243098 98186 243334
rect 98422 243098 134186 243334
rect 134422 243098 170186 243334
rect 170422 243098 206186 243334
rect 206422 243098 242186 243334
rect 242422 243098 278186 243334
rect 278422 243098 329610 243334
rect 329846 243098 566186 243334
rect 566422 243098 590202 243334
rect 590438 243098 590620 243334
rect -6696 243076 590620 243098
rect -6696 243074 -6096 243076
rect 26004 243074 26604 243076
rect 62004 243074 62604 243076
rect 98004 243074 98604 243076
rect 134004 243074 134604 243076
rect 170004 243074 170604 243076
rect 206004 243074 206604 243076
rect 242004 243074 242604 243076
rect 278004 243074 278604 243076
rect 329568 243074 329888 243076
rect 566004 243074 566604 243076
rect 590020 243074 590620 243076
rect -4816 240076 -4216 240078
rect 22404 240076 23004 240078
rect 58404 240076 59004 240078
rect 94404 240076 95004 240078
rect 130404 240076 131004 240078
rect 166404 240076 167004 240078
rect 202404 240076 203004 240078
rect 238404 240076 239004 240078
rect 274404 240076 275004 240078
rect 329568 240076 329888 240078
rect 562404 240076 563004 240078
rect 588140 240076 588740 240078
rect -4816 240054 588740 240076
rect -4816 239818 -4634 240054
rect -4398 239818 22586 240054
rect 22822 239818 58586 240054
rect 58822 239818 94586 240054
rect 94822 239818 130586 240054
rect 130822 239818 166586 240054
rect 166822 239818 202586 240054
rect 202822 239818 238586 240054
rect 238822 239818 274586 240054
rect 274822 239818 329610 240054
rect 329846 239818 562586 240054
rect 562822 239818 588322 240054
rect 588558 239818 588740 240054
rect -4816 239734 588740 239818
rect -4816 239498 -4634 239734
rect -4398 239498 22586 239734
rect 22822 239498 58586 239734
rect 58822 239498 94586 239734
rect 94822 239498 130586 239734
rect 130822 239498 166586 239734
rect 166822 239498 202586 239734
rect 202822 239498 238586 239734
rect 238822 239498 274586 239734
rect 274822 239498 329610 239734
rect 329846 239498 562586 239734
rect 562822 239498 588322 239734
rect 588558 239498 588740 239734
rect -4816 239476 588740 239498
rect -4816 239474 -4216 239476
rect 22404 239474 23004 239476
rect 58404 239474 59004 239476
rect 94404 239474 95004 239476
rect 130404 239474 131004 239476
rect 166404 239474 167004 239476
rect 202404 239474 203004 239476
rect 238404 239474 239004 239476
rect 274404 239474 275004 239476
rect 329568 239474 329888 239476
rect 562404 239474 563004 239476
rect 588140 239474 588740 239476
rect -2936 236476 -2336 236478
rect 18804 236476 19404 236478
rect 54804 236476 55404 236478
rect 90804 236476 91404 236478
rect 126804 236476 127404 236478
rect 162804 236476 163404 236478
rect 198804 236476 199404 236478
rect 234804 236476 235404 236478
rect 270804 236476 271404 236478
rect 329568 236476 329888 236478
rect 558804 236476 559404 236478
rect 586260 236476 586860 236478
rect -2936 236454 586860 236476
rect -2936 236218 -2754 236454
rect -2518 236218 18986 236454
rect 19222 236218 54986 236454
rect 55222 236218 90986 236454
rect 91222 236218 126986 236454
rect 127222 236218 162986 236454
rect 163222 236218 198986 236454
rect 199222 236218 234986 236454
rect 235222 236218 270986 236454
rect 271222 236218 329610 236454
rect 329846 236218 558986 236454
rect 559222 236218 586442 236454
rect 586678 236218 586860 236454
rect -2936 236134 586860 236218
rect -2936 235898 -2754 236134
rect -2518 235898 18986 236134
rect 19222 235898 54986 236134
rect 55222 235898 90986 236134
rect 91222 235898 126986 236134
rect 127222 235898 162986 236134
rect 163222 235898 198986 236134
rect 199222 235898 234986 236134
rect 235222 235898 270986 236134
rect 271222 235898 329610 236134
rect 329846 235898 558986 236134
rect 559222 235898 586442 236134
rect 586678 235898 586860 236134
rect -2936 235876 586860 235898
rect -2936 235874 -2336 235876
rect 18804 235874 19404 235876
rect 54804 235874 55404 235876
rect 90804 235874 91404 235876
rect 126804 235874 127404 235876
rect 162804 235874 163404 235876
rect 198804 235874 199404 235876
rect 234804 235874 235404 235876
rect 270804 235874 271404 235876
rect 329568 235874 329888 235876
rect 558804 235874 559404 235876
rect 586260 235874 586860 235876
rect -7636 229276 -7036 229278
rect 11604 229276 12204 229278
rect 47604 229276 48204 229278
rect 83604 229276 84204 229278
rect 119604 229276 120204 229278
rect 155604 229276 156204 229278
rect 191604 229276 192204 229278
rect 227604 229276 228204 229278
rect 263604 229276 264204 229278
rect 299604 229276 300204 229278
rect 314208 229276 314528 229278
rect 551604 229276 552204 229278
rect 590960 229276 591560 229278
rect -8576 229254 592500 229276
rect -8576 229018 -7454 229254
rect -7218 229018 11786 229254
rect 12022 229018 47786 229254
rect 48022 229018 83786 229254
rect 84022 229018 119786 229254
rect 120022 229018 155786 229254
rect 156022 229018 191786 229254
rect 192022 229018 227786 229254
rect 228022 229018 263786 229254
rect 264022 229018 299786 229254
rect 300022 229018 314250 229254
rect 314486 229018 551786 229254
rect 552022 229018 591142 229254
rect 591378 229018 592500 229254
rect -8576 228934 592500 229018
rect -8576 228698 -7454 228934
rect -7218 228698 11786 228934
rect 12022 228698 47786 228934
rect 48022 228698 83786 228934
rect 84022 228698 119786 228934
rect 120022 228698 155786 228934
rect 156022 228698 191786 228934
rect 192022 228698 227786 228934
rect 228022 228698 263786 228934
rect 264022 228698 299786 228934
rect 300022 228698 314250 228934
rect 314486 228698 551786 228934
rect 552022 228698 591142 228934
rect 591378 228698 592500 228934
rect -8576 228676 592500 228698
rect -7636 228674 -7036 228676
rect 11604 228674 12204 228676
rect 47604 228674 48204 228676
rect 83604 228674 84204 228676
rect 119604 228674 120204 228676
rect 155604 228674 156204 228676
rect 191604 228674 192204 228676
rect 227604 228674 228204 228676
rect 263604 228674 264204 228676
rect 299604 228674 300204 228676
rect 314208 228674 314528 228676
rect 551604 228674 552204 228676
rect 590960 228674 591560 228676
rect -5756 225676 -5156 225678
rect 8004 225676 8604 225678
rect 44004 225676 44604 225678
rect 80004 225676 80604 225678
rect 116004 225676 116604 225678
rect 152004 225676 152604 225678
rect 188004 225676 188604 225678
rect 224004 225676 224604 225678
rect 260004 225676 260604 225678
rect 296004 225676 296604 225678
rect 314208 225676 314528 225678
rect 548004 225676 548604 225678
rect 589080 225676 589680 225678
rect -6696 225654 590620 225676
rect -6696 225418 -5574 225654
rect -5338 225418 8186 225654
rect 8422 225418 44186 225654
rect 44422 225418 80186 225654
rect 80422 225418 116186 225654
rect 116422 225418 152186 225654
rect 152422 225418 188186 225654
rect 188422 225418 224186 225654
rect 224422 225418 260186 225654
rect 260422 225418 296186 225654
rect 296422 225418 314250 225654
rect 314486 225418 548186 225654
rect 548422 225418 589262 225654
rect 589498 225418 590620 225654
rect -6696 225334 590620 225418
rect -6696 225098 -5574 225334
rect -5338 225098 8186 225334
rect 8422 225098 44186 225334
rect 44422 225098 80186 225334
rect 80422 225098 116186 225334
rect 116422 225098 152186 225334
rect 152422 225098 188186 225334
rect 188422 225098 224186 225334
rect 224422 225098 260186 225334
rect 260422 225098 296186 225334
rect 296422 225098 314250 225334
rect 314486 225098 548186 225334
rect 548422 225098 589262 225334
rect 589498 225098 590620 225334
rect -6696 225076 590620 225098
rect -5756 225074 -5156 225076
rect 8004 225074 8604 225076
rect 44004 225074 44604 225076
rect 80004 225074 80604 225076
rect 116004 225074 116604 225076
rect 152004 225074 152604 225076
rect 188004 225074 188604 225076
rect 224004 225074 224604 225076
rect 260004 225074 260604 225076
rect 296004 225074 296604 225076
rect 314208 225074 314528 225076
rect 548004 225074 548604 225076
rect 589080 225074 589680 225076
rect -3876 222076 -3276 222078
rect 4404 222076 5004 222078
rect 40404 222076 41004 222078
rect 76404 222076 77004 222078
rect 112404 222076 113004 222078
rect 148404 222076 149004 222078
rect 184404 222076 185004 222078
rect 220404 222076 221004 222078
rect 256404 222076 257004 222078
rect 292404 222076 293004 222078
rect 314208 222076 314528 222078
rect 544404 222076 545004 222078
rect 580404 222076 581004 222078
rect 587200 222076 587800 222078
rect -4816 222054 588740 222076
rect -4816 221818 -3694 222054
rect -3458 221818 4586 222054
rect 4822 221818 40586 222054
rect 40822 221818 76586 222054
rect 76822 221818 112586 222054
rect 112822 221818 148586 222054
rect 148822 221818 184586 222054
rect 184822 221818 220586 222054
rect 220822 221818 256586 222054
rect 256822 221818 292586 222054
rect 292822 221818 314250 222054
rect 314486 221818 544586 222054
rect 544822 221818 580586 222054
rect 580822 221818 587382 222054
rect 587618 221818 588740 222054
rect -4816 221734 588740 221818
rect -4816 221498 -3694 221734
rect -3458 221498 4586 221734
rect 4822 221498 40586 221734
rect 40822 221498 76586 221734
rect 76822 221498 112586 221734
rect 112822 221498 148586 221734
rect 148822 221498 184586 221734
rect 184822 221498 220586 221734
rect 220822 221498 256586 221734
rect 256822 221498 292586 221734
rect 292822 221498 314250 221734
rect 314486 221498 544586 221734
rect 544822 221498 580586 221734
rect 580822 221498 587382 221734
rect 587618 221498 588740 221734
rect -4816 221476 588740 221498
rect -3876 221474 -3276 221476
rect 4404 221474 5004 221476
rect 40404 221474 41004 221476
rect 76404 221474 77004 221476
rect 112404 221474 113004 221476
rect 148404 221474 149004 221476
rect 184404 221474 185004 221476
rect 220404 221474 221004 221476
rect 256404 221474 257004 221476
rect 292404 221474 293004 221476
rect 314208 221474 314528 221476
rect 544404 221474 545004 221476
rect 580404 221474 581004 221476
rect 587200 221474 587800 221476
rect -1996 218476 -1396 218478
rect 804 218476 1404 218478
rect 36804 218476 37404 218478
rect 72804 218476 73404 218478
rect 108804 218476 109404 218478
rect 144804 218476 145404 218478
rect 180804 218476 181404 218478
rect 216804 218476 217404 218478
rect 252804 218476 253404 218478
rect 288804 218476 289404 218478
rect 314208 218476 314528 218478
rect 540804 218476 541404 218478
rect 576804 218476 577404 218478
rect 585320 218476 585920 218478
rect -2936 218454 586860 218476
rect -2936 218218 -1814 218454
rect -1578 218218 986 218454
rect 1222 218218 36986 218454
rect 37222 218218 72986 218454
rect 73222 218218 108986 218454
rect 109222 218218 144986 218454
rect 145222 218218 180986 218454
rect 181222 218218 216986 218454
rect 217222 218218 252986 218454
rect 253222 218218 288986 218454
rect 289222 218218 314250 218454
rect 314486 218218 540986 218454
rect 541222 218218 576986 218454
rect 577222 218218 585502 218454
rect 585738 218218 586860 218454
rect -2936 218134 586860 218218
rect -2936 217898 -1814 218134
rect -1578 217898 986 218134
rect 1222 217898 36986 218134
rect 37222 217898 72986 218134
rect 73222 217898 108986 218134
rect 109222 217898 144986 218134
rect 145222 217898 180986 218134
rect 181222 217898 216986 218134
rect 217222 217898 252986 218134
rect 253222 217898 288986 218134
rect 289222 217898 314250 218134
rect 314486 217898 540986 218134
rect 541222 217898 576986 218134
rect 577222 217898 585502 218134
rect 585738 217898 586860 218134
rect -2936 217876 586860 217898
rect -1996 217874 -1396 217876
rect 804 217874 1404 217876
rect 36804 217874 37404 217876
rect 72804 217874 73404 217876
rect 108804 217874 109404 217876
rect 144804 217874 145404 217876
rect 180804 217874 181404 217876
rect 216804 217874 217404 217876
rect 252804 217874 253404 217876
rect 288804 217874 289404 217876
rect 314208 217874 314528 217876
rect 540804 217874 541404 217876
rect 576804 217874 577404 217876
rect 585320 217874 585920 217876
rect -8576 211276 -7976 211278
rect 29604 211276 30204 211278
rect 65604 211276 66204 211278
rect 101604 211276 102204 211278
rect 137604 211276 138204 211278
rect 173604 211276 174204 211278
rect 209604 211276 210204 211278
rect 245604 211276 246204 211278
rect 281604 211276 282204 211278
rect 329568 211276 329888 211278
rect 533604 211276 534204 211278
rect 569604 211276 570204 211278
rect 591900 211276 592500 211278
rect -8576 211254 592500 211276
rect -8576 211018 -8394 211254
rect -8158 211018 29786 211254
rect 30022 211018 65786 211254
rect 66022 211018 101786 211254
rect 102022 211018 137786 211254
rect 138022 211018 173786 211254
rect 174022 211018 209786 211254
rect 210022 211018 245786 211254
rect 246022 211018 281786 211254
rect 282022 211018 329610 211254
rect 329846 211018 533786 211254
rect 534022 211018 569786 211254
rect 570022 211018 592082 211254
rect 592318 211018 592500 211254
rect -8576 210934 592500 211018
rect -8576 210698 -8394 210934
rect -8158 210698 29786 210934
rect 30022 210698 65786 210934
rect 66022 210698 101786 210934
rect 102022 210698 137786 210934
rect 138022 210698 173786 210934
rect 174022 210698 209786 210934
rect 210022 210698 245786 210934
rect 246022 210698 281786 210934
rect 282022 210698 329610 210934
rect 329846 210698 533786 210934
rect 534022 210698 569786 210934
rect 570022 210698 592082 210934
rect 592318 210698 592500 210934
rect -8576 210676 592500 210698
rect -8576 210674 -7976 210676
rect 29604 210674 30204 210676
rect 65604 210674 66204 210676
rect 101604 210674 102204 210676
rect 137604 210674 138204 210676
rect 173604 210674 174204 210676
rect 209604 210674 210204 210676
rect 245604 210674 246204 210676
rect 281604 210674 282204 210676
rect 329568 210674 329888 210676
rect 533604 210674 534204 210676
rect 569604 210674 570204 210676
rect 591900 210674 592500 210676
rect -6696 207676 -6096 207678
rect 26004 207676 26604 207678
rect 62004 207676 62604 207678
rect 98004 207676 98604 207678
rect 134004 207676 134604 207678
rect 170004 207676 170604 207678
rect 206004 207676 206604 207678
rect 242004 207676 242604 207678
rect 278004 207676 278604 207678
rect 329568 207676 329888 207678
rect 566004 207676 566604 207678
rect 590020 207676 590620 207678
rect -6696 207654 590620 207676
rect -6696 207418 -6514 207654
rect -6278 207418 26186 207654
rect 26422 207418 62186 207654
rect 62422 207418 98186 207654
rect 98422 207418 134186 207654
rect 134422 207418 170186 207654
rect 170422 207418 206186 207654
rect 206422 207418 242186 207654
rect 242422 207418 278186 207654
rect 278422 207418 329610 207654
rect 329846 207418 566186 207654
rect 566422 207418 590202 207654
rect 590438 207418 590620 207654
rect -6696 207334 590620 207418
rect -6696 207098 -6514 207334
rect -6278 207098 26186 207334
rect 26422 207098 62186 207334
rect 62422 207098 98186 207334
rect 98422 207098 134186 207334
rect 134422 207098 170186 207334
rect 170422 207098 206186 207334
rect 206422 207098 242186 207334
rect 242422 207098 278186 207334
rect 278422 207098 329610 207334
rect 329846 207098 566186 207334
rect 566422 207098 590202 207334
rect 590438 207098 590620 207334
rect -6696 207076 590620 207098
rect -6696 207074 -6096 207076
rect 26004 207074 26604 207076
rect 62004 207074 62604 207076
rect 98004 207074 98604 207076
rect 134004 207074 134604 207076
rect 170004 207074 170604 207076
rect 206004 207074 206604 207076
rect 242004 207074 242604 207076
rect 278004 207074 278604 207076
rect 329568 207074 329888 207076
rect 566004 207074 566604 207076
rect 590020 207074 590620 207076
rect -4816 204076 -4216 204078
rect 22404 204076 23004 204078
rect 58404 204076 59004 204078
rect 94404 204076 95004 204078
rect 130404 204076 131004 204078
rect 166404 204076 167004 204078
rect 202404 204076 203004 204078
rect 238404 204076 239004 204078
rect 274404 204076 275004 204078
rect 329568 204076 329888 204078
rect 562404 204076 563004 204078
rect 588140 204076 588740 204078
rect -4816 204054 588740 204076
rect -4816 203818 -4634 204054
rect -4398 203818 22586 204054
rect 22822 203818 58586 204054
rect 58822 203818 94586 204054
rect 94822 203818 130586 204054
rect 130822 203818 166586 204054
rect 166822 203818 202586 204054
rect 202822 203818 238586 204054
rect 238822 203818 274586 204054
rect 274822 203818 329610 204054
rect 329846 203818 562586 204054
rect 562822 203818 588322 204054
rect 588558 203818 588740 204054
rect -4816 203734 588740 203818
rect -4816 203498 -4634 203734
rect -4398 203498 22586 203734
rect 22822 203498 58586 203734
rect 58822 203498 94586 203734
rect 94822 203498 130586 203734
rect 130822 203498 166586 203734
rect 166822 203498 202586 203734
rect 202822 203498 238586 203734
rect 238822 203498 274586 203734
rect 274822 203498 329610 203734
rect 329846 203498 562586 203734
rect 562822 203498 588322 203734
rect 588558 203498 588740 203734
rect -4816 203476 588740 203498
rect -4816 203474 -4216 203476
rect 22404 203474 23004 203476
rect 58404 203474 59004 203476
rect 94404 203474 95004 203476
rect 130404 203474 131004 203476
rect 166404 203474 167004 203476
rect 202404 203474 203004 203476
rect 238404 203474 239004 203476
rect 274404 203474 275004 203476
rect 329568 203474 329888 203476
rect 562404 203474 563004 203476
rect 588140 203474 588740 203476
rect -2936 200476 -2336 200478
rect 18804 200476 19404 200478
rect 54804 200476 55404 200478
rect 90804 200476 91404 200478
rect 126804 200476 127404 200478
rect 162804 200476 163404 200478
rect 198804 200476 199404 200478
rect 234804 200476 235404 200478
rect 270804 200476 271404 200478
rect 329568 200476 329888 200478
rect 558804 200476 559404 200478
rect 586260 200476 586860 200478
rect -2936 200454 586860 200476
rect -2936 200218 -2754 200454
rect -2518 200218 18986 200454
rect 19222 200218 54986 200454
rect 55222 200218 90986 200454
rect 91222 200218 126986 200454
rect 127222 200218 162986 200454
rect 163222 200218 198986 200454
rect 199222 200218 234986 200454
rect 235222 200218 270986 200454
rect 271222 200218 329610 200454
rect 329846 200218 558986 200454
rect 559222 200218 586442 200454
rect 586678 200218 586860 200454
rect -2936 200134 586860 200218
rect -2936 199898 -2754 200134
rect -2518 199898 18986 200134
rect 19222 199898 54986 200134
rect 55222 199898 90986 200134
rect 91222 199898 126986 200134
rect 127222 199898 162986 200134
rect 163222 199898 198986 200134
rect 199222 199898 234986 200134
rect 235222 199898 270986 200134
rect 271222 199898 329610 200134
rect 329846 199898 558986 200134
rect 559222 199898 586442 200134
rect 586678 199898 586860 200134
rect -2936 199876 586860 199898
rect -2936 199874 -2336 199876
rect 18804 199874 19404 199876
rect 54804 199874 55404 199876
rect 90804 199874 91404 199876
rect 126804 199874 127404 199876
rect 162804 199874 163404 199876
rect 198804 199874 199404 199876
rect 234804 199874 235404 199876
rect 270804 199874 271404 199876
rect 329568 199874 329888 199876
rect 558804 199874 559404 199876
rect 586260 199874 586860 199876
rect -7636 193276 -7036 193278
rect 11604 193276 12204 193278
rect 47604 193276 48204 193278
rect 83604 193276 84204 193278
rect 119604 193276 120204 193278
rect 155604 193276 156204 193278
rect 191604 193276 192204 193278
rect 227604 193276 228204 193278
rect 263604 193276 264204 193278
rect 299604 193276 300204 193278
rect 314208 193276 314528 193278
rect 551604 193276 552204 193278
rect 590960 193276 591560 193278
rect -8576 193254 592500 193276
rect -8576 193018 -7454 193254
rect -7218 193018 11786 193254
rect 12022 193018 47786 193254
rect 48022 193018 83786 193254
rect 84022 193018 119786 193254
rect 120022 193018 155786 193254
rect 156022 193018 191786 193254
rect 192022 193018 227786 193254
rect 228022 193018 263786 193254
rect 264022 193018 299786 193254
rect 300022 193018 314250 193254
rect 314486 193018 551786 193254
rect 552022 193018 591142 193254
rect 591378 193018 592500 193254
rect -8576 192934 592500 193018
rect -8576 192698 -7454 192934
rect -7218 192698 11786 192934
rect 12022 192698 47786 192934
rect 48022 192698 83786 192934
rect 84022 192698 119786 192934
rect 120022 192698 155786 192934
rect 156022 192698 191786 192934
rect 192022 192698 227786 192934
rect 228022 192698 263786 192934
rect 264022 192698 299786 192934
rect 300022 192698 314250 192934
rect 314486 192698 551786 192934
rect 552022 192698 591142 192934
rect 591378 192698 592500 192934
rect -8576 192676 592500 192698
rect -7636 192674 -7036 192676
rect 11604 192674 12204 192676
rect 47604 192674 48204 192676
rect 83604 192674 84204 192676
rect 119604 192674 120204 192676
rect 155604 192674 156204 192676
rect 191604 192674 192204 192676
rect 227604 192674 228204 192676
rect 263604 192674 264204 192676
rect 299604 192674 300204 192676
rect 314208 192674 314528 192676
rect 551604 192674 552204 192676
rect 590960 192674 591560 192676
rect -5756 189676 -5156 189678
rect 8004 189676 8604 189678
rect 44004 189676 44604 189678
rect 80004 189676 80604 189678
rect 116004 189676 116604 189678
rect 152004 189676 152604 189678
rect 188004 189676 188604 189678
rect 224004 189676 224604 189678
rect 260004 189676 260604 189678
rect 296004 189676 296604 189678
rect 314208 189676 314528 189678
rect 548004 189676 548604 189678
rect 589080 189676 589680 189678
rect -6696 189654 590620 189676
rect -6696 189418 -5574 189654
rect -5338 189418 8186 189654
rect 8422 189418 44186 189654
rect 44422 189418 80186 189654
rect 80422 189418 116186 189654
rect 116422 189418 152186 189654
rect 152422 189418 188186 189654
rect 188422 189418 224186 189654
rect 224422 189418 260186 189654
rect 260422 189418 296186 189654
rect 296422 189418 314250 189654
rect 314486 189418 548186 189654
rect 548422 189418 589262 189654
rect 589498 189418 590620 189654
rect -6696 189334 590620 189418
rect -6696 189098 -5574 189334
rect -5338 189098 8186 189334
rect 8422 189098 44186 189334
rect 44422 189098 80186 189334
rect 80422 189098 116186 189334
rect 116422 189098 152186 189334
rect 152422 189098 188186 189334
rect 188422 189098 224186 189334
rect 224422 189098 260186 189334
rect 260422 189098 296186 189334
rect 296422 189098 314250 189334
rect 314486 189098 548186 189334
rect 548422 189098 589262 189334
rect 589498 189098 590620 189334
rect -6696 189076 590620 189098
rect -5756 189074 -5156 189076
rect 8004 189074 8604 189076
rect 44004 189074 44604 189076
rect 80004 189074 80604 189076
rect 116004 189074 116604 189076
rect 152004 189074 152604 189076
rect 188004 189074 188604 189076
rect 224004 189074 224604 189076
rect 260004 189074 260604 189076
rect 296004 189074 296604 189076
rect 314208 189074 314528 189076
rect 548004 189074 548604 189076
rect 589080 189074 589680 189076
rect -3876 186076 -3276 186078
rect 4404 186076 5004 186078
rect 40404 186076 41004 186078
rect 76404 186076 77004 186078
rect 112404 186076 113004 186078
rect 148404 186076 149004 186078
rect 184404 186076 185004 186078
rect 220404 186076 221004 186078
rect 256404 186076 257004 186078
rect 292404 186076 293004 186078
rect 314208 186076 314528 186078
rect 544404 186076 545004 186078
rect 580404 186076 581004 186078
rect 587200 186076 587800 186078
rect -4816 186054 588740 186076
rect -4816 185818 -3694 186054
rect -3458 185818 4586 186054
rect 4822 185818 40586 186054
rect 40822 185818 76586 186054
rect 76822 185818 112586 186054
rect 112822 185818 148586 186054
rect 148822 185818 184586 186054
rect 184822 185818 220586 186054
rect 220822 185818 256586 186054
rect 256822 185818 292586 186054
rect 292822 185818 314250 186054
rect 314486 185818 544586 186054
rect 544822 185818 580586 186054
rect 580822 185818 587382 186054
rect 587618 185818 588740 186054
rect -4816 185734 588740 185818
rect -4816 185498 -3694 185734
rect -3458 185498 4586 185734
rect 4822 185498 40586 185734
rect 40822 185498 76586 185734
rect 76822 185498 112586 185734
rect 112822 185498 148586 185734
rect 148822 185498 184586 185734
rect 184822 185498 220586 185734
rect 220822 185498 256586 185734
rect 256822 185498 292586 185734
rect 292822 185498 314250 185734
rect 314486 185498 544586 185734
rect 544822 185498 580586 185734
rect 580822 185498 587382 185734
rect 587618 185498 588740 185734
rect -4816 185476 588740 185498
rect -3876 185474 -3276 185476
rect 4404 185474 5004 185476
rect 40404 185474 41004 185476
rect 76404 185474 77004 185476
rect 112404 185474 113004 185476
rect 148404 185474 149004 185476
rect 184404 185474 185004 185476
rect 220404 185474 221004 185476
rect 256404 185474 257004 185476
rect 292404 185474 293004 185476
rect 314208 185474 314528 185476
rect 544404 185474 545004 185476
rect 580404 185474 581004 185476
rect 587200 185474 587800 185476
rect -1996 182476 -1396 182478
rect 804 182476 1404 182478
rect 36804 182476 37404 182478
rect 72804 182476 73404 182478
rect 108804 182476 109404 182478
rect 144804 182476 145404 182478
rect 180804 182476 181404 182478
rect 216804 182476 217404 182478
rect 252804 182476 253404 182478
rect 288804 182476 289404 182478
rect 314208 182476 314528 182478
rect 540804 182476 541404 182478
rect 576804 182476 577404 182478
rect 585320 182476 585920 182478
rect -2936 182454 586860 182476
rect -2936 182218 -1814 182454
rect -1578 182218 986 182454
rect 1222 182218 36986 182454
rect 37222 182218 72986 182454
rect 73222 182218 108986 182454
rect 109222 182218 144986 182454
rect 145222 182218 180986 182454
rect 181222 182218 216986 182454
rect 217222 182218 252986 182454
rect 253222 182218 288986 182454
rect 289222 182218 314250 182454
rect 314486 182218 540986 182454
rect 541222 182218 576986 182454
rect 577222 182218 585502 182454
rect 585738 182218 586860 182454
rect -2936 182134 586860 182218
rect -2936 181898 -1814 182134
rect -1578 181898 986 182134
rect 1222 181898 36986 182134
rect 37222 181898 72986 182134
rect 73222 181898 108986 182134
rect 109222 181898 144986 182134
rect 145222 181898 180986 182134
rect 181222 181898 216986 182134
rect 217222 181898 252986 182134
rect 253222 181898 288986 182134
rect 289222 181898 314250 182134
rect 314486 181898 540986 182134
rect 541222 181898 576986 182134
rect 577222 181898 585502 182134
rect 585738 181898 586860 182134
rect -2936 181876 586860 181898
rect -1996 181874 -1396 181876
rect 804 181874 1404 181876
rect 36804 181874 37404 181876
rect 72804 181874 73404 181876
rect 108804 181874 109404 181876
rect 144804 181874 145404 181876
rect 180804 181874 181404 181876
rect 216804 181874 217404 181876
rect 252804 181874 253404 181876
rect 288804 181874 289404 181876
rect 314208 181874 314528 181876
rect 540804 181874 541404 181876
rect 576804 181874 577404 181876
rect 585320 181874 585920 181876
rect -8576 175276 -7976 175278
rect 29604 175276 30204 175278
rect 65604 175276 66204 175278
rect 101604 175276 102204 175278
rect 137604 175276 138204 175278
rect 173604 175276 174204 175278
rect 209604 175276 210204 175278
rect 245604 175276 246204 175278
rect 281604 175276 282204 175278
rect 329568 175276 329888 175278
rect 533604 175276 534204 175278
rect 569604 175276 570204 175278
rect 591900 175276 592500 175278
rect -8576 175254 592500 175276
rect -8576 175018 -8394 175254
rect -8158 175018 29786 175254
rect 30022 175018 65786 175254
rect 66022 175018 101786 175254
rect 102022 175018 137786 175254
rect 138022 175018 173786 175254
rect 174022 175018 209786 175254
rect 210022 175018 245786 175254
rect 246022 175018 281786 175254
rect 282022 175018 329610 175254
rect 329846 175018 533786 175254
rect 534022 175018 569786 175254
rect 570022 175018 592082 175254
rect 592318 175018 592500 175254
rect -8576 174934 592500 175018
rect -8576 174698 -8394 174934
rect -8158 174698 29786 174934
rect 30022 174698 65786 174934
rect 66022 174698 101786 174934
rect 102022 174698 137786 174934
rect 138022 174698 173786 174934
rect 174022 174698 209786 174934
rect 210022 174698 245786 174934
rect 246022 174698 281786 174934
rect 282022 174698 329610 174934
rect 329846 174698 533786 174934
rect 534022 174698 569786 174934
rect 570022 174698 592082 174934
rect 592318 174698 592500 174934
rect -8576 174676 592500 174698
rect -8576 174674 -7976 174676
rect 29604 174674 30204 174676
rect 65604 174674 66204 174676
rect 101604 174674 102204 174676
rect 137604 174674 138204 174676
rect 173604 174674 174204 174676
rect 209604 174674 210204 174676
rect 245604 174674 246204 174676
rect 281604 174674 282204 174676
rect 329568 174674 329888 174676
rect 533604 174674 534204 174676
rect 569604 174674 570204 174676
rect 591900 174674 592500 174676
rect -6696 171676 -6096 171678
rect 26004 171676 26604 171678
rect 62004 171676 62604 171678
rect 98004 171676 98604 171678
rect 134004 171676 134604 171678
rect 170004 171676 170604 171678
rect 206004 171676 206604 171678
rect 242004 171676 242604 171678
rect 278004 171676 278604 171678
rect 329568 171676 329888 171678
rect 566004 171676 566604 171678
rect 590020 171676 590620 171678
rect -6696 171654 590620 171676
rect -6696 171418 -6514 171654
rect -6278 171418 26186 171654
rect 26422 171418 62186 171654
rect 62422 171418 98186 171654
rect 98422 171418 134186 171654
rect 134422 171418 170186 171654
rect 170422 171418 206186 171654
rect 206422 171418 242186 171654
rect 242422 171418 278186 171654
rect 278422 171418 329610 171654
rect 329846 171418 566186 171654
rect 566422 171418 590202 171654
rect 590438 171418 590620 171654
rect -6696 171334 590620 171418
rect -6696 171098 -6514 171334
rect -6278 171098 26186 171334
rect 26422 171098 62186 171334
rect 62422 171098 98186 171334
rect 98422 171098 134186 171334
rect 134422 171098 170186 171334
rect 170422 171098 206186 171334
rect 206422 171098 242186 171334
rect 242422 171098 278186 171334
rect 278422 171098 329610 171334
rect 329846 171098 566186 171334
rect 566422 171098 590202 171334
rect 590438 171098 590620 171334
rect -6696 171076 590620 171098
rect -6696 171074 -6096 171076
rect 26004 171074 26604 171076
rect 62004 171074 62604 171076
rect 98004 171074 98604 171076
rect 134004 171074 134604 171076
rect 170004 171074 170604 171076
rect 206004 171074 206604 171076
rect 242004 171074 242604 171076
rect 278004 171074 278604 171076
rect 329568 171074 329888 171076
rect 566004 171074 566604 171076
rect 590020 171074 590620 171076
rect -4816 168076 -4216 168078
rect 22404 168076 23004 168078
rect 58404 168076 59004 168078
rect 94404 168076 95004 168078
rect 130404 168076 131004 168078
rect 166404 168076 167004 168078
rect 202404 168076 203004 168078
rect 238404 168076 239004 168078
rect 274404 168076 275004 168078
rect 329568 168076 329888 168078
rect 562404 168076 563004 168078
rect 588140 168076 588740 168078
rect -4816 168054 588740 168076
rect -4816 167818 -4634 168054
rect -4398 167818 22586 168054
rect 22822 167818 58586 168054
rect 58822 167818 94586 168054
rect 94822 167818 130586 168054
rect 130822 167818 166586 168054
rect 166822 167818 202586 168054
rect 202822 167818 238586 168054
rect 238822 167818 274586 168054
rect 274822 167818 329610 168054
rect 329846 167818 562586 168054
rect 562822 167818 588322 168054
rect 588558 167818 588740 168054
rect -4816 167734 588740 167818
rect -4816 167498 -4634 167734
rect -4398 167498 22586 167734
rect 22822 167498 58586 167734
rect 58822 167498 94586 167734
rect 94822 167498 130586 167734
rect 130822 167498 166586 167734
rect 166822 167498 202586 167734
rect 202822 167498 238586 167734
rect 238822 167498 274586 167734
rect 274822 167498 329610 167734
rect 329846 167498 562586 167734
rect 562822 167498 588322 167734
rect 588558 167498 588740 167734
rect -4816 167476 588740 167498
rect -4816 167474 -4216 167476
rect 22404 167474 23004 167476
rect 58404 167474 59004 167476
rect 94404 167474 95004 167476
rect 130404 167474 131004 167476
rect 166404 167474 167004 167476
rect 202404 167474 203004 167476
rect 238404 167474 239004 167476
rect 274404 167474 275004 167476
rect 329568 167474 329888 167476
rect 562404 167474 563004 167476
rect 588140 167474 588740 167476
rect -2936 164476 -2336 164478
rect 18804 164476 19404 164478
rect 54804 164476 55404 164478
rect 90804 164476 91404 164478
rect 126804 164476 127404 164478
rect 162804 164476 163404 164478
rect 198804 164476 199404 164478
rect 234804 164476 235404 164478
rect 270804 164476 271404 164478
rect 329568 164476 329888 164478
rect 558804 164476 559404 164478
rect 586260 164476 586860 164478
rect -2936 164454 586860 164476
rect -2936 164218 -2754 164454
rect -2518 164218 18986 164454
rect 19222 164218 54986 164454
rect 55222 164218 90986 164454
rect 91222 164218 126986 164454
rect 127222 164218 162986 164454
rect 163222 164218 198986 164454
rect 199222 164218 234986 164454
rect 235222 164218 270986 164454
rect 271222 164218 329610 164454
rect 329846 164218 558986 164454
rect 559222 164218 586442 164454
rect 586678 164218 586860 164454
rect -2936 164134 586860 164218
rect -2936 163898 -2754 164134
rect -2518 163898 18986 164134
rect 19222 163898 54986 164134
rect 55222 163898 90986 164134
rect 91222 163898 126986 164134
rect 127222 163898 162986 164134
rect 163222 163898 198986 164134
rect 199222 163898 234986 164134
rect 235222 163898 270986 164134
rect 271222 163898 329610 164134
rect 329846 163898 558986 164134
rect 559222 163898 586442 164134
rect 586678 163898 586860 164134
rect -2936 163876 586860 163898
rect -2936 163874 -2336 163876
rect 18804 163874 19404 163876
rect 54804 163874 55404 163876
rect 90804 163874 91404 163876
rect 126804 163874 127404 163876
rect 162804 163874 163404 163876
rect 198804 163874 199404 163876
rect 234804 163874 235404 163876
rect 270804 163874 271404 163876
rect 329568 163874 329888 163876
rect 558804 163874 559404 163876
rect 586260 163874 586860 163876
rect -7636 157276 -7036 157278
rect 11604 157276 12204 157278
rect 47604 157276 48204 157278
rect 83604 157276 84204 157278
rect 119604 157276 120204 157278
rect 155604 157276 156204 157278
rect 191604 157276 192204 157278
rect 227604 157276 228204 157278
rect 263604 157276 264204 157278
rect 299604 157276 300204 157278
rect 314208 157276 314528 157278
rect 551604 157276 552204 157278
rect 590960 157276 591560 157278
rect -8576 157254 592500 157276
rect -8576 157018 -7454 157254
rect -7218 157018 11786 157254
rect 12022 157018 47786 157254
rect 48022 157018 83786 157254
rect 84022 157018 119786 157254
rect 120022 157018 155786 157254
rect 156022 157018 191786 157254
rect 192022 157018 227786 157254
rect 228022 157018 263786 157254
rect 264022 157018 299786 157254
rect 300022 157018 314250 157254
rect 314486 157018 551786 157254
rect 552022 157018 591142 157254
rect 591378 157018 592500 157254
rect -8576 156934 592500 157018
rect -8576 156698 -7454 156934
rect -7218 156698 11786 156934
rect 12022 156698 47786 156934
rect 48022 156698 83786 156934
rect 84022 156698 119786 156934
rect 120022 156698 155786 156934
rect 156022 156698 191786 156934
rect 192022 156698 227786 156934
rect 228022 156698 263786 156934
rect 264022 156698 299786 156934
rect 300022 156698 314250 156934
rect 314486 156698 551786 156934
rect 552022 156698 591142 156934
rect 591378 156698 592500 156934
rect -8576 156676 592500 156698
rect -7636 156674 -7036 156676
rect 11604 156674 12204 156676
rect 47604 156674 48204 156676
rect 83604 156674 84204 156676
rect 119604 156674 120204 156676
rect 155604 156674 156204 156676
rect 191604 156674 192204 156676
rect 227604 156674 228204 156676
rect 263604 156674 264204 156676
rect 299604 156674 300204 156676
rect 314208 156674 314528 156676
rect 551604 156674 552204 156676
rect 590960 156674 591560 156676
rect -5756 153676 -5156 153678
rect 8004 153676 8604 153678
rect 44004 153676 44604 153678
rect 80004 153676 80604 153678
rect 116004 153676 116604 153678
rect 152004 153676 152604 153678
rect 188004 153676 188604 153678
rect 224004 153676 224604 153678
rect 260004 153676 260604 153678
rect 296004 153676 296604 153678
rect 314208 153676 314528 153678
rect 548004 153676 548604 153678
rect 589080 153676 589680 153678
rect -6696 153654 590620 153676
rect -6696 153418 -5574 153654
rect -5338 153418 8186 153654
rect 8422 153418 44186 153654
rect 44422 153418 80186 153654
rect 80422 153418 116186 153654
rect 116422 153418 152186 153654
rect 152422 153418 188186 153654
rect 188422 153418 224186 153654
rect 224422 153418 260186 153654
rect 260422 153418 296186 153654
rect 296422 153418 314250 153654
rect 314486 153418 548186 153654
rect 548422 153418 589262 153654
rect 589498 153418 590620 153654
rect -6696 153334 590620 153418
rect -6696 153098 -5574 153334
rect -5338 153098 8186 153334
rect 8422 153098 44186 153334
rect 44422 153098 80186 153334
rect 80422 153098 116186 153334
rect 116422 153098 152186 153334
rect 152422 153098 188186 153334
rect 188422 153098 224186 153334
rect 224422 153098 260186 153334
rect 260422 153098 296186 153334
rect 296422 153098 314250 153334
rect 314486 153098 548186 153334
rect 548422 153098 589262 153334
rect 589498 153098 590620 153334
rect -6696 153076 590620 153098
rect -5756 153074 -5156 153076
rect 8004 153074 8604 153076
rect 44004 153074 44604 153076
rect 80004 153074 80604 153076
rect 116004 153074 116604 153076
rect 152004 153074 152604 153076
rect 188004 153074 188604 153076
rect 224004 153074 224604 153076
rect 260004 153074 260604 153076
rect 296004 153074 296604 153076
rect 314208 153074 314528 153076
rect 548004 153074 548604 153076
rect 589080 153074 589680 153076
rect -3876 150076 -3276 150078
rect 4404 150076 5004 150078
rect 40404 150076 41004 150078
rect 76404 150076 77004 150078
rect 112404 150076 113004 150078
rect 148404 150076 149004 150078
rect 184404 150076 185004 150078
rect 220404 150076 221004 150078
rect 256404 150076 257004 150078
rect 292404 150076 293004 150078
rect 314208 150076 314528 150078
rect 544404 150076 545004 150078
rect 580404 150076 581004 150078
rect 587200 150076 587800 150078
rect -4816 150054 588740 150076
rect -4816 149818 -3694 150054
rect -3458 149818 4586 150054
rect 4822 149818 40586 150054
rect 40822 149818 76586 150054
rect 76822 149818 112586 150054
rect 112822 149818 148586 150054
rect 148822 149818 184586 150054
rect 184822 149818 220586 150054
rect 220822 149818 256586 150054
rect 256822 149818 292586 150054
rect 292822 149818 314250 150054
rect 314486 149818 544586 150054
rect 544822 149818 580586 150054
rect 580822 149818 587382 150054
rect 587618 149818 588740 150054
rect -4816 149734 588740 149818
rect -4816 149498 -3694 149734
rect -3458 149498 4586 149734
rect 4822 149498 40586 149734
rect 40822 149498 76586 149734
rect 76822 149498 112586 149734
rect 112822 149498 148586 149734
rect 148822 149498 184586 149734
rect 184822 149498 220586 149734
rect 220822 149498 256586 149734
rect 256822 149498 292586 149734
rect 292822 149498 314250 149734
rect 314486 149498 544586 149734
rect 544822 149498 580586 149734
rect 580822 149498 587382 149734
rect 587618 149498 588740 149734
rect -4816 149476 588740 149498
rect -3876 149474 -3276 149476
rect 4404 149474 5004 149476
rect 40404 149474 41004 149476
rect 76404 149474 77004 149476
rect 112404 149474 113004 149476
rect 148404 149474 149004 149476
rect 184404 149474 185004 149476
rect 220404 149474 221004 149476
rect 256404 149474 257004 149476
rect 292404 149474 293004 149476
rect 314208 149474 314528 149476
rect 544404 149474 545004 149476
rect 580404 149474 581004 149476
rect 587200 149474 587800 149476
rect -1996 146476 -1396 146478
rect 804 146476 1404 146478
rect 36804 146476 37404 146478
rect 72804 146476 73404 146478
rect 108804 146476 109404 146478
rect 144804 146476 145404 146478
rect 180804 146476 181404 146478
rect 216804 146476 217404 146478
rect 252804 146476 253404 146478
rect 288804 146476 289404 146478
rect 314208 146476 314528 146478
rect 540804 146476 541404 146478
rect 576804 146476 577404 146478
rect 585320 146476 585920 146478
rect -2936 146454 586860 146476
rect -2936 146218 -1814 146454
rect -1578 146218 986 146454
rect 1222 146218 36986 146454
rect 37222 146218 72986 146454
rect 73222 146218 108986 146454
rect 109222 146218 144986 146454
rect 145222 146218 180986 146454
rect 181222 146218 216986 146454
rect 217222 146218 252986 146454
rect 253222 146218 288986 146454
rect 289222 146218 314250 146454
rect 314486 146218 540986 146454
rect 541222 146218 576986 146454
rect 577222 146218 585502 146454
rect 585738 146218 586860 146454
rect -2936 146134 586860 146218
rect -2936 145898 -1814 146134
rect -1578 145898 986 146134
rect 1222 145898 36986 146134
rect 37222 145898 72986 146134
rect 73222 145898 108986 146134
rect 109222 145898 144986 146134
rect 145222 145898 180986 146134
rect 181222 145898 216986 146134
rect 217222 145898 252986 146134
rect 253222 145898 288986 146134
rect 289222 145898 314250 146134
rect 314486 145898 540986 146134
rect 541222 145898 576986 146134
rect 577222 145898 585502 146134
rect 585738 145898 586860 146134
rect -2936 145876 586860 145898
rect -1996 145874 -1396 145876
rect 804 145874 1404 145876
rect 36804 145874 37404 145876
rect 72804 145874 73404 145876
rect 108804 145874 109404 145876
rect 144804 145874 145404 145876
rect 180804 145874 181404 145876
rect 216804 145874 217404 145876
rect 252804 145874 253404 145876
rect 288804 145874 289404 145876
rect 314208 145874 314528 145876
rect 540804 145874 541404 145876
rect 576804 145874 577404 145876
rect 585320 145874 585920 145876
rect -8576 139276 -7976 139278
rect 29604 139276 30204 139278
rect 65604 139276 66204 139278
rect 101604 139276 102204 139278
rect 137604 139276 138204 139278
rect 173604 139276 174204 139278
rect 209604 139276 210204 139278
rect 245604 139276 246204 139278
rect 281604 139276 282204 139278
rect 329568 139276 329888 139278
rect 533604 139276 534204 139278
rect 569604 139276 570204 139278
rect 591900 139276 592500 139278
rect -8576 139254 592500 139276
rect -8576 139018 -8394 139254
rect -8158 139018 29786 139254
rect 30022 139018 65786 139254
rect 66022 139018 101786 139254
rect 102022 139018 137786 139254
rect 138022 139018 173786 139254
rect 174022 139018 209786 139254
rect 210022 139018 245786 139254
rect 246022 139018 281786 139254
rect 282022 139018 329610 139254
rect 329846 139018 533786 139254
rect 534022 139018 569786 139254
rect 570022 139018 592082 139254
rect 592318 139018 592500 139254
rect -8576 138934 592500 139018
rect -8576 138698 -8394 138934
rect -8158 138698 29786 138934
rect 30022 138698 65786 138934
rect 66022 138698 101786 138934
rect 102022 138698 137786 138934
rect 138022 138698 173786 138934
rect 174022 138698 209786 138934
rect 210022 138698 245786 138934
rect 246022 138698 281786 138934
rect 282022 138698 329610 138934
rect 329846 138698 533786 138934
rect 534022 138698 569786 138934
rect 570022 138698 592082 138934
rect 592318 138698 592500 138934
rect -8576 138676 592500 138698
rect -8576 138674 -7976 138676
rect 29604 138674 30204 138676
rect 65604 138674 66204 138676
rect 101604 138674 102204 138676
rect 137604 138674 138204 138676
rect 173604 138674 174204 138676
rect 209604 138674 210204 138676
rect 245604 138674 246204 138676
rect 281604 138674 282204 138676
rect 329568 138674 329888 138676
rect 533604 138674 534204 138676
rect 569604 138674 570204 138676
rect 591900 138674 592500 138676
rect -6696 135676 -6096 135678
rect 26004 135676 26604 135678
rect 62004 135676 62604 135678
rect 98004 135676 98604 135678
rect 134004 135676 134604 135678
rect 170004 135676 170604 135678
rect 206004 135676 206604 135678
rect 242004 135676 242604 135678
rect 278004 135676 278604 135678
rect 329568 135676 329888 135678
rect 566004 135676 566604 135678
rect 590020 135676 590620 135678
rect -6696 135654 590620 135676
rect -6696 135418 -6514 135654
rect -6278 135418 26186 135654
rect 26422 135418 62186 135654
rect 62422 135418 98186 135654
rect 98422 135418 134186 135654
rect 134422 135418 170186 135654
rect 170422 135418 206186 135654
rect 206422 135418 242186 135654
rect 242422 135418 278186 135654
rect 278422 135418 329610 135654
rect 329846 135418 566186 135654
rect 566422 135418 590202 135654
rect 590438 135418 590620 135654
rect -6696 135334 590620 135418
rect -6696 135098 -6514 135334
rect -6278 135098 26186 135334
rect 26422 135098 62186 135334
rect 62422 135098 98186 135334
rect 98422 135098 134186 135334
rect 134422 135098 170186 135334
rect 170422 135098 206186 135334
rect 206422 135098 242186 135334
rect 242422 135098 278186 135334
rect 278422 135098 329610 135334
rect 329846 135098 566186 135334
rect 566422 135098 590202 135334
rect 590438 135098 590620 135334
rect -6696 135076 590620 135098
rect -6696 135074 -6096 135076
rect 26004 135074 26604 135076
rect 62004 135074 62604 135076
rect 98004 135074 98604 135076
rect 134004 135074 134604 135076
rect 170004 135074 170604 135076
rect 206004 135074 206604 135076
rect 242004 135074 242604 135076
rect 278004 135074 278604 135076
rect 329568 135074 329888 135076
rect 566004 135074 566604 135076
rect 590020 135074 590620 135076
rect -4816 132076 -4216 132078
rect 22404 132076 23004 132078
rect 58404 132076 59004 132078
rect 94404 132076 95004 132078
rect 130404 132076 131004 132078
rect 166404 132076 167004 132078
rect 202404 132076 203004 132078
rect 238404 132076 239004 132078
rect 274404 132076 275004 132078
rect 329568 132076 329888 132078
rect 562404 132076 563004 132078
rect 588140 132076 588740 132078
rect -4816 132054 588740 132076
rect -4816 131818 -4634 132054
rect -4398 131818 22586 132054
rect 22822 131818 58586 132054
rect 58822 131818 94586 132054
rect 94822 131818 130586 132054
rect 130822 131818 166586 132054
rect 166822 131818 202586 132054
rect 202822 131818 238586 132054
rect 238822 131818 274586 132054
rect 274822 131818 329610 132054
rect 329846 131818 562586 132054
rect 562822 131818 588322 132054
rect 588558 131818 588740 132054
rect -4816 131734 588740 131818
rect -4816 131498 -4634 131734
rect -4398 131498 22586 131734
rect 22822 131498 58586 131734
rect 58822 131498 94586 131734
rect 94822 131498 130586 131734
rect 130822 131498 166586 131734
rect 166822 131498 202586 131734
rect 202822 131498 238586 131734
rect 238822 131498 274586 131734
rect 274822 131498 329610 131734
rect 329846 131498 562586 131734
rect 562822 131498 588322 131734
rect 588558 131498 588740 131734
rect -4816 131476 588740 131498
rect -4816 131474 -4216 131476
rect 22404 131474 23004 131476
rect 58404 131474 59004 131476
rect 94404 131474 95004 131476
rect 130404 131474 131004 131476
rect 166404 131474 167004 131476
rect 202404 131474 203004 131476
rect 238404 131474 239004 131476
rect 274404 131474 275004 131476
rect 329568 131474 329888 131476
rect 562404 131474 563004 131476
rect 588140 131474 588740 131476
rect -2936 128476 -2336 128478
rect 18804 128476 19404 128478
rect 54804 128476 55404 128478
rect 90804 128476 91404 128478
rect 126804 128476 127404 128478
rect 162804 128476 163404 128478
rect 198804 128476 199404 128478
rect 234804 128476 235404 128478
rect 270804 128476 271404 128478
rect 329568 128476 329888 128478
rect 558804 128476 559404 128478
rect 586260 128476 586860 128478
rect -2936 128454 586860 128476
rect -2936 128218 -2754 128454
rect -2518 128218 18986 128454
rect 19222 128218 54986 128454
rect 55222 128218 90986 128454
rect 91222 128218 126986 128454
rect 127222 128218 162986 128454
rect 163222 128218 198986 128454
rect 199222 128218 234986 128454
rect 235222 128218 270986 128454
rect 271222 128218 329610 128454
rect 329846 128218 558986 128454
rect 559222 128218 586442 128454
rect 586678 128218 586860 128454
rect -2936 128134 586860 128218
rect -2936 127898 -2754 128134
rect -2518 127898 18986 128134
rect 19222 127898 54986 128134
rect 55222 127898 90986 128134
rect 91222 127898 126986 128134
rect 127222 127898 162986 128134
rect 163222 127898 198986 128134
rect 199222 127898 234986 128134
rect 235222 127898 270986 128134
rect 271222 127898 329610 128134
rect 329846 127898 558986 128134
rect 559222 127898 586442 128134
rect 586678 127898 586860 128134
rect -2936 127876 586860 127898
rect -2936 127874 -2336 127876
rect 18804 127874 19404 127876
rect 54804 127874 55404 127876
rect 90804 127874 91404 127876
rect 126804 127874 127404 127876
rect 162804 127874 163404 127876
rect 198804 127874 199404 127876
rect 234804 127874 235404 127876
rect 270804 127874 271404 127876
rect 329568 127874 329888 127876
rect 558804 127874 559404 127876
rect 586260 127874 586860 127876
rect -7636 121276 -7036 121278
rect 11604 121276 12204 121278
rect 47604 121276 48204 121278
rect 83604 121276 84204 121278
rect 119604 121276 120204 121278
rect 155604 121276 156204 121278
rect 191604 121276 192204 121278
rect 227604 121276 228204 121278
rect 263604 121276 264204 121278
rect 299604 121276 300204 121278
rect 314208 121276 314528 121278
rect 551604 121276 552204 121278
rect 590960 121276 591560 121278
rect -8576 121254 592500 121276
rect -8576 121018 -7454 121254
rect -7218 121018 11786 121254
rect 12022 121018 47786 121254
rect 48022 121018 83786 121254
rect 84022 121018 119786 121254
rect 120022 121018 155786 121254
rect 156022 121018 191786 121254
rect 192022 121018 227786 121254
rect 228022 121018 263786 121254
rect 264022 121018 299786 121254
rect 300022 121018 314250 121254
rect 314486 121018 551786 121254
rect 552022 121018 591142 121254
rect 591378 121018 592500 121254
rect -8576 120934 592500 121018
rect -8576 120698 -7454 120934
rect -7218 120698 11786 120934
rect 12022 120698 47786 120934
rect 48022 120698 83786 120934
rect 84022 120698 119786 120934
rect 120022 120698 155786 120934
rect 156022 120698 191786 120934
rect 192022 120698 227786 120934
rect 228022 120698 263786 120934
rect 264022 120698 299786 120934
rect 300022 120698 314250 120934
rect 314486 120698 551786 120934
rect 552022 120698 591142 120934
rect 591378 120698 592500 120934
rect -8576 120676 592500 120698
rect -7636 120674 -7036 120676
rect 11604 120674 12204 120676
rect 47604 120674 48204 120676
rect 83604 120674 84204 120676
rect 119604 120674 120204 120676
rect 155604 120674 156204 120676
rect 191604 120674 192204 120676
rect 227604 120674 228204 120676
rect 263604 120674 264204 120676
rect 299604 120674 300204 120676
rect 314208 120674 314528 120676
rect 551604 120674 552204 120676
rect 590960 120674 591560 120676
rect -5756 117676 -5156 117678
rect 8004 117676 8604 117678
rect 44004 117676 44604 117678
rect 80004 117676 80604 117678
rect 116004 117676 116604 117678
rect 152004 117676 152604 117678
rect 188004 117676 188604 117678
rect 224004 117676 224604 117678
rect 260004 117676 260604 117678
rect 296004 117676 296604 117678
rect 314208 117676 314528 117678
rect 548004 117676 548604 117678
rect 589080 117676 589680 117678
rect -6696 117654 590620 117676
rect -6696 117418 -5574 117654
rect -5338 117418 8186 117654
rect 8422 117418 44186 117654
rect 44422 117418 80186 117654
rect 80422 117418 116186 117654
rect 116422 117418 152186 117654
rect 152422 117418 188186 117654
rect 188422 117418 224186 117654
rect 224422 117418 260186 117654
rect 260422 117418 296186 117654
rect 296422 117418 314250 117654
rect 314486 117418 548186 117654
rect 548422 117418 589262 117654
rect 589498 117418 590620 117654
rect -6696 117334 590620 117418
rect -6696 117098 -5574 117334
rect -5338 117098 8186 117334
rect 8422 117098 44186 117334
rect 44422 117098 80186 117334
rect 80422 117098 116186 117334
rect 116422 117098 152186 117334
rect 152422 117098 188186 117334
rect 188422 117098 224186 117334
rect 224422 117098 260186 117334
rect 260422 117098 296186 117334
rect 296422 117098 314250 117334
rect 314486 117098 548186 117334
rect 548422 117098 589262 117334
rect 589498 117098 590620 117334
rect -6696 117076 590620 117098
rect -5756 117074 -5156 117076
rect 8004 117074 8604 117076
rect 44004 117074 44604 117076
rect 80004 117074 80604 117076
rect 116004 117074 116604 117076
rect 152004 117074 152604 117076
rect 188004 117074 188604 117076
rect 224004 117074 224604 117076
rect 260004 117074 260604 117076
rect 296004 117074 296604 117076
rect 314208 117074 314528 117076
rect 548004 117074 548604 117076
rect 589080 117074 589680 117076
rect -3876 114076 -3276 114078
rect 4404 114076 5004 114078
rect 40404 114076 41004 114078
rect 76404 114076 77004 114078
rect 112404 114076 113004 114078
rect 148404 114076 149004 114078
rect 184404 114076 185004 114078
rect 220404 114076 221004 114078
rect 256404 114076 257004 114078
rect 292404 114076 293004 114078
rect 314208 114076 314528 114078
rect 544404 114076 545004 114078
rect 580404 114076 581004 114078
rect 587200 114076 587800 114078
rect -4816 114054 588740 114076
rect -4816 113818 -3694 114054
rect -3458 113818 4586 114054
rect 4822 113818 40586 114054
rect 40822 113818 76586 114054
rect 76822 113818 112586 114054
rect 112822 113818 148586 114054
rect 148822 113818 184586 114054
rect 184822 113818 220586 114054
rect 220822 113818 256586 114054
rect 256822 113818 292586 114054
rect 292822 113818 314250 114054
rect 314486 113818 544586 114054
rect 544822 113818 580586 114054
rect 580822 113818 587382 114054
rect 587618 113818 588740 114054
rect -4816 113734 588740 113818
rect -4816 113498 -3694 113734
rect -3458 113498 4586 113734
rect 4822 113498 40586 113734
rect 40822 113498 76586 113734
rect 76822 113498 112586 113734
rect 112822 113498 148586 113734
rect 148822 113498 184586 113734
rect 184822 113498 220586 113734
rect 220822 113498 256586 113734
rect 256822 113498 292586 113734
rect 292822 113498 314250 113734
rect 314486 113498 544586 113734
rect 544822 113498 580586 113734
rect 580822 113498 587382 113734
rect 587618 113498 588740 113734
rect -4816 113476 588740 113498
rect -3876 113474 -3276 113476
rect 4404 113474 5004 113476
rect 40404 113474 41004 113476
rect 76404 113474 77004 113476
rect 112404 113474 113004 113476
rect 148404 113474 149004 113476
rect 184404 113474 185004 113476
rect 220404 113474 221004 113476
rect 256404 113474 257004 113476
rect 292404 113474 293004 113476
rect 314208 113474 314528 113476
rect 544404 113474 545004 113476
rect 580404 113474 581004 113476
rect 587200 113474 587800 113476
rect -1996 110476 -1396 110478
rect 804 110476 1404 110478
rect 36804 110476 37404 110478
rect 72804 110476 73404 110478
rect 108804 110476 109404 110478
rect 144804 110476 145404 110478
rect 180804 110476 181404 110478
rect 216804 110476 217404 110478
rect 252804 110476 253404 110478
rect 288804 110476 289404 110478
rect 314208 110476 314528 110478
rect 540804 110476 541404 110478
rect 576804 110476 577404 110478
rect 585320 110476 585920 110478
rect -2936 110454 586860 110476
rect -2936 110218 -1814 110454
rect -1578 110218 986 110454
rect 1222 110218 36986 110454
rect 37222 110218 72986 110454
rect 73222 110218 108986 110454
rect 109222 110218 144986 110454
rect 145222 110218 180986 110454
rect 181222 110218 216986 110454
rect 217222 110218 252986 110454
rect 253222 110218 288986 110454
rect 289222 110218 314250 110454
rect 314486 110218 540986 110454
rect 541222 110218 576986 110454
rect 577222 110218 585502 110454
rect 585738 110218 586860 110454
rect -2936 110134 586860 110218
rect -2936 109898 -1814 110134
rect -1578 109898 986 110134
rect 1222 109898 36986 110134
rect 37222 109898 72986 110134
rect 73222 109898 108986 110134
rect 109222 109898 144986 110134
rect 145222 109898 180986 110134
rect 181222 109898 216986 110134
rect 217222 109898 252986 110134
rect 253222 109898 288986 110134
rect 289222 109898 314250 110134
rect 314486 109898 540986 110134
rect 541222 109898 576986 110134
rect 577222 109898 585502 110134
rect 585738 109898 586860 110134
rect -2936 109876 586860 109898
rect -1996 109874 -1396 109876
rect 804 109874 1404 109876
rect 36804 109874 37404 109876
rect 72804 109874 73404 109876
rect 108804 109874 109404 109876
rect 144804 109874 145404 109876
rect 180804 109874 181404 109876
rect 216804 109874 217404 109876
rect 252804 109874 253404 109876
rect 288804 109874 289404 109876
rect 314208 109874 314528 109876
rect 540804 109874 541404 109876
rect 576804 109874 577404 109876
rect 585320 109874 585920 109876
rect -8576 103276 -7976 103278
rect 29604 103276 30204 103278
rect 65604 103276 66204 103278
rect 101604 103276 102204 103278
rect 137604 103276 138204 103278
rect 173604 103276 174204 103278
rect 209604 103276 210204 103278
rect 245604 103276 246204 103278
rect 281604 103276 282204 103278
rect 329568 103276 329888 103278
rect 533604 103276 534204 103278
rect 569604 103276 570204 103278
rect 591900 103276 592500 103278
rect -8576 103254 592500 103276
rect -8576 103018 -8394 103254
rect -8158 103018 29786 103254
rect 30022 103018 65786 103254
rect 66022 103018 101786 103254
rect 102022 103018 137786 103254
rect 138022 103018 173786 103254
rect 174022 103018 209786 103254
rect 210022 103018 245786 103254
rect 246022 103018 281786 103254
rect 282022 103018 329610 103254
rect 329846 103018 533786 103254
rect 534022 103018 569786 103254
rect 570022 103018 592082 103254
rect 592318 103018 592500 103254
rect -8576 102934 592500 103018
rect -8576 102698 -8394 102934
rect -8158 102698 29786 102934
rect 30022 102698 65786 102934
rect 66022 102698 101786 102934
rect 102022 102698 137786 102934
rect 138022 102698 173786 102934
rect 174022 102698 209786 102934
rect 210022 102698 245786 102934
rect 246022 102698 281786 102934
rect 282022 102698 329610 102934
rect 329846 102698 533786 102934
rect 534022 102698 569786 102934
rect 570022 102698 592082 102934
rect 592318 102698 592500 102934
rect -8576 102676 592500 102698
rect -8576 102674 -7976 102676
rect 29604 102674 30204 102676
rect 65604 102674 66204 102676
rect 101604 102674 102204 102676
rect 137604 102674 138204 102676
rect 173604 102674 174204 102676
rect 209604 102674 210204 102676
rect 245604 102674 246204 102676
rect 281604 102674 282204 102676
rect 329568 102674 329888 102676
rect 533604 102674 534204 102676
rect 569604 102674 570204 102676
rect 591900 102674 592500 102676
rect -6696 99676 -6096 99678
rect 26004 99676 26604 99678
rect 62004 99676 62604 99678
rect 98004 99676 98604 99678
rect 134004 99676 134604 99678
rect 170004 99676 170604 99678
rect 206004 99676 206604 99678
rect 242004 99676 242604 99678
rect 278004 99676 278604 99678
rect 329568 99676 329888 99678
rect 566004 99676 566604 99678
rect 590020 99676 590620 99678
rect -6696 99654 590620 99676
rect -6696 99418 -6514 99654
rect -6278 99418 26186 99654
rect 26422 99418 62186 99654
rect 62422 99418 98186 99654
rect 98422 99418 134186 99654
rect 134422 99418 170186 99654
rect 170422 99418 206186 99654
rect 206422 99418 242186 99654
rect 242422 99418 278186 99654
rect 278422 99418 329610 99654
rect 329846 99418 566186 99654
rect 566422 99418 590202 99654
rect 590438 99418 590620 99654
rect -6696 99334 590620 99418
rect -6696 99098 -6514 99334
rect -6278 99098 26186 99334
rect 26422 99098 62186 99334
rect 62422 99098 98186 99334
rect 98422 99098 134186 99334
rect 134422 99098 170186 99334
rect 170422 99098 206186 99334
rect 206422 99098 242186 99334
rect 242422 99098 278186 99334
rect 278422 99098 329610 99334
rect 329846 99098 566186 99334
rect 566422 99098 590202 99334
rect 590438 99098 590620 99334
rect -6696 99076 590620 99098
rect -6696 99074 -6096 99076
rect 26004 99074 26604 99076
rect 62004 99074 62604 99076
rect 98004 99074 98604 99076
rect 134004 99074 134604 99076
rect 170004 99074 170604 99076
rect 206004 99074 206604 99076
rect 242004 99074 242604 99076
rect 278004 99074 278604 99076
rect 329568 99074 329888 99076
rect 566004 99074 566604 99076
rect 590020 99074 590620 99076
rect -4816 96076 -4216 96078
rect 22404 96076 23004 96078
rect 58404 96076 59004 96078
rect 94404 96076 95004 96078
rect 130404 96076 131004 96078
rect 166404 96076 167004 96078
rect 202404 96076 203004 96078
rect 238404 96076 239004 96078
rect 274404 96076 275004 96078
rect 329568 96076 329888 96078
rect 562404 96076 563004 96078
rect 588140 96076 588740 96078
rect -4816 96054 588740 96076
rect -4816 95818 -4634 96054
rect -4398 95818 22586 96054
rect 22822 95818 58586 96054
rect 58822 95818 94586 96054
rect 94822 95818 130586 96054
rect 130822 95818 166586 96054
rect 166822 95818 202586 96054
rect 202822 95818 238586 96054
rect 238822 95818 274586 96054
rect 274822 95818 329610 96054
rect 329846 95818 562586 96054
rect 562822 95818 588322 96054
rect 588558 95818 588740 96054
rect -4816 95734 588740 95818
rect -4816 95498 -4634 95734
rect -4398 95498 22586 95734
rect 22822 95498 58586 95734
rect 58822 95498 94586 95734
rect 94822 95498 130586 95734
rect 130822 95498 166586 95734
rect 166822 95498 202586 95734
rect 202822 95498 238586 95734
rect 238822 95498 274586 95734
rect 274822 95498 329610 95734
rect 329846 95498 562586 95734
rect 562822 95498 588322 95734
rect 588558 95498 588740 95734
rect -4816 95476 588740 95498
rect -4816 95474 -4216 95476
rect 22404 95474 23004 95476
rect 58404 95474 59004 95476
rect 94404 95474 95004 95476
rect 130404 95474 131004 95476
rect 166404 95474 167004 95476
rect 202404 95474 203004 95476
rect 238404 95474 239004 95476
rect 274404 95474 275004 95476
rect 329568 95474 329888 95476
rect 562404 95474 563004 95476
rect 588140 95474 588740 95476
rect -2936 92476 -2336 92478
rect 18804 92476 19404 92478
rect 54804 92476 55404 92478
rect 90804 92476 91404 92478
rect 126804 92476 127404 92478
rect 162804 92476 163404 92478
rect 198804 92476 199404 92478
rect 234804 92476 235404 92478
rect 270804 92476 271404 92478
rect 329568 92476 329888 92478
rect 558804 92476 559404 92478
rect 586260 92476 586860 92478
rect -2936 92454 586860 92476
rect -2936 92218 -2754 92454
rect -2518 92218 18986 92454
rect 19222 92218 54986 92454
rect 55222 92218 90986 92454
rect 91222 92218 126986 92454
rect 127222 92218 162986 92454
rect 163222 92218 198986 92454
rect 199222 92218 234986 92454
rect 235222 92218 270986 92454
rect 271222 92218 329610 92454
rect 329846 92218 558986 92454
rect 559222 92218 586442 92454
rect 586678 92218 586860 92454
rect -2936 92134 586860 92218
rect -2936 91898 -2754 92134
rect -2518 91898 18986 92134
rect 19222 91898 54986 92134
rect 55222 91898 90986 92134
rect 91222 91898 126986 92134
rect 127222 91898 162986 92134
rect 163222 91898 198986 92134
rect 199222 91898 234986 92134
rect 235222 91898 270986 92134
rect 271222 91898 329610 92134
rect 329846 91898 558986 92134
rect 559222 91898 586442 92134
rect 586678 91898 586860 92134
rect -2936 91876 586860 91898
rect -2936 91874 -2336 91876
rect 18804 91874 19404 91876
rect 54804 91874 55404 91876
rect 90804 91874 91404 91876
rect 126804 91874 127404 91876
rect 162804 91874 163404 91876
rect 198804 91874 199404 91876
rect 234804 91874 235404 91876
rect 270804 91874 271404 91876
rect 329568 91874 329888 91876
rect 558804 91874 559404 91876
rect 586260 91874 586860 91876
rect -7636 85276 -7036 85278
rect 11604 85276 12204 85278
rect 47604 85276 48204 85278
rect 83604 85276 84204 85278
rect 119604 85276 120204 85278
rect 155604 85276 156204 85278
rect 191604 85276 192204 85278
rect 227604 85276 228204 85278
rect 263604 85276 264204 85278
rect 299604 85276 300204 85278
rect 314208 85276 314528 85278
rect 551604 85276 552204 85278
rect 590960 85276 591560 85278
rect -8576 85254 592500 85276
rect -8576 85018 -7454 85254
rect -7218 85018 11786 85254
rect 12022 85018 47786 85254
rect 48022 85018 83786 85254
rect 84022 85018 119786 85254
rect 120022 85018 155786 85254
rect 156022 85018 191786 85254
rect 192022 85018 227786 85254
rect 228022 85018 263786 85254
rect 264022 85018 299786 85254
rect 300022 85018 314250 85254
rect 314486 85018 551786 85254
rect 552022 85018 591142 85254
rect 591378 85018 592500 85254
rect -8576 84934 592500 85018
rect -8576 84698 -7454 84934
rect -7218 84698 11786 84934
rect 12022 84698 47786 84934
rect 48022 84698 83786 84934
rect 84022 84698 119786 84934
rect 120022 84698 155786 84934
rect 156022 84698 191786 84934
rect 192022 84698 227786 84934
rect 228022 84698 263786 84934
rect 264022 84698 299786 84934
rect 300022 84698 314250 84934
rect 314486 84698 551786 84934
rect 552022 84698 591142 84934
rect 591378 84698 592500 84934
rect -8576 84676 592500 84698
rect -7636 84674 -7036 84676
rect 11604 84674 12204 84676
rect 47604 84674 48204 84676
rect 83604 84674 84204 84676
rect 119604 84674 120204 84676
rect 155604 84674 156204 84676
rect 191604 84674 192204 84676
rect 227604 84674 228204 84676
rect 263604 84674 264204 84676
rect 299604 84674 300204 84676
rect 314208 84674 314528 84676
rect 551604 84674 552204 84676
rect 590960 84674 591560 84676
rect -5756 81676 -5156 81678
rect 8004 81676 8604 81678
rect 44004 81676 44604 81678
rect 80004 81676 80604 81678
rect 116004 81676 116604 81678
rect 152004 81676 152604 81678
rect 188004 81676 188604 81678
rect 224004 81676 224604 81678
rect 260004 81676 260604 81678
rect 296004 81676 296604 81678
rect 548004 81676 548604 81678
rect 589080 81676 589680 81678
rect -6696 81654 590620 81676
rect -6696 81418 -5574 81654
rect -5338 81418 8186 81654
rect 8422 81418 44186 81654
rect 44422 81418 80186 81654
rect 80422 81418 116186 81654
rect 116422 81418 152186 81654
rect 152422 81418 188186 81654
rect 188422 81418 224186 81654
rect 224422 81418 260186 81654
rect 260422 81418 296186 81654
rect 296422 81418 548186 81654
rect 548422 81418 589262 81654
rect 589498 81418 590620 81654
rect -6696 81334 590620 81418
rect -6696 81098 -5574 81334
rect -5338 81098 8186 81334
rect 8422 81098 44186 81334
rect 44422 81098 80186 81334
rect 80422 81098 116186 81334
rect 116422 81098 152186 81334
rect 152422 81098 188186 81334
rect 188422 81098 224186 81334
rect 224422 81098 260186 81334
rect 260422 81098 296186 81334
rect 296422 81098 548186 81334
rect 548422 81098 589262 81334
rect 589498 81098 590620 81334
rect -6696 81076 590620 81098
rect -5756 81074 -5156 81076
rect 8004 81074 8604 81076
rect 44004 81074 44604 81076
rect 80004 81074 80604 81076
rect 116004 81074 116604 81076
rect 152004 81074 152604 81076
rect 188004 81074 188604 81076
rect 224004 81074 224604 81076
rect 260004 81074 260604 81076
rect 296004 81074 296604 81076
rect 548004 81074 548604 81076
rect 589080 81074 589680 81076
rect -3876 78076 -3276 78078
rect 4404 78076 5004 78078
rect 40404 78076 41004 78078
rect 76404 78076 77004 78078
rect 112404 78076 113004 78078
rect 148404 78076 149004 78078
rect 184404 78076 185004 78078
rect 220404 78076 221004 78078
rect 256404 78076 257004 78078
rect 292404 78076 293004 78078
rect 544404 78076 545004 78078
rect 580404 78076 581004 78078
rect 587200 78076 587800 78078
rect -4816 78054 588740 78076
rect -4816 77818 -3694 78054
rect -3458 77818 4586 78054
rect 4822 77818 40586 78054
rect 40822 77818 76586 78054
rect 76822 77818 112586 78054
rect 112822 77818 148586 78054
rect 148822 77818 184586 78054
rect 184822 77818 220586 78054
rect 220822 77818 256586 78054
rect 256822 77818 292586 78054
rect 292822 77818 544586 78054
rect 544822 77818 580586 78054
rect 580822 77818 587382 78054
rect 587618 77818 588740 78054
rect -4816 77734 588740 77818
rect -4816 77498 -3694 77734
rect -3458 77498 4586 77734
rect 4822 77498 40586 77734
rect 40822 77498 76586 77734
rect 76822 77498 112586 77734
rect 112822 77498 148586 77734
rect 148822 77498 184586 77734
rect 184822 77498 220586 77734
rect 220822 77498 256586 77734
rect 256822 77498 292586 77734
rect 292822 77498 544586 77734
rect 544822 77498 580586 77734
rect 580822 77498 587382 77734
rect 587618 77498 588740 77734
rect -4816 77476 588740 77498
rect -3876 77474 -3276 77476
rect 4404 77474 5004 77476
rect 40404 77474 41004 77476
rect 76404 77474 77004 77476
rect 112404 77474 113004 77476
rect 148404 77474 149004 77476
rect 184404 77474 185004 77476
rect 220404 77474 221004 77476
rect 256404 77474 257004 77476
rect 292404 77474 293004 77476
rect 544404 77474 545004 77476
rect 580404 77474 581004 77476
rect 587200 77474 587800 77476
rect -1996 74476 -1396 74478
rect 804 74476 1404 74478
rect 36804 74476 37404 74478
rect 72804 74476 73404 74478
rect 108804 74476 109404 74478
rect 144804 74476 145404 74478
rect 180804 74476 181404 74478
rect 216804 74476 217404 74478
rect 252804 74476 253404 74478
rect 288804 74476 289404 74478
rect 324804 74476 325404 74478
rect 360804 74476 361404 74478
rect 396804 74476 397404 74478
rect 432804 74476 433404 74478
rect 468804 74476 469404 74478
rect 504804 74476 505404 74478
rect 540804 74476 541404 74478
rect 576804 74476 577404 74478
rect 585320 74476 585920 74478
rect -2936 74454 586860 74476
rect -2936 74218 -1814 74454
rect -1578 74218 986 74454
rect 1222 74218 36986 74454
rect 37222 74218 72986 74454
rect 73222 74218 108986 74454
rect 109222 74218 144986 74454
rect 145222 74218 180986 74454
rect 181222 74218 216986 74454
rect 217222 74218 252986 74454
rect 253222 74218 288986 74454
rect 289222 74218 324986 74454
rect 325222 74218 360986 74454
rect 361222 74218 396986 74454
rect 397222 74218 432986 74454
rect 433222 74218 468986 74454
rect 469222 74218 504986 74454
rect 505222 74218 540986 74454
rect 541222 74218 576986 74454
rect 577222 74218 585502 74454
rect 585738 74218 586860 74454
rect -2936 74134 586860 74218
rect -2936 73898 -1814 74134
rect -1578 73898 986 74134
rect 1222 73898 36986 74134
rect 37222 73898 72986 74134
rect 73222 73898 108986 74134
rect 109222 73898 144986 74134
rect 145222 73898 180986 74134
rect 181222 73898 216986 74134
rect 217222 73898 252986 74134
rect 253222 73898 288986 74134
rect 289222 73898 324986 74134
rect 325222 73898 360986 74134
rect 361222 73898 396986 74134
rect 397222 73898 432986 74134
rect 433222 73898 468986 74134
rect 469222 73898 504986 74134
rect 505222 73898 540986 74134
rect 541222 73898 576986 74134
rect 577222 73898 585502 74134
rect 585738 73898 586860 74134
rect -2936 73876 586860 73898
rect -1996 73874 -1396 73876
rect 804 73874 1404 73876
rect 36804 73874 37404 73876
rect 72804 73874 73404 73876
rect 108804 73874 109404 73876
rect 144804 73874 145404 73876
rect 180804 73874 181404 73876
rect 216804 73874 217404 73876
rect 252804 73874 253404 73876
rect 288804 73874 289404 73876
rect 324804 73874 325404 73876
rect 360804 73874 361404 73876
rect 396804 73874 397404 73876
rect 432804 73874 433404 73876
rect 468804 73874 469404 73876
rect 504804 73874 505404 73876
rect 540804 73874 541404 73876
rect 576804 73874 577404 73876
rect 585320 73874 585920 73876
rect -8576 67276 -7976 67278
rect 29604 67276 30204 67278
rect 65604 67276 66204 67278
rect 101604 67276 102204 67278
rect 137604 67276 138204 67278
rect 173604 67276 174204 67278
rect 209604 67276 210204 67278
rect 245604 67276 246204 67278
rect 281604 67276 282204 67278
rect 317604 67276 318204 67278
rect 353604 67276 354204 67278
rect 389604 67276 390204 67278
rect 425604 67276 426204 67278
rect 461604 67276 462204 67278
rect 497604 67276 498204 67278
rect 533604 67276 534204 67278
rect 569604 67276 570204 67278
rect 591900 67276 592500 67278
rect -8576 67254 592500 67276
rect -8576 67018 -8394 67254
rect -8158 67018 29786 67254
rect 30022 67018 65786 67254
rect 66022 67018 101786 67254
rect 102022 67018 137786 67254
rect 138022 67018 173786 67254
rect 174022 67018 209786 67254
rect 210022 67018 245786 67254
rect 246022 67018 281786 67254
rect 282022 67018 317786 67254
rect 318022 67018 353786 67254
rect 354022 67018 389786 67254
rect 390022 67018 425786 67254
rect 426022 67018 461786 67254
rect 462022 67018 497786 67254
rect 498022 67018 533786 67254
rect 534022 67018 569786 67254
rect 570022 67018 592082 67254
rect 592318 67018 592500 67254
rect -8576 66934 592500 67018
rect -8576 66698 -8394 66934
rect -8158 66698 29786 66934
rect 30022 66698 65786 66934
rect 66022 66698 101786 66934
rect 102022 66698 137786 66934
rect 138022 66698 173786 66934
rect 174022 66698 209786 66934
rect 210022 66698 245786 66934
rect 246022 66698 281786 66934
rect 282022 66698 317786 66934
rect 318022 66698 353786 66934
rect 354022 66698 389786 66934
rect 390022 66698 425786 66934
rect 426022 66698 461786 66934
rect 462022 66698 497786 66934
rect 498022 66698 533786 66934
rect 534022 66698 569786 66934
rect 570022 66698 592082 66934
rect 592318 66698 592500 66934
rect -8576 66676 592500 66698
rect -8576 66674 -7976 66676
rect 29604 66674 30204 66676
rect 65604 66674 66204 66676
rect 101604 66674 102204 66676
rect 137604 66674 138204 66676
rect 173604 66674 174204 66676
rect 209604 66674 210204 66676
rect 245604 66674 246204 66676
rect 281604 66674 282204 66676
rect 317604 66674 318204 66676
rect 353604 66674 354204 66676
rect 389604 66674 390204 66676
rect 425604 66674 426204 66676
rect 461604 66674 462204 66676
rect 497604 66674 498204 66676
rect 533604 66674 534204 66676
rect 569604 66674 570204 66676
rect 591900 66674 592500 66676
rect -6696 63676 -6096 63678
rect 26004 63676 26604 63678
rect 62004 63676 62604 63678
rect 98004 63676 98604 63678
rect 134004 63676 134604 63678
rect 170004 63676 170604 63678
rect 206004 63676 206604 63678
rect 242004 63676 242604 63678
rect 278004 63676 278604 63678
rect 314004 63676 314604 63678
rect 350004 63676 350604 63678
rect 386004 63676 386604 63678
rect 422004 63676 422604 63678
rect 458004 63676 458604 63678
rect 494004 63676 494604 63678
rect 530004 63676 530604 63678
rect 566004 63676 566604 63678
rect 590020 63676 590620 63678
rect -6696 63654 590620 63676
rect -6696 63418 -6514 63654
rect -6278 63418 26186 63654
rect 26422 63418 62186 63654
rect 62422 63418 98186 63654
rect 98422 63418 134186 63654
rect 134422 63418 170186 63654
rect 170422 63418 206186 63654
rect 206422 63418 242186 63654
rect 242422 63418 278186 63654
rect 278422 63418 314186 63654
rect 314422 63418 350186 63654
rect 350422 63418 386186 63654
rect 386422 63418 422186 63654
rect 422422 63418 458186 63654
rect 458422 63418 494186 63654
rect 494422 63418 530186 63654
rect 530422 63418 566186 63654
rect 566422 63418 590202 63654
rect 590438 63418 590620 63654
rect -6696 63334 590620 63418
rect -6696 63098 -6514 63334
rect -6278 63098 26186 63334
rect 26422 63098 62186 63334
rect 62422 63098 98186 63334
rect 98422 63098 134186 63334
rect 134422 63098 170186 63334
rect 170422 63098 206186 63334
rect 206422 63098 242186 63334
rect 242422 63098 278186 63334
rect 278422 63098 314186 63334
rect 314422 63098 350186 63334
rect 350422 63098 386186 63334
rect 386422 63098 422186 63334
rect 422422 63098 458186 63334
rect 458422 63098 494186 63334
rect 494422 63098 530186 63334
rect 530422 63098 566186 63334
rect 566422 63098 590202 63334
rect 590438 63098 590620 63334
rect -6696 63076 590620 63098
rect -6696 63074 -6096 63076
rect 26004 63074 26604 63076
rect 62004 63074 62604 63076
rect 98004 63074 98604 63076
rect 134004 63074 134604 63076
rect 170004 63074 170604 63076
rect 206004 63074 206604 63076
rect 242004 63074 242604 63076
rect 278004 63074 278604 63076
rect 314004 63074 314604 63076
rect 350004 63074 350604 63076
rect 386004 63074 386604 63076
rect 422004 63074 422604 63076
rect 458004 63074 458604 63076
rect 494004 63074 494604 63076
rect 530004 63074 530604 63076
rect 566004 63074 566604 63076
rect 590020 63074 590620 63076
rect -4816 60076 -4216 60078
rect 22404 60076 23004 60078
rect 58404 60076 59004 60078
rect 94404 60076 95004 60078
rect 130404 60076 131004 60078
rect 166404 60076 167004 60078
rect 202404 60076 203004 60078
rect 238404 60076 239004 60078
rect 274404 60076 275004 60078
rect 310404 60076 311004 60078
rect 346404 60076 347004 60078
rect 382404 60076 383004 60078
rect 418404 60076 419004 60078
rect 454404 60076 455004 60078
rect 490404 60076 491004 60078
rect 526404 60076 527004 60078
rect 562404 60076 563004 60078
rect 588140 60076 588740 60078
rect -4816 60054 588740 60076
rect -4816 59818 -4634 60054
rect -4398 59818 22586 60054
rect 22822 59818 58586 60054
rect 58822 59818 94586 60054
rect 94822 59818 130586 60054
rect 130822 59818 166586 60054
rect 166822 59818 202586 60054
rect 202822 59818 238586 60054
rect 238822 59818 274586 60054
rect 274822 59818 310586 60054
rect 310822 59818 346586 60054
rect 346822 59818 382586 60054
rect 382822 59818 418586 60054
rect 418822 59818 454586 60054
rect 454822 59818 490586 60054
rect 490822 59818 526586 60054
rect 526822 59818 562586 60054
rect 562822 59818 588322 60054
rect 588558 59818 588740 60054
rect -4816 59734 588740 59818
rect -4816 59498 -4634 59734
rect -4398 59498 22586 59734
rect 22822 59498 58586 59734
rect 58822 59498 94586 59734
rect 94822 59498 130586 59734
rect 130822 59498 166586 59734
rect 166822 59498 202586 59734
rect 202822 59498 238586 59734
rect 238822 59498 274586 59734
rect 274822 59498 310586 59734
rect 310822 59498 346586 59734
rect 346822 59498 382586 59734
rect 382822 59498 418586 59734
rect 418822 59498 454586 59734
rect 454822 59498 490586 59734
rect 490822 59498 526586 59734
rect 526822 59498 562586 59734
rect 562822 59498 588322 59734
rect 588558 59498 588740 59734
rect -4816 59476 588740 59498
rect -4816 59474 -4216 59476
rect 22404 59474 23004 59476
rect 58404 59474 59004 59476
rect 94404 59474 95004 59476
rect 130404 59474 131004 59476
rect 166404 59474 167004 59476
rect 202404 59474 203004 59476
rect 238404 59474 239004 59476
rect 274404 59474 275004 59476
rect 310404 59474 311004 59476
rect 346404 59474 347004 59476
rect 382404 59474 383004 59476
rect 418404 59474 419004 59476
rect 454404 59474 455004 59476
rect 490404 59474 491004 59476
rect 526404 59474 527004 59476
rect 562404 59474 563004 59476
rect 588140 59474 588740 59476
rect -2936 56476 -2336 56478
rect 18804 56476 19404 56478
rect 54804 56476 55404 56478
rect 90804 56476 91404 56478
rect 126804 56476 127404 56478
rect 162804 56476 163404 56478
rect 198804 56476 199404 56478
rect 234804 56476 235404 56478
rect 270804 56476 271404 56478
rect 306804 56476 307404 56478
rect 342804 56476 343404 56478
rect 378804 56476 379404 56478
rect 414804 56476 415404 56478
rect 450804 56476 451404 56478
rect 486804 56476 487404 56478
rect 522804 56476 523404 56478
rect 558804 56476 559404 56478
rect 586260 56476 586860 56478
rect -2936 56454 586860 56476
rect -2936 56218 -2754 56454
rect -2518 56218 18986 56454
rect 19222 56218 54986 56454
rect 55222 56218 90986 56454
rect 91222 56218 126986 56454
rect 127222 56218 162986 56454
rect 163222 56218 198986 56454
rect 199222 56218 234986 56454
rect 235222 56218 270986 56454
rect 271222 56218 306986 56454
rect 307222 56218 342986 56454
rect 343222 56218 378986 56454
rect 379222 56218 414986 56454
rect 415222 56218 450986 56454
rect 451222 56218 486986 56454
rect 487222 56218 522986 56454
rect 523222 56218 558986 56454
rect 559222 56218 586442 56454
rect 586678 56218 586860 56454
rect -2936 56134 586860 56218
rect -2936 55898 -2754 56134
rect -2518 55898 18986 56134
rect 19222 55898 54986 56134
rect 55222 55898 90986 56134
rect 91222 55898 126986 56134
rect 127222 55898 162986 56134
rect 163222 55898 198986 56134
rect 199222 55898 234986 56134
rect 235222 55898 270986 56134
rect 271222 55898 306986 56134
rect 307222 55898 342986 56134
rect 343222 55898 378986 56134
rect 379222 55898 414986 56134
rect 415222 55898 450986 56134
rect 451222 55898 486986 56134
rect 487222 55898 522986 56134
rect 523222 55898 558986 56134
rect 559222 55898 586442 56134
rect 586678 55898 586860 56134
rect -2936 55876 586860 55898
rect -2936 55874 -2336 55876
rect 18804 55874 19404 55876
rect 54804 55874 55404 55876
rect 90804 55874 91404 55876
rect 126804 55874 127404 55876
rect 162804 55874 163404 55876
rect 198804 55874 199404 55876
rect 234804 55874 235404 55876
rect 270804 55874 271404 55876
rect 306804 55874 307404 55876
rect 342804 55874 343404 55876
rect 378804 55874 379404 55876
rect 414804 55874 415404 55876
rect 450804 55874 451404 55876
rect 486804 55874 487404 55876
rect 522804 55874 523404 55876
rect 558804 55874 559404 55876
rect 586260 55874 586860 55876
rect -7636 49276 -7036 49278
rect 11604 49276 12204 49278
rect 47604 49276 48204 49278
rect 83604 49276 84204 49278
rect 119604 49276 120204 49278
rect 155604 49276 156204 49278
rect 191604 49276 192204 49278
rect 227604 49276 228204 49278
rect 263604 49276 264204 49278
rect 299604 49276 300204 49278
rect 335604 49276 336204 49278
rect 371604 49276 372204 49278
rect 407604 49276 408204 49278
rect 443604 49276 444204 49278
rect 479604 49276 480204 49278
rect 515604 49276 516204 49278
rect 551604 49276 552204 49278
rect 590960 49276 591560 49278
rect -8576 49254 592500 49276
rect -8576 49018 -7454 49254
rect -7218 49018 11786 49254
rect 12022 49018 47786 49254
rect 48022 49018 83786 49254
rect 84022 49018 119786 49254
rect 120022 49018 155786 49254
rect 156022 49018 191786 49254
rect 192022 49018 227786 49254
rect 228022 49018 263786 49254
rect 264022 49018 299786 49254
rect 300022 49018 335786 49254
rect 336022 49018 371786 49254
rect 372022 49018 407786 49254
rect 408022 49018 443786 49254
rect 444022 49018 479786 49254
rect 480022 49018 515786 49254
rect 516022 49018 551786 49254
rect 552022 49018 591142 49254
rect 591378 49018 592500 49254
rect -8576 48934 592500 49018
rect -8576 48698 -7454 48934
rect -7218 48698 11786 48934
rect 12022 48698 47786 48934
rect 48022 48698 83786 48934
rect 84022 48698 119786 48934
rect 120022 48698 155786 48934
rect 156022 48698 191786 48934
rect 192022 48698 227786 48934
rect 228022 48698 263786 48934
rect 264022 48698 299786 48934
rect 300022 48698 335786 48934
rect 336022 48698 371786 48934
rect 372022 48698 407786 48934
rect 408022 48698 443786 48934
rect 444022 48698 479786 48934
rect 480022 48698 515786 48934
rect 516022 48698 551786 48934
rect 552022 48698 591142 48934
rect 591378 48698 592500 48934
rect -8576 48676 592500 48698
rect -7636 48674 -7036 48676
rect 11604 48674 12204 48676
rect 47604 48674 48204 48676
rect 83604 48674 84204 48676
rect 119604 48674 120204 48676
rect 155604 48674 156204 48676
rect 191604 48674 192204 48676
rect 227604 48674 228204 48676
rect 263604 48674 264204 48676
rect 299604 48674 300204 48676
rect 335604 48674 336204 48676
rect 371604 48674 372204 48676
rect 407604 48674 408204 48676
rect 443604 48674 444204 48676
rect 479604 48674 480204 48676
rect 515604 48674 516204 48676
rect 551604 48674 552204 48676
rect 590960 48674 591560 48676
rect -5756 45676 -5156 45678
rect 8004 45676 8604 45678
rect 44004 45676 44604 45678
rect 80004 45676 80604 45678
rect 116004 45676 116604 45678
rect 152004 45676 152604 45678
rect 188004 45676 188604 45678
rect 224004 45676 224604 45678
rect 260004 45676 260604 45678
rect 296004 45676 296604 45678
rect 332004 45676 332604 45678
rect 368004 45676 368604 45678
rect 404004 45676 404604 45678
rect 440004 45676 440604 45678
rect 476004 45676 476604 45678
rect 512004 45676 512604 45678
rect 548004 45676 548604 45678
rect 589080 45676 589680 45678
rect -6696 45654 590620 45676
rect -6696 45418 -5574 45654
rect -5338 45418 8186 45654
rect 8422 45418 44186 45654
rect 44422 45418 80186 45654
rect 80422 45418 116186 45654
rect 116422 45418 152186 45654
rect 152422 45418 188186 45654
rect 188422 45418 224186 45654
rect 224422 45418 260186 45654
rect 260422 45418 296186 45654
rect 296422 45418 332186 45654
rect 332422 45418 368186 45654
rect 368422 45418 404186 45654
rect 404422 45418 440186 45654
rect 440422 45418 476186 45654
rect 476422 45418 512186 45654
rect 512422 45418 548186 45654
rect 548422 45418 589262 45654
rect 589498 45418 590620 45654
rect -6696 45334 590620 45418
rect -6696 45098 -5574 45334
rect -5338 45098 8186 45334
rect 8422 45098 44186 45334
rect 44422 45098 80186 45334
rect 80422 45098 116186 45334
rect 116422 45098 152186 45334
rect 152422 45098 188186 45334
rect 188422 45098 224186 45334
rect 224422 45098 260186 45334
rect 260422 45098 296186 45334
rect 296422 45098 332186 45334
rect 332422 45098 368186 45334
rect 368422 45098 404186 45334
rect 404422 45098 440186 45334
rect 440422 45098 476186 45334
rect 476422 45098 512186 45334
rect 512422 45098 548186 45334
rect 548422 45098 589262 45334
rect 589498 45098 590620 45334
rect -6696 45076 590620 45098
rect -5756 45074 -5156 45076
rect 8004 45074 8604 45076
rect 44004 45074 44604 45076
rect 80004 45074 80604 45076
rect 116004 45074 116604 45076
rect 152004 45074 152604 45076
rect 188004 45074 188604 45076
rect 224004 45074 224604 45076
rect 260004 45074 260604 45076
rect 296004 45074 296604 45076
rect 332004 45074 332604 45076
rect 368004 45074 368604 45076
rect 404004 45074 404604 45076
rect 440004 45074 440604 45076
rect 476004 45074 476604 45076
rect 512004 45074 512604 45076
rect 548004 45074 548604 45076
rect 589080 45074 589680 45076
rect -3876 42076 -3276 42078
rect 4404 42076 5004 42078
rect 40404 42076 41004 42078
rect 76404 42076 77004 42078
rect 112404 42076 113004 42078
rect 148404 42076 149004 42078
rect 184404 42076 185004 42078
rect 220404 42076 221004 42078
rect 256404 42076 257004 42078
rect 292404 42076 293004 42078
rect 328404 42076 329004 42078
rect 364404 42076 365004 42078
rect 400404 42076 401004 42078
rect 436404 42076 437004 42078
rect 472404 42076 473004 42078
rect 508404 42076 509004 42078
rect 544404 42076 545004 42078
rect 580404 42076 581004 42078
rect 587200 42076 587800 42078
rect -4816 42054 588740 42076
rect -4816 41818 -3694 42054
rect -3458 41818 4586 42054
rect 4822 41818 40586 42054
rect 40822 41818 76586 42054
rect 76822 41818 112586 42054
rect 112822 41818 148586 42054
rect 148822 41818 184586 42054
rect 184822 41818 220586 42054
rect 220822 41818 256586 42054
rect 256822 41818 292586 42054
rect 292822 41818 328586 42054
rect 328822 41818 364586 42054
rect 364822 41818 400586 42054
rect 400822 41818 436586 42054
rect 436822 41818 472586 42054
rect 472822 41818 508586 42054
rect 508822 41818 544586 42054
rect 544822 41818 580586 42054
rect 580822 41818 587382 42054
rect 587618 41818 588740 42054
rect -4816 41734 588740 41818
rect -4816 41498 -3694 41734
rect -3458 41498 4586 41734
rect 4822 41498 40586 41734
rect 40822 41498 76586 41734
rect 76822 41498 112586 41734
rect 112822 41498 148586 41734
rect 148822 41498 184586 41734
rect 184822 41498 220586 41734
rect 220822 41498 256586 41734
rect 256822 41498 292586 41734
rect 292822 41498 328586 41734
rect 328822 41498 364586 41734
rect 364822 41498 400586 41734
rect 400822 41498 436586 41734
rect 436822 41498 472586 41734
rect 472822 41498 508586 41734
rect 508822 41498 544586 41734
rect 544822 41498 580586 41734
rect 580822 41498 587382 41734
rect 587618 41498 588740 41734
rect -4816 41476 588740 41498
rect -3876 41474 -3276 41476
rect 4404 41474 5004 41476
rect 40404 41474 41004 41476
rect 76404 41474 77004 41476
rect 112404 41474 113004 41476
rect 148404 41474 149004 41476
rect 184404 41474 185004 41476
rect 220404 41474 221004 41476
rect 256404 41474 257004 41476
rect 292404 41474 293004 41476
rect 328404 41474 329004 41476
rect 364404 41474 365004 41476
rect 400404 41474 401004 41476
rect 436404 41474 437004 41476
rect 472404 41474 473004 41476
rect 508404 41474 509004 41476
rect 544404 41474 545004 41476
rect 580404 41474 581004 41476
rect 587200 41474 587800 41476
rect -1996 38476 -1396 38478
rect 804 38476 1404 38478
rect 36804 38476 37404 38478
rect 72804 38476 73404 38478
rect 108804 38476 109404 38478
rect 144804 38476 145404 38478
rect 180804 38476 181404 38478
rect 216804 38476 217404 38478
rect 252804 38476 253404 38478
rect 288804 38476 289404 38478
rect 324804 38476 325404 38478
rect 360804 38476 361404 38478
rect 396804 38476 397404 38478
rect 432804 38476 433404 38478
rect 468804 38476 469404 38478
rect 504804 38476 505404 38478
rect 540804 38476 541404 38478
rect 576804 38476 577404 38478
rect 585320 38476 585920 38478
rect -2936 38454 586860 38476
rect -2936 38218 -1814 38454
rect -1578 38218 986 38454
rect 1222 38218 36986 38454
rect 37222 38218 72986 38454
rect 73222 38218 108986 38454
rect 109222 38218 144986 38454
rect 145222 38218 180986 38454
rect 181222 38218 216986 38454
rect 217222 38218 252986 38454
rect 253222 38218 288986 38454
rect 289222 38218 324986 38454
rect 325222 38218 360986 38454
rect 361222 38218 396986 38454
rect 397222 38218 432986 38454
rect 433222 38218 468986 38454
rect 469222 38218 504986 38454
rect 505222 38218 540986 38454
rect 541222 38218 576986 38454
rect 577222 38218 585502 38454
rect 585738 38218 586860 38454
rect -2936 38134 586860 38218
rect -2936 37898 -1814 38134
rect -1578 37898 986 38134
rect 1222 37898 36986 38134
rect 37222 37898 72986 38134
rect 73222 37898 108986 38134
rect 109222 37898 144986 38134
rect 145222 37898 180986 38134
rect 181222 37898 216986 38134
rect 217222 37898 252986 38134
rect 253222 37898 288986 38134
rect 289222 37898 324986 38134
rect 325222 37898 360986 38134
rect 361222 37898 396986 38134
rect 397222 37898 432986 38134
rect 433222 37898 468986 38134
rect 469222 37898 504986 38134
rect 505222 37898 540986 38134
rect 541222 37898 576986 38134
rect 577222 37898 585502 38134
rect 585738 37898 586860 38134
rect -2936 37876 586860 37898
rect -1996 37874 -1396 37876
rect 804 37874 1404 37876
rect 36804 37874 37404 37876
rect 72804 37874 73404 37876
rect 108804 37874 109404 37876
rect 144804 37874 145404 37876
rect 180804 37874 181404 37876
rect 216804 37874 217404 37876
rect 252804 37874 253404 37876
rect 288804 37874 289404 37876
rect 324804 37874 325404 37876
rect 360804 37874 361404 37876
rect 396804 37874 397404 37876
rect 432804 37874 433404 37876
rect 468804 37874 469404 37876
rect 504804 37874 505404 37876
rect 540804 37874 541404 37876
rect 576804 37874 577404 37876
rect 585320 37874 585920 37876
rect -8576 31276 -7976 31278
rect 29604 31276 30204 31278
rect 65604 31276 66204 31278
rect 101604 31276 102204 31278
rect 137604 31276 138204 31278
rect 173604 31276 174204 31278
rect 209604 31276 210204 31278
rect 245604 31276 246204 31278
rect 281604 31276 282204 31278
rect 317604 31276 318204 31278
rect 353604 31276 354204 31278
rect 389604 31276 390204 31278
rect 425604 31276 426204 31278
rect 461604 31276 462204 31278
rect 497604 31276 498204 31278
rect 533604 31276 534204 31278
rect 569604 31276 570204 31278
rect 591900 31276 592500 31278
rect -8576 31254 592500 31276
rect -8576 31018 -8394 31254
rect -8158 31018 29786 31254
rect 30022 31018 65786 31254
rect 66022 31018 101786 31254
rect 102022 31018 137786 31254
rect 138022 31018 173786 31254
rect 174022 31018 209786 31254
rect 210022 31018 245786 31254
rect 246022 31018 281786 31254
rect 282022 31018 317786 31254
rect 318022 31018 353786 31254
rect 354022 31018 389786 31254
rect 390022 31018 425786 31254
rect 426022 31018 461786 31254
rect 462022 31018 497786 31254
rect 498022 31018 533786 31254
rect 534022 31018 569786 31254
rect 570022 31018 592082 31254
rect 592318 31018 592500 31254
rect -8576 30934 592500 31018
rect -8576 30698 -8394 30934
rect -8158 30698 29786 30934
rect 30022 30698 65786 30934
rect 66022 30698 101786 30934
rect 102022 30698 137786 30934
rect 138022 30698 173786 30934
rect 174022 30698 209786 30934
rect 210022 30698 245786 30934
rect 246022 30698 281786 30934
rect 282022 30698 317786 30934
rect 318022 30698 353786 30934
rect 354022 30698 389786 30934
rect 390022 30698 425786 30934
rect 426022 30698 461786 30934
rect 462022 30698 497786 30934
rect 498022 30698 533786 30934
rect 534022 30698 569786 30934
rect 570022 30698 592082 30934
rect 592318 30698 592500 30934
rect -8576 30676 592500 30698
rect -8576 30674 -7976 30676
rect 29604 30674 30204 30676
rect 65604 30674 66204 30676
rect 101604 30674 102204 30676
rect 137604 30674 138204 30676
rect 173604 30674 174204 30676
rect 209604 30674 210204 30676
rect 245604 30674 246204 30676
rect 281604 30674 282204 30676
rect 317604 30674 318204 30676
rect 353604 30674 354204 30676
rect 389604 30674 390204 30676
rect 425604 30674 426204 30676
rect 461604 30674 462204 30676
rect 497604 30674 498204 30676
rect 533604 30674 534204 30676
rect 569604 30674 570204 30676
rect 591900 30674 592500 30676
rect -6696 27676 -6096 27678
rect 26004 27676 26604 27678
rect 62004 27676 62604 27678
rect 98004 27676 98604 27678
rect 134004 27676 134604 27678
rect 170004 27676 170604 27678
rect 206004 27676 206604 27678
rect 242004 27676 242604 27678
rect 278004 27676 278604 27678
rect 314004 27676 314604 27678
rect 350004 27676 350604 27678
rect 386004 27676 386604 27678
rect 422004 27676 422604 27678
rect 458004 27676 458604 27678
rect 494004 27676 494604 27678
rect 530004 27676 530604 27678
rect 566004 27676 566604 27678
rect 590020 27676 590620 27678
rect -6696 27654 590620 27676
rect -6696 27418 -6514 27654
rect -6278 27418 26186 27654
rect 26422 27418 62186 27654
rect 62422 27418 98186 27654
rect 98422 27418 134186 27654
rect 134422 27418 170186 27654
rect 170422 27418 206186 27654
rect 206422 27418 242186 27654
rect 242422 27418 278186 27654
rect 278422 27418 314186 27654
rect 314422 27418 350186 27654
rect 350422 27418 386186 27654
rect 386422 27418 422186 27654
rect 422422 27418 458186 27654
rect 458422 27418 494186 27654
rect 494422 27418 530186 27654
rect 530422 27418 566186 27654
rect 566422 27418 590202 27654
rect 590438 27418 590620 27654
rect -6696 27334 590620 27418
rect -6696 27098 -6514 27334
rect -6278 27098 26186 27334
rect 26422 27098 62186 27334
rect 62422 27098 98186 27334
rect 98422 27098 134186 27334
rect 134422 27098 170186 27334
rect 170422 27098 206186 27334
rect 206422 27098 242186 27334
rect 242422 27098 278186 27334
rect 278422 27098 314186 27334
rect 314422 27098 350186 27334
rect 350422 27098 386186 27334
rect 386422 27098 422186 27334
rect 422422 27098 458186 27334
rect 458422 27098 494186 27334
rect 494422 27098 530186 27334
rect 530422 27098 566186 27334
rect 566422 27098 590202 27334
rect 590438 27098 590620 27334
rect -6696 27076 590620 27098
rect -6696 27074 -6096 27076
rect 26004 27074 26604 27076
rect 62004 27074 62604 27076
rect 98004 27074 98604 27076
rect 134004 27074 134604 27076
rect 170004 27074 170604 27076
rect 206004 27074 206604 27076
rect 242004 27074 242604 27076
rect 278004 27074 278604 27076
rect 314004 27074 314604 27076
rect 350004 27074 350604 27076
rect 386004 27074 386604 27076
rect 422004 27074 422604 27076
rect 458004 27074 458604 27076
rect 494004 27074 494604 27076
rect 530004 27074 530604 27076
rect 566004 27074 566604 27076
rect 590020 27074 590620 27076
rect -4816 24076 -4216 24078
rect 22404 24076 23004 24078
rect 58404 24076 59004 24078
rect 94404 24076 95004 24078
rect 130404 24076 131004 24078
rect 166404 24076 167004 24078
rect 202404 24076 203004 24078
rect 238404 24076 239004 24078
rect 274404 24076 275004 24078
rect 310404 24076 311004 24078
rect 346404 24076 347004 24078
rect 382404 24076 383004 24078
rect 418404 24076 419004 24078
rect 454404 24076 455004 24078
rect 490404 24076 491004 24078
rect 526404 24076 527004 24078
rect 562404 24076 563004 24078
rect 588140 24076 588740 24078
rect -4816 24054 588740 24076
rect -4816 23818 -4634 24054
rect -4398 23818 22586 24054
rect 22822 23818 58586 24054
rect 58822 23818 94586 24054
rect 94822 23818 130586 24054
rect 130822 23818 166586 24054
rect 166822 23818 202586 24054
rect 202822 23818 238586 24054
rect 238822 23818 274586 24054
rect 274822 23818 310586 24054
rect 310822 23818 346586 24054
rect 346822 23818 382586 24054
rect 382822 23818 418586 24054
rect 418822 23818 454586 24054
rect 454822 23818 490586 24054
rect 490822 23818 526586 24054
rect 526822 23818 562586 24054
rect 562822 23818 588322 24054
rect 588558 23818 588740 24054
rect -4816 23734 588740 23818
rect -4816 23498 -4634 23734
rect -4398 23498 22586 23734
rect 22822 23498 58586 23734
rect 58822 23498 94586 23734
rect 94822 23498 130586 23734
rect 130822 23498 166586 23734
rect 166822 23498 202586 23734
rect 202822 23498 238586 23734
rect 238822 23498 274586 23734
rect 274822 23498 310586 23734
rect 310822 23498 346586 23734
rect 346822 23498 382586 23734
rect 382822 23498 418586 23734
rect 418822 23498 454586 23734
rect 454822 23498 490586 23734
rect 490822 23498 526586 23734
rect 526822 23498 562586 23734
rect 562822 23498 588322 23734
rect 588558 23498 588740 23734
rect -4816 23476 588740 23498
rect -4816 23474 -4216 23476
rect 22404 23474 23004 23476
rect 58404 23474 59004 23476
rect 94404 23474 95004 23476
rect 130404 23474 131004 23476
rect 166404 23474 167004 23476
rect 202404 23474 203004 23476
rect 238404 23474 239004 23476
rect 274404 23474 275004 23476
rect 310404 23474 311004 23476
rect 346404 23474 347004 23476
rect 382404 23474 383004 23476
rect 418404 23474 419004 23476
rect 454404 23474 455004 23476
rect 490404 23474 491004 23476
rect 526404 23474 527004 23476
rect 562404 23474 563004 23476
rect 588140 23474 588740 23476
rect -2936 20476 -2336 20478
rect 18804 20476 19404 20478
rect 54804 20476 55404 20478
rect 90804 20476 91404 20478
rect 126804 20476 127404 20478
rect 162804 20476 163404 20478
rect 198804 20476 199404 20478
rect 234804 20476 235404 20478
rect 270804 20476 271404 20478
rect 306804 20476 307404 20478
rect 342804 20476 343404 20478
rect 378804 20476 379404 20478
rect 414804 20476 415404 20478
rect 450804 20476 451404 20478
rect 486804 20476 487404 20478
rect 522804 20476 523404 20478
rect 558804 20476 559404 20478
rect 586260 20476 586860 20478
rect -2936 20454 586860 20476
rect -2936 20218 -2754 20454
rect -2518 20218 18986 20454
rect 19222 20218 54986 20454
rect 55222 20218 90986 20454
rect 91222 20218 126986 20454
rect 127222 20218 162986 20454
rect 163222 20218 198986 20454
rect 199222 20218 234986 20454
rect 235222 20218 270986 20454
rect 271222 20218 306986 20454
rect 307222 20218 342986 20454
rect 343222 20218 378986 20454
rect 379222 20218 414986 20454
rect 415222 20218 450986 20454
rect 451222 20218 486986 20454
rect 487222 20218 522986 20454
rect 523222 20218 558986 20454
rect 559222 20218 586442 20454
rect 586678 20218 586860 20454
rect -2936 20134 586860 20218
rect -2936 19898 -2754 20134
rect -2518 19898 18986 20134
rect 19222 19898 54986 20134
rect 55222 19898 90986 20134
rect 91222 19898 126986 20134
rect 127222 19898 162986 20134
rect 163222 19898 198986 20134
rect 199222 19898 234986 20134
rect 235222 19898 270986 20134
rect 271222 19898 306986 20134
rect 307222 19898 342986 20134
rect 343222 19898 378986 20134
rect 379222 19898 414986 20134
rect 415222 19898 450986 20134
rect 451222 19898 486986 20134
rect 487222 19898 522986 20134
rect 523222 19898 558986 20134
rect 559222 19898 586442 20134
rect 586678 19898 586860 20134
rect -2936 19876 586860 19898
rect -2936 19874 -2336 19876
rect 18804 19874 19404 19876
rect 54804 19874 55404 19876
rect 90804 19874 91404 19876
rect 126804 19874 127404 19876
rect 162804 19874 163404 19876
rect 198804 19874 199404 19876
rect 234804 19874 235404 19876
rect 270804 19874 271404 19876
rect 306804 19874 307404 19876
rect 342804 19874 343404 19876
rect 378804 19874 379404 19876
rect 414804 19874 415404 19876
rect 450804 19874 451404 19876
rect 486804 19874 487404 19876
rect 522804 19874 523404 19876
rect 558804 19874 559404 19876
rect 586260 19874 586860 19876
rect -7636 13276 -7036 13278
rect 11604 13276 12204 13278
rect 47604 13276 48204 13278
rect 83604 13276 84204 13278
rect 119604 13276 120204 13278
rect 155604 13276 156204 13278
rect 191604 13276 192204 13278
rect 227604 13276 228204 13278
rect 263604 13276 264204 13278
rect 299604 13276 300204 13278
rect 335604 13276 336204 13278
rect 371604 13276 372204 13278
rect 407604 13276 408204 13278
rect 443604 13276 444204 13278
rect 479604 13276 480204 13278
rect 515604 13276 516204 13278
rect 551604 13276 552204 13278
rect 590960 13276 591560 13278
rect -8576 13254 592500 13276
rect -8576 13018 -7454 13254
rect -7218 13018 11786 13254
rect 12022 13018 47786 13254
rect 48022 13018 83786 13254
rect 84022 13018 119786 13254
rect 120022 13018 155786 13254
rect 156022 13018 191786 13254
rect 192022 13018 227786 13254
rect 228022 13018 263786 13254
rect 264022 13018 299786 13254
rect 300022 13018 335786 13254
rect 336022 13018 371786 13254
rect 372022 13018 407786 13254
rect 408022 13018 443786 13254
rect 444022 13018 479786 13254
rect 480022 13018 515786 13254
rect 516022 13018 551786 13254
rect 552022 13018 591142 13254
rect 591378 13018 592500 13254
rect -8576 12934 592500 13018
rect -8576 12698 -7454 12934
rect -7218 12698 11786 12934
rect 12022 12698 47786 12934
rect 48022 12698 83786 12934
rect 84022 12698 119786 12934
rect 120022 12698 155786 12934
rect 156022 12698 191786 12934
rect 192022 12698 227786 12934
rect 228022 12698 263786 12934
rect 264022 12698 299786 12934
rect 300022 12698 335786 12934
rect 336022 12698 371786 12934
rect 372022 12698 407786 12934
rect 408022 12698 443786 12934
rect 444022 12698 479786 12934
rect 480022 12698 515786 12934
rect 516022 12698 551786 12934
rect 552022 12698 591142 12934
rect 591378 12698 592500 12934
rect -8576 12676 592500 12698
rect -7636 12674 -7036 12676
rect 11604 12674 12204 12676
rect 47604 12674 48204 12676
rect 83604 12674 84204 12676
rect 119604 12674 120204 12676
rect 155604 12674 156204 12676
rect 191604 12674 192204 12676
rect 227604 12674 228204 12676
rect 263604 12674 264204 12676
rect 299604 12674 300204 12676
rect 335604 12674 336204 12676
rect 371604 12674 372204 12676
rect 407604 12674 408204 12676
rect 443604 12674 444204 12676
rect 479604 12674 480204 12676
rect 515604 12674 516204 12676
rect 551604 12674 552204 12676
rect 590960 12674 591560 12676
rect -5756 9676 -5156 9678
rect 8004 9676 8604 9678
rect 44004 9676 44604 9678
rect 80004 9676 80604 9678
rect 116004 9676 116604 9678
rect 152004 9676 152604 9678
rect 188004 9676 188604 9678
rect 224004 9676 224604 9678
rect 260004 9676 260604 9678
rect 296004 9676 296604 9678
rect 332004 9676 332604 9678
rect 368004 9676 368604 9678
rect 404004 9676 404604 9678
rect 440004 9676 440604 9678
rect 476004 9676 476604 9678
rect 512004 9676 512604 9678
rect 548004 9676 548604 9678
rect 589080 9676 589680 9678
rect -6696 9654 590620 9676
rect -6696 9418 -5574 9654
rect -5338 9418 8186 9654
rect 8422 9418 44186 9654
rect 44422 9418 80186 9654
rect 80422 9418 116186 9654
rect 116422 9418 152186 9654
rect 152422 9418 188186 9654
rect 188422 9418 224186 9654
rect 224422 9418 260186 9654
rect 260422 9418 296186 9654
rect 296422 9418 332186 9654
rect 332422 9418 368186 9654
rect 368422 9418 404186 9654
rect 404422 9418 440186 9654
rect 440422 9418 476186 9654
rect 476422 9418 512186 9654
rect 512422 9418 548186 9654
rect 548422 9418 589262 9654
rect 589498 9418 590620 9654
rect -6696 9334 590620 9418
rect -6696 9098 -5574 9334
rect -5338 9098 8186 9334
rect 8422 9098 44186 9334
rect 44422 9098 80186 9334
rect 80422 9098 116186 9334
rect 116422 9098 152186 9334
rect 152422 9098 188186 9334
rect 188422 9098 224186 9334
rect 224422 9098 260186 9334
rect 260422 9098 296186 9334
rect 296422 9098 332186 9334
rect 332422 9098 368186 9334
rect 368422 9098 404186 9334
rect 404422 9098 440186 9334
rect 440422 9098 476186 9334
rect 476422 9098 512186 9334
rect 512422 9098 548186 9334
rect 548422 9098 589262 9334
rect 589498 9098 590620 9334
rect -6696 9076 590620 9098
rect -5756 9074 -5156 9076
rect 8004 9074 8604 9076
rect 44004 9074 44604 9076
rect 80004 9074 80604 9076
rect 116004 9074 116604 9076
rect 152004 9074 152604 9076
rect 188004 9074 188604 9076
rect 224004 9074 224604 9076
rect 260004 9074 260604 9076
rect 296004 9074 296604 9076
rect 332004 9074 332604 9076
rect 368004 9074 368604 9076
rect 404004 9074 404604 9076
rect 440004 9074 440604 9076
rect 476004 9074 476604 9076
rect 512004 9074 512604 9076
rect 548004 9074 548604 9076
rect 589080 9074 589680 9076
rect -3876 6076 -3276 6078
rect 4404 6076 5004 6078
rect 40404 6076 41004 6078
rect 76404 6076 77004 6078
rect 112404 6076 113004 6078
rect 148404 6076 149004 6078
rect 184404 6076 185004 6078
rect 220404 6076 221004 6078
rect 256404 6076 257004 6078
rect 292404 6076 293004 6078
rect 328404 6076 329004 6078
rect 364404 6076 365004 6078
rect 400404 6076 401004 6078
rect 436404 6076 437004 6078
rect 472404 6076 473004 6078
rect 508404 6076 509004 6078
rect 544404 6076 545004 6078
rect 580404 6076 581004 6078
rect 587200 6076 587800 6078
rect -4816 6054 588740 6076
rect -4816 5818 -3694 6054
rect -3458 5818 4586 6054
rect 4822 5818 40586 6054
rect 40822 5818 76586 6054
rect 76822 5818 112586 6054
rect 112822 5818 148586 6054
rect 148822 5818 184586 6054
rect 184822 5818 220586 6054
rect 220822 5818 256586 6054
rect 256822 5818 292586 6054
rect 292822 5818 328586 6054
rect 328822 5818 364586 6054
rect 364822 5818 400586 6054
rect 400822 5818 436586 6054
rect 436822 5818 472586 6054
rect 472822 5818 508586 6054
rect 508822 5818 544586 6054
rect 544822 5818 580586 6054
rect 580822 5818 587382 6054
rect 587618 5818 588740 6054
rect -4816 5734 588740 5818
rect -4816 5498 -3694 5734
rect -3458 5498 4586 5734
rect 4822 5498 40586 5734
rect 40822 5498 76586 5734
rect 76822 5498 112586 5734
rect 112822 5498 148586 5734
rect 148822 5498 184586 5734
rect 184822 5498 220586 5734
rect 220822 5498 256586 5734
rect 256822 5498 292586 5734
rect 292822 5498 328586 5734
rect 328822 5498 364586 5734
rect 364822 5498 400586 5734
rect 400822 5498 436586 5734
rect 436822 5498 472586 5734
rect 472822 5498 508586 5734
rect 508822 5498 544586 5734
rect 544822 5498 580586 5734
rect 580822 5498 587382 5734
rect 587618 5498 588740 5734
rect -4816 5476 588740 5498
rect -3876 5474 -3276 5476
rect 4404 5474 5004 5476
rect 40404 5474 41004 5476
rect 76404 5474 77004 5476
rect 112404 5474 113004 5476
rect 148404 5474 149004 5476
rect 184404 5474 185004 5476
rect 220404 5474 221004 5476
rect 256404 5474 257004 5476
rect 292404 5474 293004 5476
rect 328404 5474 329004 5476
rect 364404 5474 365004 5476
rect 400404 5474 401004 5476
rect 436404 5474 437004 5476
rect 472404 5474 473004 5476
rect 508404 5474 509004 5476
rect 544404 5474 545004 5476
rect 580404 5474 581004 5476
rect 587200 5474 587800 5476
rect -1996 2476 -1396 2478
rect 804 2476 1404 2478
rect 36804 2476 37404 2478
rect 72804 2476 73404 2478
rect 108804 2476 109404 2478
rect 144804 2476 145404 2478
rect 180804 2476 181404 2478
rect 216804 2476 217404 2478
rect 252804 2476 253404 2478
rect 288804 2476 289404 2478
rect 324804 2476 325404 2478
rect 360804 2476 361404 2478
rect 396804 2476 397404 2478
rect 432804 2476 433404 2478
rect 468804 2476 469404 2478
rect 504804 2476 505404 2478
rect 540804 2476 541404 2478
rect 576804 2476 577404 2478
rect 585320 2476 585920 2478
rect -2936 2454 586860 2476
rect -2936 2218 -1814 2454
rect -1578 2218 986 2454
rect 1222 2218 36986 2454
rect 37222 2218 72986 2454
rect 73222 2218 108986 2454
rect 109222 2218 144986 2454
rect 145222 2218 180986 2454
rect 181222 2218 216986 2454
rect 217222 2218 252986 2454
rect 253222 2218 288986 2454
rect 289222 2218 324986 2454
rect 325222 2218 360986 2454
rect 361222 2218 396986 2454
rect 397222 2218 432986 2454
rect 433222 2218 468986 2454
rect 469222 2218 504986 2454
rect 505222 2218 540986 2454
rect 541222 2218 576986 2454
rect 577222 2218 585502 2454
rect 585738 2218 586860 2454
rect -2936 2134 586860 2218
rect -2936 1898 -1814 2134
rect -1578 1898 986 2134
rect 1222 1898 36986 2134
rect 37222 1898 72986 2134
rect 73222 1898 108986 2134
rect 109222 1898 144986 2134
rect 145222 1898 180986 2134
rect 181222 1898 216986 2134
rect 217222 1898 252986 2134
rect 253222 1898 288986 2134
rect 289222 1898 324986 2134
rect 325222 1898 360986 2134
rect 361222 1898 396986 2134
rect 397222 1898 432986 2134
rect 433222 1898 468986 2134
rect 469222 1898 504986 2134
rect 505222 1898 540986 2134
rect 541222 1898 576986 2134
rect 577222 1898 585502 2134
rect 585738 1898 586860 2134
rect -2936 1876 586860 1898
rect -1996 1874 -1396 1876
rect 804 1874 1404 1876
rect 36804 1874 37404 1876
rect 72804 1874 73404 1876
rect 108804 1874 109404 1876
rect 144804 1874 145404 1876
rect 180804 1874 181404 1876
rect 216804 1874 217404 1876
rect 252804 1874 253404 1876
rect 288804 1874 289404 1876
rect 324804 1874 325404 1876
rect 360804 1874 361404 1876
rect 396804 1874 397404 1876
rect 432804 1874 433404 1876
rect 468804 1874 469404 1876
rect 504804 1874 505404 1876
rect 540804 1874 541404 1876
rect 576804 1874 577404 1876
rect 585320 1874 585920 1876
rect -1996 -324 -1396 -322
rect 804 -324 1404 -322
rect 36804 -324 37404 -322
rect 72804 -324 73404 -322
rect 108804 -324 109404 -322
rect 144804 -324 145404 -322
rect 180804 -324 181404 -322
rect 216804 -324 217404 -322
rect 252804 -324 253404 -322
rect 288804 -324 289404 -322
rect 324804 -324 325404 -322
rect 360804 -324 361404 -322
rect 396804 -324 397404 -322
rect 432804 -324 433404 -322
rect 468804 -324 469404 -322
rect 504804 -324 505404 -322
rect 540804 -324 541404 -322
rect 576804 -324 577404 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 986 -346
rect 1222 -582 36986 -346
rect 37222 -582 72986 -346
rect 73222 -582 108986 -346
rect 109222 -582 144986 -346
rect 145222 -582 180986 -346
rect 181222 -582 216986 -346
rect 217222 -582 252986 -346
rect 253222 -582 288986 -346
rect 289222 -582 324986 -346
rect 325222 -582 360986 -346
rect 361222 -582 396986 -346
rect 397222 -582 432986 -346
rect 433222 -582 468986 -346
rect 469222 -582 504986 -346
rect 505222 -582 540986 -346
rect 541222 -582 576986 -346
rect 577222 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 986 -666
rect 1222 -902 36986 -666
rect 37222 -902 72986 -666
rect 73222 -902 108986 -666
rect 109222 -902 144986 -666
rect 145222 -902 180986 -666
rect 181222 -902 216986 -666
rect 217222 -902 252986 -666
rect 253222 -902 288986 -666
rect 289222 -902 324986 -666
rect 325222 -902 360986 -666
rect 361222 -902 396986 -666
rect 397222 -902 432986 -666
rect 433222 -902 468986 -666
rect 469222 -902 504986 -666
rect 505222 -902 540986 -666
rect 541222 -902 576986 -666
rect 577222 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 108804 -926 109404 -924
rect 144804 -926 145404 -924
rect 180804 -926 181404 -924
rect 216804 -926 217404 -924
rect 252804 -926 253404 -924
rect 288804 -926 289404 -924
rect 324804 -926 325404 -924
rect 360804 -926 361404 -924
rect 396804 -926 397404 -924
rect 432804 -926 433404 -924
rect 468804 -926 469404 -924
rect 504804 -926 505404 -924
rect 540804 -926 541404 -924
rect 576804 -926 577404 -924
rect 585320 -926 585920 -924
rect -2936 -1264 -2336 -1262
rect 18804 -1264 19404 -1262
rect 54804 -1264 55404 -1262
rect 90804 -1264 91404 -1262
rect 126804 -1264 127404 -1262
rect 162804 -1264 163404 -1262
rect 198804 -1264 199404 -1262
rect 234804 -1264 235404 -1262
rect 270804 -1264 271404 -1262
rect 306804 -1264 307404 -1262
rect 342804 -1264 343404 -1262
rect 378804 -1264 379404 -1262
rect 414804 -1264 415404 -1262
rect 450804 -1264 451404 -1262
rect 486804 -1264 487404 -1262
rect 522804 -1264 523404 -1262
rect 558804 -1264 559404 -1262
rect 586260 -1264 586860 -1262
rect -2936 -1286 586860 -1264
rect -2936 -1522 -2754 -1286
rect -2518 -1522 18986 -1286
rect 19222 -1522 54986 -1286
rect 55222 -1522 90986 -1286
rect 91222 -1522 126986 -1286
rect 127222 -1522 162986 -1286
rect 163222 -1522 198986 -1286
rect 199222 -1522 234986 -1286
rect 235222 -1522 270986 -1286
rect 271222 -1522 306986 -1286
rect 307222 -1522 342986 -1286
rect 343222 -1522 378986 -1286
rect 379222 -1522 414986 -1286
rect 415222 -1522 450986 -1286
rect 451222 -1522 486986 -1286
rect 487222 -1522 522986 -1286
rect 523222 -1522 558986 -1286
rect 559222 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect -2936 -1606 586860 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 18986 -1606
rect 19222 -1842 54986 -1606
rect 55222 -1842 90986 -1606
rect 91222 -1842 126986 -1606
rect 127222 -1842 162986 -1606
rect 163222 -1842 198986 -1606
rect 199222 -1842 234986 -1606
rect 235222 -1842 270986 -1606
rect 271222 -1842 306986 -1606
rect 307222 -1842 342986 -1606
rect 343222 -1842 378986 -1606
rect 379222 -1842 414986 -1606
rect 415222 -1842 450986 -1606
rect 451222 -1842 486986 -1606
rect 487222 -1842 522986 -1606
rect 523222 -1842 558986 -1606
rect 559222 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect -2936 -1864 586860 -1842
rect -2936 -1866 -2336 -1864
rect 18804 -1866 19404 -1864
rect 54804 -1866 55404 -1864
rect 90804 -1866 91404 -1864
rect 126804 -1866 127404 -1864
rect 162804 -1866 163404 -1864
rect 198804 -1866 199404 -1864
rect 234804 -1866 235404 -1864
rect 270804 -1866 271404 -1864
rect 306804 -1866 307404 -1864
rect 342804 -1866 343404 -1864
rect 378804 -1866 379404 -1864
rect 414804 -1866 415404 -1864
rect 450804 -1866 451404 -1864
rect 486804 -1866 487404 -1864
rect 522804 -1866 523404 -1864
rect 558804 -1866 559404 -1864
rect 586260 -1866 586860 -1864
rect -3876 -2204 -3276 -2202
rect 4404 -2204 5004 -2202
rect 40404 -2204 41004 -2202
rect 76404 -2204 77004 -2202
rect 112404 -2204 113004 -2202
rect 148404 -2204 149004 -2202
rect 184404 -2204 185004 -2202
rect 220404 -2204 221004 -2202
rect 256404 -2204 257004 -2202
rect 292404 -2204 293004 -2202
rect 328404 -2204 329004 -2202
rect 364404 -2204 365004 -2202
rect 400404 -2204 401004 -2202
rect 436404 -2204 437004 -2202
rect 472404 -2204 473004 -2202
rect 508404 -2204 509004 -2202
rect 544404 -2204 545004 -2202
rect 580404 -2204 581004 -2202
rect 587200 -2204 587800 -2202
rect -3876 -2226 587800 -2204
rect -3876 -2462 -3694 -2226
rect -3458 -2462 4586 -2226
rect 4822 -2462 40586 -2226
rect 40822 -2462 76586 -2226
rect 76822 -2462 112586 -2226
rect 112822 -2462 148586 -2226
rect 148822 -2462 184586 -2226
rect 184822 -2462 220586 -2226
rect 220822 -2462 256586 -2226
rect 256822 -2462 292586 -2226
rect 292822 -2462 328586 -2226
rect 328822 -2462 364586 -2226
rect 364822 -2462 400586 -2226
rect 400822 -2462 436586 -2226
rect 436822 -2462 472586 -2226
rect 472822 -2462 508586 -2226
rect 508822 -2462 544586 -2226
rect 544822 -2462 580586 -2226
rect 580822 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect -3876 -2546 587800 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 4586 -2546
rect 4822 -2782 40586 -2546
rect 40822 -2782 76586 -2546
rect 76822 -2782 112586 -2546
rect 112822 -2782 148586 -2546
rect 148822 -2782 184586 -2546
rect 184822 -2782 220586 -2546
rect 220822 -2782 256586 -2546
rect 256822 -2782 292586 -2546
rect 292822 -2782 328586 -2546
rect 328822 -2782 364586 -2546
rect 364822 -2782 400586 -2546
rect 400822 -2782 436586 -2546
rect 436822 -2782 472586 -2546
rect 472822 -2782 508586 -2546
rect 508822 -2782 544586 -2546
rect 544822 -2782 580586 -2546
rect 580822 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect -3876 -2804 587800 -2782
rect -3876 -2806 -3276 -2804
rect 4404 -2806 5004 -2804
rect 40404 -2806 41004 -2804
rect 76404 -2806 77004 -2804
rect 112404 -2806 113004 -2804
rect 148404 -2806 149004 -2804
rect 184404 -2806 185004 -2804
rect 220404 -2806 221004 -2804
rect 256404 -2806 257004 -2804
rect 292404 -2806 293004 -2804
rect 328404 -2806 329004 -2804
rect 364404 -2806 365004 -2804
rect 400404 -2806 401004 -2804
rect 436404 -2806 437004 -2804
rect 472404 -2806 473004 -2804
rect 508404 -2806 509004 -2804
rect 544404 -2806 545004 -2804
rect 580404 -2806 581004 -2804
rect 587200 -2806 587800 -2804
rect -4816 -3144 -4216 -3142
rect 22404 -3144 23004 -3142
rect 58404 -3144 59004 -3142
rect 94404 -3144 95004 -3142
rect 130404 -3144 131004 -3142
rect 166404 -3144 167004 -3142
rect 202404 -3144 203004 -3142
rect 238404 -3144 239004 -3142
rect 274404 -3144 275004 -3142
rect 310404 -3144 311004 -3142
rect 346404 -3144 347004 -3142
rect 382404 -3144 383004 -3142
rect 418404 -3144 419004 -3142
rect 454404 -3144 455004 -3142
rect 490404 -3144 491004 -3142
rect 526404 -3144 527004 -3142
rect 562404 -3144 563004 -3142
rect 588140 -3144 588740 -3142
rect -4816 -3166 588740 -3144
rect -4816 -3402 -4634 -3166
rect -4398 -3402 22586 -3166
rect 22822 -3402 58586 -3166
rect 58822 -3402 94586 -3166
rect 94822 -3402 130586 -3166
rect 130822 -3402 166586 -3166
rect 166822 -3402 202586 -3166
rect 202822 -3402 238586 -3166
rect 238822 -3402 274586 -3166
rect 274822 -3402 310586 -3166
rect 310822 -3402 346586 -3166
rect 346822 -3402 382586 -3166
rect 382822 -3402 418586 -3166
rect 418822 -3402 454586 -3166
rect 454822 -3402 490586 -3166
rect 490822 -3402 526586 -3166
rect 526822 -3402 562586 -3166
rect 562822 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect -4816 -3486 588740 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 22586 -3486
rect 22822 -3722 58586 -3486
rect 58822 -3722 94586 -3486
rect 94822 -3722 130586 -3486
rect 130822 -3722 166586 -3486
rect 166822 -3722 202586 -3486
rect 202822 -3722 238586 -3486
rect 238822 -3722 274586 -3486
rect 274822 -3722 310586 -3486
rect 310822 -3722 346586 -3486
rect 346822 -3722 382586 -3486
rect 382822 -3722 418586 -3486
rect 418822 -3722 454586 -3486
rect 454822 -3722 490586 -3486
rect 490822 -3722 526586 -3486
rect 526822 -3722 562586 -3486
rect 562822 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect -4816 -3744 588740 -3722
rect -4816 -3746 -4216 -3744
rect 22404 -3746 23004 -3744
rect 58404 -3746 59004 -3744
rect 94404 -3746 95004 -3744
rect 130404 -3746 131004 -3744
rect 166404 -3746 167004 -3744
rect 202404 -3746 203004 -3744
rect 238404 -3746 239004 -3744
rect 274404 -3746 275004 -3744
rect 310404 -3746 311004 -3744
rect 346404 -3746 347004 -3744
rect 382404 -3746 383004 -3744
rect 418404 -3746 419004 -3744
rect 454404 -3746 455004 -3744
rect 490404 -3746 491004 -3744
rect 526404 -3746 527004 -3744
rect 562404 -3746 563004 -3744
rect 588140 -3746 588740 -3744
rect -5756 -4084 -5156 -4082
rect 8004 -4084 8604 -4082
rect 44004 -4084 44604 -4082
rect 80004 -4084 80604 -4082
rect 116004 -4084 116604 -4082
rect 152004 -4084 152604 -4082
rect 188004 -4084 188604 -4082
rect 224004 -4084 224604 -4082
rect 260004 -4084 260604 -4082
rect 296004 -4084 296604 -4082
rect 332004 -4084 332604 -4082
rect 368004 -4084 368604 -4082
rect 404004 -4084 404604 -4082
rect 440004 -4084 440604 -4082
rect 476004 -4084 476604 -4082
rect 512004 -4084 512604 -4082
rect 548004 -4084 548604 -4082
rect 589080 -4084 589680 -4082
rect -5756 -4106 589680 -4084
rect -5756 -4342 -5574 -4106
rect -5338 -4342 8186 -4106
rect 8422 -4342 44186 -4106
rect 44422 -4342 80186 -4106
rect 80422 -4342 116186 -4106
rect 116422 -4342 152186 -4106
rect 152422 -4342 188186 -4106
rect 188422 -4342 224186 -4106
rect 224422 -4342 260186 -4106
rect 260422 -4342 296186 -4106
rect 296422 -4342 332186 -4106
rect 332422 -4342 368186 -4106
rect 368422 -4342 404186 -4106
rect 404422 -4342 440186 -4106
rect 440422 -4342 476186 -4106
rect 476422 -4342 512186 -4106
rect 512422 -4342 548186 -4106
rect 548422 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect -5756 -4426 589680 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 8186 -4426
rect 8422 -4662 44186 -4426
rect 44422 -4662 80186 -4426
rect 80422 -4662 116186 -4426
rect 116422 -4662 152186 -4426
rect 152422 -4662 188186 -4426
rect 188422 -4662 224186 -4426
rect 224422 -4662 260186 -4426
rect 260422 -4662 296186 -4426
rect 296422 -4662 332186 -4426
rect 332422 -4662 368186 -4426
rect 368422 -4662 404186 -4426
rect 404422 -4662 440186 -4426
rect 440422 -4662 476186 -4426
rect 476422 -4662 512186 -4426
rect 512422 -4662 548186 -4426
rect 548422 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect -5756 -4684 589680 -4662
rect -5756 -4686 -5156 -4684
rect 8004 -4686 8604 -4684
rect 44004 -4686 44604 -4684
rect 80004 -4686 80604 -4684
rect 116004 -4686 116604 -4684
rect 152004 -4686 152604 -4684
rect 188004 -4686 188604 -4684
rect 224004 -4686 224604 -4684
rect 260004 -4686 260604 -4684
rect 296004 -4686 296604 -4684
rect 332004 -4686 332604 -4684
rect 368004 -4686 368604 -4684
rect 404004 -4686 404604 -4684
rect 440004 -4686 440604 -4684
rect 476004 -4686 476604 -4684
rect 512004 -4686 512604 -4684
rect 548004 -4686 548604 -4684
rect 589080 -4686 589680 -4684
rect -6696 -5024 -6096 -5022
rect 26004 -5024 26604 -5022
rect 62004 -5024 62604 -5022
rect 98004 -5024 98604 -5022
rect 134004 -5024 134604 -5022
rect 170004 -5024 170604 -5022
rect 206004 -5024 206604 -5022
rect 242004 -5024 242604 -5022
rect 278004 -5024 278604 -5022
rect 314004 -5024 314604 -5022
rect 350004 -5024 350604 -5022
rect 386004 -5024 386604 -5022
rect 422004 -5024 422604 -5022
rect 458004 -5024 458604 -5022
rect 494004 -5024 494604 -5022
rect 530004 -5024 530604 -5022
rect 566004 -5024 566604 -5022
rect 590020 -5024 590620 -5022
rect -6696 -5046 590620 -5024
rect -6696 -5282 -6514 -5046
rect -6278 -5282 26186 -5046
rect 26422 -5282 62186 -5046
rect 62422 -5282 98186 -5046
rect 98422 -5282 134186 -5046
rect 134422 -5282 170186 -5046
rect 170422 -5282 206186 -5046
rect 206422 -5282 242186 -5046
rect 242422 -5282 278186 -5046
rect 278422 -5282 314186 -5046
rect 314422 -5282 350186 -5046
rect 350422 -5282 386186 -5046
rect 386422 -5282 422186 -5046
rect 422422 -5282 458186 -5046
rect 458422 -5282 494186 -5046
rect 494422 -5282 530186 -5046
rect 530422 -5282 566186 -5046
rect 566422 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect -6696 -5366 590620 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 26186 -5366
rect 26422 -5602 62186 -5366
rect 62422 -5602 98186 -5366
rect 98422 -5602 134186 -5366
rect 134422 -5602 170186 -5366
rect 170422 -5602 206186 -5366
rect 206422 -5602 242186 -5366
rect 242422 -5602 278186 -5366
rect 278422 -5602 314186 -5366
rect 314422 -5602 350186 -5366
rect 350422 -5602 386186 -5366
rect 386422 -5602 422186 -5366
rect 422422 -5602 458186 -5366
rect 458422 -5602 494186 -5366
rect 494422 -5602 530186 -5366
rect 530422 -5602 566186 -5366
rect 566422 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect -6696 -5624 590620 -5602
rect -6696 -5626 -6096 -5624
rect 26004 -5626 26604 -5624
rect 62004 -5626 62604 -5624
rect 98004 -5626 98604 -5624
rect 134004 -5626 134604 -5624
rect 170004 -5626 170604 -5624
rect 206004 -5626 206604 -5624
rect 242004 -5626 242604 -5624
rect 278004 -5626 278604 -5624
rect 314004 -5626 314604 -5624
rect 350004 -5626 350604 -5624
rect 386004 -5626 386604 -5624
rect 422004 -5626 422604 -5624
rect 458004 -5626 458604 -5624
rect 494004 -5626 494604 -5624
rect 530004 -5626 530604 -5624
rect 566004 -5626 566604 -5624
rect 590020 -5626 590620 -5624
rect -7636 -5964 -7036 -5962
rect 11604 -5964 12204 -5962
rect 47604 -5964 48204 -5962
rect 83604 -5964 84204 -5962
rect 119604 -5964 120204 -5962
rect 155604 -5964 156204 -5962
rect 191604 -5964 192204 -5962
rect 227604 -5964 228204 -5962
rect 263604 -5964 264204 -5962
rect 299604 -5964 300204 -5962
rect 335604 -5964 336204 -5962
rect 371604 -5964 372204 -5962
rect 407604 -5964 408204 -5962
rect 443604 -5964 444204 -5962
rect 479604 -5964 480204 -5962
rect 515604 -5964 516204 -5962
rect 551604 -5964 552204 -5962
rect 590960 -5964 591560 -5962
rect -7636 -5986 591560 -5964
rect -7636 -6222 -7454 -5986
rect -7218 -6222 11786 -5986
rect 12022 -6222 47786 -5986
rect 48022 -6222 83786 -5986
rect 84022 -6222 119786 -5986
rect 120022 -6222 155786 -5986
rect 156022 -6222 191786 -5986
rect 192022 -6222 227786 -5986
rect 228022 -6222 263786 -5986
rect 264022 -6222 299786 -5986
rect 300022 -6222 335786 -5986
rect 336022 -6222 371786 -5986
rect 372022 -6222 407786 -5986
rect 408022 -6222 443786 -5986
rect 444022 -6222 479786 -5986
rect 480022 -6222 515786 -5986
rect 516022 -6222 551786 -5986
rect 552022 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect -7636 -6306 591560 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 11786 -6306
rect 12022 -6542 47786 -6306
rect 48022 -6542 83786 -6306
rect 84022 -6542 119786 -6306
rect 120022 -6542 155786 -6306
rect 156022 -6542 191786 -6306
rect 192022 -6542 227786 -6306
rect 228022 -6542 263786 -6306
rect 264022 -6542 299786 -6306
rect 300022 -6542 335786 -6306
rect 336022 -6542 371786 -6306
rect 372022 -6542 407786 -6306
rect 408022 -6542 443786 -6306
rect 444022 -6542 479786 -6306
rect 480022 -6542 515786 -6306
rect 516022 -6542 551786 -6306
rect 552022 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect -7636 -6564 591560 -6542
rect -7636 -6566 -7036 -6564
rect 11604 -6566 12204 -6564
rect 47604 -6566 48204 -6564
rect 83604 -6566 84204 -6564
rect 119604 -6566 120204 -6564
rect 155604 -6566 156204 -6564
rect 191604 -6566 192204 -6564
rect 227604 -6566 228204 -6564
rect 263604 -6566 264204 -6564
rect 299604 -6566 300204 -6564
rect 335604 -6566 336204 -6564
rect 371604 -6566 372204 -6564
rect 407604 -6566 408204 -6564
rect 443604 -6566 444204 -6564
rect 479604 -6566 480204 -6564
rect 515604 -6566 516204 -6564
rect 551604 -6566 552204 -6564
rect 590960 -6566 591560 -6564
rect -8576 -6904 -7976 -6902
rect 29604 -6904 30204 -6902
rect 65604 -6904 66204 -6902
rect 101604 -6904 102204 -6902
rect 137604 -6904 138204 -6902
rect 173604 -6904 174204 -6902
rect 209604 -6904 210204 -6902
rect 245604 -6904 246204 -6902
rect 281604 -6904 282204 -6902
rect 317604 -6904 318204 -6902
rect 353604 -6904 354204 -6902
rect 389604 -6904 390204 -6902
rect 425604 -6904 426204 -6902
rect 461604 -6904 462204 -6902
rect 497604 -6904 498204 -6902
rect 533604 -6904 534204 -6902
rect 569604 -6904 570204 -6902
rect 591900 -6904 592500 -6902
rect -8576 -6926 592500 -6904
rect -8576 -7162 -8394 -6926
rect -8158 -7162 29786 -6926
rect 30022 -7162 65786 -6926
rect 66022 -7162 101786 -6926
rect 102022 -7162 137786 -6926
rect 138022 -7162 173786 -6926
rect 174022 -7162 209786 -6926
rect 210022 -7162 245786 -6926
rect 246022 -7162 281786 -6926
rect 282022 -7162 317786 -6926
rect 318022 -7162 353786 -6926
rect 354022 -7162 389786 -6926
rect 390022 -7162 425786 -6926
rect 426022 -7162 461786 -6926
rect 462022 -7162 497786 -6926
rect 498022 -7162 533786 -6926
rect 534022 -7162 569786 -6926
rect 570022 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect -8576 -7246 592500 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 29786 -7246
rect 30022 -7482 65786 -7246
rect 66022 -7482 101786 -7246
rect 102022 -7482 137786 -7246
rect 138022 -7482 173786 -7246
rect 174022 -7482 209786 -7246
rect 210022 -7482 245786 -7246
rect 246022 -7482 281786 -7246
rect 282022 -7482 317786 -7246
rect 318022 -7482 353786 -7246
rect 354022 -7482 389786 -7246
rect 390022 -7482 425786 -7246
rect 426022 -7482 461786 -7246
rect 462022 -7482 497786 -7246
rect 498022 -7482 533786 -7246
rect 534022 -7482 569786 -7246
rect 570022 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect -8576 -7504 592500 -7482
rect -8576 -7506 -7976 -7504
rect 29604 -7506 30204 -7504
rect 65604 -7506 66204 -7504
rect 101604 -7506 102204 -7504
rect 137604 -7506 138204 -7504
rect 173604 -7506 174204 -7504
rect 209604 -7506 210204 -7504
rect 245604 -7506 246204 -7504
rect 281604 -7506 282204 -7504
rect 317604 -7506 318204 -7504
rect 353604 -7506 354204 -7504
rect 389604 -7506 390204 -7504
rect 425604 -7506 426204 -7504
rect 461604 -7506 462204 -7504
rect 497604 -7506 498204 -7504
rect 533604 -7506 534204 -7504
rect 569604 -7506 570204 -7504
rect 591900 -7506 592500 -7504
use sram_1rw1r_32_256_8_sky130  sram5
timestamp 1608421104
transform 1 0 450000 0 1 320000
box 0 0 77296 91247
use sram_1rw1r_32_256_8_sky130  sram4
timestamp 1608421104
transform -1 0 417296 0 -1 411247
box 0 0 77296 91247
use sram_1rw1r_32_256_8_sky130  sram3
timestamp 1608421104
transform 1 0 440000 0 1 560000
box 0 0 77296 91247
use sram_1rw1r_32_256_8_sky130  sram2
timestamp 1608421104
transform 1 0 310000 0 1 560000
box 0 0 77296 91247
use sram_1rw1r_32_256_8_sky130  sram1
timestamp 1608421104
transform 1 0 190000 0 1 560000
box 0 0 77296 91247
use sram_1rw1r_32_256_8_sky130  sram0
timestamp 1608421104
transform 1 0 60000 0 1 560000
box 0 0 77296 91247
use hs32_core1  core1
timestamp 1608421104
transform 1 0 60000 0 1 320000
box 0 0 220000 220000
use hs32_core1  core0
timestamp 1608421104
transform 1 0 310000 0 1 80000
box 0 0 220000 220000
<< labels >>
rlabel metal3 s 583520 5796 584960 6036 6 analog_io[0]
port 0 nsew default bidirectional
rlabel metal3 s 583520 474996 584960 475236 6 analog_io[10]
port 1 nsew default bidirectional
rlabel metal3 s 583520 521916 584960 522156 6 analog_io[11]
port 2 nsew default bidirectional
rlabel metal3 s 583520 568836 584960 569076 6 analog_io[12]
port 3 nsew default bidirectional
rlabel metal3 s 583520 615756 584960 615996 6 analog_io[13]
port 4 nsew default bidirectional
rlabel metal3 s 583520 662676 584960 662916 6 analog_io[14]
port 5 nsew default bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[15]
port 6 nsew default bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[16]
port 7 nsew default bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[17]
port 8 nsew default bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[18]
port 9 nsew default bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[19]
port 10 nsew default bidirectional
rlabel metal3 s 583520 52716 584960 52956 6 analog_io[1]
port 11 nsew default bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[20]
port 12 nsew default bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[21]
port 13 nsew default bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[22]
port 14 nsew default bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[23]
port 15 nsew default bidirectional
rlabel metal3 s -960 696540 480 696780 4 analog_io[24]
port 16 nsew default bidirectional
rlabel metal3 s -960 639012 480 639252 4 analog_io[25]
port 17 nsew default bidirectional
rlabel metal3 s -960 581620 480 581860 4 analog_io[26]
port 18 nsew default bidirectional
rlabel metal3 s -960 524092 480 524332 4 analog_io[27]
port 19 nsew default bidirectional
rlabel metal3 s -960 466700 480 466940 4 analog_io[28]
port 20 nsew default bidirectional
rlabel metal3 s -960 409172 480 409412 4 analog_io[29]
port 21 nsew default bidirectional
rlabel metal3 s 583520 99636 584960 99876 6 analog_io[2]
port 22 nsew default bidirectional
rlabel metal3 s -960 351780 480 352020 4 analog_io[30]
port 23 nsew default bidirectional
rlabel metal3 s 583520 146556 584960 146796 6 analog_io[3]
port 24 nsew default bidirectional
rlabel metal3 s 583520 193476 584960 193716 6 analog_io[4]
port 25 nsew default bidirectional
rlabel metal3 s 583520 240396 584960 240636 6 analog_io[5]
port 26 nsew default bidirectional
rlabel metal3 s 583520 287316 584960 287556 6 analog_io[6]
port 27 nsew default bidirectional
rlabel metal3 s 583520 334236 584960 334476 6 analog_io[7]
port 28 nsew default bidirectional
rlabel metal3 s 583520 381156 584960 381396 6 analog_io[8]
port 29 nsew default bidirectional
rlabel metal3 s 583520 428076 584960 428316 6 analog_io[9]
port 30 nsew default bidirectional
rlabel metal3 s 583520 17492 584960 17732 6 io_in[0]
port 31 nsew default input
rlabel metal3 s 583520 486692 584960 486932 6 io_in[10]
port 32 nsew default input
rlabel metal3 s 583520 533748 584960 533988 6 io_in[11]
port 33 nsew default input
rlabel metal3 s 583520 580668 584960 580908 6 io_in[12]
port 34 nsew default input
rlabel metal3 s 583520 627588 584960 627828 6 io_in[13]
port 35 nsew default input
rlabel metal3 s 583520 674508 584960 674748 6 io_in[14]
port 36 nsew default input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 37 nsew default input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 38 nsew default input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 39 nsew default input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 40 nsew default input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 41 nsew default input
rlabel metal3 s 583520 64412 584960 64652 6 io_in[1]
port 42 nsew default input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 43 nsew default input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 44 nsew default input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 45 nsew default input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 46 nsew default input
rlabel metal3 s -960 682124 480 682364 4 io_in[24]
port 47 nsew default input
rlabel metal3 s -960 624732 480 624972 4 io_in[25]
port 48 nsew default input
rlabel metal3 s -960 567204 480 567444 4 io_in[26]
port 49 nsew default input
rlabel metal3 s -960 509812 480 510052 4 io_in[27]
port 50 nsew default input
rlabel metal3 s -960 452284 480 452524 4 io_in[28]
port 51 nsew default input
rlabel metal3 s -960 394892 480 395132 4 io_in[29]
port 52 nsew default input
rlabel metal3 s 583520 111332 584960 111572 6 io_in[2]
port 53 nsew default input
rlabel metal3 s -960 337364 480 337604 4 io_in[30]
port 54 nsew default input
rlabel metal3 s -960 294252 480 294492 4 io_in[31]
port 55 nsew default input
rlabel metal3 s -960 251140 480 251380 4 io_in[32]
port 56 nsew default input
rlabel metal3 s -960 208028 480 208268 4 io_in[33]
port 57 nsew default input
rlabel metal3 s -960 164916 480 165156 4 io_in[34]
port 58 nsew default input
rlabel metal3 s -960 121940 480 122180 4 io_in[35]
port 59 nsew default input
rlabel metal3 s -960 78828 480 79068 4 io_in[36]
port 60 nsew default input
rlabel metal3 s -960 35716 480 35956 4 io_in[37]
port 61 nsew default input
rlabel metal3 s 583520 158252 584960 158492 6 io_in[3]
port 62 nsew default input
rlabel metal3 s 583520 205172 584960 205412 6 io_in[4]
port 63 nsew default input
rlabel metal3 s 583520 252092 584960 252332 6 io_in[5]
port 64 nsew default input
rlabel metal3 s 583520 299012 584960 299252 6 io_in[6]
port 65 nsew default input
rlabel metal3 s 583520 345932 584960 346172 6 io_in[7]
port 66 nsew default input
rlabel metal3 s 583520 392852 584960 393092 6 io_in[8]
port 67 nsew default input
rlabel metal3 s 583520 439772 584960 440012 6 io_in[9]
port 68 nsew default input
rlabel metal3 s 583520 40884 584960 41124 6 io_oeb[0]
port 69 nsew default tristate
rlabel metal3 s 583520 510220 584960 510460 6 io_oeb[10]
port 70 nsew default tristate
rlabel metal3 s 583520 557140 584960 557380 6 io_oeb[11]
port 71 nsew default tristate
rlabel metal3 s 583520 604060 584960 604300 6 io_oeb[12]
port 72 nsew default tristate
rlabel metal3 s 583520 650980 584960 651220 6 io_oeb[13]
port 73 nsew default tristate
rlabel metal3 s 583520 697900 584960 698140 6 io_oeb[14]
port 74 nsew default tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 75 nsew default tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 76 nsew default tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 77 nsew default tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 78 nsew default tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 79 nsew default tristate
rlabel metal3 s 583520 87804 584960 88044 6 io_oeb[1]
port 80 nsew default tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 81 nsew default tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 82 nsew default tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 83 nsew default tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 84 nsew default tristate
rlabel metal3 s -960 653428 480 653668 4 io_oeb[24]
port 85 nsew default tristate
rlabel metal3 s -960 595900 480 596140 4 io_oeb[25]
port 86 nsew default tristate
rlabel metal3 s -960 538508 480 538748 4 io_oeb[26]
port 87 nsew default tristate
rlabel metal3 s -960 480980 480 481220 4 io_oeb[27]
port 88 nsew default tristate
rlabel metal3 s -960 423588 480 423828 4 io_oeb[28]
port 89 nsew default tristate
rlabel metal3 s -960 366060 480 366300 4 io_oeb[29]
port 90 nsew default tristate
rlabel metal3 s 583520 134724 584960 134964 6 io_oeb[2]
port 91 nsew default tristate
rlabel metal3 s -960 308668 480 308908 4 io_oeb[30]
port 92 nsew default tristate
rlabel metal3 s -960 265556 480 265796 4 io_oeb[31]
port 93 nsew default tristate
rlabel metal3 s -960 222444 480 222684 4 io_oeb[32]
port 94 nsew default tristate
rlabel metal3 s -960 179332 480 179572 4 io_oeb[33]
port 95 nsew default tristate
rlabel metal3 s -960 136220 480 136460 4 io_oeb[34]
port 96 nsew default tristate
rlabel metal3 s -960 93108 480 93348 4 io_oeb[35]
port 97 nsew default tristate
rlabel metal3 s -960 49996 480 50236 4 io_oeb[36]
port 98 nsew default tristate
rlabel metal3 s -960 7020 480 7260 4 io_oeb[37]
port 99 nsew default tristate
rlabel metal3 s 583520 181780 584960 182020 6 io_oeb[3]
port 100 nsew default tristate
rlabel metal3 s 583520 228700 584960 228940 6 io_oeb[4]
port 101 nsew default tristate
rlabel metal3 s 583520 275620 584960 275860 6 io_oeb[5]
port 102 nsew default tristate
rlabel metal3 s 583520 322540 584960 322780 6 io_oeb[6]
port 103 nsew default tristate
rlabel metal3 s 583520 369460 584960 369700 6 io_oeb[7]
port 104 nsew default tristate
rlabel metal3 s 583520 416380 584960 416620 6 io_oeb[8]
port 105 nsew default tristate
rlabel metal3 s 583520 463300 584960 463540 6 io_oeb[9]
port 106 nsew default tristate
rlabel metal3 s 583520 29188 584960 29428 6 io_out[0]
port 107 nsew default tristate
rlabel metal3 s 583520 498524 584960 498764 6 io_out[10]
port 108 nsew default tristate
rlabel metal3 s 583520 545444 584960 545684 6 io_out[11]
port 109 nsew default tristate
rlabel metal3 s 583520 592364 584960 592604 6 io_out[12]
port 110 nsew default tristate
rlabel metal3 s 583520 639284 584960 639524 6 io_out[13]
port 111 nsew default tristate
rlabel metal3 s 583520 686204 584960 686444 6 io_out[14]
port 112 nsew default tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 113 nsew default tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 114 nsew default tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 115 nsew default tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 116 nsew default tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 117 nsew default tristate
rlabel metal3 s 583520 76108 584960 76348 6 io_out[1]
port 118 nsew default tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 119 nsew default tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 120 nsew default tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 121 nsew default tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 122 nsew default tristate
rlabel metal3 s -960 667844 480 668084 4 io_out[24]
port 123 nsew default tristate
rlabel metal3 s -960 610316 480 610556 4 io_out[25]
port 124 nsew default tristate
rlabel metal3 s -960 552924 480 553164 4 io_out[26]
port 125 nsew default tristate
rlabel metal3 s -960 495396 480 495636 4 io_out[27]
port 126 nsew default tristate
rlabel metal3 s -960 437868 480 438108 4 io_out[28]
port 127 nsew default tristate
rlabel metal3 s -960 380476 480 380716 4 io_out[29]
port 128 nsew default tristate
rlabel metal3 s 583520 123028 584960 123268 6 io_out[2]
port 129 nsew default tristate
rlabel metal3 s -960 322948 480 323188 4 io_out[30]
port 130 nsew default tristate
rlabel metal3 s -960 279972 480 280212 4 io_out[31]
port 131 nsew default tristate
rlabel metal3 s -960 236860 480 237100 4 io_out[32]
port 132 nsew default tristate
rlabel metal3 s -960 193748 480 193988 4 io_out[33]
port 133 nsew default tristate
rlabel metal3 s -960 150636 480 150876 4 io_out[34]
port 134 nsew default tristate
rlabel metal3 s -960 107524 480 107764 4 io_out[35]
port 135 nsew default tristate
rlabel metal3 s -960 64412 480 64652 4 io_out[36]
port 136 nsew default tristate
rlabel metal3 s -960 21300 480 21540 4 io_out[37]
port 137 nsew default tristate
rlabel metal3 s 583520 169948 584960 170188 6 io_out[3]
port 138 nsew default tristate
rlabel metal3 s 583520 216868 584960 217108 6 io_out[4]
port 139 nsew default tristate
rlabel metal3 s 583520 263788 584960 264028 6 io_out[5]
port 140 nsew default tristate
rlabel metal3 s 583520 310708 584960 310948 6 io_out[6]
port 141 nsew default tristate
rlabel metal3 s 583520 357764 584960 358004 6 io_out[7]
port 142 nsew default tristate
rlabel metal3 s 583520 404684 584960 404924 6 io_out[8]
port 143 nsew default tristate
rlabel metal3 s 583520 451604 584960 451844 6 io_out[9]
port 144 nsew default tristate
rlabel metal2 s 126582 -960 126694 480 8 la_data_in[0]
port 145 nsew default input
rlabel metal2 s 483450 -960 483562 480 8 la_data_in[100]
port 146 nsew default input
rlabel metal2 s 486946 -960 487058 480 8 la_data_in[101]
port 147 nsew default input
rlabel metal2 s 490534 -960 490646 480 8 la_data_in[102]
port 148 nsew default input
rlabel metal2 s 494122 -960 494234 480 8 la_data_in[103]
port 149 nsew default input
rlabel metal2 s 497710 -960 497822 480 8 la_data_in[104]
port 150 nsew default input
rlabel metal2 s 501206 -960 501318 480 8 la_data_in[105]
port 151 nsew default input
rlabel metal2 s 504794 -960 504906 480 8 la_data_in[106]
port 152 nsew default input
rlabel metal2 s 508382 -960 508494 480 8 la_data_in[107]
port 153 nsew default input
rlabel metal2 s 511970 -960 512082 480 8 la_data_in[108]
port 154 nsew default input
rlabel metal2 s 515558 -960 515670 480 8 la_data_in[109]
port 155 nsew default input
rlabel metal2 s 162278 -960 162390 480 8 la_data_in[10]
port 156 nsew default input
rlabel metal2 s 519054 -960 519166 480 8 la_data_in[110]
port 157 nsew default input
rlabel metal2 s 522642 -960 522754 480 8 la_data_in[111]
port 158 nsew default input
rlabel metal2 s 526230 -960 526342 480 8 la_data_in[112]
port 159 nsew default input
rlabel metal2 s 529818 -960 529930 480 8 la_data_in[113]
port 160 nsew default input
rlabel metal2 s 533406 -960 533518 480 8 la_data_in[114]
port 161 nsew default input
rlabel metal2 s 536902 -960 537014 480 8 la_data_in[115]
port 162 nsew default input
rlabel metal2 s 540490 -960 540602 480 8 la_data_in[116]
port 163 nsew default input
rlabel metal2 s 544078 -960 544190 480 8 la_data_in[117]
port 164 nsew default input
rlabel metal2 s 547666 -960 547778 480 8 la_data_in[118]
port 165 nsew default input
rlabel metal2 s 551162 -960 551274 480 8 la_data_in[119]
port 166 nsew default input
rlabel metal2 s 165866 -960 165978 480 8 la_data_in[11]
port 167 nsew default input
rlabel metal2 s 554750 -960 554862 480 8 la_data_in[120]
port 168 nsew default input
rlabel metal2 s 558338 -960 558450 480 8 la_data_in[121]
port 169 nsew default input
rlabel metal2 s 561926 -960 562038 480 8 la_data_in[122]
port 170 nsew default input
rlabel metal2 s 565514 -960 565626 480 8 la_data_in[123]
port 171 nsew default input
rlabel metal2 s 569010 -960 569122 480 8 la_data_in[124]
port 172 nsew default input
rlabel metal2 s 572598 -960 572710 480 8 la_data_in[125]
port 173 nsew default input
rlabel metal2 s 576186 -960 576298 480 8 la_data_in[126]
port 174 nsew default input
rlabel metal2 s 579774 -960 579886 480 8 la_data_in[127]
port 175 nsew default input
rlabel metal2 s 169362 -960 169474 480 8 la_data_in[12]
port 176 nsew default input
rlabel metal2 s 172950 -960 173062 480 8 la_data_in[13]
port 177 nsew default input
rlabel metal2 s 176538 -960 176650 480 8 la_data_in[14]
port 178 nsew default input
rlabel metal2 s 180126 -960 180238 480 8 la_data_in[15]
port 179 nsew default input
rlabel metal2 s 183714 -960 183826 480 8 la_data_in[16]
port 180 nsew default input
rlabel metal2 s 187210 -960 187322 480 8 la_data_in[17]
port 181 nsew default input
rlabel metal2 s 190798 -960 190910 480 8 la_data_in[18]
port 182 nsew default input
rlabel metal2 s 194386 -960 194498 480 8 la_data_in[19]
port 183 nsew default input
rlabel metal2 s 130170 -960 130282 480 8 la_data_in[1]
port 184 nsew default input
rlabel metal2 s 197974 -960 198086 480 8 la_data_in[20]
port 185 nsew default input
rlabel metal2 s 201470 -960 201582 480 8 la_data_in[21]
port 186 nsew default input
rlabel metal2 s 205058 -960 205170 480 8 la_data_in[22]
port 187 nsew default input
rlabel metal2 s 208646 -960 208758 480 8 la_data_in[23]
port 188 nsew default input
rlabel metal2 s 212234 -960 212346 480 8 la_data_in[24]
port 189 nsew default input
rlabel metal2 s 215822 -960 215934 480 8 la_data_in[25]
port 190 nsew default input
rlabel metal2 s 219318 -960 219430 480 8 la_data_in[26]
port 191 nsew default input
rlabel metal2 s 222906 -960 223018 480 8 la_data_in[27]
port 192 nsew default input
rlabel metal2 s 226494 -960 226606 480 8 la_data_in[28]
port 193 nsew default input
rlabel metal2 s 230082 -960 230194 480 8 la_data_in[29]
port 194 nsew default input
rlabel metal2 s 133758 -960 133870 480 8 la_data_in[2]
port 195 nsew default input
rlabel metal2 s 233670 -960 233782 480 8 la_data_in[30]
port 196 nsew default input
rlabel metal2 s 237166 -960 237278 480 8 la_data_in[31]
port 197 nsew default input
rlabel metal2 s 240754 -960 240866 480 8 la_data_in[32]
port 198 nsew default input
rlabel metal2 s 244342 -960 244454 480 8 la_data_in[33]
port 199 nsew default input
rlabel metal2 s 247930 -960 248042 480 8 la_data_in[34]
port 200 nsew default input
rlabel metal2 s 251426 -960 251538 480 8 la_data_in[35]
port 201 nsew default input
rlabel metal2 s 255014 -960 255126 480 8 la_data_in[36]
port 202 nsew default input
rlabel metal2 s 258602 -960 258714 480 8 la_data_in[37]
port 203 nsew default input
rlabel metal2 s 262190 -960 262302 480 8 la_data_in[38]
port 204 nsew default input
rlabel metal2 s 265778 -960 265890 480 8 la_data_in[39]
port 205 nsew default input
rlabel metal2 s 137254 -960 137366 480 8 la_data_in[3]
port 206 nsew default input
rlabel metal2 s 269274 -960 269386 480 8 la_data_in[40]
port 207 nsew default input
rlabel metal2 s 272862 -960 272974 480 8 la_data_in[41]
port 208 nsew default input
rlabel metal2 s 276450 -960 276562 480 8 la_data_in[42]
port 209 nsew default input
rlabel metal2 s 280038 -960 280150 480 8 la_data_in[43]
port 210 nsew default input
rlabel metal2 s 283626 -960 283738 480 8 la_data_in[44]
port 211 nsew default input
rlabel metal2 s 287122 -960 287234 480 8 la_data_in[45]
port 212 nsew default input
rlabel metal2 s 290710 -960 290822 480 8 la_data_in[46]
port 213 nsew default input
rlabel metal2 s 294298 -960 294410 480 8 la_data_in[47]
port 214 nsew default input
rlabel metal2 s 297886 -960 297998 480 8 la_data_in[48]
port 215 nsew default input
rlabel metal2 s 301382 -960 301494 480 8 la_data_in[49]
port 216 nsew default input
rlabel metal2 s 140842 -960 140954 480 8 la_data_in[4]
port 217 nsew default input
rlabel metal2 s 304970 -960 305082 480 8 la_data_in[50]
port 218 nsew default input
rlabel metal2 s 308558 -960 308670 480 8 la_data_in[51]
port 219 nsew default input
rlabel metal2 s 312146 -960 312258 480 8 la_data_in[52]
port 220 nsew default input
rlabel metal2 s 315734 -960 315846 480 8 la_data_in[53]
port 221 nsew default input
rlabel metal2 s 319230 -960 319342 480 8 la_data_in[54]
port 222 nsew default input
rlabel metal2 s 322818 -960 322930 480 8 la_data_in[55]
port 223 nsew default input
rlabel metal2 s 326406 -960 326518 480 8 la_data_in[56]
port 224 nsew default input
rlabel metal2 s 329994 -960 330106 480 8 la_data_in[57]
port 225 nsew default input
rlabel metal2 s 333582 -960 333694 480 8 la_data_in[58]
port 226 nsew default input
rlabel metal2 s 337078 -960 337190 480 8 la_data_in[59]
port 227 nsew default input
rlabel metal2 s 144430 -960 144542 480 8 la_data_in[5]
port 228 nsew default input
rlabel metal2 s 340666 -960 340778 480 8 la_data_in[60]
port 229 nsew default input
rlabel metal2 s 344254 -960 344366 480 8 la_data_in[61]
port 230 nsew default input
rlabel metal2 s 347842 -960 347954 480 8 la_data_in[62]
port 231 nsew default input
rlabel metal2 s 351338 -960 351450 480 8 la_data_in[63]
port 232 nsew default input
rlabel metal2 s 354926 -960 355038 480 8 la_data_in[64]
port 233 nsew default input
rlabel metal2 s 358514 -960 358626 480 8 la_data_in[65]
port 234 nsew default input
rlabel metal2 s 362102 -960 362214 480 8 la_data_in[66]
port 235 nsew default input
rlabel metal2 s 365690 -960 365802 480 8 la_data_in[67]
port 236 nsew default input
rlabel metal2 s 369186 -960 369298 480 8 la_data_in[68]
port 237 nsew default input
rlabel metal2 s 372774 -960 372886 480 8 la_data_in[69]
port 238 nsew default input
rlabel metal2 s 148018 -960 148130 480 8 la_data_in[6]
port 239 nsew default input
rlabel metal2 s 376362 -960 376474 480 8 la_data_in[70]
port 240 nsew default input
rlabel metal2 s 379950 -960 380062 480 8 la_data_in[71]
port 241 nsew default input
rlabel metal2 s 383538 -960 383650 480 8 la_data_in[72]
port 242 nsew default input
rlabel metal2 s 387034 -960 387146 480 8 la_data_in[73]
port 243 nsew default input
rlabel metal2 s 390622 -960 390734 480 8 la_data_in[74]
port 244 nsew default input
rlabel metal2 s 394210 -960 394322 480 8 la_data_in[75]
port 245 nsew default input
rlabel metal2 s 397798 -960 397910 480 8 la_data_in[76]
port 246 nsew default input
rlabel metal2 s 401294 -960 401406 480 8 la_data_in[77]
port 247 nsew default input
rlabel metal2 s 404882 -960 404994 480 8 la_data_in[78]
port 248 nsew default input
rlabel metal2 s 408470 -960 408582 480 8 la_data_in[79]
port 249 nsew default input
rlabel metal2 s 151514 -960 151626 480 8 la_data_in[7]
port 250 nsew default input
rlabel metal2 s 412058 -960 412170 480 8 la_data_in[80]
port 251 nsew default input
rlabel metal2 s 415646 -960 415758 480 8 la_data_in[81]
port 252 nsew default input
rlabel metal2 s 419142 -960 419254 480 8 la_data_in[82]
port 253 nsew default input
rlabel metal2 s 422730 -960 422842 480 8 la_data_in[83]
port 254 nsew default input
rlabel metal2 s 426318 -960 426430 480 8 la_data_in[84]
port 255 nsew default input
rlabel metal2 s 429906 -960 430018 480 8 la_data_in[85]
port 256 nsew default input
rlabel metal2 s 433494 -960 433606 480 8 la_data_in[86]
port 257 nsew default input
rlabel metal2 s 436990 -960 437102 480 8 la_data_in[87]
port 258 nsew default input
rlabel metal2 s 440578 -960 440690 480 8 la_data_in[88]
port 259 nsew default input
rlabel metal2 s 444166 -960 444278 480 8 la_data_in[89]
port 260 nsew default input
rlabel metal2 s 155102 -960 155214 480 8 la_data_in[8]
port 261 nsew default input
rlabel metal2 s 447754 -960 447866 480 8 la_data_in[90]
port 262 nsew default input
rlabel metal2 s 451250 -960 451362 480 8 la_data_in[91]
port 263 nsew default input
rlabel metal2 s 454838 -960 454950 480 8 la_data_in[92]
port 264 nsew default input
rlabel metal2 s 458426 -960 458538 480 8 la_data_in[93]
port 265 nsew default input
rlabel metal2 s 462014 -960 462126 480 8 la_data_in[94]
port 266 nsew default input
rlabel metal2 s 465602 -960 465714 480 8 la_data_in[95]
port 267 nsew default input
rlabel metal2 s 469098 -960 469210 480 8 la_data_in[96]
port 268 nsew default input
rlabel metal2 s 472686 -960 472798 480 8 la_data_in[97]
port 269 nsew default input
rlabel metal2 s 476274 -960 476386 480 8 la_data_in[98]
port 270 nsew default input
rlabel metal2 s 479862 -960 479974 480 8 la_data_in[99]
port 271 nsew default input
rlabel metal2 s 158690 -960 158802 480 8 la_data_in[9]
port 272 nsew default input
rlabel metal2 s 127778 -960 127890 480 8 la_data_out[0]
port 273 nsew default tristate
rlabel metal2 s 484554 -960 484666 480 8 la_data_out[100]
port 274 nsew default tristate
rlabel metal2 s 488142 -960 488254 480 8 la_data_out[101]
port 275 nsew default tristate
rlabel metal2 s 491730 -960 491842 480 8 la_data_out[102]
port 276 nsew default tristate
rlabel metal2 s 495318 -960 495430 480 8 la_data_out[103]
port 277 nsew default tristate
rlabel metal2 s 498906 -960 499018 480 8 la_data_out[104]
port 278 nsew default tristate
rlabel metal2 s 502402 -960 502514 480 8 la_data_out[105]
port 279 nsew default tristate
rlabel metal2 s 505990 -960 506102 480 8 la_data_out[106]
port 280 nsew default tristate
rlabel metal2 s 509578 -960 509690 480 8 la_data_out[107]
port 281 nsew default tristate
rlabel metal2 s 513166 -960 513278 480 8 la_data_out[108]
port 282 nsew default tristate
rlabel metal2 s 516754 -960 516866 480 8 la_data_out[109]
port 283 nsew default tristate
rlabel metal2 s 163474 -960 163586 480 8 la_data_out[10]
port 284 nsew default tristate
rlabel metal2 s 520250 -960 520362 480 8 la_data_out[110]
port 285 nsew default tristate
rlabel metal2 s 523838 -960 523950 480 8 la_data_out[111]
port 286 nsew default tristate
rlabel metal2 s 527426 -960 527538 480 8 la_data_out[112]
port 287 nsew default tristate
rlabel metal2 s 531014 -960 531126 480 8 la_data_out[113]
port 288 nsew default tristate
rlabel metal2 s 534510 -960 534622 480 8 la_data_out[114]
port 289 nsew default tristate
rlabel metal2 s 538098 -960 538210 480 8 la_data_out[115]
port 290 nsew default tristate
rlabel metal2 s 541686 -960 541798 480 8 la_data_out[116]
port 291 nsew default tristate
rlabel metal2 s 545274 -960 545386 480 8 la_data_out[117]
port 292 nsew default tristate
rlabel metal2 s 548862 -960 548974 480 8 la_data_out[118]
port 293 nsew default tristate
rlabel metal2 s 552358 -960 552470 480 8 la_data_out[119]
port 294 nsew default tristate
rlabel metal2 s 167062 -960 167174 480 8 la_data_out[11]
port 295 nsew default tristate
rlabel metal2 s 555946 -960 556058 480 8 la_data_out[120]
port 296 nsew default tristate
rlabel metal2 s 559534 -960 559646 480 8 la_data_out[121]
port 297 nsew default tristate
rlabel metal2 s 563122 -960 563234 480 8 la_data_out[122]
port 298 nsew default tristate
rlabel metal2 s 566710 -960 566822 480 8 la_data_out[123]
port 299 nsew default tristate
rlabel metal2 s 570206 -960 570318 480 8 la_data_out[124]
port 300 nsew default tristate
rlabel metal2 s 573794 -960 573906 480 8 la_data_out[125]
port 301 nsew default tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[126]
port 302 nsew default tristate
rlabel metal2 s 580970 -960 581082 480 8 la_data_out[127]
port 303 nsew default tristate
rlabel metal2 s 170558 -960 170670 480 8 la_data_out[12]
port 304 nsew default tristate
rlabel metal2 s 174146 -960 174258 480 8 la_data_out[13]
port 305 nsew default tristate
rlabel metal2 s 177734 -960 177846 480 8 la_data_out[14]
port 306 nsew default tristate
rlabel metal2 s 181322 -960 181434 480 8 la_data_out[15]
port 307 nsew default tristate
rlabel metal2 s 184818 -960 184930 480 8 la_data_out[16]
port 308 nsew default tristate
rlabel metal2 s 188406 -960 188518 480 8 la_data_out[17]
port 309 nsew default tristate
rlabel metal2 s 191994 -960 192106 480 8 la_data_out[18]
port 310 nsew default tristate
rlabel metal2 s 195582 -960 195694 480 8 la_data_out[19]
port 311 nsew default tristate
rlabel metal2 s 131366 -960 131478 480 8 la_data_out[1]
port 312 nsew default tristate
rlabel metal2 s 199170 -960 199282 480 8 la_data_out[20]
port 313 nsew default tristate
rlabel metal2 s 202666 -960 202778 480 8 la_data_out[21]
port 314 nsew default tristate
rlabel metal2 s 206254 -960 206366 480 8 la_data_out[22]
port 315 nsew default tristate
rlabel metal2 s 209842 -960 209954 480 8 la_data_out[23]
port 316 nsew default tristate
rlabel metal2 s 213430 -960 213542 480 8 la_data_out[24]
port 317 nsew default tristate
rlabel metal2 s 217018 -960 217130 480 8 la_data_out[25]
port 318 nsew default tristate
rlabel metal2 s 220514 -960 220626 480 8 la_data_out[26]
port 319 nsew default tristate
rlabel metal2 s 224102 -960 224214 480 8 la_data_out[27]
port 320 nsew default tristate
rlabel metal2 s 227690 -960 227802 480 8 la_data_out[28]
port 321 nsew default tristate
rlabel metal2 s 231278 -960 231390 480 8 la_data_out[29]
port 322 nsew default tristate
rlabel metal2 s 134862 -960 134974 480 8 la_data_out[2]
port 323 nsew default tristate
rlabel metal2 s 234774 -960 234886 480 8 la_data_out[30]
port 324 nsew default tristate
rlabel metal2 s 238362 -960 238474 480 8 la_data_out[31]
port 325 nsew default tristate
rlabel metal2 s 241950 -960 242062 480 8 la_data_out[32]
port 326 nsew default tristate
rlabel metal2 s 245538 -960 245650 480 8 la_data_out[33]
port 327 nsew default tristate
rlabel metal2 s 249126 -960 249238 480 8 la_data_out[34]
port 328 nsew default tristate
rlabel metal2 s 252622 -960 252734 480 8 la_data_out[35]
port 329 nsew default tristate
rlabel metal2 s 256210 -960 256322 480 8 la_data_out[36]
port 330 nsew default tristate
rlabel metal2 s 259798 -960 259910 480 8 la_data_out[37]
port 331 nsew default tristate
rlabel metal2 s 263386 -960 263498 480 8 la_data_out[38]
port 332 nsew default tristate
rlabel metal2 s 266974 -960 267086 480 8 la_data_out[39]
port 333 nsew default tristate
rlabel metal2 s 138450 -960 138562 480 8 la_data_out[3]
port 334 nsew default tristate
rlabel metal2 s 270470 -960 270582 480 8 la_data_out[40]
port 335 nsew default tristate
rlabel metal2 s 274058 -960 274170 480 8 la_data_out[41]
port 336 nsew default tristate
rlabel metal2 s 277646 -960 277758 480 8 la_data_out[42]
port 337 nsew default tristate
rlabel metal2 s 281234 -960 281346 480 8 la_data_out[43]
port 338 nsew default tristate
rlabel metal2 s 284730 -960 284842 480 8 la_data_out[44]
port 339 nsew default tristate
rlabel metal2 s 288318 -960 288430 480 8 la_data_out[45]
port 340 nsew default tristate
rlabel metal2 s 291906 -960 292018 480 8 la_data_out[46]
port 341 nsew default tristate
rlabel metal2 s 295494 -960 295606 480 8 la_data_out[47]
port 342 nsew default tristate
rlabel metal2 s 299082 -960 299194 480 8 la_data_out[48]
port 343 nsew default tristate
rlabel metal2 s 302578 -960 302690 480 8 la_data_out[49]
port 344 nsew default tristate
rlabel metal2 s 142038 -960 142150 480 8 la_data_out[4]
port 345 nsew default tristate
rlabel metal2 s 306166 -960 306278 480 8 la_data_out[50]
port 346 nsew default tristate
rlabel metal2 s 309754 -960 309866 480 8 la_data_out[51]
port 347 nsew default tristate
rlabel metal2 s 313342 -960 313454 480 8 la_data_out[52]
port 348 nsew default tristate
rlabel metal2 s 316930 -960 317042 480 8 la_data_out[53]
port 349 nsew default tristate
rlabel metal2 s 320426 -960 320538 480 8 la_data_out[54]
port 350 nsew default tristate
rlabel metal2 s 324014 -960 324126 480 8 la_data_out[55]
port 351 nsew default tristate
rlabel metal2 s 327602 -960 327714 480 8 la_data_out[56]
port 352 nsew default tristate
rlabel metal2 s 331190 -960 331302 480 8 la_data_out[57]
port 353 nsew default tristate
rlabel metal2 s 334686 -960 334798 480 8 la_data_out[58]
port 354 nsew default tristate
rlabel metal2 s 338274 -960 338386 480 8 la_data_out[59]
port 355 nsew default tristate
rlabel metal2 s 145626 -960 145738 480 8 la_data_out[5]
port 356 nsew default tristate
rlabel metal2 s 341862 -960 341974 480 8 la_data_out[60]
port 357 nsew default tristate
rlabel metal2 s 345450 -960 345562 480 8 la_data_out[61]
port 358 nsew default tristate
rlabel metal2 s 349038 -960 349150 480 8 la_data_out[62]
port 359 nsew default tristate
rlabel metal2 s 352534 -960 352646 480 8 la_data_out[63]
port 360 nsew default tristate
rlabel metal2 s 356122 -960 356234 480 8 la_data_out[64]
port 361 nsew default tristate
rlabel metal2 s 359710 -960 359822 480 8 la_data_out[65]
port 362 nsew default tristate
rlabel metal2 s 363298 -960 363410 480 8 la_data_out[66]
port 363 nsew default tristate
rlabel metal2 s 366886 -960 366998 480 8 la_data_out[67]
port 364 nsew default tristate
rlabel metal2 s 370382 -960 370494 480 8 la_data_out[68]
port 365 nsew default tristate
rlabel metal2 s 373970 -960 374082 480 8 la_data_out[69]
port 366 nsew default tristate
rlabel metal2 s 149214 -960 149326 480 8 la_data_out[6]
port 367 nsew default tristate
rlabel metal2 s 377558 -960 377670 480 8 la_data_out[70]
port 368 nsew default tristate
rlabel metal2 s 381146 -960 381258 480 8 la_data_out[71]
port 369 nsew default tristate
rlabel metal2 s 384642 -960 384754 480 8 la_data_out[72]
port 370 nsew default tristate
rlabel metal2 s 388230 -960 388342 480 8 la_data_out[73]
port 371 nsew default tristate
rlabel metal2 s 391818 -960 391930 480 8 la_data_out[74]
port 372 nsew default tristate
rlabel metal2 s 395406 -960 395518 480 8 la_data_out[75]
port 373 nsew default tristate
rlabel metal2 s 398994 -960 399106 480 8 la_data_out[76]
port 374 nsew default tristate
rlabel metal2 s 402490 -960 402602 480 8 la_data_out[77]
port 375 nsew default tristate
rlabel metal2 s 406078 -960 406190 480 8 la_data_out[78]
port 376 nsew default tristate
rlabel metal2 s 409666 -960 409778 480 8 la_data_out[79]
port 377 nsew default tristate
rlabel metal2 s 152710 -960 152822 480 8 la_data_out[7]
port 378 nsew default tristate
rlabel metal2 s 413254 -960 413366 480 8 la_data_out[80]
port 379 nsew default tristate
rlabel metal2 s 416842 -960 416954 480 8 la_data_out[81]
port 380 nsew default tristate
rlabel metal2 s 420338 -960 420450 480 8 la_data_out[82]
port 381 nsew default tristate
rlabel metal2 s 423926 -960 424038 480 8 la_data_out[83]
port 382 nsew default tristate
rlabel metal2 s 427514 -960 427626 480 8 la_data_out[84]
port 383 nsew default tristate
rlabel metal2 s 431102 -960 431214 480 8 la_data_out[85]
port 384 nsew default tristate
rlabel metal2 s 434598 -960 434710 480 8 la_data_out[86]
port 385 nsew default tristate
rlabel metal2 s 438186 -960 438298 480 8 la_data_out[87]
port 386 nsew default tristate
rlabel metal2 s 441774 -960 441886 480 8 la_data_out[88]
port 387 nsew default tristate
rlabel metal2 s 445362 -960 445474 480 8 la_data_out[89]
port 388 nsew default tristate
rlabel metal2 s 156298 -960 156410 480 8 la_data_out[8]
port 389 nsew default tristate
rlabel metal2 s 448950 -960 449062 480 8 la_data_out[90]
port 390 nsew default tristate
rlabel metal2 s 452446 -960 452558 480 8 la_data_out[91]
port 391 nsew default tristate
rlabel metal2 s 456034 -960 456146 480 8 la_data_out[92]
port 392 nsew default tristate
rlabel metal2 s 459622 -960 459734 480 8 la_data_out[93]
port 393 nsew default tristate
rlabel metal2 s 463210 -960 463322 480 8 la_data_out[94]
port 394 nsew default tristate
rlabel metal2 s 466798 -960 466910 480 8 la_data_out[95]
port 395 nsew default tristate
rlabel metal2 s 470294 -960 470406 480 8 la_data_out[96]
port 396 nsew default tristate
rlabel metal2 s 473882 -960 473994 480 8 la_data_out[97]
port 397 nsew default tristate
rlabel metal2 s 477470 -960 477582 480 8 la_data_out[98]
port 398 nsew default tristate
rlabel metal2 s 481058 -960 481170 480 8 la_data_out[99]
port 399 nsew default tristate
rlabel metal2 s 159886 -960 159998 480 8 la_data_out[9]
port 400 nsew default tristate
rlabel metal2 s 128974 -960 129086 480 8 la_oen[0]
port 401 nsew default input
rlabel metal2 s 485750 -960 485862 480 8 la_oen[100]
port 402 nsew default input
rlabel metal2 s 489338 -960 489450 480 8 la_oen[101]
port 403 nsew default input
rlabel metal2 s 492926 -960 493038 480 8 la_oen[102]
port 404 nsew default input
rlabel metal2 s 496514 -960 496626 480 8 la_oen[103]
port 405 nsew default input
rlabel metal2 s 500102 -960 500214 480 8 la_oen[104]
port 406 nsew default input
rlabel metal2 s 503598 -960 503710 480 8 la_oen[105]
port 407 nsew default input
rlabel metal2 s 507186 -960 507298 480 8 la_oen[106]
port 408 nsew default input
rlabel metal2 s 510774 -960 510886 480 8 la_oen[107]
port 409 nsew default input
rlabel metal2 s 514362 -960 514474 480 8 la_oen[108]
port 410 nsew default input
rlabel metal2 s 517858 -960 517970 480 8 la_oen[109]
port 411 nsew default input
rlabel metal2 s 164670 -960 164782 480 8 la_oen[10]
port 412 nsew default input
rlabel metal2 s 521446 -960 521558 480 8 la_oen[110]
port 413 nsew default input
rlabel metal2 s 525034 -960 525146 480 8 la_oen[111]
port 414 nsew default input
rlabel metal2 s 528622 -960 528734 480 8 la_oen[112]
port 415 nsew default input
rlabel metal2 s 532210 -960 532322 480 8 la_oen[113]
port 416 nsew default input
rlabel metal2 s 535706 -960 535818 480 8 la_oen[114]
port 417 nsew default input
rlabel metal2 s 539294 -960 539406 480 8 la_oen[115]
port 418 nsew default input
rlabel metal2 s 542882 -960 542994 480 8 la_oen[116]
port 419 nsew default input
rlabel metal2 s 546470 -960 546582 480 8 la_oen[117]
port 420 nsew default input
rlabel metal2 s 550058 -960 550170 480 8 la_oen[118]
port 421 nsew default input
rlabel metal2 s 553554 -960 553666 480 8 la_oen[119]
port 422 nsew default input
rlabel metal2 s 168166 -960 168278 480 8 la_oen[11]
port 423 nsew default input
rlabel metal2 s 557142 -960 557254 480 8 la_oen[120]
port 424 nsew default input
rlabel metal2 s 560730 -960 560842 480 8 la_oen[121]
port 425 nsew default input
rlabel metal2 s 564318 -960 564430 480 8 la_oen[122]
port 426 nsew default input
rlabel metal2 s 567814 -960 567926 480 8 la_oen[123]
port 427 nsew default input
rlabel metal2 s 571402 -960 571514 480 8 la_oen[124]
port 428 nsew default input
rlabel metal2 s 574990 -960 575102 480 8 la_oen[125]
port 429 nsew default input
rlabel metal2 s 578578 -960 578690 480 8 la_oen[126]
port 430 nsew default input
rlabel metal2 s 582166 -960 582278 480 8 la_oen[127]
port 431 nsew default input
rlabel metal2 s 171754 -960 171866 480 8 la_oen[12]
port 432 nsew default input
rlabel metal2 s 175342 -960 175454 480 8 la_oen[13]
port 433 nsew default input
rlabel metal2 s 178930 -960 179042 480 8 la_oen[14]
port 434 nsew default input
rlabel metal2 s 182518 -960 182630 480 8 la_oen[15]
port 435 nsew default input
rlabel metal2 s 186014 -960 186126 480 8 la_oen[16]
port 436 nsew default input
rlabel metal2 s 189602 -960 189714 480 8 la_oen[17]
port 437 nsew default input
rlabel metal2 s 193190 -960 193302 480 8 la_oen[18]
port 438 nsew default input
rlabel metal2 s 196778 -960 196890 480 8 la_oen[19]
port 439 nsew default input
rlabel metal2 s 132562 -960 132674 480 8 la_oen[1]
port 440 nsew default input
rlabel metal2 s 200366 -960 200478 480 8 la_oen[20]
port 441 nsew default input
rlabel metal2 s 203862 -960 203974 480 8 la_oen[21]
port 442 nsew default input
rlabel metal2 s 207450 -960 207562 480 8 la_oen[22]
port 443 nsew default input
rlabel metal2 s 211038 -960 211150 480 8 la_oen[23]
port 444 nsew default input
rlabel metal2 s 214626 -960 214738 480 8 la_oen[24]
port 445 nsew default input
rlabel metal2 s 218122 -960 218234 480 8 la_oen[25]
port 446 nsew default input
rlabel metal2 s 221710 -960 221822 480 8 la_oen[26]
port 447 nsew default input
rlabel metal2 s 225298 -960 225410 480 8 la_oen[27]
port 448 nsew default input
rlabel metal2 s 228886 -960 228998 480 8 la_oen[28]
port 449 nsew default input
rlabel metal2 s 232474 -960 232586 480 8 la_oen[29]
port 450 nsew default input
rlabel metal2 s 136058 -960 136170 480 8 la_oen[2]
port 451 nsew default input
rlabel metal2 s 235970 -960 236082 480 8 la_oen[30]
port 452 nsew default input
rlabel metal2 s 239558 -960 239670 480 8 la_oen[31]
port 453 nsew default input
rlabel metal2 s 243146 -960 243258 480 8 la_oen[32]
port 454 nsew default input
rlabel metal2 s 246734 -960 246846 480 8 la_oen[33]
port 455 nsew default input
rlabel metal2 s 250322 -960 250434 480 8 la_oen[34]
port 456 nsew default input
rlabel metal2 s 253818 -960 253930 480 8 la_oen[35]
port 457 nsew default input
rlabel metal2 s 257406 -960 257518 480 8 la_oen[36]
port 458 nsew default input
rlabel metal2 s 260994 -960 261106 480 8 la_oen[37]
port 459 nsew default input
rlabel metal2 s 264582 -960 264694 480 8 la_oen[38]
port 460 nsew default input
rlabel metal2 s 268078 -960 268190 480 8 la_oen[39]
port 461 nsew default input
rlabel metal2 s 139646 -960 139758 480 8 la_oen[3]
port 462 nsew default input
rlabel metal2 s 271666 -960 271778 480 8 la_oen[40]
port 463 nsew default input
rlabel metal2 s 275254 -960 275366 480 8 la_oen[41]
port 464 nsew default input
rlabel metal2 s 278842 -960 278954 480 8 la_oen[42]
port 465 nsew default input
rlabel metal2 s 282430 -960 282542 480 8 la_oen[43]
port 466 nsew default input
rlabel metal2 s 285926 -960 286038 480 8 la_oen[44]
port 467 nsew default input
rlabel metal2 s 289514 -960 289626 480 8 la_oen[45]
port 468 nsew default input
rlabel metal2 s 293102 -960 293214 480 8 la_oen[46]
port 469 nsew default input
rlabel metal2 s 296690 -960 296802 480 8 la_oen[47]
port 470 nsew default input
rlabel metal2 s 300278 -960 300390 480 8 la_oen[48]
port 471 nsew default input
rlabel metal2 s 303774 -960 303886 480 8 la_oen[49]
port 472 nsew default input
rlabel metal2 s 143234 -960 143346 480 8 la_oen[4]
port 473 nsew default input
rlabel metal2 s 307362 -960 307474 480 8 la_oen[50]
port 474 nsew default input
rlabel metal2 s 310950 -960 311062 480 8 la_oen[51]
port 475 nsew default input
rlabel metal2 s 314538 -960 314650 480 8 la_oen[52]
port 476 nsew default input
rlabel metal2 s 318034 -960 318146 480 8 la_oen[53]
port 477 nsew default input
rlabel metal2 s 321622 -960 321734 480 8 la_oen[54]
port 478 nsew default input
rlabel metal2 s 325210 -960 325322 480 8 la_oen[55]
port 479 nsew default input
rlabel metal2 s 328798 -960 328910 480 8 la_oen[56]
port 480 nsew default input
rlabel metal2 s 332386 -960 332498 480 8 la_oen[57]
port 481 nsew default input
rlabel metal2 s 335882 -960 335994 480 8 la_oen[58]
port 482 nsew default input
rlabel metal2 s 339470 -960 339582 480 8 la_oen[59]
port 483 nsew default input
rlabel metal2 s 146822 -960 146934 480 8 la_oen[5]
port 484 nsew default input
rlabel metal2 s 343058 -960 343170 480 8 la_oen[60]
port 485 nsew default input
rlabel metal2 s 346646 -960 346758 480 8 la_oen[61]
port 486 nsew default input
rlabel metal2 s 350234 -960 350346 480 8 la_oen[62]
port 487 nsew default input
rlabel metal2 s 353730 -960 353842 480 8 la_oen[63]
port 488 nsew default input
rlabel metal2 s 357318 -960 357430 480 8 la_oen[64]
port 489 nsew default input
rlabel metal2 s 360906 -960 361018 480 8 la_oen[65]
port 490 nsew default input
rlabel metal2 s 364494 -960 364606 480 8 la_oen[66]
port 491 nsew default input
rlabel metal2 s 367990 -960 368102 480 8 la_oen[67]
port 492 nsew default input
rlabel metal2 s 371578 -960 371690 480 8 la_oen[68]
port 493 nsew default input
rlabel metal2 s 375166 -960 375278 480 8 la_oen[69]
port 494 nsew default input
rlabel metal2 s 150410 -960 150522 480 8 la_oen[6]
port 495 nsew default input
rlabel metal2 s 378754 -960 378866 480 8 la_oen[70]
port 496 nsew default input
rlabel metal2 s 382342 -960 382454 480 8 la_oen[71]
port 497 nsew default input
rlabel metal2 s 385838 -960 385950 480 8 la_oen[72]
port 498 nsew default input
rlabel metal2 s 389426 -960 389538 480 8 la_oen[73]
port 499 nsew default input
rlabel metal2 s 393014 -960 393126 480 8 la_oen[74]
port 500 nsew default input
rlabel metal2 s 396602 -960 396714 480 8 la_oen[75]
port 501 nsew default input
rlabel metal2 s 400190 -960 400302 480 8 la_oen[76]
port 502 nsew default input
rlabel metal2 s 403686 -960 403798 480 8 la_oen[77]
port 503 nsew default input
rlabel metal2 s 407274 -960 407386 480 8 la_oen[78]
port 504 nsew default input
rlabel metal2 s 410862 -960 410974 480 8 la_oen[79]
port 505 nsew default input
rlabel metal2 s 153906 -960 154018 480 8 la_oen[7]
port 506 nsew default input
rlabel metal2 s 414450 -960 414562 480 8 la_oen[80]
port 507 nsew default input
rlabel metal2 s 417946 -960 418058 480 8 la_oen[81]
port 508 nsew default input
rlabel metal2 s 421534 -960 421646 480 8 la_oen[82]
port 509 nsew default input
rlabel metal2 s 425122 -960 425234 480 8 la_oen[83]
port 510 nsew default input
rlabel metal2 s 428710 -960 428822 480 8 la_oen[84]
port 511 nsew default input
rlabel metal2 s 432298 -960 432410 480 8 la_oen[85]
port 512 nsew default input
rlabel metal2 s 435794 -960 435906 480 8 la_oen[86]
port 513 nsew default input
rlabel metal2 s 439382 -960 439494 480 8 la_oen[87]
port 514 nsew default input
rlabel metal2 s 442970 -960 443082 480 8 la_oen[88]
port 515 nsew default input
rlabel metal2 s 446558 -960 446670 480 8 la_oen[89]
port 516 nsew default input
rlabel metal2 s 157494 -960 157606 480 8 la_oen[8]
port 517 nsew default input
rlabel metal2 s 450146 -960 450258 480 8 la_oen[90]
port 518 nsew default input
rlabel metal2 s 453642 -960 453754 480 8 la_oen[91]
port 519 nsew default input
rlabel metal2 s 457230 -960 457342 480 8 la_oen[92]
port 520 nsew default input
rlabel metal2 s 460818 -960 460930 480 8 la_oen[93]
port 521 nsew default input
rlabel metal2 s 464406 -960 464518 480 8 la_oen[94]
port 522 nsew default input
rlabel metal2 s 467902 -960 468014 480 8 la_oen[95]
port 523 nsew default input
rlabel metal2 s 471490 -960 471602 480 8 la_oen[96]
port 524 nsew default input
rlabel metal2 s 475078 -960 475190 480 8 la_oen[97]
port 525 nsew default input
rlabel metal2 s 478666 -960 478778 480 8 la_oen[98]
port 526 nsew default input
rlabel metal2 s 482254 -960 482366 480 8 la_oen[99]
port 527 nsew default input
rlabel metal2 s 161082 -960 161194 480 8 la_oen[9]
port 528 nsew default input
rlabel metal2 s 583362 -960 583474 480 8 user_clock2
port 529 nsew default input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 530 nsew default input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 531 nsew default input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 532 nsew default tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 533 nsew default input
rlabel metal2 s 48106 -960 48218 480 8 wbs_adr_i[10]
port 534 nsew default input
rlabel metal2 s 51602 -960 51714 480 8 wbs_adr_i[11]
port 535 nsew default input
rlabel metal2 s 55190 -960 55302 480 8 wbs_adr_i[12]
port 536 nsew default input
rlabel metal2 s 58778 -960 58890 480 8 wbs_adr_i[13]
port 537 nsew default input
rlabel metal2 s 62366 -960 62478 480 8 wbs_adr_i[14]
port 538 nsew default input
rlabel metal2 s 65954 -960 66066 480 8 wbs_adr_i[15]
port 539 nsew default input
rlabel metal2 s 69450 -960 69562 480 8 wbs_adr_i[16]
port 540 nsew default input
rlabel metal2 s 73038 -960 73150 480 8 wbs_adr_i[17]
port 541 nsew default input
rlabel metal2 s 76626 -960 76738 480 8 wbs_adr_i[18]
port 542 nsew default input
rlabel metal2 s 80214 -960 80326 480 8 wbs_adr_i[19]
port 543 nsew default input
rlabel metal2 s 12410 -960 12522 480 8 wbs_adr_i[1]
port 544 nsew default input
rlabel metal2 s 83802 -960 83914 480 8 wbs_adr_i[20]
port 545 nsew default input
rlabel metal2 s 87298 -960 87410 480 8 wbs_adr_i[21]
port 546 nsew default input
rlabel metal2 s 90886 -960 90998 480 8 wbs_adr_i[22]
port 547 nsew default input
rlabel metal2 s 94474 -960 94586 480 8 wbs_adr_i[23]
port 548 nsew default input
rlabel metal2 s 98062 -960 98174 480 8 wbs_adr_i[24]
port 549 nsew default input
rlabel metal2 s 101558 -960 101670 480 8 wbs_adr_i[25]
port 550 nsew default input
rlabel metal2 s 105146 -960 105258 480 8 wbs_adr_i[26]
port 551 nsew default input
rlabel metal2 s 108734 -960 108846 480 8 wbs_adr_i[27]
port 552 nsew default input
rlabel metal2 s 112322 -960 112434 480 8 wbs_adr_i[28]
port 553 nsew default input
rlabel metal2 s 115910 -960 116022 480 8 wbs_adr_i[29]
port 554 nsew default input
rlabel metal2 s 17194 -960 17306 480 8 wbs_adr_i[2]
port 555 nsew default input
rlabel metal2 s 119406 -960 119518 480 8 wbs_adr_i[30]
port 556 nsew default input
rlabel metal2 s 122994 -960 123106 480 8 wbs_adr_i[31]
port 557 nsew default input
rlabel metal2 s 21886 -960 21998 480 8 wbs_adr_i[3]
port 558 nsew default input
rlabel metal2 s 26670 -960 26782 480 8 wbs_adr_i[4]
port 559 nsew default input
rlabel metal2 s 30258 -960 30370 480 8 wbs_adr_i[5]
port 560 nsew default input
rlabel metal2 s 33846 -960 33958 480 8 wbs_adr_i[6]
port 561 nsew default input
rlabel metal2 s 37342 -960 37454 480 8 wbs_adr_i[7]
port 562 nsew default input
rlabel metal2 s 40930 -960 41042 480 8 wbs_adr_i[8]
port 563 nsew default input
rlabel metal2 s 44518 -960 44630 480 8 wbs_adr_i[9]
port 564 nsew default input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 565 nsew default input
rlabel metal2 s 8822 -960 8934 480 8 wbs_dat_i[0]
port 566 nsew default input
rlabel metal2 s 49302 -960 49414 480 8 wbs_dat_i[10]
port 567 nsew default input
rlabel metal2 s 52798 -960 52910 480 8 wbs_dat_i[11]
port 568 nsew default input
rlabel metal2 s 56386 -960 56498 480 8 wbs_dat_i[12]
port 569 nsew default input
rlabel metal2 s 59974 -960 60086 480 8 wbs_dat_i[13]
port 570 nsew default input
rlabel metal2 s 63562 -960 63674 480 8 wbs_dat_i[14]
port 571 nsew default input
rlabel metal2 s 67150 -960 67262 480 8 wbs_dat_i[15]
port 572 nsew default input
rlabel metal2 s 70646 -960 70758 480 8 wbs_dat_i[16]
port 573 nsew default input
rlabel metal2 s 74234 -960 74346 480 8 wbs_dat_i[17]
port 574 nsew default input
rlabel metal2 s 77822 -960 77934 480 8 wbs_dat_i[18]
port 575 nsew default input
rlabel metal2 s 81410 -960 81522 480 8 wbs_dat_i[19]
port 576 nsew default input
rlabel metal2 s 13606 -960 13718 480 8 wbs_dat_i[1]
port 577 nsew default input
rlabel metal2 s 84906 -960 85018 480 8 wbs_dat_i[20]
port 578 nsew default input
rlabel metal2 s 88494 -960 88606 480 8 wbs_dat_i[21]
port 579 nsew default input
rlabel metal2 s 92082 -960 92194 480 8 wbs_dat_i[22]
port 580 nsew default input
rlabel metal2 s 95670 -960 95782 480 8 wbs_dat_i[23]
port 581 nsew default input
rlabel metal2 s 99258 -960 99370 480 8 wbs_dat_i[24]
port 582 nsew default input
rlabel metal2 s 102754 -960 102866 480 8 wbs_dat_i[25]
port 583 nsew default input
rlabel metal2 s 106342 -960 106454 480 8 wbs_dat_i[26]
port 584 nsew default input
rlabel metal2 s 109930 -960 110042 480 8 wbs_dat_i[27]
port 585 nsew default input
rlabel metal2 s 113518 -960 113630 480 8 wbs_dat_i[28]
port 586 nsew default input
rlabel metal2 s 117106 -960 117218 480 8 wbs_dat_i[29]
port 587 nsew default input
rlabel metal2 s 18298 -960 18410 480 8 wbs_dat_i[2]
port 588 nsew default input
rlabel metal2 s 120602 -960 120714 480 8 wbs_dat_i[30]
port 589 nsew default input
rlabel metal2 s 124190 -960 124302 480 8 wbs_dat_i[31]
port 590 nsew default input
rlabel metal2 s 23082 -960 23194 480 8 wbs_dat_i[3]
port 591 nsew default input
rlabel metal2 s 27866 -960 27978 480 8 wbs_dat_i[4]
port 592 nsew default input
rlabel metal2 s 31454 -960 31566 480 8 wbs_dat_i[5]
port 593 nsew default input
rlabel metal2 s 34950 -960 35062 480 8 wbs_dat_i[6]
port 594 nsew default input
rlabel metal2 s 38538 -960 38650 480 8 wbs_dat_i[7]
port 595 nsew default input
rlabel metal2 s 42126 -960 42238 480 8 wbs_dat_i[8]
port 596 nsew default input
rlabel metal2 s 45714 -960 45826 480 8 wbs_dat_i[9]
port 597 nsew default input
rlabel metal2 s 10018 -960 10130 480 8 wbs_dat_o[0]
port 598 nsew default tristate
rlabel metal2 s 50498 -960 50610 480 8 wbs_dat_o[10]
port 599 nsew default tristate
rlabel metal2 s 53994 -960 54106 480 8 wbs_dat_o[11]
port 600 nsew default tristate
rlabel metal2 s 57582 -960 57694 480 8 wbs_dat_o[12]
port 601 nsew default tristate
rlabel metal2 s 61170 -960 61282 480 8 wbs_dat_o[13]
port 602 nsew default tristate
rlabel metal2 s 64758 -960 64870 480 8 wbs_dat_o[14]
port 603 nsew default tristate
rlabel metal2 s 68254 -960 68366 480 8 wbs_dat_o[15]
port 604 nsew default tristate
rlabel metal2 s 71842 -960 71954 480 8 wbs_dat_o[16]
port 605 nsew default tristate
rlabel metal2 s 75430 -960 75542 480 8 wbs_dat_o[17]
port 606 nsew default tristate
rlabel metal2 s 79018 -960 79130 480 8 wbs_dat_o[18]
port 607 nsew default tristate
rlabel metal2 s 82606 -960 82718 480 8 wbs_dat_o[19]
port 608 nsew default tristate
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[1]
port 609 nsew default tristate
rlabel metal2 s 86102 -960 86214 480 8 wbs_dat_o[20]
port 610 nsew default tristate
rlabel metal2 s 89690 -960 89802 480 8 wbs_dat_o[21]
port 611 nsew default tristate
rlabel metal2 s 93278 -960 93390 480 8 wbs_dat_o[22]
port 612 nsew default tristate
rlabel metal2 s 96866 -960 96978 480 8 wbs_dat_o[23]
port 613 nsew default tristate
rlabel metal2 s 100454 -960 100566 480 8 wbs_dat_o[24]
port 614 nsew default tristate
rlabel metal2 s 103950 -960 104062 480 8 wbs_dat_o[25]
port 615 nsew default tristate
rlabel metal2 s 107538 -960 107650 480 8 wbs_dat_o[26]
port 616 nsew default tristate
rlabel metal2 s 111126 -960 111238 480 8 wbs_dat_o[27]
port 617 nsew default tristate
rlabel metal2 s 114714 -960 114826 480 8 wbs_dat_o[28]
port 618 nsew default tristate
rlabel metal2 s 118210 -960 118322 480 8 wbs_dat_o[29]
port 619 nsew default tristate
rlabel metal2 s 19494 -960 19606 480 8 wbs_dat_o[2]
port 620 nsew default tristate
rlabel metal2 s 121798 -960 121910 480 8 wbs_dat_o[30]
port 621 nsew default tristate
rlabel metal2 s 125386 -960 125498 480 8 wbs_dat_o[31]
port 622 nsew default tristate
rlabel metal2 s 24278 -960 24390 480 8 wbs_dat_o[3]
port 623 nsew default tristate
rlabel metal2 s 29062 -960 29174 480 8 wbs_dat_o[4]
port 624 nsew default tristate
rlabel metal2 s 32650 -960 32762 480 8 wbs_dat_o[5]
port 625 nsew default tristate
rlabel metal2 s 36146 -960 36258 480 8 wbs_dat_o[6]
port 626 nsew default tristate
rlabel metal2 s 39734 -960 39846 480 8 wbs_dat_o[7]
port 627 nsew default tristate
rlabel metal2 s 43322 -960 43434 480 8 wbs_dat_o[8]
port 628 nsew default tristate
rlabel metal2 s 46910 -960 47022 480 8 wbs_dat_o[9]
port 629 nsew default tristate
rlabel metal2 s 11214 -960 11326 480 8 wbs_sel_i[0]
port 630 nsew default input
rlabel metal2 s 15998 -960 16110 480 8 wbs_sel_i[1]
port 631 nsew default input
rlabel metal2 s 20690 -960 20802 480 8 wbs_sel_i[2]
port 632 nsew default input
rlabel metal2 s 25474 -960 25586 480 8 wbs_sel_i[3]
port 633 nsew default input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 634 nsew default input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 635 nsew default input
rlabel metal5 s -1996 -924 585920 -324 8 vccd1
port 636 nsew default input
rlabel metal5 s -2936 -1864 586860 -1264 8 vssd1
port 637 nsew default input
rlabel metal5 s -3876 -2804 587800 -2204 8 vccd2
port 638 nsew default input
rlabel metal5 s -4816 -3744 588740 -3144 8 vssd2
port 639 nsew default input
rlabel metal5 s -5756 -4684 589680 -4084 8 vdda1
port 640 nsew default input
rlabel metal5 s -6696 -5624 590620 -5024 8 vssa1
port 641 nsew default input
rlabel metal5 s -7636 -6564 591560 -5964 8 vdda2
port 642 nsew default input
rlabel metal5 s -8576 -7504 592500 -6904 8 vssa2
port 643 nsew default input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
