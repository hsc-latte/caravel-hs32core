VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO hs32_core1
  CLASS BLOCK ;
  FOREIGN hs32_core1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1100.000 BY 1100.000 ;
  PIN cpu_addr_e[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 67.360 1100.000 67.960 ;
    END
  END cpu_addr_e[0]
  PIN cpu_addr_e[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 117.680 1100.000 118.280 ;
    END
  END cpu_addr_e[10]
  PIN cpu_addr_e[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 123.120 1100.000 123.720 ;
    END
  END cpu_addr_e[11]
  PIN cpu_addr_e[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 127.880 1100.000 128.480 ;
    END
  END cpu_addr_e[12]
  PIN cpu_addr_e[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 132.640 1100.000 133.240 ;
    END
  END cpu_addr_e[13]
  PIN cpu_addr_e[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 138.080 1100.000 138.680 ;
    END
  END cpu_addr_e[14]
  PIN cpu_addr_e[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 142.840 1100.000 143.440 ;
    END
  END cpu_addr_e[15]
  PIN cpu_addr_e[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 72.120 1100.000 72.720 ;
    END
  END cpu_addr_e[1]
  PIN cpu_addr_e[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 77.560 1100.000 78.160 ;
    END
  END cpu_addr_e[2]
  PIN cpu_addr_e[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 82.320 1100.000 82.920 ;
    END
  END cpu_addr_e[3]
  PIN cpu_addr_e[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 87.760 1100.000 88.360 ;
    END
  END cpu_addr_e[4]
  PIN cpu_addr_e[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 92.520 1100.000 93.120 ;
    END
  END cpu_addr_e[5]
  PIN cpu_addr_e[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 97.960 1100.000 98.560 ;
    END
  END cpu_addr_e[6]
  PIN cpu_addr_e[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 102.720 1100.000 103.320 ;
    END
  END cpu_addr_e[7]
  PIN cpu_addr_e[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 107.480 1100.000 108.080 ;
    END
  END cpu_addr_e[8]
  PIN cpu_addr_e[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 112.920 1100.000 113.520 ;
    END
  END cpu_addr_e[9]
  PIN cpu_addr_n[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 108.650 1096.000 108.930 1100.000 ;
    END
  END cpu_addr_n[0]
  PIN cpu_addr_n[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 212.610 1096.000 212.890 1100.000 ;
    END
  END cpu_addr_n[10]
  PIN cpu_addr_n[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 222.730 1096.000 223.010 1100.000 ;
    END
  END cpu_addr_n[11]
  PIN cpu_addr_n[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 233.310 1096.000 233.590 1100.000 ;
    END
  END cpu_addr_n[12]
  PIN cpu_addr_n[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 243.430 1096.000 243.710 1100.000 ;
    END
  END cpu_addr_n[13]
  PIN cpu_addr_n[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 254.010 1096.000 254.290 1100.000 ;
    END
  END cpu_addr_n[14]
  PIN cpu_addr_n[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 264.130 1096.000 264.410 1100.000 ;
    END
  END cpu_addr_n[15]
  PIN cpu_addr_n[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 119.230 1096.000 119.510 1100.000 ;
    END
  END cpu_addr_n[1]
  PIN cpu_addr_n[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 129.350 1096.000 129.630 1100.000 ;
    END
  END cpu_addr_n[2]
  PIN cpu_addr_n[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 139.930 1096.000 140.210 1100.000 ;
    END
  END cpu_addr_n[3]
  PIN cpu_addr_n[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 150.050 1096.000 150.330 1100.000 ;
    END
  END cpu_addr_n[4]
  PIN cpu_addr_n[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 160.630 1096.000 160.910 1100.000 ;
    END
  END cpu_addr_n[5]
  PIN cpu_addr_n[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 170.750 1096.000 171.030 1100.000 ;
    END
  END cpu_addr_n[6]
  PIN cpu_addr_n[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 181.330 1096.000 181.610 1100.000 ;
    END
  END cpu_addr_n[7]
  PIN cpu_addr_n[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 191.910 1096.000 192.190 1100.000 ;
    END
  END cpu_addr_n[8]
  PIN cpu_addr_n[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 202.030 1096.000 202.310 1100.000 ;
    END
  END cpu_addr_n[9]
  PIN cpu_dtr_e0[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 228.520 1100.000 229.120 ;
    END
  END cpu_dtr_e0[0]
  PIN cpu_dtr_e0[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 279.520 1100.000 280.120 ;
    END
  END cpu_dtr_e0[10]
  PIN cpu_dtr_e0[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 284.280 1100.000 284.880 ;
    END
  END cpu_dtr_e0[11]
  PIN cpu_dtr_e0[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 289.720 1100.000 290.320 ;
    END
  END cpu_dtr_e0[12]
  PIN cpu_dtr_e0[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 294.480 1100.000 295.080 ;
    END
  END cpu_dtr_e0[13]
  PIN cpu_dtr_e0[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 299.240 1100.000 299.840 ;
    END
  END cpu_dtr_e0[14]
  PIN cpu_dtr_e0[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 304.680 1100.000 305.280 ;
    END
  END cpu_dtr_e0[15]
  PIN cpu_dtr_e0[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 309.440 1100.000 310.040 ;
    END
  END cpu_dtr_e0[16]
  PIN cpu_dtr_e0[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 314.880 1100.000 315.480 ;
    END
  END cpu_dtr_e0[17]
  PIN cpu_dtr_e0[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 319.640 1100.000 320.240 ;
    END
  END cpu_dtr_e0[18]
  PIN cpu_dtr_e0[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 325.080 1100.000 325.680 ;
    END
  END cpu_dtr_e0[19]
  PIN cpu_dtr_e0[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 233.960 1100.000 234.560 ;
    END
  END cpu_dtr_e0[1]
  PIN cpu_dtr_e0[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 329.840 1100.000 330.440 ;
    END
  END cpu_dtr_e0[20]
  PIN cpu_dtr_e0[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 334.600 1100.000 335.200 ;
    END
  END cpu_dtr_e0[21]
  PIN cpu_dtr_e0[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 340.040 1100.000 340.640 ;
    END
  END cpu_dtr_e0[22]
  PIN cpu_dtr_e0[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 344.800 1100.000 345.400 ;
    END
  END cpu_dtr_e0[23]
  PIN cpu_dtr_e0[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 350.240 1100.000 350.840 ;
    END
  END cpu_dtr_e0[24]
  PIN cpu_dtr_e0[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 355.000 1100.000 355.600 ;
    END
  END cpu_dtr_e0[25]
  PIN cpu_dtr_e0[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 359.760 1100.000 360.360 ;
    END
  END cpu_dtr_e0[26]
  PIN cpu_dtr_e0[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 365.200 1100.000 365.800 ;
    END
  END cpu_dtr_e0[27]
  PIN cpu_dtr_e0[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 369.960 1100.000 370.560 ;
    END
  END cpu_dtr_e0[28]
  PIN cpu_dtr_e0[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 375.400 1100.000 376.000 ;
    END
  END cpu_dtr_e0[29]
  PIN cpu_dtr_e0[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 238.720 1100.000 239.320 ;
    END
  END cpu_dtr_e0[2]
  PIN cpu_dtr_e0[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 380.160 1100.000 380.760 ;
    END
  END cpu_dtr_e0[30]
  PIN cpu_dtr_e0[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 385.600 1100.000 386.200 ;
    END
  END cpu_dtr_e0[31]
  PIN cpu_dtr_e0[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 244.160 1100.000 244.760 ;
    END
  END cpu_dtr_e0[3]
  PIN cpu_dtr_e0[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 248.920 1100.000 249.520 ;
    END
  END cpu_dtr_e0[4]
  PIN cpu_dtr_e0[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 254.360 1100.000 254.960 ;
    END
  END cpu_dtr_e0[5]
  PIN cpu_dtr_e0[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 259.120 1100.000 259.720 ;
    END
  END cpu_dtr_e0[6]
  PIN cpu_dtr_e0[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 263.880 1100.000 264.480 ;
    END
  END cpu_dtr_e0[7]
  PIN cpu_dtr_e0[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 269.320 1100.000 269.920 ;
    END
  END cpu_dtr_e0[8]
  PIN cpu_dtr_e0[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 274.080 1100.000 274.680 ;
    END
  END cpu_dtr_e0[9]
  PIN cpu_dtr_e1[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 390.360 1100.000 390.960 ;
    END
  END cpu_dtr_e1[0]
  PIN cpu_dtr_e1[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 440.680 1100.000 441.280 ;
    END
  END cpu_dtr_e1[10]
  PIN cpu_dtr_e1[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 446.120 1100.000 446.720 ;
    END
  END cpu_dtr_e1[11]
  PIN cpu_dtr_e1[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 450.880 1100.000 451.480 ;
    END
  END cpu_dtr_e1[12]
  PIN cpu_dtr_e1[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 455.640 1100.000 456.240 ;
    END
  END cpu_dtr_e1[13]
  PIN cpu_dtr_e1[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 461.080 1100.000 461.680 ;
    END
  END cpu_dtr_e1[14]
  PIN cpu_dtr_e1[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 465.840 1100.000 466.440 ;
    END
  END cpu_dtr_e1[15]
  PIN cpu_dtr_e1[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 471.280 1100.000 471.880 ;
    END
  END cpu_dtr_e1[16]
  PIN cpu_dtr_e1[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 476.040 1100.000 476.640 ;
    END
  END cpu_dtr_e1[17]
  PIN cpu_dtr_e1[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 481.480 1100.000 482.080 ;
    END
  END cpu_dtr_e1[18]
  PIN cpu_dtr_e1[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 486.240 1100.000 486.840 ;
    END
  END cpu_dtr_e1[19]
  PIN cpu_dtr_e1[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 395.120 1100.000 395.720 ;
    END
  END cpu_dtr_e1[1]
  PIN cpu_dtr_e1[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 491.000 1100.000 491.600 ;
    END
  END cpu_dtr_e1[20]
  PIN cpu_dtr_e1[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 496.440 1100.000 497.040 ;
    END
  END cpu_dtr_e1[21]
  PIN cpu_dtr_e1[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 501.200 1100.000 501.800 ;
    END
  END cpu_dtr_e1[22]
  PIN cpu_dtr_e1[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 506.640 1100.000 507.240 ;
    END
  END cpu_dtr_e1[23]
  PIN cpu_dtr_e1[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 511.400 1100.000 512.000 ;
    END
  END cpu_dtr_e1[24]
  PIN cpu_dtr_e1[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 516.840 1100.000 517.440 ;
    END
  END cpu_dtr_e1[25]
  PIN cpu_dtr_e1[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 521.600 1100.000 522.200 ;
    END
  END cpu_dtr_e1[26]
  PIN cpu_dtr_e1[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 526.360 1100.000 526.960 ;
    END
  END cpu_dtr_e1[27]
  PIN cpu_dtr_e1[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 531.800 1100.000 532.400 ;
    END
  END cpu_dtr_e1[28]
  PIN cpu_dtr_e1[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 536.560 1100.000 537.160 ;
    END
  END cpu_dtr_e1[29]
  PIN cpu_dtr_e1[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 400.560 1100.000 401.160 ;
    END
  END cpu_dtr_e1[2]
  PIN cpu_dtr_e1[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 542.000 1100.000 542.600 ;
    END
  END cpu_dtr_e1[30]
  PIN cpu_dtr_e1[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 546.760 1100.000 547.360 ;
    END
  END cpu_dtr_e1[31]
  PIN cpu_dtr_e1[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 405.320 1100.000 405.920 ;
    END
  END cpu_dtr_e1[3]
  PIN cpu_dtr_e1[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 410.760 1100.000 411.360 ;
    END
  END cpu_dtr_e1[4]
  PIN cpu_dtr_e1[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 415.520 1100.000 416.120 ;
    END
  END cpu_dtr_e1[5]
  PIN cpu_dtr_e1[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 420.960 1100.000 421.560 ;
    END
  END cpu_dtr_e1[6]
  PIN cpu_dtr_e1[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 425.720 1100.000 426.320 ;
    END
  END cpu_dtr_e1[7]
  PIN cpu_dtr_e1[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 430.480 1100.000 431.080 ;
    END
  END cpu_dtr_e1[8]
  PIN cpu_dtr_e1[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 435.920 1100.000 436.520 ;
    END
  END cpu_dtr_e1[9]
  PIN cpu_dtr_n0[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 440.770 1096.000 441.050 1100.000 ;
    END
  END cpu_dtr_n0[0]
  PIN cpu_dtr_n0[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 544.270 1096.000 544.550 1100.000 ;
    END
  END cpu_dtr_n0[10]
  PIN cpu_dtr_n0[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 554.850 1096.000 555.130 1100.000 ;
    END
  END cpu_dtr_n0[11]
  PIN cpu_dtr_n0[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 565.430 1096.000 565.710 1100.000 ;
    END
  END cpu_dtr_n0[12]
  PIN cpu_dtr_n0[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 575.550 1096.000 575.830 1100.000 ;
    END
  END cpu_dtr_n0[13]
  PIN cpu_dtr_n0[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 586.130 1096.000 586.410 1100.000 ;
    END
  END cpu_dtr_n0[14]
  PIN cpu_dtr_n0[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 596.250 1096.000 596.530 1100.000 ;
    END
  END cpu_dtr_n0[15]
  PIN cpu_dtr_n0[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 606.830 1096.000 607.110 1100.000 ;
    END
  END cpu_dtr_n0[16]
  PIN cpu_dtr_n0[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 616.950 1096.000 617.230 1100.000 ;
    END
  END cpu_dtr_n0[17]
  PIN cpu_dtr_n0[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 627.530 1096.000 627.810 1100.000 ;
    END
  END cpu_dtr_n0[18]
  PIN cpu_dtr_n0[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 637.650 1096.000 637.930 1100.000 ;
    END
  END cpu_dtr_n0[19]
  PIN cpu_dtr_n0[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 450.890 1096.000 451.170 1100.000 ;
    END
  END cpu_dtr_n0[1]
  PIN cpu_dtr_n0[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 648.230 1096.000 648.510 1100.000 ;
    END
  END cpu_dtr_n0[20]
  PIN cpu_dtr_n0[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 658.810 1096.000 659.090 1100.000 ;
    END
  END cpu_dtr_n0[21]
  PIN cpu_dtr_n0[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 668.930 1096.000 669.210 1100.000 ;
    END
  END cpu_dtr_n0[22]
  PIN cpu_dtr_n0[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 679.510 1096.000 679.790 1100.000 ;
    END
  END cpu_dtr_n0[23]
  PIN cpu_dtr_n0[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 689.630 1096.000 689.910 1100.000 ;
    END
  END cpu_dtr_n0[24]
  PIN cpu_dtr_n0[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 700.210 1096.000 700.490 1100.000 ;
    END
  END cpu_dtr_n0[25]
  PIN cpu_dtr_n0[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 710.330 1096.000 710.610 1100.000 ;
    END
  END cpu_dtr_n0[26]
  PIN cpu_dtr_n0[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 720.910 1096.000 721.190 1100.000 ;
    END
  END cpu_dtr_n0[27]
  PIN cpu_dtr_n0[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 731.030 1096.000 731.310 1100.000 ;
    END
  END cpu_dtr_n0[28]
  PIN cpu_dtr_n0[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 741.610 1096.000 741.890 1100.000 ;
    END
  END cpu_dtr_n0[29]
  PIN cpu_dtr_n0[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 461.470 1096.000 461.750 1100.000 ;
    END
  END cpu_dtr_n0[2]
  PIN cpu_dtr_n0[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 752.190 1096.000 752.470 1100.000 ;
    END
  END cpu_dtr_n0[30]
  PIN cpu_dtr_n0[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 762.310 1096.000 762.590 1100.000 ;
    END
  END cpu_dtr_n0[31]
  PIN cpu_dtr_n0[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 472.050 1096.000 472.330 1100.000 ;
    END
  END cpu_dtr_n0[3]
  PIN cpu_dtr_n0[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 482.170 1096.000 482.450 1100.000 ;
    END
  END cpu_dtr_n0[4]
  PIN cpu_dtr_n0[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 492.750 1096.000 493.030 1100.000 ;
    END
  END cpu_dtr_n0[5]
  PIN cpu_dtr_n0[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 502.870 1096.000 503.150 1100.000 ;
    END
  END cpu_dtr_n0[6]
  PIN cpu_dtr_n0[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 513.450 1096.000 513.730 1100.000 ;
    END
  END cpu_dtr_n0[7]
  PIN cpu_dtr_n0[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 523.570 1096.000 523.850 1100.000 ;
    END
  END cpu_dtr_n0[8]
  PIN cpu_dtr_n0[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 534.150 1096.000 534.430 1100.000 ;
    END
  END cpu_dtr_n0[9]
  PIN cpu_dtr_n1[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 772.890 1096.000 773.170 1100.000 ;
    END
  END cpu_dtr_n1[0]
  PIN cpu_dtr_n1[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 876.390 1096.000 876.670 1100.000 ;
    END
  END cpu_dtr_n1[10]
  PIN cpu_dtr_n1[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 886.970 1096.000 887.250 1100.000 ;
    END
  END cpu_dtr_n1[11]
  PIN cpu_dtr_n1[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 897.090 1096.000 897.370 1100.000 ;
    END
  END cpu_dtr_n1[12]
  PIN cpu_dtr_n1[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 907.670 1096.000 907.950 1100.000 ;
    END
  END cpu_dtr_n1[13]
  PIN cpu_dtr_n1[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 917.790 1096.000 918.070 1100.000 ;
    END
  END cpu_dtr_n1[14]
  PIN cpu_dtr_n1[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 928.370 1096.000 928.650 1100.000 ;
    END
  END cpu_dtr_n1[15]
  PIN cpu_dtr_n1[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 938.950 1096.000 939.230 1100.000 ;
    END
  END cpu_dtr_n1[16]
  PIN cpu_dtr_n1[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 949.070 1096.000 949.350 1100.000 ;
    END
  END cpu_dtr_n1[17]
  PIN cpu_dtr_n1[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 959.650 1096.000 959.930 1100.000 ;
    END
  END cpu_dtr_n1[18]
  PIN cpu_dtr_n1[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 969.770 1096.000 970.050 1100.000 ;
    END
  END cpu_dtr_n1[19]
  PIN cpu_dtr_n1[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 783.010 1096.000 783.290 1100.000 ;
    END
  END cpu_dtr_n1[1]
  PIN cpu_dtr_n1[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 980.350 1096.000 980.630 1100.000 ;
    END
  END cpu_dtr_n1[20]
  PIN cpu_dtr_n1[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 990.470 1096.000 990.750 1100.000 ;
    END
  END cpu_dtr_n1[21]
  PIN cpu_dtr_n1[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1001.050 1096.000 1001.330 1100.000 ;
    END
  END cpu_dtr_n1[22]
  PIN cpu_dtr_n1[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1011.170 1096.000 1011.450 1100.000 ;
    END
  END cpu_dtr_n1[23]
  PIN cpu_dtr_n1[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1021.750 1096.000 1022.030 1100.000 ;
    END
  END cpu_dtr_n1[24]
  PIN cpu_dtr_n1[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1032.330 1096.000 1032.610 1100.000 ;
    END
  END cpu_dtr_n1[25]
  PIN cpu_dtr_n1[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1042.450 1096.000 1042.730 1100.000 ;
    END
  END cpu_dtr_n1[26]
  PIN cpu_dtr_n1[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1053.030 1096.000 1053.310 1100.000 ;
    END
  END cpu_dtr_n1[27]
  PIN cpu_dtr_n1[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1063.150 1096.000 1063.430 1100.000 ;
    END
  END cpu_dtr_n1[28]
  PIN cpu_dtr_n1[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1073.730 1096.000 1074.010 1100.000 ;
    END
  END cpu_dtr_n1[29]
  PIN cpu_dtr_n1[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 793.590 1096.000 793.870 1100.000 ;
    END
  END cpu_dtr_n1[2]
  PIN cpu_dtr_n1[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1083.850 1096.000 1084.130 1100.000 ;
    END
  END cpu_dtr_n1[30]
  PIN cpu_dtr_n1[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1094.430 1096.000 1094.710 1100.000 ;
    END
  END cpu_dtr_n1[31]
  PIN cpu_dtr_n1[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 803.710 1096.000 803.990 1100.000 ;
    END
  END cpu_dtr_n1[3]
  PIN cpu_dtr_n1[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 814.290 1096.000 814.570 1100.000 ;
    END
  END cpu_dtr_n1[4]
  PIN cpu_dtr_n1[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 824.410 1096.000 824.690 1100.000 ;
    END
  END cpu_dtr_n1[5]
  PIN cpu_dtr_n1[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 834.990 1096.000 835.270 1100.000 ;
    END
  END cpu_dtr_n1[6]
  PIN cpu_dtr_n1[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 845.570 1096.000 845.850 1100.000 ;
    END
  END cpu_dtr_n1[7]
  PIN cpu_dtr_n1[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 855.690 1096.000 855.970 1100.000 ;
    END
  END cpu_dtr_n1[8]
  PIN cpu_dtr_n1[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 866.270 1096.000 866.550 1100.000 ;
    END
  END cpu_dtr_n1[9]
  PIN cpu_dtw_e[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 148.280 1100.000 148.880 ;
    END
  END cpu_dtw_e[0]
  PIN cpu_dtw_e[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 198.600 1100.000 199.200 ;
    END
  END cpu_dtw_e[10]
  PIN cpu_dtw_e[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 203.360 1100.000 203.960 ;
    END
  END cpu_dtw_e[11]
  PIN cpu_dtw_e[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 208.800 1100.000 209.400 ;
    END
  END cpu_dtw_e[12]
  PIN cpu_dtw_e[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 213.560 1100.000 214.160 ;
    END
  END cpu_dtw_e[13]
  PIN cpu_dtw_e[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 219.000 1100.000 219.600 ;
    END
  END cpu_dtw_e[14]
  PIN cpu_dtw_e[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 223.760 1100.000 224.360 ;
    END
  END cpu_dtw_e[15]
  PIN cpu_dtw_e[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 153.040 1100.000 153.640 ;
    END
  END cpu_dtw_e[1]
  PIN cpu_dtw_e[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 158.480 1100.000 159.080 ;
    END
  END cpu_dtw_e[2]
  PIN cpu_dtw_e[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 163.240 1100.000 163.840 ;
    END
  END cpu_dtw_e[3]
  PIN cpu_dtw_e[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 168.000 1100.000 168.600 ;
    END
  END cpu_dtw_e[4]
  PIN cpu_dtw_e[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 173.440 1100.000 174.040 ;
    END
  END cpu_dtw_e[5]
  PIN cpu_dtw_e[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 178.200 1100.000 178.800 ;
    END
  END cpu_dtw_e[6]
  PIN cpu_dtw_e[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 183.640 1100.000 184.240 ;
    END
  END cpu_dtw_e[7]
  PIN cpu_dtw_e[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 188.400 1100.000 189.000 ;
    END
  END cpu_dtw_e[8]
  PIN cpu_dtw_e[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 193.840 1100.000 194.440 ;
    END
  END cpu_dtw_e[9]
  PIN cpu_dtw_n[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 274.710 1096.000 274.990 1100.000 ;
    END
  END cpu_dtw_n[0]
  PIN cpu_dtw_n[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 378.670 1096.000 378.950 1100.000 ;
    END
  END cpu_dtw_n[10]
  PIN cpu_dtw_n[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 388.790 1096.000 389.070 1100.000 ;
    END
  END cpu_dtw_n[11]
  PIN cpu_dtw_n[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 399.370 1096.000 399.650 1100.000 ;
    END
  END cpu_dtw_n[12]
  PIN cpu_dtw_n[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 409.490 1096.000 409.770 1100.000 ;
    END
  END cpu_dtw_n[13]
  PIN cpu_dtw_n[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 420.070 1096.000 420.350 1100.000 ;
    END
  END cpu_dtw_n[14]
  PIN cpu_dtw_n[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 430.190 1096.000 430.470 1100.000 ;
    END
  END cpu_dtw_n[15]
  PIN cpu_dtw_n[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 285.290 1096.000 285.570 1100.000 ;
    END
  END cpu_dtw_n[1]
  PIN cpu_dtw_n[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 295.410 1096.000 295.690 1100.000 ;
    END
  END cpu_dtw_n[2]
  PIN cpu_dtw_n[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 305.990 1096.000 306.270 1100.000 ;
    END
  END cpu_dtw_n[3]
  PIN cpu_dtw_n[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 316.110 1096.000 316.390 1100.000 ;
    END
  END cpu_dtw_n[4]
  PIN cpu_dtw_n[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 326.690 1096.000 326.970 1100.000 ;
    END
  END cpu_dtw_n[5]
  PIN cpu_dtw_n[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 336.810 1096.000 337.090 1100.000 ;
    END
  END cpu_dtw_n[6]
  PIN cpu_dtw_n[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 347.390 1096.000 347.670 1100.000 ;
    END
  END cpu_dtw_n[7]
  PIN cpu_dtw_n[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 357.510 1096.000 357.790 1100.000 ;
    END
  END cpu_dtw_n[8]
  PIN cpu_dtw_n[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 368.090 1096.000 368.370 1100.000 ;
    END
  END cpu_dtw_n[9]
  PIN cpu_mask_e[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 17.040 1100.000 17.640 ;
    END
  END cpu_mask_e[0]
  PIN cpu_mask_e[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 21.800 1100.000 22.400 ;
    END
  END cpu_mask_e[1]
  PIN cpu_mask_e[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 27.240 1100.000 27.840 ;
    END
  END cpu_mask_e[2]
  PIN cpu_mask_e[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 32.000 1100.000 32.600 ;
    END
  END cpu_mask_e[3]
  PIN cpu_mask_e[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 36.760 1100.000 37.360 ;
    END
  END cpu_mask_e[4]
  PIN cpu_mask_e[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 42.200 1100.000 42.800 ;
    END
  END cpu_mask_e[5]
  PIN cpu_mask_e[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 46.960 1100.000 47.560 ;
    END
  END cpu_mask_e[6]
  PIN cpu_mask_e[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 52.400 1100.000 53.000 ;
    END
  END cpu_mask_e[7]
  PIN cpu_mask_n[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 5.150 1096.000 5.430 1100.000 ;
    END
  END cpu_mask_n[0]
  PIN cpu_mask_n[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 15.270 1096.000 15.550 1100.000 ;
    END
  END cpu_mask_n[1]
  PIN cpu_mask_n[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 25.850 1096.000 26.130 1100.000 ;
    END
  END cpu_mask_n[2]
  PIN cpu_mask_n[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 35.970 1096.000 36.250 1100.000 ;
    END
  END cpu_mask_n[3]
  PIN cpu_mask_n[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 46.550 1096.000 46.830 1100.000 ;
    END
  END cpu_mask_n[4]
  PIN cpu_mask_n[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 56.670 1096.000 56.950 1100.000 ;
    END
  END cpu_mask_n[5]
  PIN cpu_mask_n[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 67.250 1096.000 67.530 1100.000 ;
    END
  END cpu_mask_n[6]
  PIN cpu_mask_n[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 77.370 1096.000 77.650 1100.000 ;
    END
  END cpu_mask_n[7]
  PIN cpu_wen_e[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 57.160 1100.000 57.760 ;
    END
  END cpu_wen_e[0]
  PIN cpu_wen_e[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 62.600 1100.000 63.200 ;
    END
  END cpu_wen_e[1]
  PIN cpu_wen_n[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 87.950 1096.000 88.230 1100.000 ;
    END
  END cpu_wen_n[0]
  PIN cpu_wen_n[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 98.530 1096.000 98.810 1100.000 ;
    END
  END cpu_wen_n[1]
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.800 4.000 5.400 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 293.800 4.000 294.400 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.040 4.000 323.640 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 351.600 4.000 352.200 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 410.080 4.000 410.680 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 438.640 4.000 439.240 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 467.880 4.000 468.480 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 496.440 4.000 497.040 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 525.680 4.000 526.280 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 554.920 4.000 555.520 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 4.000 33.960 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 583.480 4.000 584.080 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 612.720 4.000 613.320 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 641.280 4.000 641.880 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 670.520 4.000 671.120 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 699.080 4.000 699.680 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 728.320 4.000 728.920 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 757.560 4.000 758.160 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 786.120 4.000 786.720 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 815.360 4.000 815.960 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 843.920 4.000 844.520 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 4.000 63.200 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 873.160 4.000 873.760 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 901.720 4.000 902.320 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 930.960 4.000 931.560 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 960.200 4.000 960.800 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 988.760 4.000 989.360 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1018.000 4.000 1018.600 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1046.560 4.000 1047.160 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1075.800 4.000 1076.400 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 4.000 91.760 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 120.400 4.000 121.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.960 4.000 149.560 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.200 4.000 178.800 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.440 4.000 208.040 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.000 4.000 236.600 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 14.320 4.000 14.920 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 303.320 4.000 303.920 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 332.560 4.000 333.160 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 361.800 4.000 362.400 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 390.360 4.000 390.960 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 419.600 4.000 420.200 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.160 4.000 448.760 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 477.400 4.000 478.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 506.640 4.000 507.240 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 535.200 4.000 535.800 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 564.440 4.000 565.040 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.880 4.000 43.480 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 593.000 4.000 593.600 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 622.240 4.000 622.840 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 650.800 4.000 651.400 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 680.040 4.000 680.640 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 709.280 4.000 709.880 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 737.840 4.000 738.440 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 767.080 4.000 767.680 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 795.640 4.000 796.240 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 824.880 4.000 825.480 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 853.440 4.000 854.040 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 4.000 72.720 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 882.680 4.000 883.280 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 911.920 4.000 912.520 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 940.480 4.000 941.080 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 969.720 4.000 970.320 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 998.280 4.000 998.880 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1027.520 4.000 1028.120 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1056.760 4.000 1057.360 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1085.320 4.000 1085.920 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 4.000 101.280 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.920 4.000 130.520 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.160 4.000 159.760 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.720 4.000 188.320 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.960 4.000 217.560 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 245.520 4.000 246.120 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.760 4.000 275.360 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 313.520 4.000 314.120 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 342.080 4.000 342.680 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 371.320 4.000 371.920 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 399.880 4.000 400.480 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 429.120 4.000 429.720 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 458.360 4.000 458.960 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.920 4.000 487.520 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 516.160 4.000 516.760 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 544.720 4.000 545.320 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 573.960 4.000 574.560 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 52.400 4.000 53.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 602.520 4.000 603.120 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 631.760 4.000 632.360 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 661.000 4.000 661.600 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 689.560 4.000 690.160 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 718.800 4.000 719.400 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 747.360 4.000 747.960 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 776.600 4.000 777.200 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 805.840 4.000 806.440 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 834.400 4.000 835.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 863.640 4.000 864.240 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 892.200 4.000 892.800 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 921.440 4.000 922.040 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 950.000 4.000 950.600 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 979.240 4.000 979.840 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1008.480 4.000 1009.080 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1037.040 4.000 1037.640 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1066.280 4.000 1066.880 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1094.840 4.000 1095.440 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.880 4.000 111.480 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.680 4.000 169.280 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 226.480 4.000 227.080 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.720 4.000 256.320 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.280 4.000 284.880 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1036.010 0.000 1036.290 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1065.450 0.000 1065.730 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1046.130 0.000 1046.410 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1075.110 0.000 1075.390 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1094.430 0.000 1094.710 4.000 ;
    END
  END la_data_out[2]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1055.790 0.000 1056.070 4.000 ;
    END
  END la_oen[0]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1084.770 0.000 1085.050 4.000 ;
    END
  END la_oen[1]
  PIN one
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 6.840 1100.000 7.440 ;
    END
  END one
  PIN ram_ce
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 11.600 1100.000 12.200 ;
    END
  END ram_ce
  PIN sr0_ce
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 552.200 1100.000 552.800 ;
    END
  END sr0_ce
  PIN sr0_dtr[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 556.960 1100.000 557.560 ;
    END
  END sr0_dtr[0]
  PIN sr0_dtr[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 607.280 1100.000 607.880 ;
    END
  END sr0_dtr[10]
  PIN sr0_dtr[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 612.720 1100.000 613.320 ;
    END
  END sr0_dtr[11]
  PIN sr0_dtr[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 617.480 1100.000 618.080 ;
    END
  END sr0_dtr[12]
  PIN sr0_dtr[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 622.240 1100.000 622.840 ;
    END
  END sr0_dtr[13]
  PIN sr0_dtr[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 627.680 1100.000 628.280 ;
    END
  END sr0_dtr[14]
  PIN sr0_dtr[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 632.440 1100.000 633.040 ;
    END
  END sr0_dtr[15]
  PIN sr0_dtr[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 637.880 1100.000 638.480 ;
    END
  END sr0_dtr[16]
  PIN sr0_dtr[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 642.640 1100.000 643.240 ;
    END
  END sr0_dtr[17]
  PIN sr0_dtr[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 648.080 1100.000 648.680 ;
    END
  END sr0_dtr[18]
  PIN sr0_dtr[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 652.840 1100.000 653.440 ;
    END
  END sr0_dtr[19]
  PIN sr0_dtr[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 561.720 1100.000 562.320 ;
    END
  END sr0_dtr[1]
  PIN sr0_dtr[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 657.600 1100.000 658.200 ;
    END
  END sr0_dtr[20]
  PIN sr0_dtr[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 663.040 1100.000 663.640 ;
    END
  END sr0_dtr[21]
  PIN sr0_dtr[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 667.800 1100.000 668.400 ;
    END
  END sr0_dtr[22]
  PIN sr0_dtr[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 673.240 1100.000 673.840 ;
    END
  END sr0_dtr[23]
  PIN sr0_dtr[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 678.000 1100.000 678.600 ;
    END
  END sr0_dtr[24]
  PIN sr0_dtr[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 682.760 1100.000 683.360 ;
    END
  END sr0_dtr[25]
  PIN sr0_dtr[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 688.200 1100.000 688.800 ;
    END
  END sr0_dtr[26]
  PIN sr0_dtr[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 692.960 1100.000 693.560 ;
    END
  END sr0_dtr[27]
  PIN sr0_dtr[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 698.400 1100.000 699.000 ;
    END
  END sr0_dtr[28]
  PIN sr0_dtr[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 703.160 1100.000 703.760 ;
    END
  END sr0_dtr[29]
  PIN sr0_dtr[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 567.160 1100.000 567.760 ;
    END
  END sr0_dtr[2]
  PIN sr0_dtr[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 708.600 1100.000 709.200 ;
    END
  END sr0_dtr[30]
  PIN sr0_dtr[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 713.360 1100.000 713.960 ;
    END
  END sr0_dtr[31]
  PIN sr0_dtr[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 571.920 1100.000 572.520 ;
    END
  END sr0_dtr[3]
  PIN sr0_dtr[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 577.360 1100.000 577.960 ;
    END
  END sr0_dtr[4]
  PIN sr0_dtr[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 582.120 1100.000 582.720 ;
    END
  END sr0_dtr[5]
  PIN sr0_dtr[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 586.880 1100.000 587.480 ;
    END
  END sr0_dtr[6]
  PIN sr0_dtr[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 592.320 1100.000 592.920 ;
    END
  END sr0_dtr[7]
  PIN sr0_dtr[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 597.080 1100.000 597.680 ;
    END
  END sr0_dtr[8]
  PIN sr0_dtr[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 602.520 1100.000 603.120 ;
    END
  END sr0_dtr[9]
  PIN sr1_ce
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 718.120 1100.000 718.720 ;
    END
  END sr1_ce
  PIN sr1_dtr[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 723.560 1100.000 724.160 ;
    END
  END sr1_dtr[0]
  PIN sr1_dtr[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 773.880 1100.000 774.480 ;
    END
  END sr1_dtr[10]
  PIN sr1_dtr[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 778.640 1100.000 779.240 ;
    END
  END sr1_dtr[11]
  PIN sr1_dtr[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 784.080 1100.000 784.680 ;
    END
  END sr1_dtr[12]
  PIN sr1_dtr[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 788.840 1100.000 789.440 ;
    END
  END sr1_dtr[13]
  PIN sr1_dtr[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 794.280 1100.000 794.880 ;
    END
  END sr1_dtr[14]
  PIN sr1_dtr[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 799.040 1100.000 799.640 ;
    END
  END sr1_dtr[15]
  PIN sr1_dtr[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 804.480 1100.000 805.080 ;
    END
  END sr1_dtr[16]
  PIN sr1_dtr[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 809.240 1100.000 809.840 ;
    END
  END sr1_dtr[17]
  PIN sr1_dtr[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 814.000 1100.000 814.600 ;
    END
  END sr1_dtr[18]
  PIN sr1_dtr[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 819.440 1100.000 820.040 ;
    END
  END sr1_dtr[19]
  PIN sr1_dtr[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 728.320 1100.000 728.920 ;
    END
  END sr1_dtr[1]
  PIN sr1_dtr[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 824.200 1100.000 824.800 ;
    END
  END sr1_dtr[20]
  PIN sr1_dtr[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 829.640 1100.000 830.240 ;
    END
  END sr1_dtr[21]
  PIN sr1_dtr[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 834.400 1100.000 835.000 ;
    END
  END sr1_dtr[22]
  PIN sr1_dtr[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 839.840 1100.000 840.440 ;
    END
  END sr1_dtr[23]
  PIN sr1_dtr[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 844.600 1100.000 845.200 ;
    END
  END sr1_dtr[24]
  PIN sr1_dtr[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 849.360 1100.000 849.960 ;
    END
  END sr1_dtr[25]
  PIN sr1_dtr[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 854.800 1100.000 855.400 ;
    END
  END sr1_dtr[26]
  PIN sr1_dtr[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 859.560 1100.000 860.160 ;
    END
  END sr1_dtr[27]
  PIN sr1_dtr[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 865.000 1100.000 865.600 ;
    END
  END sr1_dtr[28]
  PIN sr1_dtr[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 869.760 1100.000 870.360 ;
    END
  END sr1_dtr[29]
  PIN sr1_dtr[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 733.760 1100.000 734.360 ;
    END
  END sr1_dtr[2]
  PIN sr1_dtr[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 875.200 1100.000 875.800 ;
    END
  END sr1_dtr[30]
  PIN sr1_dtr[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 879.960 1100.000 880.560 ;
    END
  END sr1_dtr[31]
  PIN sr1_dtr[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 738.520 1100.000 739.120 ;
    END
  END sr1_dtr[3]
  PIN sr1_dtr[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 743.960 1100.000 744.560 ;
    END
  END sr1_dtr[4]
  PIN sr1_dtr[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 748.720 1100.000 749.320 ;
    END
  END sr1_dtr[5]
  PIN sr1_dtr[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 753.480 1100.000 754.080 ;
    END
  END sr1_dtr[6]
  PIN sr1_dtr[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 758.920 1100.000 759.520 ;
    END
  END sr1_dtr[7]
  PIN sr1_dtr[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 763.680 1100.000 764.280 ;
    END
  END sr1_dtr[8]
  PIN sr1_dtr[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1096.000 769.120 1100.000 769.720 ;
    END
  END sr1_dtr[9]
  PIN srx_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 890.160 1100.000 890.760 ;
    END
  END srx_addr[0]
  PIN srx_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 900.360 1100.000 900.960 ;
    END
  END srx_addr[1]
  PIN srx_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 909.880 1100.000 910.480 ;
    END
  END srx_addr[2]
  PIN srx_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 920.080 1100.000 920.680 ;
    END
  END srx_addr[3]
  PIN srx_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 930.280 1100.000 930.880 ;
    END
  END srx_addr[4]
  PIN srx_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 940.480 1100.000 941.080 ;
    END
  END srx_addr[5]
  PIN srx_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 950.680 1100.000 951.280 ;
    END
  END srx_addr[6]
  PIN srx_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 960.880 1100.000 961.480 ;
    END
  END srx_addr[7]
  PIN srx_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 971.080 1100.000 971.680 ;
    END
  END srx_addr[8]
  PIN srx_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 980.600 1100.000 981.200 ;
    END
  END srx_addr[9]
  PIN srx_dtw[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 894.920 1100.000 895.520 ;
    END
  END srx_dtw[0]
  PIN srx_dtw[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 990.800 1100.000 991.400 ;
    END
  END srx_dtw[10]
  PIN srx_dtw[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 996.240 1100.000 996.840 ;
    END
  END srx_dtw[11]
  PIN srx_dtw[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1001.000 1100.000 1001.600 ;
    END
  END srx_dtw[12]
  PIN srx_dtw[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1005.760 1100.000 1006.360 ;
    END
  END srx_dtw[13]
  PIN srx_dtw[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1011.200 1100.000 1011.800 ;
    END
  END srx_dtw[14]
  PIN srx_dtw[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1015.960 1100.000 1016.560 ;
    END
  END srx_dtw[15]
  PIN srx_dtw[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1021.400 1100.000 1022.000 ;
    END
  END srx_dtw[16]
  PIN srx_dtw[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1026.160 1100.000 1026.760 ;
    END
  END srx_dtw[17]
  PIN srx_dtw[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1031.600 1100.000 1032.200 ;
    END
  END srx_dtw[18]
  PIN srx_dtw[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1036.360 1100.000 1036.960 ;
    END
  END srx_dtw[19]
  PIN srx_dtw[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 905.120 1100.000 905.720 ;
    END
  END srx_dtw[1]
  PIN srx_dtw[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1041.120 1100.000 1041.720 ;
    END
  END srx_dtw[20]
  PIN srx_dtw[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1046.560 1100.000 1047.160 ;
    END
  END srx_dtw[21]
  PIN srx_dtw[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1051.320 1100.000 1051.920 ;
    END
  END srx_dtw[22]
  PIN srx_dtw[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1056.760 1100.000 1057.360 ;
    END
  END srx_dtw[23]
  PIN srx_dtw[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1061.520 1100.000 1062.120 ;
    END
  END srx_dtw[24]
  PIN srx_dtw[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1066.960 1100.000 1067.560 ;
    END
  END srx_dtw[25]
  PIN srx_dtw[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1071.720 1100.000 1072.320 ;
    END
  END srx_dtw[26]
  PIN srx_dtw[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1076.480 1100.000 1077.080 ;
    END
  END srx_dtw[27]
  PIN srx_dtw[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1081.920 1100.000 1082.520 ;
    END
  END srx_dtw[28]
  PIN srx_dtw[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1086.680 1100.000 1087.280 ;
    END
  END srx_dtw[29]
  PIN srx_dtw[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 915.320 1100.000 915.920 ;
    END
  END srx_dtw[2]
  PIN srx_dtw[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1092.120 1100.000 1092.720 ;
    END
  END srx_dtw[30]
  PIN srx_dtw[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 1096.880 1100.000 1097.480 ;
    END
  END srx_dtw[31]
  PIN srx_dtw[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 925.520 1100.000 926.120 ;
    END
  END srx_dtw[3]
  PIN srx_dtw[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 935.720 1100.000 936.320 ;
    END
  END srx_dtw[4]
  PIN srx_dtw[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 945.240 1100.000 945.840 ;
    END
  END srx_dtw[5]
  PIN srx_dtw[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 955.440 1100.000 956.040 ;
    END
  END srx_dtw[6]
  PIN srx_dtw[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 965.640 1100.000 966.240 ;
    END
  END srx_dtw[7]
  PIN srx_dtw[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 975.840 1100.000 976.440 ;
    END
  END srx_dtw[8]
  PIN srx_dtw[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 986.040 1100.000 986.640 ;
    END
  END srx_dtw[9]
  PIN srx_we
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 884.720 1100.000 885.320 ;
    END
  END srx_we
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4.690 0.000 4.970 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 14.350 0.000 14.630 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 24.010 0.000 24.290 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 393.850 0.000 394.130 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 422.830 0.000 423.110 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 452.270 0.000 452.550 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 481.250 0.000 481.530 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 510.690 0.000 510.970 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 539.670 0.000 539.950 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 569.110 0.000 569.390 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 598.090 0.000 598.370 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 627.530 0.000 627.810 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 656.510 0.000 656.790 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 101.750 0.000 102.030 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 685.950 0.000 686.230 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 714.930 0.000 715.210 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 744.370 0.000 744.650 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 773.350 0.000 773.630 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 802.790 0.000 803.070 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 831.770 0.000 832.050 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 861.210 0.000 861.490 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 890.190 0.000 890.470 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 919.170 0.000 919.450 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 948.610 0.000 948.890 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 140.850 0.000 141.130 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 977.590 0.000 977.870 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1007.030 0.000 1007.310 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 179.490 0.000 179.770 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 218.590 0.000 218.870 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 247.570 0.000 247.850 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 277.010 0.000 277.290 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 305.990 0.000 306.270 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 335.430 0.000 335.710 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 364.410 0.000 364.690 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 33.670 0.000 33.950 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 72.770 0.000 73.050 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 403.510 0.000 403.790 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 432.950 0.000 433.230 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 461.930 0.000 462.210 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 490.910 0.000 491.190 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 520.350 0.000 520.630 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 549.330 0.000 549.610 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 578.770 0.000 579.050 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 607.750 0.000 608.030 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 637.190 0.000 637.470 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 666.170 0.000 666.450 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 111.410 0.000 111.690 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 695.610 0.000 695.890 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 724.590 0.000 724.870 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 754.030 0.000 754.310 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 783.010 0.000 783.290 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 812.450 0.000 812.730 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 841.430 0.000 841.710 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 870.870 0.000 871.150 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 899.850 0.000 900.130 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 929.290 0.000 929.570 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 958.270 0.000 958.550 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 150.510 0.000 150.790 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 987.710 0.000 987.990 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1016.690 0.000 1016.970 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 189.610 0.000 189.890 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 228.250 0.000 228.530 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 316.110 0.000 316.390 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 345.090 0.000 345.370 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 374.530 0.000 374.810 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 82.430 0.000 82.710 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 413.170 0.000 413.450 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 442.610 0.000 442.890 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 471.590 0.000 471.870 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 501.030 0.000 501.310 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 530.010 0.000 530.290 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 559.450 0.000 559.730 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 588.430 0.000 588.710 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 617.870 0.000 618.150 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 646.850 0.000 647.130 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 675.830 0.000 676.110 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 121.070 0.000 121.350 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 705.270 0.000 705.550 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 734.250 0.000 734.530 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 763.690 0.000 763.970 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 792.670 0.000 792.950 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 822.110 0.000 822.390 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 851.090 0.000 851.370 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 880.530 0.000 880.810 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 909.510 0.000 909.790 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 938.950 0.000 939.230 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 967.930 0.000 968.210 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 160.170 0.000 160.450 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 997.370 0.000 997.650 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1026.350 0.000 1026.630 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 199.270 0.000 199.550 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 237.910 0.000 238.190 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 267.350 0.000 267.630 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 296.330 0.000 296.610 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 325.770 0.000 326.050 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 354.750 0.000 355.030 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 384.190 0.000 384.470 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 92.090 0.000 92.370 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 131.190 0.000 131.470 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 169.830 0.000 170.110 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 208.930 0.000 209.210 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 43.330 0.000 43.610 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.990 0.000 53.270 4.000 ;
    END
  END wbs_we_i
  PIN zero
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1096.000 2.080 1100.000 2.680 ;
    END
  END zero
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1088.240 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1088.240 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1095.115 1088.085 ;
      LAYER met1 ;
        RECT 0.070 4.460 1095.190 1095.780 ;
      LAYER met2 ;
        RECT 0.090 1095.720 4.870 1096.000 ;
        RECT 5.710 1095.720 14.990 1096.000 ;
        RECT 15.830 1095.720 25.570 1096.000 ;
        RECT 26.410 1095.720 35.690 1096.000 ;
        RECT 36.530 1095.720 46.270 1096.000 ;
        RECT 47.110 1095.720 56.390 1096.000 ;
        RECT 57.230 1095.720 66.970 1096.000 ;
        RECT 67.810 1095.720 77.090 1096.000 ;
        RECT 77.930 1095.720 87.670 1096.000 ;
        RECT 88.510 1095.720 98.250 1096.000 ;
        RECT 99.090 1095.720 108.370 1096.000 ;
        RECT 109.210 1095.720 118.950 1096.000 ;
        RECT 119.790 1095.720 129.070 1096.000 ;
        RECT 129.910 1095.720 139.650 1096.000 ;
        RECT 140.490 1095.720 149.770 1096.000 ;
        RECT 150.610 1095.720 160.350 1096.000 ;
        RECT 161.190 1095.720 170.470 1096.000 ;
        RECT 171.310 1095.720 181.050 1096.000 ;
        RECT 181.890 1095.720 191.630 1096.000 ;
        RECT 192.470 1095.720 201.750 1096.000 ;
        RECT 202.590 1095.720 212.330 1096.000 ;
        RECT 213.170 1095.720 222.450 1096.000 ;
        RECT 223.290 1095.720 233.030 1096.000 ;
        RECT 233.870 1095.720 243.150 1096.000 ;
        RECT 243.990 1095.720 253.730 1096.000 ;
        RECT 254.570 1095.720 263.850 1096.000 ;
        RECT 264.690 1095.720 274.430 1096.000 ;
        RECT 275.270 1095.720 285.010 1096.000 ;
        RECT 285.850 1095.720 295.130 1096.000 ;
        RECT 295.970 1095.720 305.710 1096.000 ;
        RECT 306.550 1095.720 315.830 1096.000 ;
        RECT 316.670 1095.720 326.410 1096.000 ;
        RECT 327.250 1095.720 336.530 1096.000 ;
        RECT 337.370 1095.720 347.110 1096.000 ;
        RECT 347.950 1095.720 357.230 1096.000 ;
        RECT 358.070 1095.720 367.810 1096.000 ;
        RECT 368.650 1095.720 378.390 1096.000 ;
        RECT 379.230 1095.720 388.510 1096.000 ;
        RECT 389.350 1095.720 399.090 1096.000 ;
        RECT 399.930 1095.720 409.210 1096.000 ;
        RECT 410.050 1095.720 419.790 1096.000 ;
        RECT 420.630 1095.720 429.910 1096.000 ;
        RECT 430.750 1095.720 440.490 1096.000 ;
        RECT 441.330 1095.720 450.610 1096.000 ;
        RECT 451.450 1095.720 461.190 1096.000 ;
        RECT 462.030 1095.720 471.770 1096.000 ;
        RECT 472.610 1095.720 481.890 1096.000 ;
        RECT 482.730 1095.720 492.470 1096.000 ;
        RECT 493.310 1095.720 502.590 1096.000 ;
        RECT 503.430 1095.720 513.170 1096.000 ;
        RECT 514.010 1095.720 523.290 1096.000 ;
        RECT 524.130 1095.720 533.870 1096.000 ;
        RECT 534.710 1095.720 543.990 1096.000 ;
        RECT 544.830 1095.720 554.570 1096.000 ;
        RECT 555.410 1095.720 565.150 1096.000 ;
        RECT 565.990 1095.720 575.270 1096.000 ;
        RECT 576.110 1095.720 585.850 1096.000 ;
        RECT 586.690 1095.720 595.970 1096.000 ;
        RECT 596.810 1095.720 606.550 1096.000 ;
        RECT 607.390 1095.720 616.670 1096.000 ;
        RECT 617.510 1095.720 627.250 1096.000 ;
        RECT 628.090 1095.720 637.370 1096.000 ;
        RECT 638.210 1095.720 647.950 1096.000 ;
        RECT 648.790 1095.720 658.530 1096.000 ;
        RECT 659.370 1095.720 668.650 1096.000 ;
        RECT 669.490 1095.720 679.230 1096.000 ;
        RECT 680.070 1095.720 689.350 1096.000 ;
        RECT 690.190 1095.720 699.930 1096.000 ;
        RECT 700.770 1095.720 710.050 1096.000 ;
        RECT 710.890 1095.720 720.630 1096.000 ;
        RECT 721.470 1095.720 730.750 1096.000 ;
        RECT 731.590 1095.720 741.330 1096.000 ;
        RECT 742.170 1095.720 751.910 1096.000 ;
        RECT 752.750 1095.720 762.030 1096.000 ;
        RECT 762.870 1095.720 772.610 1096.000 ;
        RECT 773.450 1095.720 782.730 1096.000 ;
        RECT 783.570 1095.720 793.310 1096.000 ;
        RECT 794.150 1095.720 803.430 1096.000 ;
        RECT 804.270 1095.720 814.010 1096.000 ;
        RECT 814.850 1095.720 824.130 1096.000 ;
        RECT 824.970 1095.720 834.710 1096.000 ;
        RECT 835.550 1095.720 845.290 1096.000 ;
        RECT 846.130 1095.720 855.410 1096.000 ;
        RECT 856.250 1095.720 865.990 1096.000 ;
        RECT 866.830 1095.720 876.110 1096.000 ;
        RECT 876.950 1095.720 886.690 1096.000 ;
        RECT 887.530 1095.720 896.810 1096.000 ;
        RECT 897.650 1095.720 907.390 1096.000 ;
        RECT 908.230 1095.720 917.510 1096.000 ;
        RECT 918.350 1095.720 928.090 1096.000 ;
        RECT 928.930 1095.720 938.670 1096.000 ;
        RECT 939.510 1095.720 948.790 1096.000 ;
        RECT 949.630 1095.720 959.370 1096.000 ;
        RECT 960.210 1095.720 969.490 1096.000 ;
        RECT 970.330 1095.720 980.070 1096.000 ;
        RECT 980.910 1095.720 990.190 1096.000 ;
        RECT 991.030 1095.720 1000.770 1096.000 ;
        RECT 1001.610 1095.720 1010.890 1096.000 ;
        RECT 1011.730 1095.720 1021.470 1096.000 ;
        RECT 1022.310 1095.720 1032.050 1096.000 ;
        RECT 1032.890 1095.720 1042.170 1096.000 ;
        RECT 1043.010 1095.720 1052.750 1096.000 ;
        RECT 1053.590 1095.720 1062.870 1096.000 ;
        RECT 1063.710 1095.720 1073.450 1096.000 ;
        RECT 1074.290 1095.720 1083.570 1096.000 ;
        RECT 1084.410 1095.720 1094.150 1096.000 ;
        RECT 1094.990 1095.720 1095.630 1096.000 ;
        RECT 0.090 4.280 1095.630 1095.720 ;
        RECT 0.090 2.195 4.410 4.280 ;
        RECT 5.250 2.195 14.070 4.280 ;
        RECT 14.910 2.195 23.730 4.280 ;
        RECT 24.570 2.195 33.390 4.280 ;
        RECT 34.230 2.195 43.050 4.280 ;
        RECT 43.890 2.195 52.710 4.280 ;
        RECT 53.550 2.195 62.370 4.280 ;
        RECT 63.210 2.195 72.490 4.280 ;
        RECT 73.330 2.195 82.150 4.280 ;
        RECT 82.990 2.195 91.810 4.280 ;
        RECT 92.650 2.195 101.470 4.280 ;
        RECT 102.310 2.195 111.130 4.280 ;
        RECT 111.970 2.195 120.790 4.280 ;
        RECT 121.630 2.195 130.910 4.280 ;
        RECT 131.750 2.195 140.570 4.280 ;
        RECT 141.410 2.195 150.230 4.280 ;
        RECT 151.070 2.195 159.890 4.280 ;
        RECT 160.730 2.195 169.550 4.280 ;
        RECT 170.390 2.195 179.210 4.280 ;
        RECT 180.050 2.195 189.330 4.280 ;
        RECT 190.170 2.195 198.990 4.280 ;
        RECT 199.830 2.195 208.650 4.280 ;
        RECT 209.490 2.195 218.310 4.280 ;
        RECT 219.150 2.195 227.970 4.280 ;
        RECT 228.810 2.195 237.630 4.280 ;
        RECT 238.470 2.195 247.290 4.280 ;
        RECT 248.130 2.195 257.410 4.280 ;
        RECT 258.250 2.195 267.070 4.280 ;
        RECT 267.910 2.195 276.730 4.280 ;
        RECT 277.570 2.195 286.390 4.280 ;
        RECT 287.230 2.195 296.050 4.280 ;
        RECT 296.890 2.195 305.710 4.280 ;
        RECT 306.550 2.195 315.830 4.280 ;
        RECT 316.670 2.195 325.490 4.280 ;
        RECT 326.330 2.195 335.150 4.280 ;
        RECT 335.990 2.195 344.810 4.280 ;
        RECT 345.650 2.195 354.470 4.280 ;
        RECT 355.310 2.195 364.130 4.280 ;
        RECT 364.970 2.195 374.250 4.280 ;
        RECT 375.090 2.195 383.910 4.280 ;
        RECT 384.750 2.195 393.570 4.280 ;
        RECT 394.410 2.195 403.230 4.280 ;
        RECT 404.070 2.195 412.890 4.280 ;
        RECT 413.730 2.195 422.550 4.280 ;
        RECT 423.390 2.195 432.670 4.280 ;
        RECT 433.510 2.195 442.330 4.280 ;
        RECT 443.170 2.195 451.990 4.280 ;
        RECT 452.830 2.195 461.650 4.280 ;
        RECT 462.490 2.195 471.310 4.280 ;
        RECT 472.150 2.195 480.970 4.280 ;
        RECT 481.810 2.195 490.630 4.280 ;
        RECT 491.470 2.195 500.750 4.280 ;
        RECT 501.590 2.195 510.410 4.280 ;
        RECT 511.250 2.195 520.070 4.280 ;
        RECT 520.910 2.195 529.730 4.280 ;
        RECT 530.570 2.195 539.390 4.280 ;
        RECT 540.230 2.195 549.050 4.280 ;
        RECT 549.890 2.195 559.170 4.280 ;
        RECT 560.010 2.195 568.830 4.280 ;
        RECT 569.670 2.195 578.490 4.280 ;
        RECT 579.330 2.195 588.150 4.280 ;
        RECT 588.990 2.195 597.810 4.280 ;
        RECT 598.650 2.195 607.470 4.280 ;
        RECT 608.310 2.195 617.590 4.280 ;
        RECT 618.430 2.195 627.250 4.280 ;
        RECT 628.090 2.195 636.910 4.280 ;
        RECT 637.750 2.195 646.570 4.280 ;
        RECT 647.410 2.195 656.230 4.280 ;
        RECT 657.070 2.195 665.890 4.280 ;
        RECT 666.730 2.195 675.550 4.280 ;
        RECT 676.390 2.195 685.670 4.280 ;
        RECT 686.510 2.195 695.330 4.280 ;
        RECT 696.170 2.195 704.990 4.280 ;
        RECT 705.830 2.195 714.650 4.280 ;
        RECT 715.490 2.195 724.310 4.280 ;
        RECT 725.150 2.195 733.970 4.280 ;
        RECT 734.810 2.195 744.090 4.280 ;
        RECT 744.930 2.195 753.750 4.280 ;
        RECT 754.590 2.195 763.410 4.280 ;
        RECT 764.250 2.195 773.070 4.280 ;
        RECT 773.910 2.195 782.730 4.280 ;
        RECT 783.570 2.195 792.390 4.280 ;
        RECT 793.230 2.195 802.510 4.280 ;
        RECT 803.350 2.195 812.170 4.280 ;
        RECT 813.010 2.195 821.830 4.280 ;
        RECT 822.670 2.195 831.490 4.280 ;
        RECT 832.330 2.195 841.150 4.280 ;
        RECT 841.990 2.195 850.810 4.280 ;
        RECT 851.650 2.195 860.930 4.280 ;
        RECT 861.770 2.195 870.590 4.280 ;
        RECT 871.430 2.195 880.250 4.280 ;
        RECT 881.090 2.195 889.910 4.280 ;
        RECT 890.750 2.195 899.570 4.280 ;
        RECT 900.410 2.195 909.230 4.280 ;
        RECT 910.070 2.195 918.890 4.280 ;
        RECT 919.730 2.195 929.010 4.280 ;
        RECT 929.850 2.195 938.670 4.280 ;
        RECT 939.510 2.195 948.330 4.280 ;
        RECT 949.170 2.195 957.990 4.280 ;
        RECT 958.830 2.195 967.650 4.280 ;
        RECT 968.490 2.195 977.310 4.280 ;
        RECT 978.150 2.195 987.430 4.280 ;
        RECT 988.270 2.195 997.090 4.280 ;
        RECT 997.930 2.195 1006.750 4.280 ;
        RECT 1007.590 2.195 1016.410 4.280 ;
        RECT 1017.250 2.195 1026.070 4.280 ;
        RECT 1026.910 2.195 1035.730 4.280 ;
        RECT 1036.570 2.195 1045.850 4.280 ;
        RECT 1046.690 2.195 1055.510 4.280 ;
        RECT 1056.350 2.195 1065.170 4.280 ;
        RECT 1066.010 2.195 1074.830 4.280 ;
        RECT 1075.670 2.195 1084.490 4.280 ;
        RECT 1085.330 2.195 1094.150 4.280 ;
        RECT 1094.990 2.195 1095.630 4.280 ;
      LAYER met3 ;
        RECT 0.065 1096.480 1095.600 1097.340 ;
        RECT 0.065 1095.840 1096.000 1096.480 ;
        RECT 4.400 1094.440 1096.000 1095.840 ;
        RECT 0.065 1093.120 1096.000 1094.440 ;
        RECT 0.065 1091.720 1095.600 1093.120 ;
        RECT 0.065 1087.680 1096.000 1091.720 ;
        RECT 0.065 1086.320 1095.600 1087.680 ;
        RECT 4.400 1086.280 1095.600 1086.320 ;
        RECT 4.400 1084.920 1096.000 1086.280 ;
        RECT 0.065 1082.920 1096.000 1084.920 ;
        RECT 0.065 1081.520 1095.600 1082.920 ;
        RECT 0.065 1077.480 1096.000 1081.520 ;
        RECT 0.065 1076.800 1095.600 1077.480 ;
        RECT 4.400 1076.080 1095.600 1076.800 ;
        RECT 4.400 1075.400 1096.000 1076.080 ;
        RECT 0.065 1072.720 1096.000 1075.400 ;
        RECT 0.065 1071.320 1095.600 1072.720 ;
        RECT 0.065 1067.960 1096.000 1071.320 ;
        RECT 0.065 1067.280 1095.600 1067.960 ;
        RECT 4.400 1066.560 1095.600 1067.280 ;
        RECT 4.400 1065.880 1096.000 1066.560 ;
        RECT 0.065 1062.520 1096.000 1065.880 ;
        RECT 0.065 1061.120 1095.600 1062.520 ;
        RECT 0.065 1057.760 1096.000 1061.120 ;
        RECT 4.400 1056.360 1095.600 1057.760 ;
        RECT 0.065 1052.320 1096.000 1056.360 ;
        RECT 0.065 1050.920 1095.600 1052.320 ;
        RECT 0.065 1047.560 1096.000 1050.920 ;
        RECT 4.400 1046.160 1095.600 1047.560 ;
        RECT 0.065 1042.120 1096.000 1046.160 ;
        RECT 0.065 1040.720 1095.600 1042.120 ;
        RECT 0.065 1038.040 1096.000 1040.720 ;
        RECT 4.400 1037.360 1096.000 1038.040 ;
        RECT 4.400 1036.640 1095.600 1037.360 ;
        RECT 0.065 1035.960 1095.600 1036.640 ;
        RECT 0.065 1032.600 1096.000 1035.960 ;
        RECT 0.065 1031.200 1095.600 1032.600 ;
        RECT 0.065 1028.520 1096.000 1031.200 ;
        RECT 4.400 1027.160 1096.000 1028.520 ;
        RECT 4.400 1027.120 1095.600 1027.160 ;
        RECT 0.065 1025.760 1095.600 1027.120 ;
        RECT 0.065 1022.400 1096.000 1025.760 ;
        RECT 0.065 1021.000 1095.600 1022.400 ;
        RECT 0.065 1019.000 1096.000 1021.000 ;
        RECT 4.400 1017.600 1096.000 1019.000 ;
        RECT 0.065 1016.960 1096.000 1017.600 ;
        RECT 0.065 1015.560 1095.600 1016.960 ;
        RECT 0.065 1012.200 1096.000 1015.560 ;
        RECT 0.065 1010.800 1095.600 1012.200 ;
        RECT 0.065 1009.480 1096.000 1010.800 ;
        RECT 4.400 1008.080 1096.000 1009.480 ;
        RECT 0.065 1006.760 1096.000 1008.080 ;
        RECT 0.065 1005.360 1095.600 1006.760 ;
        RECT 0.065 1002.000 1096.000 1005.360 ;
        RECT 0.065 1000.600 1095.600 1002.000 ;
        RECT 0.065 999.280 1096.000 1000.600 ;
        RECT 4.400 997.880 1096.000 999.280 ;
        RECT 0.065 997.240 1096.000 997.880 ;
        RECT 0.065 995.840 1095.600 997.240 ;
        RECT 0.065 991.800 1096.000 995.840 ;
        RECT 0.065 990.400 1095.600 991.800 ;
        RECT 0.065 989.760 1096.000 990.400 ;
        RECT 4.400 988.360 1096.000 989.760 ;
        RECT 0.065 987.040 1096.000 988.360 ;
        RECT 0.065 985.640 1095.600 987.040 ;
        RECT 0.065 981.600 1096.000 985.640 ;
        RECT 0.065 980.240 1095.600 981.600 ;
        RECT 4.400 980.200 1095.600 980.240 ;
        RECT 4.400 978.840 1096.000 980.200 ;
        RECT 0.065 976.840 1096.000 978.840 ;
        RECT 0.065 975.440 1095.600 976.840 ;
        RECT 0.065 972.080 1096.000 975.440 ;
        RECT 0.065 970.720 1095.600 972.080 ;
        RECT 4.400 970.680 1095.600 970.720 ;
        RECT 4.400 969.320 1096.000 970.680 ;
        RECT 0.065 966.640 1096.000 969.320 ;
        RECT 0.065 965.240 1095.600 966.640 ;
        RECT 0.065 961.880 1096.000 965.240 ;
        RECT 0.065 961.200 1095.600 961.880 ;
        RECT 4.400 960.480 1095.600 961.200 ;
        RECT 4.400 959.800 1096.000 960.480 ;
        RECT 0.065 956.440 1096.000 959.800 ;
        RECT 0.065 955.040 1095.600 956.440 ;
        RECT 0.065 951.680 1096.000 955.040 ;
        RECT 0.065 951.000 1095.600 951.680 ;
        RECT 4.400 950.280 1095.600 951.000 ;
        RECT 4.400 949.600 1096.000 950.280 ;
        RECT 0.065 946.240 1096.000 949.600 ;
        RECT 0.065 944.840 1095.600 946.240 ;
        RECT 0.065 941.480 1096.000 944.840 ;
        RECT 4.400 940.080 1095.600 941.480 ;
        RECT 0.065 936.720 1096.000 940.080 ;
        RECT 0.065 935.320 1095.600 936.720 ;
        RECT 0.065 931.960 1096.000 935.320 ;
        RECT 4.400 931.280 1096.000 931.960 ;
        RECT 4.400 930.560 1095.600 931.280 ;
        RECT 0.065 929.880 1095.600 930.560 ;
        RECT 0.065 926.520 1096.000 929.880 ;
        RECT 0.065 925.120 1095.600 926.520 ;
        RECT 0.065 922.440 1096.000 925.120 ;
        RECT 4.400 921.080 1096.000 922.440 ;
        RECT 4.400 921.040 1095.600 921.080 ;
        RECT 0.065 919.680 1095.600 921.040 ;
        RECT 0.065 916.320 1096.000 919.680 ;
        RECT 0.065 914.920 1095.600 916.320 ;
        RECT 0.065 912.920 1096.000 914.920 ;
        RECT 4.400 911.520 1096.000 912.920 ;
        RECT 0.065 910.880 1096.000 911.520 ;
        RECT 0.065 909.480 1095.600 910.880 ;
        RECT 0.065 906.120 1096.000 909.480 ;
        RECT 0.065 904.720 1095.600 906.120 ;
        RECT 0.065 902.720 1096.000 904.720 ;
        RECT 4.400 901.360 1096.000 902.720 ;
        RECT 4.400 901.320 1095.600 901.360 ;
        RECT 0.065 899.960 1095.600 901.320 ;
        RECT 0.065 895.920 1096.000 899.960 ;
        RECT 0.065 894.520 1095.600 895.920 ;
        RECT 0.065 893.200 1096.000 894.520 ;
        RECT 4.400 891.800 1096.000 893.200 ;
        RECT 0.065 891.160 1096.000 891.800 ;
        RECT 0.065 889.760 1095.600 891.160 ;
        RECT 0.065 885.720 1096.000 889.760 ;
        RECT 0.065 884.320 1095.600 885.720 ;
        RECT 0.065 883.680 1096.000 884.320 ;
        RECT 4.400 882.280 1096.000 883.680 ;
        RECT 0.065 880.960 1096.000 882.280 ;
        RECT 0.065 879.560 1095.600 880.960 ;
        RECT 0.065 876.200 1096.000 879.560 ;
        RECT 0.065 874.800 1095.600 876.200 ;
        RECT 0.065 874.160 1096.000 874.800 ;
        RECT 4.400 872.760 1096.000 874.160 ;
        RECT 0.065 870.760 1096.000 872.760 ;
        RECT 0.065 869.360 1095.600 870.760 ;
        RECT 0.065 866.000 1096.000 869.360 ;
        RECT 0.065 864.640 1095.600 866.000 ;
        RECT 4.400 864.600 1095.600 864.640 ;
        RECT 4.400 863.240 1096.000 864.600 ;
        RECT 0.065 860.560 1096.000 863.240 ;
        RECT 0.065 859.160 1095.600 860.560 ;
        RECT 0.065 855.800 1096.000 859.160 ;
        RECT 0.065 854.440 1095.600 855.800 ;
        RECT 4.400 854.400 1095.600 854.440 ;
        RECT 4.400 853.040 1096.000 854.400 ;
        RECT 0.065 850.360 1096.000 853.040 ;
        RECT 0.065 848.960 1095.600 850.360 ;
        RECT 0.065 845.600 1096.000 848.960 ;
        RECT 0.065 844.920 1095.600 845.600 ;
        RECT 4.400 844.200 1095.600 844.920 ;
        RECT 4.400 843.520 1096.000 844.200 ;
        RECT 0.065 840.840 1096.000 843.520 ;
        RECT 0.065 839.440 1095.600 840.840 ;
        RECT 0.065 835.400 1096.000 839.440 ;
        RECT 4.400 834.000 1095.600 835.400 ;
        RECT 0.065 830.640 1096.000 834.000 ;
        RECT 0.065 829.240 1095.600 830.640 ;
        RECT 0.065 825.880 1096.000 829.240 ;
        RECT 4.400 825.200 1096.000 825.880 ;
        RECT 4.400 824.480 1095.600 825.200 ;
        RECT 0.065 823.800 1095.600 824.480 ;
        RECT 0.065 820.440 1096.000 823.800 ;
        RECT 0.065 819.040 1095.600 820.440 ;
        RECT 0.065 816.360 1096.000 819.040 ;
        RECT 4.400 815.000 1096.000 816.360 ;
        RECT 4.400 814.960 1095.600 815.000 ;
        RECT 0.065 813.600 1095.600 814.960 ;
        RECT 0.065 810.240 1096.000 813.600 ;
        RECT 0.065 808.840 1095.600 810.240 ;
        RECT 0.065 806.840 1096.000 808.840 ;
        RECT 4.400 805.480 1096.000 806.840 ;
        RECT 4.400 805.440 1095.600 805.480 ;
        RECT 0.065 804.080 1095.600 805.440 ;
        RECT 0.065 800.040 1096.000 804.080 ;
        RECT 0.065 798.640 1095.600 800.040 ;
        RECT 0.065 796.640 1096.000 798.640 ;
        RECT 4.400 795.280 1096.000 796.640 ;
        RECT 4.400 795.240 1095.600 795.280 ;
        RECT 0.065 793.880 1095.600 795.240 ;
        RECT 0.065 789.840 1096.000 793.880 ;
        RECT 0.065 788.440 1095.600 789.840 ;
        RECT 0.065 787.120 1096.000 788.440 ;
        RECT 4.400 785.720 1096.000 787.120 ;
        RECT 0.065 785.080 1096.000 785.720 ;
        RECT 0.065 783.680 1095.600 785.080 ;
        RECT 0.065 779.640 1096.000 783.680 ;
        RECT 0.065 778.240 1095.600 779.640 ;
        RECT 0.065 777.600 1096.000 778.240 ;
        RECT 4.400 776.200 1096.000 777.600 ;
        RECT 0.065 774.880 1096.000 776.200 ;
        RECT 0.065 773.480 1095.600 774.880 ;
        RECT 0.065 770.120 1096.000 773.480 ;
        RECT 0.065 768.720 1095.600 770.120 ;
        RECT 0.065 768.080 1096.000 768.720 ;
        RECT 4.400 766.680 1096.000 768.080 ;
        RECT 0.065 764.680 1096.000 766.680 ;
        RECT 0.065 763.280 1095.600 764.680 ;
        RECT 0.065 759.920 1096.000 763.280 ;
        RECT 0.065 758.560 1095.600 759.920 ;
        RECT 4.400 758.520 1095.600 758.560 ;
        RECT 4.400 757.160 1096.000 758.520 ;
        RECT 0.065 754.480 1096.000 757.160 ;
        RECT 0.065 753.080 1095.600 754.480 ;
        RECT 0.065 749.720 1096.000 753.080 ;
        RECT 0.065 748.360 1095.600 749.720 ;
        RECT 4.400 748.320 1095.600 748.360 ;
        RECT 4.400 746.960 1096.000 748.320 ;
        RECT 0.065 744.960 1096.000 746.960 ;
        RECT 0.065 743.560 1095.600 744.960 ;
        RECT 0.065 739.520 1096.000 743.560 ;
        RECT 0.065 738.840 1095.600 739.520 ;
        RECT 4.400 738.120 1095.600 738.840 ;
        RECT 4.400 737.440 1096.000 738.120 ;
        RECT 0.065 734.760 1096.000 737.440 ;
        RECT 0.065 733.360 1095.600 734.760 ;
        RECT 0.065 729.320 1096.000 733.360 ;
        RECT 4.400 727.920 1095.600 729.320 ;
        RECT 0.065 724.560 1096.000 727.920 ;
        RECT 0.065 723.160 1095.600 724.560 ;
        RECT 0.065 719.800 1096.000 723.160 ;
        RECT 4.400 719.120 1096.000 719.800 ;
        RECT 4.400 718.400 1095.600 719.120 ;
        RECT 0.065 717.720 1095.600 718.400 ;
        RECT 0.065 714.360 1096.000 717.720 ;
        RECT 0.065 712.960 1095.600 714.360 ;
        RECT 0.065 710.280 1096.000 712.960 ;
        RECT 4.400 709.600 1096.000 710.280 ;
        RECT 4.400 708.880 1095.600 709.600 ;
        RECT 0.065 708.200 1095.600 708.880 ;
        RECT 0.065 704.160 1096.000 708.200 ;
        RECT 0.065 702.760 1095.600 704.160 ;
        RECT 0.065 700.080 1096.000 702.760 ;
        RECT 4.400 699.400 1096.000 700.080 ;
        RECT 4.400 698.680 1095.600 699.400 ;
        RECT 0.065 698.000 1095.600 698.680 ;
        RECT 0.065 693.960 1096.000 698.000 ;
        RECT 0.065 692.560 1095.600 693.960 ;
        RECT 0.065 690.560 1096.000 692.560 ;
        RECT 4.400 689.200 1096.000 690.560 ;
        RECT 4.400 689.160 1095.600 689.200 ;
        RECT 0.065 687.800 1095.600 689.160 ;
        RECT 0.065 683.760 1096.000 687.800 ;
        RECT 0.065 682.360 1095.600 683.760 ;
        RECT 0.065 681.040 1096.000 682.360 ;
        RECT 4.400 679.640 1096.000 681.040 ;
        RECT 0.065 679.000 1096.000 679.640 ;
        RECT 0.065 677.600 1095.600 679.000 ;
        RECT 0.065 674.240 1096.000 677.600 ;
        RECT 0.065 672.840 1095.600 674.240 ;
        RECT 0.065 671.520 1096.000 672.840 ;
        RECT 4.400 670.120 1096.000 671.520 ;
        RECT 0.065 668.800 1096.000 670.120 ;
        RECT 0.065 667.400 1095.600 668.800 ;
        RECT 0.065 664.040 1096.000 667.400 ;
        RECT 0.065 662.640 1095.600 664.040 ;
        RECT 0.065 662.000 1096.000 662.640 ;
        RECT 4.400 660.600 1096.000 662.000 ;
        RECT 0.065 658.600 1096.000 660.600 ;
        RECT 0.065 657.200 1095.600 658.600 ;
        RECT 0.065 653.840 1096.000 657.200 ;
        RECT 0.065 652.440 1095.600 653.840 ;
        RECT 0.065 651.800 1096.000 652.440 ;
        RECT 4.400 650.400 1096.000 651.800 ;
        RECT 0.065 649.080 1096.000 650.400 ;
        RECT 0.065 647.680 1095.600 649.080 ;
        RECT 0.065 643.640 1096.000 647.680 ;
        RECT 0.065 642.280 1095.600 643.640 ;
        RECT 4.400 642.240 1095.600 642.280 ;
        RECT 4.400 640.880 1096.000 642.240 ;
        RECT 0.065 638.880 1096.000 640.880 ;
        RECT 0.065 637.480 1095.600 638.880 ;
        RECT 0.065 633.440 1096.000 637.480 ;
        RECT 0.065 632.760 1095.600 633.440 ;
        RECT 4.400 632.040 1095.600 632.760 ;
        RECT 4.400 631.360 1096.000 632.040 ;
        RECT 0.065 628.680 1096.000 631.360 ;
        RECT 0.065 627.280 1095.600 628.680 ;
        RECT 0.065 623.240 1096.000 627.280 ;
        RECT 4.400 621.840 1095.600 623.240 ;
        RECT 0.065 618.480 1096.000 621.840 ;
        RECT 0.065 617.080 1095.600 618.480 ;
        RECT 0.065 613.720 1096.000 617.080 ;
        RECT 4.400 612.320 1095.600 613.720 ;
        RECT 0.065 608.280 1096.000 612.320 ;
        RECT 0.065 606.880 1095.600 608.280 ;
        RECT 0.065 603.520 1096.000 606.880 ;
        RECT 4.400 602.120 1095.600 603.520 ;
        RECT 0.065 598.080 1096.000 602.120 ;
        RECT 0.065 596.680 1095.600 598.080 ;
        RECT 0.065 594.000 1096.000 596.680 ;
        RECT 4.400 593.320 1096.000 594.000 ;
        RECT 4.400 592.600 1095.600 593.320 ;
        RECT 0.065 591.920 1095.600 592.600 ;
        RECT 0.065 587.880 1096.000 591.920 ;
        RECT 0.065 586.480 1095.600 587.880 ;
        RECT 0.065 584.480 1096.000 586.480 ;
        RECT 4.400 583.120 1096.000 584.480 ;
        RECT 4.400 583.080 1095.600 583.120 ;
        RECT 0.065 581.720 1095.600 583.080 ;
        RECT 0.065 578.360 1096.000 581.720 ;
        RECT 0.065 576.960 1095.600 578.360 ;
        RECT 0.065 574.960 1096.000 576.960 ;
        RECT 4.400 573.560 1096.000 574.960 ;
        RECT 0.065 572.920 1096.000 573.560 ;
        RECT 0.065 571.520 1095.600 572.920 ;
        RECT 0.065 568.160 1096.000 571.520 ;
        RECT 0.065 566.760 1095.600 568.160 ;
        RECT 0.065 565.440 1096.000 566.760 ;
        RECT 4.400 564.040 1096.000 565.440 ;
        RECT 0.065 562.720 1096.000 564.040 ;
        RECT 0.065 561.320 1095.600 562.720 ;
        RECT 0.065 557.960 1096.000 561.320 ;
        RECT 0.065 556.560 1095.600 557.960 ;
        RECT 0.065 555.920 1096.000 556.560 ;
        RECT 4.400 554.520 1096.000 555.920 ;
        RECT 0.065 553.200 1096.000 554.520 ;
        RECT 0.065 551.800 1095.600 553.200 ;
        RECT 0.065 547.760 1096.000 551.800 ;
        RECT 0.065 546.360 1095.600 547.760 ;
        RECT 0.065 545.720 1096.000 546.360 ;
        RECT 4.400 544.320 1096.000 545.720 ;
        RECT 0.065 543.000 1096.000 544.320 ;
        RECT 0.065 541.600 1095.600 543.000 ;
        RECT 0.065 537.560 1096.000 541.600 ;
        RECT 0.065 536.200 1095.600 537.560 ;
        RECT 4.400 536.160 1095.600 536.200 ;
        RECT 4.400 534.800 1096.000 536.160 ;
        RECT 0.065 532.800 1096.000 534.800 ;
        RECT 0.065 531.400 1095.600 532.800 ;
        RECT 0.065 527.360 1096.000 531.400 ;
        RECT 0.065 526.680 1095.600 527.360 ;
        RECT 4.400 525.960 1095.600 526.680 ;
        RECT 4.400 525.280 1096.000 525.960 ;
        RECT 0.065 522.600 1096.000 525.280 ;
        RECT 0.065 521.200 1095.600 522.600 ;
        RECT 0.065 517.840 1096.000 521.200 ;
        RECT 0.065 517.160 1095.600 517.840 ;
        RECT 4.400 516.440 1095.600 517.160 ;
        RECT 4.400 515.760 1096.000 516.440 ;
        RECT 0.065 512.400 1096.000 515.760 ;
        RECT 0.065 511.000 1095.600 512.400 ;
        RECT 0.065 507.640 1096.000 511.000 ;
        RECT 4.400 506.240 1095.600 507.640 ;
        RECT 0.065 502.200 1096.000 506.240 ;
        RECT 0.065 500.800 1095.600 502.200 ;
        RECT 0.065 497.440 1096.000 500.800 ;
        RECT 4.400 496.040 1095.600 497.440 ;
        RECT 0.065 492.000 1096.000 496.040 ;
        RECT 0.065 490.600 1095.600 492.000 ;
        RECT 0.065 487.920 1096.000 490.600 ;
        RECT 4.400 487.240 1096.000 487.920 ;
        RECT 4.400 486.520 1095.600 487.240 ;
        RECT 0.065 485.840 1095.600 486.520 ;
        RECT 0.065 482.480 1096.000 485.840 ;
        RECT 0.065 481.080 1095.600 482.480 ;
        RECT 0.065 478.400 1096.000 481.080 ;
        RECT 4.400 477.040 1096.000 478.400 ;
        RECT 4.400 477.000 1095.600 477.040 ;
        RECT 0.065 475.640 1095.600 477.000 ;
        RECT 0.065 472.280 1096.000 475.640 ;
        RECT 0.065 470.880 1095.600 472.280 ;
        RECT 0.065 468.880 1096.000 470.880 ;
        RECT 4.400 467.480 1096.000 468.880 ;
        RECT 0.065 466.840 1096.000 467.480 ;
        RECT 0.065 465.440 1095.600 466.840 ;
        RECT 0.065 462.080 1096.000 465.440 ;
        RECT 0.065 460.680 1095.600 462.080 ;
        RECT 0.065 459.360 1096.000 460.680 ;
        RECT 4.400 457.960 1096.000 459.360 ;
        RECT 0.065 456.640 1096.000 457.960 ;
        RECT 0.065 455.240 1095.600 456.640 ;
        RECT 0.065 451.880 1096.000 455.240 ;
        RECT 0.065 450.480 1095.600 451.880 ;
        RECT 0.065 449.160 1096.000 450.480 ;
        RECT 4.400 447.760 1096.000 449.160 ;
        RECT 0.065 447.120 1096.000 447.760 ;
        RECT 0.065 445.720 1095.600 447.120 ;
        RECT 0.065 441.680 1096.000 445.720 ;
        RECT 0.065 440.280 1095.600 441.680 ;
        RECT 0.065 439.640 1096.000 440.280 ;
        RECT 4.400 438.240 1096.000 439.640 ;
        RECT 0.065 436.920 1096.000 438.240 ;
        RECT 0.065 435.520 1095.600 436.920 ;
        RECT 0.065 431.480 1096.000 435.520 ;
        RECT 0.065 430.120 1095.600 431.480 ;
        RECT 4.400 430.080 1095.600 430.120 ;
        RECT 4.400 428.720 1096.000 430.080 ;
        RECT 0.065 426.720 1096.000 428.720 ;
        RECT 0.065 425.320 1095.600 426.720 ;
        RECT 0.065 421.960 1096.000 425.320 ;
        RECT 0.065 420.600 1095.600 421.960 ;
        RECT 4.400 420.560 1095.600 420.600 ;
        RECT 4.400 419.200 1096.000 420.560 ;
        RECT 0.065 416.520 1096.000 419.200 ;
        RECT 0.065 415.120 1095.600 416.520 ;
        RECT 0.065 411.760 1096.000 415.120 ;
        RECT 0.065 411.080 1095.600 411.760 ;
        RECT 4.400 410.360 1095.600 411.080 ;
        RECT 4.400 409.680 1096.000 410.360 ;
        RECT 0.065 406.320 1096.000 409.680 ;
        RECT 0.065 404.920 1095.600 406.320 ;
        RECT 0.065 401.560 1096.000 404.920 ;
        RECT 0.065 400.880 1095.600 401.560 ;
        RECT 4.400 400.160 1095.600 400.880 ;
        RECT 4.400 399.480 1096.000 400.160 ;
        RECT 0.065 396.120 1096.000 399.480 ;
        RECT 0.065 394.720 1095.600 396.120 ;
        RECT 0.065 391.360 1096.000 394.720 ;
        RECT 4.400 389.960 1095.600 391.360 ;
        RECT 0.065 386.600 1096.000 389.960 ;
        RECT 0.065 385.200 1095.600 386.600 ;
        RECT 0.065 381.840 1096.000 385.200 ;
        RECT 4.400 381.160 1096.000 381.840 ;
        RECT 4.400 380.440 1095.600 381.160 ;
        RECT 0.065 379.760 1095.600 380.440 ;
        RECT 0.065 376.400 1096.000 379.760 ;
        RECT 0.065 375.000 1095.600 376.400 ;
        RECT 0.065 372.320 1096.000 375.000 ;
        RECT 4.400 370.960 1096.000 372.320 ;
        RECT 4.400 370.920 1095.600 370.960 ;
        RECT 0.065 369.560 1095.600 370.920 ;
        RECT 0.065 366.200 1096.000 369.560 ;
        RECT 0.065 364.800 1095.600 366.200 ;
        RECT 0.065 362.800 1096.000 364.800 ;
        RECT 4.400 361.400 1096.000 362.800 ;
        RECT 0.065 360.760 1096.000 361.400 ;
        RECT 0.065 359.360 1095.600 360.760 ;
        RECT 0.065 356.000 1096.000 359.360 ;
        RECT 0.065 354.600 1095.600 356.000 ;
        RECT 0.065 352.600 1096.000 354.600 ;
        RECT 4.400 351.240 1096.000 352.600 ;
        RECT 4.400 351.200 1095.600 351.240 ;
        RECT 0.065 349.840 1095.600 351.200 ;
        RECT 0.065 345.800 1096.000 349.840 ;
        RECT 0.065 344.400 1095.600 345.800 ;
        RECT 0.065 343.080 1096.000 344.400 ;
        RECT 4.400 341.680 1096.000 343.080 ;
        RECT 0.065 341.040 1096.000 341.680 ;
        RECT 0.065 339.640 1095.600 341.040 ;
        RECT 0.065 335.600 1096.000 339.640 ;
        RECT 0.065 334.200 1095.600 335.600 ;
        RECT 0.065 333.560 1096.000 334.200 ;
        RECT 4.400 332.160 1096.000 333.560 ;
        RECT 0.065 330.840 1096.000 332.160 ;
        RECT 0.065 329.440 1095.600 330.840 ;
        RECT 0.065 326.080 1096.000 329.440 ;
        RECT 0.065 324.680 1095.600 326.080 ;
        RECT 0.065 324.040 1096.000 324.680 ;
        RECT 4.400 322.640 1096.000 324.040 ;
        RECT 0.065 320.640 1096.000 322.640 ;
        RECT 0.065 319.240 1095.600 320.640 ;
        RECT 0.065 315.880 1096.000 319.240 ;
        RECT 0.065 314.520 1095.600 315.880 ;
        RECT 4.400 314.480 1095.600 314.520 ;
        RECT 4.400 313.120 1096.000 314.480 ;
        RECT 0.065 310.440 1096.000 313.120 ;
        RECT 0.065 309.040 1095.600 310.440 ;
        RECT 0.065 305.680 1096.000 309.040 ;
        RECT 0.065 304.320 1095.600 305.680 ;
        RECT 4.400 304.280 1095.600 304.320 ;
        RECT 4.400 302.920 1096.000 304.280 ;
        RECT 0.065 300.240 1096.000 302.920 ;
        RECT 0.065 298.840 1095.600 300.240 ;
        RECT 0.065 295.480 1096.000 298.840 ;
        RECT 0.065 294.800 1095.600 295.480 ;
        RECT 4.400 294.080 1095.600 294.800 ;
        RECT 4.400 293.400 1096.000 294.080 ;
        RECT 0.065 290.720 1096.000 293.400 ;
        RECT 0.065 289.320 1095.600 290.720 ;
        RECT 0.065 285.280 1096.000 289.320 ;
        RECT 4.400 283.880 1095.600 285.280 ;
        RECT 0.065 280.520 1096.000 283.880 ;
        RECT 0.065 279.120 1095.600 280.520 ;
        RECT 0.065 275.760 1096.000 279.120 ;
        RECT 4.400 275.080 1096.000 275.760 ;
        RECT 4.400 274.360 1095.600 275.080 ;
        RECT 0.065 273.680 1095.600 274.360 ;
        RECT 0.065 270.320 1096.000 273.680 ;
        RECT 0.065 268.920 1095.600 270.320 ;
        RECT 0.065 266.240 1096.000 268.920 ;
        RECT 4.400 264.880 1096.000 266.240 ;
        RECT 4.400 264.840 1095.600 264.880 ;
        RECT 0.065 263.480 1095.600 264.840 ;
        RECT 0.065 260.120 1096.000 263.480 ;
        RECT 0.065 258.720 1095.600 260.120 ;
        RECT 0.065 256.720 1096.000 258.720 ;
        RECT 4.400 255.360 1096.000 256.720 ;
        RECT 4.400 255.320 1095.600 255.360 ;
        RECT 0.065 253.960 1095.600 255.320 ;
        RECT 0.065 249.920 1096.000 253.960 ;
        RECT 0.065 248.520 1095.600 249.920 ;
        RECT 0.065 246.520 1096.000 248.520 ;
        RECT 4.400 245.160 1096.000 246.520 ;
        RECT 4.400 245.120 1095.600 245.160 ;
        RECT 0.065 243.760 1095.600 245.120 ;
        RECT 0.065 239.720 1096.000 243.760 ;
        RECT 0.065 238.320 1095.600 239.720 ;
        RECT 0.065 237.000 1096.000 238.320 ;
        RECT 4.400 235.600 1096.000 237.000 ;
        RECT 0.065 234.960 1096.000 235.600 ;
        RECT 0.065 233.560 1095.600 234.960 ;
        RECT 0.065 229.520 1096.000 233.560 ;
        RECT 0.065 228.120 1095.600 229.520 ;
        RECT 0.065 227.480 1096.000 228.120 ;
        RECT 4.400 226.080 1096.000 227.480 ;
        RECT 0.065 224.760 1096.000 226.080 ;
        RECT 0.065 223.360 1095.600 224.760 ;
        RECT 0.065 220.000 1096.000 223.360 ;
        RECT 0.065 218.600 1095.600 220.000 ;
        RECT 0.065 217.960 1096.000 218.600 ;
        RECT 4.400 216.560 1096.000 217.960 ;
        RECT 0.065 214.560 1096.000 216.560 ;
        RECT 0.065 213.160 1095.600 214.560 ;
        RECT 0.065 209.800 1096.000 213.160 ;
        RECT 0.065 208.440 1095.600 209.800 ;
        RECT 4.400 208.400 1095.600 208.440 ;
        RECT 4.400 207.040 1096.000 208.400 ;
        RECT 0.065 204.360 1096.000 207.040 ;
        RECT 0.065 202.960 1095.600 204.360 ;
        RECT 0.065 199.600 1096.000 202.960 ;
        RECT 0.065 198.240 1095.600 199.600 ;
        RECT 4.400 198.200 1095.600 198.240 ;
        RECT 4.400 196.840 1096.000 198.200 ;
        RECT 0.065 194.840 1096.000 196.840 ;
        RECT 0.065 193.440 1095.600 194.840 ;
        RECT 0.065 189.400 1096.000 193.440 ;
        RECT 0.065 188.720 1095.600 189.400 ;
        RECT 4.400 188.000 1095.600 188.720 ;
        RECT 4.400 187.320 1096.000 188.000 ;
        RECT 0.065 184.640 1096.000 187.320 ;
        RECT 0.065 183.240 1095.600 184.640 ;
        RECT 0.065 179.200 1096.000 183.240 ;
        RECT 4.400 177.800 1095.600 179.200 ;
        RECT 0.065 174.440 1096.000 177.800 ;
        RECT 0.065 173.040 1095.600 174.440 ;
        RECT 0.065 169.680 1096.000 173.040 ;
        RECT 4.400 169.000 1096.000 169.680 ;
        RECT 4.400 168.280 1095.600 169.000 ;
        RECT 0.065 167.600 1095.600 168.280 ;
        RECT 0.065 164.240 1096.000 167.600 ;
        RECT 0.065 162.840 1095.600 164.240 ;
        RECT 0.065 160.160 1096.000 162.840 ;
        RECT 4.400 159.480 1096.000 160.160 ;
        RECT 4.400 158.760 1095.600 159.480 ;
        RECT 0.065 158.080 1095.600 158.760 ;
        RECT 0.065 154.040 1096.000 158.080 ;
        RECT 0.065 152.640 1095.600 154.040 ;
        RECT 0.065 149.960 1096.000 152.640 ;
        RECT 4.400 149.280 1096.000 149.960 ;
        RECT 4.400 148.560 1095.600 149.280 ;
        RECT 0.065 147.880 1095.600 148.560 ;
        RECT 0.065 143.840 1096.000 147.880 ;
        RECT 0.065 142.440 1095.600 143.840 ;
        RECT 0.065 140.440 1096.000 142.440 ;
        RECT 4.400 139.080 1096.000 140.440 ;
        RECT 4.400 139.040 1095.600 139.080 ;
        RECT 0.065 137.680 1095.600 139.040 ;
        RECT 0.065 133.640 1096.000 137.680 ;
        RECT 0.065 132.240 1095.600 133.640 ;
        RECT 0.065 130.920 1096.000 132.240 ;
        RECT 4.400 129.520 1096.000 130.920 ;
        RECT 0.065 128.880 1096.000 129.520 ;
        RECT 0.065 127.480 1095.600 128.880 ;
        RECT 0.065 124.120 1096.000 127.480 ;
        RECT 0.065 122.720 1095.600 124.120 ;
        RECT 0.065 121.400 1096.000 122.720 ;
        RECT 4.400 120.000 1096.000 121.400 ;
        RECT 0.065 118.680 1096.000 120.000 ;
        RECT 0.065 117.280 1095.600 118.680 ;
        RECT 0.065 113.920 1096.000 117.280 ;
        RECT 0.065 112.520 1095.600 113.920 ;
        RECT 0.065 111.880 1096.000 112.520 ;
        RECT 4.400 110.480 1096.000 111.880 ;
        RECT 0.065 108.480 1096.000 110.480 ;
        RECT 0.065 107.080 1095.600 108.480 ;
        RECT 0.065 103.720 1096.000 107.080 ;
        RECT 0.065 102.320 1095.600 103.720 ;
        RECT 0.065 101.680 1096.000 102.320 ;
        RECT 4.400 100.280 1096.000 101.680 ;
        RECT 0.065 98.960 1096.000 100.280 ;
        RECT 0.065 97.560 1095.600 98.960 ;
        RECT 0.065 93.520 1096.000 97.560 ;
        RECT 0.065 92.160 1095.600 93.520 ;
        RECT 4.400 92.120 1095.600 92.160 ;
        RECT 4.400 90.760 1096.000 92.120 ;
        RECT 0.065 88.760 1096.000 90.760 ;
        RECT 0.065 87.360 1095.600 88.760 ;
        RECT 0.065 83.320 1096.000 87.360 ;
        RECT 0.065 82.640 1095.600 83.320 ;
        RECT 4.400 81.920 1095.600 82.640 ;
        RECT 4.400 81.240 1096.000 81.920 ;
        RECT 0.065 78.560 1096.000 81.240 ;
        RECT 0.065 77.160 1095.600 78.560 ;
        RECT 0.065 73.120 1096.000 77.160 ;
        RECT 4.400 71.720 1095.600 73.120 ;
        RECT 0.065 68.360 1096.000 71.720 ;
        RECT 0.065 66.960 1095.600 68.360 ;
        RECT 0.065 63.600 1096.000 66.960 ;
        RECT 4.400 62.200 1095.600 63.600 ;
        RECT 0.065 58.160 1096.000 62.200 ;
        RECT 0.065 56.760 1095.600 58.160 ;
        RECT 0.065 53.400 1096.000 56.760 ;
        RECT 4.400 52.000 1095.600 53.400 ;
        RECT 0.065 47.960 1096.000 52.000 ;
        RECT 0.065 46.560 1095.600 47.960 ;
        RECT 0.065 43.880 1096.000 46.560 ;
        RECT 4.400 43.200 1096.000 43.880 ;
        RECT 4.400 42.480 1095.600 43.200 ;
        RECT 0.065 41.800 1095.600 42.480 ;
        RECT 0.065 37.760 1096.000 41.800 ;
        RECT 0.065 36.360 1095.600 37.760 ;
        RECT 0.065 34.360 1096.000 36.360 ;
        RECT 4.400 33.000 1096.000 34.360 ;
        RECT 4.400 32.960 1095.600 33.000 ;
        RECT 0.065 31.600 1095.600 32.960 ;
        RECT 0.065 28.240 1096.000 31.600 ;
        RECT 0.065 26.840 1095.600 28.240 ;
        RECT 0.065 24.840 1096.000 26.840 ;
        RECT 4.400 23.440 1096.000 24.840 ;
        RECT 0.065 22.800 1096.000 23.440 ;
        RECT 0.065 21.400 1095.600 22.800 ;
        RECT 0.065 18.040 1096.000 21.400 ;
        RECT 0.065 16.640 1095.600 18.040 ;
        RECT 0.065 15.320 1096.000 16.640 ;
        RECT 4.400 13.920 1096.000 15.320 ;
        RECT 0.065 12.600 1096.000 13.920 ;
        RECT 0.065 11.200 1095.600 12.600 ;
        RECT 0.065 7.840 1096.000 11.200 ;
        RECT 0.065 6.440 1095.600 7.840 ;
        RECT 0.065 5.800 1096.000 6.440 ;
        RECT 4.400 4.400 1096.000 5.800 ;
        RECT 0.065 3.080 1096.000 4.400 ;
        RECT 0.065 2.215 1095.600 3.080 ;
      LAYER met4 ;
        RECT 23.295 1088.640 1089.905 1097.345 ;
        RECT 23.295 10.240 97.440 1088.640 ;
        RECT 99.840 10.240 1089.905 1088.640 ;
        RECT 23.295 6.975 1089.905 10.240 ;
  END
END hs32_core1
END LIBRARY

